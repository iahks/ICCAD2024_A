 module top_809568696_809776567_809698999_863110837_1234615 (a, b, o);

      input a, b; output o; nor_6 g0(a,b,o); endmodule