 module top_810026173_843396535_809698999_829556405_809567927 (a, o);

      input a, b; output o; buf_5 g0(a,o); endmodule