// Benchmark "top_810222779_843330999_776144567_776418743_1234615" written by ABC on Mon Aug 12 17:39:42 2024

module top_810222779_843330999_776144567_776418743_1234615 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107;
  wire new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n551, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1068, new_n1069, new_n1070, new_n1071, new_n1073,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1126, new_n1127, new_n1128, new_n1130, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1311, new_n1312, new_n1313, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1320, new_n1321, new_n1324,
    new_n1326, new_n1328, new_n1329, new_n1332, new_n1333, new_n1334,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1356, new_n1357, new_n1358, new_n1359, new_n1360,
    new_n1361, new_n1362, new_n1363, new_n1364, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369, new_n1370, new_n1371, new_n1377,
    new_n1380, new_n1381, new_n1385;
  nand_5 g0000(.A(pi123), .B(pi000), .Y(new_n316));
  not_8  g0001(.A(pi150), .Y(new_n317));
  or_6   g0002(.A(new_n317), .B(pi026), .Y(new_n318));
  nand_5 g0003(.A(new_n318), .B(new_n316), .Y(new_n319));
  xor_4  g0004(.A(new_n319), .B(pi153), .Y(new_n320));
  not_8  g0005(.A(new_n320), .Y(new_n321));
  or_6   g0006(.A(new_n317), .B(pi054), .Y(new_n322));
  nand_5 g0007(.A(new_n322), .B(new_n316), .Y(new_n323));
  nand_5 g0008(.A(new_n323), .B(pi050), .Y(new_n324));
  xor_4  g0009(.A(new_n323), .B(pi050), .Y(new_n325));
  not_8  g0010(.A(new_n325), .Y(new_n326));
  or_6   g0011(.A(new_n317), .B(pi115), .Y(new_n327));
  nand_5 g0012(.A(new_n327), .B(new_n316), .Y(new_n328));
  or_6   g0013(.A(new_n328), .B(pi056), .Y(new_n329));
  xor_4  g0014(.A(new_n328), .B(pi056), .Y(new_n330));
  or_6   g0015(.A(pi154), .B(new_n317), .Y(new_n331));
  nand_5 g0016(.A(new_n331), .B(new_n316), .Y(new_n332));
  nor_5  g0017(.A(new_n332), .B(pi122), .Y(new_n333));
  not_8  g0018(.A(new_n333), .Y(new_n334));
  nand_5 g0019(.A(new_n332), .B(pi122), .Y(new_n335));
  not_8  g0020(.A(new_n335), .Y(new_n336));
  nor_5  g0021(.A(new_n336), .B(new_n333), .Y(new_n337));
  or_6   g0022(.A(pi175), .B(new_n317), .Y(new_n338));
  nand_5 g0023(.A(new_n338), .B(new_n316), .Y(new_n339));
  nand_5 g0024(.A(new_n339), .B(pi047), .Y(new_n340));
  not_8  g0025(.A(new_n340), .Y(new_n341));
  nor_5  g0026(.A(new_n339), .B(pi047), .Y(new_n342));
  or_6   g0027(.A(pi182), .B(new_n317), .Y(new_n343));
  or_6   g0028(.A(pi186), .B(pi150), .Y(new_n344));
  nand_5 g0029(.A(new_n344), .B(new_n343), .Y(new_n345));
  nand_5 g0030(.A(new_n345), .B(pi196), .Y(new_n346));
  or_6   g0031(.A(new_n345), .B(pi196), .Y(new_n347));
  or_6   g0032(.A(pi177), .B(pi150), .Y(new_n348));
  or_6   g0033(.A(new_n317), .B(pi009), .Y(new_n349));
  nand_5 g0034(.A(new_n349), .B(new_n348), .Y(new_n350));
  nand_5 g0035(.A(new_n350), .B(pi199), .Y(new_n351));
  or_6   g0036(.A(new_n350), .B(pi199), .Y(new_n352));
  or_6   g0037(.A(pi203), .B(pi150), .Y(new_n353));
  or_6   g0038(.A(new_n317), .B(pi080), .Y(new_n354));
  nand_5 g0039(.A(new_n354), .B(new_n353), .Y(new_n355));
  nand_5 g0040(.A(new_n355), .B(pi178), .Y(new_n356));
  or_6   g0041(.A(new_n355), .B(pi178), .Y(new_n357));
  or_6   g0042(.A(pi151), .B(pi150), .Y(new_n358));
  or_6   g0043(.A(pi172), .B(new_n317), .Y(new_n359));
  nand_5 g0044(.A(new_n359), .B(new_n358), .Y(new_n360));
  or_6   g0045(.A(new_n360), .B(pi162), .Y(new_n361));
  nand_5 g0046(.A(new_n361), .B(new_n357), .Y(new_n362));
  nand_5 g0047(.A(new_n362), .B(new_n356), .Y(new_n363));
  nand_5 g0048(.A(new_n363), .B(new_n352), .Y(new_n364));
  nand_5 g0049(.A(new_n364), .B(new_n351), .Y(new_n365));
  nand_5 g0050(.A(new_n365), .B(new_n347), .Y(new_n366));
  nand_5 g0051(.A(new_n366), .B(new_n346), .Y(new_n367));
  nand_5 g0052(.A(new_n357), .B(new_n356), .Y(new_n368));
  not_8  g0053(.A(new_n368), .Y(new_n369));
  nand_5 g0054(.A(new_n352), .B(new_n351), .Y(new_n370));
  not_8  g0055(.A(new_n370), .Y(new_n371));
  nand_5 g0056(.A(new_n371), .B(new_n369), .Y(new_n372));
  nand_5 g0057(.A(new_n360), .B(pi162), .Y(new_n373));
  nand_5 g0058(.A(new_n373), .B(new_n361), .Y(new_n374));
  nor_5  g0059(.A(new_n374), .B(new_n372), .Y(new_n375));
  nand_5 g0060(.A(new_n375), .B(new_n346), .Y(new_n376));
  or_6   g0061(.A(pi164), .B(new_n317), .Y(new_n377));
  or_6   g0062(.A(pi150), .B(pi034), .Y(new_n378));
  nand_5 g0063(.A(new_n378), .B(new_n377), .Y(new_n379));
  nor_5  g0064(.A(new_n379), .B(pi160), .Y(new_n380));
  not_8  g0065(.A(pi160), .Y(new_n381));
  xor_4  g0066(.A(new_n379), .B(new_n381), .Y(new_n382));
  or_6   g0067(.A(pi150), .B(pi139), .Y(new_n383));
  or_6   g0068(.A(new_n317), .B(pi090), .Y(new_n384));
  nand_5 g0069(.A(new_n384), .B(new_n383), .Y(new_n385));
  nand_5 g0070(.A(new_n385), .B(pi192), .Y(new_n386));
  or_6   g0071(.A(new_n385), .B(pi192), .Y(new_n387));
  or_6   g0072(.A(pi158), .B(new_n317), .Y(new_n388));
  or_6   g0073(.A(pi150), .B(pi146), .Y(new_n389));
  nand_5 g0074(.A(new_n389), .B(new_n388), .Y(new_n390));
  nand_5 g0075(.A(new_n390), .B(pi116), .Y(new_n391));
  not_8  g0076(.A(pi116), .Y(new_n392));
  not_8  g0077(.A(new_n390), .Y(new_n393));
  nand_5 g0078(.A(new_n393), .B(new_n392), .Y(new_n394));
  or_6   g0079(.A(pi150), .B(pi086), .Y(new_n395));
  or_6   g0080(.A(new_n317), .B(pi030), .Y(new_n396));
  nand_5 g0081(.A(new_n396), .B(new_n395), .Y(new_n397));
  nor_5  g0082(.A(new_n397), .B(pi039), .Y(new_n398));
  not_8  g0083(.A(new_n398), .Y(new_n399));
  nand_5 g0084(.A(new_n399), .B(new_n394), .Y(new_n400));
  nand_5 g0085(.A(new_n400), .B(new_n391), .Y(new_n401));
  nand_5 g0086(.A(new_n401), .B(new_n387), .Y(new_n402));
  not_8  g0087(.A(new_n402), .Y(new_n403));
  nand_5 g0088(.A(new_n397), .B(pi039), .Y(new_n404));
  nand_5 g0089(.A(new_n404), .B(new_n399), .Y(new_n405));
  nand_5 g0090(.A(new_n394), .B(new_n391), .Y(new_n406));
  nor_5  g0091(.A(new_n406), .B(new_n405), .Y(new_n407));
  not_8  g0092(.A(new_n407), .Y(new_n408));
  not_8  g0093(.A(pi057), .Y(new_n409));
  nand_5 g0094(.A(new_n317), .B(pi142), .Y(new_n410));
  nand_5 g0095(.A(pi150), .B(pi032), .Y(new_n411));
  nand_5 g0096(.A(new_n411), .B(new_n410), .Y(new_n412));
  or_6   g0097(.A(new_n412), .B(new_n409), .Y(new_n413));
  nand_5 g0098(.A(new_n412), .B(new_n409), .Y(new_n414));
  or_6   g0099(.A(pi187), .B(new_n317), .Y(new_n415));
  or_6   g0100(.A(pi150), .B(pi094), .Y(new_n416));
  nand_5 g0101(.A(new_n416), .B(new_n415), .Y(new_n417));
  nand_5 g0102(.A(new_n417), .B(pi183), .Y(new_n418));
  nor_5  g0103(.A(new_n417), .B(pi183), .Y(new_n419));
  or_6   g0104(.A(pi189), .B(pi150), .Y(new_n420));
  or_6   g0105(.A(new_n317), .B(pi106), .Y(new_n421));
  nand_5 g0106(.A(new_n421), .B(new_n420), .Y(new_n422));
  nand_5 g0107(.A(new_n422), .B(pi107), .Y(new_n423));
  or_6   g0108(.A(new_n422), .B(pi107), .Y(new_n424));
  or_6   g0109(.A(pi156), .B(pi150), .Y(new_n425));
  or_6   g0110(.A(pi194), .B(new_n317), .Y(new_n426));
  nand_5 g0111(.A(new_n426), .B(new_n425), .Y(new_n427));
  nand_5 g0112(.A(new_n427), .B(pi020), .Y(new_n428));
  or_6   g0113(.A(pi150), .B(pi131), .Y(new_n429));
  or_6   g0114(.A(new_n317), .B(pi012), .Y(new_n430));
  nand_5 g0115(.A(new_n430), .B(new_n429), .Y(new_n431));
  or_6   g0116(.A(new_n431), .B(pi170), .Y(new_n432));
  or_6   g0117(.A(new_n427), .B(pi020), .Y(new_n433));
  nand_5 g0118(.A(new_n433), .B(new_n432), .Y(new_n434));
  nand_5 g0119(.A(new_n434), .B(new_n428), .Y(new_n435));
  nand_5 g0120(.A(new_n435), .B(new_n424), .Y(new_n436));
  nand_5 g0121(.A(new_n436), .B(new_n423), .Y(new_n437));
  not_8  g0122(.A(new_n437), .Y(new_n438));
  nor_5  g0123(.A(new_n438), .B(new_n419), .Y(new_n439));
  nand_5 g0124(.A(new_n424), .B(new_n423), .Y(new_n440));
  not_8  g0125(.A(new_n440), .Y(new_n441));
  nand_5 g0126(.A(new_n433), .B(new_n428), .Y(new_n442));
  nand_5 g0127(.A(new_n431), .B(pi170), .Y(new_n443));
  nand_5 g0128(.A(new_n443), .B(new_n432), .Y(new_n444));
  not_8  g0129(.A(new_n444), .Y(new_n445));
  or_6   g0130(.A(new_n317), .B(pi087), .Y(new_n446));
  or_6   g0131(.A(pi150), .B(pi014), .Y(new_n447));
  nand_5 g0132(.A(new_n447), .B(new_n446), .Y(new_n448));
  nor_5  g0133(.A(new_n448), .B(pi051), .Y(new_n449));
  xnor_4 g0134(.A(new_n448), .B(pi051), .Y(new_n450));
  or_6   g0135(.A(pi150), .B(pi081), .Y(new_n451));
  or_6   g0136(.A(new_n317), .B(pi035), .Y(new_n452));
  nand_5 g0137(.A(new_n452), .B(new_n451), .Y(new_n453));
  nand_5 g0138(.A(new_n453), .B(pi074), .Y(new_n454));
  or_6   g0139(.A(new_n453), .B(pi074), .Y(new_n455));
  nand_5 g0140(.A(new_n455), .B(new_n454), .Y(new_n456));
  not_8  g0141(.A(new_n456), .Y(new_n457));
  or_6   g0142(.A(pi169), .B(new_n317), .Y(new_n458));
  or_6   g0143(.A(pi150), .B(pi033), .Y(new_n459));
  nand_5 g0144(.A(new_n459), .B(new_n458), .Y(new_n460));
  nand_5 g0145(.A(new_n460), .B(pi180), .Y(new_n461));
  not_8  g0146(.A(new_n461), .Y(new_n462));
  nor_5  g0147(.A(new_n460), .B(pi180), .Y(new_n463));
  or_6   g0148(.A(new_n317), .B(pi044), .Y(new_n464));
  or_6   g0149(.A(pi150), .B(pi042), .Y(new_n465));
  nand_5 g0150(.A(new_n465), .B(new_n464), .Y(new_n466));
  nand_5 g0151(.A(new_n466), .B(pi027), .Y(new_n467));
  nor_5  g0152(.A(new_n467), .B(new_n463), .Y(new_n468));
  nor_5  g0153(.A(new_n468), .B(new_n462), .Y(new_n469));
  nor_5  g0154(.A(new_n466), .B(pi027), .Y(new_n470));
  nor_5  g0155(.A(new_n470), .B(new_n463), .Y(new_n471));
  or_6   g0156(.A(pi197), .B(new_n317), .Y(new_n472));
  or_6   g0157(.A(pi150), .B(pi007), .Y(new_n473));
  nand_5 g0158(.A(new_n473), .B(new_n472), .Y(new_n474));
  nand_5 g0159(.A(new_n474), .B(pi083), .Y(new_n475));
  xor_4  g0160(.A(new_n474), .B(pi083), .Y(new_n476));
  not_8  g0161(.A(pi132), .Y(new_n477));
  or_6   g0162(.A(pi150), .B(pi143), .Y(new_n478));
  or_6   g0163(.A(new_n317), .B(pi043), .Y(new_n479));
  nand_5 g0164(.A(new_n479), .B(new_n478), .Y(new_n480));
  not_8  g0165(.A(new_n480), .Y(new_n481));
  nand_5 g0166(.A(new_n481), .B(new_n477), .Y(new_n482));
  not_8  g0167(.A(new_n482), .Y(new_n483));
  nand_5 g0168(.A(new_n480), .B(pi132), .Y(new_n484));
  nand_5 g0169(.A(new_n484), .B(new_n482), .Y(new_n485));
  or_6   g0170(.A(pi150), .B(pi058), .Y(new_n486));
  or_6   g0171(.A(new_n317), .B(pi025), .Y(new_n487));
  nand_5 g0172(.A(new_n487), .B(new_n486), .Y(new_n488));
  nand_5 g0173(.A(new_n488), .B(pi004), .Y(new_n489));
  nor_5  g0174(.A(new_n488), .B(pi004), .Y(new_n490));
  not_8  g0175(.A(new_n490), .Y(new_n491));
  nand_5 g0176(.A(new_n491), .B(new_n489), .Y(new_n492));
  not_8  g0177(.A(new_n492), .Y(new_n493));
  or_6   g0178(.A(pi152), .B(pi150), .Y(new_n494));
  or_6   g0179(.A(pi193), .B(new_n317), .Y(new_n495));
  nand_5 g0180(.A(new_n495), .B(new_n494), .Y(new_n496));
  nand_5 g0181(.A(new_n496), .B(pi092), .Y(new_n497));
  or_6   g0182(.A(new_n496), .B(pi092), .Y(new_n498));
  nand_5 g0183(.A(new_n498), .B(new_n497), .Y(new_n499));
  not_8  g0184(.A(pi147), .Y(new_n500));
  nand_5 g0185(.A(new_n500), .B(pi069), .Y(new_n501));
  nor_5  g0186(.A(new_n501), .B(pi150), .Y(new_n502));
  not_8  g0187(.A(new_n502), .Y(new_n503));
  nor_5  g0188(.A(pi150), .B(pi069), .Y(new_n504));
  nand_5 g0189(.A(new_n504), .B(pi147), .Y(new_n505));
  nand_5 g0190(.A(new_n505), .B(new_n503), .Y(new_n506));
  not_8  g0191(.A(new_n506), .Y(new_n507));
  nand_5 g0192(.A(new_n507), .B(pi070), .Y(new_n508));
  nand_5 g0193(.A(new_n508), .B(new_n503), .Y(new_n509));
  or_6   g0194(.A(new_n509), .B(new_n499), .Y(new_n510));
  nand_5 g0195(.A(new_n510), .B(new_n497), .Y(new_n511));
  nand_5 g0196(.A(new_n511), .B(new_n493), .Y(new_n512));
  nand_5 g0197(.A(new_n512), .B(new_n489), .Y(new_n513));
  nor_5  g0198(.A(new_n513), .B(new_n485), .Y(new_n514));
  nor_5  g0199(.A(new_n514), .B(new_n483), .Y(new_n515));
  nand_5 g0200(.A(new_n515), .B(new_n476), .Y(new_n516));
  nand_5 g0201(.A(new_n516), .B(new_n475), .Y(new_n517));
  nand_5 g0202(.A(new_n517), .B(new_n471), .Y(new_n518));
  nand_5 g0203(.A(new_n518), .B(new_n469), .Y(new_n519));
  nand_5 g0204(.A(new_n519), .B(new_n457), .Y(new_n520));
  nand_5 g0205(.A(new_n520), .B(new_n454), .Y(new_n521));
  nor_5  g0206(.A(new_n521), .B(new_n450), .Y(new_n522));
  nor_5  g0207(.A(new_n522), .B(new_n449), .Y(new_n523));
  not_8  g0208(.A(new_n523), .Y(new_n524));
  nand_5 g0209(.A(new_n524), .B(new_n445), .Y(new_n525));
  nor_5  g0210(.A(new_n525), .B(new_n442), .Y(new_n526));
  nand_5 g0211(.A(new_n526), .B(new_n441), .Y(new_n527));
  nand_5 g0212(.A(new_n527), .B(new_n439), .Y(new_n528));
  nand_5 g0213(.A(new_n528), .B(new_n418), .Y(new_n529));
  nand_5 g0214(.A(new_n529), .B(new_n414), .Y(new_n530));
  nand_5 g0215(.A(new_n530), .B(new_n413), .Y(new_n531));
  or_6   g0216(.A(new_n531), .B(new_n408), .Y(new_n532));
  nand_5 g0217(.A(new_n532), .B(new_n403), .Y(new_n533));
  nand_5 g0218(.A(new_n533), .B(new_n386), .Y(new_n534));
  nor_5  g0219(.A(new_n534), .B(new_n382), .Y(new_n535));
  nor_5  g0220(.A(new_n535), .B(new_n380), .Y(new_n536));
  or_6   g0221(.A(new_n536), .B(new_n376), .Y(new_n537));
  nand_5 g0222(.A(new_n537), .B(new_n367), .Y(new_n538));
  nor_5  g0223(.A(new_n538), .B(new_n342), .Y(new_n539));
  nor_5  g0224(.A(new_n539), .B(new_n341), .Y(new_n540));
  nand_5 g0225(.A(new_n540), .B(new_n337), .Y(new_n541));
  nand_5 g0226(.A(new_n541), .B(new_n334), .Y(new_n542));
  nand_5 g0227(.A(new_n542), .B(new_n330), .Y(new_n543));
  nand_5 g0228(.A(new_n543), .B(new_n329), .Y(new_n544));
  or_6   g0229(.A(new_n544), .B(new_n326), .Y(new_n545));
  nand_5 g0230(.A(new_n545), .B(new_n324), .Y(new_n546));
  xor_4  g0231(.A(new_n546), .B(new_n321), .Y(po000));
  not_8  g0232(.A(pi165), .Y(new_n548));
  nand_5 g0233(.A(pi167), .B(new_n548), .Y(po003));
  xor_4  g0234(.A(new_n531), .B(new_n405), .Y(po005));
  nand_5 g0235(.A(pi075), .B(pi037), .Y(new_n551));
  nand_5 g0236(.A(pi198), .B(pi188), .Y(new_n552));
  nor_5  g0237(.A(new_n552), .B(new_n551), .Y(new_n553));
  not_8  g0238(.A(new_n553), .Y(po006));
  or_6   g0239(.A(new_n317), .B(pi052), .Y(new_n555));
  nand_5 g0240(.A(new_n555), .B(new_n378), .Y(new_n556));
  not_8  g0241(.A(new_n556), .Y(new_n557));
  nand_5 g0242(.A(new_n381), .B(pi150), .Y(new_n558));
  nand_5 g0243(.A(new_n317), .B(pi104), .Y(new_n559));
  nand_5 g0244(.A(new_n559), .B(new_n558), .Y(new_n560));
  or_6   g0245(.A(new_n560), .B(new_n557), .Y(new_n561));
  nand_5 g0246(.A(new_n560), .B(new_n557), .Y(new_n562));
  or_6   g0247(.A(pi192), .B(new_n317), .Y(new_n563));
  nand_5 g0248(.A(new_n317), .B(pi068), .Y(new_n564));
  nand_5 g0249(.A(new_n564), .B(new_n563), .Y(new_n565));
  or_6   g0250(.A(new_n317), .B(pi036), .Y(new_n566));
  nand_5 g0251(.A(new_n566), .B(new_n383), .Y(new_n567));
  not_8  g0252(.A(new_n567), .Y(new_n568));
  or_6   g0253(.A(new_n317), .B(pi002), .Y(new_n569));
  nand_5 g0254(.A(new_n569), .B(new_n486), .Y(new_n570));
  nand_5 g0255(.A(pi150), .B(pi004), .Y(new_n571));
  not_8  g0256(.A(new_n571), .Y(new_n572));
  nor_5  g0257(.A(pi150), .B(pi111), .Y(new_n573));
  nor_5  g0258(.A(new_n573), .B(new_n572), .Y(new_n574));
  not_8  g0259(.A(new_n574), .Y(new_n575));
  or_6   g0260(.A(new_n575), .B(new_n570), .Y(new_n576));
  nand_5 g0261(.A(new_n317), .B(pi066), .Y(new_n577));
  or_6   g0262(.A(new_n317), .B(pi092), .Y(new_n578));
  nand_5 g0263(.A(new_n578), .B(new_n577), .Y(new_n579));
  or_6   g0264(.A(new_n317), .B(pi103), .Y(new_n580));
  nand_5 g0265(.A(new_n580), .B(new_n494), .Y(new_n581));
  nand_5 g0266(.A(new_n317), .B(pi096), .Y(new_n582));
  nor_5  g0267(.A(pi091), .B(pi069), .Y(new_n583));
  nor_5  g0268(.A(new_n583), .B(new_n582), .Y(new_n584));
  not_8  g0269(.A(new_n504), .Y(new_n585));
  nand_5 g0270(.A(new_n585), .B(pi091), .Y(new_n586));
  not_8  g0271(.A(new_n586), .Y(new_n587));
  nor_5  g0272(.A(new_n587), .B(new_n584), .Y(new_n588));
  nor_5  g0273(.A(new_n588), .B(new_n581), .Y(new_n589));
  or_6   g0274(.A(new_n589), .B(new_n579), .Y(new_n590));
  nand_5 g0275(.A(new_n588), .B(new_n581), .Y(new_n591));
  nand_5 g0276(.A(new_n591), .B(new_n590), .Y(new_n592));
  nand_5 g0277(.A(new_n592), .B(new_n576), .Y(new_n593));
  nand_5 g0278(.A(new_n575), .B(new_n570), .Y(new_n594));
  or_6   g0279(.A(new_n317), .B(pi089), .Y(new_n595));
  nand_5 g0280(.A(new_n595), .B(new_n478), .Y(new_n596));
  nand_5 g0281(.A(new_n317), .B(pi048), .Y(new_n597));
  nand_5 g0282(.A(pi150), .B(new_n477), .Y(new_n598));
  nand_5 g0283(.A(new_n598), .B(new_n597), .Y(new_n599));
  not_8  g0284(.A(new_n599), .Y(new_n600));
  nand_5 g0285(.A(new_n600), .B(new_n596), .Y(new_n601));
  and_6  g0286(.A(new_n601), .B(new_n594), .Y(new_n602));
  nand_5 g0287(.A(new_n602), .B(new_n593), .Y(new_n603));
  or_6   g0288(.A(new_n317), .B(pi055), .Y(new_n604));
  nand_5 g0289(.A(new_n604), .B(new_n473), .Y(new_n605));
  nand_5 g0290(.A(pi150), .B(pi083), .Y(new_n606));
  or_6   g0291(.A(pi150), .B(pi098), .Y(new_n607));
  nand_5 g0292(.A(new_n607), .B(new_n606), .Y(new_n608));
  nor_5  g0293(.A(new_n608), .B(new_n605), .Y(new_n609));
  nor_5  g0294(.A(new_n600), .B(new_n596), .Y(new_n610));
  nor_5  g0295(.A(new_n610), .B(new_n609), .Y(new_n611));
  nand_5 g0296(.A(new_n611), .B(new_n603), .Y(new_n612));
  or_6   g0297(.A(new_n317), .B(pi067), .Y(new_n613));
  nand_5 g0298(.A(new_n613), .B(new_n465), .Y(new_n614));
  nand_5 g0299(.A(pi150), .B(pi027), .Y(new_n615));
  or_6   g0300(.A(pi150), .B(pi029), .Y(new_n616));
  nand_5 g0301(.A(new_n616), .B(new_n615), .Y(new_n617));
  nand_5 g0302(.A(new_n617), .B(new_n614), .Y(new_n618));
  nand_5 g0303(.A(new_n608), .B(new_n605), .Y(new_n619));
  and_6  g0304(.A(new_n619), .B(new_n618), .Y(new_n620));
  nand_5 g0305(.A(new_n620), .B(new_n612), .Y(new_n621));
  nor_5  g0306(.A(new_n617), .B(new_n614), .Y(new_n622));
  or_6   g0307(.A(new_n317), .B(pi059), .Y(new_n623));
  nand_5 g0308(.A(new_n623), .B(new_n459), .Y(new_n624));
  not_8  g0309(.A(new_n624), .Y(new_n625));
  or_6   g0310(.A(pi180), .B(new_n317), .Y(new_n626));
  nand_5 g0311(.A(new_n317), .B(pi023), .Y(new_n627));
  nand_5 g0312(.A(new_n627), .B(new_n626), .Y(new_n628));
  and_6  g0313(.A(new_n628), .B(new_n625), .Y(new_n629));
  nor_5  g0314(.A(new_n629), .B(new_n622), .Y(new_n630));
  nand_5 g0315(.A(new_n630), .B(new_n621), .Y(new_n631));
  nor_5  g0316(.A(new_n628), .B(new_n625), .Y(new_n632));
  or_6   g0317(.A(new_n317), .B(pi038), .Y(new_n633));
  nand_5 g0318(.A(new_n633), .B(new_n451), .Y(new_n634));
  nand_5 g0319(.A(pi150), .B(pi074), .Y(new_n635));
  not_8  g0320(.A(new_n635), .Y(new_n636));
  nor_5  g0321(.A(pi150), .B(pi117), .Y(new_n637));
  nor_5  g0322(.A(new_n637), .B(new_n636), .Y(new_n638));
  not_8  g0323(.A(new_n638), .Y(new_n639));
  and_6  g0324(.A(new_n639), .B(new_n634), .Y(new_n640));
  nor_5  g0325(.A(new_n640), .B(new_n632), .Y(new_n641));
  nand_5 g0326(.A(new_n641), .B(new_n631), .Y(new_n642));
  nor_5  g0327(.A(new_n639), .B(new_n634), .Y(new_n643));
  or_6   g0328(.A(pi206), .B(new_n317), .Y(new_n644));
  nand_5 g0329(.A(new_n644), .B(new_n447), .Y(new_n645));
  nand_5 g0330(.A(pi150), .B(pi051), .Y(new_n646));
  or_6   g0331(.A(pi150), .B(pi100), .Y(new_n647));
  nand_5 g0332(.A(new_n647), .B(new_n646), .Y(new_n648));
  nor_5  g0333(.A(new_n648), .B(new_n645), .Y(new_n649));
  nor_5  g0334(.A(new_n649), .B(new_n643), .Y(new_n650));
  nand_5 g0335(.A(new_n650), .B(new_n642), .Y(new_n651));
  or_6   g0336(.A(new_n317), .B(pi135), .Y(new_n652));
  nand_5 g0337(.A(new_n652), .B(new_n425), .Y(new_n653));
  nor_5  g0338(.A(pi201), .B(pi150), .Y(new_n654));
  nand_5 g0339(.A(pi150), .B(pi020), .Y(new_n655));
  not_8  g0340(.A(new_n655), .Y(new_n656));
  nor_5  g0341(.A(new_n656), .B(new_n654), .Y(new_n657));
  not_8  g0342(.A(new_n657), .Y(new_n658));
  nand_5 g0343(.A(new_n658), .B(new_n653), .Y(new_n659));
  or_6   g0344(.A(new_n317), .B(pi049), .Y(new_n660));
  nand_5 g0345(.A(new_n660), .B(new_n429), .Y(new_n661));
  not_8  g0346(.A(new_n661), .Y(new_n662));
  or_6   g0347(.A(pi170), .B(new_n317), .Y(new_n663));
  nand_5 g0348(.A(new_n317), .B(pi149), .Y(new_n664));
  nand_5 g0349(.A(new_n664), .B(new_n663), .Y(new_n665));
  or_6   g0350(.A(new_n665), .B(new_n662), .Y(new_n666));
  nand_5 g0351(.A(new_n666), .B(new_n659), .Y(new_n667));
  or_6   g0352(.A(new_n658), .B(new_n653), .Y(new_n668));
  nand_5 g0353(.A(new_n648), .B(new_n645), .Y(new_n669));
  nand_5 g0354(.A(new_n669), .B(new_n668), .Y(new_n670));
  nor_5  g0355(.A(new_n670), .B(new_n667), .Y(new_n671));
  nand_5 g0356(.A(new_n671), .B(new_n651), .Y(new_n672));
  and_6  g0357(.A(new_n665), .B(new_n662), .Y(new_n673));
  and_6  g0358(.A(new_n673), .B(new_n659), .Y(new_n674));
  or_6   g0359(.A(new_n317), .B(pi011), .Y(new_n675));
  nand_5 g0360(.A(new_n675), .B(new_n420), .Y(new_n676));
  not_8  g0361(.A(new_n676), .Y(new_n677));
  nand_5 g0362(.A(pi150), .B(pi107), .Y(new_n678));
  not_8  g0363(.A(new_n678), .Y(new_n679));
  nor_5  g0364(.A(pi150), .B(pi113), .Y(new_n680));
  nor_5  g0365(.A(new_n680), .B(new_n679), .Y(new_n681));
  nand_5 g0366(.A(new_n681), .B(new_n677), .Y(new_n682));
  nand_5 g0367(.A(new_n682), .B(new_n668), .Y(new_n683));
  nor_5  g0368(.A(new_n683), .B(new_n674), .Y(new_n684));
  nand_5 g0369(.A(new_n684), .B(new_n672), .Y(new_n685));
  or_6   g0370(.A(pi195), .B(new_n317), .Y(new_n686));
  nand_5 g0371(.A(new_n686), .B(new_n416), .Y(new_n687));
  or_6   g0372(.A(pi183), .B(new_n317), .Y(new_n688));
  nand_5 g0373(.A(pi166), .B(new_n317), .Y(new_n689));
  nand_5 g0374(.A(new_n689), .B(new_n688), .Y(new_n690));
  not_8  g0375(.A(new_n690), .Y(new_n691));
  and_6  g0376(.A(new_n691), .B(new_n687), .Y(new_n692));
  nor_5  g0377(.A(new_n681), .B(new_n677), .Y(new_n693));
  nor_5  g0378(.A(new_n693), .B(new_n692), .Y(new_n694));
  nand_5 g0379(.A(new_n694), .B(new_n685), .Y(new_n695));
  nand_5 g0380(.A(pi150), .B(pi097), .Y(new_n696));
  nand_5 g0381(.A(new_n696), .B(new_n410), .Y(new_n697));
  nand_5 g0382(.A(pi150), .B(pi057), .Y(new_n698));
  not_8  g0383(.A(new_n698), .Y(new_n699));
  nor_5  g0384(.A(pi150), .B(pi138), .Y(new_n700));
  nor_5  g0385(.A(new_n700), .B(new_n699), .Y(new_n701));
  and_6  g0386(.A(new_n701), .B(new_n697), .Y(new_n702));
  nor_5  g0387(.A(new_n691), .B(new_n687), .Y(new_n703));
  nor_5  g0388(.A(new_n703), .B(new_n702), .Y(new_n704));
  nand_5 g0389(.A(new_n704), .B(new_n695), .Y(new_n705));
  or_6   g0390(.A(new_n317), .B(pi114), .Y(new_n706));
  nand_5 g0391(.A(new_n706), .B(new_n389), .Y(new_n707));
  nand_5 g0392(.A(new_n317), .B(pi016), .Y(new_n708));
  nand_5 g0393(.A(pi150), .B(new_n392), .Y(new_n709));
  nand_5 g0394(.A(new_n709), .B(new_n708), .Y(new_n710));
  not_8  g0395(.A(new_n710), .Y(new_n711));
  nand_5 g0396(.A(new_n711), .B(new_n707), .Y(new_n712));
  or_6   g0397(.A(new_n317), .B(pi005), .Y(new_n713));
  nand_5 g0398(.A(new_n713), .B(new_n395), .Y(new_n714));
  or_6   g0399(.A(pi179), .B(pi150), .Y(new_n715));
  nand_5 g0400(.A(pi150), .B(pi039), .Y(new_n716));
  nand_5 g0401(.A(new_n716), .B(new_n715), .Y(new_n717));
  or_6   g0402(.A(new_n717), .B(new_n714), .Y(new_n718));
  nand_5 g0403(.A(new_n718), .B(new_n712), .Y(new_n719));
  or_6   g0404(.A(new_n701), .B(new_n697), .Y(new_n720));
  nor_5  g0405(.A(new_n711), .B(new_n707), .Y(new_n721));
  and_6  g0406(.A(new_n717), .B(new_n714), .Y(new_n722));
  nor_5  g0407(.A(new_n722), .B(new_n721), .Y(new_n723));
  nand_5 g0408(.A(new_n723), .B(new_n720), .Y(new_n724));
  nor_5  g0409(.A(new_n724), .B(new_n719), .Y(new_n725));
  nand_5 g0410(.A(new_n725), .B(new_n705), .Y(new_n726));
  not_8  g0411(.A(new_n712), .Y(new_n727));
  nor_5  g0412(.A(new_n718), .B(new_n727), .Y(new_n728));
  nor_5  g0413(.A(new_n728), .B(new_n721), .Y(new_n729));
  nand_5 g0414(.A(new_n729), .B(new_n726), .Y(new_n730));
  and_6  g0415(.A(new_n730), .B(new_n568), .Y(new_n731));
  nor_5  g0416(.A(new_n731), .B(new_n565), .Y(new_n732));
  nor_5  g0417(.A(new_n730), .B(new_n568), .Y(new_n733));
  or_6   g0418(.A(new_n733), .B(new_n732), .Y(new_n734));
  nand_5 g0419(.A(new_n734), .B(new_n562), .Y(new_n735));
  nand_5 g0420(.A(new_n735), .B(new_n561), .Y(new_n736));
  or_6   g0421(.A(new_n317), .B(pi095), .Y(new_n737));
  nand_5 g0422(.A(new_n737), .B(new_n316), .Y(new_n738));
  or_6   g0423(.A(pi153), .B(new_n317), .Y(new_n739));
  nand_5 g0424(.A(new_n317), .B(pi003), .Y(new_n740));
  nand_5 g0425(.A(new_n740), .B(new_n739), .Y(new_n741));
  not_8  g0426(.A(new_n741), .Y(new_n742));
  nand_5 g0427(.A(new_n742), .B(new_n738), .Y(new_n743));
  not_8  g0428(.A(pi015), .Y(new_n744));
  nand_5 g0429(.A(pi150), .B(new_n744), .Y(new_n745));
  nand_5 g0430(.A(new_n745), .B(new_n316), .Y(new_n746));
  not_8  g0431(.A(new_n746), .Y(new_n747));
  nand_5 g0432(.A(pi150), .B(pi050), .Y(new_n748));
  not_8  g0433(.A(new_n748), .Y(new_n749));
  nor_5  g0434(.A(pi150), .B(pi065), .Y(new_n750));
  nor_5  g0435(.A(new_n750), .B(new_n749), .Y(new_n751));
  nand_5 g0436(.A(new_n751), .B(new_n747), .Y(new_n752));
  nand_5 g0437(.A(new_n752), .B(new_n743), .Y(new_n753));
  or_6   g0438(.A(new_n317), .B(pi105), .Y(new_n754));
  nand_5 g0439(.A(new_n754), .B(new_n316), .Y(new_n755));
  nand_5 g0440(.A(pi150), .B(pi056), .Y(new_n756));
  or_6   g0441(.A(pi150), .B(pi141), .Y(new_n757));
  nand_5 g0442(.A(new_n757), .B(new_n756), .Y(new_n758));
  nand_5 g0443(.A(new_n758), .B(new_n755), .Y(new_n759));
  nor_5  g0444(.A(new_n742), .B(new_n738), .Y(new_n760));
  nor_5  g0445(.A(new_n751), .B(new_n747), .Y(new_n761));
  nor_5  g0446(.A(new_n761), .B(new_n760), .Y(new_n762));
  nand_5 g0447(.A(new_n762), .B(new_n759), .Y(new_n763));
  nor_5  g0448(.A(new_n763), .B(new_n753), .Y(new_n764));
  or_6   g0449(.A(new_n317), .B(pi006), .Y(new_n765));
  nand_5 g0450(.A(new_n765), .B(new_n348), .Y(new_n766));
  or_6   g0451(.A(pi199), .B(new_n317), .Y(new_n767));
  nand_5 g0452(.A(pi173), .B(new_n317), .Y(new_n768));
  nand_5 g0453(.A(new_n768), .B(new_n767), .Y(new_n769));
  not_8  g0454(.A(new_n769), .Y(new_n770));
  nand_5 g0455(.A(new_n770), .B(new_n766), .Y(new_n771));
  or_6   g0456(.A(new_n317), .B(pi119), .Y(new_n772));
  nand_5 g0457(.A(new_n772), .B(new_n344), .Y(new_n773));
  or_6   g0458(.A(pi196), .B(new_n317), .Y(new_n774));
  nand_5 g0459(.A(pi161), .B(new_n317), .Y(new_n775));
  nand_5 g0460(.A(new_n775), .B(new_n774), .Y(new_n776));
  not_8  g0461(.A(new_n776), .Y(new_n777));
  nand_5 g0462(.A(new_n777), .B(new_n773), .Y(new_n778));
  nand_5 g0463(.A(new_n778), .B(new_n771), .Y(new_n779));
  or_6   g0464(.A(pi174), .B(new_n317), .Y(new_n780));
  nand_5 g0465(.A(new_n780), .B(new_n353), .Y(new_n781));
  or_6   g0466(.A(pi178), .B(new_n317), .Y(new_n782));
  nand_5 g0467(.A(new_n317), .B(pi140), .Y(new_n783));
  nand_5 g0468(.A(new_n783), .B(new_n782), .Y(new_n784));
  not_8  g0469(.A(new_n784), .Y(new_n785));
  nand_5 g0470(.A(new_n785), .B(new_n781), .Y(new_n786));
  or_6   g0471(.A(new_n317), .B(pi082), .Y(new_n787));
  nand_5 g0472(.A(new_n787), .B(new_n358), .Y(new_n788));
  nor_5  g0473(.A(pi162), .B(new_n317), .Y(new_n789));
  and_6  g0474(.A(new_n317), .B(pi121), .Y(new_n790));
  nor_5  g0475(.A(new_n790), .B(new_n789), .Y(new_n791));
  nand_5 g0476(.A(new_n791), .B(new_n788), .Y(new_n792));
  nand_5 g0477(.A(new_n792), .B(new_n786), .Y(new_n793));
  or_6   g0478(.A(new_n793), .B(new_n779), .Y(new_n794));
  or_6   g0479(.A(new_n317), .B(pi110), .Y(new_n795));
  nand_5 g0480(.A(new_n795), .B(new_n316), .Y(new_n796));
  or_6   g0481(.A(pi190), .B(pi150), .Y(new_n797));
  nand_5 g0482(.A(pi150), .B(pi047), .Y(new_n798));
  nand_5 g0483(.A(new_n798), .B(new_n797), .Y(new_n799));
  nand_5 g0484(.A(new_n799), .B(new_n796), .Y(new_n800));
  not_8  g0485(.A(pi084), .Y(new_n801));
  nand_5 g0486(.A(pi150), .B(new_n801), .Y(new_n802));
  nand_5 g0487(.A(new_n802), .B(new_n316), .Y(new_n803));
  nand_5 g0488(.A(new_n317), .B(pi010), .Y(new_n804));
  or_6   g0489(.A(new_n317), .B(pi122), .Y(new_n805));
  nand_5 g0490(.A(new_n805), .B(new_n804), .Y(new_n806));
  not_8  g0491(.A(new_n806), .Y(new_n807));
  nand_5 g0492(.A(new_n807), .B(new_n803), .Y(new_n808));
  nand_5 g0493(.A(new_n808), .B(new_n800), .Y(new_n809));
  nor_5  g0494(.A(new_n777), .B(new_n773), .Y(new_n810));
  nor_5  g0495(.A(new_n799), .B(new_n796), .Y(new_n811));
  nor_5  g0496(.A(new_n811), .B(new_n810), .Y(new_n812));
  nor_5  g0497(.A(new_n770), .B(new_n766), .Y(new_n813));
  nor_5  g0498(.A(new_n785), .B(new_n781), .Y(new_n814));
  nor_5  g0499(.A(new_n814), .B(new_n813), .Y(new_n815));
  nand_5 g0500(.A(new_n815), .B(new_n812), .Y(new_n816));
  or_6   g0501(.A(new_n816), .B(new_n809), .Y(new_n817));
  nor_5  g0502(.A(new_n817), .B(new_n794), .Y(new_n818));
  nand_5 g0503(.A(new_n818), .B(new_n764), .Y(new_n819));
  nor_5  g0504(.A(new_n819), .B(new_n736), .Y(new_n820));
  nor_5  g0505(.A(new_n791), .B(new_n788), .Y(new_n821));
  nand_5 g0506(.A(new_n821), .B(new_n786), .Y(new_n822));
  and_6  g0507(.A(new_n822), .B(new_n815), .Y(new_n823));
  or_6   g0508(.A(new_n823), .B(new_n779), .Y(new_n824));
  and_6  g0509(.A(new_n824), .B(new_n812), .Y(new_n825));
  or_6   g0510(.A(new_n825), .B(new_n809), .Y(new_n826));
  nor_5  g0511(.A(new_n758), .B(new_n755), .Y(new_n827));
  nor_5  g0512(.A(new_n807), .B(new_n803), .Y(new_n828));
  nor_5  g0513(.A(new_n828), .B(new_n827), .Y(new_n829));
  nand_5 g0514(.A(new_n829), .B(new_n826), .Y(new_n830));
  nand_5 g0515(.A(new_n830), .B(new_n764), .Y(new_n831));
  not_8  g0516(.A(new_n743), .Y(new_n832));
  nor_5  g0517(.A(new_n752), .B(new_n832), .Y(new_n833));
  nor_5  g0518(.A(new_n833), .B(new_n760), .Y(new_n834));
  nand_5 g0519(.A(new_n834), .B(new_n831), .Y(new_n835));
  nor_5  g0520(.A(new_n835), .B(new_n820), .Y(new_n836));
  or_6   g0521(.A(pi204), .B(new_n317), .Y(new_n837));
  nand_5 g0522(.A(new_n317), .B(pi088), .Y(new_n838));
  nand_5 g0523(.A(new_n838), .B(new_n837), .Y(new_n839));
  or_6   g0524(.A(new_n839), .B(new_n316), .Y(new_n840));
  or_6   g0525(.A(new_n317), .B(pi028), .Y(new_n841));
  nand_5 g0526(.A(new_n841), .B(new_n316), .Y(new_n842));
  or_6   g0527(.A(pi181), .B(new_n317), .Y(new_n843));
  nand_5 g0528(.A(new_n317), .B(pi041), .Y(new_n844));
  nand_5 g0529(.A(new_n844), .B(new_n843), .Y(new_n845));
  not_8  g0530(.A(new_n845), .Y(new_n846));
  nand_5 g0531(.A(new_n846), .B(new_n842), .Y(new_n847));
  nand_5 g0532(.A(new_n847), .B(new_n840), .Y(new_n848));
  nor_5  g0533(.A(new_n846), .B(new_n842), .Y(new_n849));
  not_8  g0534(.A(new_n849), .Y(new_n850));
  or_6   g0535(.A(pi185), .B(new_n317), .Y(new_n851));
  and_6  g0536(.A(new_n851), .B(new_n316), .Y(new_n852));
  nand_5 g0537(.A(new_n317), .B(pi019), .Y(new_n853));
  or_6   g0538(.A(new_n317), .B(pi085), .Y(new_n854));
  nand_5 g0539(.A(new_n854), .B(new_n853), .Y(new_n855));
  or_6   g0540(.A(new_n855), .B(new_n852), .Y(new_n856));
  nand_5 g0541(.A(new_n856), .B(new_n850), .Y(new_n857));
  nor_5  g0542(.A(new_n857), .B(new_n848), .Y(new_n858));
  or_6   g0543(.A(new_n317), .B(pi013), .Y(new_n859));
  nand_5 g0544(.A(new_n859), .B(new_n316), .Y(new_n860));
  nand_5 g0545(.A(pi150), .B(pi018), .Y(new_n861));
  or_6   g0546(.A(pi150), .B(pi073), .Y(new_n862));
  nand_5 g0547(.A(new_n862), .B(new_n861), .Y(new_n863));
  nand_5 g0548(.A(new_n863), .B(new_n860), .Y(new_n864));
  or_6   g0549(.A(pi159), .B(new_n317), .Y(new_n865));
  nand_5 g0550(.A(new_n865), .B(new_n316), .Y(new_n866));
  nand_5 g0551(.A(pi150), .B(pi101), .Y(new_n867));
  or_6   g0552(.A(pi150), .B(pi112), .Y(new_n868));
  nand_5 g0553(.A(new_n868), .B(new_n867), .Y(new_n869));
  nand_5 g0554(.A(new_n869), .B(new_n866), .Y(new_n870));
  nand_5 g0555(.A(new_n870), .B(new_n864), .Y(new_n871));
  not_8  g0556(.A(pi124), .Y(new_n872));
  nand_5 g0557(.A(pi078), .B(pi071), .Y(new_n873));
  nand_5 g0558(.A(new_n873), .B(pi022), .Y(new_n874));
  and_6  g0559(.A(new_n874), .B(new_n872), .Y(new_n875));
  not_8  g0560(.A(pi071), .Y(new_n876));
  nand_5 g0561(.A(new_n876), .B(pi022), .Y(new_n877));
  nor_5  g0562(.A(new_n877), .B(new_n872), .Y(new_n878));
  nor_5  g0563(.A(new_n878), .B(new_n875), .Y(new_n879));
  nor_5  g0564(.A(new_n879), .B(new_n871), .Y(new_n880));
  nand_5 g0565(.A(new_n880), .B(new_n858), .Y(new_n881));
  nor_5  g0566(.A(new_n881), .B(new_n836), .Y(new_n882));
  nor_5  g0567(.A(pi078), .B(pi071), .Y(new_n883));
  nand_5 g0568(.A(new_n883), .B(pi022), .Y(new_n884));
  nand_5 g0569(.A(new_n884), .B(pi124), .Y(new_n885));
  nor_5  g0570(.A(new_n869), .B(new_n866), .Y(new_n886));
  and_6  g0571(.A(new_n855), .B(new_n851), .Y(new_n887));
  nor_5  g0572(.A(new_n887), .B(new_n839), .Y(new_n888));
  nand_5 g0573(.A(new_n856), .B(new_n316), .Y(new_n889));
  nor_5  g0574(.A(new_n889), .B(new_n888), .Y(new_n890));
  nor_5  g0575(.A(new_n890), .B(new_n886), .Y(new_n891));
  or_6   g0576(.A(new_n891), .B(new_n871), .Y(new_n892));
  nor_5  g0577(.A(new_n863), .B(new_n860), .Y(new_n893));
  nor_5  g0578(.A(new_n893), .B(new_n849), .Y(new_n894));
  nand_5 g0579(.A(new_n894), .B(new_n892), .Y(new_n895));
  not_8  g0580(.A(new_n847), .Y(new_n896));
  nor_5  g0581(.A(new_n879), .B(new_n896), .Y(new_n897));
  nand_5 g0582(.A(new_n897), .B(new_n895), .Y(new_n898));
  nand_5 g0583(.A(new_n898), .B(new_n885), .Y(new_n899));
  or_6   g0584(.A(new_n899), .B(new_n882), .Y(po008));
  nor_5  g0585(.A(new_n342), .B(new_n341), .Y(new_n901));
  xor_4  g0586(.A(new_n901), .B(new_n538), .Y(po009));
  xor_4  g0587(.A(new_n540), .B(new_n337), .Y(po011));
  or_6   g0588(.A(new_n317), .B(pi062), .Y(new_n904));
  nand_5 g0589(.A(new_n904), .B(new_n316), .Y(new_n905));
  nand_5 g0590(.A(new_n905), .B(pi101), .Y(new_n906));
  or_6   g0591(.A(new_n905), .B(pi101), .Y(new_n907));
  nand_5 g0592(.A(new_n907), .B(new_n906), .Y(new_n908));
  or_6   g0593(.A(new_n317), .B(pi145), .Y(new_n909));
  nand_5 g0594(.A(new_n909), .B(new_n316), .Y(new_n910));
  or_6   g0595(.A(new_n910), .B(pi085), .Y(new_n911));
  nand_5 g0596(.A(new_n910), .B(pi085), .Y(new_n912));
  or_6   g0597(.A(new_n317), .B(pi061), .Y(new_n913));
  nand_5 g0598(.A(new_n913), .B(new_n316), .Y(new_n914));
  nor_5  g0599(.A(new_n914), .B(pi204), .Y(new_n915));
  not_8  g0600(.A(new_n915), .Y(new_n916));
  nand_5 g0601(.A(new_n319), .B(pi153), .Y(new_n917));
  nand_5 g0602(.A(new_n546), .B(new_n320), .Y(new_n918));
  nand_5 g0603(.A(new_n918), .B(new_n917), .Y(new_n919));
  nand_5 g0604(.A(new_n914), .B(pi204), .Y(new_n920));
  nand_5 g0605(.A(new_n920), .B(new_n916), .Y(new_n921));
  or_6   g0606(.A(new_n921), .B(new_n919), .Y(new_n922));
  nand_5 g0607(.A(new_n922), .B(new_n916), .Y(new_n923));
  nand_5 g0608(.A(new_n923), .B(new_n912), .Y(new_n924));
  nand_5 g0609(.A(new_n924), .B(new_n911), .Y(new_n925));
  xnor_4 g0610(.A(new_n925), .B(new_n908), .Y(po013));
  nand_5 g0611(.A(new_n469), .B(new_n454), .Y(new_n927));
  not_8  g0612(.A(new_n469), .Y(new_n928));
  nand_5 g0613(.A(new_n928), .B(new_n455), .Y(new_n929));
  nand_5 g0614(.A(new_n929), .B(new_n927), .Y(new_n930));
  xor_4  g0615(.A(new_n930), .B(new_n470), .Y(new_n931));
  or_6   g0616(.A(new_n931), .B(new_n517), .Y(new_n932));
  nor_5  g0617(.A(new_n471), .B(new_n462), .Y(new_n933));
  nand_5 g0618(.A(new_n933), .B(new_n454), .Y(new_n934));
  not_8  g0619(.A(new_n933), .Y(new_n935));
  nand_5 g0620(.A(new_n935), .B(new_n455), .Y(new_n936));
  nand_5 g0621(.A(new_n936), .B(new_n934), .Y(new_n937));
  xor_4  g0622(.A(new_n937), .B(new_n467), .Y(new_n938));
  nand_5 g0623(.A(new_n938), .B(new_n517), .Y(new_n939));
  nand_5 g0624(.A(new_n939), .B(new_n932), .Y(new_n940));
  not_8  g0625(.A(new_n505), .Y(new_n941));
  nand_5 g0626(.A(new_n941), .B(new_n498), .Y(new_n942));
  nand_5 g0627(.A(new_n942), .B(new_n497), .Y(new_n943));
  not_8  g0628(.A(new_n499), .Y(new_n944));
  xor_4  g0629(.A(new_n506), .B(new_n492), .Y(new_n945));
  xor_4  g0630(.A(new_n945), .B(new_n476), .Y(new_n946));
  xor_4  g0631(.A(new_n946), .B(new_n485), .Y(new_n947));
  xor_4  g0632(.A(new_n947), .B(new_n944), .Y(new_n948));
  xor_4  g0633(.A(new_n948), .B(new_n943), .Y(new_n949));
  nand_5 g0634(.A(new_n507), .B(new_n493), .Y(new_n950));
  nor_5  g0635(.A(new_n950), .B(new_n499), .Y(new_n951));
  and_6  g0636(.A(new_n951), .B(new_n484), .Y(new_n952));
  not_8  g0637(.A(new_n951), .Y(new_n953));
  not_8  g0638(.A(new_n489), .Y(new_n954));
  nor_5  g0639(.A(new_n943), .B(new_n954), .Y(new_n955));
  nand_5 g0640(.A(new_n955), .B(new_n953), .Y(new_n956));
  nand_5 g0641(.A(new_n956), .B(new_n491), .Y(new_n957));
  nand_5 g0642(.A(new_n957), .B(new_n484), .Y(new_n958));
  nand_5 g0643(.A(new_n958), .B(new_n482), .Y(new_n959));
  or_6   g0644(.A(new_n959), .B(new_n952), .Y(new_n960));
  xor_4  g0645(.A(new_n960), .B(new_n949), .Y(new_n961));
  nand_5 g0646(.A(new_n957), .B(new_n505), .Y(new_n962));
  nor_5  g0647(.A(new_n951), .B(new_n941), .Y(new_n963));
  or_6   g0648(.A(new_n963), .B(new_n957), .Y(new_n964));
  nand_5 g0649(.A(new_n964), .B(new_n962), .Y(new_n965));
  nor_5  g0650(.A(new_n965), .B(new_n961), .Y(new_n966));
  nand_5 g0651(.A(new_n965), .B(new_n961), .Y(new_n967));
  nand_5 g0652(.A(new_n967), .B(pi070), .Y(new_n968));
  or_6   g0653(.A(new_n968), .B(new_n966), .Y(new_n969));
  nand_5 g0654(.A(new_n502), .B(new_n497), .Y(new_n970));
  nand_5 g0655(.A(new_n503), .B(new_n498), .Y(new_n971));
  nand_5 g0656(.A(new_n971), .B(new_n970), .Y(new_n972));
  xor_4  g0657(.A(new_n972), .B(new_n957), .Y(new_n973));
  xor_4  g0658(.A(new_n959), .B(new_n948), .Y(new_n974));
  nand_5 g0659(.A(new_n974), .B(new_n973), .Y(new_n975));
  nor_5  g0660(.A(new_n974), .B(new_n973), .Y(new_n976));
  nor_5  g0661(.A(new_n976), .B(pi070), .Y(new_n977));
  nand_5 g0662(.A(new_n977), .B(new_n975), .Y(new_n978));
  nand_5 g0663(.A(new_n978), .B(new_n969), .Y(new_n979));
  or_6   g0664(.A(new_n463), .B(new_n462), .Y(new_n980));
  xor_4  g0665(.A(new_n457), .B(new_n450), .Y(new_n981));
  xor_4  g0666(.A(new_n981), .B(new_n980), .Y(new_n982));
  xor_4  g0667(.A(new_n982), .B(new_n979), .Y(new_n983));
  xor_4  g0668(.A(new_n983), .B(new_n940), .Y(po015));
  xor_4  g0669(.A(new_n417), .B(pi183), .Y(new_n985));
  nand_5 g0670(.A(new_n527), .B(new_n437), .Y(new_n986));
  xor_4  g0671(.A(new_n986), .B(new_n985), .Y(po016));
  not_8  g0672(.A(pi125), .Y(po017));
  and_6  g0673(.A(pi109), .B(pi060), .Y(po020));
  xor_4  g0674(.A(new_n544), .B(new_n325), .Y(po024));
  nand_5 g0675(.A(new_n414), .B(new_n413), .Y(new_n991));
  xor_4  g0676(.A(new_n991), .B(new_n529), .Y(po025));
  nand_5 g0677(.A(new_n916), .B(new_n911), .Y(new_n993));
  nand_5 g0678(.A(new_n993), .B(new_n912), .Y(new_n994));
  nand_5 g0679(.A(new_n994), .B(new_n907), .Y(new_n995));
  nand_5 g0680(.A(new_n995), .B(new_n906), .Y(new_n996));
  not_8  g0681(.A(new_n921), .Y(new_n997));
  nand_5 g0682(.A(new_n912), .B(new_n911), .Y(new_n998));
  not_8  g0683(.A(new_n998), .Y(new_n999));
  nand_5 g0684(.A(new_n999), .B(new_n997), .Y(new_n1000));
  nor_5  g0685(.A(new_n1000), .B(new_n908), .Y(new_n1001));
  not_8  g0686(.A(new_n1001), .Y(new_n1002));
  nand_5 g0687(.A(new_n1002), .B(new_n920), .Y(new_n1003));
  nand_5 g0688(.A(new_n1003), .B(new_n996), .Y(new_n1004));
  not_8  g0689(.A(new_n996), .Y(new_n1005));
  nand_5 g0690(.A(new_n1005), .B(new_n920), .Y(new_n1006));
  nand_5 g0691(.A(new_n1006), .B(new_n1004), .Y(new_n1007));
  nor_5  g0692(.A(new_n999), .B(new_n997), .Y(new_n1008));
  or_6   g0693(.A(pi184), .B(new_n317), .Y(new_n1009));
  nand_5 g0694(.A(new_n1009), .B(new_n316), .Y(new_n1010));
  nand_5 g0695(.A(new_n1010), .B(pi018), .Y(new_n1011));
  nor_5  g0696(.A(new_n1010), .B(pi018), .Y(new_n1012));
  nor_5  g0697(.A(new_n1012), .B(new_n1005), .Y(new_n1013));
  not_8  g0698(.A(new_n1013), .Y(new_n1014));
  nand_5 g0699(.A(new_n1014), .B(new_n1011), .Y(new_n1015));
  nand_5 g0700(.A(new_n1011), .B(new_n1001), .Y(new_n1016));
  nand_5 g0701(.A(new_n1016), .B(new_n1015), .Y(new_n1017));
  xor_4  g0702(.A(new_n1017), .B(new_n1008), .Y(new_n1018));
  xor_4  g0703(.A(new_n1018), .B(new_n1007), .Y(new_n1019));
  or_6   g0704(.A(new_n1019), .B(new_n919), .Y(new_n1020));
  xor_4  g0705(.A(new_n998), .B(new_n921), .Y(new_n1021));
  xor_4  g0706(.A(new_n1021), .B(new_n1015), .Y(new_n1022));
  xor_4  g0707(.A(new_n996), .B(new_n915), .Y(new_n1023));
  xor_4  g0708(.A(new_n1023), .B(new_n1022), .Y(new_n1024));
  nand_5 g0709(.A(new_n1024), .B(new_n919), .Y(new_n1025));
  nand_5 g0710(.A(new_n1025), .B(new_n1020), .Y(new_n1026));
  nand_5 g0711(.A(pi024), .B(pi022), .Y(new_n1027));
  nand_5 g0712(.A(new_n1027), .B(new_n872), .Y(new_n1028));
  xor_4  g0713(.A(new_n1027), .B(pi124), .Y(new_n1029));
  not_8  g0714(.A(pi077), .Y(new_n1030));
  nand_5 g0715(.A(pi150), .B(new_n1030), .Y(new_n1031));
  nand_5 g0716(.A(new_n1031), .B(new_n316), .Y(new_n1032));
  nand_5 g0717(.A(new_n1032), .B(pi181), .Y(new_n1033));
  or_6   g0718(.A(new_n1032), .B(pi181), .Y(new_n1034));
  or_6   g0719(.A(new_n1002), .B(new_n919), .Y(new_n1035));
  nand_5 g0720(.A(new_n1035), .B(new_n1013), .Y(new_n1036));
  nand_5 g0721(.A(new_n1036), .B(new_n1011), .Y(new_n1037));
  nand_5 g0722(.A(new_n1037), .B(new_n1034), .Y(new_n1038));
  nand_5 g0723(.A(new_n1038), .B(new_n1033), .Y(new_n1039));
  or_6   g0724(.A(new_n1039), .B(new_n1029), .Y(new_n1040));
  nand_5 g0725(.A(new_n1040), .B(new_n1028), .Y(new_n1041));
  nand_5 g0726(.A(new_n1034), .B(new_n1033), .Y(new_n1042));
  xor_4  g0727(.A(new_n1042), .B(new_n994), .Y(new_n1043));
  xor_4  g0728(.A(new_n1043), .B(new_n908), .Y(new_n1044));
  nand_5 g0729(.A(pi064), .B(pi022), .Y(new_n1045));
  xor_4  g0730(.A(new_n1010), .B(pi018), .Y(new_n1046));
  xor_4  g0731(.A(new_n1046), .B(new_n1045), .Y(new_n1047));
  xor_4  g0732(.A(new_n1047), .B(new_n1044), .Y(new_n1048));
  xor_4  g0733(.A(new_n1048), .B(new_n1041), .Y(new_n1049));
  xor_4  g0734(.A(new_n1049), .B(new_n1026), .Y(po026));
  nor_5  g0735(.A(new_n333), .B(new_n330), .Y(new_n1051));
  nand_5 g0736(.A(new_n1051), .B(new_n541), .Y(new_n1052));
  nand_5 g0737(.A(new_n335), .B(new_n330), .Y(new_n1053));
  not_8  g0738(.A(new_n1053), .Y(new_n1054));
  nand_5 g0739(.A(new_n1054), .B(new_n542), .Y(new_n1055));
  and_6  g0740(.A(new_n1055), .B(new_n1052), .Y(po027));
  nand_5 g0741(.A(new_n1039), .B(new_n1029), .Y(new_n1057));
  and_6  g0742(.A(new_n1045), .B(pi124), .Y(new_n1058));
  nand_5 g0743(.A(pi064), .B(pi024), .Y(new_n1059));
  nor_5  g0744(.A(pi064), .B(pi024), .Y(new_n1060));
  nand_5 g0745(.A(new_n872), .B(pi022), .Y(new_n1061));
  nor_5  g0746(.A(new_n1061), .B(new_n1060), .Y(new_n1062));
  and_6  g0747(.A(new_n1062), .B(new_n1059), .Y(new_n1063));
  nor_5  g0748(.A(new_n1063), .B(new_n1058), .Y(new_n1064));
  xor_4  g0749(.A(new_n1064), .B(new_n1057), .Y(po029));
  nand_5 g0750(.A(new_n1057), .B(new_n1040), .Y(po030));
  xor_4  g0751(.A(new_n534), .B(new_n382), .Y(po038));
  not_8  g0752(.A(new_n374), .Y(new_n1068));
  nand_5 g0753(.A(new_n1068), .B(new_n356), .Y(new_n1069));
  or_6   g0754(.A(new_n1069), .B(new_n536), .Y(new_n1070));
  nand_5 g0755(.A(new_n1070), .B(new_n363), .Y(new_n1071));
  xor_4  g0756(.A(new_n1071), .B(new_n371), .Y(po039));
  nor_5  g0757(.A(new_n1058), .B(new_n1057), .Y(new_n1073));
  nor_5  g0758(.A(new_n1073), .B(new_n1062), .Y(po040));
  xor_4  g0759(.A(new_n507), .B(pi070), .Y(po043));
  xnor_4 g0760(.A(new_n985), .B(new_n435), .Y(new_n1076));
  xor_4  g0761(.A(new_n1076), .B(new_n991), .Y(new_n1077));
  not_8  g0762(.A(new_n442), .Y(new_n1078));
  xor_4  g0763(.A(new_n443), .B(new_n1078), .Y(new_n1079));
  not_8  g0764(.A(new_n439), .Y(new_n1080));
  nand_5 g0765(.A(new_n1080), .B(new_n418), .Y(new_n1081));
  xor_4  g0766(.A(new_n1081), .B(new_n441), .Y(new_n1082));
  xor_4  g0767(.A(new_n1082), .B(new_n437), .Y(new_n1083));
  xor_4  g0768(.A(new_n1083), .B(new_n1079), .Y(new_n1084));
  xor_4  g0769(.A(new_n1084), .B(new_n1077), .Y(new_n1085));
  nand_5 g0770(.A(new_n1085), .B(new_n523), .Y(new_n1086));
  nand_5 g0771(.A(new_n1078), .B(new_n441), .Y(new_n1087));
  nor_5  g0772(.A(new_n1087), .B(new_n444), .Y(new_n1088));
  and_6  g0773(.A(new_n1088), .B(new_n418), .Y(new_n1089));
  or_6   g0774(.A(new_n1089), .B(new_n1082), .Y(new_n1090));
  nor_5  g0775(.A(new_n445), .B(new_n1078), .Y(new_n1091));
  xor_4  g0776(.A(new_n1091), .B(new_n1077), .Y(new_n1092));
  xor_4  g0777(.A(new_n1092), .B(new_n1090), .Y(new_n1093));
  not_8  g0778(.A(new_n1088), .Y(new_n1094));
  nand_5 g0779(.A(new_n1094), .B(new_n443), .Y(new_n1095));
  nor_5  g0780(.A(new_n1095), .B(new_n438), .Y(new_n1096));
  nor_5  g0781(.A(new_n443), .B(new_n437), .Y(new_n1097));
  nor_5  g0782(.A(new_n1097), .B(new_n1096), .Y(new_n1098));
  xor_4  g0783(.A(new_n1098), .B(new_n1093), .Y(new_n1099));
  nand_5 g0784(.A(new_n1099), .B(new_n524), .Y(new_n1100));
  nand_5 g0785(.A(new_n1100), .B(new_n1086), .Y(new_n1101));
  nand_5 g0786(.A(new_n402), .B(new_n386), .Y(new_n1102));
  nand_5 g0787(.A(new_n407), .B(new_n386), .Y(new_n1103));
  nand_5 g0788(.A(new_n1103), .B(new_n1102), .Y(new_n1104));
  nor_5  g0789(.A(new_n404), .B(pi116), .Y(new_n1105));
  nand_5 g0790(.A(new_n399), .B(new_n392), .Y(new_n1106));
  nand_5 g0791(.A(new_n1106), .B(new_n404), .Y(new_n1107));
  nand_5 g0792(.A(new_n1107), .B(new_n393), .Y(new_n1108));
  nand_5 g0793(.A(new_n398), .B(new_n394), .Y(new_n1109));
  nand_5 g0794(.A(new_n1109), .B(new_n1108), .Y(new_n1110));
  nor_5  g0795(.A(new_n1110), .B(new_n1105), .Y(new_n1111));
  and_6  g0796(.A(new_n387), .B(new_n386), .Y(new_n1112));
  xor_4  g0797(.A(new_n1112), .B(new_n382), .Y(new_n1113));
  xor_4  g0798(.A(new_n1113), .B(new_n1111), .Y(new_n1114));
  xor_4  g0799(.A(new_n1114), .B(new_n1104), .Y(new_n1115));
  or_6   g0800(.A(new_n1115), .B(new_n531), .Y(new_n1116));
  nand_5 g0801(.A(new_n1110), .B(pi116), .Y(new_n1117));
  nor_5  g0802(.A(new_n1107), .B(new_n393), .Y(new_n1118));
  nor_5  g0803(.A(new_n1118), .B(new_n1105), .Y(new_n1119));
  nand_5 g0804(.A(new_n1119), .B(new_n1117), .Y(new_n1120));
  xor_4  g0805(.A(new_n1113), .B(new_n1102), .Y(new_n1121));
  xor_4  g0806(.A(new_n1121), .B(new_n1120), .Y(new_n1122));
  nand_5 g0807(.A(new_n1122), .B(new_n531), .Y(new_n1123));
  nand_5 g0808(.A(new_n1123), .B(new_n1116), .Y(new_n1124));
  xor_4  g0809(.A(new_n1124), .B(new_n1101), .Y(po044));
  nand_5 g0810(.A(pi126), .B(pi046), .Y(new_n1126));
  nand_5 g0811(.A(pi191), .B(pi176), .Y(new_n1127));
  nor_5  g0812(.A(new_n1127), .B(new_n1126), .Y(new_n1128));
  not_8  g0813(.A(new_n1128), .Y(po047));
  nand_5 g0814(.A(new_n525), .B(new_n432), .Y(new_n1130));
  xor_4  g0815(.A(new_n1130), .B(new_n1078), .Y(po048));
  xor_4  g0816(.A(new_n521), .B(new_n450), .Y(po049));
  or_6   g0817(.A(pi165), .B(pi148), .Y(po050));
  xor_4  g0818(.A(new_n511), .B(new_n492), .Y(po054));
  and_6  g0819(.A(new_n347), .B(new_n346), .Y(new_n1135));
  not_8  g0820(.A(new_n536), .Y(new_n1136));
  nand_5 g0821(.A(new_n1136), .B(new_n375), .Y(new_n1137));
  nand_5 g0822(.A(new_n1137), .B(new_n365), .Y(new_n1138));
  xor_4  g0823(.A(new_n1138), .B(new_n1135), .Y(po057));
  xor_4  g0824(.A(new_n921), .B(new_n919), .Y(po058));
  xnor_4 g0825(.A(new_n799), .B(new_n758), .Y(new_n1141));
  xor_4  g0826(.A(new_n1141), .B(new_n751), .Y(new_n1142));
  or_6   g0827(.A(pi202), .B(pi150), .Y(new_n1143));
  nand_5 g0828(.A(pi150), .B(pi001), .Y(new_n1144));
  nand_5 g0829(.A(new_n1144), .B(new_n1143), .Y(new_n1145));
  xor_4  g0830(.A(new_n791), .B(new_n784), .Y(new_n1146));
  xor_4  g0831(.A(new_n1146), .B(new_n776), .Y(new_n1147));
  xor_4  g0832(.A(new_n1147), .B(new_n741), .Y(new_n1148));
  xor_4  g0833(.A(new_n1148), .B(new_n1145), .Y(new_n1149));
  xor_4  g0834(.A(new_n1149), .B(new_n1142), .Y(new_n1150));
  xor_4  g0835(.A(new_n1150), .B(new_n806), .Y(new_n1151));
  xor_4  g0836(.A(new_n1151), .B(new_n769), .Y(new_n1152));
  xor_4  g0837(.A(new_n639), .B(new_n628), .Y(new_n1153));
  xor_4  g0838(.A(new_n1153), .B(new_n617), .Y(new_n1154));
  nand_5 g0839(.A(pi150), .B(new_n500), .Y(new_n1155));
  nand_5 g0840(.A(new_n1155), .B(new_n582), .Y(new_n1156));
  xor_4  g0841(.A(new_n608), .B(new_n599), .Y(new_n1157));
  xor_4  g0842(.A(new_n1157), .B(new_n1156), .Y(new_n1158));
  xor_4  g0843(.A(new_n1158), .B(new_n579), .Y(new_n1159));
  or_6   g0844(.A(pi150), .B(pi021), .Y(new_n1160));
  nand_5 g0845(.A(pi150), .B(pi137), .Y(new_n1161));
  nand_5 g0846(.A(new_n1161), .B(new_n1160), .Y(new_n1162));
  xor_4  g0847(.A(new_n1162), .B(new_n575), .Y(new_n1163));
  xor_4  g0848(.A(new_n1163), .B(new_n648), .Y(new_n1164));
  xor_4  g0849(.A(new_n1164), .B(new_n1159), .Y(new_n1165));
  nand_5 g0850(.A(new_n1165), .B(new_n1154), .Y(new_n1166));
  nor_5  g0851(.A(new_n1165), .B(new_n1154), .Y(new_n1167));
  or_6   g0852(.A(new_n317), .B(pi108), .Y(new_n1168));
  nand_5 g0853(.A(pi163), .B(new_n317), .Y(new_n1169));
  nand_5 g0854(.A(new_n1169), .B(new_n1168), .Y(new_n1170));
  xor_4  g0855(.A(new_n1170), .B(new_n863), .Y(new_n1171));
  xor_4  g0856(.A(new_n855), .B(new_n839), .Y(new_n1172));
  xor_4  g0857(.A(new_n869), .B(new_n845), .Y(new_n1173));
  xor_4  g0858(.A(new_n1173), .B(new_n1172), .Y(new_n1174));
  xor_4  g0859(.A(pi064), .B(pi024), .Y(new_n1175));
  nor_5  g0860(.A(new_n1175), .B(new_n317), .Y(new_n1176));
  xor_4  g0861(.A(pi078), .B(pi071), .Y(new_n1177));
  nor_5  g0862(.A(new_n1177), .B(pi150), .Y(new_n1178));
  nor_5  g0863(.A(new_n1178), .B(new_n1176), .Y(new_n1179));
  xor_4  g0864(.A(new_n1179), .B(new_n1174), .Y(new_n1180));
  xor_4  g0865(.A(new_n1180), .B(new_n1171), .Y(new_n1181));
  xor_4  g0866(.A(new_n565), .B(new_n560), .Y(new_n1182));
  xor_4  g0867(.A(new_n717), .B(new_n710), .Y(new_n1183));
  xor_4  g0868(.A(new_n1183), .B(new_n1182), .Y(new_n1184));
  xor_4  g0869(.A(new_n681), .B(new_n657), .Y(new_n1185));
  xor_4  g0870(.A(new_n1185), .B(new_n665), .Y(new_n1186));
  or_6   g0871(.A(pi205), .B(pi150), .Y(new_n1187));
  nand_5 g0872(.A(pi150), .B(pi118), .Y(new_n1188));
  nand_5 g0873(.A(new_n1188), .B(new_n1187), .Y(new_n1189));
  xor_4  g0874(.A(new_n1189), .B(new_n690), .Y(new_n1190));
  xor_4  g0875(.A(new_n1190), .B(new_n701), .Y(new_n1191));
  xor_4  g0876(.A(new_n1191), .B(new_n1186), .Y(new_n1192));
  xor_4  g0877(.A(new_n1192), .B(new_n1184), .Y(new_n1193));
  nand_5 g0878(.A(new_n1193), .B(new_n1181), .Y(new_n1194));
  nor_5  g0879(.A(new_n1194), .B(new_n1167), .Y(new_n1195));
  nand_5 g0880(.A(new_n1195), .B(new_n1166), .Y(new_n1196));
  nor_5  g0881(.A(new_n1196), .B(new_n1152), .Y(new_n1197));
  or_6   g0882(.A(new_n317), .B(pi120), .Y(new_n1198));
  nand_5 g0883(.A(new_n1198), .B(new_n585), .Y(new_n1199));
  xor_4  g0884(.A(new_n1199), .B(new_n448), .Y(new_n1200));
  xor_4  g0885(.A(new_n1200), .B(new_n466), .Y(new_n1201));
  or_6   g0886(.A(pi150), .B(pi040), .Y(new_n1202));
  or_6   g0887(.A(pi155), .B(new_n317), .Y(new_n1203));
  nand_5 g0888(.A(new_n1203), .B(new_n1202), .Y(new_n1204));
  xor_4  g0889(.A(new_n488), .B(new_n474), .Y(new_n1205));
  xor_4  g0890(.A(new_n1205), .B(new_n480), .Y(new_n1206));
  xor_4  g0891(.A(new_n1206), .B(new_n460), .Y(new_n1207));
  xor_4  g0892(.A(new_n1207), .B(new_n1204), .Y(new_n1208));
  xor_4  g0893(.A(new_n1208), .B(new_n1201), .Y(new_n1209));
  xor_4  g0894(.A(new_n1209), .B(new_n453), .Y(new_n1210));
  or_6   g0895(.A(new_n1210), .B(new_n496), .Y(new_n1211));
  xor_4  g0896(.A(new_n412), .B(new_n379), .Y(new_n1212));
  nand_5 g0897(.A(new_n317), .B(pi136), .Y(new_n1213));
  nand_5 g0898(.A(pi150), .B(pi045), .Y(new_n1214));
  nand_5 g0899(.A(new_n1214), .B(new_n1213), .Y(new_n1215));
  xor_4  g0900(.A(new_n1215), .B(new_n427), .Y(new_n1216));
  xor_4  g0901(.A(new_n1216), .B(new_n390), .Y(new_n1217));
  xor_4  g0902(.A(new_n1217), .B(new_n1212), .Y(new_n1218));
  xnor_4 g0903(.A(new_n431), .B(new_n417), .Y(new_n1219));
  xor_4  g0904(.A(new_n1219), .B(new_n422), .Y(new_n1220));
  xor_4  g0905(.A(new_n1220), .B(new_n385), .Y(new_n1221));
  xor_4  g0906(.A(new_n1221), .B(new_n397), .Y(new_n1222));
  xor_4  g0907(.A(new_n1222), .B(new_n1218), .Y(new_n1223));
  xor_4  g0908(.A(pi200), .B(pi102), .Y(new_n1224));
  xor_4  g0909(.A(new_n1224), .B(pi061), .Y(new_n1225));
  xor_4  g0910(.A(pi145), .B(pi062), .Y(new_n1226));
  xor_4  g0911(.A(pi184), .B(new_n1030), .Y(new_n1227));
  xor_4  g0912(.A(new_n1227), .B(new_n1226), .Y(new_n1228));
  nor_5  g0913(.A(new_n1228), .B(new_n1225), .Y(new_n1229));
  nand_5 g0914(.A(new_n316), .B(pi150), .Y(new_n1230));
  and_6  g0915(.A(new_n1228), .B(new_n1225), .Y(new_n1231));
  or_6   g0916(.A(new_n1231), .B(new_n1230), .Y(new_n1232));
  nor_5  g0917(.A(new_n1232), .B(new_n1229), .Y(new_n1233));
  nor_5  g0918(.A(new_n1233), .B(new_n1223), .Y(new_n1234));
  nand_5 g0919(.A(new_n1234), .B(new_n1211), .Y(new_n1235));
  nand_5 g0920(.A(new_n1210), .B(new_n496), .Y(new_n1236));
  nand_5 g0921(.A(new_n317), .B(pi134), .Y(new_n1237));
  nand_5 g0922(.A(pi150), .B(pi017), .Y(new_n1238));
  nand_5 g0923(.A(new_n1238), .B(new_n1237), .Y(new_n1239));
  xor_4  g0924(.A(new_n1239), .B(new_n355), .Y(new_n1240));
  xor_4  g0925(.A(pi154), .B(pi115), .Y(new_n1241));
  xor_4  g0926(.A(pi054), .B(pi026), .Y(new_n1242));
  nand_5 g0927(.A(new_n1242), .B(new_n1241), .Y(new_n1243));
  nor_5  g0928(.A(new_n1242), .B(new_n1241), .Y(new_n1244));
  nor_5  g0929(.A(new_n1244), .B(new_n1230), .Y(new_n1245));
  nand_5 g0930(.A(new_n1245), .B(new_n1243), .Y(new_n1246));
  xor_4  g0931(.A(new_n1246), .B(new_n345), .Y(new_n1247));
  xor_4  g0932(.A(new_n1247), .B(new_n339), .Y(new_n1248));
  xor_4  g0933(.A(new_n1248), .B(new_n350), .Y(new_n1249));
  xor_4  g0934(.A(new_n1249), .B(new_n360), .Y(new_n1250));
  xor_4  g0935(.A(new_n1250), .B(new_n1240), .Y(new_n1251));
  nand_5 g0936(.A(new_n1251), .B(new_n1236), .Y(new_n1252));
  or_6   g0937(.A(new_n1252), .B(new_n1235), .Y(po080));
  or_6   g0938(.A(pi171), .B(new_n317), .Y(new_n1254));
  nand_5 g0939(.A(new_n1254), .B(new_n585), .Y(new_n1255));
  xor_4  g0940(.A(new_n605), .B(new_n570), .Y(new_n1256));
  xor_4  g0941(.A(new_n1256), .B(new_n1255), .Y(new_n1257));
  xor_4  g0942(.A(new_n1257), .B(new_n624), .Y(new_n1258));
  xor_4  g0943(.A(new_n1258), .B(new_n634), .Y(new_n1259));
  or_6   g0944(.A(new_n317), .B(pi129), .Y(new_n1260));
  nand_5 g0945(.A(new_n1260), .B(new_n1202), .Y(new_n1261));
  xor_4  g0946(.A(new_n596), .B(new_n581), .Y(new_n1262));
  xor_4  g0947(.A(new_n1262), .B(new_n1261), .Y(new_n1263));
  xor_4  g0948(.A(new_n1263), .B(new_n614), .Y(new_n1264));
  xor_4  g0949(.A(new_n1264), .B(new_n645), .Y(new_n1265));
  xor_4  g0950(.A(new_n1265), .B(new_n1259), .Y(new_n1266));
  xor_4  g0951(.A(pi185), .B(pi159), .Y(new_n1267));
  xnor_4 g0952(.A(pi168), .B(pi031), .Y(new_n1268));
  xor_4  g0953(.A(new_n1268), .B(pi008), .Y(new_n1269));
  xor_4  g0954(.A(pi028), .B(pi013), .Y(new_n1270));
  xor_4  g0955(.A(new_n1270), .B(new_n1269), .Y(new_n1271));
  nand_5 g0956(.A(new_n1271), .B(new_n1267), .Y(new_n1272));
  nor_5  g0957(.A(new_n1271), .B(new_n1267), .Y(new_n1273));
  nor_5  g0958(.A(new_n1273), .B(new_n1230), .Y(new_n1274));
  nand_5 g0959(.A(new_n1274), .B(new_n1272), .Y(new_n1275));
  nand_5 g0960(.A(new_n1275), .B(new_n1266), .Y(new_n1276));
  xor_4  g0961(.A(pi105), .B(new_n801), .Y(new_n1277));
  nor_5  g0962(.A(new_n1277), .B(new_n1230), .Y(new_n1278));
  xor_4  g0963(.A(new_n1278), .B(new_n788), .Y(new_n1279));
  xor_4  g0964(.A(new_n1279), .B(new_n773), .Y(new_n1280));
  nand_5 g0965(.A(pi150), .B(pi127), .Y(new_n1281));
  nand_5 g0966(.A(new_n1281), .B(new_n1237), .Y(new_n1282));
  xor_4  g0967(.A(pi095), .B(new_n744), .Y(new_n1283));
  nor_5  g0968(.A(new_n1283), .B(new_n1230), .Y(new_n1284));
  nor_5  g0969(.A(new_n1284), .B(new_n796), .Y(new_n1285));
  not_8  g0970(.A(new_n1284), .Y(new_n1286));
  nor_5  g0971(.A(new_n1286), .B(pi110), .Y(new_n1287));
  nor_5  g0972(.A(new_n1287), .B(new_n1285), .Y(new_n1288));
  xor_4  g0973(.A(new_n1288), .B(new_n1282), .Y(new_n1289));
  xor_4  g0974(.A(new_n1289), .B(new_n1280), .Y(new_n1290));
  xor_4  g0975(.A(new_n1290), .B(new_n781), .Y(new_n1291));
  xor_4  g0976(.A(new_n1291), .B(new_n766), .Y(new_n1292));
  nor_5  g0977(.A(new_n1292), .B(new_n1276), .Y(new_n1293));
  xor_4  g0978(.A(new_n697), .B(new_n661), .Y(new_n1294));
  xor_4  g0979(.A(new_n677), .B(new_n653), .Y(new_n1295));
  xor_4  g0980(.A(new_n1295), .B(new_n687), .Y(new_n1296));
  xor_4  g0981(.A(new_n1296), .B(new_n568), .Y(new_n1297));
  nand_5 g0982(.A(pi150), .B(pi072), .Y(new_n1298));
  nand_5 g0983(.A(new_n1298), .B(new_n1213), .Y(new_n1299));
  xor_4  g0984(.A(new_n1299), .B(new_n556), .Y(new_n1300));
  xor_4  g0985(.A(new_n1300), .B(new_n707), .Y(new_n1301));
  xor_4  g0986(.A(new_n1301), .B(new_n1297), .Y(new_n1302));
  xor_4  g0987(.A(new_n1302), .B(new_n714), .Y(new_n1303));
  xor_4  g0988(.A(new_n1303), .B(new_n1294), .Y(new_n1304));
  nand_5 g0989(.A(new_n1304), .B(new_n1293), .Y(po090));
  nor_5  g0990(.A(po047), .B(po006), .Y(new_n1306));
  nand_5 g0991(.A(pi128), .B(pi079), .Y(new_n1307));
  nand_5 g0992(.A(pi157), .B(pi130), .Y(new_n1308));
  nor_5  g0993(.A(new_n1308), .B(new_n1307), .Y(new_n1309));
  not_8  g0994(.A(new_n1309), .Y(po100));
  nand_5 g0995(.A(pi076), .B(pi063), .Y(new_n1311));
  nand_5 g0996(.A(pi133), .B(pi099), .Y(new_n1312));
  nor_5  g0997(.A(new_n1312), .B(new_n1311), .Y(new_n1313));
  not_8  g0998(.A(new_n1313), .Y(po107));
  nor_5  g0999(.A(po107), .B(po100), .Y(new_n1315));
  nand_5 g1000(.A(new_n1315), .B(new_n1306), .Y(new_n1316));
  or_6   g1001(.A(new_n1316), .B(po090), .Y(new_n1317));
  nor_5  g1002(.A(new_n1317), .B(po080), .Y(new_n1318));
  nand_5 g1003(.A(new_n1318), .B(new_n1197), .Y(po059));
  not_8  g1004(.A(new_n526), .Y(new_n1320));
  nand_5 g1005(.A(new_n1320), .B(new_n435), .Y(new_n1321));
  xor_4  g1006(.A(new_n1321), .B(new_n441), .Y(po060));
  xor_4  g1007(.A(new_n1042), .B(new_n1037), .Y(po061));
  xor_4  g1008(.A(new_n466), .B(pi027), .Y(new_n1324));
  xnor_4 g1009(.A(new_n1324), .B(new_n517), .Y(po062));
  nand_5 g1010(.A(pi093), .B(pi053), .Y(new_n1326));
  or_6   g1011(.A(new_n1326), .B(pi165), .Y(po065));
  nand_5 g1012(.A(new_n1136), .B(new_n1068), .Y(new_n1328));
  nand_5 g1013(.A(new_n1328), .B(new_n361), .Y(new_n1329));
  xor_4  g1014(.A(new_n1329), .B(new_n369), .Y(po066));
  xor_4  g1015(.A(new_n513), .B(new_n485), .Y(po067));
  not_8  g1016(.A(new_n405), .Y(new_n1332));
  nand_5 g1017(.A(new_n531), .B(new_n1332), .Y(new_n1333));
  nand_5 g1018(.A(new_n1333), .B(new_n404), .Y(new_n1334));
  xor_4  g1019(.A(new_n1334), .B(new_n406), .Y(po068));
  xor_4  g1020(.A(new_n523), .B(new_n444), .Y(po069));
  xor_4  g1021(.A(new_n1135), .B(new_n325), .Y(new_n1337));
  xor_4  g1022(.A(new_n333), .B(new_n330), .Y(new_n1338));
  nor_5  g1023(.A(new_n323), .B(pi050), .Y(new_n1339));
  nand_5 g1024(.A(new_n1053), .B(new_n329), .Y(new_n1340));
  or_6   g1025(.A(new_n1340), .B(new_n1339), .Y(new_n1341));
  nand_5 g1026(.A(new_n1340), .B(new_n324), .Y(new_n1342));
  nand_5 g1027(.A(new_n1342), .B(new_n1341), .Y(new_n1343));
  xor_4  g1028(.A(new_n1343), .B(new_n1338), .Y(new_n1344));
  nand_5 g1029(.A(new_n1344), .B(new_n540), .Y(new_n1345));
  nand_5 g1030(.A(new_n333), .B(new_n330), .Y(new_n1346));
  nand_5 g1031(.A(new_n1346), .B(new_n329), .Y(new_n1347));
  or_6   g1032(.A(new_n1347), .B(new_n1339), .Y(new_n1348));
  nand_5 g1033(.A(new_n1347), .B(new_n324), .Y(new_n1349));
  nand_5 g1034(.A(new_n1349), .B(new_n1348), .Y(new_n1350));
  xor_4  g1035(.A(new_n335), .B(new_n330), .Y(new_n1351));
  xor_4  g1036(.A(new_n1351), .B(new_n1350), .Y(new_n1352));
  or_6   g1037(.A(new_n1352), .B(new_n540), .Y(new_n1353));
  nand_5 g1038(.A(new_n1353), .B(new_n1345), .Y(new_n1354));
  xor_4  g1039(.A(new_n1354), .B(new_n321), .Y(new_n1355));
  nand_5 g1040(.A(new_n374), .B(new_n363), .Y(new_n1356));
  nand_5 g1041(.A(new_n1356), .B(new_n1069), .Y(new_n1357));
  xor_4  g1042(.A(new_n373), .B(new_n365), .Y(new_n1358));
  xor_4  g1043(.A(new_n370), .B(new_n368), .Y(new_n1359));
  xor_4  g1044(.A(new_n1359), .B(new_n367), .Y(new_n1360));
  xor_4  g1045(.A(new_n1360), .B(new_n1358), .Y(new_n1361));
  not_8  g1046(.A(new_n1361), .Y(new_n1362));
  or_6   g1047(.A(new_n1362), .B(new_n375), .Y(new_n1363));
  nand_5 g1048(.A(new_n1363), .B(new_n376), .Y(new_n1364));
  xor_4  g1049(.A(new_n1364), .B(new_n1357), .Y(new_n1365));
  nand_5 g1050(.A(new_n1365), .B(new_n1136), .Y(new_n1366));
  xor_4  g1051(.A(new_n1362), .B(new_n363), .Y(new_n1367));
  nand_5 g1052(.A(new_n1367), .B(new_n536), .Y(new_n1368));
  nand_5 g1053(.A(new_n1368), .B(new_n1366), .Y(new_n1369));
  xor_4  g1054(.A(new_n1369), .B(new_n901), .Y(new_n1370));
  xor_4  g1055(.A(new_n1370), .B(new_n1355), .Y(new_n1371));
  xor_4  g1056(.A(new_n1371), .B(new_n1337), .Y(po070));
  xor_4  g1057(.A(new_n519), .B(new_n456), .Y(po073));
  xor_4  g1058(.A(new_n999), .B(new_n923), .Y(po083));
  not_8  g1059(.A(new_n736), .Y(po084));
  not_8  g1060(.A(new_n1197), .Y(po086));
  nand_5 g1061(.A(new_n1035), .B(new_n996), .Y(new_n1377));
  xor_4  g1062(.A(new_n1377), .B(new_n1046), .Y(po091));
  xor_4  g1063(.A(new_n509), .B(new_n944), .Y(po092));
  nand_5 g1064(.A(new_n1324), .B(new_n517), .Y(new_n1380));
  nand_5 g1065(.A(new_n1380), .B(new_n467), .Y(new_n1381));
  xor_4  g1066(.A(new_n1381), .B(new_n980), .Y(po094));
  xor_4  g1067(.A(new_n536), .B(new_n374), .Y(po095));
  xnor_4 g1068(.A(new_n515), .B(new_n476), .Y(po102));
  nand_5 g1069(.A(new_n532), .B(new_n401), .Y(new_n1385));
  xor_4  g1070(.A(new_n1385), .B(new_n1112), .Y(po104));
  buf_8  g1071(.A(pi050), .Y(po001));
  buf_8  g1072(.A(pi118), .Y(po002));
  buf_8  g1073(.A(pi020), .Y(po004));
  buf_8  g1074(.A(pi196), .Y(po007));
  buf_8  g1075(.A(pi107), .Y(po010));
  buf_8  g1076(.A(pi060), .Y(po012));
  buf_8  g1077(.A(pi108), .Y(po014));
  buf_8  g1078(.A(pi057), .Y(po018));
  buf_8  g1079(.A(pi047), .Y(po019));
  buf_8  g1080(.A(pi085), .Y(po021));
  buf_8  g1081(.A(pi180), .Y(po022));
  buf_8  g1082(.A(po003), .Y(po023));
  buf_8  g1083(.A(pi056), .Y(po028));
  buf_8  g1084(.A(po008), .Y(po031));
  buf_8  g1085(.A(pi001), .Y(po032));
  buf_8  g1086(.A(pi204), .Y(po033));
  buf_8  g1087(.A(pi039), .Y(po034));
  buf_8  g1088(.A(pi024), .Y(po035));
  buf_8  g1089(.A(pi101), .Y(po036));
  buf_8  g1090(.A(pi144), .Y(po037));
  buf_8  g1091(.A(po040), .Y(po041));
  buf_8  g1092(.A(pi160), .Y(po042));
  buf_8  g1093(.A(pi060), .Y(po045));
  buf_8  g1094(.A(pi162), .Y(po046));
  buf_8  g1095(.A(po017), .Y(po051));
  buf_8  g1096(.A(pi122), .Y(po052));
  buf_8  g1097(.A(pi027), .Y(po053));
  buf_8  g1098(.A(pi051), .Y(po055));
  buf_8  g1099(.A(pi147), .Y(po056));
  buf_8  g1100(.A(pi183), .Y(po063));
  buf_8  g1101(.A(pi192), .Y(po064));
  buf_8  g1102(.A(pi064), .Y(po071));
  buf_8  g1103(.A(po040), .Y(po072));
  buf_8  g1104(.A(pi132), .Y(po074));
  buf_8  g1105(.A(po008), .Y(po075));
  buf_8  g1106(.A(pi181), .Y(po076));
  buf_8  g1107(.A(pi083), .Y(po077));
  buf_8  g1108(.A(po065), .Y(po078));
  buf_8  g1109(.A(pi170), .Y(po079));
  buf_8  g1110(.A(pi199), .Y(po081));
  buf_8  g1111(.A(po017), .Y(po082));
  buf_8  g1112(.A(pi153), .Y(po085));
  buf_8  g1113(.A(pi137), .Y(po087));
  buf_8  g1114(.A(po030), .Y(po088));
  buf_8  g1115(.A(pi060), .Y(po089));
  buf_8  g1116(.A(pi092), .Y(po093));
  buf_8  g1117(.A(pi116), .Y(po096));
  buf_8  g1118(.A(pi060), .Y(po097));
  buf_8  g1119(.A(pi074), .Y(po098));
  buf_8  g1120(.A(po029), .Y(po099));
  buf_8  g1121(.A(po040), .Y(po101));
  buf_8  g1122(.A(pi178), .Y(po103));
  buf_8  g1123(.A(pi018), .Y(po105));
  buf_8  g1124(.A(pi004), .Y(po106));
endmodule


