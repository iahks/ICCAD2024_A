// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Mon Jul 15 23:49:29 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604,
    n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112,
    n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288,
    n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558,
    n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738,
    n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088,
    n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272,
    n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479,
    n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816,
    n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136,
    n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349,
    n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618,
    n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952,
    n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319,
    n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722,
    n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031,
    n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213,
    n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443,
    n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822,
    n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379,
    n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590,
    n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790,
    n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305,
    n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566,
    n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731,
    n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963,
    n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305,
    n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614,
    n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827,
    n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251,
    n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493,
    n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926,
    n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117,
    n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514,
    n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763,
    n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220,
    n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479,
    n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667,
    n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121,
    n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398,
    n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650,
    n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900,
    n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263,
    n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494,
    n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783,
    n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230,
    n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603,
    n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899,
    n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271,
    n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546,
    n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918,
    n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247,
    n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524,
    n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968,
    n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095,
    n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954,
    n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227,
    n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496,
    n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880,
    n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107,
    n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327,
    n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531,
    n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770,
    n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040,
    n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259,
    n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478,
    n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946,
    n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287,
    n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674,
    n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898,
    n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068,
    n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309,
    n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492,
    n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764,
    n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068,
    n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333,
    n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657,
    n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912,
    n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129,
    n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485,
    n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023,
    n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240,
    n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435,
    n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643,
    n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926,
    n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191,
    n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512,
    n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752,
    n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089,
    n27104, n27120, n27134, n27188,
    n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194  );
  input  n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583,
    n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099,
    n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279,
    n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536,
    n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689,
    n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035,
    n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210,
    n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421,
    n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809,
    n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030,
    n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324,
    n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582,
    n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945,
    n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306,
    n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665,
    n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026,
    n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211,
    n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438,
    n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752,
    n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369,
    n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556,
    n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785,
    n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149,
    n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524,
    n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721,
    n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949,
    n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285,
    n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581,
    n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806,
    n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246,
    n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460,
    n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872,
    n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096,
    n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411,
    n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739,
    n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201,
    n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473,
    n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630,
    n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113,
    n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384,
    n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626,
    n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892,
    n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190,
    n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490,
    n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781,
    n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148,
    n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576,
    n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826,
    n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258,
    n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539,
    n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884,
    n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223,
    n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521,
    n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911,
    n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090,
    n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911,
    n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171,
    n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483,
    n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745,
    n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081,
    n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282,
    n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515,
    n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701,
    n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036,
    n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250,
    n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470,
    n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929,
    n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276,
    n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654,
    n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839,
    n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043,
    n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290,
    n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470,
    n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660,
    n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065,
    n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304,
    n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586,
    n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895,
    n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093,
    n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374,
    n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937,
    n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168,
    n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381,
    n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629,
    n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923,
    n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180,
    n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510,
    n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748,
    n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037,
    n27089, n27104, n27120, n27134, n27188;
  output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355_1, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361_1, new_n2362, new_n2363_1, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374_1, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387_1, new_n2388_1, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409_1, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416_1, new_n2417, new_n2418, new_n2419, new_n2420_1,
    new_n2421_1, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440_1, new_n2441, new_n2442, new_n2443, new_n2444_1,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479_1, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513_1, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533_1, new_n2534,
    new_n2535_1, new_n2536, new_n2537_1, new_n2538, new_n2539, new_n2540,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2548,
    new_n2549, new_n2550, new_n2551, new_n2552, new_n2554, new_n2555_1,
    new_n2556, new_n2557, new_n2558, new_n2559, new_n2560_1, new_n2561_1,
    new_n2562, new_n2563, new_n2564, new_n2565, new_n2566, new_n2567,
    new_n2568, new_n2569, new_n2570_1, new_n2571, new_n2572, new_n2573_1,
    new_n2574, new_n2575, new_n2576, new_n2577, new_n2578_1, new_n2579,
    new_n2580, new_n2581, new_n2582_1, new_n2583, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602_1, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619_1, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646_1, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659_1, new_n2660, new_n2661_1, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680_1, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693_1,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703_1, new_n2704, new_n2705,
    new_n2706_1, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711_1,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731_1, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743_1, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761_1, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774_1, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779_1, new_n2780, new_n2781, new_n2782, new_n2783_1,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809_1, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816_1, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826_1, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853_1, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858_1, new_n2859, new_n2860_1, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886_1,
    new_n2887_1, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929_1, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944_1, new_n2945, new_n2946,
    new_n2947, new_n2948_1, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961_1, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971_1, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978_1, new_n2979_1, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985_1, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999_1, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010_1, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017_1, new_n3018_1,
    new_n3019, new_n3020_1, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030_1,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067_1, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076_1, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3086, new_n3087, new_n3088, new_n3089_1, new_n3090, new_n3091,
    new_n3092, new_n3093, new_n3094, new_n3095, new_n3096, new_n3097,
    new_n3098, new_n3099, new_n3100, new_n3101, new_n3102, new_n3103,
    new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125_1, new_n3126_1, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136_1, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161_1, new_n3162, new_n3163,
    new_n3164_1, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208_1, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219_1, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228_1, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235_1,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244_1, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253_1,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260_1, new_n3261, new_n3262, new_n3263_1, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279_1, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289_1,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301_1,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306_1, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316_1, new_n3317, new_n3318, new_n3319,
    new_n3320_1, new_n3321, new_n3322, new_n3323, new_n3324_1, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332_1, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343_1,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349_1,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366_1, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390_1, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425_1, new_n3426_1, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451_1, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459_1, new_n3460_1, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468_1, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480_1, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502_1, new_n3503, new_n3504, new_n3505, new_n3506_1,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516_1, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528_1, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541_1, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555_1, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561_1, new_n3562, new_n3563_1, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570_1, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582_1, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617_1, new_n3618_1, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642_1, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649_1, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665_1, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679_1, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710_1,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3725_1, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733_1, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740_1, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755_1, new_n3756, new_n3757, new_n3758_1, new_n3759,
    new_n3760_1, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781_1, new_n3782, new_n3783,
    new_n3784, new_n3785_1, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794_1, new_n3795_1,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828_1, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850_1, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869_1, new_n3870, new_n3871_1, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891_1,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909_1,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918_1, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925_1, new_n3926, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933, new_n3934_1,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945_1, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952_1,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959_1, new_n3960, new_n3961, new_n3962_1, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971_1, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983_1, new_n3984_1, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000_1,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010_1, new_n4011, new_n4012,
    new_n4013, new_n4014_1, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071_1, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085_1, new_n4086, new_n4087, new_n4088_1, new_n4089_1, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100_1, new_n4101, new_n4102,
    new_n4103_1, new_n4104, new_n4106, new_n4107, new_n4108, new_n4109,
    new_n4110, new_n4111, new_n4112, new_n4113, new_n4114, new_n4115,
    new_n4116, new_n4117, new_n4118, new_n4119_1, new_n4120, new_n4121,
    new_n4122, new_n4123_1, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134_1, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146_1, new_n4147, new_n4148, new_n4149, new_n4150_1, new_n4151_1,
    new_n4152_1, new_n4153_1, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4165_1, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172_1, new_n4173_1, new_n4174, new_n4175, new_n4176_1,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186_1, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204_1, new_n4205_1, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215_1, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221_1, new_n4222, new_n4223, new_n4224_1,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231_1, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256_1, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266_1,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272_1,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306_1, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4312, new_n4313, new_n4314, new_n4315,
    new_n4316, new_n4317, new_n4318, new_n4319_1, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325_1, new_n4326_1, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340_1, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374_1, new_n4375,
    new_n4376_1, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401_1, new_n4402, new_n4403, new_n4404, new_n4405,
    new_n4406, new_n4407, new_n4408, new_n4409_1, new_n4410, new_n4411,
    new_n4412, new_n4413, new_n4414, new_n4415, new_n4416, new_n4417,
    new_n4418, new_n4419, new_n4420, new_n4421, new_n4422, new_n4423,
    new_n4424_1, new_n4425, new_n4426_1, new_n4427, new_n4428, new_n4429,
    new_n4430, new_n4431, new_n4432_1, new_n4433, new_n4434, new_n4435,
    new_n4436, new_n4437, new_n4438, new_n4439, new_n4440, new_n4441_1,
    new_n4442, new_n4443, new_n4444, new_n4445, new_n4446, new_n4447,
    new_n4448, new_n4449, new_n4450, new_n4451_1, new_n4452, new_n4453,
    new_n4454, new_n4455, new_n4456, new_n4457, new_n4458, new_n4459,
    new_n4460, new_n4461, new_n4462, new_n4463, new_n4464, new_n4465,
    new_n4466, new_n4467, new_n4468, new_n4469, new_n4470, new_n4471,
    new_n4472, new_n4473, new_n4474, new_n4475, new_n4476_1, new_n4477,
    new_n4478_1, new_n4479, new_n4480, new_n4481, new_n4482, new_n4483,
    new_n4484, new_n4485, new_n4486, new_n4487, new_n4488, new_n4489,
    new_n4490, new_n4491, new_n4492, new_n4493, new_n4494, new_n4495,
    new_n4496, new_n4497, new_n4498, new_n4499, new_n4500, new_n4501,
    new_n4502, new_n4503, new_n4504, new_n4505, new_n4506, new_n4507,
    new_n4508, new_n4509, new_n4510, new_n4511, new_n4512, new_n4513,
    new_n4514_1, new_n4515, new_n4516, new_n4517, new_n4518, new_n4519,
    new_n4520, new_n4521, new_n4522, new_n4523, new_n4524, new_n4525,
    new_n4526, new_n4527, new_n4528, new_n4529_1, new_n4530, new_n4531,
    new_n4532, new_n4533, new_n4534, new_n4535, new_n4536, new_n4537,
    new_n4538, new_n4539, new_n4540, new_n4541, new_n4542, new_n4543,
    new_n4544, new_n4545, new_n4546, new_n4547, new_n4548, new_n4549,
    new_n4550, new_n4551, new_n4552_1, new_n4553, new_n4554, new_n4555,
    new_n4556, new_n4557, new_n4558, new_n4559, new_n4560, new_n4561,
    new_n4562, new_n4563, new_n4564, new_n4565, new_n4566, new_n4567,
    new_n4568, new_n4569, new_n4570, new_n4571, new_n4572, new_n4573,
    new_n4574, new_n4575, new_n4576, new_n4577, new_n4578, new_n4579,
    new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585,
    new_n4586, new_n4587, new_n4588_1, new_n4589, new_n4590_1, new_n4591,
    new_n4592, new_n4593, new_n4594, new_n4595_1, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4611, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624_1, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646_1,
    new_n4647, new_n4648, new_n4649, new_n4650, new_n4651, new_n4652,
    new_n4653, new_n4654, new_n4655, new_n4656, new_n4657, new_n4658,
    new_n4659, new_n4660, new_n4661, new_n4662, new_n4663, new_n4664,
    new_n4665_1, new_n4666, new_n4667, new_n4668, new_n4669, new_n4670,
    new_n4671, new_n4672, new_n4673, new_n4674_1, new_n4675, new_n4676,
    new_n4677, new_n4678, new_n4679, new_n4680, new_n4681, new_n4682,
    new_n4683, new_n4684, new_n4685, new_n4686, new_n4687, new_n4688,
    new_n4689, new_n4690, new_n4691, new_n4692, new_n4693_1, new_n4694,
    new_n4695, new_n4696, new_n4697, new_n4698, new_n4699, new_n4700,
    new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706,
    new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712,
    new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718,
    new_n4719, new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731_1, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745_1, new_n4746, new_n4747_1, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755, new_n4756, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766_1, new_n4767,
    new_n4768, new_n4769, new_n4770_1, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777_1, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785_1,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804_1, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810_1, new_n4811, new_n4812_1, new_n4813, new_n4814_1, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850_1, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858_1, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891_1, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913_1, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921, new_n4922, new_n4923,
    new_n4924, new_n4925_1, new_n4926, new_n4927, new_n4928, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938, new_n4939_1, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947_1,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952_1, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957_1, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964_1, new_n4965,
    new_n4966_1, new_n4967_1, new_n4968, new_n4969, new_n4970, new_n4971,
    new_n4972_1, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011_1, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020_1, new_n5021, new_n5022, new_n5023, new_n5024_1, new_n5025_1,
    new_n5026_1, new_n5027, new_n5028, new_n5030, new_n5031_1, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046_1, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060_1, new_n5061, new_n5062_1,
    new_n5063, new_n5064_1, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077_1, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082_1, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5090, new_n5091, new_n5092, new_n5093,
    new_n5094, new_n5095, new_n5096, new_n5097, new_n5098_1, new_n5099,
    new_n5100, new_n5101_1, new_n5102, new_n5103, new_n5104, new_n5105,
    new_n5106, new_n5107, new_n5108, new_n5109, new_n5110, new_n5111,
    new_n5112, new_n5113, new_n5114, new_n5115_1, new_n5116, new_n5117,
    new_n5118, new_n5119, new_n5120_1, new_n5121, new_n5122, new_n5123,
    new_n5124, new_n5125, new_n5126, new_n5127, new_n5128_1, new_n5129,
    new_n5130, new_n5131_1, new_n5132, new_n5133, new_n5134, new_n5135,
    new_n5136, new_n5137, new_n5138, new_n5139, new_n5140_1, new_n5141,
    new_n5142, new_n5143, new_n5144, new_n5145, new_n5146, new_n5147,
    new_n5148, new_n5149, new_n5150, new_n5151, new_n5152, new_n5153,
    new_n5154, new_n5155, new_n5156, new_n5157, new_n5158_1, new_n5159,
    new_n5160, new_n5161, new_n5162, new_n5163, new_n5164, new_n5165,
    new_n5166, new_n5167, new_n5168_1, new_n5169, new_n5170, new_n5171,
    new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177,
    new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183,
    new_n5184_1, new_n5185, new_n5186, new_n5187, new_n5188, new_n5189,
    new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195,
    new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201,
    new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207,
    new_n5208, new_n5209, new_n5210, new_n5211_1, new_n5212, new_n5213_1,
    new_n5214, new_n5215, new_n5216, new_n5217, new_n5219, new_n5220,
    new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226_1,
    new_n5227, new_n5228_1, new_n5229, new_n5230, new_n5231, new_n5232,
    new_n5233, new_n5234, new_n5235, new_n5236, new_n5237, new_n5238,
    new_n5239, new_n5240, new_n5241, new_n5242, new_n5243, new_n5244,
    new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255_1, new_n5256_1,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265_1, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273_1, new_n5274_1,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300_1, new_n5301, new_n5302_1, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310,
    new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316,
    new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322,
    new_n5323, new_n5324, new_n5325_1, new_n5326, new_n5327, new_n5328,
    new_n5329, new_n5330_1, new_n5331, new_n5332, new_n5333, new_n5334,
    new_n5335, new_n5336, new_n5337_1, new_n5338, new_n5339, new_n5340,
    new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346,
    new_n5347, new_n5348, new_n5349, new_n5350, new_n5351_1, new_n5352,
    new_n5353_1, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358,
    new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376_1,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386_1, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399_1, new_n5400_1,
    new_n5401, new_n5402, new_n5403_1, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430_1,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438_1, new_n5439_1, new_n5440, new_n5441, new_n5442,
    new_n5443_1, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451_1, new_n5453, new_n5454, new_n5455,
    new_n5456, new_n5457, new_n5458, new_n5459, new_n5460, new_n5461,
    new_n5462, new_n5463, new_n5464, new_n5465, new_n5466, new_n5467,
    new_n5468, new_n5469, new_n5470, new_n5471, new_n5472_1, new_n5473,
    new_n5474, new_n5475, new_n5476, new_n5477, new_n5478, new_n5479,
    new_n5480, new_n5481, new_n5482, new_n5483, new_n5484, new_n5485_1,
    new_n5486, new_n5487, new_n5488, new_n5489, new_n5490, new_n5491,
    new_n5492, new_n5493, new_n5494, new_n5495, new_n5496, new_n5497,
    new_n5498, new_n5499, new_n5500, new_n5501, new_n5502, new_n5503,
    new_n5504, new_n5505, new_n5506, new_n5507, new_n5508, new_n5509,
    new_n5510, new_n5511, new_n5512, new_n5513, new_n5514, new_n5515,
    new_n5516, new_n5517_1, new_n5518, new_n5519, new_n5520, new_n5521_1,
    new_n5522, new_n5523, new_n5524_1, new_n5525, new_n5526, new_n5527,
    new_n5528, new_n5529, new_n5530, new_n5531, new_n5532_1, new_n5533,
    new_n5534, new_n5535, new_n5536, new_n5537, new_n5538, new_n5539,
    new_n5540, new_n5541, new_n5542, new_n5543, new_n5544, new_n5545,
    new_n5546, new_n5547, new_n5548, new_n5549, new_n5550, new_n5551,
    new_n5552, new_n5553, new_n5554, new_n5555, new_n5556, new_n5557,
    new_n5558, new_n5559, new_n5560, new_n5561, new_n5562, new_n5563,
    new_n5564_1, new_n5565, new_n5566, new_n5567, new_n5568, new_n5569,
    new_n5570, new_n5571, new_n5572, new_n5573, new_n5574, new_n5575,
    new_n5576, new_n5577, new_n5578, new_n5579_1, new_n5580, new_n5581,
    new_n5582, new_n5583, new_n5584, new_n5585, new_n5586, new_n5587,
    new_n5588, new_n5589, new_n5590, new_n5591, new_n5592, new_n5593_1,
    new_n5594, new_n5595, new_n5596, new_n5597, new_n5598, new_n5599,
    new_n5600, new_n5601, new_n5602, new_n5603_1, new_n5604, new_n5605_1,
    new_n5606, new_n5607, new_n5608, new_n5609_1, new_n5610, new_n5611,
    new_n5612, new_n5613, new_n5614, new_n5615, new_n5616, new_n5617,
    new_n5618, new_n5619, new_n5620, new_n5621, new_n5622, new_n5623,
    new_n5624, new_n5625, new_n5626, new_n5627, new_n5628, new_n5629,
    new_n5630, new_n5631, new_n5632, new_n5633, new_n5634_1, new_n5635,
    new_n5636, new_n5637, new_n5638, new_n5639, new_n5640, new_n5641,
    new_n5642, new_n5643_1, new_n5644, new_n5645, new_n5646, new_n5647,
    new_n5648, new_n5649, new_n5650, new_n5651, new_n5652, new_n5653,
    new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659,
    new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665,
    new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671,
    new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677,
    new_n5678, new_n5679, new_n5680_1, new_n5681, new_n5682, new_n5683,
    new_n5684, new_n5685, new_n5686, new_n5687_1, new_n5688, new_n5689,
    new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695,
    new_n5696_1, new_n5697, new_n5698, new_n5699, new_n5700_1, new_n5701,
    new_n5702, new_n5703, new_n5704_1, new_n5705, new_n5706, new_n5707,
    new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713,
    new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719,
    new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725,
    new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731,
    new_n5732_1, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5742_1, new_n5743,
    new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749,
    new_n5750, new_n5751, new_n5752_1, new_n5753, new_n5754, new_n5755,
    new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761,
    new_n5762, new_n5763, new_n5764, new_n5765_1, new_n5766, new_n5767,
    new_n5769, new_n5770, new_n5771, new_n5772, new_n5773, new_n5774,
    new_n5775, new_n5776_1, new_n5777, new_n5778, new_n5779, new_n5780,
    new_n5781, new_n5782_1, new_n5783, new_n5784, new_n5785, new_n5786,
    new_n5787, new_n5788, new_n5789, new_n5790, new_n5792, new_n5793,
    new_n5794, new_n5795, new_n5798, new_n5799, new_n5800, new_n5801,
    new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807,
    new_n5808, new_n5809, new_n5810, new_n5811, new_n5812, new_n5813,
    new_n5814, new_n5815, new_n5816, new_n5817, new_n5818, new_n5819,
    new_n5820, new_n5821, new_n5822_1, new_n5823, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833_1, new_n5834_1, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840_1, new_n5841_1, new_n5842_1, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850_1,
    new_n5851, new_n5853, new_n5856, new_n5857, new_n5858, new_n5859,
    new_n5860, new_n5861, new_n5862, new_n5863, new_n5864, new_n5865,
    new_n5866, new_n5867, new_n5868, new_n5869, new_n5870, new_n5871,
    new_n5872, new_n5873, new_n5874, new_n5875, new_n5876, new_n5877,
    new_n5878, new_n5879, new_n5880, new_n5881, new_n5882_1, new_n5883,
    new_n5884, new_n5885, new_n5886, new_n5887, new_n5888, new_n5889,
    new_n5890, new_n5891, new_n5892, new_n5893, new_n5894, new_n5895,
    new_n5896, new_n5897, new_n5898, new_n5899, new_n5900, new_n5901,
    new_n5902, new_n5903_1, new_n5904_1, new_n5905, new_n5906, new_n5907,
    new_n5908, new_n5909, new_n5910, new_n5911_1, new_n5912, new_n5913,
    new_n5914, new_n5915, new_n5916, new_n5917, new_n5918, new_n5919,
    new_n5920, new_n5921, new_n5922, new_n5923, new_n5924, new_n5925,
    new_n5926, new_n5927, new_n5928, new_n5929, new_n5930, new_n5931,
    new_n5932, new_n5933, new_n5934, new_n5935, new_n5936_1, new_n5937,
    new_n5938, new_n5939, new_n5940, new_n5941, new_n5942, new_n5943_1,
    new_n5944, new_n5945, new_n5946, new_n5947, new_n5948, new_n5949,
    new_n5950, new_n5951, new_n5952, new_n5953, new_n5954, new_n5955,
    new_n5956, new_n5957, new_n5958, new_n5959, new_n5960, new_n5961,
    new_n5962, new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967,
    new_n5968, new_n5969, new_n5970, new_n5971, new_n5972, new_n5973,
    new_n5974, new_n5975, new_n5976, new_n5977, new_n5978, new_n5979,
    new_n5980_1, new_n5981, new_n5982, new_n5983, new_n5984, new_n5985,
    new_n5986, new_n5987, new_n5988, new_n5989, new_n5990, new_n5991,
    new_n5992, new_n5993, new_n5994, new_n5995, new_n5996, new_n5997,
    new_n5998, new_n5999, new_n6000, new_n6001, new_n6002, new_n6003,
    new_n6004, new_n6005, new_n6006, new_n6007, new_n6008, new_n6009,
    new_n6010, new_n6011, new_n6012_1, new_n6013, new_n6014, new_n6015,
    new_n6016, new_n6017, new_n6018, new_n6019, new_n6020, new_n6021,
    new_n6022_1, new_n6023, new_n6024, new_n6025, new_n6026, new_n6027,
    new_n6028, new_n6029, new_n6030, new_n6031_1, new_n6032, new_n6033,
    new_n6034, new_n6035, new_n6036, new_n6037, new_n6038, new_n6039,
    new_n6040, new_n6041, new_n6042, new_n6043, new_n6044_1, new_n6045,
    new_n6046_1, new_n6047, new_n6048, new_n6049, new_n6050, new_n6051,
    new_n6052, new_n6053, new_n6054, new_n6055, new_n6056, new_n6057,
    new_n6058, new_n6059, new_n6060, new_n6061, new_n6062, new_n6063,
    new_n6064, new_n6065, new_n6066, new_n6067, new_n6068, new_n6069,
    new_n6070, new_n6071, new_n6072, new_n6073, new_n6074, new_n6075,
    new_n6076, new_n6077, new_n6078, new_n6079, new_n6080, new_n6081,
    new_n6082, new_n6083, new_n6084_1, new_n6085, new_n6086, new_n6087,
    new_n6088, new_n6089, new_n6090, new_n6091, new_n6092, new_n6093,
    new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099,
    new_n6100, new_n6101, new_n6102, new_n6103, new_n6104_1, new_n6105_1,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123,
    new_n6124, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6151, new_n6152, new_n6153, new_n6154,
    new_n6155, new_n6156, new_n6157, new_n6158, new_n6159, new_n6160_1,
    new_n6161, new_n6162, new_n6163, new_n6164, new_n6165, new_n6166,
    new_n6167, new_n6168, new_n6169, new_n6170, new_n6171_1, new_n6172,
    new_n6173, new_n6174, new_n6175, new_n6176, new_n6177, new_n6178,
    new_n6179, new_n6180, new_n6181, new_n6182, new_n6183_1, new_n6184,
    new_n6185, new_n6186, new_n6187, new_n6188, new_n6189_1, new_n6190,
    new_n6191, new_n6192, new_n6193, new_n6194, new_n6195, new_n6196,
    new_n6197, new_n6198, new_n6199, new_n6200, new_n6201, new_n6202,
    new_n6203, new_n6204_1, new_n6205, new_n6206, new_n6207, new_n6208,
    new_n6209, new_n6210, new_n6211, new_n6212, new_n6213, new_n6214,
    new_n6215, new_n6216, new_n6217, new_n6218_1, new_n6219, new_n6220,
    new_n6221, new_n6222, new_n6223_1, new_n6224, new_n6225, new_n6226,
    new_n6227, new_n6228, new_n6229, new_n6230, new_n6231, new_n6232,
    new_n6233_1, new_n6234, new_n6235, new_n6236, new_n6237, new_n6238,
    new_n6239, new_n6240, new_n6241, new_n6242, new_n6243, new_n6244,
    new_n6245_1, new_n6246, new_n6247, new_n6248_1, new_n6249, new_n6250,
    new_n6251, new_n6252, new_n6253, new_n6254, new_n6255, new_n6256_1,
    new_n6257, new_n6258, new_n6259, new_n6260, new_n6261, new_n6262,
    new_n6263, new_n6264, new_n6265, new_n6266, new_n6267, new_n6268,
    new_n6269, new_n6270, new_n6271_1, new_n6272, new_n6273, new_n6274,
    new_n6275, new_n6276_1, new_n6277, new_n6278, new_n6279, new_n6280,
    new_n6281, new_n6282, new_n6283, new_n6284, new_n6285, new_n6286,
    new_n6287, new_n6288, new_n6289, new_n6290, new_n6291, new_n6292,
    new_n6293, new_n6294, new_n6295, new_n6296, new_n6297, new_n6298,
    new_n6299, new_n6300, new_n6301, new_n6302, new_n6303, new_n6304,
    new_n6305, new_n6306, new_n6307, new_n6308_1, new_n6309, new_n6310,
    new_n6311_1, new_n6312, new_n6313, new_n6314, new_n6315, new_n6316,
    new_n6317, new_n6318, new_n6319, new_n6320, new_n6321, new_n6322,
    new_n6323_1, new_n6324, new_n6325, new_n6326, new_n6327, new_n6328,
    new_n6329, new_n6330_1, new_n6331, new_n6332, new_n6333, new_n6334,
    new_n6335, new_n6336, new_n6337, new_n6338, new_n6339_1, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354_1, new_n6355, new_n6356_1, new_n6357, new_n6358,
    new_n6359, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364,
    new_n6365, new_n6366, new_n6367, new_n6368, new_n6369_1, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375_1, new_n6376,
    new_n6377, new_n6378, new_n6379_1, new_n6380, new_n6381_1, new_n6382,
    new_n6383_1, new_n6384, new_n6385_1, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397_1, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407_1, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6425,
    new_n6426, new_n6427_1, new_n6428, new_n6429, new_n6430, new_n6431_1,
    new_n6432, new_n6433, new_n6434, new_n6435, new_n6436, new_n6437_1,
    new_n6438, new_n6439, new_n6440, new_n6441, new_n6442, new_n6443,
    new_n6444, new_n6445, new_n6446, new_n6447, new_n6448, new_n6449,
    new_n6450, new_n6451, new_n6452, new_n6453, new_n6454, new_n6455,
    new_n6456_1, new_n6457_1, new_n6458, new_n6459, new_n6460, new_n6461,
    new_n6462, new_n6463, new_n6464, new_n6465_1, new_n6466, new_n6467,
    new_n6468, new_n6469, new_n6470_1, new_n6471, new_n6472, new_n6473,
    new_n6474, new_n6475, new_n6476_1, new_n6477, new_n6478, new_n6479,
    new_n6480, new_n6481, new_n6482, new_n6483, new_n6484, new_n6485_1,
    new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491,
    new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497,
    new_n6498, new_n6499, new_n6500, new_n6501, new_n6502_1, new_n6503,
    new_n6504, new_n6505, new_n6506_1, new_n6507, new_n6508, new_n6509,
    new_n6510, new_n6511, new_n6512, new_n6513_1, new_n6514_1, new_n6515,
    new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521,
    new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542_1, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556_1, new_n6557,
    new_n6558_1, new_n6559, new_n6560_1, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567_1, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576_1, new_n6577, new_n6578, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6585, new_n6586, new_n6587_1, new_n6589,
    new_n6590_1, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595,
    new_n6596_1, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601,
    new_n6602, new_n6603, new_n6604, new_n6605, new_n6606, new_n6607,
    new_n6608, new_n6609, new_n6610, new_n6611_1, new_n6612_1, new_n6613,
    new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619,
    new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6625,
    new_n6626, new_n6627, new_n6628_1, new_n6629, new_n6630_1, new_n6631_1,
    new_n6632, new_n6633, new_n6634_1, new_n6635, new_n6636, new_n6637,
    new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643,
    new_n6644, new_n6645, new_n6646, new_n6647, new_n6648, new_n6649,
    new_n6650, new_n6651, new_n6652_1, new_n6653, new_n6654, new_n6655_1,
    new_n6656, new_n6657, new_n6658, new_n6659_1, new_n6660, new_n6661,
    new_n6662, new_n6663, new_n6664, new_n6665, new_n6666, new_n6667,
    new_n6668, new_n6669_1, new_n6670, new_n6671_1, new_n6672, new_n6673_1,
    new_n6675, new_n6676, new_n6677, new_n6678, new_n6679, new_n6680,
    new_n6681, new_n6682, new_n6683, new_n6684_1, new_n6685, new_n6686,
    new_n6687, new_n6688, new_n6689, new_n6690, new_n6691_1, new_n6692,
    new_n6693, new_n6694, new_n6695, new_n6696, new_n6697, new_n6698,
    new_n6699, new_n6700, new_n6701, new_n6702, new_n6703, new_n6704,
    new_n6705, new_n6706_1, new_n6707_1, new_n6708, new_n6709, new_n6710,
    new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716,
    new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722,
    new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728,
    new_n6729_1, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734,
    new_n6735, new_n6736_1, new_n6737, new_n6738, new_n6739, new_n6740,
    new_n6741, new_n6742, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6772, new_n6773_1, new_n6774, new_n6775_1, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785_1, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790_1, new_n6791_1, new_n6792, new_n6793, new_n6794_1, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802_1, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814_1, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826_1, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835_1, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853_1, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861_1,
    new_n6862_1, new_n6863_1, new_n6864, new_n6865, new_n6866, new_n6867_1,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6966, new_n6967_1, new_n6968, new_n6969, new_n6970,
    new_n6971_1, new_n6972, new_n6973, new_n6974, new_n6975_1, new_n6976,
    new_n6977, new_n6978, new_n6979, new_n6980, new_n6981, new_n6982,
    new_n6983_1, new_n6984, new_n6985_1, new_n6986, new_n6987, new_n6988,
    new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994,
    new_n6995, new_n6996, new_n6997, new_n6998_1, new_n6999, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026_1, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032_1, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038_1, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054,
    new_n7055, new_n7056, new_n7057_1, new_n7058, new_n7059, new_n7060,
    new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066,
    new_n7067, new_n7068, new_n7069, new_n7070, new_n7071, new_n7072,
    new_n7073, new_n7074, new_n7075, new_n7076, new_n7077, new_n7078,
    new_n7079_1, new_n7080, new_n7081, new_n7082, new_n7083, new_n7084,
    new_n7085, new_n7086, new_n7087, new_n7088, new_n7089, new_n7090,
    new_n7091, new_n7092, new_n7093, new_n7094, new_n7095, new_n7096,
    new_n7097, new_n7098, new_n7099_1, new_n7100, new_n7101, new_n7102,
    new_n7103, new_n7104, new_n7105, new_n7106, new_n7107, new_n7108,
    new_n7109, new_n7110, new_n7111, new_n7112, new_n7113, new_n7114,
    new_n7115, new_n7116, new_n7117, new_n7118, new_n7119, new_n7120,
    new_n7121, new_n7122, new_n7123, new_n7124, new_n7125, new_n7126,
    new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132,
    new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138,
    new_n7139_1, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144,
    new_n7145, new_n7146, new_n7147, new_n7148, new_n7149_1, new_n7150,
    new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156,
    new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7188, new_n7189, new_n7190_1, new_n7191, new_n7192,
    new_n7193, new_n7194, new_n7195, new_n7196, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229_1, new_n7230_1,
    new_n7231, new_n7232, new_n7233_1, new_n7234, new_n7235, new_n7236_1,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253_1, new_n7254,
    new_n7255, new_n7256_1, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268_1, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277_1, new_n7278,
    new_n7279, new_n7280_1, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298_1, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305_1, new_n7306, new_n7307, new_n7308_1,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313_1, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330_1, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335_1, new_n7336, new_n7337, new_n7338,
    new_n7339_1, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346_1, new_n7347, new_n7348, new_n7349_1, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363_1, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377_1, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390_1, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403_1, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408_1, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421_1, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7429,
    new_n7430, new_n7431, new_n7432_1, new_n7433, new_n7434, new_n7435,
    new_n7436, new_n7437_1, new_n7438, new_n7439, new_n7440, new_n7441,
    new_n7442, new_n7443, new_n7444, new_n7445, new_n7446, new_n7447,
    new_n7448, new_n7449, new_n7450, new_n7451, new_n7452, new_n7453,
    new_n7454, new_n7455, new_n7456, new_n7457, new_n7458, new_n7459,
    new_n7460_1, new_n7461, new_n7462, new_n7463, new_n7464, new_n7465,
    new_n7466, new_n7467, new_n7468, new_n7469, new_n7470, new_n7471,
    new_n7472, new_n7473, new_n7474, new_n7475_1, new_n7476, new_n7477_1,
    new_n7478, new_n7479, new_n7480, new_n7481, new_n7482, new_n7483,
    new_n7484, new_n7485, new_n7486, new_n7487, new_n7488, new_n7489,
    new_n7490, new_n7491, new_n7492, new_n7493, new_n7494, new_n7495,
    new_n7496, new_n7497, new_n7498, new_n7499, new_n7500, new_n7501,
    new_n7502, new_n7503, new_n7504, new_n7505, new_n7506, new_n7507_1,
    new_n7508, new_n7509, new_n7510, new_n7511, new_n7512, new_n7513,
    new_n7514_1, new_n7515, new_n7516, new_n7517, new_n7518, new_n7519,
    new_n7520, new_n7521, new_n7522, new_n7523, new_n7524_1, new_n7525,
    new_n7526, new_n7527, new_n7528, new_n7529, new_n7530, new_n7531,
    new_n7532, new_n7533, new_n7534, new_n7535, new_n7536, new_n7537,
    new_n7538, new_n7539, new_n7540, new_n7541, new_n7542, new_n7543,
    new_n7544, new_n7545, new_n7546, new_n7547, new_n7548, new_n7549,
    new_n7550, new_n7551, new_n7552, new_n7553, new_n7554, new_n7555,
    new_n7556, new_n7557, new_n7558_1, new_n7559, new_n7560, new_n7561,
    new_n7562, new_n7563, new_n7564, new_n7565, new_n7566_1, new_n7567,
    new_n7568, new_n7569_1, new_n7570, new_n7571, new_n7572_1, new_n7573,
    new_n7574, new_n7575_1, new_n7576, new_n7577, new_n7578, new_n7579,
    new_n7580, new_n7581, new_n7582, new_n7583, new_n7584, new_n7585_1,
    new_n7586, new_n7587, new_n7588_1, new_n7589, new_n7590, new_n7591,
    new_n7592, new_n7593_1, new_n7594, new_n7595, new_n7596, new_n7597,
    new_n7598_1, new_n7599, new_n7600, new_n7601, new_n7602, new_n7603,
    new_n7604, new_n7605, new_n7606, new_n7608, new_n7609, new_n7610_1,
    new_n7611, new_n7612, new_n7613, new_n7614, new_n7615, new_n7616_1,
    new_n7617, new_n7618, new_n7619, new_n7620, new_n7621, new_n7622,
    new_n7623, new_n7624, new_n7625, new_n7626, new_n7627, new_n7628,
    new_n7629, new_n7630_1, new_n7631, new_n7632, new_n7633, new_n7634,
    new_n7635, new_n7636, new_n7637, new_n7638, new_n7639, new_n7640,
    new_n7641, new_n7642, new_n7643_1, new_n7644, new_n7645, new_n7646,
    new_n7647_1, new_n7648, new_n7649, new_n7650, new_n7651, new_n7652,
    new_n7653, new_n7654, new_n7655, new_n7656, new_n7657_1, new_n7658,
    new_n7659, new_n7660, new_n7661, new_n7662, new_n7663, new_n7664,
    new_n7665, new_n7666, new_n7667, new_n7668, new_n7669, new_n7670_1,
    new_n7671, new_n7672, new_n7673, new_n7674_1, new_n7675, new_n7676,
    new_n7677, new_n7678_1, new_n7679_1, new_n7680, new_n7681, new_n7682,
    new_n7683, new_n7684, new_n7685, new_n7686_1, new_n7687, new_n7688,
    new_n7689, new_n7690, new_n7691, new_n7692_1, new_n7693_1, new_n7694,
    new_n7695, new_n7696, new_n7697, new_n7698_1, new_n7699, new_n7700,
    new_n7701, new_n7702, new_n7703, new_n7704, new_n7705, new_n7706,
    new_n7707, new_n7708_1, new_n7709, new_n7710, new_n7711, new_n7712,
    new_n7713, new_n7714, new_n7715, new_n7716, new_n7717, new_n7718,
    new_n7719, new_n7720, new_n7721_1, new_n7722, new_n7723, new_n7724,
    new_n7725, new_n7726, new_n7727, new_n7728, new_n7729, new_n7730,
    new_n7731_1, new_n7732, new_n7733, new_n7734, new_n7735, new_n7736,
    new_n7737, new_n7738, new_n7739, new_n7740, new_n7741, new_n7742,
    new_n7743, new_n7744, new_n7745, new_n7746, new_n7747, new_n7748,
    new_n7749, new_n7750, new_n7751_1, new_n7752, new_n7753, new_n7754,
    new_n7755, new_n7756, new_n7757, new_n7758, new_n7759_1, new_n7760,
    new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766,
    new_n7767, new_n7768, new_n7769_1, new_n7770, new_n7771, new_n7772,
    new_n7773_1, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778,
    new_n7779, new_n7780_1, new_n7781, new_n7782, new_n7783, new_n7784,
    new_n7785, new_n7786, new_n7787, new_n7788_1, new_n7789, new_n7790,
    new_n7791, new_n7792, new_n7793, new_n7794_1, new_n7795, new_n7796,
    new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802,
    new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808,
    new_n7809, new_n7810, new_n7811_1, new_n7812, new_n7813, new_n7814,
    new_n7815, new_n7816, new_n7817, new_n7818, new_n7819, new_n7820,
    new_n7821, new_n7822, new_n7823, new_n7824, new_n7825, new_n7826,
    new_n7827, new_n7828, new_n7829, new_n7830_1, new_n7831, new_n7832,
    new_n7833, new_n7834_1, new_n7835, new_n7836, new_n7837, new_n7838,
    new_n7839, new_n7840, new_n7841_1, new_n7842, new_n7843, new_n7844,
    new_n7845, new_n7846, new_n7847, new_n7848, new_n7849, new_n7850,
    new_n7851, new_n7852, new_n7853, new_n7854, new_n7855, new_n7856,
    new_n7857, new_n7858, new_n7859, new_n7860, new_n7861, new_n7862,
    new_n7863, new_n7864, new_n7865, new_n7866, new_n7867, new_n7868,
    new_n7869, new_n7870, new_n7871, new_n7872, new_n7873, new_n7874,
    new_n7875, new_n7876_1, new_n7877, new_n7878, new_n7879, new_n7880,
    new_n7881, new_n7882, new_n7883, new_n7884_1, new_n7885, new_n7886,
    new_n7887, new_n7888, new_n7889, new_n7890, new_n7891, new_n7892,
    new_n7893, new_n7894, new_n7895, new_n7896, new_n7897, new_n7898,
    new_n7899, new_n7900, new_n7901, new_n7902, new_n7903, new_n7904,
    new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7918, new_n7919, new_n7920, new_n7921, new_n7922, new_n7923,
    new_n7924, new_n7925, new_n7926, new_n7927, new_n7928, new_n7929,
    new_n7930, new_n7931, new_n7932, new_n7933, new_n7934, new_n7935,
    new_n7936, new_n7937_1, new_n7938, new_n7939, new_n7940, new_n7941,
    new_n7942, new_n7943_1, new_n7944, new_n7945, new_n7946, new_n7947,
    new_n7948, new_n7949_1, new_n7950_1, new_n7951, new_n7952, new_n7953,
    new_n7954, new_n7955, new_n7956, new_n7957, new_n7958, new_n7959_1,
    new_n7960, new_n7961, new_n7962, new_n7963_1, new_n7964, new_n7965,
    new_n7966, new_n7967, new_n7968_1, new_n7969, new_n7970, new_n7971,
    new_n7972, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977,
    new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983,
    new_n7984, new_n7985, new_n7986, new_n7987, new_n7988, new_n7989,
    new_n7990, new_n7991, new_n7992_1, new_n7993, new_n7994, new_n7995,
    new_n7996, new_n7997, new_n7998, new_n7999_1, new_n8000, new_n8001,
    new_n8002, new_n8003, new_n8004, new_n8005, new_n8006_1, new_n8007,
    new_n8008, new_n8009, new_n8010, new_n8011, new_n8012, new_n8013,
    new_n8014, new_n8015, new_n8016, new_n8017, new_n8018, new_n8019,
    new_n8020, new_n8021, new_n8022, new_n8023, new_n8024, new_n8025,
    new_n8026, new_n8027_1, new_n8028, new_n8029, new_n8030, new_n8031_1,
    new_n8032, new_n8033, new_n8034, new_n8035, new_n8036, new_n8037,
    new_n8038, new_n8039, new_n8040, new_n8041, new_n8042_1, new_n8043,
    new_n8044, new_n8045, new_n8046, new_n8047, new_n8048, new_n8049,
    new_n8050, new_n8051, new_n8052_1, new_n8053, new_n8054, new_n8055,
    new_n8056, new_n8057, new_n8058, new_n8059, new_n8060, new_n8061,
    new_n8062, new_n8063, new_n8064, new_n8065, new_n8066, new_n8067_1,
    new_n8068, new_n8069, new_n8070, new_n8071, new_n8072, new_n8073,
    new_n8074, new_n8075, new_n8076, new_n8077, new_n8078, new_n8079,
    new_n8080, new_n8081, new_n8082, new_n8083, new_n8084, new_n8085,
    new_n8086, new_n8087, new_n8088, new_n8089, new_n8090, new_n8091,
    new_n8092, new_n8093, new_n8094, new_n8095_1, new_n8096, new_n8097,
    new_n8098, new_n8099, new_n8100, new_n8101, new_n8102, new_n8103_1,
    new_n8104, new_n8105, new_n8106, new_n8107, new_n8108, new_n8109_1,
    new_n8110, new_n8111, new_n8112, new_n8113, new_n8114, new_n8115,
    new_n8116, new_n8117, new_n8118, new_n8119, new_n8120, new_n8121,
    new_n8122, new_n8123, new_n8124, new_n8125, new_n8126, new_n8127_1,
    new_n8128, new_n8129, new_n8130_1, new_n8131, new_n8132, new_n8133,
    new_n8134, new_n8135_1, new_n8136, new_n8137, new_n8138, new_n8139_1,
    new_n8140, new_n8141, new_n8142, new_n8143, new_n8144, new_n8145,
    new_n8146, new_n8147, new_n8148_1, new_n8149_1, new_n8150, new_n8151,
    new_n8152, new_n8153, new_n8154, new_n8155, new_n8156, new_n8157,
    new_n8158, new_n8159_1, new_n8160, new_n8161, new_n8162, new_n8163,
    new_n8164, new_n8165, new_n8166, new_n8167, new_n8168, new_n8169,
    new_n8170, new_n8171, new_n8172, new_n8173, new_n8174, new_n8175,
    new_n8176, new_n8177, new_n8178, new_n8179_1, new_n8180, new_n8181,
    new_n8182, new_n8183, new_n8184, new_n8185, new_n8186, new_n8187,
    new_n8188, new_n8189, new_n8190, new_n8191, new_n8192, new_n8193,
    new_n8194_1, new_n8195, new_n8196, new_n8197, new_n8198, new_n8199,
    new_n8200, new_n8201, new_n8202, new_n8203, new_n8204, new_n8205,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215_1, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244_1, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255_1,
    new_n8256_1, new_n8257, new_n8258, new_n8259_1, new_n8260, new_n8261,
    new_n8262, new_n8263, new_n8264, new_n8265, new_n8266, new_n8267_1,
    new_n8268, new_n8269, new_n8270, new_n8271, new_n8272, new_n8273,
    new_n8274, new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279,
    new_n8280, new_n8281, new_n8282, new_n8283, new_n8284, new_n8285_1,
    new_n8286, new_n8287, new_n8288_1, new_n8289, new_n8290, new_n8291,
    new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297,
    new_n8298, new_n8299, new_n8300, new_n8301, new_n8302, new_n8303,
    new_n8304, new_n8305_1, new_n8306_1, new_n8307, new_n8308, new_n8309_1,
    new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320_1, new_n8321_1,
    new_n8322, new_n8323, new_n8324_1, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336, new_n8337, new_n8338, new_n8339_1,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363_1,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376_1, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381_1,
    new_n8382, new_n8383, new_n8384, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398, new_n8399_1, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405_1, new_n8406,
    new_n8407, new_n8408_1, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417_1, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8432_1, new_n8433, new_n8434, new_n8435, new_n8436, new_n8437,
    new_n8438, new_n8439_1, new_n8440, new_n8441, new_n8442, new_n8443,
    new_n8444, new_n8445, new_n8446, new_n8447, new_n8448, new_n8449,
    new_n8450, new_n8451, new_n8452, new_n8453_1, new_n8454, new_n8455,
    new_n8456, new_n8457, new_n8458, new_n8459, new_n8460, new_n8461,
    new_n8462, new_n8463, new_n8464, new_n8465, new_n8466, new_n8467,
    new_n8468, new_n8469, new_n8470, new_n8471, new_n8472, new_n8473,
    new_n8474, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480_1,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489_1, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505_1, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510_1,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519_1, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526_1, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535_1, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550_1, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563_1, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577,
    new_n8578, new_n8579, new_n8580, new_n8581_1, new_n8582, new_n8583,
    new_n8584, new_n8585, new_n8586, new_n8587, new_n8588, new_n8589,
    new_n8590, new_n8591, new_n8592, new_n8593, new_n8594_1, new_n8595,
    new_n8596, new_n8597, new_n8598, new_n8599, new_n8600, new_n8601,
    new_n8602, new_n8603, new_n8604, new_n8605, new_n8606, new_n8607,
    new_n8608_1, new_n8609, new_n8610, new_n8611, new_n8612, new_n8613,
    new_n8614_1, new_n8615, new_n8616, new_n8617, new_n8618, new_n8619,
    new_n8620_1, new_n8621, new_n8622, new_n8623, new_n8624, new_n8625,
    new_n8626, new_n8627, new_n8628, new_n8629, new_n8630, new_n8631,
    new_n8632, new_n8633, new_n8634, new_n8635, new_n8636, new_n8637_1,
    new_n8638_1, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8645, new_n8646, new_n8647, new_n8648, new_n8649, new_n8650,
    new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656_1,
    new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662_1,
    new_n8663, new_n8664, new_n8665, new_n8666, new_n8667, new_n8668,
    new_n8669, new_n8670, new_n8671, new_n8672, new_n8673, new_n8674,
    new_n8675, new_n8676, new_n8677, new_n8678_1, new_n8679, new_n8680,
    new_n8681, new_n8682, new_n8683, new_n8684, new_n8685, new_n8686,
    new_n8687_1, new_n8688, new_n8689, new_n8690, new_n8691, new_n8692,
    new_n8693, new_n8694_1, new_n8695, new_n8696, new_n8697, new_n8698,
    new_n8699, new_n8700, new_n8701, new_n8702, new_n8703, new_n8704,
    new_n8705, new_n8706, new_n8707, new_n8708, new_n8709, new_n8710,
    new_n8711, new_n8712, new_n8713, new_n8714, new_n8715, new_n8716_1,
    new_n8717, new_n8718, new_n8719, new_n8720, new_n8721_1, new_n8722,
    new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728,
    new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734,
    new_n8735, new_n8736, new_n8737, new_n8738, new_n8739, new_n8740,
    new_n8741, new_n8742, new_n8743, new_n8744_1, new_n8745_1, new_n8746,
    new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752,
    new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758,
    new_n8759, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764,
    new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770,
    new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776,
    new_n8777, new_n8778, new_n8779, new_n8780, new_n8781, new_n8782_1,
    new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788,
    new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794,
    new_n8795, new_n8796, new_n8797, new_n8798, new_n8799, new_n8800,
    new_n8801, new_n8802, new_n8803_1, new_n8804, new_n8805, new_n8806_1,
    new_n8807, new_n8808, new_n8809_1, new_n8810, new_n8811, new_n8812,
    new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818,
    new_n8819, new_n8820, new_n8821_1, new_n8822, new_n8823, new_n8824_1,
    new_n8825, new_n8826, new_n8827_1, new_n8828, new_n8829, new_n8830,
    new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836,
    new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842,
    new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848,
    new_n8849_1, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854,
    new_n8855, new_n8856_1, new_n8857, new_n8858, new_n8859, new_n8860,
    new_n8861_1, new_n8862_1, new_n8863, new_n8864, new_n8865, new_n8866,
    new_n8867, new_n8868, new_n8869_1, new_n8870, new_n8871, new_n8872,
    new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878,
    new_n8879, new_n8880, new_n8881, new_n8882, new_n8883, new_n8884_1,
    new_n8885, new_n8886, new_n8887, new_n8888, new_n8889, new_n8890,
    new_n8891, new_n8892, new_n8893, new_n8894, new_n8895, new_n8896,
    new_n8897, new_n8898, new_n8899, new_n8900, new_n8901, new_n8902,
    new_n8903, new_n8904, new_n8905, new_n8906, new_n8907, new_n8908,
    new_n8909_1, new_n8911_1, new_n8912, new_n8913, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920_1, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943_1, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964_1,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971_1, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982_1,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993_1, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003_1, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012_1,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032_1, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042_1,
    new_n9043, new_n9044, new_n9045, new_n9046_1, new_n9047_1, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9061,
    new_n9062, new_n9063, new_n9064, new_n9065, new_n9066, new_n9067,
    new_n9068, new_n9069, new_n9070, new_n9071, new_n9072, new_n9073,
    new_n9074, new_n9075, new_n9076, new_n9077, new_n9078, new_n9079,
    new_n9080, new_n9081, new_n9082, new_n9083, new_n9084, new_n9085,
    new_n9086, new_n9087, new_n9088, new_n9089, new_n9090_1, new_n9091,
    new_n9092, new_n9093, new_n9094, new_n9095, new_n9096, new_n9097,
    new_n9098, new_n9099, new_n9100, new_n9101, new_n9102, new_n9103,
    new_n9104_1, new_n9105, new_n9106, new_n9107, new_n9108, new_n9109,
    new_n9110, new_n9111, new_n9112, new_n9113, new_n9114, new_n9115,
    new_n9116, new_n9117, new_n9118, new_n9119, new_n9120, new_n9121,
    new_n9122, new_n9123, new_n9124, new_n9125, new_n9126, new_n9127,
    new_n9128, new_n9129_1, new_n9130, new_n9131, new_n9132, new_n9133,
    new_n9134, new_n9135, new_n9136, new_n9137, new_n9138, new_n9139,
    new_n9140, new_n9141, new_n9142, new_n9143, new_n9144, new_n9145,
    new_n9146_1, new_n9147, new_n9148, new_n9149, new_n9150, new_n9151,
    new_n9152, new_n9153, new_n9154, new_n9155, new_n9156, new_n9157,
    new_n9158, new_n9159, new_n9160, new_n9161, new_n9162, new_n9163,
    new_n9164_1, new_n9165, new_n9166_1, new_n9167, new_n9168, new_n9169,
    new_n9170, new_n9171, new_n9172_1, new_n9173, new_n9174, new_n9175,
    new_n9176, new_n9177, new_n9178, new_n9179, new_n9180, new_n9181,
    new_n9182_1, new_n9183, new_n9184, new_n9185, new_n9186, new_n9187,
    new_n9188, new_n9189, new_n9190, new_n9191_1, new_n9192, new_n9193,
    new_n9194, new_n9195, new_n9196, new_n9197, new_n9198, new_n9199,
    new_n9200, new_n9201, new_n9202, new_n9203, new_n9204, new_n9205,
    new_n9206, new_n9207, new_n9208, new_n9209, new_n9210, new_n9211,
    new_n9212, new_n9213, new_n9214, new_n9215, new_n9216, new_n9217_1,
    new_n9218, new_n9219, new_n9220_1, new_n9221, new_n9226, new_n9227,
    new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233,
    new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239,
    new_n9240, new_n9241, new_n9242, new_n9243, new_n9244, new_n9245,
    new_n9246_1, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251_1,
    new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259_1, new_n9260, new_n9261_1, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287_1,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308_1, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318_1, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323_1,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344_1, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364_1, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371_1,
    new_n9372_1, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380_1, new_n9381, new_n9382_1, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9393, new_n9394, new_n9395, new_n9396_1,
    new_n9397, new_n9398, new_n9399_1, new_n9400, new_n9401, new_n9402,
    new_n9403_1, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419_1, new_n9420,
    new_n9421, new_n9422, new_n9423_1, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430_1, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435_1, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445_1, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451_1, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458_1, new_n9459_1, new_n9460_1, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493_1, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507_1, new_n9508_1, new_n9509, new_n9510, new_n9511, new_n9512_1,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552_1, new_n9553, new_n9554_1,
    new_n9555, new_n9556_1, new_n9557_1, new_n9558_1, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9569, new_n9570, new_n9571, new_n9572, new_n9573,
    new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579,
    new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585,
    new_n9586, new_n9587, new_n9588, new_n9589, new_n9590, new_n9591,
    new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597,
    new_n9598_1, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603,
    new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609,
    new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615,
    new_n9616_1, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621,
    new_n9622_1, new_n9623, new_n9624, new_n9625, new_n9626_1, new_n9627,
    new_n9628, new_n9629, new_n9630, new_n9631, new_n9632, new_n9633_1,
    new_n9634, new_n9635_1, new_n9636, new_n9637, new_n9638, new_n9639,
    new_n9640, new_n9641, new_n9642, new_n9643, new_n9644, new_n9645,
    new_n9646_1, new_n9647, new_n9648_1, new_n9649, new_n9650, new_n9651,
    new_n9652, new_n9653, new_n9654, new_n9655_1, new_n9656, new_n9657,
    new_n9658, new_n9659, new_n9660, new_n9661, new_n9662, new_n9663,
    new_n9664, new_n9665, new_n9666, new_n9667, new_n9668, new_n9669,
    new_n9670, new_n9671, new_n9672, new_n9673, new_n9674, new_n9675,
    new_n9676, new_n9677, new_n9678, new_n9679, new_n9680, new_n9681,
    new_n9682, new_n9683, new_n9684, new_n9685, new_n9686, new_n9687,
    new_n9688, new_n9689_1, new_n9690, new_n9691, new_n9692, new_n9693,
    new_n9694, new_n9695_1, new_n9696, new_n9697, new_n9698, new_n9699_1,
    new_n9700, new_n9701, new_n9702, new_n9703, new_n9705, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726_1,
    new_n9727, new_n9729, new_n9731, new_n9732, new_n9733, new_n9734,
    new_n9735, new_n9736, new_n9737, new_n9738, new_n9739, new_n9740,
    new_n9741, new_n9742, new_n9743, new_n9744, new_n9745, new_n9746,
    new_n9747, new_n9748, new_n9749, new_n9750, new_n9751, new_n9752,
    new_n9753_1, new_n9754, new_n9755, new_n9756, new_n9757, new_n9758,
    new_n9759, new_n9760, new_n9761_1, new_n9762, new_n9763_1, new_n9764,
    new_n9765, new_n9766, new_n9767_1, new_n9768, new_n9769, new_n9770,
    new_n9771_1, new_n9772, new_n9773, new_n9774, new_n9775, new_n9776,
    new_n9777, new_n9778_1, new_n9779, new_n9780, new_n9781, new_n9782,
    new_n9783_1, new_n9784, new_n9785, new_n9786, new_n9787, new_n9788,
    new_n9789, new_n9790, new_n9791, new_n9792, new_n9793, new_n9794,
    new_n9795, new_n9796, new_n9797, new_n9798, new_n9799, new_n9800,
    new_n9801, new_n9802, new_n9803_1, new_n9804, new_n9805, new_n9806,
    new_n9807, new_n9808, new_n9809, new_n9810, new_n9811, new_n9812,
    new_n9813, new_n9814, new_n9815, new_n9816, new_n9817, new_n9818,
    new_n9819, new_n9820, new_n9821, new_n9822, new_n9823, new_n9824,
    new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830,
    new_n9831, new_n9832_1, new_n9833_1, new_n9834, new_n9835, new_n9836,
    new_n9837, new_n9838_1, new_n9839, new_n9840, new_n9841, new_n9842,
    new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9848,
    new_n9849, new_n9850, new_n9851, new_n9852, new_n9853, new_n9854,
    new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860,
    new_n9861, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866,
    new_n9867_1, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872_1,
    new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878,
    new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884,
    new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890_1,
    new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9896,
    new_n9897, new_n9898, new_n9899, new_n9900, new_n9901, new_n9902,
    new_n9903, new_n9904, new_n9905, new_n9906, new_n9907, new_n9908,
    new_n9909, new_n9910, new_n9911, new_n9912, new_n9913, new_n9914,
    new_n9915, new_n9916, new_n9917_1, new_n9918, new_n9919_1, new_n9920,
    new_n9921, new_n9922, new_n9923, new_n9924, new_n9925, new_n9926_1,
    new_n9927, new_n9928, new_n9929, new_n9930, new_n9931, new_n9932,
    new_n9933, new_n9934_1, new_n9935, new_n9936, new_n9937, new_n9938_1,
    new_n9939, new_n9940, new_n9941, new_n9942_1, new_n9943, new_n9944,
    new_n9945, new_n9946_1, new_n9947, new_n9948, new_n9949, new_n9950,
    new_n9951, new_n9952, new_n9953, new_n9954, new_n9955, new_n9956,
    new_n9957, new_n9958, new_n9959, new_n9960, new_n9961, new_n9962,
    new_n9963, new_n9964, new_n9965, new_n9966, new_n9967_1, new_n9968_1,
    new_n9969, new_n9970, new_n9971, new_n9972, new_n9973, new_n9974,
    new_n9975, new_n9976, new_n9977, new_n9978, new_n9979, new_n9980,
    new_n9981, new_n9982, new_n9983, new_n9984, new_n9985, new_n9986,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009_1, new_n10010_1,
    new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017_1, new_n10018_1, new_n10019_1, new_n10020, new_n10021_1,
    new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027,
    new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033,
    new_n10034, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039,
    new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045,
    new_n10046, new_n10047, new_n10048, new_n10049, new_n10050, new_n10051,
    new_n10052, new_n10053_1, new_n10054, new_n10055_1, new_n10056,
    new_n10057_1, new_n10058, new_n10059, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096_1,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101_1,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111_1, new_n10112,
    new_n10113, new_n10114, new_n10115, new_n10116, new_n10117_1,
    new_n10118, new_n10119, new_n10120, new_n10121, new_n10122, new_n10123,
    new_n10124, new_n10125_1, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157,
    new_n10158_1, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10165_1, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173, new_n10174,
    new_n10175, new_n10176, new_n10177, new_n10178, new_n10179, new_n10180,
    new_n10181, new_n10182, new_n10183, new_n10184, new_n10185, new_n10186,
    new_n10187, new_n10188, new_n10189, new_n10190, new_n10191, new_n10192,
    new_n10193, new_n10194, new_n10195, new_n10196, new_n10197, new_n10198,
    new_n10199, new_n10200, new_n10201_1, new_n10202, new_n10203,
    new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209,
    new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215,
    new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236_1, new_n10237, new_n10238,
    new_n10239_1, new_n10240, new_n10241, new_n10242, new_n10243,
    new_n10244_1, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250_1, new_n10251, new_n10252, new_n10253,
    new_n10254, new_n10255, new_n10256, new_n10257, new_n10258, new_n10259,
    new_n10260, new_n10261_1, new_n10262_1, new_n10263, new_n10264,
    new_n10265, new_n10266, new_n10267, new_n10268, new_n10269, new_n10270,
    new_n10271, new_n10272, new_n10273, new_n10274, new_n10275_1,
    new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283, new_n10284, new_n10285, new_n10286,
    new_n10287_1, new_n10288, new_n10289, new_n10290, new_n10291,
    new_n10292, new_n10293, new_n10294, new_n10295_1, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321_1, new_n10322, new_n10323, new_n10324, new_n10325,
    new_n10326_1, new_n10327_1, new_n10328, new_n10329, new_n10330_1,
    new_n10331, new_n10332, new_n10333, new_n10334, new_n10335, new_n10336,
    new_n10337, new_n10338, new_n10339, new_n10340_1, new_n10341,
    new_n10342, new_n10343, new_n10344, new_n10345_1, new_n10346,
    new_n10347, new_n10348, new_n10349, new_n10350, new_n10351, new_n10352,
    new_n10353, new_n10354, new_n10355, new_n10356_1, new_n10357,
    new_n10358, new_n10359, new_n10360, new_n10361, new_n10362, new_n10363,
    new_n10364, new_n10365, new_n10366, new_n10367, new_n10368, new_n10369,
    new_n10370, new_n10371, new_n10372_1, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385_1,
    new_n10386, new_n10387_1, new_n10388_1, new_n10389, new_n10390_1,
    new_n10391, new_n10392, new_n10393, new_n10394, new_n10395, new_n10396,
    new_n10397, new_n10398, new_n10399, new_n10400, new_n10401, new_n10402,
    new_n10403, new_n10404_1, new_n10405_1, new_n10406, new_n10407,
    new_n10408, new_n10409_1, new_n10410, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420_1, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432_1, new_n10433, new_n10434, new_n10435,
    new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476, new_n10477,
    new_n10478, new_n10479, new_n10480, new_n10481, new_n10482, new_n10483,
    new_n10484_1, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489_1, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514_1, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525_1, new_n10526, new_n10527, new_n10528,
    new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534,
    new_n10535, new_n10536, new_n10537, new_n10538, new_n10539,
    new_n10540_1, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561_1,
    new_n10562, new_n10563, new_n10564_1, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577_1,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588_1,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593_1,
    new_n10594, new_n10595_1, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611_1, new_n10612, new_n10613, new_n10614_1, new_n10615,
    new_n10616, new_n10617_1, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628_1, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647_1, new_n10648,
    new_n10649, new_n10650_1, new_n10651, new_n10652, new_n10653_1,
    new_n10654, new_n10655, new_n10656, new_n10657, new_n10658, new_n10659,
    new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665,
    new_n10666, new_n10667, new_n10668, new_n10669, new_n10670, new_n10671,
    new_n10672, new_n10673, new_n10674, new_n10675, new_n10676, new_n10677,
    new_n10678, new_n10679, new_n10680, new_n10681, new_n10682, new_n10683,
    new_n10684, new_n10685, new_n10686, new_n10687, new_n10688, new_n10689,
    new_n10690, new_n10691, new_n10692_1, new_n10693, new_n10694_1,
    new_n10695, new_n10696, new_n10697, new_n10698, new_n10699, new_n10700,
    new_n10701_1, new_n10702, new_n10703, new_n10704, new_n10705,
    new_n10706, new_n10707, new_n10708, new_n10709, new_n10710_1,
    new_n10711, new_n10712_1, new_n10713, new_n10714, new_n10715,
    new_n10716, new_n10717, new_n10718, new_n10719, new_n10720, new_n10721,
    new_n10722, new_n10723, new_n10724, new_n10725, new_n10726, new_n10727,
    new_n10728, new_n10729, new_n10730, new_n10731, new_n10732, new_n10733,
    new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739_1, new_n10740, new_n10741, new_n10742, new_n10743,
    new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749,
    new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755,
    new_n10756_1, new_n10757, new_n10758, new_n10759, new_n10760,
    new_n10761, new_n10762, new_n10763_1, new_n10764, new_n10765,
    new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771,
    new_n10772, new_n10773, new_n10774, new_n10775_1, new_n10777,
    new_n10778, new_n10779, new_n10781, new_n10782, new_n10783, new_n10784,
    new_n10785, new_n10786, new_n10787, new_n10788, new_n10789, new_n10790,
    new_n10791, new_n10792_1, new_n10793, new_n10794, new_n10795,
    new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807,
    new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817_1, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834_1, new_n10835,
    new_n10836, new_n10837, new_n10838, new_n10839, new_n10840, new_n10841,
    new_n10842, new_n10843, new_n10844, new_n10845, new_n10846, new_n10847,
    new_n10848, new_n10849, new_n10850, new_n10851_1, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10870, new_n10871,
    new_n10872, new_n10873, new_n10874_1, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923,
    new_n10924_1, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943_1, new_n10944, new_n10945,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961_1, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005_1, new_n11006, new_n11007, new_n11008, new_n11009,
    new_n11010, new_n11011_1, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023_1, new_n11024, new_n11025_1,
    new_n11026, new_n11027, new_n11028, new_n11029, new_n11030, new_n11031,
    new_n11032, new_n11033, new_n11034, new_n11035, new_n11036, new_n11037,
    new_n11038, new_n11039, new_n11040, new_n11041, new_n11042, new_n11043,
    new_n11044_1, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056_1, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063_1, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078_1, new_n11079, new_n11080_1, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11092, new_n11093,
    new_n11094_1, new_n11095, new_n11096, new_n11097, new_n11098,
    new_n11099, new_n11100, new_n11101_1, new_n11102, new_n11103_1,
    new_n11104, new_n11105, new_n11106, new_n11107, new_n11108, new_n11109,
    new_n11110, new_n11111, new_n11112, new_n11113, new_n11114, new_n11115,
    new_n11116, new_n11117, new_n11118, new_n11119, new_n11120_1,
    new_n11121_1, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127_1, new_n11128, new_n11129, new_n11130,
    new_n11131, new_n11132_1, new_n11133, new_n11134_1, new_n11135,
    new_n11136, new_n11137, new_n11138_1, new_n11139, new_n11140,
    new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178,
    new_n11179, new_n11180, new_n11181, new_n11182_1, new_n11183,
    new_n11184_1, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192_1, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201_1, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220_1, new_n11221,
    new_n11222, new_n11223_1, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234_1, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245_1, new_n11246, new_n11247, new_n11248,
    new_n11249, new_n11250, new_n11251, new_n11252, new_n11253, new_n11254,
    new_n11255, new_n11256, new_n11257, new_n11258, new_n11259, new_n11260,
    new_n11261_1, new_n11262, new_n11263, new_n11264, new_n11265,
    new_n11266_1, new_n11267, new_n11272, new_n11273_1, new_n11274,
    new_n11275_1, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290_1,
    new_n11291, new_n11292, new_n11293, new_n11294, new_n11295, new_n11296,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301,
    new_n11302_1, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313_1, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323,
    new_n11324, new_n11325_1, new_n11326_1, new_n11327, new_n11328,
    new_n11329, new_n11330_1, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345,
    new_n11346, new_n11347_1, new_n11348_1, new_n11349, new_n11350,
    new_n11351, new_n11352_1, new_n11353, new_n11354, new_n11355,
    new_n11356_1, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375_1, new_n11376, new_n11377,
    new_n11378, new_n11379_1, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386_1, new_n11387,
    new_n11388, new_n11389, new_n11390, new_n11391_1, new_n11392,
    new_n11393, new_n11394, new_n11395, new_n11396, new_n11397,
    new_n11398_1, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403_1, new_n11404, new_n11405, new_n11406, new_n11407,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11415, new_n11416, new_n11417, new_n11418, new_n11419_1,
    new_n11420, new_n11421, new_n11422, new_n11423, new_n11424_1,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439_1, new_n11440, new_n11441,
    new_n11442, new_n11443, new_n11444, new_n11445, new_n11446, new_n11447,
    new_n11448, new_n11449, new_n11450, new_n11451, new_n11452, new_n11453,
    new_n11454, new_n11455_1, new_n11456, new_n11457, new_n11458,
    new_n11459, new_n11460, new_n11461, new_n11462_1, new_n11463,
    new_n11464, new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470_1, new_n11471, new_n11472_1, new_n11473_1, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479_1,
    new_n11480, new_n11481_1, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486_1, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496_1, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503_1, new_n11504, new_n11505,
    new_n11506_1, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515_1,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536, new_n11537, new_n11538_1,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548_1, new_n11549,
    new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555,
    new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561,
    new_n11562, new_n11563, new_n11564_1, new_n11565, new_n11566_1,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579_1, new_n11580_1, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11590, new_n11591_1,
    new_n11592, new_n11593, new_n11594, new_n11595, new_n11596, new_n11597,
    new_n11598, new_n11599, new_n11600, new_n11603, new_n11605, new_n11606,
    new_n11607_1, new_n11608, new_n11609, new_n11610, new_n11611,
    new_n11612, new_n11613, new_n11614, new_n11615_1, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630_1, new_n11631, new_n11634, new_n11635,
    new_n11636, new_n11637, new_n11638, new_n11639, new_n11640, new_n11641,
    new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647_1, new_n11648, new_n11649, new_n11650, new_n11651,
    new_n11652, new_n11653, new_n11654, new_n11655, new_n11656, new_n11657,
    new_n11658, new_n11659, new_n11660, new_n11661, new_n11662, new_n11663,
    new_n11664, new_n11665, new_n11666, new_n11667_1, new_n11668,
    new_n11669, new_n11670, new_n11671, new_n11672, new_n11673,
    new_n11674_1, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682_1, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706, new_n11707,
    new_n11708, new_n11709, new_n11710_1, new_n11711, new_n11712_1,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724_1, new_n11725, new_n11726, new_n11727, new_n11728,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736_1, new_n11737, new_n11738, new_n11739,
    new_n11740, new_n11741_1, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749_1,
    new_n11750, new_n11751, new_n11752, new_n11753, new_n11754, new_n11755,
    new_n11756, new_n11757, new_n11758, new_n11759, new_n11760, new_n11761,
    new_n11762, new_n11763, new_n11764, new_n11765, new_n11766, new_n11767,
    new_n11768, new_n11769, new_n11770_1, new_n11771_1, new_n11772,
    new_n11773, new_n11774, new_n11775_1, new_n11776, new_n11777,
    new_n11778, new_n11779, new_n11780, new_n11781, new_n11782, new_n11783,
    new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789,
    new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818_1, new_n11819, new_n11820,
    new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826,
    new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832,
    new_n11833, new_n11834, new_n11835, new_n11836, new_n11837_1,
    new_n11838, new_n11839, new_n11840, new_n11841_1, new_n11842_1,
    new_n11843_1, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898_1, new_n11899, new_n11900,
    new_n11901, new_n11902, new_n11903, new_n11904, new_n11905_1,
    new_n11906, new_n11907, new_n11909, new_n11910, new_n11911, new_n11912,
    new_n11913, new_n11914, new_n11915, new_n11916, new_n11917, new_n11918,
    new_n11919, new_n11920, new_n11921, new_n11922, new_n11923, new_n11924,
    new_n11925, new_n11926_1, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964,
    new_n11965_1, new_n11966, new_n11967, new_n11968, new_n11969,
    new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975,
    new_n11976, new_n11977, new_n11978, new_n11979, new_n11980_1,
    new_n11981, new_n11982, new_n11983, new_n11984, new_n11985, new_n11986,
    new_n11987, new_n11988, new_n11989, new_n11990, new_n11991, new_n11992,
    new_n11993, new_n11994, new_n11995, new_n11996, new_n11997, new_n11998,
    new_n11999, new_n12000_1, new_n12001, new_n12002, new_n12003_1,
    new_n12004, new_n12005, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011_1, new_n12012, new_n12013, new_n12014,
    new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021,
    new_n12022, new_n12023, new_n12024, new_n12025, new_n12026, new_n12027,
    new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033,
    new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039,
    new_n12040, new_n12041, new_n12045, new_n12046, new_n12047, new_n12048,
    new_n12049, new_n12050, new_n12051, new_n12052, new_n12053, new_n12054,
    new_n12055, new_n12056, new_n12057, new_n12058, new_n12059, new_n12060,
    new_n12061, new_n12062, new_n12063, new_n12064, new_n12065, new_n12066,
    new_n12067, new_n12068, new_n12069, new_n12070, new_n12071,
    new_n12072_1, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12110, new_n12111, new_n12112, new_n12113_1,
    new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119,
    new_n12120, new_n12121_1, new_n12122, new_n12123, new_n12124,
    new_n12125, new_n12126, new_n12127, new_n12128, new_n12129, new_n12130,
    new_n12131_1, new_n12132, new_n12133, new_n12134, new_n12135,
    new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141,
    new_n12142, new_n12143, new_n12144, new_n12145, new_n12146_1,
    new_n12147, new_n12148, new_n12149, new_n12150, new_n12151,
    new_n12152_1, new_n12153_1, new_n12154, new_n12155, new_n12156,
    new_n12157_1, new_n12158_1, new_n12159, new_n12160, new_n12161_1,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12172, new_n12173,
    new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179_1, new_n12180, new_n12181, new_n12182, new_n12183,
    new_n12184, new_n12185, new_n12186, new_n12187, new_n12188, new_n12189,
    new_n12190, new_n12191, new_n12192_1, new_n12193, new_n12194,
    new_n12195, new_n12196, new_n12197, new_n12198, new_n12199, new_n12200,
    new_n12201, new_n12202, new_n12203, new_n12204, new_n12205, new_n12206,
    new_n12207, new_n12208, new_n12209_1, new_n12210, new_n12211,
    new_n12212, new_n12213, new_n12214, new_n12215, new_n12216, new_n12217,
    new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223_1, new_n12224, new_n12225_1, new_n12226, new_n12227,
    new_n12228_1, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235_1, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247, new_n12248, new_n12249,
    new_n12250, new_n12251, new_n12252, new_n12253, new_n12254, new_n12255,
    new_n12256, new_n12257, new_n12258, new_n12259, new_n12260, new_n12261,
    new_n12262, new_n12263, new_n12264, new_n12265, new_n12266, new_n12267,
    new_n12268, new_n12269, new_n12270, new_n12271, new_n12272, new_n12273,
    new_n12274, new_n12275, new_n12276, new_n12277, new_n12278, new_n12279,
    new_n12280, new_n12281, new_n12282, new_n12283, new_n12284, new_n12285,
    new_n12286, new_n12287, new_n12288, new_n12289, new_n12290, new_n12291,
    new_n12292, new_n12293, new_n12294, new_n12295, new_n12296, new_n12297,
    new_n12298, new_n12299, new_n12300, new_n12301, new_n12302_1,
    new_n12303, new_n12304_1, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315_1, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12324_1, new_n12325_1,
    new_n12326, new_n12327, new_n12328, new_n12329_1, new_n12330_1,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12336,
    new_n12337, new_n12338, new_n12339, new_n12340, new_n12341_1,
    new_n12342, new_n12343, new_n12344, new_n12345, new_n12346_1,
    new_n12347, new_n12348, new_n12349_1, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12355, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363,
    new_n12364_1, new_n12365, new_n12366, new_n12367, new_n12368,
    new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374,
    new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380_1, new_n12381, new_n12382, new_n12383_1, new_n12384_1,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397_1, new_n12398_1, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408_1, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446_1, new_n12447,
    new_n12448, new_n12449_1, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461_1, new_n12462_1, new_n12463,
    new_n12464, new_n12465, new_n12466, new_n12467_1, new_n12468,
    new_n12469_1, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495_1, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507_1,
    new_n12508, new_n12509, new_n12510, new_n12511, new_n12512, new_n12513,
    new_n12514, new_n12515_1, new_n12516_1, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540_1, new_n12541,
    new_n12542, new_n12543, new_n12544, new_n12545_1, new_n12546_1,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552_1, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561,
    new_n12562_1, new_n12563, new_n12564, new_n12565, new_n12566_1,
    new_n12567, new_n12568, new_n12569_1, new_n12570, new_n12571,
    new_n12572, new_n12573, new_n12574, new_n12575, new_n12576, new_n12577,
    new_n12578, new_n12579, new_n12580, new_n12581, new_n12582, new_n12583,
    new_n12584, new_n12585, new_n12586, new_n12587_1, new_n12588,
    new_n12589, new_n12590, new_n12591, new_n12592, new_n12593_1,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607_1, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620_1, new_n12621_1,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626_1,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649,
    new_n12650_1, new_n12651, new_n12652, new_n12653, new_n12654_1,
    new_n12655, new_n12656, new_n12657_1, new_n12658, new_n12659,
    new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665_1, new_n12666, new_n12667, new_n12670_1, new_n12671,
    new_n12672, new_n12673, new_n12674, new_n12675, new_n12676, new_n12677,
    new_n12678, new_n12679, new_n12680, new_n12681, new_n12682, new_n12683,
    new_n12684, new_n12685, new_n12686, new_n12687, new_n12688, new_n12689,
    new_n12690, new_n12691, new_n12692, new_n12693, new_n12694, new_n12695,
    new_n12696, new_n12697, new_n12698, new_n12699, new_n12700, new_n12701,
    new_n12702_1, new_n12703, new_n12704, new_n12705, new_n12706,
    new_n12707_1, new_n12708, new_n12709, new_n12710, new_n12711,
    new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717,
    new_n12718, new_n12719, new_n12720, new_n12721, new_n12722, new_n12723,
    new_n12724, new_n12725_1, new_n12726, new_n12727_1, new_n12728,
    new_n12729, new_n12730, new_n12731, new_n12732, new_n12737, new_n12738,
    new_n12739, new_n12740_1, new_n12741, new_n12742_1, new_n12743,
    new_n12744, new_n12745, new_n12746_1, new_n12747, new_n12748,
    new_n12749, new_n12750, new_n12754, new_n12755, new_n12756_1,
    new_n12757, new_n12758, new_n12759, new_n12760, new_n12761, new_n12762,
    new_n12763, new_n12764, new_n12765, new_n12766, new_n12767, new_n12768,
    new_n12769, new_n12770, new_n12771, new_n12772, new_n12773, new_n12774,
    new_n12778, new_n12779, new_n12780, new_n12781, new_n12782,
    new_n12783_1, new_n12784, new_n12785, new_n12786, new_n12787,
    new_n12788, new_n12789, new_n12790, new_n12791, new_n12792, new_n12793,
    new_n12794, new_n12795, new_n12796, new_n12797, new_n12798, new_n12799,
    new_n12800, new_n12801_1, new_n12802, new_n12803, new_n12804,
    new_n12805, new_n12806, new_n12808, new_n12809, new_n12810,
    new_n12811_1, new_n12812_1, new_n12813, new_n12814, new_n12815,
    new_n12816_1, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821_1, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12840,
    new_n12841, new_n12842, new_n12843_1, new_n12844, new_n12845,
    new_n12846, new_n12847, new_n12848, new_n12849, new_n12850, new_n12851,
    new_n12852, new_n12853, new_n12854, new_n12855, new_n12856, new_n12857,
    new_n12858, new_n12859, new_n12860, new_n12861_1, new_n12862,
    new_n12863, new_n12864_1, new_n12865_1, new_n12866, new_n12867,
    new_n12868, new_n12869, new_n12870_1, new_n12871_1, new_n12872,
    new_n12873_1, new_n12874, new_n12875_1, new_n12876, new_n12877,
    new_n12878, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892_1, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900_1, new_n12901,
    new_n12902, new_n12903, new_n12904_1, new_n12905, new_n12906,
    new_n12907, new_n12908, new_n12909, new_n12910, new_n12911, new_n12912,
    new_n12913, new_n12914, new_n12915, new_n12916, new_n12917_1,
    new_n12918, new_n12919, new_n12920, new_n12921, new_n12922, new_n12923,
    new_n12924, new_n12925, new_n12926, new_n12927, new_n12928, new_n12929,
    new_n12930, new_n12931, new_n12932, new_n12933, new_n12934, new_n12935,
    new_n12936, new_n12937, new_n12938, new_n12939, new_n12940,
    new_n12941_1, new_n12942_1, new_n12943, new_n12944, new_n12945,
    new_n12946, new_n12947, new_n12948, new_n12949, new_n12950, new_n12951,
    new_n12952, new_n12953, new_n12954, new_n12955, new_n12956_1,
    new_n12957, new_n12958, new_n12959, new_n12960, new_n12961, new_n12962,
    new_n12963, new_n12964, new_n12965, new_n12966, new_n12967, new_n12968,
    new_n12969, new_n12970, new_n12971, new_n12972, new_n12973, new_n12974,
    new_n12975, new_n12976, new_n12977, new_n12978_1, new_n12979,
    new_n12980_1, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985_1, new_n12986, new_n12987_1, new_n12988, new_n12989,
    new_n12991, new_n12992_1, new_n12993, new_n12994, new_n12995,
    new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001,
    new_n13002, new_n13003, new_n13004, new_n13005_1, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026_1, new_n13027, new_n13028, new_n13029,
    new_n13030, new_n13031, new_n13032, new_n13033, new_n13034, new_n13035,
    new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041,
    new_n13042, new_n13043_1, new_n13044_1, new_n13045, new_n13046,
    new_n13047, new_n13048_1, new_n13049, new_n13050, new_n13051,
    new_n13052, new_n13053, new_n13054_1, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073,
    new_n13074_1, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082_1, new_n13083,
    new_n13084, new_n13085, new_n13086, new_n13087, new_n13088, new_n13089,
    new_n13090, new_n13091, new_n13092, new_n13093, new_n13094, new_n13095,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110_1, new_n13111, new_n13112, new_n13113,
    new_n13114, new_n13115, new_n13116_1, new_n13117, new_n13118,
    new_n13119, new_n13120, new_n13121, new_n13122_1, new_n13123,
    new_n13124, new_n13125, new_n13126, new_n13127, new_n13128, new_n13129,
    new_n13130, new_n13131, new_n13132, new_n13133, new_n13134, new_n13135,
    new_n13136, new_n13137_1, new_n13138, new_n13139, new_n13142,
    new_n13143, new_n13144_1, new_n13145, new_n13146, new_n13147,
    new_n13148, new_n13149, new_n13150, new_n13151, new_n13153, new_n13154,
    new_n13155, new_n13156, new_n13157, new_n13158, new_n13159, new_n13160,
    new_n13161, new_n13162, new_n13163, new_n13164, new_n13165, new_n13166,
    new_n13167, new_n13168_1, new_n13169, new_n13170, new_n13171,
    new_n13172, new_n13173, new_n13174, new_n13175, new_n13176, new_n13177,
    new_n13178, new_n13179, new_n13180, new_n13181, new_n13182, new_n13183,
    new_n13184, new_n13185, new_n13186, new_n13187, new_n13188, new_n13189,
    new_n13190_1, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198_1, new_n13199_1,
    new_n13200, new_n13201, new_n13202, new_n13203, new_n13204_1,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209_1,
    new_n13210, new_n13211, new_n13212, new_n13213, new_n13214, new_n13215,
    new_n13216, new_n13217, new_n13218, new_n13219, new_n13220, new_n13221,
    new_n13222, new_n13223, new_n13224, new_n13225, new_n13226, new_n13227,
    new_n13228, new_n13229, new_n13230, new_n13231, new_n13232, new_n13233,
    new_n13234, new_n13235, new_n13236, new_n13237, new_n13238, new_n13239,
    new_n13240, new_n13241, new_n13242, new_n13243, new_n13244, new_n13245,
    new_n13246, new_n13247, new_n13248, new_n13249, new_n13250, new_n13251,
    new_n13252, new_n13253, new_n13254, new_n13255, new_n13256, new_n13257,
    new_n13258, new_n13259, new_n13260, new_n13261, new_n13262,
    new_n13263_1, new_n13264, new_n13265, new_n13266, new_n13267,
    new_n13268, new_n13269, new_n13270_1, new_n13271, new_n13272,
    new_n13273_1, new_n13274, new_n13275, new_n13276, new_n13277,
    new_n13278, new_n13279, new_n13280, new_n13281, new_n13282, new_n13283,
    new_n13284, new_n13285_1, new_n13286, new_n13287, new_n13288,
    new_n13289, new_n13290, new_n13291, new_n13292, new_n13293, new_n13294,
    new_n13295, new_n13296, new_n13297, new_n13298, new_n13299, new_n13300,
    new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306,
    new_n13307, new_n13308, new_n13309, new_n13310, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319_1,
    new_n13320, new_n13321, new_n13322, new_n13323, new_n13324, new_n13325,
    new_n13326, new_n13327, new_n13328, new_n13329, new_n13330, new_n13331,
    new_n13332, new_n13333_1, new_n13334, new_n13335, new_n13336,
    new_n13337, new_n13338_1, new_n13339, new_n13340, new_n13341,
    new_n13342, new_n13343, new_n13344, new_n13345, new_n13346, new_n13347,
    new_n13348, new_n13349, new_n13350, new_n13351, new_n13352, new_n13353,
    new_n13354, new_n13355, new_n13356, new_n13357, new_n13358, new_n13359,
    new_n13360, new_n13361, new_n13362, new_n13363, new_n13364, new_n13365,
    new_n13366, new_n13367_1, new_n13368, new_n13369, new_n13370,
    new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13376,
    new_n13377, new_n13378, new_n13379, new_n13380, new_n13381, new_n13382,
    new_n13383, new_n13384, new_n13385, new_n13386, new_n13387, new_n13388,
    new_n13389, new_n13390, new_n13392, new_n13393, new_n13394, new_n13395,
    new_n13396, new_n13397, new_n13398, new_n13399, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407_1, new_n13408,
    new_n13409_1, new_n13410, new_n13411, new_n13412, new_n13413,
    new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419_1, new_n13420, new_n13421, new_n13422, new_n13423,
    new_n13424_1, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453_1, new_n13454, new_n13455, new_n13456_1, new_n13457_1,
    new_n13458, new_n13459, new_n13460_1, new_n13461, new_n13462,
    new_n13463, new_n13464, new_n13465, new_n13466, new_n13467, new_n13468,
    new_n13469, new_n13470, new_n13471, new_n13472, new_n13473, new_n13474,
    new_n13475, new_n13476, new_n13477_1, new_n13478, new_n13479,
    new_n13480, new_n13481, new_n13482, new_n13484_1, new_n13485,
    new_n13486_1, new_n13487_1, new_n13488, new_n13489, new_n13490_1,
    new_n13491, new_n13492, new_n13493, new_n13494_1, new_n13495,
    new_n13496, new_n13497, new_n13498, new_n13499, new_n13500_1,
    new_n13501_1, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506_1, new_n13507, new_n13508, new_n13509, new_n13510,
    new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13532, new_n13533, new_n13534,
    new_n13535, new_n13536, new_n13537, new_n13538, new_n13539, new_n13540,
    new_n13541, new_n13542, new_n13543, new_n13544, new_n13545, new_n13546,
    new_n13547, new_n13548_1, new_n13549_1, new_n13550, new_n13551_1,
    new_n13552, new_n13553, new_n13554, new_n13555, new_n13556, new_n13557,
    new_n13558, new_n13559, new_n13560, new_n13561, new_n13562, new_n13563,
    new_n13564, new_n13565, new_n13566, new_n13567, new_n13568, new_n13569,
    new_n13570, new_n13571, new_n13572, new_n13573, new_n13574, new_n13575,
    new_n13576, new_n13577, new_n13578, new_n13579, new_n13580, new_n13581,
    new_n13582, new_n13583, new_n13584, new_n13585, new_n13586, new_n13587,
    new_n13588, new_n13589, new_n13590, new_n13591, new_n13592, new_n13593,
    new_n13594, new_n13595, new_n13598, new_n13599, new_n13600, new_n13601,
    new_n13602_1, new_n13603, new_n13604, new_n13605, new_n13606,
    new_n13607, new_n13608, new_n13609, new_n13610, new_n13611, new_n13612,
    new_n13613, new_n13614, new_n13615, new_n13616, new_n13617, new_n13618,
    new_n13619, new_n13620, new_n13621, new_n13622, new_n13623, new_n13624,
    new_n13625, new_n13626_1, new_n13627, new_n13628, new_n13629,
    new_n13630, new_n13631, new_n13632, new_n13633, new_n13634, new_n13635,
    new_n13636, new_n13637, new_n13638, new_n13639, new_n13640, new_n13643,
    new_n13644, new_n13645, new_n13646, new_n13647, new_n13648, new_n13649,
    new_n13650, new_n13651, new_n13652, new_n13653, new_n13654, new_n13655,
    new_n13656, new_n13657, new_n13658, new_n13659, new_n13660, new_n13661,
    new_n13662, new_n13663, new_n13664, new_n13665, new_n13666, new_n13667,
    new_n13668_1, new_n13669, new_n13670, new_n13671, new_n13672,
    new_n13673, new_n13674, new_n13675, new_n13676, new_n13677_1,
    new_n13678, new_n13679, new_n13680, new_n13681, new_n13682,
    new_n13683_1, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708_1, new_n13709, new_n13710_1,
    new_n13711, new_n13712, new_n13713, new_n13714_1, new_n13715,
    new_n13716, new_n13717, new_n13718, new_n13719_1, new_n13720,
    new_n13721, new_n13722_1, new_n13723, new_n13724, new_n13725,
    new_n13726, new_n13727, new_n13728, new_n13729, new_n13730, new_n13731,
    new_n13732, new_n13733, new_n13734, new_n13735, new_n13736, new_n13737,
    new_n13738, new_n13739, new_n13740, new_n13741, new_n13742, new_n13743,
    new_n13744, new_n13745, new_n13746, new_n13747, new_n13748, new_n13749,
    new_n13750, new_n13751, new_n13752, new_n13753, new_n13754_1,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764_1, new_n13765,
    new_n13766, new_n13767, new_n13768, new_n13769, new_n13770, new_n13771,
    new_n13772, new_n13773, new_n13774, new_n13775_1, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781_1,
    new_n13783_1, new_n13784, new_n13785, new_n13786, new_n13787,
    new_n13788, new_n13789, new_n13790, new_n13791, new_n13792, new_n13793,
    new_n13794, new_n13795, new_n13796, new_n13797, new_n13798_1,
    new_n13799, new_n13800, new_n13801, new_n13802, new_n13803, new_n13804,
    new_n13805, new_n13806, new_n13807, new_n13808, new_n13810, new_n13811,
    new_n13812, new_n13813, new_n13814, new_n13815, new_n13816, new_n13817,
    new_n13818, new_n13819, new_n13820, new_n13821, new_n13822, new_n13823,
    new_n13824, new_n13825, new_n13826, new_n13827, new_n13828, new_n13829,
    new_n13830, new_n13831, new_n13832, new_n13833, new_n13834,
    new_n13835_1, new_n13836, new_n13837, new_n13838, new_n13839,
    new_n13840, new_n13841, new_n13842, new_n13843, new_n13844, new_n13845,
    new_n13846, new_n13847, new_n13848, new_n13849, new_n13850_1,
    new_n13851_1, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912_1, new_n13913, new_n13914_1,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922_1, new_n13923_1, new_n13924, new_n13925,
    new_n13926, new_n13927, new_n13928, new_n13929, new_n13930, new_n13931,
    new_n13932, new_n13933, new_n13934, new_n13935, new_n13936, new_n13937,
    new_n13938, new_n13939, new_n13940, new_n13941, new_n13942, new_n13943,
    new_n13944, new_n13945, new_n13946, new_n13947, new_n13948, new_n13949,
    new_n13950, new_n13951_1, new_n13952, new_n13953, new_n13954,
    new_n13955, new_n13956, new_n13957, new_n13958, new_n13959, new_n13960,
    new_n13961, new_n13962, new_n13963, new_n13964, new_n13965, new_n13966,
    new_n13967, new_n13968, new_n13969, new_n13970, new_n13971, new_n13972,
    new_n13973, new_n13974, new_n13975, new_n13976, new_n13977, new_n13978,
    new_n13979, new_n13980, new_n13981, new_n13982, new_n13983, new_n13984,
    new_n13985, new_n13986, new_n13987, new_n13988, new_n13989, new_n13990,
    new_n13991, new_n13992, new_n13993, new_n13994, new_n13996, new_n13997,
    new_n13998, new_n13999, new_n14000, new_n14001, new_n14002, new_n14003,
    new_n14004_1, new_n14005, new_n14006, new_n14007, new_n14008,
    new_n14009, new_n14010, new_n14011, new_n14012, new_n14013, new_n14014,
    new_n14015, new_n14016, new_n14017, new_n14018, new_n14019, new_n14020,
    new_n14021, new_n14022, new_n14023, new_n14024, new_n14025, new_n14026,
    new_n14027, new_n14028, new_n14029, new_n14030, new_n14031, new_n14032,
    new_n14033, new_n14034, new_n14035, new_n14036_1, new_n14037,
    new_n14038, new_n14039, new_n14040, new_n14041, new_n14042, new_n14043,
    new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049,
    new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055,
    new_n14056, new_n14057, new_n14058, new_n14059_1, new_n14060,
    new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066,
    new_n14067, new_n14068, new_n14069, new_n14070, new_n14071_1,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081_1, new_n14082,
    new_n14083, new_n14084, new_n14085, new_n14086, new_n14087, new_n14088,
    new_n14089, new_n14090_1, new_n14091, new_n14092, new_n14093,
    new_n14094, new_n14095_1, new_n14096, new_n14097, new_n14098,
    new_n14099, new_n14100, new_n14101, new_n14102, new_n14103, new_n14104,
    new_n14105, new_n14106, new_n14107_1, new_n14108, new_n14109,
    new_n14110, new_n14111, new_n14112, new_n14113, new_n14114, new_n14115,
    new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121_1, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126_1, new_n14127, new_n14128, new_n14129, new_n14130_1,
    new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136_1, new_n14137, new_n14138, new_n14139, new_n14140,
    new_n14141, new_n14142, new_n14143, new_n14144, new_n14145, new_n14146,
    new_n14147_1, new_n14148_1, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14164,
    new_n14165, new_n14166, new_n14167, new_n14168, new_n14169, new_n14170,
    new_n14171, new_n14172, new_n14173, new_n14174_1, new_n14175,
    new_n14176, new_n14177, new_n14178, new_n14179, new_n14180, new_n14181,
    new_n14182, new_n14183, new_n14184, new_n14185, new_n14186, new_n14187,
    new_n14188, new_n14189, new_n14190_1, new_n14191, new_n14192,
    new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198,
    new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204,
    new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210,
    new_n14211_1, new_n14212, new_n14213, new_n14214, new_n14215,
    new_n14216, new_n14217, new_n14218, new_n14219, new_n14220, new_n14221,
    new_n14222_1, new_n14223, new_n14224, new_n14225, new_n14226,
    new_n14227, new_n14228, new_n14229, new_n14230_1, new_n14231,
    new_n14232, new_n14233, new_n14234, new_n14235, new_n14236, new_n14237,
    new_n14238, new_n14239, new_n14240, new_n14241, new_n14242, new_n14243,
    new_n14244, new_n14245, new_n14246, new_n14247, new_n14248, new_n14249,
    new_n14250, new_n14251, new_n14252, new_n14253, new_n14254, new_n14255,
    new_n14256, new_n14257, new_n14258, new_n14259, new_n14260, new_n14261,
    new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267_1, new_n14268, new_n14269, new_n14270, new_n14271_1,
    new_n14272, new_n14273, new_n14274, new_n14275_1, new_n14276,
    new_n14277_1, new_n14278, new_n14279, new_n14280, new_n14281,
    new_n14282, new_n14283, new_n14284, new_n14285, new_n14286, new_n14287,
    new_n14288, new_n14289, new_n14290, new_n14291, new_n14292, new_n14293,
    new_n14294_1, new_n14295, new_n14296, new_n14297, new_n14298,
    new_n14299, new_n14300, new_n14301, new_n14302, new_n14303, new_n14304,
    new_n14305, new_n14306, new_n14307, new_n14309, new_n14310_1,
    new_n14311, new_n14312, new_n14313, new_n14314, new_n14315, new_n14316,
    new_n14317, new_n14318, new_n14319, new_n14320, new_n14321, new_n14322,
    new_n14323_1, new_n14324, new_n14325, new_n14326_1, new_n14327,
    new_n14328, new_n14329, new_n14330, new_n14331, new_n14332, new_n14333,
    new_n14334, new_n14335, new_n14336, new_n14337, new_n14338, new_n14339,
    new_n14340, new_n14341, new_n14342_1, new_n14343, new_n14344,
    new_n14345_1, new_n14346, new_n14347, new_n14348, new_n14349,
    new_n14350, new_n14351, new_n14352, new_n14353_1, new_n14354,
    new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360,
    new_n14361, new_n14362, new_n14363, new_n14364_1, new_n14365,
    new_n14366, new_n14367, new_n14368, new_n14369, new_n14370, new_n14371,
    new_n14372, new_n14373, new_n14374, new_n14375_1, new_n14376,
    new_n14377, new_n14378, new_n14379, new_n14380, new_n14381, new_n14382,
    new_n14383, new_n14384, new_n14385, new_n14386, new_n14387, new_n14388,
    new_n14389, new_n14390, new_n14391, new_n14392, new_n14393, new_n14394,
    new_n14395, new_n14396, new_n14397, new_n14398, new_n14399, new_n14400,
    new_n14401, new_n14402, new_n14403, new_n14404, new_n14405, new_n14406,
    new_n14407, new_n14408, new_n14409, new_n14410, new_n14411,
    new_n14412_1, new_n14413, new_n14415, new_n14416, new_n14417,
    new_n14418, new_n14419, new_n14420, new_n14421, new_n14422, new_n14423,
    new_n14424, new_n14425, new_n14426, new_n14427, new_n14428, new_n14429,
    new_n14430, new_n14431, new_n14432, new_n14433, new_n14434, new_n14435,
    new_n14436, new_n14437, new_n14438, new_n14439, new_n14440_1,
    new_n14441, new_n14442, new_n14443, new_n14444, new_n14445, new_n14446,
    new_n14447, new_n14448, new_n14449, new_n14450, new_n14451, new_n14452,
    new_n14453, new_n14454, new_n14455, new_n14456, new_n14457_1,
    new_n14458, new_n14459, new_n14460, new_n14461, new_n14462, new_n14463,
    new_n14464_1, new_n14465, new_n14466, new_n14467, new_n14468,
    new_n14469, new_n14470, new_n14471_1, new_n14472, new_n14473,
    new_n14474, new_n14475_1, new_n14476, new_n14477, new_n14478,
    new_n14481, new_n14482, new_n14483, new_n14484, new_n14485, new_n14486,
    new_n14487, new_n14488, new_n14489, new_n14490, new_n14491, new_n14492,
    new_n14493, new_n14494, new_n14495, new_n14496, new_n14497, new_n14498,
    new_n14499, new_n14500, new_n14501, new_n14502, new_n14503, new_n14504,
    new_n14505, new_n14506, new_n14507, new_n14508, new_n14509,
    new_n14510_1, new_n14511, new_n14512, new_n14513, new_n14514,
    new_n14515, new_n14516, new_n14517, new_n14518, new_n14519, new_n14520,
    new_n14521, new_n14522, new_n14523, new_n14524, new_n14525, new_n14526,
    new_n14527, new_n14528, new_n14529, new_n14530, new_n14531, new_n14532,
    new_n14533, new_n14534, new_n14535, new_n14536, new_n14537, new_n14538,
    new_n14539, new_n14540, new_n14541_1, new_n14542, new_n14543,
    new_n14544, new_n14545, new_n14546_1, new_n14547_1, new_n14548,
    new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554,
    new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560,
    new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566,
    new_n14567, new_n14568, new_n14569, new_n14570_1, new_n14571,
    new_n14572, new_n14573, new_n14574, new_n14575_1, new_n14576_1,
    new_n14577, new_n14578, new_n14579, new_n14580, new_n14581, new_n14582,
    new_n14583, new_n14584, new_n14585, new_n14586, new_n14587, new_n14588,
    new_n14589, new_n14590, new_n14591, new_n14592, new_n14593_1,
    new_n14594, new_n14595, new_n14596, new_n14597, new_n14598, new_n14599,
    new_n14600, new_n14601, new_n14602, new_n14603_1, new_n14604,
    new_n14605, new_n14606, new_n14607, new_n14608, new_n14609, new_n14610,
    new_n14611, new_n14612, new_n14613, new_n14614, new_n14615, new_n14616,
    new_n14617, new_n14618, new_n14619, new_n14620, new_n14621, new_n14622,
    new_n14623, new_n14624, new_n14625, new_n14626, new_n14628, new_n14629,
    new_n14630, new_n14631, new_n14632, new_n14633_1, new_n14634,
    new_n14635, new_n14636_1, new_n14637, new_n14638, new_n14639,
    new_n14640, new_n14641, new_n14642, new_n14643, new_n14644, new_n14645,
    new_n14646, new_n14647, new_n14648, new_n14649, new_n14650, new_n14651,
    new_n14652, new_n14653, new_n14654, new_n14655, new_n14656, new_n14657,
    new_n14658, new_n14659, new_n14660, new_n14661, new_n14662, new_n14663,
    new_n14664, new_n14665, new_n14666, new_n14667, new_n14668, new_n14669,
    new_n14670, new_n14671, new_n14672, new_n14673, new_n14674, new_n14675,
    new_n14676, new_n14677, new_n14678, new_n14679, new_n14680_1,
    new_n14681, new_n14682, new_n14683, new_n14684_1, new_n14685,
    new_n14686, new_n14687, new_n14688, new_n14689, new_n14690, new_n14691,
    new_n14692_1, new_n14693, new_n14694, new_n14695, new_n14696,
    new_n14697, new_n14698, new_n14699, new_n14700, new_n14701_1,
    new_n14702_1, new_n14703, new_n14704_1, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724,
    new_n14725, new_n14726, new_n14727, new_n14728, new_n14729, new_n14730,
    new_n14731, new_n14732, new_n14733, new_n14734_1, new_n14740,
    new_n14743, new_n14744, new_n14745, new_n14747, new_n14748, new_n14749,
    new_n14750, new_n14751, new_n14752, new_n14753, new_n14754, new_n14755,
    new_n14756, new_n14757, new_n14758, new_n14759, new_n14760, new_n14761,
    new_n14762, new_n14763_1, new_n14764, new_n14765, new_n14766,
    new_n14767, new_n14768, new_n14769, new_n14770, new_n14771,
    new_n14772_1, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14780, new_n14781, new_n14782, new_n14783, new_n14784,
    new_n14785, new_n14786, new_n14787, new_n14788, new_n14789,
    new_n14790_1, new_n14791, new_n14792, new_n14793, new_n14794,
    new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14800,
    new_n14801_1, new_n14802, new_n14803, new_n14804, new_n14805,
    new_n14806, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811,
    new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817,
    new_n14818, new_n14819_1, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826_1, new_n14827_1,
    new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833,
    new_n14834, new_n14835, new_n14836, new_n14837, new_n14838,
    new_n14839_1, new_n14840, new_n14841, new_n14842, new_n14843,
    new_n14844, new_n14845, new_n14846, new_n14847, new_n14853, new_n14854,
    new_n14855, new_n14856, new_n14857, new_n14858, new_n14859, new_n14860,
    new_n14861, new_n14862, new_n14863, new_n14864, new_n14865, new_n14866,
    new_n14867, new_n14868, new_n14869, new_n14870, new_n14871, new_n14872,
    new_n14873, new_n14874, new_n14875, new_n14876, new_n14877, new_n14878,
    new_n14879, new_n14880, new_n14881, new_n14882, new_n14883, new_n14884,
    new_n14885, new_n14886, new_n14887, new_n14888, new_n14889, new_n14890,
    new_n14891_1, new_n14892, new_n14893, new_n14894, new_n14895,
    new_n14896, new_n14897, new_n14898, new_n14899_1, new_n14900,
    new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906,
    new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912,
    new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918,
    new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924,
    new_n14925, new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931_1, new_n14932, new_n14933, new_n14934, new_n14935,
    new_n14936, new_n14937, new_n14938, new_n14939, new_n14940, new_n14941,
    new_n14942, new_n14943, new_n14944_1, new_n14945, new_n14946,
    new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952,
    new_n14953, new_n14954_1, new_n14955, new_n14956, new_n14957,
    new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963,
    new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969,
    new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975,
    new_n14976, new_n14977_1, new_n14978, new_n14979, new_n14982,
    new_n14983, new_n14984, new_n14985, new_n14986, new_n14987, new_n14988,
    new_n14989_1, new_n14990, new_n14991, new_n14992, new_n14993,
    new_n14994, new_n14995, new_n14996, new_n14997, new_n14998, new_n14999,
    new_n15000, new_n15001, new_n15002_1, new_n15003, new_n15004_1,
    new_n15005, new_n15006, new_n15007, new_n15008, new_n15009, new_n15010,
    new_n15011_1, new_n15012, new_n15013, new_n15014, new_n15015,
    new_n15016, new_n15017, new_n15018, new_n15019_1, new_n15020,
    new_n15021, new_n15022, new_n15023, new_n15024, new_n15025, new_n15026,
    new_n15027, new_n15028, new_n15029, new_n15030, new_n15031_1,
    new_n15032, new_n15033_1, new_n15034, new_n15035, new_n15036,
    new_n15037, new_n15038, new_n15039, new_n15040, new_n15041, new_n15042,
    new_n15044, new_n15045, new_n15046, new_n15047, new_n15048, new_n15049,
    new_n15050, new_n15051, new_n15052_1, new_n15053_1, new_n15054,
    new_n15055, new_n15056, new_n15057, new_n15058, new_n15059, new_n15060,
    new_n15061, new_n15062, new_n15063, new_n15064, new_n15065, new_n15066,
    new_n15067, new_n15068, new_n15069, new_n15070, new_n15071, new_n15072,
    new_n15073, new_n15074, new_n15075, new_n15076, new_n15079, new_n15080,
    new_n15081, new_n15082_1, new_n15083, new_n15084, new_n15085,
    new_n15086, new_n15087, new_n15088, new_n15089, new_n15090, new_n15091,
    new_n15092, new_n15093, new_n15094_1, new_n15095, new_n15096,
    new_n15097, new_n15098, new_n15099, new_n15100, new_n15101, new_n15102,
    new_n15103, new_n15104, new_n15105, new_n15106, new_n15107, new_n15108,
    new_n15109, new_n15110, new_n15111, new_n15112, new_n15113, new_n15114,
    new_n15115, new_n15116, new_n15117, new_n15118_1, new_n15119,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128_1, new_n15129, new_n15130, new_n15131,
    new_n15132, new_n15133, new_n15134, new_n15135, new_n15136, new_n15137,
    new_n15138, new_n15139_1, new_n15140, new_n15141, new_n15142,
    new_n15143, new_n15144, new_n15145_1, new_n15146_1, new_n15147,
    new_n15148, new_n15149, new_n15150, new_n15151, new_n15152, new_n15153,
    new_n15154, new_n15155, new_n15156, new_n15157, new_n15158, new_n15159,
    new_n15161, new_n15162, new_n15163, new_n15164, new_n15165_1,
    new_n15166, new_n15167_1, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175,
    new_n15176_1, new_n15177, new_n15178, new_n15179, new_n15180_1,
    new_n15181, new_n15182_1, new_n15183, new_n15184, new_n15185,
    new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191,
    new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197,
    new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203,
    new_n15204, new_n15205_1, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230_1, new_n15231,
    new_n15232, new_n15233, new_n15234, new_n15235, new_n15236, new_n15237,
    new_n15238, new_n15239, new_n15240, new_n15241_1, new_n15242,
    new_n15243, new_n15244, new_n15245, new_n15246, new_n15247, new_n15248,
    new_n15249, new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15255_1, new_n15256, new_n15257, new_n15258_1, new_n15259,
    new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265,
    new_n15266, new_n15267, new_n15268, new_n15269, new_n15270,
    new_n15271_1, new_n15272, new_n15273, new_n15274, new_n15275_1,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289_1, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300_1, new_n15301, new_n15302, new_n15303,
    new_n15304, new_n15305, new_n15306, new_n15307_1, new_n15308,
    new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314,
    new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320,
    new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326,
    new_n15327_1, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332_1, new_n15333, new_n15334, new_n15335, new_n15336,
    new_n15337, new_n15338, new_n15341, new_n15344, new_n15345_1,
    new_n15346, new_n15347, new_n15348, new_n15349, new_n15350, new_n15351,
    new_n15352, new_n15353_1, new_n15354, new_n15355, new_n15356,
    new_n15357, new_n15360, new_n15361, new_n15362, new_n15363, new_n15364,
    new_n15365, new_n15366_1, new_n15367, new_n15368, new_n15369,
    new_n15370, new_n15371, new_n15372, new_n15373, new_n15374, new_n15375,
    new_n15376, new_n15377, new_n15378_1, new_n15379, new_n15380,
    new_n15381, new_n15382_1, new_n15383, new_n15384, new_n15385,
    new_n15386, new_n15387, new_n15388, new_n15389, new_n15390, new_n15391,
    new_n15392, new_n15393, new_n15394, new_n15395, new_n15396, new_n15397,
    new_n15398, new_n15399, new_n15400, new_n15401, new_n15402, new_n15403,
    new_n15404, new_n15405, new_n15406, new_n15407_1, new_n15408,
    new_n15409, new_n15410, new_n15411, new_n15412, new_n15413, new_n15414,
    new_n15415, new_n15416, new_n15417, new_n15418, new_n15419, new_n15420,
    new_n15421, new_n15422, new_n15423, new_n15424_1, new_n15425,
    new_n15426, new_n15427, new_n15428_1, new_n15429, new_n15430,
    new_n15431, new_n15432, new_n15433, new_n15434, new_n15435_1,
    new_n15436, new_n15437, new_n15438_1, new_n15439, new_n15440,
    new_n15441, new_n15442, new_n15443, new_n15444, new_n15445, new_n15446,
    new_n15447, new_n15448, new_n15449, new_n15450, new_n15451, new_n15452,
    new_n15453, new_n15454, new_n15455, new_n15458, new_n15459, new_n15460,
    new_n15461, new_n15462, new_n15463, new_n15464, new_n15465_1,
    new_n15466, new_n15467_1, new_n15468, new_n15469, new_n15470_1,
    new_n15471, new_n15472, new_n15473, new_n15474, new_n15475, new_n15476,
    new_n15477_1, new_n15478, new_n15479, new_n15480, new_n15482,
    new_n15483, new_n15484, new_n15485, new_n15486, new_n15487, new_n15488,
    new_n15489, new_n15490_1, new_n15491, new_n15492, new_n15493,
    new_n15494, new_n15495, new_n15496_1, new_n15497, new_n15498,
    new_n15499, new_n15500, new_n15501_1, new_n15502, new_n15505,
    new_n15506_1, new_n15507, new_n15508_1, new_n15509, new_n15510,
    new_n15511, new_n15512, new_n15513, new_n15514, new_n15515, new_n15516,
    new_n15517, new_n15518, new_n15519, new_n15520, new_n15521, new_n15522,
    new_n15523, new_n15524, new_n15525, new_n15526, new_n15527, new_n15528,
    new_n15529, new_n15530, new_n15531, new_n15532, new_n15533, new_n15534,
    new_n15535, new_n15536, new_n15537, new_n15538, new_n15539_1,
    new_n15540, new_n15541, new_n15543, new_n15544, new_n15545,
    new_n15546_1, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555_1,
    new_n15556, new_n15557, new_n15558_1, new_n15559_1, new_n15560,
    new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566,
    new_n15567, new_n15568, new_n15569, new_n15570_1, new_n15571,
    new_n15572, new_n15573_1, new_n15574, new_n15575, new_n15576,
    new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582,
    new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588_1, new_n15589, new_n15590_1, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597,
    new_n15598_1, new_n15599, new_n15600, new_n15601, new_n15602_1,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613,
    new_n15614_1, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635,
    new_n15636_1, new_n15637, new_n15638, new_n15639, new_n15640,
    new_n15641, new_n15642, new_n15643, new_n15644, new_n15645, new_n15646,
    new_n15647, new_n15648, new_n15649, new_n15650, new_n15651,
    new_n15652_1, new_n15653, new_n15654, new_n15655, new_n15656,
    new_n15657, new_n15658, new_n15659, new_n15660, new_n15661,
    new_n15662_1, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714,
    new_n15715, new_n15717, new_n15718, new_n15719, new_n15720, new_n15721,
    new_n15722, new_n15723, new_n15724, new_n15725, new_n15726, new_n15727,
    new_n15728, new_n15729, new_n15730, new_n15731, new_n15732, new_n15733,
    new_n15734, new_n15735, new_n15736, new_n15737, new_n15738, new_n15739,
    new_n15740, new_n15741, new_n15742, new_n15743_1, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749_1,
    new_n15750, new_n15751, new_n15752, new_n15753, new_n15754, new_n15755,
    new_n15756, new_n15757, new_n15758, new_n15759, new_n15760,
    new_n15761_1, new_n15762_1, new_n15763, new_n15764, new_n15765,
    new_n15766_1, new_n15767, new_n15768, new_n15769, new_n15770,
    new_n15771, new_n15772, new_n15773, new_n15774, new_n15775, new_n15776,
    new_n15777, new_n15778, new_n15779, new_n15780_1, new_n15781,
    new_n15782, new_n15783, new_n15784, new_n15785, new_n15786, new_n15787,
    new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793_1, new_n15794, new_n15795, new_n15796, new_n15797,
    new_n15798, new_n15799, new_n15800, new_n15801, new_n15802, new_n15803,
    new_n15804, new_n15805, new_n15806, new_n15807, new_n15808, new_n15809,
    new_n15810, new_n15811, new_n15812_1, new_n15813, new_n15814,
    new_n15815_1, new_n15816_1, new_n15817, new_n15818, new_n15821,
    new_n15822, new_n15823, new_n15824, new_n15825, new_n15826, new_n15827,
    new_n15828, new_n15829, new_n15830, new_n15831_1, new_n15832,
    new_n15833, new_n15834, new_n15835, new_n15836, new_n15837, new_n15838,
    new_n15839, new_n15840, new_n15841, new_n15842, new_n15843, new_n15844,
    new_n15845, new_n15846_1, new_n15847, new_n15848, new_n15849,
    new_n15850, new_n15851, new_n15852, new_n15853, new_n15854, new_n15855,
    new_n15856, new_n15857, new_n15858, new_n15859_1, new_n15860,
    new_n15861, new_n15862, new_n15863, new_n15864, new_n15865, new_n15866,
    new_n15867, new_n15868, new_n15869_1, new_n15870, new_n15871,
    new_n15872, new_n15873, new_n15874, new_n15875, new_n15876, new_n15877,
    new_n15878, new_n15879, new_n15880, new_n15881, new_n15882, new_n15883,
    new_n15884_1, new_n15885_1, new_n15886, new_n15887, new_n15888,
    new_n15889_1, new_n15890, new_n15891, new_n15892, new_n15893,
    new_n15894, new_n15895, new_n15896, new_n15897, new_n15898, new_n15899,
    new_n15900, new_n15901, new_n15902, new_n15903, new_n15904, new_n15905,
    new_n15906, new_n15907, new_n15908, new_n15909, new_n15910, new_n15911,
    new_n15912, new_n15913, new_n15914, new_n15915, new_n15916,
    new_n15917_1, new_n15918_1, new_n15919, new_n15920, new_n15921,
    new_n15922_1, new_n15923, new_n15925, new_n15926, new_n15927,
    new_n15928, new_n15929, new_n15930, new_n15931, new_n15932, new_n15933,
    new_n15934, new_n15935, new_n15936_1, new_n15937, new_n15938,
    new_n15939, new_n15940, new_n15941, new_n15942, new_n15943, new_n15944,
    new_n15945, new_n15946, new_n15947_1, new_n15948, new_n15949,
    new_n15950, new_n15951, new_n15952, new_n15953, new_n15954, new_n15955,
    new_n15956_1, new_n15957, new_n15958_1, new_n15959, new_n15960,
    new_n15961, new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967_1, new_n15968, new_n15969, new_n15970, new_n15971,
    new_n15972, new_n15973, new_n15974, new_n15975, new_n15977, new_n15978,
    new_n15979_1, new_n15980, new_n15981, new_n15982, new_n15983,
    new_n15984, new_n15985, new_n15986_1, new_n15987, new_n15988,
    new_n15989, new_n15990, new_n15991, new_n15992, new_n15993, new_n15994,
    new_n15995, new_n15996, new_n15997, new_n15998, new_n16001, new_n16002,
    new_n16003, new_n16004, new_n16005, new_n16006, new_n16007, new_n16008,
    new_n16009, new_n16010, new_n16011, new_n16012, new_n16013_1,
    new_n16014, new_n16015, new_n16016, new_n16017, new_n16018, new_n16019,
    new_n16020, new_n16021, new_n16022, new_n16023, new_n16024, new_n16025,
    new_n16026, new_n16027, new_n16028, new_n16029_1, new_n16030,
    new_n16031, new_n16032, new_n16033, new_n16034, new_n16035, new_n16036,
    new_n16037, new_n16038, new_n16039, new_n16040, new_n16041, new_n16042,
    new_n16043, new_n16044, new_n16045, new_n16046, new_n16047, new_n16048,
    new_n16049, new_n16050, new_n16051, new_n16052, new_n16053, new_n16054,
    new_n16055, new_n16056, new_n16057, new_n16058, new_n16059,
    new_n16060_1, new_n16061, new_n16062_1, new_n16063, new_n16064,
    new_n16065, new_n16066, new_n16067, new_n16068_1, new_n16069,
    new_n16070, new_n16071, new_n16072, new_n16073, new_n16074, new_n16075,
    new_n16076, new_n16077, new_n16081, new_n16082, new_n16083, new_n16084,
    new_n16085, new_n16086, new_n16087, new_n16088, new_n16089, new_n16090,
    new_n16091, new_n16095, new_n16096, new_n16097, new_n16098_1,
    new_n16099, new_n16100, new_n16101, new_n16102, new_n16103, new_n16104,
    new_n16105, new_n16106, new_n16107, new_n16108, new_n16109,
    new_n16110_1, new_n16111, new_n16112, new_n16113, new_n16114,
    new_n16115, new_n16116, new_n16117, new_n16118, new_n16119, new_n16122,
    new_n16123, new_n16124, new_n16125, new_n16126, new_n16127, new_n16128,
    new_n16129, new_n16130, new_n16131, new_n16132, new_n16133, new_n16134,
    new_n16135, new_n16136, new_n16137, new_n16138, new_n16139, new_n16140,
    new_n16141, new_n16142_1, new_n16143, new_n16144, new_n16145,
    new_n16146, new_n16147, new_n16148, new_n16149, new_n16150, new_n16151,
    new_n16152, new_n16153, new_n16154, new_n16155, new_n16156, new_n16157,
    new_n16158_1, new_n16159, new_n16160, new_n16161, new_n16162,
    new_n16163, new_n16164, new_n16165, new_n16166, new_n16167_1,
    new_n16168, new_n16169, new_n16170, new_n16171, new_n16172, new_n16173,
    new_n16174, new_n16175, new_n16176, new_n16177, new_n16178, new_n16179,
    new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185_1, new_n16186, new_n16187, new_n16188, new_n16189,
    new_n16190, new_n16191, new_n16192, new_n16193, new_n16194, new_n16195,
    new_n16196_1, new_n16197, new_n16198, new_n16199, new_n16200,
    new_n16201, new_n16202, new_n16203, new_n16204, new_n16205,
    new_n16206_1, new_n16207, new_n16208, new_n16209, new_n16210,
    new_n16211, new_n16212, new_n16213, new_n16214, new_n16215_1,
    new_n16216, new_n16217_1, new_n16218_1, new_n16219_1, new_n16220,
    new_n16221, new_n16222, new_n16223_1, new_n16224, new_n16225,
    new_n16229, new_n16230_1, new_n16231, new_n16232, new_n16233,
    new_n16234, new_n16235, new_n16236, new_n16237, new_n16238, new_n16239,
    new_n16240, new_n16241, new_n16242, new_n16243_1, new_n16244,
    new_n16245, new_n16246, new_n16247_1, new_n16248, new_n16249,
    new_n16250, new_n16251, new_n16252, new_n16253, new_n16254, new_n16255,
    new_n16256, new_n16257, new_n16258, new_n16259, new_n16260, new_n16261,
    new_n16262, new_n16263, new_n16264, new_n16265, new_n16266, new_n16267,
    new_n16268, new_n16269, new_n16270, new_n16271, new_n16272, new_n16273,
    new_n16274, new_n16275_1, new_n16276, new_n16277, new_n16278,
    new_n16279_1, new_n16280, new_n16281, new_n16282, new_n16283,
    new_n16284, new_n16285, new_n16286, new_n16287, new_n16288, new_n16289,
    new_n16290, new_n16291, new_n16292, new_n16293, new_n16294, new_n16295,
    new_n16296, new_n16297, new_n16298, new_n16299, new_n16300, new_n16301,
    new_n16302, new_n16303, new_n16304, new_n16305, new_n16306, new_n16307,
    new_n16308, new_n16309, new_n16310, new_n16311, new_n16312, new_n16313,
    new_n16314, new_n16315, new_n16316, new_n16317, new_n16318, new_n16319,
    new_n16320, new_n16321, new_n16322_1, new_n16323, new_n16324,
    new_n16325, new_n16326, new_n16327_1, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350_1, new_n16351, new_n16352,
    new_n16353, new_n16354, new_n16355, new_n16356, new_n16357, new_n16358,
    new_n16359, new_n16360, new_n16361, new_n16362, new_n16363, new_n16365,
    new_n16366, new_n16367_1, new_n16368, new_n16369, new_n16370,
    new_n16371, new_n16372, new_n16373, new_n16374, new_n16375, new_n16377,
    new_n16378, new_n16379_1, new_n16380, new_n16381, new_n16382,
    new_n16383, new_n16384, new_n16385, new_n16386, new_n16387, new_n16388,
    new_n16389, new_n16390, new_n16391, new_n16392, new_n16393, new_n16394,
    new_n16395, new_n16396_1, new_n16397, new_n16398_1, new_n16399,
    new_n16400, new_n16401, new_n16402, new_n16403, new_n16404, new_n16405,
    new_n16406_1, new_n16407_1, new_n16408, new_n16409, new_n16410,
    new_n16411, new_n16412, new_n16413, new_n16414, new_n16416, new_n16417,
    new_n16418, new_n16419_1, new_n16420, new_n16421, new_n16422,
    new_n16423, new_n16424_1, new_n16425, new_n16426, new_n16427,
    new_n16428_1, new_n16429, new_n16430, new_n16431, new_n16432,
    new_n16433_1, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439_1, new_n16440_1, new_n16441, new_n16442,
    new_n16443, new_n16444, new_n16445_1, new_n16446, new_n16447,
    new_n16448, new_n16449, new_n16450, new_n16451, new_n16452, new_n16454,
    new_n16455, new_n16456, new_n16457, new_n16458, new_n16459,
    new_n16460_1, new_n16461, new_n16462, new_n16463, new_n16464,
    new_n16465, new_n16466, new_n16467, new_n16468, new_n16469, new_n16470,
    new_n16471, new_n16472, new_n16473, new_n16474, new_n16475,
    new_n16476_1, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481_1, new_n16482_1, new_n16483, new_n16484, new_n16485,
    new_n16488, new_n16489, new_n16490, new_n16491, new_n16492,
    new_n16493_1, new_n16494, new_n16495, new_n16496, new_n16497,
    new_n16498, new_n16499, new_n16500, new_n16501, new_n16502_1,
    new_n16503, new_n16504, new_n16505, new_n16506_1, new_n16507_1,
    new_n16508, new_n16509, new_n16510, new_n16511, new_n16512, new_n16513,
    new_n16515, new_n16516_1, new_n16517_1, new_n16518, new_n16519,
    new_n16520, new_n16521_1, new_n16522, new_n16523, new_n16524_1,
    new_n16525, new_n16526, new_n16527_1, new_n16528, new_n16529,
    new_n16530, new_n16531, new_n16532, new_n16533, new_n16534, new_n16535,
    new_n16536, new_n16537, new_n16538, new_n16539, new_n16540, new_n16541,
    new_n16542, new_n16543, new_n16544_1, new_n16545, new_n16546,
    new_n16547, new_n16548, new_n16549, new_n16550, new_n16551, new_n16552,
    new_n16553, new_n16554_1, new_n16555, new_n16556, new_n16557,
    new_n16558, new_n16559, new_n16560, new_n16561, new_n16562, new_n16563,
    new_n16564, new_n16565, new_n16566, new_n16567, new_n16568, new_n16569,
    new_n16570, new_n16571, new_n16572, new_n16573, new_n16574, new_n16575,
    new_n16576, new_n16577, new_n16578, new_n16579, new_n16580, new_n16581,
    new_n16583_1, new_n16584_1, new_n16585, new_n16586, new_n16587,
    new_n16588, new_n16589_1, new_n16590, new_n16591, new_n16592,
    new_n16593, new_n16594, new_n16595, new_n16596_1, new_n16597,
    new_n16598, new_n16599, new_n16600, new_n16601, new_n16602, new_n16603,
    new_n16604, new_n16605, new_n16606, new_n16607, new_n16608_1,
    new_n16609, new_n16610, new_n16611, new_n16612, new_n16613, new_n16614,
    new_n16615, new_n16616, new_n16617_1, new_n16618, new_n16619,
    new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16626, new_n16627, new_n16628, new_n16629, new_n16630_1,
    new_n16631, new_n16632, new_n16633, new_n16634, new_n16635, new_n16636,
    new_n16637, new_n16638, new_n16639, new_n16640_1, new_n16641,
    new_n16642, new_n16643, new_n16644, new_n16645, new_n16646, new_n16647,
    new_n16648, new_n16649, new_n16650, new_n16651, new_n16652, new_n16653,
    new_n16654, new_n16655, new_n16656_1, new_n16657, new_n16658,
    new_n16659, new_n16660, new_n16661, new_n16662, new_n16663, new_n16664,
    new_n16665, new_n16666, new_n16667, new_n16668, new_n16669, new_n16670,
    new_n16671, new_n16672, new_n16673, new_n16674_1, new_n16675,
    new_n16676, new_n16677, new_n16678, new_n16679, new_n16680, new_n16681,
    new_n16682_1, new_n16683, new_n16684_1, new_n16685, new_n16686,
    new_n16687, new_n16688_1, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697,
    new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703,
    new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709,
    new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715,
    new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722_1, new_n16723, new_n16724, new_n16725, new_n16726,
    new_n16727, new_n16728, new_n16729, new_n16730, new_n16731, new_n16732,
    new_n16733_1, new_n16734, new_n16735, new_n16736, new_n16737,
    new_n16738, new_n16739, new_n16741, new_n16742, new_n16743_1,
    new_n16744, new_n16745, new_n16746, new_n16747, new_n16748, new_n16749,
    new_n16750, new_n16751, new_n16752, new_n16753, new_n16754, new_n16755,
    new_n16758, new_n16759, new_n16760, new_n16761, new_n16762, new_n16763,
    new_n16764, new_n16765, new_n16766, new_n16767, new_n16772, new_n16773,
    new_n16774, new_n16775, new_n16776, new_n16777, new_n16778, new_n16779,
    new_n16780, new_n16781, new_n16782, new_n16783, new_n16790, new_n16791,
    new_n16792, new_n16793, new_n16794, new_n16795, new_n16796, new_n16797,
    new_n16798_1, new_n16799, new_n16800, new_n16801, new_n16802,
    new_n16803, new_n16804, new_n16805, new_n16806, new_n16807, new_n16808,
    new_n16809, new_n16810, new_n16811, new_n16812_1, new_n16813,
    new_n16814, new_n16815, new_n16816, new_n16817, new_n16818_1,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823,
    new_n16824_1, new_n16825, new_n16826, new_n16827, new_n16828,
    new_n16829, new_n16830, new_n16831, new_n16832, new_n16833,
    new_n16834_1, new_n16835, new_n16836, new_n16837_1, new_n16838,
    new_n16839, new_n16840, new_n16841_1, new_n16842, new_n16843,
    new_n16844, new_n16845, new_n16846, new_n16847, new_n16848, new_n16849,
    new_n16850, new_n16851, new_n16852, new_n16853, new_n16854, new_n16855,
    new_n16856, new_n16857, new_n16858, new_n16859, new_n16860, new_n16861,
    new_n16862, new_n16863, new_n16864, new_n16865, new_n16866, new_n16867,
    new_n16868, new_n16869, new_n16870, new_n16871, new_n16872, new_n16873,
    new_n16874, new_n16875, new_n16876, new_n16877, new_n16878, new_n16879,
    new_n16880, new_n16881, new_n16883, new_n16884, new_n16885_1,
    new_n16886, new_n16887, new_n16888, new_n16889, new_n16890, new_n16891,
    new_n16892, new_n16893, new_n16894, new_n16895, new_n16896, new_n16897,
    new_n16898, new_n16899, new_n16900, new_n16901, new_n16902, new_n16903,
    new_n16904, new_n16905_1, new_n16906, new_n16907, new_n16908,
    new_n16909, new_n16910, new_n16911_1, new_n16912, new_n16913,
    new_n16914, new_n16915, new_n16916, new_n16917, new_n16918, new_n16919,
    new_n16920, new_n16921, new_n16922, new_n16923, new_n16924, new_n16925,
    new_n16926, new_n16927, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951_1, new_n16952, new_n16953, new_n16954_1, new_n16955,
    new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961,
    new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967,
    new_n16968_1, new_n16969, new_n16970, new_n16971_1, new_n16972,
    new_n16973, new_n16974, new_n16975, new_n16976, new_n16977, new_n16978,
    new_n16979, new_n16980, new_n16981, new_n16982, new_n16983, new_n16984,
    new_n16985, new_n16986, new_n16987, new_n16988_1, new_n16989_1,
    new_n16990, new_n16991, new_n16992, new_n16993, new_n16994_1,
    new_n16995, new_n16996, new_n16997, new_n16998, new_n16999, new_n17000,
    new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006_1, new_n17007, new_n17008, new_n17009, new_n17010,
    new_n17011, new_n17012, new_n17013, new_n17014, new_n17015, new_n17016,
    new_n17017, new_n17018, new_n17019, new_n17020, new_n17021, new_n17022,
    new_n17023, new_n17024, new_n17025, new_n17026, new_n17027, new_n17028,
    new_n17029, new_n17030, new_n17031, new_n17032, new_n17033, new_n17034,
    new_n17035_1, new_n17036, new_n17037_1, new_n17038, new_n17039,
    new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17045,
    new_n17046, new_n17047, new_n17048, new_n17049, new_n17050, new_n17051,
    new_n17052, new_n17053, new_n17054, new_n17055, new_n17056, new_n17057,
    new_n17058, new_n17059, new_n17060, new_n17061, new_n17062, new_n17063,
    new_n17064, new_n17065, new_n17066, new_n17067, new_n17068_1,
    new_n17069_1, new_n17070_1, new_n17071, new_n17072, new_n17073,
    new_n17074, new_n17075_1, new_n17076, new_n17077_1, new_n17078,
    new_n17079, new_n17080, new_n17082, new_n17083, new_n17084_1,
    new_n17085, new_n17086, new_n17087, new_n17088, new_n17089,
    new_n17090_1, new_n17091, new_n17092, new_n17093, new_n17094,
    new_n17095_1, new_n17096, new_n17097, new_n17098, new_n17099,
    new_n17100, new_n17101, new_n17102, new_n17103, new_n17104_1,
    new_n17105, new_n17106_1, new_n17107, new_n17108, new_n17109,
    new_n17110, new_n17111, new_n17112, new_n17113, new_n17114, new_n17115,
    new_n17116, new_n17117, new_n17118, new_n17119_1, new_n17120,
    new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126,
    new_n17127, new_n17128, new_n17131, new_n17132, new_n17133, new_n17134,
    new_n17135, new_n17136, new_n17137, new_n17138_1, new_n17139,
    new_n17140, new_n17141, new_n17142, new_n17143, new_n17144, new_n17145,
    new_n17146, new_n17149, new_n17150, new_n17151, new_n17152, new_n17153,
    new_n17154, new_n17155, new_n17156, new_n17157, new_n17161, new_n17162,
    new_n17163_1, new_n17164, new_n17165, new_n17166, new_n17167,
    new_n17168_1, new_n17169, new_n17170, new_n17171, new_n17172,
    new_n17173, new_n17174, new_n17175, new_n17176, new_n17177, new_n17178,
    new_n17179, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184,
    new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190,
    new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196,
    new_n17197, new_n17198, new_n17199, new_n17200, new_n17201,
    new_n17202_1, new_n17203, new_n17204, new_n17207, new_n17208,
    new_n17209, new_n17210, new_n17211, new_n17212, new_n17213, new_n17214,
    new_n17215, new_n17216, new_n17217, new_n17218, new_n17219_1,
    new_n17220, new_n17221, new_n17222, new_n17223, new_n17224, new_n17225,
    new_n17226, new_n17227, new_n17228, new_n17229, new_n17230, new_n17231,
    new_n17232_1, new_n17233, new_n17234, new_n17235, new_n17236_1,
    new_n17237, new_n17238, new_n17239, new_n17240, new_n17241, new_n17242,
    new_n17243_1, new_n17244, new_n17245, new_n17246, new_n17247,
    new_n17248, new_n17249, new_n17250_1, new_n17251_1, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263_1,
    new_n17264, new_n17265, new_n17266, new_n17267, new_n17268, new_n17269,
    new_n17270, new_n17271, new_n17272, new_n17273, new_n17274, new_n17275,
    new_n17276, new_n17277, new_n17278, new_n17279, new_n17280, new_n17281,
    new_n17282, new_n17283, new_n17284, new_n17285_1, new_n17286,
    new_n17287, new_n17288, new_n17289, new_n17290, new_n17291, new_n17293,
    new_n17294, new_n17295, new_n17296, new_n17297, new_n17298, new_n17299,
    new_n17300, new_n17301, new_n17302_1, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320_1, new_n17321,
    new_n17322, new_n17323, new_n17324, new_n17325, new_n17326, new_n17327,
    new_n17328, new_n17329, new_n17331, new_n17332, new_n17333, new_n17334,
    new_n17335, new_n17336, new_n17337_1, new_n17338, new_n17339,
    new_n17340, new_n17341, new_n17342, new_n17343, new_n17344_1,
    new_n17345, new_n17346, new_n17347, new_n17348, new_n17349, new_n17350,
    new_n17351_1, new_n17352, new_n17353, new_n17354, new_n17355,
    new_n17356, new_n17357, new_n17358, new_n17359_1, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366,
    new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372,
    new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378,
    new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384,
    new_n17385, new_n17386, new_n17387_1, new_n17388, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418,
    new_n17419, new_n17420, new_n17421_1, new_n17422, new_n17423,
    new_n17424, new_n17425, new_n17426, new_n17427, new_n17428, new_n17429,
    new_n17430, new_n17431, new_n17432_1, new_n17433, new_n17434,
    new_n17435, new_n17436_1, new_n17437, new_n17438, new_n17439,
    new_n17440_1, new_n17441, new_n17442, new_n17443, new_n17444,
    new_n17445, new_n17446, new_n17447, new_n17448, new_n17449,
    new_n17450_1, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17460, new_n17461_1,
    new_n17462, new_n17463, new_n17464, new_n17465, new_n17466_1,
    new_n17467, new_n17468, new_n17469, new_n17470, new_n17471, new_n17472,
    new_n17473, new_n17474, new_n17475, new_n17476, new_n17477, new_n17478,
    new_n17479, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484,
    new_n17485, new_n17488, new_n17489, new_n17490, new_n17491, new_n17492,
    new_n17493_1, new_n17494, new_n17495, new_n17496, new_n17497,
    new_n17498, new_n17499, new_n17500_1, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17509,
    new_n17514, new_n17515, new_n17516, new_n17517, new_n17518, new_n17519,
    new_n17520, new_n17521, new_n17522, new_n17523, new_n17524_1,
    new_n17525, new_n17526, new_n17527, new_n17528, new_n17529_1,
    new_n17530, new_n17531, new_n17532, new_n17533, new_n17534, new_n17535,
    new_n17536, new_n17537, new_n17538, new_n17539, new_n17540, new_n17541,
    new_n17542, new_n17543, new_n17544, new_n17545, new_n17546, new_n17547,
    new_n17548, new_n17549, new_n17550, new_n17551, new_n17552, new_n17553,
    new_n17554, new_n17555, new_n17556, new_n17557_1, new_n17558,
    new_n17559, new_n17560, new_n17561, new_n17562, new_n17563, new_n17564,
    new_n17565, new_n17566, new_n17567, new_n17568, new_n17569, new_n17570,
    new_n17571, new_n17572, new_n17573, new_n17574, new_n17575, new_n17576,
    new_n17577, new_n17578, new_n17579, new_n17580, new_n17581, new_n17582,
    new_n17583_1, new_n17584, new_n17585, new_n17586, new_n17587,
    new_n17588, new_n17589, new_n17590, new_n17591, new_n17592_1,
    new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17598,
    new_n17599, new_n17600, new_n17601, new_n17602, new_n17603, new_n17604,
    new_n17605, new_n17606, new_n17607, new_n17608, new_n17609, new_n17610,
    new_n17611, new_n17612, new_n17613, new_n17614, new_n17615, new_n17616,
    new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17625,
    new_n17626, new_n17627, new_n17628, new_n17629, new_n17630, new_n17631,
    new_n17632, new_n17633, new_n17634, new_n17635, new_n17636, new_n17637,
    new_n17638_1, new_n17639, new_n17640, new_n17641, new_n17642,
    new_n17643, new_n17644, new_n17645, new_n17646, new_n17647, new_n17648,
    new_n17649, new_n17650, new_n17651, new_n17658, new_n17659, new_n17660,
    new_n17661, new_n17662, new_n17663, new_n17664_1, new_n17665,
    new_n17666, new_n17667, new_n17668, new_n17669, new_n17670, new_n17671,
    new_n17672, new_n17673, new_n17674, new_n17675, new_n17676, new_n17677,
    new_n17678, new_n17679, new_n17680, new_n17681, new_n17682, new_n17683,
    new_n17684, new_n17685, new_n17686, new_n17687_1, new_n17688,
    new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694,
    new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700,
    new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706,
    new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712,
    new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718,
    new_n17719, new_n17720, new_n17721_1, new_n17722, new_n17723,
    new_n17724, new_n17725, new_n17726, new_n17727, new_n17728, new_n17729,
    new_n17732, new_n17733, new_n17734, new_n17735_1, new_n17736,
    new_n17737, new_n17738_1, new_n17739, new_n17740, new_n17741,
    new_n17742, new_n17743, new_n17744, new_n17745, new_n17746_1,
    new_n17747, new_n17748, new_n17749_1, new_n17750, new_n17751,
    new_n17752, new_n17753, new_n17754, new_n17755, new_n17756, new_n17757,
    new_n17758, new_n17759, new_n17760, new_n17761, new_n17762, new_n17763,
    new_n17764, new_n17765, new_n17766, new_n17767, new_n17768, new_n17769,
    new_n17770, new_n17771, new_n17772, new_n17773, new_n17774, new_n17775,
    new_n17776, new_n17777, new_n17778, new_n17779, new_n17780, new_n17781,
    new_n17782, new_n17783, new_n17784_1, new_n17785, new_n17786,
    new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792,
    new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798,
    new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17806, new_n17808, new_n17809, new_n17810, new_n17811,
    new_n17812, new_n17813, new_n17814, new_n17815, new_n17816, new_n17817,
    new_n17818, new_n17819, new_n17820_1, new_n17821, new_n17822,
    new_n17823, new_n17824, new_n17825, new_n17826, new_n17827, new_n17828,
    new_n17829, new_n17830, new_n17831, new_n17832, new_n17833, new_n17834,
    new_n17835, new_n17836, new_n17837, new_n17838, new_n17839, new_n17840,
    new_n17841, new_n17842, new_n17843, new_n17844, new_n17845, new_n17846,
    new_n17847, new_n17848, new_n17849, new_n17850, new_n17851, new_n17852,
    new_n17853, new_n17854, new_n17855_1, new_n17856, new_n17857,
    new_n17858, new_n17859, new_n17861, new_n17862, new_n17863, new_n17864,
    new_n17865, new_n17866, new_n17867, new_n17868, new_n17869, new_n17870,
    new_n17871, new_n17872, new_n17873, new_n17874, new_n17875, new_n17876,
    new_n17877_1, new_n17878, new_n17879, new_n17880, new_n17881,
    new_n17882, new_n17883, new_n17884, new_n17885, new_n17886, new_n17887,
    new_n17888, new_n17889_1, new_n17890, new_n17891, new_n17892,
    new_n17893, new_n17894, new_n17895, new_n17896, new_n17897, new_n17898,
    new_n17899, new_n17900, new_n17901, new_n17902, new_n17903, new_n17908,
    new_n17909, new_n17910, new_n17911_1, new_n17912_1, new_n17913,
    new_n17914, new_n17915, new_n17916, new_n17917, new_n17918, new_n17919,
    new_n17920, new_n17921, new_n17922, new_n17923, new_n17928, new_n17929,
    new_n17930, new_n17931_1, new_n17932, new_n17933, new_n17934,
    new_n17935, new_n17936, new_n17937, new_n17938, new_n17939, new_n17940,
    new_n17941, new_n17942, new_n17943, new_n17944, new_n17945, new_n17946,
    new_n17947, new_n17948_1, new_n17949, new_n17950, new_n17951,
    new_n17952, new_n17953, new_n17954_1, new_n17955, new_n17956_1,
    new_n17957, new_n17958, new_n17959_1, new_n17960, new_n17961,
    new_n17962, new_n17963_1, new_n17964, new_n17965, new_n17966,
    new_n17967, new_n17968_1, new_n17969, new_n17970, new_n17971,
    new_n17972, new_n17973, new_n17974, new_n17976_1, new_n17977,
    new_n17978, new_n17979, new_n17981, new_n17982, new_n17983, new_n17984,
    new_n17985, new_n17986, new_n17987, new_n17988, new_n17989, new_n17990,
    new_n17991, new_n17992, new_n17996, new_n17997, new_n17998_1,
    new_n17999, new_n18000, new_n18001, new_n18002, new_n18003, new_n18004,
    new_n18005, new_n18006, new_n18007, new_n18008, new_n18009, new_n18010,
    new_n18011, new_n18012, new_n18013, new_n18015, new_n18016, new_n18017,
    new_n18018, new_n18019, new_n18020, new_n18021, new_n18022, new_n18023,
    new_n18024, new_n18025_1, new_n18026, new_n18027, new_n18028,
    new_n18029, new_n18030, new_n18031, new_n18032, new_n18033, new_n18034,
    new_n18035_1, new_n18036, new_n18037, new_n18038, new_n18039,
    new_n18040, new_n18041, new_n18042, new_n18043_1, new_n18044,
    new_n18045_1, new_n18046, new_n18047, new_n18048, new_n18049,
    new_n18050, new_n18051, new_n18052, new_n18053, new_n18054, new_n18055,
    new_n18056, new_n18057, new_n18058, new_n18059_1, new_n18060,
    new_n18061_1, new_n18062, new_n18063, new_n18064, new_n18065,
    new_n18066, new_n18067, new_n18068, new_n18069, new_n18070,
    new_n18071_1, new_n18072, new_n18073, new_n18074, new_n18075,
    new_n18076, new_n18077, new_n18079, new_n18080, new_n18081, new_n18082,
    new_n18083, new_n18084, new_n18085, new_n18086, new_n18087, new_n18088,
    new_n18090, new_n18091, new_n18092, new_n18093, new_n18094, new_n18095,
    new_n18096, new_n18097, new_n18098, new_n18099, new_n18100, new_n18101,
    new_n18102, new_n18103, new_n18104, new_n18105_1, new_n18106,
    new_n18107, new_n18108, new_n18109, new_n18110, new_n18111, new_n18112,
    new_n18113, new_n18114, new_n18115, new_n18116, new_n18117, new_n18118,
    new_n18119, new_n18120, new_n18121, new_n18122, new_n18123, new_n18124,
    new_n18125, new_n18126, new_n18127, new_n18128, new_n18129, new_n18130,
    new_n18131, new_n18132, new_n18133, new_n18134, new_n18135, new_n18136,
    new_n18137, new_n18138, new_n18139, new_n18140, new_n18141, new_n18142,
    new_n18143_1, new_n18144, new_n18145_1, new_n18146, new_n18147,
    new_n18148, new_n18149, new_n18150, new_n18151_1, new_n18152_1,
    new_n18153, new_n18154, new_n18155, new_n18156, new_n18157_1,
    new_n18158, new_n18159, new_n18160, new_n18161, new_n18162, new_n18163,
    new_n18164, new_n18165, new_n18166, new_n18167, new_n18168, new_n18169,
    new_n18170, new_n18171_1, new_n18172, new_n18173, new_n18174,
    new_n18175, new_n18176, new_n18177, new_n18178, new_n18179, new_n18180,
    new_n18181, new_n18182, new_n18183, new_n18184, new_n18185, new_n18186,
    new_n18187, new_n18188, new_n18189, new_n18190, new_n18191, new_n18192,
    new_n18193_1, new_n18194, new_n18195, new_n18196, new_n18197,
    new_n18198, new_n18199, new_n18200, new_n18201, new_n18202, new_n18203,
    new_n18204, new_n18205, new_n18206, new_n18207, new_n18208, new_n18209,
    new_n18210, new_n18211, new_n18212, new_n18213, new_n18214, new_n18215,
    new_n18216, new_n18217, new_n18218, new_n18219, new_n18220, new_n18221,
    new_n18222, new_n18223, new_n18224, new_n18225, new_n18226,
    new_n18227_1, new_n18228, new_n18229, new_n18230, new_n18231,
    new_n18232_1, new_n18233, new_n18234, new_n18235, new_n18236,
    new_n18237, new_n18238_1, new_n18239, new_n18240, new_n18241_1,
    new_n18242, new_n18243, new_n18244, new_n18245, new_n18246, new_n18247,
    new_n18248, new_n18249, new_n18250, new_n18251, new_n18252, new_n18253,
    new_n18254_1, new_n18255, new_n18256, new_n18257, new_n18258,
    new_n18259, new_n18260, new_n18261, new_n18262, new_n18263, new_n18264,
    new_n18265, new_n18266, new_n18267, new_n18268, new_n18269, new_n18270,
    new_n18271, new_n18272, new_n18273, new_n18274_1, new_n18275,
    new_n18276, new_n18277, new_n18278, new_n18279, new_n18280, new_n18281,
    new_n18282, new_n18283, new_n18284, new_n18287, new_n18288_1,
    new_n18289, new_n18290_1, new_n18291, new_n18292, new_n18293,
    new_n18294, new_n18295_1, new_n18296, new_n18297, new_n18298,
    new_n18299, new_n18300, new_n18301_1, new_n18302, new_n18303,
    new_n18304_1, new_n18305, new_n18306, new_n18307, new_n18308,
    new_n18309, new_n18310_1, new_n18311_1, new_n18312, new_n18313,
    new_n18315, new_n18316, new_n18317, new_n18318, new_n18319, new_n18320,
    new_n18321, new_n18322, new_n18323_1, new_n18324, new_n18325,
    new_n18326, new_n18327, new_n18328, new_n18329, new_n18330, new_n18331,
    new_n18332_1, new_n18333, new_n18336, new_n18337, new_n18338,
    new_n18339, new_n18340, new_n18341, new_n18346, new_n18347, new_n18348,
    new_n18349, new_n18350_1, new_n18351, new_n18352, new_n18353,
    new_n18354, new_n18355, new_n18356, new_n18357, new_n18358, new_n18359,
    new_n18360, new_n18361, new_n18362_1, new_n18363, new_n18364,
    new_n18365, new_n18366, new_n18367, new_n18368, new_n18369, new_n18370,
    new_n18371, new_n18372, new_n18373, new_n18374, new_n18375, new_n18376,
    new_n18377_1, new_n18378, new_n18379, new_n18380, new_n18381,
    new_n18382, new_n18383, new_n18384, new_n18385, new_n18386, new_n18387,
    new_n18388, new_n18389, new_n18390, new_n18391, new_n18392, new_n18393,
    new_n18394, new_n18395, new_n18396, new_n18397, new_n18398, new_n18399,
    new_n18400, new_n18401, new_n18402, new_n18403, new_n18404,
    new_n18405_1, new_n18406, new_n18407, new_n18408, new_n18409_1,
    new_n18410, new_n18411, new_n18412, new_n18413, new_n18414_1,
    new_n18415, new_n18416, new_n18417, new_n18418_1, new_n18419,
    new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425,
    new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431,
    new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437_1, new_n18438, new_n18439_1, new_n18440, new_n18441,
    new_n18442, new_n18443, new_n18444_1, new_n18445_1, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451, new_n18454,
    new_n18455, new_n18456, new_n18457, new_n18458, new_n18459, new_n18460,
    new_n18461, new_n18462, new_n18463, new_n18464, new_n18465, new_n18466,
    new_n18467_1, new_n18468, new_n18469, new_n18471, new_n18472,
    new_n18473, new_n18474, new_n18475, new_n18476, new_n18477, new_n18478,
    new_n18479, new_n18480, new_n18481, new_n18482_1, new_n18483_1,
    new_n18484, new_n18485, new_n18486, new_n18487, new_n18488, new_n18489,
    new_n18490, new_n18491, new_n18492, new_n18493, new_n18494, new_n18495,
    new_n18496_1, new_n18497, new_n18498, new_n18499, new_n18500,
    new_n18501, new_n18502, new_n18503, new_n18504, new_n18505, new_n18506,
    new_n18507, new_n18508, new_n18509_1, new_n18510, new_n18511,
    new_n18512, new_n18513_1, new_n18514, new_n18515_1, new_n18516,
    new_n18517, new_n18518, new_n18521, new_n18522, new_n18523, new_n18524,
    new_n18525, new_n18526, new_n18527, new_n18528, new_n18529, new_n18530,
    new_n18531, new_n18532, new_n18533, new_n18534, new_n18535, new_n18536,
    new_n18537_1, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18556, new_n18557, new_n18558_1, new_n18559,
    new_n18560, new_n18561, new_n18562, new_n18563, new_n18564, new_n18565,
    new_n18566, new_n18567, new_n18568, new_n18569, new_n18570, new_n18571,
    new_n18572_1, new_n18573, new_n18574_1, new_n18575, new_n18576_1,
    new_n18577, new_n18578_1, new_n18579, new_n18580, new_n18581,
    new_n18582_1, new_n18583_1, new_n18584_1, new_n18585, new_n18586,
    new_n18587, new_n18588, new_n18589, new_n18590, new_n18595, new_n18596,
    new_n18597, new_n18598, new_n18599, new_n18600, new_n18601, new_n18602,
    new_n18603, new_n18604, new_n18605, new_n18606, new_n18607, new_n18608,
    new_n18609, new_n18610_1, new_n18611, new_n18612, new_n18613,
    new_n18618, new_n18619, new_n18620, new_n18621, new_n18622, new_n18623,
    new_n18624, new_n18625, new_n18626, new_n18627, new_n18628, new_n18629,
    new_n18630, new_n18631, new_n18632, new_n18633, new_n18634,
    new_n18635_1, new_n18636, new_n18637, new_n18638, new_n18639,
    new_n18640, new_n18641, new_n18642, new_n18643, new_n18644, new_n18645,
    new_n18646, new_n18647, new_n18648, new_n18649_1, new_n18650,
    new_n18651, new_n18652, new_n18653_1, new_n18654, new_n18655,
    new_n18656, new_n18657, new_n18658, new_n18659, new_n18660, new_n18661,
    new_n18662, new_n18663, new_n18664, new_n18665, new_n18666, new_n18667,
    new_n18668, new_n18669, new_n18670, new_n18671, new_n18672, new_n18673,
    new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679_1, new_n18680, new_n18681, new_n18682, new_n18683,
    new_n18684, new_n18685, new_n18686, new_n18687, new_n18688, new_n18689,
    new_n18690_1, new_n18691, new_n18692, new_n18693_1, new_n18694,
    new_n18695, new_n18701, new_n18702, new_n18703, new_n18704, new_n18705,
    new_n18706, new_n18707, new_n18708_1, new_n18709, new_n18710,
    new_n18711, new_n18712, new_n18713, new_n18714, new_n18715, new_n18716,
    new_n18717, new_n18719, new_n18720, new_n18721_1, new_n18722,
    new_n18723, new_n18724, new_n18725_1, new_n18726, new_n18727,
    new_n18728, new_n18729, new_n18730, new_n18731, new_n18732, new_n18733,
    new_n18734, new_n18735, new_n18736, new_n18737_1, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745_1, new_n18746, new_n18747, new_n18748, new_n18749,
    new_n18750, new_n18751_1, new_n18752, new_n18753, new_n18754,
    new_n18755, new_n18756, new_n18757, new_n18758, new_n18759, new_n18760,
    new_n18761, new_n18762, new_n18763, new_n18764, new_n18765, new_n18766,
    new_n18767, new_n18768, new_n18769, new_n18770, new_n18771, new_n18772,
    new_n18773, new_n18774, new_n18775, new_n18776, new_n18777, new_n18778,
    new_n18779, new_n18780_1, new_n18781, new_n18782_1, new_n18783,
    new_n18784, new_n18785, new_n18786, new_n18787, new_n18788, new_n18789,
    new_n18790, new_n18791, new_n18796, new_n18797, new_n18798, new_n18799,
    new_n18800, new_n18801, new_n18802_1, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822,
    new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828,
    new_n18829, new_n18830_1, new_n18831_1, new_n18832, new_n18833,
    new_n18834, new_n18835, new_n18836, new_n18837, new_n18838, new_n18839,
    new_n18840, new_n18841, new_n18842, new_n18843_1, new_n18844,
    new_n18845, new_n18846, new_n18847, new_n18848, new_n18849, new_n18850,
    new_n18851, new_n18852, new_n18853, new_n18854, new_n18855, new_n18856,
    new_n18857, new_n18858_1, new_n18859_1, new_n18860, new_n18863,
    new_n18864_1, new_n18865_1, new_n18866, new_n18867, new_n18868,
    new_n18869, new_n18870, new_n18871, new_n18872, new_n18873, new_n18874,
    new_n18875, new_n18876, new_n18877, new_n18878, new_n18879,
    new_n18880_1, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18885, new_n18886_1, new_n18887_1, new_n18888, new_n18889,
    new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895,
    new_n18896, new_n18897, new_n18898, new_n18899, new_n18900,
    new_n18901_1, new_n18902, new_n18903, new_n18904, new_n18905,
    new_n18906, new_n18907_1, new_n18908, new_n18909, new_n18910,
    new_n18911, new_n18912, new_n18913, new_n18914, new_n18915, new_n18916,
    new_n18917, new_n18918, new_n18919_1, new_n18920, new_n18921,
    new_n18922, new_n18923, new_n18924, new_n18925, new_n18928, new_n18929,
    new_n18930, new_n18931, new_n18932, new_n18933, new_n18934, new_n18935,
    new_n18936, new_n18937, new_n18938, new_n18939, new_n18940_1,
    new_n18941, new_n18942, new_n18943, new_n18944, new_n18946, new_n18947,
    new_n18948, new_n18949, new_n18950, new_n18951, new_n18952, new_n18953,
    new_n18954, new_n18955, new_n18956, new_n18957, new_n18958, new_n18959,
    new_n18960, new_n18961, new_n18962_1, new_n18963, new_n18964,
    new_n18965, new_n18967, new_n18968, new_n18969, new_n18970_1,
    new_n18971, new_n18972, new_n18973, new_n18974, new_n18975, new_n18976,
    new_n18977_1, new_n18978, new_n18979, new_n18980, new_n18981,
    new_n18982_1, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999_1, new_n19000, new_n19001, new_n19002, new_n19003,
    new_n19004, new_n19005_1, new_n19006, new_n19007, new_n19011,
    new_n19012, new_n19013, new_n19014, new_n19015, new_n19016, new_n19017,
    new_n19018, new_n19019, new_n19020, new_n19021, new_n19022, new_n19023,
    new_n19024, new_n19025, new_n19026, new_n19027, new_n19028, new_n19029,
    new_n19030, new_n19031, new_n19032, new_n19033_1, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042_1, new_n19043, new_n19044_1, new_n19045,
    new_n19046, new_n19047, new_n19048, new_n19049, new_n19050, new_n19051,
    new_n19052, new_n19053, new_n19054, new_n19055, new_n19056, new_n19057,
    new_n19058, new_n19059, new_n19061, new_n19062, new_n19063, new_n19064,
    new_n19065, new_n19066, new_n19067, new_n19068, new_n19069, new_n19070,
    new_n19071, new_n19072, new_n19073, new_n19074, new_n19075, new_n19076,
    new_n19077, new_n19078, new_n19079, new_n19080, new_n19081_1,
    new_n19082, new_n19083, new_n19084, new_n19085, new_n19086, new_n19087,
    new_n19088, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19110,
    new_n19111, new_n19112, new_n19113, new_n19114, new_n19115,
    new_n19116_1, new_n19117, new_n19118, new_n19121, new_n19122,
    new_n19123, new_n19124, new_n19125_1, new_n19126, new_n19127,
    new_n19128, new_n19129, new_n19130, new_n19131, new_n19132, new_n19133,
    new_n19134, new_n19135, new_n19136, new_n19137, new_n19138, new_n19139,
    new_n19140, new_n19141_1, new_n19142, new_n19143, new_n19144_1,
    new_n19145, new_n19146, new_n19147, new_n19148, new_n19149, new_n19150,
    new_n19151, new_n19152, new_n19153, new_n19154, new_n19155, new_n19156,
    new_n19157, new_n19158, new_n19159, new_n19160, new_n19161, new_n19162,
    new_n19163_1, new_n19164_1, new_n19165, new_n19166, new_n19167,
    new_n19168, new_n19169, new_n19170, new_n19171, new_n19172, new_n19173,
    new_n19174_1, new_n19175, new_n19176_1, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19191, new_n19192, new_n19193, new_n19194,
    new_n19195, new_n19196_1, new_n19197, new_n19198, new_n19199,
    new_n19200, new_n19201, new_n19202_1, new_n19203, new_n19204,
    new_n19205, new_n19206, new_n19207, new_n19208, new_n19209, new_n19210,
    new_n19211, new_n19212, new_n19216, new_n19217, new_n19218, new_n19219,
    new_n19220_1, new_n19221_1, new_n19222, new_n19223_1, new_n19224_1,
    new_n19225, new_n19226, new_n19227, new_n19228_1, new_n19229,
    new_n19230, new_n19231, new_n19232, new_n19233_1, new_n19234_1,
    new_n19235, new_n19236, new_n19237, new_n19238, new_n19239, new_n19240,
    new_n19241, new_n19242, new_n19243, new_n19244_1, new_n19245,
    new_n19246, new_n19247, new_n19248, new_n19249, new_n19250, new_n19251,
    new_n19252, new_n19253, new_n19254, new_n19255, new_n19256, new_n19257,
    new_n19258, new_n19259, new_n19260, new_n19261, new_n19262, new_n19263,
    new_n19264, new_n19265, new_n19266, new_n19267, new_n19268, new_n19269,
    new_n19270_1, new_n19271, new_n19272, new_n19273, new_n19274,
    new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280,
    new_n19281, new_n19282_1, new_n19283, new_n19284, new_n19285,
    new_n19286, new_n19287, new_n19288, new_n19289, new_n19290, new_n19291,
    new_n19292, new_n19293, new_n19294, new_n19295, new_n19296, new_n19297,
    new_n19298, new_n19299, new_n19300, new_n19301, new_n19302, new_n19303,
    new_n19304, new_n19305, new_n19306, new_n19307, new_n19308, new_n19309,
    new_n19310, new_n19318, new_n19319, new_n19320, new_n19321, new_n19322,
    new_n19323_1, new_n19324, new_n19325, new_n19326, new_n19327_1,
    new_n19328, new_n19329, new_n19330, new_n19331, new_n19332,
    new_n19333_1, new_n19334, new_n19335, new_n19336, new_n19337,
    new_n19338, new_n19339, new_n19340, new_n19341, new_n19342, new_n19343,
    new_n19344, new_n19345, new_n19346, new_n19347, new_n19348_1,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353,
    new_n19354_1, new_n19355, new_n19356, new_n19357_1, new_n19358,
    new_n19359, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367_1, new_n19368, new_n19369, new_n19370, new_n19371,
    new_n19372, new_n19373, new_n19374, new_n19375, new_n19376, new_n19377,
    new_n19378, new_n19379, new_n19380, new_n19381, new_n19382, new_n19383,
    new_n19384, new_n19385_1, new_n19386, new_n19387, new_n19388,
    new_n19389_1, new_n19390, new_n19391, new_n19392, new_n19393,
    new_n19394, new_n19395, new_n19396, new_n19397, new_n19398, new_n19399,
    new_n19400, new_n19401_1, new_n19402, new_n19403, new_n19404,
    new_n19405, new_n19406, new_n19407, new_n19408, new_n19409, new_n19410,
    new_n19411, new_n19412, new_n19413, new_n19414_1, new_n19415,
    new_n19416, new_n19417, new_n19418, new_n19419, new_n19420, new_n19421,
    new_n19422, new_n19423, new_n19424_1, new_n19425, new_n19426,
    new_n19427, new_n19428, new_n19429, new_n19430, new_n19431, new_n19432,
    new_n19433, new_n19434, new_n19435, new_n19436, new_n19437, new_n19438,
    new_n19439, new_n19440, new_n19441, new_n19442, new_n19443, new_n19444,
    new_n19445, new_n19446, new_n19447, new_n19448, new_n19449,
    new_n19450_1, new_n19451, new_n19452, new_n19453, new_n19454_1,
    new_n19455, new_n19457, new_n19458_1, new_n19459, new_n19460,
    new_n19461, new_n19462, new_n19463, new_n19464, new_n19465, new_n19466,
    new_n19470, new_n19471, new_n19472_1, new_n19473, new_n19474,
    new_n19475, new_n19476, new_n19477_1, new_n19478, new_n19479,
    new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485,
    new_n19486, new_n19487, new_n19488, new_n19489, new_n19490, new_n19491,
    new_n19492, new_n19494_1, new_n19495, new_n19496_1, new_n19497,
    new_n19498, new_n19499, new_n19500, new_n19501, new_n19502, new_n19503,
    new_n19504, new_n19505, new_n19506, new_n19507, new_n19508, new_n19509,
    new_n19510, new_n19511, new_n19512, new_n19513, new_n19514_1,
    new_n19515_1, new_n19516, new_n19517, new_n19518, new_n19519,
    new_n19520, new_n19521, new_n19522, new_n19523_1, new_n19524,
    new_n19525, new_n19526, new_n19527, new_n19528, new_n19529, new_n19530,
    new_n19531_1, new_n19532, new_n19533, new_n19534, new_n19535,
    new_n19536, new_n19537, new_n19538, new_n19539_1, new_n19540,
    new_n19541, new_n19542, new_n19543, new_n19544, new_n19545, new_n19546,
    new_n19547, new_n19548, new_n19549, new_n19550, new_n19551, new_n19552,
    new_n19553, new_n19554, new_n19555, new_n19556, new_n19557, new_n19558,
    new_n19559, new_n19560, new_n19561, new_n19562, new_n19564, new_n19567,
    new_n19568, new_n19569, new_n19570_1, new_n19571, new_n19572,
    new_n19573, new_n19574, new_n19575_1, new_n19576, new_n19577,
    new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584_1, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602_1, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608_1, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617_1, new_n19618_1, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623_1, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641_1, new_n19642, new_n19643,
    new_n19644, new_n19645, new_n19646, new_n19647, new_n19648_1,
    new_n19649, new_n19650, new_n19651, new_n19652_1, new_n19653,
    new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659,
    new_n19660, new_n19661, new_n19662, new_n19663, new_n19664_1,
    new_n19665, new_n19668, new_n19669, new_n19670, new_n19671, new_n19672,
    new_n19673, new_n19674, new_n19675, new_n19676, new_n19677, new_n19678,
    new_n19679, new_n19680_1, new_n19681, new_n19682, new_n19683,
    new_n19684, new_n19685, new_n19686, new_n19687, new_n19688, new_n19689,
    new_n19690, new_n19691, new_n19692, new_n19693, new_n19694, new_n19695,
    new_n19696, new_n19697, new_n19698, new_n19699, new_n19700,
    new_n19701_1, new_n19702, new_n19703, new_n19704, new_n19705,
    new_n19706, new_n19707, new_n19708, new_n19709, new_n19710, new_n19711,
    new_n19712, new_n19713, new_n19714, new_n19715, new_n19716, new_n19717,
    new_n19718, new_n19719, new_n19720, new_n19721, new_n19722, new_n19723,
    new_n19724, new_n19725, new_n19726, new_n19727, new_n19728, new_n19729,
    new_n19730, new_n19731, new_n19732, new_n19733, new_n19740, new_n19741,
    new_n19742, new_n19746, new_n19747, new_n19748, new_n19749_1,
    new_n19750, new_n19751, new_n19752, new_n19753, new_n19754, new_n19755,
    new_n19756_1, new_n19757, new_n19758, new_n19759, new_n19760,
    new_n19761, new_n19762, new_n19763, new_n19764, new_n19765, new_n19766,
    new_n19767_1, new_n19768, new_n19769, new_n19770_1, new_n19771,
    new_n19772, new_n19773, new_n19774, new_n19775, new_n19776, new_n19777,
    new_n19778, new_n19779, new_n19780_1, new_n19781, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789_1, new_n19790, new_n19791, new_n19792_1, new_n19793,
    new_n19794, new_n19795, new_n19796, new_n19797, new_n19798_1,
    new_n19799, new_n19800, new_n19801, new_n19802, new_n19803_1,
    new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809,
    new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815,
    new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821,
    new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827,
    new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833,
    new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839,
    new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845,
    new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851,
    new_n19852, new_n19853, new_n19854, new_n19855, new_n19856, new_n19857,
    new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863,
    new_n19864, new_n19865, new_n19866, new_n19867, new_n19868, new_n19869,
    new_n19870, new_n19871, new_n19872, new_n19873_1, new_n19874,
    new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19882,
    new_n19883, new_n19884, new_n19885, new_n19886, new_n19887, new_n19888,
    new_n19889, new_n19890, new_n19891, new_n19892, new_n19893, new_n19894,
    new_n19895, new_n19896, new_n19897, new_n19898, new_n19899, new_n19900,
    new_n19901, new_n19902, new_n19903, new_n19904, new_n19905_1,
    new_n19906, new_n19907, new_n19908, new_n19909_1, new_n19910,
    new_n19911_1, new_n19912, new_n19913, new_n19914, new_n19915,
    new_n19916_1, new_n19917, new_n19918, new_n19919, new_n19920,
    new_n19921, new_n19922_1, new_n19923_1, new_n19924, new_n19925,
    new_n19926, new_n19927, new_n19928, new_n19929, new_n19930_1,
    new_n19931, new_n19932, new_n19933, new_n19934, new_n19935, new_n19936,
    new_n19937, new_n19938, new_n19939, new_n19940, new_n19941_1,
    new_n19942, new_n19943, new_n19944, new_n19945, new_n19946, new_n19947,
    new_n19948, new_n19949, new_n19950, new_n19951, new_n19952, new_n19953,
    new_n19954, new_n19955, new_n19956, new_n19957, new_n19958, new_n19959,
    new_n19960, new_n19961, new_n19962, new_n19963, new_n19964, new_n19965,
    new_n19966, new_n19967, new_n19968_1, new_n19969, new_n19970,
    new_n19971, new_n19972, new_n19977, new_n19978, new_n19979, new_n19980,
    new_n19981, new_n19982, new_n19983, new_n19984, new_n19985, new_n19986,
    new_n19987, new_n19988_1, new_n19989, new_n19990, new_n19991,
    new_n19992, new_n19993, new_n19994, new_n19995, new_n19996, new_n19997,
    new_n19998, new_n19999, new_n20000, new_n20001, new_n20002, new_n20003,
    new_n20004_1, new_n20005, new_n20006, new_n20007, new_n20008,
    new_n20009, new_n20010, new_n20011, new_n20012, new_n20013_1,
    new_n20014, new_n20015, new_n20016, new_n20017_1, new_n20018,
    new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024,
    new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030,
    new_n20031, new_n20032, new_n20033_1, new_n20034, new_n20035,
    new_n20036_1, new_n20037, new_n20038, new_n20039, new_n20040_1,
    new_n20041, new_n20042, new_n20043, new_n20044, new_n20045, new_n20046,
    new_n20047, new_n20048, new_n20049, new_n20050, new_n20051, new_n20052,
    new_n20053, new_n20054, new_n20055, new_n20056, new_n20057, new_n20058,
    new_n20059, new_n20060, new_n20061_1, new_n20062, new_n20063,
    new_n20064, new_n20065, new_n20066, new_n20067, new_n20068,
    new_n20069_1, new_n20071, new_n20072, new_n20073, new_n20074,
    new_n20075, new_n20076, new_n20077_1, new_n20078, new_n20080,
    new_n20081, new_n20082, new_n20083, new_n20084, new_n20085,
    new_n20086_1, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095,
    new_n20096_1, new_n20097, new_n20098, new_n20099, new_n20100,
    new_n20101, new_n20102, new_n20103_1, new_n20104, new_n20105,
    new_n20106, new_n20113, new_n20114, new_n20115, new_n20116, new_n20117,
    new_n20118, new_n20119, new_n20120, new_n20121, new_n20122, new_n20123,
    new_n20124, new_n20125, new_n20126_1, new_n20127, new_n20128,
    new_n20129, new_n20132, new_n20142, new_n20143, new_n20144, new_n20145,
    new_n20146, new_n20147, new_n20148, new_n20149_1, new_n20150,
    new_n20151_1, new_n20152, new_n20153, new_n20154, new_n20155,
    new_n20156, new_n20157, new_n20158, new_n20159, new_n20160, new_n20161,
    new_n20162, new_n20163, new_n20164, new_n20165, new_n20166, new_n20167,
    new_n20168, new_n20169_1, new_n20170, new_n20171, new_n20172,
    new_n20173, new_n20174, new_n20175, new_n20176, new_n20177, new_n20178,
    new_n20179_1, new_n20180, new_n20181, new_n20182, new_n20183,
    new_n20185, new_n20186, new_n20187_1, new_n20188, new_n20189,
    new_n20190, new_n20191, new_n20192, new_n20193, new_n20194, new_n20195,
    new_n20196, new_n20197, new_n20198, new_n20199, new_n20200, new_n20201,
    new_n20202, new_n20203, new_n20204, new_n20205, new_n20206, new_n20207,
    new_n20208, new_n20209, new_n20210, new_n20211, new_n20212, new_n20214,
    new_n20215, new_n20216, new_n20217, new_n20218, new_n20219, new_n20220,
    new_n20221, new_n20222, new_n20223, new_n20224, new_n20225, new_n20226,
    new_n20227, new_n20228, new_n20229, new_n20230, new_n20231, new_n20232,
    new_n20233, new_n20234, new_n20235_1, new_n20236, new_n20237,
    new_n20238, new_n20239, new_n20240, new_n20241, new_n20242, new_n20243,
    new_n20244, new_n20245, new_n20246, new_n20247, new_n20248, new_n20249,
    new_n20250_1, new_n20251, new_n20252, new_n20253, new_n20254,
    new_n20255, new_n20256, new_n20257, new_n20258, new_n20259_1,
    new_n20260, new_n20261, new_n20262, new_n20263, new_n20264, new_n20265,
    new_n20266, new_n20267, new_n20268, new_n20269, new_n20270, new_n20271,
    new_n20272, new_n20273, new_n20274, new_n20275, new_n20276, new_n20277,
    new_n20278, new_n20279_1, new_n20280, new_n20281, new_n20282,
    new_n20283, new_n20284, new_n20285, new_n20286, new_n20287_1,
    new_n20288, new_n20289, new_n20290, new_n20291, new_n20292, new_n20293,
    new_n20294, new_n20295, new_n20296, new_n20297, new_n20298, new_n20299,
    new_n20300, new_n20301_1, new_n20302, new_n20303, new_n20304,
    new_n20305, new_n20306, new_n20307, new_n20308, new_n20309, new_n20310,
    new_n20311, new_n20312, new_n20313, new_n20314, new_n20315, new_n20316,
    new_n20317, new_n20318, new_n20319, new_n20320, new_n20321, new_n20322,
    new_n20323, new_n20324, new_n20325, new_n20326, new_n20327, new_n20328,
    new_n20329, new_n20330_1, new_n20331, new_n20332, new_n20333_1,
    new_n20334, new_n20335, new_n20336, new_n20337, new_n20338, new_n20339,
    new_n20340, new_n20341, new_n20342, new_n20343, new_n20344, new_n20345,
    new_n20346, new_n20347, new_n20348, new_n20349_1, new_n20350,
    new_n20351, new_n20352, new_n20353, new_n20354, new_n20355_1,
    new_n20356, new_n20357, new_n20358, new_n20359_1, new_n20360,
    new_n20361, new_n20362, new_n20363, new_n20364, new_n20365,
    new_n20366_1, new_n20367, new_n20368, new_n20369, new_n20370,
    new_n20371, new_n20372, new_n20373, new_n20374, new_n20375, new_n20376,
    new_n20377, new_n20378, new_n20379, new_n20380, new_n20381, new_n20382,
    new_n20383, new_n20384, new_n20385_1, new_n20386, new_n20387,
    new_n20392, new_n20393, new_n20394, new_n20395, new_n20396, new_n20397,
    new_n20398, new_n20399, new_n20400, new_n20401, new_n20402_1,
    new_n20403_1, new_n20404, new_n20405, new_n20406, new_n20407,
    new_n20408, new_n20409_1, new_n20410, new_n20411_1, new_n20414,
    new_n20415, new_n20416, new_n20417, new_n20418, new_n20419, new_n20420,
    new_n20421, new_n20422, new_n20423, new_n20424_1, new_n20425,
    new_n20426, new_n20427, new_n20428, new_n20429_1, new_n20430,
    new_n20431, new_n20432, new_n20433, new_n20436_1, new_n20437,
    new_n20438, new_n20439, new_n20440, new_n20441_1, new_n20442,
    new_n20447, new_n20448, new_n20452, new_n20453, new_n20454,
    new_n20455_1, new_n20456, new_n20457, new_n20458, new_n20459,
    new_n20460, new_n20461, new_n20462, new_n20463, new_n20464, new_n20465,
    new_n20466, new_n20467, new_n20468, new_n20472, new_n20473, new_n20474,
    new_n20475, new_n20476, new_n20477, new_n20478_1, new_n20479,
    new_n20480, new_n20482, new_n20483, new_n20484, new_n20485, new_n20486,
    new_n20487, new_n20488, new_n20489_1, new_n20490_1, new_n20491,
    new_n20492, new_n20493, new_n20494, new_n20495_1, new_n20496,
    new_n20497, new_n20498, new_n20499, new_n20501, new_n20502, new_n20503,
    new_n20504, new_n20505, new_n20506, new_n20507, new_n20508, new_n20509,
    new_n20510, new_n20511, new_n20512, new_n20513, new_n20514,
    new_n20515_1, new_n20516, new_n20517, new_n20518, new_n20519,
    new_n20520, new_n20521, new_n20522, new_n20523, new_n20524, new_n20525,
    new_n20526, new_n20527, new_n20528, new_n20529, new_n20530, new_n20531,
    new_n20532, new_n20533_1, new_n20534, new_n20535, new_n20536,
    new_n20538, new_n20539, new_n20540, new_n20541, new_n20542, new_n20543,
    new_n20544, new_n20545, new_n20546, new_n20547, new_n20548, new_n20549,
    new_n20550, new_n20551, new_n20552, new_n20553, new_n20554, new_n20555,
    new_n20556, new_n20557, new_n20558, new_n20559, new_n20560, new_n20561,
    new_n20562, new_n20563, new_n20564, new_n20565, new_n20566, new_n20567,
    new_n20568, new_n20569, new_n20570, new_n20571, new_n20572, new_n20573,
    new_n20574, new_n20575, new_n20576, new_n20577, new_n20578, new_n20579,
    new_n20580, new_n20581, new_n20582_1, new_n20583, new_n20584,
    new_n20585, new_n20586, new_n20587, new_n20588, new_n20589,
    new_n20590_1, new_n20591, new_n20592, new_n20593, new_n20594,
    new_n20595, new_n20596, new_n20597, new_n20598, new_n20599, new_n20600,
    new_n20601, new_n20602_1, new_n20603, new_n20604_1, new_n20605,
    new_n20606, new_n20607, new_n20608, new_n20609_1, new_n20610,
    new_n20611, new_n20612, new_n20613, new_n20614, new_n20615, new_n20616,
    new_n20617, new_n20618, new_n20619, new_n20620, new_n20621, new_n20626,
    new_n20627, new_n20628, new_n20629_1, new_n20630, new_n20631,
    new_n20632, new_n20633, new_n20634, new_n20635, new_n20636, new_n20637,
    new_n20638, new_n20639, new_n20640, new_n20641, new_n20642, new_n20643,
    new_n20644, new_n20645, new_n20646, new_n20647, new_n20648, new_n20649,
    new_n20650, new_n20651, new_n20652, new_n20653, new_n20654, new_n20655,
    new_n20656, new_n20657, new_n20658_1, new_n20659, new_n20660,
    new_n20661_1, new_n20662, new_n20663, new_n20664, new_n20665,
    new_n20666, new_n20667, new_n20668, new_n20669, new_n20670, new_n20671,
    new_n20672, new_n20673_1, new_n20674, new_n20675, new_n20676,
    new_n20677, new_n20678_1, new_n20679, new_n20680_1, new_n20681,
    new_n20682, new_n20683, new_n20684, new_n20685_1, new_n20686,
    new_n20687, new_n20688, new_n20689, new_n20690, new_n20691_1,
    new_n20692, new_n20693, new_n20694, new_n20695, new_n20696_1,
    new_n20697, new_n20698, new_n20699, new_n20700_1, new_n20701,
    new_n20702, new_n20703, new_n20704_1, new_n20705_1, new_n20706,
    new_n20707, new_n20708, new_n20709_1, new_n20710, new_n20711,
    new_n20712, new_n20713_1, new_n20714, new_n20715, new_n20716,
    new_n20717, new_n20718, new_n20719, new_n20720, new_n20721,
    new_n20722_1, new_n20723_1, new_n20724, new_n20725, new_n20726,
    new_n20727, new_n20728, new_n20729, new_n20730, new_n20731, new_n20732,
    new_n20733, new_n20734, new_n20735, new_n20736, new_n20737, new_n20738,
    new_n20739, new_n20740, new_n20742, new_n20743, new_n20748_1,
    new_n20751, new_n20752, new_n20753, new_n20754, new_n20755, new_n20756,
    new_n20757, new_n20758, new_n20759, new_n20760, new_n20761_1,
    new_n20762, new_n20763, new_n20764, new_n20765, new_n20766, new_n20767,
    new_n20768, new_n20769, new_n20770, new_n20771, new_n20772, new_n20773,
    new_n20774_1, new_n20775, new_n20776, new_n20777, new_n20778,
    new_n20779, new_n20780, new_n20781, new_n20782, new_n20783, new_n20784,
    new_n20786, new_n20787, new_n20788_1, new_n20789, new_n20790,
    new_n20791, new_n20792, new_n20793, new_n20794_1, new_n20795_1,
    new_n20796, new_n20797, new_n20798, new_n20799, new_n20800, new_n20801,
    new_n20802, new_n20803_1, new_n20804, new_n20805, new_n20806,
    new_n20807, new_n20808, new_n20809, new_n20810, new_n20811, new_n20812,
    new_n20813, new_n20814, new_n20815, new_n20824, new_n20825,
    new_n20826_1, new_n20827, new_n20828, new_n20829, new_n20830,
    new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20839,
    new_n20840, new_n20841, new_n20842, new_n20843, new_n20844, new_n20845,
    new_n20846, new_n20847, new_n20848, new_n20849, new_n20850, new_n20851,
    new_n20852, new_n20853, new_n20854, new_n20855, new_n20856, new_n20857,
    new_n20858, new_n20859, new_n20860, new_n20861, new_n20862, new_n20863,
    new_n20864, new_n20865, new_n20866, new_n20867, new_n20868,
    new_n20869_1, new_n20872, new_n20873, new_n20874, new_n20875,
    new_n20876, new_n20877, new_n20878, new_n20879_1, new_n20880,
    new_n20881, new_n20882, new_n20883, new_n20884, new_n20885, new_n20886,
    new_n20887, new_n20888, new_n20889, new_n20890, new_n20891, new_n20892,
    new_n20893, new_n20894, new_n20895, new_n20896, new_n20897, new_n20898,
    new_n20899, new_n20900, new_n20901, new_n20902, new_n20903, new_n20904,
    new_n20905, new_n20906, new_n20907, new_n20908, new_n20909, new_n20910,
    new_n20911, new_n20912, new_n20913, new_n20914, new_n20915_1,
    new_n20916, new_n20917, new_n20918, new_n20919, new_n20920, new_n20921,
    new_n20922, new_n20923_1, new_n20924, new_n20925, new_n20926,
    new_n20927, new_n20928, new_n20929_1, new_n20930, new_n20931,
    new_n20932, new_n20933, new_n20934, new_n20936_1, new_n20937,
    new_n20938, new_n20939, new_n20940, new_n20941, new_n20942, new_n20943,
    new_n20944, new_n20945, new_n20946_1, new_n20947, new_n20948,
    new_n20949, new_n20950, new_n20951, new_n20952, new_n20953, new_n20954,
    new_n20955, new_n20956, new_n20957, new_n20958, new_n20959, new_n20960,
    new_n20961, new_n20962, new_n20963, new_n20964, new_n20965, new_n20966,
    new_n20967, new_n20968, new_n20970, new_n20971, new_n20973, new_n20974,
    new_n20975, new_n20976, new_n20977, new_n20978, new_n20979, new_n20980,
    new_n20981, new_n20982, new_n20983, new_n20984, new_n20985,
    new_n20986_1, new_n20987, new_n20988, new_n20989, new_n20990,
    new_n20991, new_n20992, new_n20993, new_n20994, new_n20995, new_n20996,
    new_n20997, new_n20998, new_n20999, new_n21000, new_n21001, new_n21002,
    new_n21003, new_n21004, new_n21005, new_n21006, new_n21007, new_n21010,
    new_n21011, new_n21014, new_n21015, new_n21016, new_n21017_1,
    new_n21018, new_n21019, new_n21020, new_n21021, new_n21022, new_n21023,
    new_n21024, new_n21025, new_n21026, new_n21027, new_n21028, new_n21029,
    new_n21030, new_n21031, new_n21032, new_n21033, new_n21034_1,
    new_n21035, new_n21036, new_n21037, new_n21038, new_n21039, new_n21040,
    new_n21041, new_n21042, new_n21043, new_n21044, new_n21045,
    new_n21046_1, new_n21047, new_n21048, new_n21049, new_n21050,
    new_n21051, new_n21052, new_n21055, new_n21056, new_n21057, new_n21058,
    new_n21059, new_n21060, new_n21061, new_n21062_1, new_n21063,
    new_n21064, new_n21065, new_n21066, new_n21067, new_n21068, new_n21069,
    new_n21070, new_n21071, new_n21072, new_n21073, new_n21074, new_n21075,
    new_n21076, new_n21077, new_n21078_1, new_n21086, new_n21087,
    new_n21088, new_n21089, new_n21090, new_n21091, new_n21092,
    new_n21093_1, new_n21094_1, new_n21095_1, new_n21096, new_n21097,
    new_n21098, new_n21099, new_n21100, new_n21101, new_n21102, new_n21103,
    new_n21104, new_n21105, new_n21106, new_n21107, new_n21108, new_n21109,
    new_n21110, new_n21111, new_n21112, new_n21113, new_n21114, new_n21115,
    new_n21116, new_n21117, new_n21118, new_n21119, new_n21120, new_n21121,
    new_n21122, new_n21123_1, new_n21124, new_n21125, new_n21126,
    new_n21127, new_n21128, new_n21129, new_n21130, new_n21131, new_n21132,
    new_n21133, new_n21134_1, new_n21135, new_n21136, new_n21137,
    new_n21138_1, new_n21139, new_n21140, new_n21141, new_n21142,
    new_n21143, new_n21150, new_n21154_1, new_n21155, new_n21156,
    new_n21157_1, new_n21158, new_n21159, new_n21160, new_n21161,
    new_n21162, new_n21163, new_n21164, new_n21180, new_n21182_1,
    new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193_1,
    new_n21194, new_n21195, new_n21196, new_n21197, new_n21198, new_n21199,
    new_n21200, new_n21201, new_n21202, new_n21203_1, new_n21204,
    new_n21206, new_n21207, new_n21208, new_n21209, new_n21210, new_n21211,
    new_n21212, new_n21213, new_n21214, new_n21215, new_n21216, new_n21217,
    new_n21218, new_n21219, new_n21220, new_n21221, new_n21222_1,
    new_n21223, new_n21224, new_n21226_1, new_n21227, new_n21228,
    new_n21229, new_n21230, new_n21231, new_n21232, new_n21233, new_n21234,
    new_n21235, new_n21236, new_n21237, new_n21238_1, new_n21239,
    new_n21240, new_n21241, new_n21246, new_n21247, new_n21248, new_n21249,
    new_n21250, new_n21251, new_n21252, new_n21253, new_n21254_1,
    new_n21255, new_n21256, new_n21257, new_n21258, new_n21259, new_n21260,
    new_n21261, new_n21262, new_n21263, new_n21264, new_n21267, new_n21274,
    new_n21275, new_n21276_1, new_n21277, new_n21278, new_n21279,
    new_n21280, new_n21286, new_n21287_1, new_n21288, new_n21289,
    new_n21290, new_n21291, new_n21292, new_n21293, new_n21294, new_n21295,
    new_n21300, new_n21306, new_n21307, new_n21308, new_n21309, new_n21310,
    new_n21311, new_n21312, new_n21313, new_n21314, new_n21315, new_n21316,
    new_n21317_1, new_n21318, new_n21319, new_n21320, new_n21321,
    new_n21322, new_n21327, new_n21328, new_n21329, new_n21330, new_n21331,
    new_n21332, new_n21339, new_n21340, new_n21341, new_n21342, new_n21343,
    new_n21344, new_n21345, new_n21346, new_n21347, new_n21348,
    new_n21349_1, new_n21350, new_n21351, new_n21352, new_n21353,
    new_n21354, new_n21355, new_n21356, new_n21357, new_n21358, new_n21359,
    new_n21360, new_n21361, new_n21362, new_n21363, new_n21364,
    new_n21365_1, new_n21366, new_n21367_1, new_n21368, new_n21369,
    new_n21370, new_n21371, new_n21372, new_n21373, new_n21374, new_n21375,
    new_n21376, new_n21377, new_n21378, new_n21379, new_n21380, new_n21381,
    new_n21382, new_n21385, new_n21386, new_n21387, new_n21388, new_n21389,
    new_n21390, new_n21391, new_n21392, new_n21393, new_n21395,
    new_n21396_1, new_n21397, new_n21398_1, new_n21399_1, new_n21400,
    new_n21401, new_n21402, new_n21403, new_n21404_1, new_n21405,
    new_n21406, new_n21407, new_n21408, new_n21409, new_n21410, new_n21411,
    new_n21421, new_n21422, new_n21423, new_n21424, new_n21425, new_n21426,
    new_n21427, new_n21428, new_n21429, new_n21430, new_n21431, new_n21432,
    new_n21433, new_n21434, new_n21435, new_n21436, new_n21437, new_n21438,
    new_n21439, new_n21440, new_n21441, new_n21442, new_n21443, new_n21444,
    new_n21445, new_n21446_1, new_n21447, new_n21448, new_n21449,
    new_n21450, new_n21451, new_n21452, new_n21453, new_n21459, new_n21460,
    new_n21461, new_n21462, new_n21472_1, new_n21473, new_n21474,
    new_n21475, new_n21476, new_n21477, new_n21478, new_n21479, new_n21480,
    new_n21481, new_n21482, new_n21483, new_n21484, new_n21485, new_n21486,
    new_n21487, new_n21488, new_n21489_1, new_n21490, new_n21491,
    new_n21492, new_n21493, new_n21494, new_n21495, new_n21496, new_n21497,
    new_n21498, new_n21499, new_n21500, new_n21501, new_n21502, new_n21503,
    new_n21504, new_n21505, new_n21506, new_n21507, new_n21508, new_n21509,
    new_n21510, new_n21511, new_n21512, new_n21513, new_n21514, new_n21515,
    new_n21516, new_n21517, new_n21518, new_n21519, new_n21520, new_n21521,
    new_n21522, new_n21523, new_n21524, new_n21525_1, new_n21526,
    new_n21527, new_n21528, new_n21529, new_n21530, new_n21531, new_n21532,
    new_n21533, new_n21534, new_n21535, new_n21536, new_n21537,
    new_n21538_1, new_n21539, new_n21540, new_n21541, new_n21542,
    new_n21543, new_n21544, new_n21546, new_n21547, new_n21548,
    new_n21549_1, new_n21550, new_n21551, new_n21552, new_n21553,
    new_n21554, new_n21555, new_n21556, new_n21557, new_n21558, new_n21559,
    new_n21560, new_n21561, new_n21562, new_n21563, new_n21564, new_n21565,
    new_n21566, new_n21567, new_n21568, new_n21569, new_n21570, new_n21571,
    new_n21572, new_n21573, new_n21574, new_n21575, new_n21576, new_n21577,
    new_n21578, new_n21579, new_n21580, new_n21581, new_n21582, new_n21583,
    new_n21584, new_n21585, new_n21586, new_n21587, new_n21588, new_n21589,
    new_n21590, new_n21591, new_n21592, new_n21593, new_n21594, new_n21595,
    new_n21596, new_n21597, new_n21598, new_n21599_1, new_n21600,
    new_n21601, new_n21602, new_n21603, new_n21604, new_n21605, new_n21606,
    new_n21607, new_n21608, new_n21609, new_n21610, new_n21611, new_n21612,
    new_n21613, new_n21614, new_n21617, new_n21618, new_n21619, new_n21620,
    new_n21621, new_n21622, new_n21623, new_n21624, new_n21625, new_n21626,
    new_n21627, new_n21628_1, new_n21629, new_n21635, new_n21636,
    new_n21637_1, new_n21638, new_n21639, new_n21640, new_n21641,
    new_n21642, new_n21643, new_n21644, new_n21645_1, new_n21646,
    new_n21647, new_n21648, new_n21649_1, new_n21650, new_n21651,
    new_n21652, new_n21653, new_n21654_1, new_n21655, new_n21656,
    new_n21657, new_n21658, new_n21659, new_n21660, new_n21661, new_n21662,
    new_n21663, new_n21664, new_n21665_1, new_n21666, new_n21667,
    new_n21668, new_n21669, new_n21670, new_n21671, new_n21672, new_n21673,
    new_n21674_1, new_n21675, new_n21676, new_n21677, new_n21678,
    new_n21679, new_n21680_1, new_n21681, new_n21682, new_n21683,
    new_n21684, new_n21685_1, new_n21686, new_n21687_1, new_n21688,
    new_n21689, new_n21690, new_n21691, new_n21692, new_n21693, new_n21694,
    new_n21695, new_n21696, new_n21697, new_n21698, new_n21699, new_n21700,
    new_n21701, new_n21702, new_n21703, new_n21704, new_n21705, new_n21706,
    new_n21708, new_n21709, new_n21710, new_n21711, new_n21712, new_n21713,
    new_n21714, new_n21715, new_n21716, new_n21717_1, new_n21720,
    new_n21721, new_n21722, new_n21723, new_n21724, new_n21725, new_n21726,
    new_n21727, new_n21728, new_n21729, new_n21735_1, new_n21736,
    new_n21737, new_n21738, new_n21739, new_n21740, new_n21741, new_n21742,
    new_n21743, new_n21744, new_n21745, new_n21746, new_n21747, new_n21748,
    new_n21749_1, new_n21750_1, new_n21751, new_n21752, new_n21753_1,
    new_n21754, new_n21755, new_n21756, new_n21757, new_n21758, new_n21759,
    new_n21760, new_n21761, new_n21762, new_n21763, new_n21764,
    new_n21765_1, new_n21766, new_n21767, new_n21768, new_n21769,
    new_n21770, new_n21771, new_n21772, new_n21773, new_n21774, new_n21775,
    new_n21776, new_n21777, new_n21778, new_n21779_1, new_n21780,
    new_n21781, new_n21782, new_n21783, new_n21784_1, new_n21785,
    new_n21786, new_n21787, new_n21788, new_n21789, new_n21790, new_n21791,
    new_n21792, new_n21793, new_n21794, new_n21795, new_n21796, new_n21797,
    new_n21798, new_n21799, new_n21800_1, new_n21801, new_n21802,
    new_n21810, new_n21811, new_n21812, new_n21813, new_n21814, new_n21819,
    new_n21822, new_n21824, new_n21825, new_n21826, new_n21827, new_n21828,
    new_n21829, new_n21830, new_n21831, new_n21832_1, new_n21833,
    new_n21834, new_n21835, new_n21836, new_n21837, new_n21838,
    new_n21839_1, new_n21840, new_n21841, new_n21842, new_n21843,
    new_n21844, new_n21845, new_n21846, new_n21847, new_n21848, new_n21849,
    new_n21850, new_n21851, new_n21852, new_n21853, new_n21854, new_n21855,
    new_n21856, new_n21857, new_n21858, new_n21859, new_n21860, new_n21861,
    new_n21862, new_n21863, new_n21864, new_n21865, new_n21866, new_n21867,
    new_n21868, new_n21869, new_n21872, new_n21873, new_n21874_1,
    new_n21875, new_n21883, new_n21884, new_n21885, new_n21886, new_n21887,
    new_n21888, new_n21889, new_n21890, new_n21891, new_n21895, new_n21903,
    new_n21904, new_n21905_1, new_n21906, new_n21907, new_n21908,
    new_n21909, new_n21910, new_n21911, new_n21912, new_n21913, new_n21914,
    new_n21915_1, new_n21916, new_n21918, new_n21919, new_n21920,
    new_n21921, new_n21922, new_n21923, new_n21924, new_n21925, new_n21926,
    new_n21927, new_n21928, new_n21929, new_n21930, new_n21931, new_n21932,
    new_n21933, new_n21934_1, new_n21940, new_n21941, new_n21942,
    new_n21943_1, new_n21944, new_n21945, new_n21946, new_n21947,
    new_n21948, new_n21949, new_n21950, new_n21951, new_n21952, new_n21953,
    new_n21954, new_n21955, new_n21956, new_n21957_1, new_n21958,
    new_n21959, new_n21960_1, new_n21961, new_n21962, new_n21963,
    new_n21964, new_n21965, new_n21966, new_n21967, new_n21968, new_n21969,
    new_n21972, new_n21973, new_n21974, new_n21975, new_n21976_1,
    new_n21977, new_n21978, new_n21979, new_n21980, new_n21981_1,
    new_n21982, new_n21983, new_n21984, new_n21985, new_n21986_1,
    new_n21987, new_n21988, new_n21989, new_n21990, new_n21991, new_n21992,
    new_n21993_1, new_n21994, new_n21996, new_n21997_1, new_n21998,
    new_n21999, new_n22000, new_n22001, new_n22002, new_n22003, new_n22004,
    new_n22005, new_n22006, new_n22007, new_n22008, new_n22009, new_n22013,
    new_n22015, new_n22016_1, new_n22021, new_n22022, new_n22023,
    new_n22024, new_n22025, new_n22026, new_n22027_1, new_n22028,
    new_n22029, new_n22030, new_n22031, new_n22032, new_n22033, new_n22034,
    new_n22035, new_n22036, new_n22037, new_n22038, new_n22039, new_n22040,
    new_n22041, new_n22042, new_n22043_1, new_n22044, new_n22045,
    new_n22046, new_n22047, new_n22048, new_n22049, new_n22050_1,
    new_n22051, new_n22052, new_n22053, new_n22054, new_n22055, new_n22056,
    new_n22057, new_n22058, new_n22059, new_n22060, new_n22061, new_n22062,
    new_n22063_1, new_n22064, new_n22065, new_n22067, new_n22068_1,
    new_n22069, new_n22070, new_n22071, new_n22072_1, new_n22073,
    new_n22074, new_n22075, new_n22076_1, new_n22077, new_n22078,
    new_n22079, new_n22080, new_n22081, new_n22082, new_n22083, new_n22084,
    new_n22085, new_n22086, new_n22087, new_n22088, new_n22089,
    new_n22090_1, new_n22091, new_n22092, new_n22093, new_n22094,
    new_n22095, new_n22096, new_n22097, new_n22098, new_n22099, new_n22100,
    new_n22101, new_n22102, new_n22103, new_n22104, new_n22105, new_n22106,
    new_n22107_1, new_n22108, new_n22109, new_n22110, new_n22111,
    new_n22112, new_n22113_1, new_n22114, new_n22115, new_n22116,
    new_n22117, new_n22123, new_n22132, new_n22133, new_n22134, new_n22135,
    new_n22141, new_n22148, new_n22149, new_n22150_1, new_n22151,
    new_n22152, new_n22153, new_n22154, new_n22155, new_n22156,
    new_n22157_1, new_n22158, new_n22159, new_n22160, new_n22161,
    new_n22162, new_n22163, new_n22164, new_n22165, new_n22166, new_n22167,
    new_n22168, new_n22169, new_n22170, new_n22171, new_n22172,
    new_n22173_1, new_n22174, new_n22175, new_n22176, new_n22177,
    new_n22178, new_n22179, new_n22180, new_n22181, new_n22182, new_n22183,
    new_n22184, new_n22187, new_n22188, new_n22189, new_n22190, new_n22191,
    new_n22192, new_n22193, new_n22194, new_n22195, new_n22196, new_n22197,
    new_n22198_1, new_n22205, new_n22206, new_n22207, new_n22208,
    new_n22209, new_n22210, new_n22211, new_n22212, new_n22213_1,
    new_n22214, new_n22215, new_n22216, new_n22217, new_n22218, new_n22219,
    new_n22220, new_n22221, new_n22222, new_n22223, new_n22224, new_n22225,
    new_n22226, new_n22227, new_n22228, new_n22229, new_n22230, new_n22231,
    new_n22232, new_n22233, new_n22234, new_n22235, new_n22236, new_n22237,
    new_n22238, new_n22239, new_n22240, new_n22241, new_n22242, new_n22243,
    new_n22244, new_n22245, new_n22246, new_n22247, new_n22248, new_n22249,
    new_n22250, new_n22251, new_n22252, new_n22253_1, new_n22254,
    new_n22255, new_n22256, new_n22257, new_n22258, new_n22259, new_n22260,
    new_n22261, new_n22262, new_n22263, new_n22264, new_n22265, new_n22266,
    new_n22267, new_n22268, new_n22269, new_n22270_1, new_n22271,
    new_n22272, new_n22273, new_n22274_1, new_n22275, new_n22276,
    new_n22277, new_n22278, new_n22279, new_n22280, new_n22281, new_n22282,
    new_n22283_1, new_n22284, new_n22285, new_n22286, new_n22287,
    new_n22288, new_n22289, new_n22290_1, new_n22291, new_n22292,
    new_n22293, new_n22294, new_n22295, new_n22296, new_n22297, new_n22298,
    new_n22299, new_n22300, new_n22301, new_n22302, new_n22303, new_n22304,
    new_n22305, new_n22306, new_n22307, new_n22308, new_n22309_1,
    new_n22310, new_n22311_1, new_n22312, new_n22313, new_n22314,
    new_n22315, new_n22316, new_n22317_1, new_n22318, new_n22319,
    new_n22320, new_n22321, new_n22322, new_n22323, new_n22324, new_n22325,
    new_n22326, new_n22327, new_n22328, new_n22329, new_n22330, new_n22331,
    new_n22332_1, new_n22333, new_n22337, new_n22340, new_n22341_1,
    new_n22342, new_n22343, new_n22344, new_n22345, new_n22346, new_n22347,
    new_n22348, new_n22349, new_n22350, new_n22351, new_n22352,
    new_n22353_1, new_n22354, new_n22355, new_n22360, new_n22361,
    new_n22362, new_n22363, new_n22364, new_n22365, new_n22366, new_n22367,
    new_n22368, new_n22369, new_n22370, new_n22371, new_n22372, new_n22373,
    new_n22374, new_n22375, new_n22376, new_n22377, new_n22378,
    new_n22379_1, new_n22380, new_n22381, new_n22382, new_n22383,
    new_n22384, new_n22386, new_n22387, new_n22388, new_n22389, new_n22390,
    new_n22391, new_n22395, new_n22396, new_n22397, new_n22398, new_n22404,
    new_n22409, new_n22410, new_n22411, new_n22412, new_n22413, new_n22414,
    new_n22415, new_n22416, new_n22417, new_n22418, new_n22419, new_n22420,
    new_n22421, new_n22422, new_n22423, new_n22424, new_n22425, new_n22426,
    new_n22427, new_n22428, new_n22429, new_n22430, new_n22431, new_n22452,
    new_n22453, new_n22454, new_n22455, new_n22456, new_n22457, new_n22458,
    new_n22459, new_n22460, new_n22461, new_n22462, new_n22463, new_n22464,
    new_n22465, new_n22466, new_n22467_1, new_n22468, new_n22469,
    new_n22470_1, new_n22471, new_n22472, new_n22473, new_n22474,
    new_n22475, new_n22476, new_n22477, new_n22478, new_n22479, new_n22480,
    new_n22481, new_n22482, new_n22483, new_n22484_1, new_n22485,
    new_n22486, new_n22487, new_n22495, new_n22496, new_n22497, new_n22498,
    new_n22499, new_n22500, new_n22501, new_n22502, new_n22503, new_n22504,
    new_n22505, new_n22506, new_n22507, new_n22508, new_n22512, new_n22513,
    new_n22516, new_n22517, new_n22518, new_n22519, new_n22520, new_n22521,
    new_n22522, new_n22523, new_n22526, new_n22527, new_n22528, new_n22529,
    new_n22530, new_n22531, new_n22532, new_n22533_1, new_n22534,
    new_n22535, new_n22536, new_n22537, new_n22538, new_n22539, new_n22540,
    new_n22541, new_n22542, new_n22543, new_n22544, new_n22545, new_n22546,
    new_n22547, new_n22550, new_n22551, new_n22552, new_n22553,
    new_n22554_1, new_n22555, new_n22556, new_n22557, new_n22558,
    new_n22559, new_n22560, new_n22561, new_n22562, new_n22563, new_n22564,
    new_n22565, new_n22566, new_n22567, new_n22568, new_n22569, new_n22570,
    new_n22571, new_n22572, new_n22573, new_n22574, new_n22575, new_n22576,
    new_n22577, new_n22578, new_n22579, new_n22580, new_n22581, new_n22582,
    new_n22583, new_n22584_1, new_n22585, new_n22586, new_n22587,
    new_n22608, new_n22612, new_n22613, new_n22614, new_n22615, new_n22616,
    new_n22617, new_n22618, new_n22619_1, new_n22620_1, new_n22621,
    new_n22622, new_n22623_1, new_n22624, new_n22625, new_n22628,
    new_n22629, new_n22630, new_n22631_1, new_n22632, new_n22633,
    new_n22634, new_n22635, new_n22636, new_n22637, new_n22638, new_n22639,
    new_n22640, new_n22641, new_n22642, new_n22643, new_n22644, new_n22645,
    new_n22646, new_n22647, new_n22651, new_n22652, new_n22653, new_n22654,
    new_n22655, new_n22656, new_n22657, new_n22661, new_n22664, new_n22667,
    new_n22668, new_n22669, new_n22670, new_n22671, new_n22672, new_n22673,
    new_n22675, new_n22676, new_n22677, new_n22678, new_n22679, new_n22680,
    new_n22681, new_n22682, new_n22683, new_n22684, new_n22685, new_n22686,
    new_n22687, new_n22688, new_n22689, new_n22690, new_n22691, new_n22692,
    new_n22693, new_n22714_1, new_n22717, new_n22718, new_n22719,
    new_n22720, new_n22721, new_n22722, new_n22723, new_n22724, new_n22725,
    new_n22726, new_n22727, new_n22728, new_n22729, new_n22730, new_n22731,
    new_n22732, new_n22733, new_n22734, new_n22735, new_n22736, new_n22737,
    new_n22742, new_n22743, new_n22744, new_n22745, new_n22757, new_n22760,
    new_n22775, new_n22776, new_n22777, new_n22778, new_n22779_1,
    new_n22780, new_n22794, new_n22795, new_n22796, new_n22797, new_n22798,
    new_n22799, new_n22800, new_n22804, new_n22805, new_n22806, new_n22807,
    new_n22808, new_n22809, new_n22810, new_n22815, new_n22816, new_n22817,
    new_n22818, new_n22819_1, new_n22820, new_n22821, new_n22822,
    new_n22823, new_n22826, new_n22827, new_n22842, new_n22843_1,
    new_n22844, new_n22847, new_n22848, new_n22849, new_n22850,
    new_n22858_1, new_n22859, new_n22868, new_n22874, new_n22879_1,
    new_n22880, new_n22881, new_n22882, new_n22883, new_n22884, new_n22885,
    new_n22886, new_n22887, new_n22888, new_n22896, new_n22898, new_n22899,
    new_n22900, new_n22901, new_n22902, new_n22903_1, new_n22904,
    new_n22905, new_n22906, new_n22907_1, new_n22909, new_n22910_1,
    new_n22911, new_n22912, new_n22923, new_n22924, new_n22926, new_n22927,
    new_n22928, new_n22929, new_n22930, new_n22931, new_n22932, new_n22933,
    new_n22934, new_n22935, new_n22936, new_n22937, new_n22938,
    new_n22939_1, new_n22957, new_n22958, new_n22959, new_n22960,
    new_n22961, new_n22962, new_n22963, new_n22964, new_n22965, new_n22966,
    new_n22967, new_n22968, new_n22969, new_n22972, new_n22973, new_n22974,
    new_n22975, new_n22979, new_n22981, new_n22982, new_n22983, new_n22984,
    new_n22985, new_n22986, new_n22987, new_n22988, new_n22991, new_n22992,
    new_n22993, new_n22994, new_n22995, new_n22998_1, new_n22999,
    new_n23000, new_n23001, new_n23002, new_n23004, new_n23005,
    new_n23006_1, new_n23007_1, new_n23008, new_n23009_1, new_n23010,
    new_n23011, new_n23012, new_n23013, new_n23014_1, new_n23015,
    new_n23016, new_n23017, new_n23018, new_n23019, new_n23020, new_n23021,
    new_n23022, new_n23023, new_n23024, new_n23025, new_n23026, new_n23030,
    new_n23031, new_n23032, new_n23033, new_n23034, new_n23035_1,
    new_n23049, new_n23050, new_n23061, new_n23068_1, new_n23069,
    new_n23070, new_n23071, new_n23072, new_n23073, new_n23081, new_n23100,
    new_n23122, new_n23123, new_n23137, new_n23138, new_n23139, new_n23140,
    new_n23141, new_n23142, new_n23143, new_n23144, new_n23151, new_n23159,
    new_n23160_1, new_n23161, new_n23162, new_n23163, new_n23164,
    new_n23165, new_n23166_1, new_n23167, new_n23168, new_n23169,
    new_n23170, new_n23176, new_n23177, new_n23178, new_n23179, new_n23180,
    new_n23181, new_n23182, new_n23183, new_n23184, new_n23187, new_n23188,
    new_n23189, new_n23190, new_n23196, new_n23197, new_n23198, new_n23199,
    new_n23201, new_n23202, new_n23203, new_n23204, new_n23205, new_n23206,
    new_n23207, new_n23208, new_n23209, new_n23210, new_n23211, new_n23212,
    new_n23213, new_n23214, new_n23215, new_n23227, new_n23255, new_n23256,
    new_n23257, new_n23258, new_n23269, new_n23275, new_n23276, new_n23277,
    new_n23278, new_n23279, new_n23294, new_n23301, new_n23302, new_n23303,
    new_n23304_1, new_n23305_1, new_n23306, new_n23307, new_n23308,
    new_n23323, new_n23324, new_n23325, new_n23326, new_n23327, new_n23328,
    new_n23329, new_n23330, new_n23335, new_n23341_1, new_n23342_1,
    new_n23343, new_n23344, new_n23345, new_n23346, new_n23347, new_n23348,
    new_n23349, new_n23350, new_n23363, new_n23364, new_n23365,
    new_n23369_1, new_n23374, new_n23375, new_n23376, new_n23377,
    new_n23384, new_n23385, new_n23386, new_n23387, new_n23388, new_n23389,
    new_n23390, new_n23396, new_n23397, new_n23405, new_n23406, new_n23407,
    new_n23408, new_n23409, new_n23412, new_n23415, new_n23416, new_n23417,
    new_n23418, new_n23431, new_n23432, new_n23433_1, new_n23434_1,
    new_n23436, new_n23447, new_n23448, new_n23449, new_n23450_1,
    new_n23453, new_n23461, new_n23462, new_n23463_1, new_n23464,
    new_n23465, new_n23466, new_n23467, new_n23468, new_n23469,
    new_n23471_1, new_n23476, new_n23477, new_n23478, new_n23479,
    new_n23481, new_n23482, new_n23483, new_n23484, new_n23489, new_n23490,
    new_n23491, new_n23492, new_n23493_1, new_n23494, new_n23495,
    new_n23496, new_n23497, new_n23498, new_n23499, new_n23500, new_n23501,
    new_n23502, new_n23503, new_n23504, new_n23505, new_n23506, new_n23507,
    new_n23508, new_n23509, new_n23510, new_n23515, new_n23516, new_n23517,
    new_n23518, new_n23522, new_n23532, new_n23533, new_n23534, new_n23535,
    new_n23536, new_n23555, new_n23556, new_n23557, new_n23558, new_n23559,
    new_n23560, new_n23562, new_n23563, new_n23564, new_n23565, new_n23566,
    new_n23567, new_n23578, new_n23590, new_n23591, new_n23595, new_n23596,
    new_n23597, new_n23598, new_n23600, new_n23601, new_n23603, new_n23613,
    new_n23614, new_n23615, new_n23616, new_n23617, new_n23626,
    new_n23637_1, new_n23646, new_n23655, new_n23656, new_n23666,
    new_n23667, new_n23668, new_n23669_1, new_n23675, new_n23676,
    new_n23677, new_n23678, new_n23681, new_n23682, new_n23683,
    new_n23684_1, new_n23705, new_n23725, new_n23735, new_n23736,
    new_n23737, new_n23751, new_n23752, new_n23767, new_n23783, new_n23788,
    new_n23791, new_n23792, new_n23798, new_n23799, new_n23800, new_n23804,
    new_n23805, new_n23806, new_n23807, new_n23809, new_n23822, new_n23825,
    new_n23826, new_n23827, new_n23828, new_n23831_1, new_n23834,
    new_n23835, new_n23836, new_n23837, new_n23851, new_n23852, new_n23855,
    new_n23867, new_n23869, new_n23870, new_n23871, new_n23872, new_n23875,
    new_n23876, new_n23886, new_n23888_1, new_n23893, new_n23894,
    new_n23895_1, new_n23896, new_n23902, new_n23903_1, new_n23913_1,
    new_n23927, new_n23936, new_n23937, new_n23940;
xnor g00000 ( new_n2349 , n9942 , n10739 );
not  g00001 ( new_n2350 , n21753 );
nor  g00002 ( new_n2351 , new_n2350 , n25643 );
xnor g00003 ( new_n2352 , n21753 , n25643 );
not  g00004 ( new_n2353 , n21832 );
nor  g00005 ( new_n2354 , n9557 , new_n2353 );
xnor g00006 ( new_n2355_1 , n9557 , n21832 );
not  g00007 ( new_n2356 , n26913 );
nor  g00008 ( new_n2357 , n3136 , new_n2356 );
xnor g00009 ( new_n2358 , n3136 , n26913 );
not  g00010 ( new_n2359 , n6385 );
nor  g00011 ( new_n2360 , new_n2359 , n16223 );
not  g00012 ( new_n2361_1 , n16223 );
nor  g00013 ( new_n2362 , n6385 , new_n2361_1 );
not  g00014 ( new_n2363_1 , n20138 );
nor  g00015 ( new_n2364 , n19494 , new_n2363_1 );
not  g00016 ( new_n2365 , n19494 );
nor  g00017 ( new_n2366 , new_n2365 , n20138 );
not  g00018 ( new_n2367 , n9251 );
nor  g00019 ( new_n2368 , n2387 , new_n2367 );
not  g00020 ( new_n2369 , new_n2368 );
nor  g00021 ( new_n2370 , new_n2366 , new_n2369 );
nor  g00022 ( new_n2371 , new_n2364 , new_n2370 );
nor  g00023 ( new_n2372 , new_n2362 , new_n2371 );
nor  g00024 ( new_n2373 , new_n2360 , new_n2372 );
and  g00025 ( new_n2374_1 , new_n2358 , new_n2373 );
or   g00026 ( new_n2375 , new_n2357 , new_n2374_1 );
and  g00027 ( new_n2376 , new_n2355_1 , new_n2375 );
or   g00028 ( new_n2377 , new_n2354 , new_n2376 );
and  g00029 ( new_n2378 , new_n2352 , new_n2377 );
or   g00030 ( new_n2379 , new_n2351 , new_n2378 );
xor  g00031 ( new_n2380 , new_n2349 , new_n2379 );
not  g00032 ( new_n2381 , n5704 );
xnor g00033 ( new_n2382 , new_n2381 , n13781 );
not  g00034 ( new_n2383 , n13781 );
nor  g00035 ( new_n2384 , new_n2381 , new_n2383 );
xnor g00036 ( new_n2385 , n11486 , n18409 );
xnor g00037 ( new_n2386 , new_n2384 , new_n2385 );
nor  g00038 ( new_n2387_1 , new_n2382 , new_n2386 );
not  g00039 ( new_n2388_1 , new_n2387_1 );
not  g00040 ( new_n2389 , n13708 );
xnor g00041 ( new_n2390 , new_n2389 , n16722 );
nor  g00042 ( new_n2391 , n11486 , n18409 );
nor  g00043 ( new_n2392 , new_n2384 , new_n2385 );
nor  g00044 ( new_n2393 , new_n2391 , new_n2392 );
xnor g00045 ( new_n2394 , new_n2390 , new_n2393 );
not  g00046 ( new_n2395 , new_n2394 );
nor  g00047 ( new_n2396 , new_n2388_1 , new_n2395 );
not  g00048 ( new_n2397 , new_n2396 );
not  g00049 ( new_n2398 , n3480 );
xnor g00050 ( new_n2399 , new_n2398 , n19911 );
nor  g00051 ( new_n2400 , n13708 , n16722 );
or   g00052 ( new_n2401 , new_n2391 , new_n2392 );
and  g00053 ( new_n2402 , new_n2390 , new_n2401 );
nor  g00054 ( new_n2403 , new_n2400 , new_n2402 );
xnor g00055 ( new_n2404 , new_n2399 , new_n2403 );
not  g00056 ( new_n2405 , new_n2404 );
nor  g00057 ( new_n2406 , new_n2397 , new_n2405 );
not  g00058 ( new_n2407 , new_n2406 );
not  g00059 ( new_n2408 , n2731 );
xnor g00060 ( new_n2409_1 , new_n2408 , n3018 );
nor  g00061 ( new_n2410 , n3480 , n19911 );
or   g00062 ( new_n2411 , new_n2400 , new_n2402 );
and  g00063 ( new_n2412 , new_n2399 , new_n2411 );
nor  g00064 ( new_n2413 , new_n2410 , new_n2412 );
xnor g00065 ( new_n2414 , new_n2409_1 , new_n2413 );
not  g00066 ( new_n2415 , new_n2414 );
nor  g00067 ( new_n2416_1 , new_n2407 , new_n2415 );
not  g00068 ( new_n2417 , new_n2416_1 );
xnor g00069 ( new_n2418 , n18907 , n26660 );
nor  g00070 ( new_n2419 , n2731 , n3018 );
or   g00071 ( new_n2420_1 , new_n2410 , new_n2412 );
and  g00072 ( new_n2421_1 , new_n2409_1 , new_n2420_1 );
nor  g00073 ( new_n2422 , new_n2419 , new_n2421_1 );
xnor g00074 ( new_n2423 , new_n2418 , new_n2422 );
nor  g00075 ( new_n2424 , new_n2417 , new_n2423 );
not  g00076 ( new_n2425 , n13783 );
xnor g00077 ( new_n2426 , new_n2425 , n22332 );
nor  g00078 ( new_n2427 , n18907 , n26660 );
nor  g00079 ( new_n2428 , new_n2418 , new_n2422 );
nor  g00080 ( new_n2429 , new_n2427 , new_n2428 );
xnor g00081 ( new_n2430 , new_n2426 , new_n2429 );
not  g00082 ( new_n2431 , new_n2430 );
xnor g00083 ( new_n2432 , new_n2424 , new_n2431 );
xnor g00084 ( new_n2433 , n7751 , n13490 );
nor  g00085 ( new_n2434 , n22660 , n26823 );
xnor g00086 ( new_n2435 , n22660 , n26823 );
nor  g00087 ( new_n2436 , n1777 , n4812 );
xnor g00088 ( new_n2437 , n1777 , n4812 );
nor  g00089 ( new_n2438 , n8745 , n24278 );
xnor g00090 ( new_n2439 , n8745 , n24278 );
nor  g00091 ( new_n2440_1 , n15636 , n24618 );
not  g00092 ( new_n2441 , n15636 );
xnor g00093 ( new_n2442 , new_n2441 , n24618 );
not  g00094 ( new_n2443 , n3952 );
not  g00095 ( new_n2444_1 , n20077 );
nor  g00096 ( new_n2445 , new_n2443 , new_n2444_1 );
or   g00097 ( new_n2446 , n3952 , n20077 );
not  g00098 ( new_n2447 , n6794 );
not  g00099 ( new_n2448 , n12315 );
nor  g00100 ( new_n2449 , new_n2447 , new_n2448 );
and  g00101 ( new_n2450 , new_n2446 , new_n2449 );
nor  g00102 ( new_n2451 , new_n2445 , new_n2450 );
and  g00103 ( new_n2452 , new_n2442 , new_n2451 );
nor  g00104 ( new_n2453 , new_n2440_1 , new_n2452 );
nor  g00105 ( new_n2454 , new_n2439 , new_n2453 );
nor  g00106 ( new_n2455 , new_n2438 , new_n2454 );
nor  g00107 ( new_n2456 , new_n2437 , new_n2455 );
nor  g00108 ( new_n2457 , new_n2436 , new_n2456 );
nor  g00109 ( new_n2458 , new_n2435 , new_n2457 );
nor  g00110 ( new_n2459 , new_n2434 , new_n2458 );
xnor g00111 ( new_n2460 , new_n2433 , new_n2459 );
xnor g00112 ( new_n2461 , new_n2432 , new_n2460 );
xnor g00113 ( new_n2462 , new_n2416_1 , new_n2423 );
xnor g00114 ( new_n2463 , new_n2435 , new_n2457 );
nor  g00115 ( new_n2464 , new_n2462 , new_n2463 );
xnor g00116 ( new_n2465 , new_n2406 , new_n2415 );
xnor g00117 ( new_n2466 , new_n2437 , new_n2455 );
nor  g00118 ( new_n2467 , new_n2465 , new_n2466 );
xnor g00119 ( new_n2468 , new_n2465 , new_n2466 );
xnor g00120 ( new_n2469 , new_n2396 , new_n2405 );
xnor g00121 ( new_n2470 , new_n2439 , new_n2453 );
nor  g00122 ( new_n2471 , new_n2469 , new_n2470 );
xnor g00123 ( new_n2472 , new_n2387_1 , new_n2395 );
xnor g00124 ( new_n2473 , new_n2442 , new_n2451 );
nor  g00125 ( new_n2474 , new_n2472 , new_n2473 );
not  g00126 ( new_n2475 , new_n2473 );
xnor g00127 ( new_n2476 , new_n2472 , new_n2475 );
not  g00128 ( new_n2477 , new_n2382 );
xnor g00129 ( new_n2478 , n6794 , n12315 );
nor  g00130 ( new_n2479_1 , new_n2477 , new_n2478 );
xnor g00131 ( new_n2480 , n3952 , n20077 );
xnor g00132 ( new_n2481 , new_n2449 , new_n2480 );
nor  g00133 ( new_n2482 , new_n2479_1 , new_n2481 );
or   g00134 ( new_n2483 , n5704 , n13781 );
and  g00135 ( new_n2484 , new_n2483 , new_n2392 );
or   g00136 ( new_n2485 , new_n2387_1 , new_n2484 );
not  g00137 ( new_n2486 , new_n2479_1 );
nor  g00138 ( new_n2487 , new_n2486 , new_n2480 );
nor  g00139 ( new_n2488 , new_n2482 , new_n2487 );
and  g00140 ( new_n2489 , new_n2485 , new_n2488 );
or   g00141 ( new_n2490 , new_n2482 , new_n2489 );
and  g00142 ( new_n2491 , new_n2476 , new_n2490 );
nor  g00143 ( new_n2492 , new_n2474 , new_n2491 );
xnor g00144 ( new_n2493 , new_n2469 , new_n2470 );
nor  g00145 ( new_n2494 , new_n2492 , new_n2493 );
nor  g00146 ( new_n2495 , new_n2471 , new_n2494 );
nor  g00147 ( new_n2496 , new_n2468 , new_n2495 );
nor  g00148 ( new_n2497 , new_n2467 , new_n2496 );
xnor g00149 ( new_n2498 , new_n2462 , new_n2463 );
nor  g00150 ( new_n2499 , new_n2497 , new_n2498 );
nor  g00151 ( new_n2500 , new_n2464 , new_n2499 );
xnor g00152 ( new_n2501 , new_n2461 , new_n2500 );
xor  g00153 ( new_n2502 , new_n2380 , new_n2501 );
xor  g00154 ( new_n2503 , new_n2352 , new_n2377 );
xnor g00155 ( new_n2504 , new_n2497 , new_n2498 );
nor  g00156 ( new_n2505 , new_n2503 , new_n2504 );
xnor g00157 ( new_n2506 , new_n2503 , new_n2504 );
xor  g00158 ( new_n2507 , new_n2355_1 , new_n2375 );
xnor g00159 ( new_n2508 , new_n2468 , new_n2495 );
nor  g00160 ( new_n2509 , new_n2507 , new_n2508 );
xnor g00161 ( new_n2510 , new_n2507 , new_n2508 );
xnor g00162 ( new_n2511 , new_n2358 , new_n2373 );
xnor g00163 ( new_n2512 , new_n2492 , new_n2493 );
not  g00164 ( new_n2513_1 , new_n2512 );
and  g00165 ( new_n2514 , new_n2511 , new_n2513_1 );
xnor g00166 ( new_n2515_1 , new_n2511 , new_n2513_1 );
xor  g00167 ( new_n2516 , new_n2476 , new_n2490 );
xnor g00168 ( new_n2517 , n6385 , n16223 );
xnor g00169 ( new_n2518 , new_n2371 , new_n2517 );
and  g00170 ( new_n2519 , new_n2516 , new_n2518 );
xnor g00171 ( new_n2520 , new_n2516 , new_n2518 );
xnor g00172 ( new_n2521 , n2387 , n9251 );
xnor g00173 ( new_n2522 , new_n2382 , new_n2478 );
not  g00174 ( new_n2523 , new_n2522 );
or   g00175 ( new_n2524 , new_n2521 , new_n2523 );
xnor g00176 ( new_n2525 , n19494 , n20138 );
xnor g00177 ( new_n2526 , new_n2369 , new_n2525 );
and  g00178 ( new_n2527 , new_n2524 , new_n2526 );
xnor g00179 ( new_n2528 , new_n2485 , new_n2488 );
not  g00180 ( new_n2529 , new_n2528 );
xor  g00181 ( new_n2530 , new_n2524 , new_n2526 );
and  g00182 ( new_n2531 , new_n2529 , new_n2530 );
nor  g00183 ( new_n2532 , new_n2527 , new_n2531 );
nor  g00184 ( new_n2533_1 , new_n2520 , new_n2532 );
nor  g00185 ( new_n2534 , new_n2519 , new_n2533_1 );
nor  g00186 ( new_n2535_1 , new_n2515_1 , new_n2534 );
nor  g00187 ( new_n2536 , new_n2514 , new_n2535_1 );
nor  g00188 ( new_n2537_1 , new_n2510 , new_n2536 );
nor  g00189 ( new_n2538 , new_n2509 , new_n2537_1 );
nor  g00190 ( new_n2539 , new_n2506 , new_n2538 );
nor  g00191 ( new_n2540 , new_n2505 , new_n2539 );
xor  g00192 ( n7 , new_n2502 , new_n2540 );
not  g00193 ( new_n2542 , n4588 );
xnor g00194 ( new_n2543 , n1681 , n3618 );
xnor g00195 ( new_n2544 , new_n2542 , new_n2543 );
xnor g00196 ( new_n2545 , n583 , n22843 );
xnor g00197 ( new_n2546 , n22201 , new_n2545 );
xnor g00198 ( n50 , new_n2544 , new_n2546 );
not  g00199 ( new_n2548 , n21687 );
xnor g00200 ( new_n2549 , n6773 , n19922 );
xnor g00201 ( new_n2550 , new_n2548 , new_n2549 );
xnor g00202 ( new_n2551 , n14090 , n21398 );
xnor g00203 ( new_n2552 , n25926 , new_n2551 );
xnor g00204 ( n55 , new_n2550 , new_n2552 );
not  g00205 ( new_n2554 , n9396 );
xnor g00206 ( new_n2555_1 , new_n2554 , n20040 );
not  g00207 ( new_n2556 , new_n2555_1 );
nor  g00208 ( new_n2557 , n1999 , n19531 );
not  g00209 ( new_n2558 , n19531 );
xnor g00210 ( new_n2559 , n1999 , new_n2558 );
not  g00211 ( new_n2560_1 , new_n2559 );
nor  g00212 ( new_n2561_1 , n18345 , n25168 );
not  g00213 ( new_n2562 , n18345 );
xnor g00214 ( new_n2563 , new_n2562 , n25168 );
not  g00215 ( new_n2564 , new_n2563 );
nor  g00216 ( new_n2565 , n9318 , n13190 );
not  g00217 ( new_n2566 , n13190 );
xnor g00218 ( new_n2567 , n9318 , new_n2566 );
not  g00219 ( new_n2568 , new_n2567 );
nor  g00220 ( new_n2569 , n3460 , n19477 );
xnor g00221 ( new_n2570_1 , n3460 , n19477 );
nor  g00222 ( new_n2571 , n5226 , n11223 );
xnor g00223 ( new_n2572 , n5226 , n11223 );
nor  g00224 ( new_n2573_1 , n5115 , n17664 );
not  g00225 ( new_n2574 , n17664 );
xnor g00226 ( new_n2575 , n5115 , new_n2574 );
not  g00227 ( new_n2576 , new_n2575 );
nor  g00228 ( new_n2577 , n23369 , n26572 );
not  g00229 ( new_n2578_1 , n23369 );
xnor g00230 ( new_n2579 , new_n2578_1 , n26572 );
not  g00231 ( new_n2580 , new_n2579 );
nor  g00232 ( new_n2581 , n1136 , n11667 );
not  g00233 ( new_n2582_1 , n19234 );
not  g00234 ( new_n2583 , n21398 );
nor  g00235 ( new_n2584 , new_n2582_1 , new_n2583 );
xnor g00236 ( new_n2585 , n1136 , n11667 );
nor  g00237 ( new_n2586 , new_n2584 , new_n2585 );
nor  g00238 ( new_n2587 , new_n2581 , new_n2586 );
nor  g00239 ( new_n2588 , new_n2580 , new_n2587 );
nor  g00240 ( new_n2589 , new_n2577 , new_n2588 );
nor  g00241 ( new_n2590 , new_n2576 , new_n2589 );
nor  g00242 ( new_n2591 , new_n2573_1 , new_n2590 );
nor  g00243 ( new_n2592 , new_n2572 , new_n2591 );
nor  g00244 ( new_n2593 , new_n2571 , new_n2592 );
nor  g00245 ( new_n2594 , new_n2570_1 , new_n2593 );
nor  g00246 ( new_n2595 , new_n2569 , new_n2594 );
nor  g00247 ( new_n2596 , new_n2568 , new_n2595 );
nor  g00248 ( new_n2597 , new_n2565 , new_n2596 );
nor  g00249 ( new_n2598 , new_n2564 , new_n2597 );
nor  g00250 ( new_n2599 , new_n2561_1 , new_n2598 );
nor  g00251 ( new_n2600 , new_n2560_1 , new_n2599 );
nor  g00252 ( new_n2601 , new_n2557 , new_n2600 );
xnor g00253 ( new_n2602_1 , new_n2556 , new_n2601 );
not  g00254 ( new_n2603 , new_n2602_1 );
xnor g00255 ( new_n2604 , n25365 , new_n2603 );
xnor g00256 ( new_n2605 , new_n2560_1 , new_n2599 );
and  g00257 ( new_n2606 , n14704 , new_n2605 );
not  g00258 ( new_n2607 , new_n2605 );
xnor g00259 ( new_n2608 , n14704 , new_n2607 );
xnor g00260 ( new_n2609 , new_n2564 , new_n2597 );
and  g00261 ( new_n2610 , n19270 , new_n2609 );
not  g00262 ( new_n2611 , new_n2609 );
xnor g00263 ( new_n2612 , n19270 , new_n2611 );
xnor g00264 ( new_n2613 , new_n2568 , new_n2595 );
and  g00265 ( new_n2614 , n8687 , new_n2613 );
xnor g00266 ( new_n2615 , new_n2570_1 , new_n2593 );
nor  g00267 ( new_n2616 , n24768 , new_n2615 );
xnor g00268 ( new_n2617 , n24768 , new_n2615 );
xnor g00269 ( new_n2618 , new_n2572 , new_n2591 );
nor  g00270 ( new_n2619_1 , n26483 , new_n2618 );
xnor g00271 ( new_n2620 , n26483 , new_n2618 );
xnor g00272 ( new_n2621 , new_n2576 , new_n2589 );
and  g00273 ( new_n2622 , n15979 , new_n2621 );
not  g00274 ( new_n2623 , new_n2621 );
xnor g00275 ( new_n2624 , n15979 , new_n2623 );
xnor g00276 ( new_n2625 , new_n2580 , new_n2587 );
and  g00277 ( new_n2626 , n8638 , new_n2625 );
xnor g00278 ( new_n2627 , new_n2584 , new_n2585 );
nor  g00279 ( new_n2628 , n16247 , new_n2627 );
not  g00280 ( new_n2629 , n23541 );
xnor g00281 ( new_n2630 , n19234 , n21398 );
or   g00282 ( new_n2631 , new_n2629 , new_n2630 );
not  g00283 ( new_n2632 , n16247 );
xnor g00284 ( new_n2633 , new_n2632 , new_n2627 );
and  g00285 ( new_n2634 , new_n2631 , new_n2633 );
nor  g00286 ( new_n2635 , new_n2628 , new_n2634 );
not  g00287 ( new_n2636 , new_n2625 );
xnor g00288 ( new_n2637 , n8638 , new_n2636 );
and  g00289 ( new_n2638 , new_n2635 , new_n2637 );
or   g00290 ( new_n2639 , new_n2626 , new_n2638 );
and  g00291 ( new_n2640 , new_n2624 , new_n2639 );
nor  g00292 ( new_n2641 , new_n2622 , new_n2640 );
not  g00293 ( new_n2642 , new_n2641 );
nor  g00294 ( new_n2643 , new_n2620 , new_n2642 );
nor  g00295 ( new_n2644 , new_n2619_1 , new_n2643 );
nor  g00296 ( new_n2645 , new_n2617 , new_n2644 );
nor  g00297 ( new_n2646_1 , new_n2616 , new_n2645 );
not  g00298 ( new_n2647 , new_n2613 );
xnor g00299 ( new_n2648 , n8687 , new_n2647 );
and  g00300 ( new_n2649 , new_n2646_1 , new_n2648 );
or   g00301 ( new_n2650 , new_n2614 , new_n2649 );
and  g00302 ( new_n2651 , new_n2612 , new_n2650 );
or   g00303 ( new_n2652 , new_n2610 , new_n2651 );
and  g00304 ( new_n2653 , new_n2608 , new_n2652 );
nor  g00305 ( new_n2654 , new_n2606 , new_n2653 );
xnor g00306 ( new_n2655 , new_n2604 , new_n2654 );
not  g00307 ( new_n2656 , new_n2655 );
nor  g00308 ( new_n2657 , n11503 , n18151 );
not  g00309 ( new_n2658 , new_n2657 );
nor  g00310 ( new_n2659_1 , n16971 , new_n2658 );
not  g00311 ( new_n2660 , new_n2659_1 );
nor  g00312 ( new_n2661_1 , n10411 , new_n2660 );
not  g00313 ( new_n2662 , new_n2661_1 );
nor  g00314 ( new_n2663 , n23430 , new_n2662 );
not  g00315 ( new_n2664 , new_n2663 );
nor  g00316 ( new_n2665 , n5579 , new_n2664 );
not  g00317 ( new_n2666 , new_n2665 );
nor  g00318 ( new_n2667 , n25523 , new_n2666 );
not  g00319 ( new_n2668 , new_n2667 );
nor  g00320 ( new_n2669 , n8439 , new_n2668 );
not  g00321 ( new_n2670 , new_n2669 );
nor  g00322 ( new_n2671 , n22793 , new_n2670 );
not  g00323 ( new_n2672 , new_n2671 );
xnor g00324 ( new_n2673 , n13951 , new_n2672 );
not  g00325 ( new_n2674 , n2944 );
xnor g00326 ( new_n2675 , new_n2674 , n22270 );
nor  g00327 ( new_n2676 , n767 , n8806 );
not  g00328 ( new_n2677 , n767 );
xnor g00329 ( new_n2678 , new_n2677 , n8806 );
nor  g00330 ( new_n2679 , n2479 , n7330 );
not  g00331 ( new_n2680_1 , n2479 );
xnor g00332 ( new_n2681 , new_n2680_1 , n7330 );
nor  g00333 ( new_n2682 , n9372 , n22492 );
not  g00334 ( new_n2683 , n22492 );
xnor g00335 ( new_n2684 , n9372 , new_n2683 );
nor  g00336 ( new_n2685 , n6596 , n12821 );
not  g00337 ( new_n2686 , n6596 );
xnor g00338 ( new_n2687 , new_n2686 , n12821 );
nor  g00339 ( new_n2688 , n3468 , n15289 );
not  g00340 ( new_n2689 , n3468 );
xnor g00341 ( new_n2690 , new_n2689 , n15289 );
nor  g00342 ( new_n2691 , n6556 , n18558 );
not  g00343 ( new_n2692 , n6556 );
xnor g00344 ( new_n2693_1 , new_n2692 , n18558 );
nor  g00345 ( new_n2694 , n7149 , n22871 );
not  g00346 ( new_n2695 , n7149 );
xnor g00347 ( new_n2696 , new_n2695 , n22871 );
nor  g00348 ( new_n2697 , n14148 , n14275 );
not  g00349 ( new_n2698 , n1152 );
not  g00350 ( new_n2699 , n25023 );
or   g00351 ( new_n2700 , new_n2698 , new_n2699 );
not  g00352 ( new_n2701 , n14148 );
xnor g00353 ( new_n2702 , new_n2701 , n14275 );
and  g00354 ( new_n2703_1 , new_n2700 , new_n2702 );
or   g00355 ( new_n2704 , new_n2697 , new_n2703_1 );
and  g00356 ( new_n2705 , new_n2696 , new_n2704 );
or   g00357 ( new_n2706_1 , new_n2694 , new_n2705 );
and  g00358 ( new_n2707 , new_n2693_1 , new_n2706_1 );
or   g00359 ( new_n2708 , new_n2691 , new_n2707 );
and  g00360 ( new_n2709 , new_n2690 , new_n2708 );
or   g00361 ( new_n2710 , new_n2688 , new_n2709 );
and  g00362 ( new_n2711_1 , new_n2687 , new_n2710 );
or   g00363 ( new_n2712 , new_n2685 , new_n2711_1 );
and  g00364 ( new_n2713 , new_n2684 , new_n2712 );
or   g00365 ( new_n2714 , new_n2682 , new_n2713 );
and  g00366 ( new_n2715 , new_n2681 , new_n2714 );
or   g00367 ( new_n2716 , new_n2679 , new_n2715 );
and  g00368 ( new_n2717 , new_n2678 , new_n2716 );
nor  g00369 ( new_n2718 , new_n2676 , new_n2717 );
xnor g00370 ( new_n2719 , new_n2675 , new_n2718 );
xnor g00371 ( new_n2720 , new_n2673 , new_n2719 );
xnor g00372 ( new_n2721 , n22793 , new_n2669 );
nor  g00373 ( new_n2722 , new_n2679 , new_n2715 );
xnor g00374 ( new_n2723 , new_n2678 , new_n2722 );
and  g00375 ( new_n2724 , new_n2721 , new_n2723 );
not  g00376 ( new_n2725 , new_n2723 );
xnor g00377 ( new_n2726 , new_n2721 , new_n2725 );
xnor g00378 ( new_n2727 , n8439 , new_n2667 );
nor  g00379 ( new_n2728 , new_n2682 , new_n2713 );
xnor g00380 ( new_n2729 , new_n2681 , new_n2728 );
nor  g00381 ( new_n2730 , new_n2727 , new_n2729 );
xnor g00382 ( new_n2731_1 , new_n2727 , new_n2729 );
xnor g00383 ( new_n2732 , n25523 , new_n2665 );
xor  g00384 ( new_n2733 , new_n2684 , new_n2712 );
nor  g00385 ( new_n2734 , new_n2732 , new_n2733 );
xnor g00386 ( new_n2735 , new_n2732 , new_n2733 );
xnor g00387 ( new_n2736 , n5579 , new_n2663 );
nor  g00388 ( new_n2737 , new_n2688 , new_n2709 );
xnor g00389 ( new_n2738 , new_n2687 , new_n2737 );
nor  g00390 ( new_n2739 , new_n2736 , new_n2738 );
not  g00391 ( new_n2740 , new_n2738 );
xnor g00392 ( new_n2741 , new_n2736 , new_n2740 );
xnor g00393 ( new_n2742 , n23430 , new_n2661_1 );
nor  g00394 ( new_n2743_1 , new_n2691 , new_n2707 );
xnor g00395 ( new_n2744 , new_n2690 , new_n2743_1 );
nor  g00396 ( new_n2745 , new_n2742 , new_n2744 );
xnor g00397 ( new_n2746 , n10411 , new_n2659_1 );
nor  g00398 ( new_n2747 , new_n2694 , new_n2705 );
xnor g00399 ( new_n2748 , new_n2693_1 , new_n2747 );
nor  g00400 ( new_n2749 , new_n2746 , new_n2748 );
xnor g00401 ( new_n2750 , new_n2746 , new_n2748 );
xnor g00402 ( new_n2751 , n16971 , new_n2657 );
nor  g00403 ( new_n2752 , new_n2697 , new_n2703_1 );
xnor g00404 ( new_n2753 , new_n2696 , new_n2752 );
nor  g00405 ( new_n2754 , new_n2751 , new_n2753 );
xnor g00406 ( new_n2755 , new_n2751 , new_n2753 );
not  g00407 ( new_n2756 , n11503 );
xnor g00408 ( new_n2757 , new_n2756 , n18151 );
nor  g00409 ( new_n2758 , new_n2698 , new_n2699 );
xnor g00410 ( new_n2759 , new_n2758 , new_n2702 );
nor  g00411 ( new_n2760 , new_n2757 , new_n2759 );
xnor g00412 ( new_n2761_1 , n1152 , n25023 );
nor  g00413 ( new_n2762 , n18151 , new_n2761_1 );
not  g00414 ( new_n2763 , new_n2759 );
xnor g00415 ( new_n2764 , new_n2757 , new_n2763 );
and  g00416 ( new_n2765 , new_n2762 , new_n2764 );
nor  g00417 ( new_n2766 , new_n2760 , new_n2765 );
nor  g00418 ( new_n2767 , new_n2755 , new_n2766 );
nor  g00419 ( new_n2768 , new_n2754 , new_n2767 );
nor  g00420 ( new_n2769 , new_n2750 , new_n2768 );
or   g00421 ( new_n2770 , new_n2749 , new_n2769 );
not  g00422 ( new_n2771 , new_n2744 );
xnor g00423 ( new_n2772 , new_n2742 , new_n2771 );
and  g00424 ( new_n2773 , new_n2770 , new_n2772 );
or   g00425 ( new_n2774_1 , new_n2745 , new_n2773 );
and  g00426 ( new_n2775 , new_n2741 , new_n2774_1 );
nor  g00427 ( new_n2776 , new_n2739 , new_n2775 );
nor  g00428 ( new_n2777 , new_n2735 , new_n2776 );
nor  g00429 ( new_n2778 , new_n2734 , new_n2777 );
nor  g00430 ( new_n2779_1 , new_n2731_1 , new_n2778 );
nor  g00431 ( new_n2780 , new_n2730 , new_n2779_1 );
and  g00432 ( new_n2781 , new_n2726 , new_n2780 );
or   g00433 ( new_n2782 , new_n2724 , new_n2781 );
xor  g00434 ( new_n2783_1 , new_n2720 , new_n2782 );
xnor g00435 ( new_n2784 , new_n2656 , new_n2783_1 );
nor  g00436 ( new_n2785 , new_n2610 , new_n2651 );
xnor g00437 ( new_n2786 , new_n2608 , new_n2785 );
not  g00438 ( new_n2787 , new_n2786 );
xnor g00439 ( new_n2788 , new_n2726 , new_n2780 );
nor  g00440 ( new_n2789 , new_n2787 , new_n2788 );
xnor g00441 ( new_n2790 , new_n2786 , new_n2788 );
nor  g00442 ( new_n2791 , new_n2614 , new_n2649 );
xnor g00443 ( new_n2792 , new_n2612 , new_n2791 );
xnor g00444 ( new_n2793 , new_n2731_1 , new_n2778 );
nor  g00445 ( new_n2794 , new_n2792 , new_n2793 );
xnor g00446 ( new_n2795 , new_n2792 , new_n2793 );
xnor g00447 ( new_n2796 , new_n2646_1 , new_n2648 );
not  g00448 ( new_n2797 , new_n2796 );
xnor g00449 ( new_n2798 , new_n2735 , new_n2776 );
nor  g00450 ( new_n2799 , new_n2797 , new_n2798 );
xnor g00451 ( new_n2800 , new_n2796 , new_n2798 );
xnor g00452 ( new_n2801 , new_n2617 , new_n2644 );
not  g00453 ( new_n2802 , new_n2801 );
xor  g00454 ( new_n2803 , new_n2741 , new_n2774_1 );
nor  g00455 ( new_n2804 , new_n2802 , new_n2803 );
xnor g00456 ( new_n2805 , new_n2801 , new_n2803 );
xnor g00457 ( new_n2806 , new_n2620 , new_n2641 );
xor  g00458 ( new_n2807 , new_n2770 , new_n2772 );
and  g00459 ( new_n2808 , new_n2806 , new_n2807 );
xnor g00460 ( new_n2809_1 , new_n2806 , new_n2807 );
xnor g00461 ( new_n2810 , new_n2750 , new_n2768 );
nor  g00462 ( new_n2811 , new_n2626 , new_n2638 );
xnor g00463 ( new_n2812 , new_n2624 , new_n2811 );
nor  g00464 ( new_n2813 , new_n2810 , new_n2812 );
not  g00465 ( new_n2814 , new_n2812 );
xnor g00466 ( new_n2815 , new_n2810 , new_n2814 );
xnor g00467 ( new_n2816_1 , new_n2755 , new_n2766 );
xnor g00468 ( new_n2817 , new_n2635 , new_n2637 );
not  g00469 ( new_n2818 , new_n2817 );
and  g00470 ( new_n2819 , new_n2816_1 , new_n2818 );
xnor g00471 ( new_n2820 , new_n2816_1 , new_n2817 );
xnor g00472 ( new_n2821 , new_n2762 , new_n2764 );
nor  g00473 ( new_n2822 , new_n2629 , new_n2630 );
xnor g00474 ( new_n2823 , new_n2822 , new_n2633 );
not  g00475 ( new_n2824 , new_n2823 );
nor  g00476 ( new_n2825 , new_n2821 , new_n2824 );
xnor g00477 ( new_n2826_1 , n23541 , new_n2630 );
not  g00478 ( new_n2827 , new_n2826_1 );
not  g00479 ( new_n2828 , n18151 );
xnor g00480 ( new_n2829 , new_n2828 , new_n2761_1 );
nor  g00481 ( new_n2830 , new_n2827 , new_n2829 );
xnor g00482 ( new_n2831 , new_n2821 , new_n2824 );
nor  g00483 ( new_n2832 , new_n2830 , new_n2831 );
nor  g00484 ( new_n2833 , new_n2825 , new_n2832 );
and  g00485 ( new_n2834 , new_n2820 , new_n2833 );
nor  g00486 ( new_n2835 , new_n2819 , new_n2834 );
and  g00487 ( new_n2836 , new_n2815 , new_n2835 );
nor  g00488 ( new_n2837 , new_n2813 , new_n2836 );
nor  g00489 ( new_n2838 , new_n2809_1 , new_n2837 );
nor  g00490 ( new_n2839 , new_n2808 , new_n2838 );
and  g00491 ( new_n2840 , new_n2805 , new_n2839 );
nor  g00492 ( new_n2841 , new_n2804 , new_n2840 );
and  g00493 ( new_n2842 , new_n2800 , new_n2841 );
nor  g00494 ( new_n2843 , new_n2799 , new_n2842 );
nor  g00495 ( new_n2844 , new_n2795 , new_n2843 );
nor  g00496 ( new_n2845 , new_n2794 , new_n2844 );
and  g00497 ( new_n2846 , new_n2790 , new_n2845 );
nor  g00498 ( new_n2847 , new_n2789 , new_n2846 );
xnor g00499 ( n108 , new_n2784 , new_n2847 );
xnor g00500 ( new_n2849 , n767 , n22379 );
not  g00501 ( new_n2850 , n1662 );
nor  g00502 ( new_n2851 , new_n2850 , n7330 );
xnor g00503 ( new_n2852 , n1662 , n7330 );
not  g00504 ( new_n2853_1 , n12875 );
nor  g00505 ( new_n2854 , new_n2853_1 , n22492 );
xnor g00506 ( new_n2855 , n12875 , n22492 );
not  g00507 ( new_n2856 , n2035 );
nor  g00508 ( new_n2857 , new_n2856 , n12821 );
xnor g00509 ( new_n2858_1 , n2035 , n12821 );
not  g00510 ( new_n2859 , n5213 );
nor  g00511 ( new_n2860_1 , n3468 , new_n2859 );
xnor g00512 ( new_n2861 , n3468 , n5213 );
not  g00513 ( new_n2862 , n4665 );
nor  g00514 ( new_n2863 , new_n2862 , n18558 );
xnor g00515 ( new_n2864 , n4665 , n18558 );
nor  g00516 ( new_n2865 , new_n2695 , n19005 );
not  g00517 ( new_n2866 , n19005 );
nor  g00518 ( new_n2867 , n7149 , new_n2866 );
nor  g00519 ( new_n2868 , n4326 , new_n2701 );
not  g00520 ( new_n2869 , n4326 );
or   g00521 ( new_n2870 , new_n2869 , n14148 );
nor  g00522 ( new_n2871 , new_n2698 , n5438 );
and  g00523 ( new_n2872 , new_n2870 , new_n2871 );
nor  g00524 ( new_n2873 , new_n2868 , new_n2872 );
nor  g00525 ( new_n2874 , new_n2867 , new_n2873 );
nor  g00526 ( new_n2875 , new_n2865 , new_n2874 );
and  g00527 ( new_n2876 , new_n2864 , new_n2875 );
or   g00528 ( new_n2877 , new_n2863 , new_n2876 );
and  g00529 ( new_n2878 , new_n2861 , new_n2877 );
or   g00530 ( new_n2879 , new_n2860_1 , new_n2878 );
and  g00531 ( new_n2880 , new_n2858_1 , new_n2879 );
or   g00532 ( new_n2881 , new_n2857 , new_n2880 );
and  g00533 ( new_n2882 , new_n2855 , new_n2881 );
or   g00534 ( new_n2883 , new_n2854 , new_n2882 );
and  g00535 ( new_n2884 , new_n2852 , new_n2883 );
or   g00536 ( new_n2885 , new_n2851 , new_n2884 );
xor  g00537 ( new_n2886_1 , new_n2849 , new_n2885 );
not  g00538 ( new_n2887_1 , n6814 );
xnor g00539 ( new_n2888 , new_n2887_1 , n10763 );
nor  g00540 ( new_n2889 , n7437 , n19701 );
not  g00541 ( new_n2890 , n7437 );
xnor g00542 ( new_n2891 , new_n2890 , n19701 );
nor  g00543 ( new_n2892 , n20700 , n23529 );
not  g00544 ( new_n2893 , n20700 );
xnor g00545 ( new_n2894 , new_n2893 , n23529 );
nor  g00546 ( new_n2895 , n7099 , n24620 );
not  g00547 ( new_n2896 , n7099 );
xnor g00548 ( new_n2897 , new_n2896 , n24620 );
nor  g00549 ( new_n2898 , n5211 , n12811 );
xnor g00550 ( new_n2899 , n5211 , n12811 );
nor  g00551 ( new_n2900 , n1118 , n12956 );
xnor g00552 ( new_n2901 , n1118 , n12956 );
nor  g00553 ( new_n2902 , n18295 , n25974 );
not  g00554 ( new_n2903 , n18295 );
xnor g00555 ( new_n2904 , new_n2903 , n25974 );
nor  g00556 ( new_n2905 , n1630 , n6502 );
not  g00557 ( new_n2906 , n1451 );
not  g00558 ( new_n2907 , n15780 );
or   g00559 ( new_n2908 , new_n2906 , new_n2907 );
not  g00560 ( new_n2909 , n1630 );
xnor g00561 ( new_n2910 , new_n2909 , n6502 );
and  g00562 ( new_n2911 , new_n2908 , new_n2910 );
or   g00563 ( new_n2912 , new_n2905 , new_n2911 );
and  g00564 ( new_n2913 , new_n2904 , new_n2912 );
nor  g00565 ( new_n2914 , new_n2902 , new_n2913 );
nor  g00566 ( new_n2915 , new_n2901 , new_n2914 );
nor  g00567 ( new_n2916 , new_n2900 , new_n2915 );
nor  g00568 ( new_n2917 , new_n2899 , new_n2916 );
or   g00569 ( new_n2918 , new_n2898 , new_n2917 );
and  g00570 ( new_n2919 , new_n2897 , new_n2918 );
or   g00571 ( new_n2920 , new_n2895 , new_n2919 );
and  g00572 ( new_n2921 , new_n2894 , new_n2920 );
or   g00573 ( new_n2922 , new_n2892 , new_n2921 );
and  g00574 ( new_n2923 , new_n2891 , new_n2922 );
or   g00575 ( new_n2924 , new_n2889 , new_n2923 );
xor  g00576 ( new_n2925 , new_n2888 , new_n2924 );
not  g00577 ( new_n2926 , n12657 );
xnor g00578 ( new_n2927 , new_n2926 , n27089 );
nor  g00579 ( new_n2928 , n11841 , n17077 );
not  g00580 ( new_n2929_1 , n11841 );
xnor g00581 ( new_n2930 , new_n2929_1 , n17077 );
not  g00582 ( new_n2931 , new_n2930 );
nor  g00583 ( new_n2932 , n10710 , n26510 );
not  g00584 ( new_n2933 , n10710 );
xnor g00585 ( new_n2934 , new_n2933 , n26510 );
not  g00586 ( new_n2935 , new_n2934 );
nor  g00587 ( new_n2936 , n20929 , n23068 );
not  g00588 ( new_n2937 , n20929 );
xnor g00589 ( new_n2938 , new_n2937 , n23068 );
not  g00590 ( new_n2939 , new_n2938 );
nor  g00591 ( new_n2940 , n8006 , n19514 );
not  g00592 ( new_n2941 , n8006 );
xnor g00593 ( new_n2942 , new_n2941 , n19514 );
nor  g00594 ( new_n2943 , n10053 , n25074 );
not  g00595 ( new_n2944_1 , n10053 );
xnor g00596 ( new_n2945 , new_n2944_1 , n25074 );
nor  g00597 ( new_n2946 , n8399 , n16396 );
not  g00598 ( new_n2947 , n8399 );
xnor g00599 ( new_n2948_1 , new_n2947 , n16396 );
not  g00600 ( new_n2949 , new_n2948_1 );
nor  g00601 ( new_n2950 , n9399 , n9507 );
not  g00602 ( new_n2951 , n2088 );
not  g00603 ( new_n2952 , n26979 );
nor  g00604 ( new_n2953 , new_n2951 , new_n2952 );
xnor g00605 ( new_n2954 , n9399 , n9507 );
nor  g00606 ( new_n2955 , new_n2953 , new_n2954 );
nor  g00607 ( new_n2956 , new_n2950 , new_n2955 );
nor  g00608 ( new_n2957 , new_n2949 , new_n2956 );
or   g00609 ( new_n2958 , new_n2946 , new_n2957 );
and  g00610 ( new_n2959 , new_n2945 , new_n2958 );
or   g00611 ( new_n2960 , new_n2943 , new_n2959 );
and  g00612 ( new_n2961_1 , new_n2942 , new_n2960 );
nor  g00613 ( new_n2962 , new_n2940 , new_n2961_1 );
nor  g00614 ( new_n2963 , new_n2939 , new_n2962 );
nor  g00615 ( new_n2964 , new_n2936 , new_n2963 );
nor  g00616 ( new_n2965 , new_n2935 , new_n2964 );
nor  g00617 ( new_n2966 , new_n2932 , new_n2965 );
nor  g00618 ( new_n2967 , new_n2931 , new_n2966 );
nor  g00619 ( new_n2968 , new_n2928 , new_n2967 );
xnor g00620 ( new_n2969 , new_n2927 , new_n2968 );
xnor g00621 ( new_n2970 , new_n2925 , new_n2969 );
nor  g00622 ( new_n2971_1 , new_n2892 , new_n2921 );
xnor g00623 ( new_n2972 , new_n2891 , new_n2971_1 );
xnor g00624 ( new_n2973 , new_n2930 , new_n2966 );
not  g00625 ( new_n2974 , new_n2973 );
nor  g00626 ( new_n2975 , new_n2972 , new_n2974 );
not  g00627 ( new_n2976 , new_n2972 );
xnor g00628 ( new_n2977 , new_n2976 , new_n2974 );
nor  g00629 ( new_n2978_1 , new_n2895 , new_n2919 );
xnor g00630 ( new_n2979_1 , new_n2894 , new_n2978_1 );
not  g00631 ( new_n2980 , new_n2979_1 );
xnor g00632 ( new_n2981 , new_n2934 , new_n2964 );
nor  g00633 ( new_n2982 , new_n2980 , new_n2981 );
xnor g00634 ( new_n2983 , new_n2980 , new_n2981 );
nor  g00635 ( new_n2984 , new_n2898 , new_n2917 );
xnor g00636 ( new_n2985_1 , new_n2897 , new_n2984 );
not  g00637 ( new_n2986 , new_n2985_1 );
xnor g00638 ( new_n2987 , new_n2938 , new_n2962 );
nor  g00639 ( new_n2988 , new_n2986 , new_n2987 );
xnor g00640 ( new_n2989 , new_n2986 , new_n2987 );
xnor g00641 ( new_n2990 , new_n2899 , new_n2916 );
nor  g00642 ( new_n2991 , new_n2943 , new_n2959 );
xnor g00643 ( new_n2992 , new_n2942 , new_n2991 );
nor  g00644 ( new_n2993 , new_n2990 , new_n2992 );
not  g00645 ( new_n2994 , new_n2992 );
xnor g00646 ( new_n2995 , new_n2990 , new_n2994 );
xnor g00647 ( new_n2996 , new_n2901 , new_n2914 );
nor  g00648 ( new_n2997 , new_n2946 , new_n2957 );
xnor g00649 ( new_n2998 , new_n2945 , new_n2997 );
nor  g00650 ( new_n2999_1 , new_n2996 , new_n2998 );
not  g00651 ( new_n3000 , new_n2998 );
xnor g00652 ( new_n3001 , new_n2996 , new_n3000 );
xor  g00653 ( new_n3002 , new_n2904 , new_n2912 );
xnor g00654 ( new_n3003 , new_n2948_1 , new_n2956 );
not  g00655 ( new_n3004 , new_n3003 );
nor  g00656 ( new_n3005 , new_n3002 , new_n3004 );
xnor g00657 ( new_n3006 , new_n3002 , new_n3003 );
nor  g00658 ( new_n3007 , new_n2906 , new_n2907 );
xnor g00659 ( new_n3008 , new_n3007 , new_n2910 );
not  g00660 ( new_n3009 , new_n3008 );
xnor g00661 ( new_n3010_1 , new_n2953 , new_n2954 );
not  g00662 ( new_n3011 , new_n3010_1 );
nor  g00663 ( new_n3012 , new_n3009 , new_n3011 );
xnor g00664 ( new_n3013 , new_n2906 , n15780 );
xnor g00665 ( new_n3014 , new_n2951 , n26979 );
not  g00666 ( new_n3015 , new_n3014 );
nor  g00667 ( new_n3016 , new_n3013 , new_n3015 );
xnor g00668 ( new_n3017_1 , new_n3009 , new_n3010_1 );
and  g00669 ( new_n3018_1 , new_n3016 , new_n3017_1 );
nor  g00670 ( new_n3019 , new_n3012 , new_n3018_1 );
and  g00671 ( new_n3020_1 , new_n3006 , new_n3019 );
nor  g00672 ( new_n3021 , new_n3005 , new_n3020_1 );
and  g00673 ( new_n3022 , new_n3001 , new_n3021 );
or   g00674 ( new_n3023 , new_n2999_1 , new_n3022 );
and  g00675 ( new_n3024 , new_n2995 , new_n3023 );
nor  g00676 ( new_n3025 , new_n2993 , new_n3024 );
nor  g00677 ( new_n3026 , new_n2989 , new_n3025 );
nor  g00678 ( new_n3027 , new_n2988 , new_n3026 );
nor  g00679 ( new_n3028 , new_n2983 , new_n3027 );
nor  g00680 ( new_n3029 , new_n2982 , new_n3028 );
and  g00681 ( new_n3030_1 , new_n2977 , new_n3029 );
or   g00682 ( new_n3031 , new_n2975 , new_n3030_1 );
xor  g00683 ( new_n3032 , new_n2970 , new_n3031 );
xnor g00684 ( new_n3033 , new_n2886_1 , new_n3032 );
xor  g00685 ( new_n3034 , new_n2852 , new_n2883 );
xor  g00686 ( new_n3035 , new_n2977 , new_n3029 );
nor  g00687 ( new_n3036 , new_n3034 , new_n3035 );
xnor g00688 ( new_n3037 , new_n3034 , new_n3035 );
xor  g00689 ( new_n3038 , new_n2855 , new_n2881 );
xnor g00690 ( new_n3039 , new_n2983 , new_n3027 );
nor  g00691 ( new_n3040 , new_n3038 , new_n3039 );
xnor g00692 ( new_n3041 , new_n3038 , new_n3039 );
xor  g00693 ( new_n3042 , new_n2858_1 , new_n2879 );
xnor g00694 ( new_n3043 , new_n2989 , new_n3025 );
nor  g00695 ( new_n3044 , new_n3042 , new_n3043 );
xnor g00696 ( new_n3045 , new_n3042 , new_n3043 );
xor  g00697 ( new_n3046 , new_n2861 , new_n2877 );
nor  g00698 ( new_n3047 , new_n2999_1 , new_n3022 );
xnor g00699 ( new_n3048 , new_n2995 , new_n3047 );
not  g00700 ( new_n3049 , new_n3048 );
nor  g00701 ( new_n3050 , new_n3046 , new_n3049 );
xnor g00702 ( new_n3051 , new_n3046 , new_n3049 );
xnor g00703 ( new_n3052 , new_n3001 , new_n3021 );
not  g00704 ( new_n3053 , new_n3052 );
xnor g00705 ( new_n3054 , new_n2864 , new_n2875 );
and  g00706 ( new_n3055 , new_n3053 , new_n3054 );
xnor g00707 ( new_n3056 , new_n3053 , new_n3054 );
xnor g00708 ( new_n3057 , new_n3006 , new_n3019 );
xnor g00709 ( new_n3058 , n7149 , n19005 );
xnor g00710 ( new_n3059 , new_n2873 , new_n3058 );
and  g00711 ( new_n3060 , new_n3057 , new_n3059 );
xnor g00712 ( new_n3061 , new_n3057 , new_n3059 );
xnor g00713 ( new_n3062 , n1152 , n5438 );
not  g00714 ( new_n3063 , new_n3013 );
xnor g00715 ( new_n3064 , new_n3063 , new_n3015 );
nor  g00716 ( new_n3065 , new_n3062 , new_n3064 );
xnor g00717 ( new_n3066 , n4326 , n14148 );
xnor g00718 ( new_n3067_1 , new_n2871 , new_n3066 );
nor  g00719 ( new_n3068 , new_n3065 , new_n3067_1 );
xnor g00720 ( new_n3069 , new_n3016 , new_n3017_1 );
xnor g00721 ( new_n3070 , new_n3065 , new_n3067_1 );
nor  g00722 ( new_n3071 , new_n3069 , new_n3070 );
nor  g00723 ( new_n3072 , new_n3068 , new_n3071 );
nor  g00724 ( new_n3073 , new_n3061 , new_n3072 );
nor  g00725 ( new_n3074 , new_n3060 , new_n3073 );
nor  g00726 ( new_n3075 , new_n3056 , new_n3074 );
nor  g00727 ( new_n3076_1 , new_n3055 , new_n3075 );
nor  g00728 ( new_n3077 , new_n3051 , new_n3076_1 );
nor  g00729 ( new_n3078 , new_n3050 , new_n3077 );
nor  g00730 ( new_n3079 , new_n3045 , new_n3078 );
nor  g00731 ( new_n3080 , new_n3044 , new_n3079 );
nor  g00732 ( new_n3081 , new_n3041 , new_n3080 );
nor  g00733 ( new_n3082 , new_n3040 , new_n3081 );
nor  g00734 ( new_n3083 , new_n3037 , new_n3082 );
nor  g00735 ( new_n3084 , new_n3036 , new_n3083 );
xnor g00736 ( n142 , new_n3033 , new_n3084 );
not  g00737 ( new_n3086 , n5025 );
not  g00738 ( new_n3087 , n4319 );
xnor g00739 ( new_n3088 , new_n3087 , n7335 );
not  g00740 ( new_n3089_1 , new_n3088 );
nor  g00741 ( new_n3090 , n5696 , n23463 );
not  g00742 ( new_n3091 , n5696 );
xnor g00743 ( new_n3092 , new_n3091 , n23463 );
not  g00744 ( new_n3093 , new_n3092 );
nor  g00745 ( new_n3094 , n13074 , n13367 );
not  g00746 ( new_n3095 , n13074 );
xnor g00747 ( new_n3096 , new_n3095 , n13367 );
not  g00748 ( new_n3097 , new_n3096 );
nor  g00749 ( new_n3098 , n932 , n10739 );
not  g00750 ( new_n3099 , n10739 );
xnor g00751 ( new_n3100 , n932 , new_n3099 );
not  g00752 ( new_n3101 , new_n3100 );
nor  g00753 ( new_n3102 , n6691 , n21753 );
xnor g00754 ( new_n3103 , n6691 , new_n2350 );
not  g00755 ( new_n3104 , new_n3103 );
nor  g00756 ( new_n3105 , n3260 , n21832 );
not  g00757 ( new_n3106 , n3260 );
xnor g00758 ( new_n3107 , new_n3106 , n21832 );
not  g00759 ( new_n3108 , new_n3107 );
nor  g00760 ( new_n3109 , n20489 , n26913 );
not  g00761 ( new_n3110 , n20489 );
xnor g00762 ( new_n3111 , new_n3110 , n26913 );
not  g00763 ( new_n3112 , new_n3111 );
nor  g00764 ( new_n3113 , n2355 , n16223 );
xnor g00765 ( new_n3114 , n2355 , n16223 );
nor  g00766 ( new_n3115 , n11121 , n19494 );
not  g00767 ( new_n3116 , n2387 );
not  g00768 ( new_n3117 , n16217 );
nor  g00769 ( new_n3118 , new_n3116 , new_n3117 );
xnor g00770 ( new_n3119 , n11121 , new_n2365 );
not  g00771 ( new_n3120 , new_n3119 );
nor  g00772 ( new_n3121 , new_n3118 , new_n3120 );
nor  g00773 ( new_n3122 , new_n3115 , new_n3121 );
nor  g00774 ( new_n3123 , new_n3114 , new_n3122 );
nor  g00775 ( new_n3124 , new_n3113 , new_n3123 );
nor  g00776 ( new_n3125_1 , new_n3112 , new_n3124 );
nor  g00777 ( new_n3126_1 , new_n3109 , new_n3125_1 );
nor  g00778 ( new_n3127 , new_n3108 , new_n3126_1 );
nor  g00779 ( new_n3128 , new_n3105 , new_n3127 );
nor  g00780 ( new_n3129 , new_n3104 , new_n3128 );
nor  g00781 ( new_n3130 , new_n3102 , new_n3129 );
nor  g00782 ( new_n3131 , new_n3101 , new_n3130 );
nor  g00783 ( new_n3132 , new_n3098 , new_n3131 );
nor  g00784 ( new_n3133 , new_n3097 , new_n3132 );
nor  g00785 ( new_n3134 , new_n3094 , new_n3133 );
nor  g00786 ( new_n3135 , new_n3093 , new_n3134 );
nor  g00787 ( new_n3136_1 , new_n3090 , new_n3135 );
xnor g00788 ( new_n3137 , new_n3089_1 , new_n3136_1 );
and  g00789 ( new_n3138 , new_n3086 , new_n3137 );
xnor g00790 ( new_n3139 , new_n3086 , new_n3137 );
not  g00791 ( new_n3140 , n6485 );
xnor g00792 ( new_n3141 , new_n3093 , new_n3134 );
and  g00793 ( new_n3142 , new_n3140 , new_n3141 );
xnor g00794 ( new_n3143 , new_n3140 , new_n3141 );
not  g00795 ( new_n3144 , n26036 );
xnor g00796 ( new_n3145 , new_n3097 , new_n3132 );
and  g00797 ( new_n3146 , new_n3144 , new_n3145 );
xnor g00798 ( new_n3147 , new_n3144 , new_n3145 );
not  g00799 ( new_n3148 , n19770 );
xnor g00800 ( new_n3149 , new_n3101 , new_n3130 );
and  g00801 ( new_n3150 , new_n3148 , new_n3149 );
xnor g00802 ( new_n3151 , new_n3148 , new_n3149 );
not  g00803 ( new_n3152 , n8782 );
xnor g00804 ( new_n3153 , new_n3104 , new_n3128 );
and  g00805 ( new_n3154 , new_n3152 , new_n3153 );
xnor g00806 ( new_n3155 , new_n3152 , new_n3153 );
not  g00807 ( new_n3156 , n8678 );
xnor g00808 ( new_n3157 , new_n3108 , new_n3126_1 );
and  g00809 ( new_n3158 , new_n3156 , new_n3157 );
xnor g00810 ( new_n3159 , new_n3156 , new_n3157 );
xnor g00811 ( new_n3160 , new_n3111 , new_n3124 );
nor  g00812 ( new_n3161_1 , n1432 , new_n3160 );
not  g00813 ( new_n3162 , n1432 );
not  g00814 ( new_n3163 , new_n3160 );
xnor g00815 ( new_n3164_1 , new_n3162 , new_n3163 );
xnor g00816 ( new_n3165 , new_n3114 , new_n3122 );
not  g00817 ( new_n3166 , new_n3165 );
nor  g00818 ( new_n3167 , n21599 , new_n3166 );
xnor g00819 ( new_n3168 , n21599 , new_n3166 );
not  g00820 ( new_n3169 , n25336 );
xnor g00821 ( new_n3170 , n2387 , n16217 );
nor  g00822 ( new_n3171 , n11424 , new_n3170 );
and  g00823 ( new_n3172 , new_n3169 , new_n3171 );
xnor g00824 ( new_n3173 , new_n3169 , new_n3171 );
xnor g00825 ( new_n3174 , new_n3118 , new_n3119 );
nor  g00826 ( new_n3175 , new_n3173 , new_n3174 );
nor  g00827 ( new_n3176 , new_n3172 , new_n3175 );
nor  g00828 ( new_n3177 , new_n3168 , new_n3176 );
nor  g00829 ( new_n3178 , new_n3167 , new_n3177 );
nor  g00830 ( new_n3179 , new_n3164_1 , new_n3178 );
nor  g00831 ( new_n3180 , new_n3161_1 , new_n3179 );
nor  g00832 ( new_n3181 , new_n3159 , new_n3180 );
nor  g00833 ( new_n3182 , new_n3158 , new_n3181 );
nor  g00834 ( new_n3183 , new_n3155 , new_n3182 );
nor  g00835 ( new_n3184 , new_n3154 , new_n3183 );
nor  g00836 ( new_n3185 , new_n3151 , new_n3184 );
nor  g00837 ( new_n3186 , new_n3150 , new_n3185 );
nor  g00838 ( new_n3187 , new_n3147 , new_n3186 );
nor  g00839 ( new_n3188 , new_n3146 , new_n3187 );
nor  g00840 ( new_n3189 , new_n3143 , new_n3188 );
nor  g00841 ( new_n3190 , new_n3142 , new_n3189 );
nor  g00842 ( new_n3191 , new_n3139 , new_n3190 );
nor  g00843 ( new_n3192 , new_n3138 , new_n3191 );
nor  g00844 ( new_n3193 , n4319 , n7335 );
nor  g00845 ( new_n3194 , new_n3089_1 , new_n3136_1 );
nor  g00846 ( new_n3195 , new_n3193 , new_n3194 );
not  g00847 ( new_n3196 , new_n3195 );
nand g00848 ( new_n3197 , new_n3192 , new_n3196 );
not  g00849 ( new_n3198 , n9967 );
nor  g00850 ( new_n3199 , n3952 , n12315 );
not  g00851 ( new_n3200 , new_n3199 );
nor  g00852 ( new_n3201 , n24618 , new_n3200 );
not  g00853 ( new_n3202 , new_n3201 );
nor  g00854 ( new_n3203 , n24278 , new_n3202 );
not  g00855 ( new_n3204 , new_n3203 );
nor  g00856 ( new_n3205 , n4812 , new_n3204 );
not  g00857 ( new_n3206 , new_n3205 );
nor  g00858 ( new_n3207 , n26823 , new_n3206 );
not  g00859 ( new_n3208_1 , new_n3207 );
nor  g00860 ( new_n3209 , n7751 , new_n3208_1 );
not  g00861 ( new_n3210 , new_n3209 );
nor  g00862 ( new_n3211 , n20946 , new_n3210 );
and  g00863 ( new_n3212 , new_n3198 , new_n3211 );
xnor g00864 ( new_n3213 , n3425 , new_n3212 );
not  g00865 ( new_n3214 , new_n3213 );
xor  g00866 ( new_n3215 , new_n3139 , new_n3190 );
nor  g00867 ( new_n3216 , new_n3214 , new_n3215 );
not  g00868 ( new_n3217 , n3425 );
and  g00869 ( new_n3218 , new_n3217 , new_n3212 );
xnor g00870 ( new_n3219_1 , new_n3214 , new_n3215 );
xnor g00871 ( new_n3220 , n9967 , new_n3211 );
not  g00872 ( new_n3221 , new_n3220 );
xor  g00873 ( new_n3222 , new_n3143 , new_n3188 );
nor  g00874 ( new_n3223 , new_n3221 , new_n3222 );
not  g00875 ( new_n3224 , new_n3222 );
xnor g00876 ( new_n3225 , new_n3220 , new_n3224 );
xnor g00877 ( new_n3226 , n20946 , new_n3209 );
not  g00878 ( new_n3227 , new_n3226 );
xor  g00879 ( new_n3228_1 , new_n3147 , new_n3186 );
nor  g00880 ( new_n3229 , new_n3227 , new_n3228_1 );
xnor g00881 ( new_n3230 , new_n3227 , new_n3228_1 );
xnor g00882 ( new_n3231 , n7751 , new_n3207 );
not  g00883 ( new_n3232 , new_n3231 );
xor  g00884 ( new_n3233 , new_n3151 , new_n3184 );
nor  g00885 ( new_n3234 , new_n3232 , new_n3233 );
xnor g00886 ( new_n3235_1 , new_n3232 , new_n3233 );
xnor g00887 ( new_n3236 , n26823 , new_n3205 );
not  g00888 ( new_n3237 , new_n3236 );
xor  g00889 ( new_n3238 , new_n3155 , new_n3182 );
nor  g00890 ( new_n3239 , new_n3237 , new_n3238 );
xnor g00891 ( new_n3240 , new_n3237 , new_n3238 );
xnor g00892 ( new_n3241 , n4812 , new_n3203 );
not  g00893 ( new_n3242 , new_n3241 );
xor  g00894 ( new_n3243 , new_n3159 , new_n3180 );
nor  g00895 ( new_n3244_1 , new_n3242 , new_n3243 );
xnor g00896 ( new_n3245 , new_n3242 , new_n3243 );
xnor g00897 ( new_n3246 , n24278 , new_n3201 );
not  g00898 ( new_n3247 , new_n3246 );
xor  g00899 ( new_n3248 , new_n3164_1 , new_n3178 );
nor  g00900 ( new_n3249 , new_n3247 , new_n3248 );
xnor g00901 ( new_n3250 , new_n3247 , new_n3248 );
xnor g00902 ( new_n3251 , n24618 , new_n3199 );
not  g00903 ( new_n3252 , new_n3251 );
xor  g00904 ( new_n3253_1 , new_n3168 , new_n3176 );
nor  g00905 ( new_n3254 , new_n3252 , new_n3253_1 );
xnor g00906 ( new_n3255 , new_n3252 , new_n3253_1 );
not  g00907 ( new_n3256 , n11424 );
xnor g00908 ( new_n3257 , new_n3256 , new_n3170 );
nor  g00909 ( new_n3258 , new_n2448 , new_n3257 );
and  g00910 ( new_n3259 , new_n2443 , new_n3258 );
xnor g00911 ( new_n3260_1 , new_n3118 , new_n3120 );
xnor g00912 ( new_n3261 , new_n3173 , new_n3260_1 );
xnor g00913 ( new_n3262 , new_n2443 , n12315 );
nor  g00914 ( new_n3263_1 , new_n3258 , new_n3262 );
or   g00915 ( new_n3264 , new_n3259 , new_n3263_1 );
nor  g00916 ( new_n3265 , new_n3261 , new_n3264 );
nor  g00917 ( new_n3266 , new_n3259 , new_n3265 );
nor  g00918 ( new_n3267 , new_n3255 , new_n3266 );
nor  g00919 ( new_n3268 , new_n3254 , new_n3267 );
nor  g00920 ( new_n3269 , new_n3250 , new_n3268 );
nor  g00921 ( new_n3270 , new_n3249 , new_n3269 );
nor  g00922 ( new_n3271 , new_n3245 , new_n3270 );
nor  g00923 ( new_n3272 , new_n3244_1 , new_n3271 );
nor  g00924 ( new_n3273 , new_n3240 , new_n3272 );
nor  g00925 ( new_n3274 , new_n3239 , new_n3273 );
nor  g00926 ( new_n3275 , new_n3235_1 , new_n3274 );
nor  g00927 ( new_n3276 , new_n3234 , new_n3275 );
nor  g00928 ( new_n3277 , new_n3230 , new_n3276 );
nor  g00929 ( new_n3278 , new_n3229 , new_n3277 );
nor  g00930 ( new_n3279_1 , new_n3225 , new_n3278 );
nor  g00931 ( new_n3280 , new_n3223 , new_n3279_1 );
nor  g00932 ( new_n3281 , new_n3219_1 , new_n3280 );
or   g00933 ( new_n3282 , new_n3218 , new_n3281 );
nor  g00934 ( new_n3283 , new_n3216 , new_n3282 );
not  g00935 ( new_n3284 , new_n3283 );
nor  g00936 ( new_n3285 , new_n3197 , new_n3284 );
nor  g00937 ( new_n3286 , n5101 , n7593 );
xnor g00938 ( new_n3287 , n5101 , n7593 );
nor  g00939 ( new_n3288 , n337 , n16507 );
xnor g00940 ( new_n3289_1 , n337 , n16507 );
nor  g00941 ( new_n3290 , n3228 , n22470 );
xnor g00942 ( new_n3291 , n3228 , n22470 );
nor  g00943 ( new_n3292 , n5302 , n19116 );
xnor g00944 ( new_n3293 , n5302 , n19116 );
nor  g00945 ( new_n3294 , n6861 , n25738 );
xnor g00946 ( new_n3295 , n6861 , n25738 );
nor  g00947 ( new_n3296 , n19357 , n21471 );
xnor g00948 ( new_n3297 , n19357 , n21471 );
nor  g00949 ( new_n3298 , n2328 , n18737 );
xnor g00950 ( new_n3299 , n2328 , n18737 );
nor  g00951 ( new_n3300 , n14603 , n15053 );
not  g00952 ( new_n3301_1 , n14603 );
xnor g00953 ( new_n3302 , new_n3301_1 , n15053 );
nor  g00954 ( new_n3303 , n20794 , n25471 );
not  g00955 ( new_n3304 , n16502 );
not  g00956 ( new_n3305 , n23333 );
nor  g00957 ( new_n3306_1 , new_n3304 , new_n3305 );
not  g00958 ( new_n3307 , n20794 );
xnor g00959 ( new_n3308 , new_n3307 , n25471 );
not  g00960 ( new_n3309 , new_n3308 );
nor  g00961 ( new_n3310 , new_n3306_1 , new_n3309 );
or   g00962 ( new_n3311 , new_n3303 , new_n3310 );
and  g00963 ( new_n3312 , new_n3302 , new_n3311 );
nor  g00964 ( new_n3313 , new_n3300 , new_n3312 );
nor  g00965 ( new_n3314 , new_n3299 , new_n3313 );
nor  g00966 ( new_n3315 , new_n3298 , new_n3314 );
nor  g00967 ( new_n3316_1 , new_n3297 , new_n3315 );
nor  g00968 ( new_n3317 , new_n3296 , new_n3316_1 );
nor  g00969 ( new_n3318 , new_n3295 , new_n3317 );
nor  g00970 ( new_n3319 , new_n3294 , new_n3318 );
nor  g00971 ( new_n3320_1 , new_n3293 , new_n3319 );
nor  g00972 ( new_n3321 , new_n3292 , new_n3320_1 );
nor  g00973 ( new_n3322 , new_n3291 , new_n3321 );
nor  g00974 ( new_n3323 , new_n3290 , new_n3322 );
nor  g00975 ( new_n3324_1 , new_n3289_1 , new_n3323 );
nor  g00976 ( new_n3325 , new_n3288 , new_n3324_1 );
nor  g00977 ( new_n3326 , new_n3287 , new_n3325 );
nor  g00978 ( new_n3327 , new_n3286 , new_n3326 );
xnor g00979 ( new_n3328 , new_n3192 , new_n3196 );
not  g00980 ( new_n3329 , new_n3328 );
xnor g00981 ( new_n3330 , new_n3284 , new_n3329 );
and  g00982 ( new_n3331 , new_n3327 , new_n3330 );
nor  g00983 ( new_n3332_1 , new_n3327 , new_n3330 );
xor  g00984 ( new_n3333 , new_n3219_1 , new_n3280 );
xnor g00985 ( new_n3334 , new_n3287 , new_n3325 );
nor  g00986 ( new_n3335 , new_n3333 , new_n3334 );
xnor g00987 ( new_n3336 , new_n3333 , new_n3334 );
xor  g00988 ( new_n3337 , new_n3225 , new_n3278 );
xnor g00989 ( new_n3338 , new_n3289_1 , new_n3323 );
nor  g00990 ( new_n3339 , new_n3337 , new_n3338 );
xnor g00991 ( new_n3340_1 , new_n3337 , new_n3338 );
xor  g00992 ( new_n3341 , new_n3230 , new_n3276 );
xnor g00993 ( new_n3342 , new_n3291 , new_n3321 );
nor  g00994 ( new_n3343_1 , new_n3341 , new_n3342 );
xnor g00995 ( new_n3344 , new_n3341 , new_n3342 );
xor  g00996 ( new_n3345 , new_n3235_1 , new_n3274 );
xnor g00997 ( new_n3346 , new_n3293 , new_n3319 );
nor  g00998 ( new_n3347 , new_n3345 , new_n3346 );
xnor g00999 ( new_n3348 , new_n3345 , new_n3346 );
xor  g01000 ( new_n3349_1 , new_n3240 , new_n3272 );
xnor g01001 ( new_n3350 , new_n3295 , new_n3317 );
nor  g01002 ( new_n3351 , new_n3349_1 , new_n3350 );
xnor g01003 ( new_n3352 , new_n3349_1 , new_n3350 );
xor  g01004 ( new_n3353 , new_n3245 , new_n3270 );
xnor g01005 ( new_n3354 , new_n3297 , new_n3315 );
nor  g01006 ( new_n3355 , new_n3353 , new_n3354 );
xnor g01007 ( new_n3356 , new_n3353 , new_n3354 );
xor  g01008 ( new_n3357 , new_n3250 , new_n3268 );
xnor g01009 ( new_n3358 , new_n3299 , new_n3313 );
nor  g01010 ( new_n3359 , new_n3357 , new_n3358 );
xnor g01011 ( new_n3360 , new_n3357 , new_n3358 );
xor  g01012 ( new_n3361 , new_n3255 , new_n3266 );
nor  g01013 ( new_n3362 , new_n3303 , new_n3310 );
xnor g01014 ( new_n3363 , new_n3302 , new_n3362 );
not  g01015 ( new_n3364 , new_n3363 );
nor  g01016 ( new_n3365 , new_n3361 , new_n3364 );
xnor g01017 ( new_n3366_1 , new_n3361 , new_n3364 );
xnor g01018 ( new_n3367 , new_n3304 , n23333 );
xnor g01019 ( new_n3368 , n12315 , new_n3257 );
and  g01020 ( new_n3369 , new_n3367 , new_n3368 );
xnor g01021 ( new_n3370 , new_n3306_1 , new_n3309 );
nor  g01022 ( new_n3371 , new_n3369 , new_n3370 );
xor  g01023 ( new_n3372 , new_n3261 , new_n3264 );
not  g01024 ( new_n3373 , new_n3372 );
and  g01025 ( new_n3374 , new_n3308 , new_n3369 );
nor  g01026 ( new_n3375 , new_n3371 , new_n3374 );
and  g01027 ( new_n3376 , new_n3373 , new_n3375 );
nor  g01028 ( new_n3377 , new_n3371 , new_n3376 );
nor  g01029 ( new_n3378 , new_n3366_1 , new_n3377 );
nor  g01030 ( new_n3379 , new_n3365 , new_n3378 );
nor  g01031 ( new_n3380 , new_n3360 , new_n3379 );
nor  g01032 ( new_n3381 , new_n3359 , new_n3380 );
nor  g01033 ( new_n3382 , new_n3356 , new_n3381 );
nor  g01034 ( new_n3383 , new_n3355 , new_n3382 );
nor  g01035 ( new_n3384 , new_n3352 , new_n3383 );
nor  g01036 ( new_n3385 , new_n3351 , new_n3384 );
nor  g01037 ( new_n3386 , new_n3348 , new_n3385 );
nor  g01038 ( new_n3387 , new_n3347 , new_n3386 );
nor  g01039 ( new_n3388 , new_n3344 , new_n3387 );
nor  g01040 ( new_n3389 , new_n3343_1 , new_n3388 );
nor  g01041 ( new_n3390_1 , new_n3340_1 , new_n3389 );
nor  g01042 ( new_n3391 , new_n3339 , new_n3390_1 );
nor  g01043 ( new_n3392 , new_n3336 , new_n3391 );
or   g01044 ( new_n3393 , new_n3335 , new_n3392 );
nor  g01045 ( new_n3394 , new_n3332_1 , new_n3393 );
nor  g01046 ( new_n3395 , new_n3331 , new_n3394 );
not  g01047 ( new_n3396 , new_n3395 );
and  g01048 ( new_n3397 , new_n3285 , new_n3396 );
nor  g01049 ( new_n3398 , new_n3197 , new_n3283 );
or   g01050 ( new_n3399 , new_n3192 , new_n3196 );
nor  g01051 ( new_n3400 , new_n3284 , new_n3399 );
or   g01052 ( new_n3401 , new_n3398 , new_n3400 );
nor  g01053 ( new_n3402 , new_n3395 , new_n3401 );
nor  g01054 ( new_n3403 , new_n3285 , new_n3402 );
nor  g01055 ( n175 , new_n3397 , new_n3403 );
not  g01056 ( new_n3405 , n14130 );
nor  g01057 ( new_n3406 , n9251 , n20138 );
not  g01058 ( new_n3407 , new_n3406 );
nor  g01059 ( new_n3408 , n6385 , new_n3407 );
not  g01060 ( new_n3409 , new_n3408 );
nor  g01061 ( new_n3410 , n3136 , new_n3409 );
not  g01062 ( new_n3411 , new_n3410 );
nor  g01063 ( new_n3412 , n9557 , new_n3411 );
not  g01064 ( new_n3413 , new_n3412 );
nor  g01065 ( new_n3414 , n25643 , new_n3413 );
not  g01066 ( new_n3415 , new_n3414 );
nor  g01067 ( new_n3416 , n9942 , new_n3415 );
not  g01068 ( new_n3417 , new_n3416 );
nor  g01069 ( new_n3418 , n16482 , new_n3417 );
and  g01070 ( new_n3419 , new_n3405 , new_n3418 );
xnor g01071 ( new_n3420 , n8856 , new_n3419 );
xnor g01072 ( new_n3421 , n25494 , new_n3420 );
xnor g01073 ( new_n3422 , n14130 , new_n3418 );
nor  g01074 ( new_n3423 , n10117 , new_n3422 );
not  g01075 ( new_n3424 , n10117 );
xnor g01076 ( new_n3425_1 , new_n3424 , new_n3422 );
xnor g01077 ( new_n3426_1 , n16482 , new_n3416 );
nor  g01078 ( new_n3427 , n13460 , new_n3426_1 );
not  g01079 ( new_n3428 , n13460 );
xnor g01080 ( new_n3429 , new_n3428 , new_n3426_1 );
xnor g01081 ( new_n3430 , n9942 , new_n3414 );
nor  g01082 ( new_n3431 , n6104 , new_n3430 );
not  g01083 ( new_n3432 , n6104 );
xnor g01084 ( new_n3433 , new_n3432 , new_n3430 );
xnor g01085 ( new_n3434 , n25643 , new_n3412 );
nor  g01086 ( new_n3435 , n4119 , new_n3434 );
not  g01087 ( new_n3436 , n4119 );
xnor g01088 ( new_n3437 , new_n3436 , new_n3434 );
xnor g01089 ( new_n3438 , n9557 , new_n3410 );
nor  g01090 ( new_n3439 , n14510 , new_n3438 );
not  g01091 ( new_n3440 , n14510 );
xnor g01092 ( new_n3441 , new_n3440 , new_n3438 );
xnor g01093 ( new_n3442 , n3136 , new_n3408 );
nor  g01094 ( new_n3443 , n13263 , new_n3442 );
xnor g01095 ( new_n3444 , n6385 , new_n3406 );
nor  g01096 ( new_n3445 , n20455 , new_n3444 );
not  g01097 ( new_n3446 , n20455 );
xnor g01098 ( new_n3447 , new_n3446 , new_n3444 );
not  g01099 ( new_n3448 , n1639 );
xnor g01100 ( new_n3449 , n9251 , n20138 );
and  g01101 ( new_n3450 , new_n3448 , new_n3449 );
not  g01102 ( new_n3451_1 , n16968 );
or   g01103 ( new_n3452 , new_n2367 , new_n3451_1 );
xnor g01104 ( new_n3453 , n1639 , new_n3449 );
and  g01105 ( new_n3454 , new_n3452 , new_n3453 );
or   g01106 ( new_n3455 , new_n3450 , new_n3454 );
and  g01107 ( new_n3456 , new_n3447 , new_n3455 );
or   g01108 ( new_n3457 , new_n3445 , new_n3456 );
not  g01109 ( new_n3458 , n13263 );
xnor g01110 ( new_n3459_1 , new_n3458 , new_n3442 );
and  g01111 ( new_n3460_1 , new_n3457 , new_n3459_1 );
or   g01112 ( new_n3461 , new_n3443 , new_n3460_1 );
and  g01113 ( new_n3462 , new_n3441 , new_n3461 );
or   g01114 ( new_n3463 , new_n3439 , new_n3462 );
and  g01115 ( new_n3464 , new_n3437 , new_n3463 );
or   g01116 ( new_n3465 , new_n3435 , new_n3464 );
and  g01117 ( new_n3466 , new_n3433 , new_n3465 );
or   g01118 ( new_n3467 , new_n3431 , new_n3466 );
and  g01119 ( new_n3468_1 , new_n3429 , new_n3467 );
or   g01120 ( new_n3469 , new_n3427 , new_n3468_1 );
and  g01121 ( new_n3470 , new_n3425_1 , new_n3469 );
nor  g01122 ( new_n3471 , new_n3423 , new_n3470 );
xnor g01123 ( new_n3472 , new_n3421 , new_n3471 );
xnor g01124 ( new_n3473 , n26180 , new_n3472 );
nor  g01125 ( new_n3474 , new_n3427 , new_n3468_1 );
xnor g01126 ( new_n3475 , new_n3425_1 , new_n3474 );
not  g01127 ( new_n3476 , new_n3475 );
nor  g01128 ( new_n3477 , n24004 , new_n3476 );
xnor g01129 ( new_n3478 , n24004 , new_n3475 );
nor  g01130 ( new_n3479 , new_n3431 , new_n3466 );
xnor g01131 ( new_n3480_1 , new_n3429 , new_n3479 );
not  g01132 ( new_n3481 , new_n3480_1 );
nor  g01133 ( new_n3482 , n12871 , new_n3481 );
xnor g01134 ( new_n3483 , n12871 , new_n3480_1 );
nor  g01135 ( new_n3484 , new_n3435 , new_n3464 );
xnor g01136 ( new_n3485 , new_n3433 , new_n3484 );
not  g01137 ( new_n3486 , new_n3485 );
nor  g01138 ( new_n3487 , n23304 , new_n3486 );
xnor g01139 ( new_n3488 , n23304 , new_n3485 );
nor  g01140 ( new_n3489 , new_n3439 , new_n3462 );
xnor g01141 ( new_n3490 , new_n3437 , new_n3489 );
not  g01142 ( new_n3491 , new_n3490 );
nor  g01143 ( new_n3492 , n19361 , new_n3491 );
xnor g01144 ( new_n3493 , n19361 , new_n3490 );
xor  g01145 ( new_n3494 , new_n3441 , new_n3461 );
not  g01146 ( new_n3495 , new_n3494 );
nor  g01147 ( new_n3496 , n1437 , new_n3495 );
not  g01148 ( new_n3497 , n1437 );
xnor g01149 ( new_n3498 , new_n3497 , new_n3495 );
nor  g01150 ( new_n3499 , new_n3445 , new_n3456 );
xnor g01151 ( new_n3500 , new_n3499 , new_n3459_1 );
not  g01152 ( new_n3501 , new_n3500 );
nor  g01153 ( new_n3502_1 , n4722 , new_n3501 );
not  g01154 ( new_n3503 , n4722 );
xnor g01155 ( new_n3504 , new_n3503 , new_n3501 );
not  g01156 ( new_n3505 , n14633 );
nor  g01157 ( new_n3506_1 , new_n3450 , new_n3454 );
xnor g01158 ( new_n3507 , new_n3447 , new_n3506_1 );
nor  g01159 ( new_n3508 , new_n3505 , new_n3507 );
not  g01160 ( new_n3509 , new_n3507 );
xnor g01161 ( new_n3510 , new_n3505 , new_n3509 );
not  g01162 ( new_n3511 , n8721 );
nor  g01163 ( new_n3512 , new_n2367 , new_n3451_1 );
xnor g01164 ( new_n3513 , new_n3512 , new_n3453 );
nor  g01165 ( new_n3514 , new_n3511 , new_n3513 );
not  g01166 ( new_n3515 , n18578 );
xnor g01167 ( new_n3516_1 , n9251 , n16968 );
nor  g01168 ( new_n3517 , new_n3515 , new_n3516_1 );
xnor g01169 ( new_n3518 , n8721 , new_n3513 );
and  g01170 ( new_n3519 , new_n3517 , new_n3518 );
or   g01171 ( new_n3520 , new_n3514 , new_n3519 );
and  g01172 ( new_n3521 , new_n3510 , new_n3520 );
nor  g01173 ( new_n3522 , new_n3508 , new_n3521 );
and  g01174 ( new_n3523 , new_n3504 , new_n3522 );
or   g01175 ( new_n3524 , new_n3502_1 , new_n3523 );
and  g01176 ( new_n3525 , new_n3498 , new_n3524 );
or   g01177 ( new_n3526 , new_n3496 , new_n3525 );
and  g01178 ( new_n3527 , new_n3493 , new_n3526 );
or   g01179 ( new_n3528_1 , new_n3492 , new_n3527 );
and  g01180 ( new_n3529 , new_n3488 , new_n3528_1 );
or   g01181 ( new_n3530 , new_n3487 , new_n3529 );
and  g01182 ( new_n3531 , new_n3483 , new_n3530 );
or   g01183 ( new_n3532 , new_n3482 , new_n3531 );
and  g01184 ( new_n3533 , new_n3478 , new_n3532 );
nor  g01185 ( new_n3534 , new_n3477 , new_n3533 );
xnor g01186 ( new_n3535 , new_n3473 , new_n3534 );
xnor g01187 ( new_n3536 , n2743 , n3506 );
not  g01188 ( new_n3537 , n7026 );
nor  g01189 ( new_n3538 , new_n3537 , n14899 );
xnor g01190 ( new_n3539 , n7026 , n14899 );
not  g01191 ( new_n3540 , n13719 );
nor  g01192 ( new_n3541_1 , new_n3540 , n18444 );
xnor g01193 ( new_n3542 , n13719 , n18444 );
not  g01194 ( new_n3543 , n442 );
nor  g01195 ( new_n3544 , new_n3543 , n24638 );
xnor g01196 ( new_n3545 , n442 , n24638 );
not  g01197 ( new_n3546 , n9172 );
nor  g01198 ( new_n3547 , new_n3546 , n21674 );
xnor g01199 ( new_n3548 , n9172 , n21674 );
not  g01200 ( new_n3549 , n4913 );
nor  g01201 ( new_n3550 , new_n3549 , n17251 );
xnor g01202 ( new_n3551 , n4913 , n17251 );
not  g01203 ( new_n3552 , n604 );
nor  g01204 ( new_n3553 , new_n3552 , n14790 );
xnor g01205 ( new_n3554 , n604 , n14790 );
not  g01206 ( new_n3555_1 , n10096 );
nor  g01207 ( new_n3556 , new_n3555_1 , n16824 );
and  g01208 ( new_n3557 , new_n3555_1 , n16824 );
not  g01209 ( new_n3558 , n16994 );
nor  g01210 ( new_n3559 , n16521 , new_n3558 );
not  g01211 ( new_n3560 , n16521 );
nor  g01212 ( new_n3561_1 , new_n3560 , n16994 );
not  g01213 ( new_n3562 , n9246 );
nor  g01214 ( new_n3563_1 , n7139 , new_n3562 );
not  g01215 ( new_n3564 , new_n3563_1 );
nor  g01216 ( new_n3565 , new_n3561_1 , new_n3564 );
nor  g01217 ( new_n3566 , new_n3559 , new_n3565 );
nor  g01218 ( new_n3567 , new_n3557 , new_n3566 );
nor  g01219 ( new_n3568 , new_n3556 , new_n3567 );
and  g01220 ( new_n3569 , new_n3554 , new_n3568 );
or   g01221 ( new_n3570_1 , new_n3553 , new_n3569 );
and  g01222 ( new_n3571 , new_n3551 , new_n3570_1 );
or   g01223 ( new_n3572 , new_n3550 , new_n3571 );
and  g01224 ( new_n3573 , new_n3548 , new_n3572 );
or   g01225 ( new_n3574 , new_n3547 , new_n3573 );
and  g01226 ( new_n3575 , new_n3545 , new_n3574 );
or   g01227 ( new_n3576 , new_n3544 , new_n3575 );
and  g01228 ( new_n3577 , new_n3542 , new_n3576 );
or   g01229 ( new_n3578 , new_n3541_1 , new_n3577 );
and  g01230 ( new_n3579 , new_n3539 , new_n3578 );
or   g01231 ( new_n3580 , new_n3538 , new_n3579 );
xor  g01232 ( new_n3581 , new_n3536 , new_n3580 );
not  g01233 ( new_n3582_1 , new_n3581 );
not  g01234 ( new_n3583 , n21489 );
nor  g01235 ( new_n3584 , n21993 , n25565 );
not  g01236 ( new_n3585 , new_n3584 );
nor  g01237 ( new_n3586 , n11273 , new_n3585 );
not  g01238 ( new_n3587 , new_n3586 );
nor  g01239 ( new_n3588 , n22290 , new_n3587 );
not  g01240 ( new_n3589 , new_n3588 );
nor  g01241 ( new_n3590 , n9598 , new_n3589 );
not  g01242 ( new_n3591 , new_n3590 );
nor  g01243 ( new_n3592 , n7670 , new_n3591 );
not  g01244 ( new_n3593 , new_n3592 );
nor  g01245 ( new_n3594 , n13912 , new_n3593 );
not  g01246 ( new_n3595 , new_n3594 );
nor  g01247 ( new_n3596 , n20213 , new_n3595 );
and  g01248 ( new_n3597 , new_n3583 , new_n3596 );
xnor g01249 ( new_n3598 , n9259 , new_n3597 );
xnor g01250 ( new_n3599 , new_n3582_1 , new_n3598 );
xor  g01251 ( new_n3600 , new_n3539 , new_n3578 );
not  g01252 ( new_n3601 , new_n3600 );
xnor g01253 ( new_n3602 , n21489 , new_n3596 );
not  g01254 ( new_n3603 , new_n3602 );
nor  g01255 ( new_n3604 , new_n3601 , new_n3603 );
xnor g01256 ( new_n3605 , new_n3601 , new_n3602 );
nor  g01257 ( new_n3606 , new_n3544 , new_n3575 );
xnor g01258 ( new_n3607 , new_n3542 , new_n3606 );
xnor g01259 ( new_n3608 , n20213 , new_n3594 );
nor  g01260 ( new_n3609 , new_n3607 , new_n3608 );
not  g01261 ( new_n3610 , new_n3607 );
not  g01262 ( new_n3611 , new_n3608 );
xnor g01263 ( new_n3612 , new_n3610 , new_n3611 );
xor  g01264 ( new_n3613 , new_n3545 , new_n3574 );
xnor g01265 ( new_n3614 , n13912 , new_n3592 );
nor  g01266 ( new_n3615 , new_n3613 , new_n3614 );
xnor g01267 ( new_n3616 , new_n3613 , new_n3614 );
xor  g01268 ( new_n3617_1 , new_n3548 , new_n3572 );
xnor g01269 ( new_n3618_1 , n7670 , new_n3590 );
nor  g01270 ( new_n3619 , new_n3617_1 , new_n3618_1 );
xnor g01271 ( new_n3620 , new_n3617_1 , new_n3618_1 );
xnor g01272 ( new_n3621 , n9598 , new_n3588 );
xor  g01273 ( new_n3622 , new_n3551 , new_n3570_1 );
nor  g01274 ( new_n3623 , new_n3621 , new_n3622 );
xnor g01275 ( new_n3624 , new_n3621 , new_n3622 );
xnor g01276 ( new_n3625 , n22290 , new_n3586 );
not  g01277 ( new_n3626 , new_n3625 );
xnor g01278 ( new_n3627 , new_n3554 , new_n3568 );
and  g01279 ( new_n3628 , new_n3626 , new_n3627 );
xnor g01280 ( new_n3629 , n11273 , new_n3584 );
not  g01281 ( new_n3630 , new_n3629 );
xnor g01282 ( new_n3631 , n10096 , n16824 );
xnor g01283 ( new_n3632 , new_n3566 , new_n3631 );
and  g01284 ( new_n3633 , new_n3630 , new_n3632 );
xnor g01285 ( new_n3634 , new_n3629 , new_n3632 );
not  g01286 ( new_n3635 , n21993 );
xnor g01287 ( new_n3636 , new_n3635 , n25565 );
xnor g01288 ( new_n3637 , n16521 , n16994 );
xnor g01289 ( new_n3638 , new_n3564 , new_n3637 );
not  g01290 ( new_n3639 , new_n3638 );
nor  g01291 ( new_n3640 , new_n3636 , new_n3639 );
xnor g01292 ( new_n3641 , n7139 , n9246 );
nor  g01293 ( new_n3642_1 , new_n3635 , new_n3641 );
not  g01294 ( new_n3643 , new_n3636 );
xnor g01295 ( new_n3644 , new_n3643 , new_n3638 );
nor  g01296 ( new_n3645 , new_n3642_1 , new_n3644 );
or   g01297 ( new_n3646 , new_n3640 , new_n3645 );
and  g01298 ( new_n3647 , new_n3634 , new_n3646 );
or   g01299 ( new_n3648 , new_n3633 , new_n3647 );
xnor g01300 ( new_n3649_1 , new_n3625 , new_n3627 );
and  g01301 ( new_n3650 , new_n3648 , new_n3649_1 );
nor  g01302 ( new_n3651 , new_n3628 , new_n3650 );
nor  g01303 ( new_n3652 , new_n3624 , new_n3651 );
nor  g01304 ( new_n3653 , new_n3623 , new_n3652 );
nor  g01305 ( new_n3654 , new_n3620 , new_n3653 );
nor  g01306 ( new_n3655 , new_n3619 , new_n3654 );
nor  g01307 ( new_n3656 , new_n3616 , new_n3655 );
nor  g01308 ( new_n3657 , new_n3615 , new_n3656 );
nor  g01309 ( new_n3658 , new_n3612 , new_n3657 );
nor  g01310 ( new_n3659 , new_n3609 , new_n3658 );
and  g01311 ( new_n3660 , new_n3605 , new_n3659 );
or   g01312 ( new_n3661 , new_n3604 , new_n3660 );
xor  g01313 ( new_n3662 , new_n3599 , new_n3661 );
xnor g01314 ( new_n3663 , new_n3535 , new_n3662 );
nor  g01315 ( new_n3664 , new_n3482 , new_n3531 );
xnor g01316 ( new_n3665_1 , new_n3478 , new_n3664 );
not  g01317 ( new_n3666 , new_n3665_1 );
xor  g01318 ( new_n3667 , new_n3605 , new_n3659 );
nor  g01319 ( new_n3668 , new_n3666 , new_n3667 );
xnor g01320 ( new_n3669 , new_n3666 , new_n3667 );
xor  g01321 ( new_n3670 , new_n3483 , new_n3530 );
not  g01322 ( new_n3671 , new_n3670 );
xnor g01323 ( new_n3672 , new_n3612 , new_n3657 );
nor  g01324 ( new_n3673 , new_n3671 , new_n3672 );
xnor g01325 ( new_n3674 , new_n3671 , new_n3672 );
xor  g01326 ( new_n3675 , new_n3488 , new_n3528_1 );
not  g01327 ( new_n3676 , new_n3675 );
xnor g01328 ( new_n3677 , new_n3616 , new_n3655 );
nor  g01329 ( new_n3678 , new_n3676 , new_n3677 );
xnor g01330 ( new_n3679_1 , new_n3676 , new_n3677 );
xor  g01331 ( new_n3680 , new_n3493 , new_n3526 );
not  g01332 ( new_n3681 , new_n3680 );
xnor g01333 ( new_n3682 , new_n3620 , new_n3653 );
nor  g01334 ( new_n3683 , new_n3681 , new_n3682 );
xnor g01335 ( new_n3684 , new_n3681 , new_n3682 );
xor  g01336 ( new_n3685 , new_n3498 , new_n3524 );
not  g01337 ( new_n3686 , new_n3685 );
xnor g01338 ( new_n3687 , new_n3624 , new_n3651 );
nor  g01339 ( new_n3688 , new_n3686 , new_n3687 );
xnor g01340 ( new_n3689 , new_n3686 , new_n3687 );
xnor g01341 ( new_n3690 , new_n3504 , new_n3522 );
not  g01342 ( new_n3691 , new_n3690 );
xor  g01343 ( new_n3692 , new_n3648 , new_n3649_1 );
and  g01344 ( new_n3693 , new_n3691 , new_n3692 );
xnor g01345 ( new_n3694 , new_n3691 , new_n3692 );
nor  g01346 ( new_n3695 , new_n3514 , new_n3519 );
xnor g01347 ( new_n3696 , new_n3510 , new_n3695 );
not  g01348 ( new_n3697 , new_n3696 );
xor  g01349 ( new_n3698 , new_n3634 , new_n3646 );
and  g01350 ( new_n3699 , new_n3697 , new_n3698 );
xnor g01351 ( new_n3700 , new_n3697 , new_n3698 );
xnor g01352 ( new_n3701 , new_n3642_1 , new_n3644 );
xor  g01353 ( new_n3702 , new_n3517 , new_n3518 );
nor  g01354 ( new_n3703 , new_n3701 , new_n3702 );
xnor g01355 ( new_n3704 , n18578 , new_n3516_1 );
xnor g01356 ( new_n3705 , n21993 , new_n3641 );
and  g01357 ( new_n3706 , new_n3704 , new_n3705 );
xnor g01358 ( new_n3707 , new_n3701 , new_n3702 );
nor  g01359 ( new_n3708 , new_n3706 , new_n3707 );
nor  g01360 ( new_n3709 , new_n3703 , new_n3708 );
nor  g01361 ( new_n3710_1 , new_n3700 , new_n3709 );
nor  g01362 ( new_n3711 , new_n3699 , new_n3710_1 );
nor  g01363 ( new_n3712 , new_n3694 , new_n3711 );
nor  g01364 ( new_n3713 , new_n3693 , new_n3712 );
nor  g01365 ( new_n3714 , new_n3689 , new_n3713 );
nor  g01366 ( new_n3715 , new_n3688 , new_n3714 );
nor  g01367 ( new_n3716 , new_n3684 , new_n3715 );
nor  g01368 ( new_n3717 , new_n3683 , new_n3716 );
nor  g01369 ( new_n3718 , new_n3679_1 , new_n3717 );
nor  g01370 ( new_n3719 , new_n3678 , new_n3718 );
nor  g01371 ( new_n3720 , new_n3674 , new_n3719 );
nor  g01372 ( new_n3721 , new_n3673 , new_n3720 );
nor  g01373 ( new_n3722 , new_n3669 , new_n3721 );
nor  g01374 ( new_n3723 , new_n3668 , new_n3722 );
xnor g01375 ( n235 , new_n3663 , new_n3723 );
not  g01376 ( new_n3725_1 , n25749 );
not  g01377 ( new_n3726 , n19327 );
nor  g01378 ( new_n3727 , n13319 , n25435 );
not  g01379 ( new_n3728 , new_n3727 );
nor  g01380 ( new_n3729 , n15967 , new_n3728 );
not  g01381 ( new_n3730 , new_n3729 );
nor  g01382 ( new_n3731 , n25797 , new_n3730 );
not  g01383 ( new_n3732 , new_n3731 );
nor  g01384 ( new_n3733_1 , n6369 , new_n3732 );
not  g01385 ( new_n3734 , new_n3733_1 );
nor  g01386 ( new_n3735 , n21134 , new_n3734 );
xnor g01387 ( new_n3736 , n2113 , new_n3735 );
xnor g01388 ( new_n3737 , new_n3726 , new_n3736 );
xnor g01389 ( new_n3738 , n21134 , new_n3733_1 );
nor  g01390 ( new_n3739 , n22597 , new_n3738 );
not  g01391 ( new_n3740_1 , n22597 );
xnor g01392 ( new_n3741 , new_n3740_1 , new_n3738 );
xnor g01393 ( new_n3742 , n6369 , new_n3731 );
nor  g01394 ( new_n3743 , n26107 , new_n3742 );
not  g01395 ( new_n3744 , n26107 );
xnor g01396 ( new_n3745 , new_n3744 , new_n3742 );
xnor g01397 ( new_n3746 , n25797 , new_n3729 );
nor  g01398 ( new_n3747 , n342 , new_n3746 );
xnor g01399 ( new_n3748 , n15967 , new_n3727 );
nor  g01400 ( new_n3749 , n26553 , new_n3748 );
not  g01401 ( new_n3750 , new_n3748 );
xnor g01402 ( new_n3751 , n26553 , new_n3750 );
not  g01403 ( new_n3752 , n13319 );
xnor g01404 ( new_n3753 , new_n3752 , n25435 );
nor  g01405 ( new_n3754 , n4964 , new_n3753 );
not  g01406 ( new_n3755_1 , n7876 );
not  g01407 ( new_n3756 , n25435 );
or   g01408 ( new_n3757 , new_n3755_1 , new_n3756 );
not  g01409 ( new_n3758_1 , new_n3753 );
xnor g01410 ( new_n3759 , n4964 , new_n3758_1 );
and  g01411 ( new_n3760_1 , new_n3757 , new_n3759 );
or   g01412 ( new_n3761 , new_n3754 , new_n3760_1 );
and  g01413 ( new_n3762 , new_n3751 , new_n3761 );
or   g01414 ( new_n3763 , new_n3749 , new_n3762 );
xor  g01415 ( new_n3764 , n342 , new_n3746 );
and  g01416 ( new_n3765 , new_n3763 , new_n3764 );
or   g01417 ( new_n3766 , new_n3747 , new_n3765 );
and  g01418 ( new_n3767 , new_n3745 , new_n3766 );
or   g01419 ( new_n3768 , new_n3743 , new_n3767 );
and  g01420 ( new_n3769 , new_n3741 , new_n3768 );
nor  g01421 ( new_n3770 , new_n3739 , new_n3769 );
xnor g01422 ( new_n3771 , new_n3737 , new_n3770 );
not  g01423 ( new_n3772 , new_n3771 );
xnor g01424 ( new_n3773 , new_n3725_1 , new_n3772 );
not  g01425 ( new_n3774 , n3161 );
xor  g01426 ( new_n3775 , new_n3741 , new_n3768 );
nor  g01427 ( new_n3776 , new_n3774 , new_n3775 );
xnor g01428 ( new_n3777 , n3161 , new_n3775 );
not  g01429 ( new_n3778 , n9003 );
nor  g01430 ( new_n3779 , new_n3747 , new_n3765 );
xnor g01431 ( new_n3780 , new_n3745 , new_n3779 );
nor  g01432 ( new_n3781_1 , new_n3778 , new_n3780 );
not  g01433 ( new_n3782 , new_n3780 );
xnor g01434 ( new_n3783 , new_n3778 , new_n3782 );
not  g01435 ( new_n3784 , n4957 );
xor  g01436 ( new_n3785_1 , new_n3763 , new_n3764 );
nor  g01437 ( new_n3786 , new_n3784 , new_n3785_1 );
xnor g01438 ( new_n3787 , n4957 , new_n3785_1 );
not  g01439 ( new_n3788 , n7524 );
nor  g01440 ( new_n3789 , new_n3754 , new_n3760_1 );
xnor g01441 ( new_n3790 , new_n3751 , new_n3789 );
nor  g01442 ( new_n3791 , new_n3788 , new_n3790 );
not  g01443 ( new_n3792 , new_n3790 );
xnor g01444 ( new_n3793 , new_n3788 , new_n3792 );
not  g01445 ( new_n3794_1 , n15743 );
nor  g01446 ( new_n3795_1 , new_n3755_1 , new_n3756 );
xnor g01447 ( new_n3796 , new_n3795_1 , new_n3759 );
nor  g01448 ( new_n3797 , new_n3794_1 , new_n3796 );
not  g01449 ( new_n3798 , n20658 );
xnor g01450 ( new_n3799 , new_n3755_1 , n25435 );
not  g01451 ( new_n3800 , new_n3799 );
nor  g01452 ( new_n3801 , new_n3798 , new_n3800 );
xnor g01453 ( new_n3802 , n15743 , new_n3796 );
and  g01454 ( new_n3803 , new_n3801 , new_n3802 );
or   g01455 ( new_n3804 , new_n3797 , new_n3803 );
and  g01456 ( new_n3805 , new_n3793 , new_n3804 );
or   g01457 ( new_n3806 , new_n3791 , new_n3805 );
and  g01458 ( new_n3807 , new_n3787 , new_n3806 );
or   g01459 ( new_n3808 , new_n3786 , new_n3807 );
and  g01460 ( new_n3809 , new_n3783 , new_n3808 );
or   g01461 ( new_n3810 , new_n3781_1 , new_n3809 );
and  g01462 ( new_n3811 , new_n3777 , new_n3810 );
or   g01463 ( new_n3812 , new_n3776 , new_n3811 );
xor  g01464 ( new_n3813 , new_n3773 , new_n3812 );
xnor g01465 ( new_n3814 , n22332 , n26510 );
not  g01466 ( new_n3815 , n23068 );
and  g01467 ( new_n3816 , n18907 , new_n3815 );
xnor g01468 ( new_n3817 , n18907 , n23068 );
nor  g01469 ( new_n3818 , new_n2408 , n19514 );
xnor g01470 ( new_n3819 , n2731 , n19514 );
and  g01471 ( new_n3820 , new_n2944_1 , n19911 );
xnor g01472 ( new_n3821 , n10053 , n19911 );
nor  g01473 ( new_n3822 , new_n2947 , n13708 );
nor  g01474 ( new_n3823 , n8399 , new_n2389 );
not  g01475 ( new_n3824 , n9507 );
nor  g01476 ( new_n3825 , new_n3824 , n18409 );
not  g01477 ( new_n3826 , n18409 );
nor  g01478 ( new_n3827 , n9507 , new_n3826 );
nor  g01479 ( new_n3828_1 , n5704 , new_n2952 );
not  g01480 ( new_n3829 , new_n3828_1 );
nor  g01481 ( new_n3830 , new_n3827 , new_n3829 );
nor  g01482 ( new_n3831 , new_n3825 , new_n3830 );
nor  g01483 ( new_n3832 , new_n3823 , new_n3831 );
nor  g01484 ( new_n3833 , new_n3822 , new_n3832 );
and  g01485 ( new_n3834 , new_n3821 , new_n3833 );
or   g01486 ( new_n3835 , new_n3820 , new_n3834 );
and  g01487 ( new_n3836 , new_n3819 , new_n3835 );
or   g01488 ( new_n3837 , new_n3818 , new_n3836 );
and  g01489 ( new_n3838 , new_n3817 , new_n3837 );
or   g01490 ( new_n3839 , new_n3816 , new_n3838 );
xor  g01491 ( new_n3840 , new_n3814 , new_n3839 );
nor  g01492 ( new_n3841 , n12121 , n22043 );
not  g01493 ( new_n3842_1 , new_n3841 );
nor  g01494 ( new_n3843 , n19618 , new_n3842_1 );
not  g01495 ( new_n3844 , new_n3843 );
nor  g01496 ( new_n3845 , n1204 , new_n3844 );
not  g01497 ( new_n3846 , new_n3845 );
nor  g01498 ( new_n3847 , n626 , new_n3846 );
not  g01499 ( new_n3848 , new_n3847 );
nor  g01500 ( new_n3849 , n5337 , new_n3848 );
xnor g01501 ( new_n3850_1 , n4325 , new_n3849 );
xnor g01502 ( new_n3851 , new_n3840 , new_n3850_1 );
xor  g01503 ( new_n3852 , new_n3817 , new_n3837 );
xnor g01504 ( new_n3853 , n5337 , new_n3847 );
nor  g01505 ( new_n3854 , new_n3852 , new_n3853 );
xnor g01506 ( new_n3855 , new_n3852 , new_n3853 );
xor  g01507 ( new_n3856 , new_n3819 , new_n3835 );
xnor g01508 ( new_n3857 , n626 , new_n3845 );
nor  g01509 ( new_n3858 , new_n3856 , new_n3857 );
xnor g01510 ( new_n3859 , new_n3856 , new_n3857 );
xnor g01511 ( new_n3860 , n1204 , new_n3843 );
xnor g01512 ( new_n3861 , new_n3821 , new_n3833 );
not  g01513 ( new_n3862 , new_n3861 );
nor  g01514 ( new_n3863 , new_n3860 , new_n3862 );
xnor g01515 ( new_n3864 , new_n3860 , new_n3861 );
xnor g01516 ( new_n3865 , n19618 , new_n3841 );
xnor g01517 ( new_n3866 , n8399 , n13708 );
xnor g01518 ( new_n3867 , new_n3831 , new_n3866 );
not  g01519 ( new_n3868 , new_n3867 );
nor  g01520 ( new_n3869_1 , new_n3865 , new_n3868 );
xnor g01521 ( new_n3870 , new_n3865 , new_n3867 );
xnor g01522 ( new_n3871_1 , n12121 , n22043 );
xnor g01523 ( new_n3872 , n9507 , n18409 );
xnor g01524 ( new_n3873 , new_n3829 , new_n3872 );
nor  g01525 ( new_n3874 , new_n3871_1 , new_n3873 );
not  g01526 ( new_n3875 , n12121 );
xnor g01527 ( new_n3876 , n5704 , n26979 );
nor  g01528 ( new_n3877 , new_n3875 , new_n3876 );
xor  g01529 ( new_n3878 , new_n3871_1 , new_n3873 );
and  g01530 ( new_n3879 , new_n3877 , new_n3878 );
nor  g01531 ( new_n3880 , new_n3874 , new_n3879 );
and  g01532 ( new_n3881 , new_n3870 , new_n3880 );
or   g01533 ( new_n3882 , new_n3869_1 , new_n3881 );
and  g01534 ( new_n3883 , new_n3864 , new_n3882 );
nor  g01535 ( new_n3884 , new_n3863 , new_n3883 );
nor  g01536 ( new_n3885 , new_n3859 , new_n3884 );
nor  g01537 ( new_n3886 , new_n3858 , new_n3885 );
nor  g01538 ( new_n3887 , new_n3855 , new_n3886 );
nor  g01539 ( new_n3888 , new_n3854 , new_n3887 );
xnor g01540 ( new_n3889 , new_n3851 , new_n3888 );
xnor g01541 ( new_n3890 , new_n3813 , new_n3889 );
xnor g01542 ( new_n3891_1 , new_n3855 , new_n3886 );
xor  g01543 ( new_n3892 , new_n3777 , new_n3810 );
nor  g01544 ( new_n3893 , new_n3891_1 , new_n3892 );
xnor g01545 ( new_n3894 , new_n3891_1 , new_n3892 );
xnor g01546 ( new_n3895 , new_n3859 , new_n3884 );
xor  g01547 ( new_n3896 , new_n3783 , new_n3808 );
nor  g01548 ( new_n3897 , new_n3895 , new_n3896 );
xnor g01549 ( new_n3898 , new_n3895 , new_n3896 );
xor  g01550 ( new_n3899 , new_n3864 , new_n3882 );
not  g01551 ( new_n3900 , new_n3899 );
xor  g01552 ( new_n3901 , new_n3787 , new_n3806 );
nor  g01553 ( new_n3902 , new_n3900 , new_n3901 );
xnor g01554 ( new_n3903 , new_n3900 , new_n3901 );
xnor g01555 ( new_n3904 , new_n3870 , new_n3880 );
xor  g01556 ( new_n3905 , new_n3793 , new_n3804 );
nor  g01557 ( new_n3906 , new_n3904 , new_n3905 );
xnor g01558 ( new_n3907 , new_n3904 , new_n3905 );
xnor g01559 ( new_n3908 , new_n3877 , new_n3878 );
not  g01560 ( new_n3909_1 , new_n3908 );
xor  g01561 ( new_n3910 , new_n3801 , new_n3802 );
nor  g01562 ( new_n3911 , new_n3909_1 , new_n3910 );
xnor g01563 ( new_n3912 , new_n3798 , new_n3800 );
xnor g01564 ( new_n3913 , n12121 , new_n3876 );
not  g01565 ( new_n3914 , new_n3913 );
nor  g01566 ( new_n3915 , new_n3912 , new_n3914 );
xnor g01567 ( new_n3916 , new_n3909_1 , new_n3910 );
nor  g01568 ( new_n3917 , new_n3915 , new_n3916 );
nor  g01569 ( new_n3918_1 , new_n3911 , new_n3917 );
nor  g01570 ( new_n3919 , new_n3907 , new_n3918_1 );
nor  g01571 ( new_n3920 , new_n3906 , new_n3919 );
nor  g01572 ( new_n3921 , new_n3903 , new_n3920 );
nor  g01573 ( new_n3922 , new_n3902 , new_n3921 );
nor  g01574 ( new_n3923 , new_n3898 , new_n3922 );
nor  g01575 ( new_n3924 , new_n3897 , new_n3923 );
nor  g01576 ( new_n3925_1 , new_n3894 , new_n3924 );
nor  g01577 ( new_n3926 , new_n3893 , new_n3925_1 );
xnor g01578 ( n242 , new_n3890 , new_n3926 );
nor  g01579 ( new_n3928 , n11667 , n21398 );
not  g01580 ( new_n3929 , new_n3928 );
nor  g01581 ( new_n3930 , n26572 , new_n3929 );
not  g01582 ( new_n3931 , new_n3930 );
nor  g01583 ( new_n3932_1 , n5115 , new_n3931 );
not  g01584 ( new_n3933 , new_n3932_1 );
nor  g01585 ( new_n3934_1 , n11223 , new_n3933 );
xnor g01586 ( new_n3935 , n19477 , new_n3934_1 );
xnor g01587 ( new_n3936 , n11011 , new_n3935 );
xnor g01588 ( new_n3937 , n11223 , new_n3932_1 );
nor  g01589 ( new_n3938 , n16029 , new_n3937 );
not  g01590 ( new_n3939 , n16029 );
xnor g01591 ( new_n3940 , new_n3939 , new_n3937 );
xnor g01592 ( new_n3941 , n5115 , new_n3930 );
and  g01593 ( new_n3942 , n16476 , new_n3941 );
not  g01594 ( new_n3943 , n16476 );
xnor g01595 ( new_n3944 , new_n3943 , new_n3941 );
xnor g01596 ( new_n3945_1 , n26572 , new_n3928 );
nor  g01597 ( new_n3946 , n11615 , new_n3945_1 );
not  g01598 ( new_n3947 , n11615 );
xnor g01599 ( new_n3948 , new_n3947 , new_n3945_1 );
not  g01600 ( new_n3949 , n22433 );
xnor g01601 ( new_n3950 , n11667 , n21398 );
and  g01602 ( new_n3951 , new_n3949 , new_n3950 );
not  g01603 ( new_n3952_1 , n14090 );
or   g01604 ( new_n3953 , new_n3952_1 , new_n2583 );
xnor g01605 ( new_n3954 , n22433 , new_n3950 );
and  g01606 ( new_n3955 , new_n3953 , new_n3954 );
or   g01607 ( new_n3956 , new_n3951 , new_n3955 );
and  g01608 ( new_n3957 , new_n3948 , new_n3956 );
nor  g01609 ( new_n3958 , new_n3946 , new_n3957 );
and  g01610 ( new_n3959_1 , new_n3944 , new_n3958 );
nor  g01611 ( new_n3960 , new_n3942 , new_n3959_1 );
and  g01612 ( new_n3961 , new_n3940 , new_n3960 );
nor  g01613 ( new_n3962_1 , new_n3938 , new_n3961 );
xnor g01614 ( new_n3963 , new_n3936 , new_n3962_1 );
xnor g01615 ( new_n3964 , n13677 , new_n3963 );
xnor g01616 ( new_n3965 , new_n3940 , new_n3960 );
nor  g01617 ( new_n3966 , n18926 , new_n3965 );
not  g01618 ( new_n3967 , n5451 );
xnor g01619 ( new_n3968 , new_n3944 , new_n3958 );
nor  g01620 ( new_n3969 , new_n3967 , new_n3968 );
not  g01621 ( new_n3970 , new_n3968 );
xnor g01622 ( new_n3971_1 , new_n3967 , new_n3970 );
not  g01623 ( new_n3972 , n5330 );
nor  g01624 ( new_n3973 , new_n3951 , new_n3955 );
xnor g01625 ( new_n3974 , new_n3948 , new_n3973 );
nor  g01626 ( new_n3975 , new_n3972 , new_n3974 );
not  g01627 ( new_n3976 , new_n3974 );
xnor g01628 ( new_n3977 , new_n3972 , new_n3976 );
not  g01629 ( new_n3978 , n7657 );
nor  g01630 ( new_n3979 , new_n3952_1 , new_n2583 );
xnor g01631 ( new_n3980 , new_n3979 , new_n3954 );
nor  g01632 ( new_n3981 , new_n3978 , new_n3980 );
not  g01633 ( new_n3982 , n25926 );
nor  g01634 ( new_n3983_1 , new_n3982 , new_n2551 );
not  g01635 ( new_n3984_1 , new_n3980 );
xnor g01636 ( new_n3985 , new_n3978 , new_n3984_1 );
and  g01637 ( new_n3986 , new_n3983_1 , new_n3985 );
or   g01638 ( new_n3987 , new_n3981 , new_n3986 );
and  g01639 ( new_n3988 , new_n3977 , new_n3987 );
or   g01640 ( new_n3989 , new_n3975 , new_n3988 );
and  g01641 ( new_n3990 , new_n3971_1 , new_n3989 );
nor  g01642 ( new_n3991 , new_n3969 , new_n3990 );
not  g01643 ( new_n3992 , new_n3991 );
xnor g01644 ( new_n3993 , n18926 , new_n3965 );
nor  g01645 ( new_n3994 , new_n3992 , new_n3993 );
nor  g01646 ( new_n3995 , new_n3966 , new_n3994 );
xnor g01647 ( new_n3996 , new_n3964 , new_n3995 );
nor  g01648 ( new_n3997 , n6729 , n21687 );
not  g01649 ( new_n3998 , new_n3997 );
nor  g01650 ( new_n3999 , n8285 , new_n3998 );
not  g01651 ( new_n4000_1 , new_n3999 );
nor  g01652 ( new_n4001 , n20169 , new_n4000_1 );
not  g01653 ( new_n4002 , new_n4001 );
nor  g01654 ( new_n4003 , n19789 , new_n4002 );
xnor g01655 ( new_n4004 , n12398 , new_n4003 );
nor  g01656 ( new_n4005 , n10792 , n19922 );
not  g01657 ( new_n4006 , new_n4005 );
nor  g01658 ( new_n4007 , n9323 , new_n4006 );
not  g01659 ( new_n4008 , new_n4007 );
nor  g01660 ( new_n4009 , n1949 , new_n4008 );
not  g01661 ( new_n4010_1 , new_n4009 );
nor  g01662 ( new_n4011 , n15424 , new_n4010_1 );
xnor g01663 ( new_n4012 , n25694 , new_n4011 );
not  g01664 ( new_n4013 , new_n4012 );
xnor g01665 ( new_n4014_1 , n20151 , new_n4013 );
not  g01666 ( new_n4015 , n7693 );
xnor g01667 ( new_n4016 , n15424 , new_n4009 );
not  g01668 ( new_n4017 , new_n4016 );
nor  g01669 ( new_n4018 , new_n4015 , new_n4017 );
xnor g01670 ( new_n4019 , n1949 , new_n4007 );
and  g01671 ( new_n4020 , n10405 , new_n4019 );
not  g01672 ( new_n4021 , n10405 );
xnor g01673 ( new_n4022 , new_n4021 , new_n4019 );
xnor g01674 ( new_n4023 , n9323 , new_n4005 );
nor  g01675 ( new_n4024 , n11302 , new_n4023 );
not  g01676 ( new_n4025 , new_n4023 );
xnor g01677 ( new_n4026 , n11302 , new_n4025 );
xnor g01678 ( new_n4027 , n10792 , n19922 );
not  g01679 ( new_n4028 , new_n4027 );
nor  g01680 ( new_n4029 , n17090 , new_n4028 );
not  g01681 ( new_n4030 , n6773 );
not  g01682 ( new_n4031 , n19922 );
or   g01683 ( new_n4032 , new_n4030 , new_n4031 );
xnor g01684 ( new_n4033 , n17090 , new_n4027 );
and  g01685 ( new_n4034 , new_n4032 , new_n4033 );
or   g01686 ( new_n4035 , new_n4029 , new_n4034 );
and  g01687 ( new_n4036 , new_n4026 , new_n4035 );
nor  g01688 ( new_n4037 , new_n4024 , new_n4036 );
and  g01689 ( new_n4038 , new_n4022 , new_n4037 );
or   g01690 ( new_n4039 , new_n4020 , new_n4038 );
xnor g01691 ( new_n4040 , n7693 , new_n4017 );
and  g01692 ( new_n4041 , new_n4039 , new_n4040 );
nor  g01693 ( new_n4042 , new_n4018 , new_n4041 );
xnor g01694 ( new_n4043 , new_n4014_1 , new_n4042 );
not  g01695 ( new_n4044 , new_n4043 );
xnor g01696 ( new_n4045 , new_n4004 , new_n4044 );
xnor g01697 ( new_n4046 , n19789 , new_n4001 );
xor  g01698 ( new_n4047 , new_n4039 , new_n4040 );
and  g01699 ( new_n4048 , new_n4046 , new_n4047 );
not  g01700 ( new_n4049 , new_n4047 );
xnor g01701 ( new_n4050 , new_n4046 , new_n4049 );
xnor g01702 ( new_n4051 , new_n4022 , new_n4037 );
not  g01703 ( new_n4052 , new_n4051 );
xnor g01704 ( new_n4053 , n20169 , new_n3999 );
nor  g01705 ( new_n4054 , new_n4052 , new_n4053 );
xnor g01706 ( new_n4055 , new_n4051 , new_n4053 );
nor  g01707 ( new_n4056 , new_n4029 , new_n4034 );
xnor g01708 ( new_n4057 , new_n4026 , new_n4056 );
not  g01709 ( new_n4058 , new_n4057 );
xnor g01710 ( new_n4059 , n8285 , new_n3997 );
and  g01711 ( new_n4060 , new_n4058 , new_n4059 );
xnor g01712 ( new_n4061 , new_n4057 , new_n4059 );
xnor g01713 ( new_n4062 , n6729 , n21687 );
nor  g01714 ( new_n4063 , new_n4030 , new_n4031 );
xnor g01715 ( new_n4064 , new_n4063 , new_n4033 );
nor  g01716 ( new_n4065 , new_n4062 , new_n4064 );
nor  g01717 ( new_n4066 , new_n2548 , new_n2549 );
not  g01718 ( new_n4067 , new_n4064 );
xnor g01719 ( new_n4068 , new_n4062 , new_n4067 );
and  g01720 ( new_n4069 , new_n4066 , new_n4068 );
or   g01721 ( new_n4070 , new_n4065 , new_n4069 );
and  g01722 ( new_n4071_1 , new_n4061 , new_n4070 );
nor  g01723 ( new_n4072 , new_n4060 , new_n4071_1 );
and  g01724 ( new_n4073 , new_n4055 , new_n4072 );
nor  g01725 ( new_n4074 , new_n4054 , new_n4073 );
and  g01726 ( new_n4075 , new_n4050 , new_n4074 );
or   g01727 ( new_n4076 , new_n4048 , new_n4075 );
xor  g01728 ( new_n4077 , new_n4045 , new_n4076 );
xnor g01729 ( new_n4078 , new_n3996 , new_n4077 );
xnor g01730 ( new_n4079 , new_n4050 , new_n4074 );
xnor g01731 ( new_n4080 , new_n3991 , new_n3993 );
and  g01732 ( new_n4081 , new_n4079 , new_n4080 );
xnor g01733 ( new_n4082 , new_n4079 , new_n4080 );
xnor g01734 ( new_n4083 , new_n4055 , new_n4072 );
xor  g01735 ( new_n4084 , new_n3971_1 , new_n3989 );
nor  g01736 ( new_n4085_1 , new_n4083 , new_n4084 );
xnor g01737 ( new_n4086 , new_n4083 , new_n4084 );
xor  g01738 ( new_n4087 , new_n3977 , new_n3987 );
xor  g01739 ( new_n4088_1 , new_n4061 , new_n4070 );
nor  g01740 ( new_n4089_1 , new_n4087 , new_n4088_1 );
xnor g01741 ( new_n4090 , new_n4087 , new_n4088_1 );
xor  g01742 ( new_n4091 , new_n4066 , new_n4068 );
xor  g01743 ( new_n4092 , new_n3983_1 , new_n3985 );
nor  g01744 ( new_n4093 , new_n4091 , new_n4092 );
not  g01745 ( new_n4094 , new_n2552 );
nor  g01746 ( new_n4095 , new_n2550 , new_n4094 );
xnor g01747 ( new_n4096 , new_n4091 , new_n4092 );
nor  g01748 ( new_n4097 , new_n4095 , new_n4096 );
nor  g01749 ( new_n4098 , new_n4093 , new_n4097 );
nor  g01750 ( new_n4099 , new_n4090 , new_n4098 );
nor  g01751 ( new_n4100_1 , new_n4089_1 , new_n4099 );
nor  g01752 ( new_n4101 , new_n4086 , new_n4100_1 );
nor  g01753 ( new_n4102 , new_n4085_1 , new_n4101 );
nor  g01754 ( new_n4103_1 , new_n4082 , new_n4102 );
nor  g01755 ( new_n4104 , new_n4081 , new_n4103_1 );
xnor g01756 ( n243 , new_n4078 , new_n4104 );
not  g01757 ( new_n4106 , n11302 );
xnor g01758 ( new_n4107 , new_n4106 , n24786 );
nor  g01759 ( new_n4108 , n17090 , n27120 );
not  g01760 ( new_n4109 , n23065 );
or   g01761 ( new_n4110 , new_n4030 , new_n4109 );
not  g01762 ( new_n4111 , n17090 );
xnor g01763 ( new_n4112 , new_n4111 , n27120 );
and  g01764 ( new_n4113 , new_n4110 , new_n4112 );
nor  g01765 ( new_n4114 , new_n4108 , new_n4113 );
xnor g01766 ( new_n4115 , new_n4107 , new_n4114 );
not  g01767 ( new_n4116 , new_n4115 );
xnor g01768 ( new_n4117 , n1689 , n20036 );
not  g01769 ( new_n4118 , n22274 );
nor  g01770 ( new_n4119_1 , n11192 , new_n4118 );
not  g01771 ( new_n4120 , n11192 );
nor  g01772 ( new_n4121 , new_n4120 , n22274 );
not  g01773 ( new_n4122 , n24129 );
nor  g01774 ( new_n4123_1 , n9380 , new_n4122 );
not  g01775 ( new_n4124 , new_n4123_1 );
nor  g01776 ( new_n4125 , new_n4121 , new_n4124 );
nor  g01777 ( new_n4126 , new_n4119_1 , new_n4125 );
xnor g01778 ( new_n4127 , new_n4117 , new_n4126 );
xnor g01779 ( new_n4128 , new_n4116 , new_n4127 );
nor  g01780 ( new_n4129 , new_n4030 , new_n4109 );
xnor g01781 ( new_n4130 , new_n4129 , new_n4112 );
xnor g01782 ( new_n4131 , n11192 , n22274 );
xnor g01783 ( new_n4132 , new_n4124 , new_n4131 );
nor  g01784 ( new_n4133 , new_n4130 , new_n4132 );
xnor g01785 ( new_n4134_1 , new_n4030 , n23065 );
not  g01786 ( new_n4135 , new_n4134_1 );
xnor g01787 ( new_n4136 , n9380 , n24129 );
nor  g01788 ( new_n4137 , new_n4135 , new_n4136 );
not  g01789 ( new_n4138 , new_n4130 );
xnor g01790 ( new_n4139 , new_n4138 , new_n4132 );
and  g01791 ( new_n4140 , new_n4137 , new_n4139 );
nor  g01792 ( new_n4141 , new_n4133 , new_n4140 );
xnor g01793 ( new_n4142 , new_n4128 , new_n4141 );
not  g01794 ( new_n4143 , n919 );
xnor g01795 ( new_n4144 , new_n4143 , n5330 );
nor  g01796 ( new_n4145 , n7657 , n25316 );
not  g01797 ( new_n4146_1 , n20385 );
or   g01798 ( new_n4147 , new_n4146_1 , new_n3982 );
xnor g01799 ( new_n4148 , new_n3978 , n25316 );
and  g01800 ( new_n4149 , new_n4147 , new_n4148 );
nor  g01801 ( new_n4150_1 , new_n4145 , new_n4149 );
xnor g01802 ( new_n4151_1 , new_n4144 , new_n4150_1 );
xnor g01803 ( new_n4152_1 , new_n4142 , new_n4151_1 );
xor  g01804 ( new_n4153_1 , new_n4137 , new_n4139 );
nor  g01805 ( new_n4154 , new_n4146_1 , new_n3982 );
xnor g01806 ( new_n4155 , new_n4154 , new_n4148 );
nor  g01807 ( new_n4156 , new_n4153_1 , new_n4155 );
xnor g01808 ( new_n4157 , n20385 , n25926 );
xnor g01809 ( new_n4158 , new_n4134_1 , new_n4136 );
nor  g01810 ( new_n4159 , new_n4157 , new_n4158 );
not  g01811 ( new_n4160 , new_n4155 );
xnor g01812 ( new_n4161 , new_n4153_1 , new_n4160 );
and  g01813 ( new_n4162 , new_n4159 , new_n4161 );
nor  g01814 ( new_n4163 , new_n4156 , new_n4162 );
xnor g01815 ( n248 , new_n4152_1 , new_n4163 );
not  g01816 ( new_n4165_1 , n6369 );
nor  g01817 ( new_n4166 , n6631 , n24732 );
not  g01818 ( new_n4167 , new_n4166 );
nor  g01819 ( new_n4168 , n14684 , new_n4167 );
not  g01820 ( new_n4169 , new_n4168 );
nor  g01821 ( new_n4170 , n17035 , new_n4169 );
xnor g01822 ( new_n4171 , n19905 , new_n4170 );
xnor g01823 ( new_n4172_1 , new_n4165_1 , new_n4171 );
xnor g01824 ( new_n4173_1 , n17035 , new_n4168 );
and  g01825 ( new_n4174 , n25797 , new_n4173_1 );
xnor g01826 ( new_n4175 , n25797 , new_n4173_1 );
xnor g01827 ( new_n4176_1 , n14684 , new_n4166 );
nor  g01828 ( new_n4177 , n15967 , new_n4176_1 );
not  g01829 ( new_n4178 , n15967 );
xnor g01830 ( new_n4179 , new_n4178 , new_n4176_1 );
not  g01831 ( new_n4180 , n6631 );
xnor g01832 ( new_n4181 , new_n4180 , n24732 );
nor  g01833 ( new_n4182 , n13319 , new_n4181 );
not  g01834 ( new_n4183 , n24732 );
or   g01835 ( new_n4184 , new_n4183 , new_n3756 );
not  g01836 ( new_n4185 , new_n4181 );
xnor g01837 ( new_n4186_1 , n13319 , new_n4185 );
and  g01838 ( new_n4187 , new_n4184 , new_n4186_1 );
or   g01839 ( new_n4188 , new_n4182 , new_n4187 );
and  g01840 ( new_n4189 , new_n4179 , new_n4188 );
nor  g01841 ( new_n4190 , new_n4177 , new_n4189 );
not  g01842 ( new_n4191 , new_n4190 );
nor  g01843 ( new_n4192 , new_n4175 , new_n4191 );
nor  g01844 ( new_n4193 , new_n4174 , new_n4192 );
xnor g01845 ( new_n4194 , new_n4172_1 , new_n4193 );
not  g01846 ( new_n4195 , new_n4194 );
nor  g01847 ( new_n4196 , n1152 , n14148 );
not  g01848 ( new_n4197 , new_n4196 );
nor  g01849 ( new_n4198 , n7149 , new_n4197 );
not  g01850 ( new_n4199 , new_n4198 );
nor  g01851 ( new_n4200 , n18558 , new_n4199 );
xnor g01852 ( new_n4201 , n3468 , new_n4200 );
not  g01853 ( new_n4202 , new_n4201 );
xnor g01854 ( new_n4203 , n19514 , new_n4202 );
xnor g01855 ( new_n4204_1 , n18558 , new_n4198 );
and  g01856 ( new_n4205_1 , n10053 , new_n4204_1 );
xnor g01857 ( new_n4206 , new_n2944_1 , new_n4204_1 );
xnor g01858 ( new_n4207 , n7149 , new_n4196 );
not  g01859 ( new_n4208 , new_n4207 );
nor  g01860 ( new_n4209 , new_n2947 , new_n4208 );
xnor g01861 ( new_n4210 , n8399 , new_n4208 );
xnor g01862 ( new_n4211 , n1152 , n14148 );
nor  g01863 ( new_n4212 , new_n3824 , new_n4211 );
nor  g01864 ( new_n4213 , new_n2698 , new_n2952 );
xnor g01865 ( new_n4214 , n9507 , new_n4211 );
and  g01866 ( new_n4215_1 , new_n4213 , new_n4214 );
or   g01867 ( new_n4216 , new_n4212 , new_n4215_1 );
and  g01868 ( new_n4217 , new_n4210 , new_n4216 );
or   g01869 ( new_n4218 , new_n4209 , new_n4217 );
and  g01870 ( new_n4219 , new_n4206 , new_n4218 );
nor  g01871 ( new_n4220 , new_n4205_1 , new_n4219 );
xnor g01872 ( new_n4221_1 , new_n4203 , new_n4220 );
not  g01873 ( new_n4222 , new_n4221_1 );
not  g01874 ( new_n4223 , n626 );
nor  g01875 ( new_n4224_1 , n8920 , n10057 );
not  g01876 ( new_n4225 , new_n4224_1 );
nor  g01877 ( new_n4226 , n26748 , new_n4225 );
not  g01878 ( new_n4227 , new_n4226 );
nor  g01879 ( new_n4228 , n21276 , new_n4227 );
xnor g01880 ( new_n4229 , n13668 , new_n4228 );
xnor g01881 ( new_n4230 , new_n4223 , new_n4229 );
xnor g01882 ( new_n4231_1 , n21276 , new_n4226 );
and  g01883 ( new_n4232 , n1204 , new_n4231_1 );
not  g01884 ( new_n4233 , n1204 );
xnor g01885 ( new_n4234 , new_n4233 , new_n4231_1 );
xnor g01886 ( new_n4235 , n26748 , new_n4224_1 );
and  g01887 ( new_n4236 , n19618 , new_n4235 );
not  g01888 ( new_n4237 , n19618 );
xnor g01889 ( new_n4238 , new_n4237 , new_n4235 );
xnor g01890 ( new_n4239 , n8920 , n10057 );
not  g01891 ( new_n4240 , new_n4239 );
nor  g01892 ( new_n4241 , n22043 , new_n4240 );
not  g01893 ( new_n4242 , n8920 );
or   g01894 ( new_n4243 , new_n4242 , new_n3875 );
xnor g01895 ( new_n4244 , n22043 , new_n4239 );
and  g01896 ( new_n4245 , new_n4243 , new_n4244 );
nor  g01897 ( new_n4246 , new_n4241 , new_n4245 );
and  g01898 ( new_n4247 , new_n4238 , new_n4246 );
or   g01899 ( new_n4248 , new_n4236 , new_n4247 );
and  g01900 ( new_n4249 , new_n4234 , new_n4248 );
nor  g01901 ( new_n4250 , new_n4232 , new_n4249 );
xnor g01902 ( new_n4251 , new_n4230 , new_n4250 );
xnor g01903 ( new_n4252 , new_n4222 , new_n4251 );
nor  g01904 ( new_n4253 , new_n4209 , new_n4217 );
xnor g01905 ( new_n4254 , new_n4206 , new_n4253 );
not  g01906 ( new_n4255 , new_n4254 );
nor  g01907 ( new_n4256_1 , new_n4236 , new_n4247 );
xnor g01908 ( new_n4257 , new_n4234 , new_n4256_1 );
not  g01909 ( new_n4258 , new_n4257 );
nor  g01910 ( new_n4259 , new_n4255 , new_n4258 );
xnor g01911 ( new_n4260 , new_n4255 , new_n4258 );
xnor g01912 ( new_n4261 , new_n4238 , new_n4246 );
xnor g01913 ( new_n4262 , new_n4213 , new_n4214 );
nor  g01914 ( new_n4263 , new_n4242 , new_n3875 );
xnor g01915 ( new_n4264 , new_n4263 , new_n4244 );
nor  g01916 ( new_n4265 , new_n4262 , new_n4264 );
xnor g01917 ( new_n4266_1 , n8920 , n12121 );
xnor g01918 ( new_n4267 , new_n2698 , n26979 );
not  g01919 ( new_n4268 , new_n4267 );
nor  g01920 ( new_n4269 , new_n4266_1 , new_n4268 );
not  g01921 ( new_n4270 , new_n4262 );
xnor g01922 ( new_n4271 , new_n4270 , new_n4264 );
and  g01923 ( new_n4272_1 , new_n4269 , new_n4271 );
nor  g01924 ( new_n4273 , new_n4265 , new_n4272_1 );
nor  g01925 ( new_n4274 , new_n4261 , new_n4273 );
nor  g01926 ( new_n4275 , new_n4212 , new_n4215_1 );
xnor g01927 ( new_n4276 , new_n4210 , new_n4275 );
not  g01928 ( new_n4277 , new_n4261 );
xnor g01929 ( new_n4278 , new_n4277 , new_n4273 );
and  g01930 ( new_n4279 , new_n4276 , new_n4278 );
nor  g01931 ( new_n4280 , new_n4274 , new_n4279 );
nor  g01932 ( new_n4281 , new_n4260 , new_n4280 );
or   g01933 ( new_n4282 , new_n4259 , new_n4281 );
xor  g01934 ( new_n4283 , new_n4252 , new_n4282 );
xnor g01935 ( new_n4284 , new_n4195 , new_n4283 );
xnor g01936 ( new_n4285 , new_n4175 , new_n4190 );
not  g01937 ( new_n4286 , new_n4285 );
xnor g01938 ( new_n4287 , new_n4260 , new_n4280 );
nor  g01939 ( new_n4288 , new_n4286 , new_n4287 );
xnor g01940 ( new_n4289 , new_n4285 , new_n4287 );
not  g01941 ( new_n4290 , new_n4276 );
xnor g01942 ( new_n4291 , new_n4290 , new_n4278 );
not  g01943 ( new_n4292 , new_n4291 );
xor  g01944 ( new_n4293 , new_n4179 , new_n4188 );
nor  g01945 ( new_n4294 , new_n4292 , new_n4293 );
xnor g01946 ( new_n4295 , new_n4291 , new_n4293 );
xnor g01947 ( new_n4296 , new_n4269 , new_n4271 );
not  g01948 ( new_n4297 , new_n4296 );
nor  g01949 ( new_n4298 , new_n4186_1 , new_n4297 );
xor  g01950 ( new_n4299 , new_n4184 , new_n4186_1 );
nor  g01951 ( new_n4300 , new_n4296 , new_n4299 );
xnor g01952 ( new_n4301 , n24732 , n25435 );
xnor g01953 ( new_n4302 , new_n4266_1 , new_n4267 );
not  g01954 ( new_n4303 , new_n4302 );
nor  g01955 ( new_n4304 , new_n4301 , new_n4303 );
nor  g01956 ( new_n4305 , new_n4300 , new_n4304 );
nor  g01957 ( new_n4306_1 , new_n4298 , new_n4305 );
and  g01958 ( new_n4307 , new_n4295 , new_n4306_1 );
or   g01959 ( new_n4308 , new_n4294 , new_n4307 );
and  g01960 ( new_n4309 , new_n4289 , new_n4308 );
nor  g01961 ( new_n4310 , new_n4288 , new_n4309 );
xnor g01962 ( n266 , new_n4284 , new_n4310 );
not  g01963 ( new_n4312 , n21839 );
nor  g01964 ( new_n4313 , new_n4312 , n22270 );
xnor g01965 ( new_n4314 , n21839 , n22270 );
not  g01966 ( new_n4315 , n27089 );
nor  g01967 ( new_n4316 , n8806 , new_n4315 );
xnor g01968 ( new_n4317 , n8806 , n27089 );
nor  g01969 ( new_n4318 , n2479 , new_n2929_1 );
xnor g01970 ( new_n4319_1 , n2479 , n11841 );
nor  g01971 ( new_n4320 , n9372 , new_n2933 );
xnor g01972 ( new_n4321 , n9372 , n10710 );
nor  g01973 ( new_n4322 , n6596 , new_n2937 );
xnor g01974 ( new_n4323 , n6596 , n20929 );
nor  g01975 ( new_n4324 , new_n2941 , n15289 );
xnor g01976 ( new_n4325_1 , n8006 , n15289 );
and  g01977 ( new_n4326_1 , new_n2692 , n25074 );
xnor g01978 ( new_n4327 , n6556 , n25074 );
not  g01979 ( new_n4328 , n16396 );
and  g01980 ( new_n4329 , new_n4328 , n22871 );
nor  g01981 ( new_n4330 , new_n4328 , n22871 );
not  g01982 ( new_n4331 , n9399 );
and  g01983 ( new_n4332 , new_n4331 , n14275 );
nor  g01984 ( new_n4333 , new_n4331 , n14275 );
nor  g01985 ( new_n4334 , n2088 , new_n2699 );
not  g01986 ( new_n4335 , new_n4334 );
nor  g01987 ( new_n4336 , new_n4333 , new_n4335 );
nor  g01988 ( new_n4337 , new_n4332 , new_n4336 );
nor  g01989 ( new_n4338 , new_n4330 , new_n4337 );
nor  g01990 ( new_n4339 , new_n4329 , new_n4338 );
and  g01991 ( new_n4340_1 , new_n4327 , new_n4339 );
or   g01992 ( new_n4341 , new_n4326_1 , new_n4340_1 );
and  g01993 ( new_n4342 , new_n4325_1 , new_n4341 );
or   g01994 ( new_n4343 , new_n4324 , new_n4342 );
and  g01995 ( new_n4344 , new_n4323 , new_n4343 );
or   g01996 ( new_n4345 , new_n4322 , new_n4344 );
and  g01997 ( new_n4346 , new_n4321 , new_n4345 );
or   g01998 ( new_n4347 , new_n4320 , new_n4346 );
and  g01999 ( new_n4348 , new_n4319_1 , new_n4347 );
or   g02000 ( new_n4349 , new_n4318 , new_n4348 );
and  g02001 ( new_n4350 , new_n4317 , new_n4349 );
or   g02002 ( new_n4351 , new_n4316 , new_n4350 );
and  g02003 ( new_n4352 , new_n4314 , new_n4351 );
nor  g02004 ( new_n4353 , new_n4313 , new_n4352 );
nor  g02005 ( new_n4354 , new_n4316 , new_n4350 );
xnor g02006 ( new_n4355 , new_n4314 , new_n4354 );
nor  g02007 ( new_n4356 , n23272 , new_n4355 );
not  g02008 ( new_n4357 , new_n4355 );
xnor g02009 ( new_n4358 , n23272 , new_n4357 );
xor  g02010 ( new_n4359 , new_n4317 , new_n4349 );
nor  g02011 ( new_n4360 , n11481 , new_n4359 );
not  g02012 ( new_n4361 , n11481 );
xnor g02013 ( new_n4362 , new_n4361 , new_n4359 );
xor  g02014 ( new_n4363 , new_n4319_1 , new_n4347 );
nor  g02015 ( new_n4364 , n16439 , new_n4363 );
not  g02016 ( new_n4365 , n16439 );
xnor g02017 ( new_n4366 , new_n4365 , new_n4363 );
xor  g02018 ( new_n4367 , new_n4321 , new_n4345 );
nor  g02019 ( new_n4368 , n15241 , new_n4367 );
not  g02020 ( new_n4369 , n15241 );
xnor g02021 ( new_n4370 , new_n4369 , new_n4367 );
xor  g02022 ( new_n4371 , new_n4323 , new_n4343 );
nor  g02023 ( new_n4372 , n7678 , new_n4371 );
not  g02024 ( new_n4373 , n7678 );
xnor g02025 ( new_n4374_1 , new_n4373 , new_n4371 );
xor  g02026 ( new_n4375 , new_n4325_1 , new_n4341 );
nor  g02027 ( new_n4376_1 , n3785 , new_n4375 );
not  g02028 ( new_n4377 , n3785 );
xnor g02029 ( new_n4378 , new_n4377 , new_n4375 );
xnor g02030 ( new_n4379 , new_n4327 , new_n4339 );
not  g02031 ( new_n4380 , new_n4379 );
nor  g02032 ( new_n4381 , n20250 , new_n4380 );
not  g02033 ( new_n4382 , n20250 );
xnor g02034 ( new_n4383 , new_n4382 , new_n4380 );
not  g02035 ( new_n4384 , n5822 );
xnor g02036 ( new_n4385 , n16396 , n22871 );
xnor g02037 ( new_n4386 , new_n4337 , new_n4385 );
nor  g02038 ( new_n4387 , new_n4384 , new_n4386 );
not  g02039 ( new_n4388 , new_n4386 );
or   g02040 ( new_n4389 , n5822 , new_n4388 );
xnor g02041 ( new_n4390 , n9399 , n14275 );
xnor g02042 ( new_n4391 , new_n4335 , new_n4390 );
not  g02043 ( new_n4392 , new_n4391 );
nor  g02044 ( new_n4393 , n26443 , new_n4392 );
not  g02045 ( new_n4394 , n1681 );
xnor g02046 ( new_n4395 , n2088 , n25023 );
or   g02047 ( new_n4396 , new_n4394 , new_n4395 );
xnor g02048 ( new_n4397 , n26443 , new_n4391 );
and  g02049 ( new_n4398 , new_n4396 , new_n4397 );
nor  g02050 ( new_n4399 , new_n4393 , new_n4398 );
and  g02051 ( new_n4400 , new_n4389 , new_n4399 );
nor  g02052 ( new_n4401_1 , new_n4387 , new_n4400 );
and  g02053 ( new_n4402 , new_n4383 , new_n4401_1 );
or   g02054 ( new_n4403 , new_n4381 , new_n4402 );
and  g02055 ( new_n4404 , new_n4378 , new_n4403 );
or   g02056 ( new_n4405 , new_n4376_1 , new_n4404 );
and  g02057 ( new_n4406 , new_n4374_1 , new_n4405 );
or   g02058 ( new_n4407 , new_n4372 , new_n4406 );
and  g02059 ( new_n4408 , new_n4370 , new_n4407 );
or   g02060 ( new_n4409_1 , new_n4368 , new_n4408 );
and  g02061 ( new_n4410 , new_n4366 , new_n4409_1 );
or   g02062 ( new_n4411 , new_n4364 , new_n4410 );
and  g02063 ( new_n4412 , new_n4362 , new_n4411 );
or   g02064 ( new_n4413 , new_n4360 , new_n4412 );
and  g02065 ( new_n4414 , new_n4358 , new_n4413 );
nor  g02066 ( new_n4415 , new_n4356 , new_n4414 );
and  g02067 ( new_n4416 , new_n4353 , new_n4415 );
not  g02068 ( new_n4417 , new_n4416 );
not  g02069 ( new_n4418 , new_n3934_1 );
nor  g02070 ( new_n4419 , n19477 , new_n4418 );
not  g02071 ( new_n4420 , new_n4419 );
nor  g02072 ( new_n4421 , n9318 , new_n4420 );
not  g02073 ( new_n4422 , new_n4421 );
nor  g02074 ( new_n4423 , n25168 , new_n4422 );
not  g02075 ( new_n4424_1 , new_n4423 );
nor  g02076 ( new_n4425 , n1999 , new_n4424_1 );
and  g02077 ( new_n4426_1 , new_n2554 , new_n4425 );
xnor g02078 ( new_n4427 , n9396 , new_n4425 );
nor  g02079 ( new_n4428 , n18880 , new_n4427 );
xnor g02080 ( new_n4429 , n1999 , new_n4423 );
nor  g02081 ( new_n4430 , n25475 , new_n4429 );
not  g02082 ( new_n4431 , n25475 );
xnor g02083 ( new_n4432_1 , new_n4431 , new_n4429 );
xnor g02084 ( new_n4433 , n25168 , new_n4421 );
nor  g02085 ( new_n4434 , n23849 , new_n4433 );
not  g02086 ( new_n4435 , n23849 );
xnor g02087 ( new_n4436 , new_n4435 , new_n4433 );
xnor g02088 ( new_n4437 , n9318 , new_n4419 );
nor  g02089 ( new_n4438 , n12446 , new_n4437 );
nor  g02090 ( new_n4439 , n11011 , new_n3935 );
nor  g02091 ( new_n4440 , new_n3936 , new_n3962_1 );
or   g02092 ( new_n4441_1 , new_n4439 , new_n4440 );
not  g02093 ( new_n4442 , n12446 );
xnor g02094 ( new_n4443 , new_n4442 , new_n4437 );
and  g02095 ( new_n4444 , new_n4441_1 , new_n4443 );
or   g02096 ( new_n4445 , new_n4438 , new_n4444 );
and  g02097 ( new_n4446 , new_n4436 , new_n4445 );
or   g02098 ( new_n4447 , new_n4434 , new_n4446 );
and  g02099 ( new_n4448 , new_n4432_1 , new_n4447 );
nor  g02100 ( new_n4449 , new_n4430 , new_n4448 );
and  g02101 ( new_n4450 , n18880 , new_n4427 );
nor  g02102 ( new_n4451_1 , new_n4449 , new_n4450 );
nor  g02103 ( new_n4452 , new_n4428 , new_n4451_1 );
nor  g02104 ( new_n4453 , new_n4426_1 , new_n4452 );
nor  g02105 ( new_n4454 , n22843 , n24032 );
not  g02106 ( new_n4455 , new_n4454 );
nor  g02107 ( new_n4456 , n6785 , new_n4455 );
not  g02108 ( new_n4457 , new_n4456 );
nor  g02109 ( new_n4458 , n24879 , new_n4457 );
not  g02110 ( new_n4459 , new_n4458 );
nor  g02111 ( new_n4460 , n268 , new_n4459 );
not  g02112 ( new_n4461 , new_n4460 );
nor  g02113 ( new_n4462 , n12587 , new_n4461 );
not  g02114 ( new_n4463 , new_n4462 );
nor  g02115 ( new_n4464 , n25381 , new_n4463 );
not  g02116 ( new_n4465 , new_n4464 );
nor  g02117 ( new_n4466 , n16376 , new_n4465 );
not  g02118 ( new_n4467 , new_n4466 );
nor  g02119 ( new_n4468 , n24196 , new_n4467 );
xnor g02120 ( new_n4469 , n18105 , new_n4468 );
not  g02121 ( new_n4470 , new_n4469 );
not  g02122 ( new_n4471 , n18880 );
xnor g02123 ( new_n4472 , new_n4471 , new_n4427 );
xnor g02124 ( new_n4473 , new_n4449 , new_n4472 );
nor  g02125 ( new_n4474 , new_n4470 , new_n4473 );
not  g02126 ( new_n4475 , new_n4468 );
nor  g02127 ( new_n4476_1 , n18105 , new_n4475 );
not  g02128 ( new_n4477 , new_n4473 );
xnor g02129 ( new_n4478_1 , new_n4470 , new_n4477 );
xnor g02130 ( new_n4479 , n24196 , new_n4466 );
nor  g02131 ( new_n4480 , new_n4434 , new_n4446 );
xnor g02132 ( new_n4481 , new_n4432_1 , new_n4480 );
not  g02133 ( new_n4482 , new_n4481 );
nor  g02134 ( new_n4483 , new_n4479 , new_n4482 );
xnor g02135 ( new_n4484 , new_n4479 , new_n4482 );
xnor g02136 ( new_n4485 , n16376 , new_n4464 );
nor  g02137 ( new_n4486 , new_n4438 , new_n4444 );
xnor g02138 ( new_n4487 , new_n4436 , new_n4486 );
not  g02139 ( new_n4488 , new_n4487 );
nor  g02140 ( new_n4489 , new_n4485 , new_n4488 );
xnor g02141 ( new_n4490 , new_n4485 , new_n4488 );
xnor g02142 ( new_n4491 , n25381 , new_n4462 );
xor  g02143 ( new_n4492 , new_n4441_1 , new_n4443 );
not  g02144 ( new_n4493 , new_n4492 );
nor  g02145 ( new_n4494 , new_n4491 , new_n4493 );
xnor g02146 ( new_n4495 , new_n4491 , new_n4493 );
xnor g02147 ( new_n4496 , n12587 , new_n4460 );
nor  g02148 ( new_n4497 , new_n3963 , new_n4496 );
xnor g02149 ( new_n4498 , new_n3963 , new_n4496 );
xnor g02150 ( new_n4499 , n268 , new_n4458 );
nor  g02151 ( new_n4500 , new_n3965 , new_n4499 );
xnor g02152 ( new_n4501 , n24879 , new_n4456 );
nor  g02153 ( new_n4502 , new_n3970 , new_n4501 );
xnor g02154 ( new_n4503 , new_n3968 , new_n4501 );
xnor g02155 ( new_n4504 , n6785 , new_n4454 );
and  g02156 ( new_n4505 , new_n3976 , new_n4504 );
xnor g02157 ( new_n4506 , new_n3974 , new_n4504 );
not  g02158 ( new_n4507 , n22843 );
xnor g02159 ( new_n4508 , new_n4507 , n24032 );
nor  g02160 ( new_n4509 , new_n3984_1 , new_n4508 );
or   g02161 ( new_n4510 , new_n4507 , new_n2551 );
xnor g02162 ( new_n4511 , new_n3980 , new_n4508 );
and  g02163 ( new_n4512 , new_n4510 , new_n4511 );
nor  g02164 ( new_n4513 , new_n4509 , new_n4512 );
and  g02165 ( new_n4514_1 , new_n4506 , new_n4513 );
nor  g02166 ( new_n4515 , new_n4505 , new_n4514_1 );
and  g02167 ( new_n4516 , new_n4503 , new_n4515 );
nor  g02168 ( new_n4517 , new_n4502 , new_n4516 );
xnor g02169 ( new_n4518 , new_n3965 , new_n4499 );
nor  g02170 ( new_n4519 , new_n4517 , new_n4518 );
nor  g02171 ( new_n4520 , new_n4500 , new_n4519 );
nor  g02172 ( new_n4521 , new_n4498 , new_n4520 );
nor  g02173 ( new_n4522 , new_n4497 , new_n4521 );
nor  g02174 ( new_n4523 , new_n4495 , new_n4522 );
nor  g02175 ( new_n4524 , new_n4494 , new_n4523 );
nor  g02176 ( new_n4525 , new_n4490 , new_n4524 );
nor  g02177 ( new_n4526 , new_n4489 , new_n4525 );
nor  g02178 ( new_n4527 , new_n4484 , new_n4526 );
nor  g02179 ( new_n4528 , new_n4483 , new_n4527 );
and  g02180 ( new_n4529_1 , new_n4478_1 , new_n4528 );
or   g02181 ( new_n4530 , new_n4476_1 , new_n4529_1 );
nor  g02182 ( new_n4531 , new_n4474 , new_n4530 );
not  g02183 ( new_n4532 , new_n4531 );
nor  g02184 ( new_n4533 , new_n4453 , new_n4532 );
xnor g02185 ( new_n4534 , new_n4417 , new_n4533 );
not  g02186 ( new_n4535 , new_n4415 );
xnor g02187 ( new_n4536 , new_n4353 , new_n4535 );
not  g02188 ( new_n4537 , new_n4536 );
not  g02189 ( new_n4538 , new_n4453 );
xnor g02190 ( new_n4539 , new_n4538 , new_n4532 );
and  g02191 ( new_n4540 , new_n4537 , new_n4539 );
xnor g02192 ( new_n4541 , new_n4537 , new_n4539 );
xnor g02193 ( new_n4542 , new_n4478_1 , new_n4528 );
nor  g02194 ( new_n4543 , new_n4360 , new_n4412 );
xnor g02195 ( new_n4544 , new_n4358 , new_n4543 );
and  g02196 ( new_n4545 , new_n4542 , new_n4544 );
xnor g02197 ( new_n4546 , new_n4542 , new_n4544 );
xnor g02198 ( new_n4547 , new_n4484 , new_n4526 );
xor  g02199 ( new_n4548 , new_n4362 , new_n4411 );
not  g02200 ( new_n4549 , new_n4548 );
nor  g02201 ( new_n4550 , new_n4547 , new_n4549 );
xnor g02202 ( new_n4551 , new_n4547 , new_n4549 );
xnor g02203 ( new_n4552_1 , new_n4490 , new_n4524 );
xor  g02204 ( new_n4553 , new_n4366 , new_n4409_1 );
not  g02205 ( new_n4554 , new_n4553 );
nor  g02206 ( new_n4555 , new_n4552_1 , new_n4554 );
xnor g02207 ( new_n4556 , new_n4552_1 , new_n4554 );
xnor g02208 ( new_n4557 , new_n4495 , new_n4522 );
xor  g02209 ( new_n4558 , new_n4370 , new_n4407 );
not  g02210 ( new_n4559 , new_n4558 );
nor  g02211 ( new_n4560 , new_n4557 , new_n4559 );
xnor g02212 ( new_n4561 , new_n4557 , new_n4559 );
xnor g02213 ( new_n4562 , new_n4498 , new_n4520 );
xor  g02214 ( new_n4563 , new_n4374_1 , new_n4405 );
not  g02215 ( new_n4564 , new_n4563 );
nor  g02216 ( new_n4565 , new_n4562 , new_n4564 );
xnor g02217 ( new_n4566 , new_n4562 , new_n4564 );
xor  g02218 ( new_n4567 , new_n4378 , new_n4403 );
not  g02219 ( new_n4568 , new_n4567 );
xnor g02220 ( new_n4569 , new_n4517 , new_n4518 );
nor  g02221 ( new_n4570 , new_n4568 , new_n4569 );
xnor g02222 ( new_n4571 , new_n4568 , new_n4569 );
xnor g02223 ( new_n4572 , new_n4503 , new_n4515 );
xnor g02224 ( new_n4573 , new_n4383 , new_n4401_1 );
nor  g02225 ( new_n4574 , new_n4572 , new_n4573 );
not  g02226 ( new_n4575 , new_n4573 );
xnor g02227 ( new_n4576 , new_n4572 , new_n4575 );
xnor g02228 ( new_n4577 , new_n4506 , new_n4513 );
xnor g02229 ( new_n4578 , new_n4384 , new_n4388 );
xnor g02230 ( new_n4579 , new_n4399 , new_n4578 );
nor  g02231 ( new_n4580 , new_n4577 , new_n4579 );
xor  g02232 ( new_n4581 , new_n4396 , new_n4397 );
xor  g02233 ( new_n4582 , new_n4510 , new_n4511 );
and  g02234 ( new_n4583 , new_n4581 , new_n4582 );
xnor g02235 ( new_n4584 , new_n4507 , new_n2551 );
xnor g02236 ( new_n4585 , n1681 , new_n4395 );
not  g02237 ( new_n4586 , new_n4585 );
nor  g02238 ( new_n4587 , new_n4584 , new_n4586 );
xnor g02239 ( new_n4588_1 , new_n4581 , new_n4582 );
nor  g02240 ( new_n4589 , new_n4587 , new_n4588_1 );
nor  g02241 ( new_n4590_1 , new_n4583 , new_n4589 );
not  g02242 ( new_n4591 , new_n4579 );
xnor g02243 ( new_n4592 , new_n4577 , new_n4591 );
and  g02244 ( new_n4593 , new_n4590_1 , new_n4592 );
nor  g02245 ( new_n4594 , new_n4580 , new_n4593 );
and  g02246 ( new_n4595_1 , new_n4576 , new_n4594 );
nor  g02247 ( new_n4596 , new_n4574 , new_n4595_1 );
nor  g02248 ( new_n4597 , new_n4571 , new_n4596 );
nor  g02249 ( new_n4598 , new_n4570 , new_n4597 );
nor  g02250 ( new_n4599 , new_n4566 , new_n4598 );
nor  g02251 ( new_n4600 , new_n4565 , new_n4599 );
nor  g02252 ( new_n4601 , new_n4561 , new_n4600 );
nor  g02253 ( new_n4602 , new_n4560 , new_n4601 );
nor  g02254 ( new_n4603 , new_n4556 , new_n4602 );
nor  g02255 ( new_n4604 , new_n4555 , new_n4603 );
nor  g02256 ( new_n4605 , new_n4551 , new_n4604 );
nor  g02257 ( new_n4606 , new_n4550 , new_n4605 );
nor  g02258 ( new_n4607 , new_n4546 , new_n4606 );
nor  g02259 ( new_n4608 , new_n4545 , new_n4607 );
nor  g02260 ( new_n4609 , new_n4541 , new_n4608 );
nor  g02261 ( new_n4610 , new_n4540 , new_n4609 );
not  g02262 ( new_n4611 , new_n4610 );
xnor g02263 ( n298 , new_n4534 , new_n4611 );
xnor g02264 ( new_n4613 , n20604 , n21735 );
not  g02265 ( new_n4614 , n16158 );
and  g02266 ( new_n4615 , new_n4614 , n24085 );
xnor g02267 ( new_n4616 , n16158 , n24085 );
not  g02268 ( new_n4617 , n5752 );
and  g02269 ( new_n4618 , new_n4617 , n14071 );
xnor g02270 ( new_n4619 , n5752 , n14071 );
not  g02271 ( new_n4620 , n18171 );
nor  g02272 ( new_n4621 , n1738 , new_n4620 );
and  g02273 ( new_n4622 , n1738 , new_n4620 );
not  g02274 ( new_n4623 , n25073 );
nor  g02275 ( new_n4624_1 , n12152 , new_n4623 );
nand g02276 ( new_n4625 , n12152 , new_n4623 );
not  g02277 ( new_n4626 , n22309 );
nor  g02278 ( new_n4627 , n19107 , new_n4626 );
and  g02279 ( new_n4628 , new_n4625 , new_n4627 );
nor  g02280 ( new_n4629 , new_n4624_1 , new_n4628 );
nor  g02281 ( new_n4630 , new_n4622 , new_n4629 );
nor  g02282 ( new_n4631 , new_n4621 , new_n4630 );
and  g02283 ( new_n4632 , new_n4619 , new_n4631 );
or   g02284 ( new_n4633 , new_n4618 , new_n4632 );
and  g02285 ( new_n4634 , new_n4616 , new_n4633 );
or   g02286 ( new_n4635 , new_n4615 , new_n4634 );
xor  g02287 ( new_n4636 , new_n4613 , new_n4635 );
xnor g02288 ( new_n4637 , n1525 , n4119 );
not  g02289 ( new_n4638 , n16988 );
nor  g02290 ( new_n4639 , n14510 , new_n4638 );
xnor g02291 ( new_n4640 , n14510 , n16988 );
not  g02292 ( new_n4641 , n21779 );
nor  g02293 ( new_n4642 , n13263 , new_n4641 );
xnor g02294 ( new_n4643 , n13263 , n21779 );
nor  g02295 ( new_n4644 , n5376 , new_n3446 );
not  g02296 ( new_n4645 , n5376 );
nor  g02297 ( new_n4646_1 , new_n4645 , n20455 );
nor  g02298 ( new_n4647 , new_n3448 , n5128 );
not  g02299 ( new_n4648 , n5128 );
nor  g02300 ( new_n4649 , n1639 , new_n4648 );
nor  g02301 ( new_n4650 , new_n3451_1 , n23120 );
not  g02302 ( new_n4651 , new_n4650 );
nor  g02303 ( new_n4652 , new_n4649 , new_n4651 );
nor  g02304 ( new_n4653 , new_n4647 , new_n4652 );
nor  g02305 ( new_n4654 , new_n4646_1 , new_n4653 );
nor  g02306 ( new_n4655 , new_n4644 , new_n4654 );
and  g02307 ( new_n4656 , new_n4643 , new_n4655 );
or   g02308 ( new_n4657 , new_n4642 , new_n4656 );
and  g02309 ( new_n4658 , new_n4640 , new_n4657 );
or   g02310 ( new_n4659 , new_n4639 , new_n4658 );
xor  g02311 ( new_n4660 , new_n4637 , new_n4659 );
xnor g02312 ( new_n4661 , n4272 , n12626 );
not  g02313 ( new_n4662 , n24319 );
nor  g02314 ( new_n4663 , n6971 , new_n4662 );
xnor g02315 ( new_n4664 , n6971 , n24319 );
not  g02316 ( new_n4665_1 , n7460 );
nor  g02317 ( new_n4666 , new_n4665_1 , n22068 );
xnor g02318 ( new_n4667 , n7460 , n22068 );
not  g02319 ( new_n4668 , n196 );
and  g02320 ( new_n4669 , new_n4668 , n9460 );
nor  g02321 ( new_n4670 , new_n4668 , n9460 );
not  g02322 ( new_n4671 , n11749 );
and  g02323 ( new_n4672 , new_n4671 , n14954 );
nor  g02324 ( new_n4673 , new_n4671 , n14954 );
not  g02325 ( new_n4674_1 , n23831 );
nor  g02326 ( new_n4675 , n13424 , new_n4674_1 );
not  g02327 ( new_n4676 , new_n4675 );
nor  g02328 ( new_n4677 , new_n4673 , new_n4676 );
nor  g02329 ( new_n4678 , new_n4672 , new_n4677 );
nor  g02330 ( new_n4679 , new_n4670 , new_n4678 );
nor  g02331 ( new_n4680 , new_n4669 , new_n4679 );
and  g02332 ( new_n4681 , new_n4667 , new_n4680 );
or   g02333 ( new_n4682 , new_n4666 , new_n4681 );
and  g02334 ( new_n4683 , new_n4664 , new_n4682 );
or   g02335 ( new_n4684 , new_n4663 , new_n4683 );
xor  g02336 ( new_n4685 , new_n4661 , new_n4684 );
xnor g02337 ( new_n4686 , new_n4660 , new_n4685 );
xor  g02338 ( new_n4687 , new_n4640 , new_n4657 );
xor  g02339 ( new_n4688 , new_n4664 , new_n4682 );
and  g02340 ( new_n4689 , new_n4687 , new_n4688 );
xor  g02341 ( new_n4690 , new_n4687 , new_n4688 );
xnor g02342 ( new_n4691 , new_n4643 , new_n4655 );
not  g02343 ( new_n4692 , new_n4691 );
xnor g02344 ( new_n4693_1 , new_n4667 , new_n4680 );
not  g02345 ( new_n4694 , new_n4693_1 );
nor  g02346 ( new_n4695 , new_n4692 , new_n4694 );
xnor g02347 ( new_n4696 , new_n4692 , new_n4694 );
xnor g02348 ( new_n4697 , n5376 , n20455 );
xnor g02349 ( new_n4698 , new_n4653 , new_n4697 );
not  g02350 ( new_n4699 , new_n4698 );
xnor g02351 ( new_n4700 , n196 , n9460 );
xnor g02352 ( new_n4701 , new_n4678 , new_n4700 );
not  g02353 ( new_n4702 , new_n4701 );
nor  g02354 ( new_n4703 , new_n4699 , new_n4702 );
xnor g02355 ( new_n4704 , new_n4699 , new_n4701 );
xnor g02356 ( new_n4705 , n1639 , n5128 );
xnor g02357 ( new_n4706 , new_n4651 , new_n4705 );
xnor g02358 ( new_n4707 , n11749 , n14954 );
xnor g02359 ( new_n4708 , new_n4676 , new_n4707 );
nor  g02360 ( new_n4709 , new_n4706 , new_n4708 );
xnor g02361 ( new_n4710 , n16968 , n23120 );
xnor g02362 ( new_n4711 , n13424 , n23831 );
nor  g02363 ( new_n4712 , new_n4710 , new_n4711 );
not  g02364 ( new_n4713 , new_n4706 );
xnor g02365 ( new_n4714 , new_n4713 , new_n4708 );
and  g02366 ( new_n4715 , new_n4712 , new_n4714 );
nor  g02367 ( new_n4716 , new_n4709 , new_n4715 );
and  g02368 ( new_n4717 , new_n4704 , new_n4716 );
nor  g02369 ( new_n4718 , new_n4703 , new_n4717 );
nor  g02370 ( new_n4719 , new_n4696 , new_n4718 );
nor  g02371 ( new_n4720 , new_n4695 , new_n4719 );
and  g02372 ( new_n4721 , new_n4690 , new_n4720 );
nor  g02373 ( new_n4722_1 , new_n4689 , new_n4721 );
xnor g02374 ( new_n4723 , new_n4686 , new_n4722_1 );
xnor g02375 ( new_n4724 , new_n4636 , new_n4723 );
xor  g02376 ( new_n4725 , new_n4616 , new_n4633 );
xor  g02377 ( new_n4726 , new_n4690 , new_n4720 );
nor  g02378 ( new_n4727 , new_n4725 , new_n4726 );
xnor g02379 ( new_n4728 , new_n4725 , new_n4726 );
xnor g02380 ( new_n4729 , new_n4696 , new_n4718 );
not  g02381 ( new_n4730 , new_n4729 );
xnor g02382 ( new_n4731_1 , new_n4619 , new_n4631 );
and  g02383 ( new_n4732 , new_n4730 , new_n4731_1 );
xnor g02384 ( new_n4733 , new_n4704 , new_n4716 );
not  g02385 ( new_n4734 , new_n4733 );
xnor g02386 ( new_n4735 , n1738 , n18171 );
xnor g02387 ( new_n4736 , new_n4629 , new_n4735 );
and  g02388 ( new_n4737 , new_n4734 , new_n4736 );
xnor g02389 ( new_n4738 , new_n4734 , new_n4736 );
xnor g02390 ( new_n4739 , n19107 , n22309 );
xnor g02391 ( new_n4740 , new_n4710 , new_n4711 );
nor  g02392 ( new_n4741 , new_n4739 , new_n4740 );
xnor g02393 ( new_n4742 , n12152 , n25073 );
xnor g02394 ( new_n4743 , new_n4627 , new_n4742 );
nor  g02395 ( new_n4744 , new_n4741 , new_n4743 );
xnor g02396 ( new_n4745_1 , new_n4712 , new_n4714 );
not  g02397 ( new_n4746 , new_n4745_1 );
xnor g02398 ( new_n4747_1 , new_n4741 , new_n4743 );
nor  g02399 ( new_n4748 , new_n4746 , new_n4747_1 );
nor  g02400 ( new_n4749 , new_n4744 , new_n4748 );
nor  g02401 ( new_n4750 , new_n4738 , new_n4749 );
nor  g02402 ( new_n4751 , new_n4737 , new_n4750 );
xnor g02403 ( new_n4752 , new_n4730 , new_n4731_1 );
nor  g02404 ( new_n4753 , new_n4751 , new_n4752 );
nor  g02405 ( new_n4754 , new_n4732 , new_n4753 );
nor  g02406 ( new_n4755 , new_n4728 , new_n4754 );
nor  g02407 ( new_n4756 , new_n4727 , new_n4755 );
xor  g02408 ( n317 , new_n4724 , new_n4756 );
nor  g02409 ( new_n4758 , n3506 , n9934 );
xnor g02410 ( new_n4759 , n3506 , n9934 );
nor  g02411 ( new_n4760 , n14899 , n18496 );
xnor g02412 ( new_n4761 , n14899 , n18496 );
nor  g02413 ( new_n4762 , n18444 , n26224 );
xnor g02414 ( new_n4763 , n18444 , n26224 );
nor  g02415 ( new_n4764 , n19327 , n24638 );
xnor g02416 ( new_n4765 , n19327 , n24638 );
nor  g02417 ( new_n4766_1 , n21674 , n22597 );
xnor g02418 ( new_n4767 , n21674 , n22597 );
nor  g02419 ( new_n4768 , n17251 , n26107 );
xnor g02420 ( new_n4769 , n17251 , n26107 );
nor  g02421 ( new_n4770_1 , n342 , n14790 );
xnor g02422 ( new_n4771 , n342 , n14790 );
nor  g02423 ( new_n4772 , n10096 , n26553 );
xnor g02424 ( new_n4773 , new_n3555_1 , n26553 );
nor  g02425 ( new_n4774 , n4964 , n16994 );
nor  g02426 ( new_n4775 , new_n3755_1 , new_n3562 );
not  g02427 ( new_n4776 , n4964 );
xnor g02428 ( new_n4777_1 , new_n4776 , n16994 );
not  g02429 ( new_n4778 , new_n4777_1 );
nor  g02430 ( new_n4779 , new_n4775 , new_n4778 );
or   g02431 ( new_n4780 , new_n4774 , new_n4779 );
and  g02432 ( new_n4781 , new_n4773 , new_n4780 );
nor  g02433 ( new_n4782 , new_n4772 , new_n4781 );
nor  g02434 ( new_n4783 , new_n4771 , new_n4782 );
nor  g02435 ( new_n4784 , new_n4770_1 , new_n4783 );
nor  g02436 ( new_n4785_1 , new_n4769 , new_n4784 );
nor  g02437 ( new_n4786 , new_n4768 , new_n4785_1 );
nor  g02438 ( new_n4787 , new_n4767 , new_n4786 );
nor  g02439 ( new_n4788 , new_n4766_1 , new_n4787 );
nor  g02440 ( new_n4789 , new_n4765 , new_n4788 );
nor  g02441 ( new_n4790 , new_n4764 , new_n4789 );
nor  g02442 ( new_n4791 , new_n4763 , new_n4790 );
nor  g02443 ( new_n4792 , new_n4762 , new_n4791 );
nor  g02444 ( new_n4793 , new_n4761 , new_n4792 );
nor  g02445 ( new_n4794 , new_n4760 , new_n4793 );
nor  g02446 ( new_n4795 , new_n4759 , new_n4794 );
nor  g02447 ( new_n4796 , new_n4758 , new_n4795 );
not  g02448 ( new_n4797 , n9259 );
not  g02449 ( new_n4798 , n2979 );
xnor g02450 ( new_n4799 , new_n4798 , n9554 );
nor  g02451 ( new_n4800 , n647 , n26408 );
not  g02452 ( new_n4801 , n647 );
xnor g02453 ( new_n4802 , new_n4801 , n26408 );
nor  g02454 ( new_n4803 , n18227 , n20409 );
not  g02455 ( new_n4804_1 , n18227 );
xnor g02456 ( new_n4805 , new_n4804_1 , n20409 );
nor  g02457 ( new_n4806 , n7377 , n25749 );
not  g02458 ( new_n4807 , n7377 );
xnor g02459 ( new_n4808 , new_n4807 , n25749 );
nor  g02460 ( new_n4809 , n3161 , n11630 );
xnor g02461 ( new_n4810_1 , new_n3774 , n11630 );
nor  g02462 ( new_n4811 , n9003 , n13453 );
xnor g02463 ( new_n4812_1 , new_n3778 , n13453 );
nor  g02464 ( new_n4813 , n4957 , n7421 );
xnor g02465 ( new_n4814_1 , new_n3784 , n7421 );
nor  g02466 ( new_n4815 , n7524 , n19680 );
xnor g02467 ( new_n4816 , new_n3788 , n19680 );
nor  g02468 ( new_n4817 , n2809 , n15743 );
not  g02469 ( new_n4818 , n15508 );
nor  g02470 ( new_n4819 , new_n4818 , new_n3798 );
xnor g02471 ( new_n4820 , n2809 , n15743 );
nor  g02472 ( new_n4821 , new_n4819 , new_n4820 );
or   g02473 ( new_n4822 , new_n4817 , new_n4821 );
and  g02474 ( new_n4823 , new_n4816 , new_n4822 );
or   g02475 ( new_n4824 , new_n4815 , new_n4823 );
and  g02476 ( new_n4825 , new_n4814_1 , new_n4824 );
or   g02477 ( new_n4826 , new_n4813 , new_n4825 );
and  g02478 ( new_n4827 , new_n4812_1 , new_n4826 );
or   g02479 ( new_n4828 , new_n4811 , new_n4827 );
and  g02480 ( new_n4829 , new_n4810_1 , new_n4828 );
or   g02481 ( new_n4830 , new_n4809 , new_n4829 );
and  g02482 ( new_n4831 , new_n4808 , new_n4830 );
or   g02483 ( new_n4832 , new_n4806 , new_n4831 );
and  g02484 ( new_n4833 , new_n4805 , new_n4832 );
or   g02485 ( new_n4834 , new_n4803 , new_n4833 );
and  g02486 ( new_n4835 , new_n4802 , new_n4834 );
nor  g02487 ( new_n4836 , new_n4800 , new_n4835 );
xnor g02488 ( new_n4837 , new_n4799 , new_n4836 );
nor  g02489 ( new_n4838 , new_n4797 , new_n4837 );
not  g02490 ( new_n4839 , new_n4837 );
xnor g02491 ( new_n4840 , new_n4797 , new_n4839 );
xor  g02492 ( new_n4841 , new_n4802 , new_n4834 );
nor  g02493 ( new_n4842 , new_n3583 , new_n4841 );
xnor g02494 ( new_n4843 , new_n3583 , new_n4841 );
not  g02495 ( new_n4844 , n20213 );
xor  g02496 ( new_n4845 , new_n4805 , new_n4832 );
nor  g02497 ( new_n4846 , new_n4844 , new_n4845 );
xnor g02498 ( new_n4847 , new_n4844 , new_n4845 );
not  g02499 ( new_n4848 , n13912 );
nor  g02500 ( new_n4849 , new_n4809 , new_n4829 );
xnor g02501 ( new_n4850_1 , new_n4808 , new_n4849 );
nor  g02502 ( new_n4851 , new_n4848 , new_n4850_1 );
xnor g02503 ( new_n4852 , new_n4848 , new_n4850_1 );
not  g02504 ( new_n4853 , n7670 );
xor  g02505 ( new_n4854 , new_n4810_1 , new_n4828 );
nor  g02506 ( new_n4855 , new_n4853 , new_n4854 );
xnor g02507 ( new_n4856 , new_n4853 , new_n4854 );
not  g02508 ( new_n4857 , n9598 );
nor  g02509 ( new_n4858_1 , new_n4813 , new_n4825 );
xnor g02510 ( new_n4859 , new_n4812_1 , new_n4858_1 );
nor  g02511 ( new_n4860 , new_n4857 , new_n4859 );
not  g02512 ( new_n4861 , new_n4859 );
xnor g02513 ( new_n4862 , n9598 , new_n4861 );
not  g02514 ( new_n4863 , n22290 );
xor  g02515 ( new_n4864 , new_n4814_1 , new_n4824 );
nor  g02516 ( new_n4865 , new_n4863 , new_n4864 );
xnor g02517 ( new_n4866 , new_n4863 , new_n4864 );
not  g02518 ( new_n4867 , n11273 );
nor  g02519 ( new_n4868 , new_n4817 , new_n4821 );
xnor g02520 ( new_n4869 , new_n4816 , new_n4868 );
nor  g02521 ( new_n4870 , new_n4867 , new_n4869 );
xor  g02522 ( new_n4871 , new_n4819 , new_n4820 );
not  g02523 ( new_n4872 , new_n4871 );
nor  g02524 ( new_n4873 , n25565 , new_n4872 );
xnor g02525 ( new_n4874 , n15508 , n20658 );
nor  g02526 ( new_n4875 , new_n3635 , new_n4874 );
xnor g02527 ( new_n4876 , n25565 , new_n4872 );
nor  g02528 ( new_n4877 , new_n4875 , new_n4876 );
nor  g02529 ( new_n4878 , new_n4873 , new_n4877 );
not  g02530 ( new_n4879 , new_n4878 );
not  g02531 ( new_n4880 , new_n4869 );
xnor g02532 ( new_n4881 , n11273 , new_n4880 );
nor  g02533 ( new_n4882 , new_n4879 , new_n4881 );
nor  g02534 ( new_n4883 , new_n4870 , new_n4882 );
nor  g02535 ( new_n4884 , new_n4866 , new_n4883 );
nor  g02536 ( new_n4885 , new_n4865 , new_n4884 );
nor  g02537 ( new_n4886 , new_n4862 , new_n4885 );
nor  g02538 ( new_n4887 , new_n4860 , new_n4886 );
nor  g02539 ( new_n4888 , new_n4856 , new_n4887 );
nor  g02540 ( new_n4889 , new_n4855 , new_n4888 );
nor  g02541 ( new_n4890 , new_n4852 , new_n4889 );
nor  g02542 ( new_n4891_1 , new_n4851 , new_n4890 );
nor  g02543 ( new_n4892 , new_n4847 , new_n4891_1 );
nor  g02544 ( new_n4893 , new_n4846 , new_n4892 );
nor  g02545 ( new_n4894 , new_n4843 , new_n4893 );
or   g02546 ( new_n4895 , new_n4842 , new_n4894 );
and  g02547 ( new_n4896 , new_n4840 , new_n4895 );
nor  g02548 ( new_n4897 , new_n4838 , new_n4896 );
nor  g02549 ( new_n4898 , n2979 , n9554 );
or   g02550 ( new_n4899 , new_n4800 , new_n4835 );
and  g02551 ( new_n4900 , new_n4799 , new_n4899 );
nor  g02552 ( new_n4901 , new_n4898 , new_n4900 );
xnor g02553 ( new_n4902 , new_n4897 , new_n4901 );
nor  g02554 ( new_n4903 , new_n4842 , new_n4894 );
xnor g02555 ( new_n4904 , new_n4840 , new_n4903 );
not  g02556 ( new_n4905 , new_n4904 );
nor  g02557 ( new_n4906 , n3740 , new_n4905 );
not  g02558 ( new_n4907 , n3740 );
xnor g02559 ( new_n4908 , new_n4907 , new_n4905 );
not  g02560 ( new_n4909 , n2858 );
xor  g02561 ( new_n4910 , new_n4843 , new_n4893 );
nor  g02562 ( new_n4911 , new_n4909 , new_n4910 );
xnor g02563 ( new_n4912 , new_n4909 , new_n4910 );
not  g02564 ( new_n4913_1 , n2659 );
xor  g02565 ( new_n4914 , new_n4847 , new_n4891_1 );
nor  g02566 ( new_n4915 , new_n4913_1 , new_n4914 );
xnor g02567 ( new_n4916 , new_n4913_1 , new_n4914 );
not  g02568 ( new_n4917 , n24327 );
xor  g02569 ( new_n4918 , new_n4852 , new_n4889 );
nor  g02570 ( new_n4919 , new_n4917 , new_n4918 );
not  g02571 ( new_n4920 , new_n4918 );
xnor g02572 ( new_n4921 , n24327 , new_n4920 );
not  g02573 ( new_n4922 , n22198 );
xor  g02574 ( new_n4923 , new_n4856 , new_n4887 );
nor  g02575 ( new_n4924 , new_n4922 , new_n4923 );
not  g02576 ( new_n4925_1 , new_n4923 );
xnor g02577 ( new_n4926 , n22198 , new_n4925_1 );
not  g02578 ( new_n4927 , n20826 );
xor  g02579 ( new_n4928 , new_n4862 , new_n4885 );
nor  g02580 ( new_n4929 , new_n4927 , new_n4928 );
not  g02581 ( new_n4930 , new_n4928 );
xnor g02582 ( new_n4931 , n20826 , new_n4930 );
not  g02583 ( new_n4932 , n7305 );
xor  g02584 ( new_n4933 , new_n4866 , new_n4883 );
nor  g02585 ( new_n4934 , new_n4932 , new_n4933 );
xnor g02586 ( new_n4935 , new_n4878 , new_n4881 );
not  g02587 ( new_n4936 , new_n4935 );
nor  g02588 ( new_n4937 , n25872 , new_n4936 );
xnor g02589 ( new_n4938 , n25872 , new_n4935 );
not  g02590 ( new_n4939_1 , n20259 );
xnor g02591 ( new_n4940 , new_n4875 , new_n4876 );
nor  g02592 ( new_n4941 , new_n4939_1 , new_n4940 );
xnor g02593 ( new_n4942 , n21993 , new_n4874 );
not  g02594 ( new_n4943 , new_n4942 );
nor  g02595 ( new_n4944 , n3925 , new_n4943 );
xnor g02596 ( new_n4945 , new_n4939_1 , new_n4940 );
nor  g02597 ( new_n4946 , new_n4944 , new_n4945 );
nor  g02598 ( new_n4947_1 , new_n4941 , new_n4946 );
and  g02599 ( new_n4948 , new_n4938 , new_n4947_1 );
nor  g02600 ( new_n4949 , new_n4937 , new_n4948 );
not  g02601 ( new_n4950 , new_n4933 );
xnor g02602 ( new_n4951 , new_n4932 , new_n4950 );
and  g02603 ( new_n4952_1 , new_n4949 , new_n4951 );
nor  g02604 ( new_n4953 , new_n4934 , new_n4952_1 );
nor  g02605 ( new_n4954 , new_n4931 , new_n4953 );
nor  g02606 ( new_n4955 , new_n4929 , new_n4954 );
nor  g02607 ( new_n4956 , new_n4926 , new_n4955 );
nor  g02608 ( new_n4957_1 , new_n4924 , new_n4956 );
nor  g02609 ( new_n4958 , new_n4921 , new_n4957_1 );
nor  g02610 ( new_n4959 , new_n4919 , new_n4958 );
nor  g02611 ( new_n4960 , new_n4916 , new_n4959 );
nor  g02612 ( new_n4961 , new_n4915 , new_n4960 );
nor  g02613 ( new_n4962 , new_n4912 , new_n4961 );
nor  g02614 ( new_n4963 , new_n4911 , new_n4962 );
and  g02615 ( new_n4964_1 , new_n4908 , new_n4963 );
nor  g02616 ( new_n4965 , new_n4906 , new_n4964_1 );
xnor g02617 ( new_n4966_1 , new_n4902 , new_n4965 );
xor  g02618 ( new_n4967_1 , new_n4796 , new_n4966_1 );
xnor g02619 ( new_n4968 , new_n4759 , new_n4794 );
xnor g02620 ( new_n4969 , new_n4908 , new_n4963 );
nor  g02621 ( new_n4970 , new_n4968 , new_n4969 );
xnor g02622 ( new_n4971 , new_n4968 , new_n4969 );
xnor g02623 ( new_n4972_1 , new_n4761 , new_n4792 );
xor  g02624 ( new_n4973 , new_n4912 , new_n4961 );
nor  g02625 ( new_n4974 , new_n4972_1 , new_n4973 );
xnor g02626 ( new_n4975 , new_n4972_1 , new_n4973 );
xnor g02627 ( new_n4976 , new_n4763 , new_n4790 );
xor  g02628 ( new_n4977 , new_n4916 , new_n4959 );
nor  g02629 ( new_n4978 , new_n4976 , new_n4977 );
xnor g02630 ( new_n4979 , new_n4976 , new_n4977 );
xnor g02631 ( new_n4980 , new_n4765 , new_n4788 );
xor  g02632 ( new_n4981 , new_n4921 , new_n4957_1 );
nor  g02633 ( new_n4982 , new_n4980 , new_n4981 );
xnor g02634 ( new_n4983 , new_n4980 , new_n4981 );
xnor g02635 ( new_n4984 , new_n4767 , new_n4786 );
xor  g02636 ( new_n4985 , new_n4926 , new_n4955 );
nor  g02637 ( new_n4986 , new_n4984 , new_n4985 );
xnor g02638 ( new_n4987 , new_n4984 , new_n4985 );
xnor g02639 ( new_n4988 , new_n4769 , new_n4784 );
xor  g02640 ( new_n4989 , new_n4931 , new_n4953 );
nor  g02641 ( new_n4990 , new_n4988 , new_n4989 );
xnor g02642 ( new_n4991 , new_n4988 , new_n4989 );
xnor g02643 ( new_n4992 , new_n4771 , new_n4782 );
xor  g02644 ( new_n4993 , new_n4949 , new_n4951 );
nor  g02645 ( new_n4994 , new_n4992 , new_n4993 );
xnor g02646 ( new_n4995 , new_n4992 , new_n4993 );
xnor g02647 ( new_n4996 , new_n4938 , new_n4947_1 );
nor  g02648 ( new_n4997 , new_n4774 , new_n4779 );
xnor g02649 ( new_n4998 , new_n4773 , new_n4997 );
not  g02650 ( new_n4999 , new_n4998 );
nor  g02651 ( new_n5000 , new_n4996 , new_n4999 );
xnor g02652 ( new_n5001 , new_n4996 , new_n4998 );
not  g02653 ( new_n5002 , n3925 );
xnor g02654 ( new_n5003 , new_n5002 , new_n4943 );
xnor g02655 ( new_n5004 , n7876 , n9246 );
nor  g02656 ( new_n5005 , new_n5003 , new_n5004 );
and  g02657 ( new_n5006 , new_n4777_1 , new_n5005 );
xor  g02658 ( new_n5007 , new_n4944 , new_n4945 );
xnor g02659 ( new_n5008 , new_n4775 , new_n4778 );
nor  g02660 ( new_n5009 , new_n5005 , new_n5008 );
nor  g02661 ( new_n5010 , new_n5006 , new_n5009 );
and  g02662 ( new_n5011_1 , new_n5007 , new_n5010 );
nor  g02663 ( new_n5012 , new_n5006 , new_n5011_1 );
and  g02664 ( new_n5013 , new_n5001 , new_n5012 );
nor  g02665 ( new_n5014 , new_n5000 , new_n5013 );
nor  g02666 ( new_n5015 , new_n4995 , new_n5014 );
nor  g02667 ( new_n5016 , new_n4994 , new_n5015 );
nor  g02668 ( new_n5017 , new_n4991 , new_n5016 );
nor  g02669 ( new_n5018 , new_n4990 , new_n5017 );
nor  g02670 ( new_n5019 , new_n4987 , new_n5018 );
nor  g02671 ( new_n5020_1 , new_n4986 , new_n5019 );
nor  g02672 ( new_n5021 , new_n4983 , new_n5020_1 );
nor  g02673 ( new_n5022 , new_n4982 , new_n5021 );
nor  g02674 ( new_n5023 , new_n4979 , new_n5022 );
nor  g02675 ( new_n5024_1 , new_n4978 , new_n5023 );
nor  g02676 ( new_n5025_1 , new_n4975 , new_n5024_1 );
nor  g02677 ( new_n5026_1 , new_n4974 , new_n5025_1 );
nor  g02678 ( new_n5027 , new_n4971 , new_n5026_1 );
nor  g02679 ( new_n5028 , new_n4970 , new_n5027 );
xor  g02680 ( n332 , new_n4967_1 , new_n5028 );
xnor g02681 ( new_n5030 , new_n2361_1 , n18295 );
nor  g02682 ( new_n5031_1 , n6502 , n19494 );
or   g02683 ( new_n5032 , new_n3116 , new_n2907 );
not  g02684 ( new_n5033 , n6502 );
xnor g02685 ( new_n5034 , new_n5033 , n19494 );
and  g02686 ( new_n5035 , new_n5032 , new_n5034 );
nor  g02687 ( new_n5036 , new_n5031_1 , new_n5035 );
xnor g02688 ( new_n5037 , new_n5030 , new_n5036 );
not  g02689 ( new_n5038 , new_n5037 );
xnor g02690 ( new_n5039 , n8381 , new_n5038 );
not  g02691 ( new_n5040 , n20235 );
xnor g02692 ( new_n5041 , new_n3116 , n15780 );
not  g02693 ( new_n5042 , new_n5041 );
nor  g02694 ( new_n5043 , n12495 , new_n5042 );
and  g02695 ( new_n5044 , new_n5040 , new_n5043 );
xnor g02696 ( new_n5045 , n20235 , new_n5043 );
not  g02697 ( new_n5046_1 , new_n5045 );
nor  g02698 ( new_n5047 , new_n3116 , new_n2907 );
xnor g02699 ( new_n5048 , new_n5047 , new_n5034 );
nor  g02700 ( new_n5049 , new_n5046_1 , new_n5048 );
nor  g02701 ( new_n5050 , new_n5044 , new_n5049 );
xnor g02702 ( new_n5051 , new_n5039 , new_n5050 );
not  g02703 ( new_n5052 , new_n5051 );
not  g02704 ( new_n5053 , n23146 );
nor  g02705 ( new_n5054 , new_n3304 , n21654 );
xnor g02706 ( new_n5055 , n23842 , n25471 );
xnor g02707 ( new_n5056 , new_n5054 , new_n5055 );
not  g02708 ( new_n5057 , new_n5056 );
nor  g02709 ( new_n5058 , new_n5053 , new_n5057 );
xnor g02710 ( new_n5059 , new_n3304 , n21654 );
and  g02711 ( new_n5060_1 , n17968 , new_n5059 );
xnor g02712 ( new_n5061 , n23146 , new_n5057 );
and  g02713 ( new_n5062_1 , new_n5060_1 , new_n5061 );
nor  g02714 ( new_n5063 , new_n5058 , new_n5062_1 );
not  g02715 ( new_n5064_1 , n3828 );
xnor g02716 ( new_n5065 , new_n5064_1 , n15053 );
not  g02717 ( new_n5066 , n25471 );
nor  g02718 ( new_n5067 , n23842 , new_n5066 );
and  g02719 ( new_n5068 , new_n5054 , new_n5055 );
nor  g02720 ( new_n5069 , new_n5067 , new_n5068 );
xor  g02721 ( new_n5070 , new_n5065 , new_n5069 );
xnor g02722 ( new_n5071 , n11184 , new_n5070 );
xnor g02723 ( new_n5072 , new_n5063 , new_n5071 );
xnor g02724 ( new_n5073 , new_n5052 , new_n5072 );
not  g02725 ( new_n5074 , new_n5061 );
xnor g02726 ( new_n5075 , new_n5060_1 , new_n5074 );
not  g02727 ( new_n5076 , new_n5048 );
xnor g02728 ( new_n5077_1 , new_n5046_1 , new_n5076 );
not  g02729 ( new_n5078 , new_n5077_1 );
nor  g02730 ( new_n5079 , new_n5075 , new_n5078 );
not  g02731 ( new_n5080 , n12495 );
xnor g02732 ( new_n5081 , new_n5080 , new_n5042 );
xnor g02733 ( new_n5082_1 , n16502 , n21654 );
xnor g02734 ( new_n5083 , n17968 , new_n5082_1 );
not  g02735 ( new_n5084 , new_n5083 );
nor  g02736 ( new_n5085 , new_n5081 , new_n5084 );
xnor g02737 ( new_n5086 , new_n5075 , new_n5078 );
nor  g02738 ( new_n5087 , new_n5085 , new_n5086 );
nor  g02739 ( new_n5088 , new_n5079 , new_n5087 );
xnor g02740 ( n357 , new_n5073 , new_n5088 );
xnor g02741 ( new_n5090 , new_n2367 , n22309 );
nor  g02742 ( new_n5091 , new_n2367 , new_n4626 );
xnor g02743 ( new_n5092 , new_n2363_1 , n25073 );
xnor g02744 ( new_n5093 , new_n5091 , new_n5092 );
not  g02745 ( new_n5094 , new_n5093 );
nor  g02746 ( new_n5095 , new_n5090 , new_n5094 );
not  g02747 ( new_n5096 , new_n5095 );
xnor g02748 ( new_n5097 , new_n2359 , n18171 );
nor  g02749 ( new_n5098_1 , n20138 , n25073 );
or   g02750 ( new_n5099 , new_n2367 , new_n4626 );
and  g02751 ( new_n5100 , new_n5099 , new_n5092 );
nor  g02752 ( new_n5101_1 , new_n5098_1 , new_n5100 );
xnor g02753 ( new_n5102 , new_n5097 , new_n5101_1 );
not  g02754 ( new_n5103 , new_n5102 );
nor  g02755 ( new_n5104 , new_n5096 , new_n5103 );
not  g02756 ( new_n5105 , new_n5104 );
not  g02757 ( new_n5106 , n3136 );
xnor g02758 ( new_n5107 , new_n5106 , n5752 );
nor  g02759 ( new_n5108 , n6385 , n18171 );
or   g02760 ( new_n5109 , new_n5098_1 , new_n5100 );
and  g02761 ( new_n5110 , new_n5097 , new_n5109 );
nor  g02762 ( new_n5111 , new_n5108 , new_n5110 );
xnor g02763 ( new_n5112 , new_n5107 , new_n5111 );
not  g02764 ( new_n5113 , new_n5112 );
nor  g02765 ( new_n5114 , new_n5105 , new_n5113 );
not  g02766 ( new_n5115_1 , new_n5114 );
not  g02767 ( new_n5116 , n9557 );
xnor g02768 ( new_n5117 , new_n5116 , n16158 );
nor  g02769 ( new_n5118 , n3136 , n5752 );
or   g02770 ( new_n5119 , new_n5108 , new_n5110 );
and  g02771 ( new_n5120_1 , new_n5107 , new_n5119 );
nor  g02772 ( new_n5121 , new_n5118 , new_n5120_1 );
xnor g02773 ( new_n5122 , new_n5117 , new_n5121 );
not  g02774 ( new_n5123 , new_n5122 );
nor  g02775 ( new_n5124 , new_n5115_1 , new_n5123 );
not  g02776 ( new_n5125 , n20604 );
xnor g02777 ( new_n5126 , new_n5125 , n25643 );
nor  g02778 ( new_n5127 , n9557 , n16158 );
or   g02779 ( new_n5128_1 , new_n5118 , new_n5120_1 );
and  g02780 ( new_n5129 , new_n5117 , new_n5128_1 );
nor  g02781 ( new_n5130 , new_n5127 , new_n5129 );
xnor g02782 ( new_n5131_1 , new_n5126 , new_n5130 );
not  g02783 ( new_n5132 , new_n5131_1 );
xnor g02784 ( new_n5133 , new_n5124 , new_n5132 );
xnor g02785 ( new_n5134 , new_n3153 , new_n5133 );
xnor g02786 ( new_n5135 , new_n5114 , new_n5123 );
nor  g02787 ( new_n5136 , new_n3157 , new_n5135 );
xnor g02788 ( new_n5137 , new_n3157 , new_n5135 );
xnor g02789 ( new_n5138 , new_n5104 , new_n5113 );
nor  g02790 ( new_n5139 , new_n3163 , new_n5138 );
xnor g02791 ( new_n5140_1 , new_n3160 , new_n5138 );
xnor g02792 ( new_n5141 , new_n5095 , new_n5103 );
and  g02793 ( new_n5142 , new_n3165 , new_n5141 );
not  g02794 ( new_n5143 , new_n5090 );
nor  g02795 ( new_n5144 , new_n3170 , new_n5143 );
nor  g02796 ( new_n5145 , new_n3260_1 , new_n5144 );
or   g02797 ( new_n5146 , n9251 , n22309 );
and  g02798 ( new_n5147 , new_n5146 , new_n5100 );
or   g02799 ( new_n5148 , new_n5095 , new_n5147 );
and  g02800 ( new_n5149 , new_n3119 , new_n5144 );
nor  g02801 ( new_n5150 , new_n5145 , new_n5149 );
and  g02802 ( new_n5151 , new_n5148 , new_n5150 );
nor  g02803 ( new_n5152 , new_n5145 , new_n5151 );
xnor g02804 ( new_n5153 , new_n3166 , new_n5141 );
and  g02805 ( new_n5154 , new_n5152 , new_n5153 );
nor  g02806 ( new_n5155 , new_n5142 , new_n5154 );
and  g02807 ( new_n5156 , new_n5140_1 , new_n5155 );
nor  g02808 ( new_n5157 , new_n5139 , new_n5156 );
nor  g02809 ( new_n5158_1 , new_n5137 , new_n5157 );
nor  g02810 ( new_n5159 , new_n5136 , new_n5158_1 );
xnor g02811 ( new_n5160 , new_n5134 , new_n5159 );
not  g02812 ( new_n5161 , new_n5160 );
xnor g02813 ( new_n5162 , n4119 , n5255 );
not  g02814 ( new_n5163 , n21649 );
nor  g02815 ( new_n5164 , n14510 , new_n5163 );
xnor g02816 ( new_n5165 , n14510 , n21649 );
not  g02817 ( new_n5166 , n18274 );
nor  g02818 ( new_n5167 , n13263 , new_n5166 );
xnor g02819 ( new_n5168_1 , n13263 , n18274 );
nor  g02820 ( new_n5169 , n3828 , new_n3446 );
nor  g02821 ( new_n5170 , new_n5064_1 , n20455 );
nor  g02822 ( new_n5171 , new_n3448 , n23842 );
not  g02823 ( new_n5172 , n23842 );
nor  g02824 ( new_n5173 , n1639 , new_n5172 );
nor  g02825 ( new_n5174 , new_n3451_1 , n21654 );
not  g02826 ( new_n5175 , new_n5174 );
nor  g02827 ( new_n5176 , new_n5173 , new_n5175 );
nor  g02828 ( new_n5177 , new_n5171 , new_n5176 );
nor  g02829 ( new_n5178 , new_n5170 , new_n5177 );
nor  g02830 ( new_n5179 , new_n5169 , new_n5178 );
and  g02831 ( new_n5180 , new_n5168_1 , new_n5179 );
or   g02832 ( new_n5181 , new_n5167 , new_n5180 );
and  g02833 ( new_n5182 , new_n5165 , new_n5181 );
or   g02834 ( new_n5183 , new_n5164 , new_n5182 );
xor  g02835 ( new_n5184_1 , new_n5162 , new_n5183 );
xnor g02836 ( new_n5185 , new_n5161 , new_n5184_1 );
xor  g02837 ( new_n5186 , new_n5165 , new_n5181 );
xnor g02838 ( new_n5187 , new_n5137 , new_n5157 );
nor  g02839 ( new_n5188 , new_n5186 , new_n5187 );
xnor g02840 ( new_n5189 , new_n5186 , new_n5187 );
xnor g02841 ( new_n5190 , new_n5140_1 , new_n5155 );
not  g02842 ( new_n5191 , new_n5190 );
xnor g02843 ( new_n5192 , new_n5168_1 , new_n5179 );
and  g02844 ( new_n5193 , new_n5191 , new_n5192 );
xnor g02845 ( new_n5194 , new_n5191 , new_n5192 );
xnor g02846 ( new_n5195 , new_n5152 , new_n5153 );
xnor g02847 ( new_n5196 , n3828 , n20455 );
xnor g02848 ( new_n5197 , new_n5177 , new_n5196 );
and  g02849 ( new_n5198 , new_n5195 , new_n5197 );
xnor g02850 ( new_n5199 , new_n5195 , new_n5197 );
xnor g02851 ( new_n5200 , n16968 , n21654 );
xnor g02852 ( new_n5201 , new_n3170 , new_n5090 );
not  g02853 ( new_n5202 , new_n5201 );
or   g02854 ( new_n5203 , new_n5200 , new_n5202 );
xnor g02855 ( new_n5204 , n1639 , n23842 );
xnor g02856 ( new_n5205 , new_n5175 , new_n5204 );
and  g02857 ( new_n5206 , new_n5203 , new_n5205 );
xnor g02858 ( new_n5207 , new_n5148 , new_n5150 );
not  g02859 ( new_n5208 , new_n5207 );
xor  g02860 ( new_n5209 , new_n5203 , new_n5205 );
and  g02861 ( new_n5210 , new_n5208 , new_n5209 );
nor  g02862 ( new_n5211_1 , new_n5206 , new_n5210 );
nor  g02863 ( new_n5212 , new_n5199 , new_n5211_1 );
nor  g02864 ( new_n5213_1 , new_n5198 , new_n5212 );
nor  g02865 ( new_n5214 , new_n5194 , new_n5213_1 );
nor  g02866 ( new_n5215 , new_n5193 , new_n5214 );
nor  g02867 ( new_n5216 , new_n5189 , new_n5215 );
nor  g02868 ( new_n5217 , new_n5188 , new_n5216 );
xor  g02869 ( n422 , new_n5185 , new_n5217 );
nor  g02870 ( new_n5219 , n20794 , n23333 );
not  g02871 ( new_n5220 , new_n5219 );
nor  g02872 ( new_n5221 , n14603 , new_n5220 );
not  g02873 ( new_n5222 , new_n5221 );
nor  g02874 ( new_n5223 , n18737 , new_n5222 );
not  g02875 ( new_n5224 , new_n5223 );
nor  g02876 ( new_n5225 , n21471 , new_n5224 );
not  g02877 ( new_n5226_1 , new_n5225 );
nor  g02878 ( new_n5227 , n25738 , new_n5226_1 );
not  g02879 ( new_n5228_1 , new_n5227 );
nor  g02880 ( new_n5229 , n5302 , new_n5228_1 );
not  g02881 ( new_n5230 , new_n5229 );
nor  g02882 ( new_n5231 , n3228 , new_n5230 );
xnor g02883 ( new_n5232 , n337 , new_n5231 );
xnor g02884 ( new_n5233 , new_n3140 , new_n5232 );
xnor g02885 ( new_n5234 , n3228 , new_n5229 );
nor  g02886 ( new_n5235 , n26036 , new_n5234 );
xnor g02887 ( new_n5236 , n26036 , new_n5234 );
xnor g02888 ( new_n5237 , n5302 , new_n5227 );
nor  g02889 ( new_n5238 , n19770 , new_n5237 );
xnor g02890 ( new_n5239 , new_n3148 , new_n5237 );
xnor g02891 ( new_n5240 , n25738 , new_n5225 );
nor  g02892 ( new_n5241 , n8782 , new_n5240 );
xnor g02893 ( new_n5242 , new_n3152 , new_n5240 );
xnor g02894 ( new_n5243 , n21471 , new_n5223 );
nor  g02895 ( new_n5244 , n8678 , new_n5243 );
xnor g02896 ( new_n5245 , n8678 , new_n5243 );
xnor g02897 ( new_n5246 , n18737 , new_n5221 );
nor  g02898 ( new_n5247 , n1432 , new_n5246 );
xnor g02899 ( new_n5248 , n14603 , new_n5219 );
nor  g02900 ( new_n5249 , n21599 , new_n5248 );
xor  g02901 ( new_n5250 , n21599 , new_n5248 );
xnor g02902 ( new_n5251 , new_n3307 , n23333 );
nor  g02903 ( new_n5252 , n25336 , new_n5251 );
or   g02904 ( new_n5253 , new_n3256 , new_n3305 );
xnor g02905 ( new_n5254 , new_n3169 , new_n5251 );
and  g02906 ( new_n5255_1 , new_n5253 , new_n5254 );
or   g02907 ( new_n5256_1 , new_n5252 , new_n5255_1 );
and  g02908 ( new_n5257 , new_n5250 , new_n5256_1 );
or   g02909 ( new_n5258 , new_n5249 , new_n5257 );
xnor g02910 ( new_n5259 , new_n3162 , new_n5246 );
and  g02911 ( new_n5260 , new_n5258 , new_n5259 );
nor  g02912 ( new_n5261 , new_n5247 , new_n5260 );
nor  g02913 ( new_n5262 , new_n5245 , new_n5261 );
or   g02914 ( new_n5263 , new_n5244 , new_n5262 );
and  g02915 ( new_n5264 , new_n5242 , new_n5263 );
or   g02916 ( new_n5265_1 , new_n5241 , new_n5264 );
and  g02917 ( new_n5266 , new_n5239 , new_n5265_1 );
nor  g02918 ( new_n5267 , new_n5238 , new_n5266 );
nor  g02919 ( new_n5268 , new_n5236 , new_n5267 );
or   g02920 ( new_n5269 , new_n5235 , new_n5268 );
xor  g02921 ( new_n5270 , new_n5233 , new_n5269 );
xnor g02922 ( new_n5271 , n9967 , n22379 );
nor  g02923 ( new_n5272 , n1662 , n20946 );
xnor g02924 ( new_n5273_1 , new_n2850 , n20946 );
nor  g02925 ( new_n5274_1 , n7751 , n12875 );
not  g02926 ( new_n5275 , n7751 );
xnor g02927 ( new_n5276 , new_n5275 , n12875 );
nor  g02928 ( new_n5277 , n2035 , n26823 );
xnor g02929 ( new_n5278 , new_n2856 , n26823 );
nor  g02930 ( new_n5279 , n4812 , n5213 );
not  g02931 ( new_n5280 , n4812 );
xnor g02932 ( new_n5281 , new_n5280 , n5213 );
nor  g02933 ( new_n5282 , n4665 , n24278 );
xnor g02934 ( new_n5283 , new_n2862 , n24278 );
nor  g02935 ( new_n5284 , n19005 , n24618 );
xnor g02936 ( new_n5285 , new_n2866 , n24618 );
nor  g02937 ( new_n5286 , n3952 , n4326 );
not  g02938 ( new_n5287 , n5438 );
or   g02939 ( new_n5288 , new_n5287 , new_n2448 );
xnor g02940 ( new_n5289 , new_n2443 , n4326 );
and  g02941 ( new_n5290 , new_n5288 , new_n5289 );
or   g02942 ( new_n5291 , new_n5286 , new_n5290 );
and  g02943 ( new_n5292 , new_n5285 , new_n5291 );
or   g02944 ( new_n5293 , new_n5284 , new_n5292 );
and  g02945 ( new_n5294 , new_n5283 , new_n5293 );
or   g02946 ( new_n5295 , new_n5282 , new_n5294 );
and  g02947 ( new_n5296 , new_n5281 , new_n5295 );
or   g02948 ( new_n5297 , new_n5279 , new_n5296 );
and  g02949 ( new_n5298 , new_n5278 , new_n5297 );
or   g02950 ( new_n5299 , new_n5277 , new_n5298 );
and  g02951 ( new_n5300_1 , new_n5276 , new_n5299 );
or   g02952 ( new_n5301 , new_n5274_1 , new_n5300_1 );
and  g02953 ( new_n5302_1 , new_n5273_1 , new_n5301 );
nor  g02954 ( new_n5303 , new_n5272 , new_n5302_1 );
xnor g02955 ( new_n5304 , new_n5271 , new_n5303 );
xnor g02956 ( new_n5305 , new_n3091 , n10763 );
nor  g02957 ( new_n5306 , n7437 , n13367 );
xnor g02958 ( new_n5307 , new_n2890 , n13367 );
nor  g02959 ( new_n5308 , n932 , n20700 );
xnor g02960 ( new_n5309 , n932 , n20700 );
nor  g02961 ( new_n5310 , n6691 , n7099 );
xnor g02962 ( new_n5311 , n6691 , n7099 );
nor  g02963 ( new_n5312 , n3260 , n12811 );
xnor g02964 ( new_n5313 , new_n3106 , n12811 );
nor  g02965 ( new_n5314 , n1118 , n20489 );
xnor g02966 ( new_n5315 , n1118 , n20489 );
nor  g02967 ( new_n5316 , n2355 , n25974 );
xnor g02968 ( new_n5317 , n2355 , n25974 );
nor  g02969 ( new_n5318 , n1630 , n11121 );
nor  g02970 ( new_n5319 , new_n2906 , new_n3117 );
xnor g02971 ( new_n5320 , n1630 , n11121 );
nor  g02972 ( new_n5321 , new_n5319 , new_n5320 );
nor  g02973 ( new_n5322 , new_n5318 , new_n5321 );
nor  g02974 ( new_n5323 , new_n5317 , new_n5322 );
nor  g02975 ( new_n5324 , new_n5316 , new_n5323 );
nor  g02976 ( new_n5325_1 , new_n5315 , new_n5324 );
or   g02977 ( new_n5326 , new_n5314 , new_n5325_1 );
and  g02978 ( new_n5327 , new_n5313 , new_n5326 );
nor  g02979 ( new_n5328 , new_n5312 , new_n5327 );
nor  g02980 ( new_n5329 , new_n5311 , new_n5328 );
nor  g02981 ( new_n5330_1 , new_n5310 , new_n5329 );
nor  g02982 ( new_n5331 , new_n5309 , new_n5330_1 );
or   g02983 ( new_n5332 , new_n5308 , new_n5331 );
and  g02984 ( new_n5333 , new_n5307 , new_n5332 );
or   g02985 ( new_n5334 , new_n5306 , new_n5333 );
xor  g02986 ( new_n5335 , new_n5305 , new_n5334 );
xnor g02987 ( new_n5336 , new_n5304 , new_n5335 );
nor  g02988 ( new_n5337_1 , new_n5308 , new_n5331 );
xnor g02989 ( new_n5338 , new_n5307 , new_n5337_1 );
nor  g02990 ( new_n5339 , new_n5274_1 , new_n5300_1 );
xnor g02991 ( new_n5340 , new_n5273_1 , new_n5339 );
not  g02992 ( new_n5341 , new_n5340 );
nor  g02993 ( new_n5342 , new_n5338 , new_n5341 );
xnor g02994 ( new_n5343 , new_n5338 , new_n5340 );
xnor g02995 ( new_n5344 , new_n5309 , new_n5330_1 );
nor  g02996 ( new_n5345 , new_n5277 , new_n5298 );
xnor g02997 ( new_n5346 , new_n5276 , new_n5345 );
nor  g02998 ( new_n5347 , new_n5344 , new_n5346 );
not  g02999 ( new_n5348 , new_n5346 );
xnor g03000 ( new_n5349 , new_n5344 , new_n5348 );
xnor g03001 ( new_n5350 , new_n5311 , new_n5328 );
nor  g03002 ( new_n5351_1 , new_n5279 , new_n5296 );
xnor g03003 ( new_n5352 , new_n5278 , new_n5351_1 );
nor  g03004 ( new_n5353_1 , new_n5350 , new_n5352 );
xnor g03005 ( new_n5354 , new_n5315 , new_n5324 );
nor  g03006 ( new_n5355 , new_n5284 , new_n5292 );
xnor g03007 ( new_n5356 , new_n5283 , new_n5355 );
nor  g03008 ( new_n5357 , new_n5354 , new_n5356 );
not  g03009 ( new_n5358 , new_n5356 );
xnor g03010 ( new_n5359 , new_n5354 , new_n5358 );
xnor g03011 ( new_n5360 , new_n5317 , new_n5322 );
nor  g03012 ( new_n5361 , new_n5286 , new_n5290 );
xnor g03013 ( new_n5362 , new_n5285 , new_n5361 );
nor  g03014 ( new_n5363 , new_n5360 , new_n5362 );
nor  g03015 ( new_n5364 , new_n5287 , new_n2448 );
xnor g03016 ( new_n5365 , new_n5364 , new_n5289 );
xnor g03017 ( new_n5366 , new_n5319 , new_n5320 );
nor  g03018 ( new_n5367 , new_n5365 , new_n5366 );
xnor g03019 ( new_n5368 , new_n5287 , n12315 );
not  g03020 ( new_n5369 , new_n5368 );
xnor g03021 ( new_n5370 , new_n2906 , n16217 );
nor  g03022 ( new_n5371 , new_n5369 , new_n5370 );
not  g03023 ( new_n5372 , new_n5365 );
xnor g03024 ( new_n5373 , new_n5372 , new_n5366 );
and  g03025 ( new_n5374 , new_n5371 , new_n5373 );
or   g03026 ( new_n5375 , new_n5367 , new_n5374 );
not  g03027 ( new_n5376_1 , new_n5362 );
xnor g03028 ( new_n5377 , new_n5360 , new_n5376_1 );
and  g03029 ( new_n5378 , new_n5375 , new_n5377 );
or   g03030 ( new_n5379 , new_n5363 , new_n5378 );
and  g03031 ( new_n5380 , new_n5359 , new_n5379 );
nor  g03032 ( new_n5381 , new_n5357 , new_n5380 );
xor  g03033 ( new_n5382 , new_n5313 , new_n5326 );
not  g03034 ( new_n5383 , new_n5382 );
and  g03035 ( new_n5384 , new_n5381 , new_n5383 );
xnor g03036 ( new_n5385 , new_n5381 , new_n5383 );
nor  g03037 ( new_n5386_1 , new_n5282 , new_n5294 );
xnor g03038 ( new_n5387 , new_n5281 , new_n5386_1 );
not  g03039 ( new_n5388 , new_n5387 );
nor  g03040 ( new_n5389 , new_n5385 , new_n5388 );
nor  g03041 ( new_n5390 , new_n5384 , new_n5389 );
not  g03042 ( new_n5391 , new_n5352 );
xnor g03043 ( new_n5392 , new_n5350 , new_n5391 );
and  g03044 ( new_n5393 , new_n5390 , new_n5392 );
or   g03045 ( new_n5394 , new_n5353_1 , new_n5393 );
and  g03046 ( new_n5395 , new_n5349 , new_n5394 );
nor  g03047 ( new_n5396 , new_n5347 , new_n5395 );
and  g03048 ( new_n5397 , new_n5343 , new_n5396 );
nor  g03049 ( new_n5398 , new_n5342 , new_n5397 );
xnor g03050 ( new_n5399_1 , new_n5336 , new_n5398 );
not  g03051 ( new_n5400_1 , new_n5399_1 );
xnor g03052 ( new_n5401 , new_n5270 , new_n5400_1 );
xnor g03053 ( new_n5402 , new_n5236 , new_n5267 );
xnor g03054 ( new_n5403_1 , new_n5343 , new_n5396 );
not  g03055 ( new_n5404 , new_n5403_1 );
nor  g03056 ( new_n5405 , new_n5402 , new_n5404 );
xnor g03057 ( new_n5406 , new_n5402 , new_n5404 );
xor  g03058 ( new_n5407 , new_n5239 , new_n5265_1 );
nor  g03059 ( new_n5408 , new_n5353_1 , new_n5393 );
xnor g03060 ( new_n5409 , new_n5349 , new_n5408 );
and  g03061 ( new_n5410 , new_n5407 , new_n5409 );
xnor g03062 ( new_n5411 , new_n5407 , new_n5409 );
xor  g03063 ( new_n5412 , new_n5242 , new_n5263 );
xnor g03064 ( new_n5413 , new_n5390 , new_n5392 );
not  g03065 ( new_n5414 , new_n5413 );
and  g03066 ( new_n5415 , new_n5412 , new_n5414 );
xnor g03067 ( new_n5416 , new_n5412 , new_n5414 );
xnor g03068 ( new_n5417 , new_n5245 , new_n5261 );
xnor g03069 ( new_n5418 , new_n5385 , new_n5387 );
nor  g03070 ( new_n5419 , new_n5417 , new_n5418 );
xnor g03071 ( new_n5420 , new_n5417 , new_n5418 );
xor  g03072 ( new_n5421 , new_n5359 , new_n5379 );
xor  g03073 ( new_n5422 , new_n5258 , new_n5259 );
and  g03074 ( new_n5423 , new_n5421 , new_n5422 );
xnor g03075 ( new_n5424 , new_n5421 , new_n5422 );
not  g03076 ( new_n5425 , new_n5424 );
xor  g03077 ( new_n5426 , new_n5250 , new_n5256_1 );
xor  g03078 ( new_n5427 , new_n5375 , new_n5377 );
nor  g03079 ( new_n5428 , new_n5426 , new_n5427 );
xor  g03080 ( new_n5429 , new_n5426 , new_n5427 );
xnor g03081 ( new_n5430_1 , new_n5371 , new_n5373 );
nor  g03082 ( new_n5431 , new_n5254 , new_n5430_1 );
not  g03083 ( new_n5432 , new_n5430_1 );
xor  g03084 ( new_n5433 , new_n5253 , new_n5254 );
nor  g03085 ( new_n5434 , new_n5432 , new_n5433 );
xnor g03086 ( new_n5435 , n11424 , n23333 );
xnor g03087 ( new_n5436 , new_n5368 , new_n5370 );
nor  g03088 ( new_n5437 , new_n5435 , new_n5436 );
nor  g03089 ( new_n5438_1 , new_n5434 , new_n5437 );
nor  g03090 ( new_n5439_1 , new_n5431 , new_n5438_1 );
and  g03091 ( new_n5440 , new_n5429 , new_n5439_1 );
nor  g03092 ( new_n5441 , new_n5428 , new_n5440 );
and  g03093 ( new_n5442 , new_n5425 , new_n5441 );
nor  g03094 ( new_n5443_1 , new_n5423 , new_n5442 );
nor  g03095 ( new_n5444 , new_n5420 , new_n5443_1 );
nor  g03096 ( new_n5445 , new_n5419 , new_n5444 );
nor  g03097 ( new_n5446 , new_n5416 , new_n5445 );
nor  g03098 ( new_n5447 , new_n5415 , new_n5446 );
nor  g03099 ( new_n5448 , new_n5411 , new_n5447 );
nor  g03100 ( new_n5449 , new_n5410 , new_n5448 );
nor  g03101 ( new_n5450 , new_n5406 , new_n5449 );
nor  g03102 ( new_n5451_1 , new_n5405 , new_n5450 );
xor  g03103 ( n431 , new_n5401 , new_n5451_1 );
not  g03104 ( new_n5453 , n23895 );
nor  g03105 ( new_n5454 , n8614 , new_n5453 );
xnor g03106 ( new_n5455 , n8614 , n23895 );
not  g03107 ( new_n5456 , n17351 );
nor  g03108 ( new_n5457 , n15182 , new_n5456 );
xnor g03109 ( new_n5458 , n15182 , n17351 );
not  g03110 ( new_n5459 , n11736 );
nor  g03111 ( new_n5460 , new_n5459 , n27037 );
xnor g03112 ( new_n5461 , n11736 , n27037 );
not  g03113 ( new_n5462 , n23200 );
nor  g03114 ( new_n5463 , n8964 , new_n5462 );
xnor g03115 ( new_n5464 , n8964 , n23200 );
not  g03116 ( new_n5465 , n17959 );
nor  g03117 ( new_n5466 , new_n5465 , n20151 );
xnor g03118 ( new_n5467 , n17959 , n20151 );
not  g03119 ( new_n5468 , n7566 );
nor  g03120 ( new_n5469 , new_n5468 , n7693 );
xnor g03121 ( new_n5470 , n7566 , n7693 );
not  g03122 ( new_n5471 , n7731 );
nor  g03123 ( new_n5472_1 , new_n5471 , n10405 );
xnor g03124 ( new_n5473 , n7731 , n10405 );
nor  g03125 ( new_n5474 , new_n4106 , n12341 );
not  g03126 ( new_n5475 , n12341 );
nor  g03127 ( new_n5476 , n11302 , new_n5475 );
nor  g03128 ( new_n5477 , new_n4111 , n20986 );
not  g03129 ( new_n5478 , n20986 );
or   g03130 ( new_n5479 , n17090 , new_n5478 );
nor  g03131 ( new_n5480 , new_n4030 , n12384 );
and  g03132 ( new_n5481 , new_n5479 , new_n5480 );
nor  g03133 ( new_n5482 , new_n5477 , new_n5481 );
nor  g03134 ( new_n5483 , new_n5476 , new_n5482 );
nor  g03135 ( new_n5484 , new_n5474 , new_n5483 );
and  g03136 ( new_n5485_1 , new_n5473 , new_n5484 );
or   g03137 ( new_n5486 , new_n5472_1 , new_n5485_1 );
and  g03138 ( new_n5487 , new_n5470 , new_n5486 );
or   g03139 ( new_n5488 , new_n5469 , new_n5487 );
and  g03140 ( new_n5489 , new_n5467 , new_n5488 );
or   g03141 ( new_n5490 , new_n5466 , new_n5489 );
and  g03142 ( new_n5491 , new_n5464 , new_n5490 );
or   g03143 ( new_n5492 , new_n5463 , new_n5491 );
and  g03144 ( new_n5493 , new_n5461 , new_n5492 );
or   g03145 ( new_n5494 , new_n5460 , new_n5493 );
and  g03146 ( new_n5495 , new_n5458 , new_n5494 );
or   g03147 ( new_n5496 , new_n5457 , new_n5495 );
and  g03148 ( new_n5497 , new_n5455 , new_n5496 );
nor  g03149 ( new_n5498 , new_n5454 , new_n5497 );
not  g03150 ( new_n5499 , new_n5498 );
not  g03151 ( new_n5500 , n13494 );
nor  g03152 ( new_n5501 , new_n5500 , n18880 );
xnor g03153 ( new_n5502 , n13494 , n18880 );
not  g03154 ( new_n5503 , n25345 );
nor  g03155 ( new_n5504 , new_n5503 , n25475 );
xnor g03156 ( new_n5505 , n25345 , n25475 );
not  g03157 ( new_n5506 , n9655 );
nor  g03158 ( new_n5507 , new_n5506 , n23849 );
xnor g03159 ( new_n5508 , n9655 , n23849 );
and  g03160 ( new_n5509 , new_n4442 , n13490 );
xnor g03161 ( new_n5510 , n12446 , n13490 );
not  g03162 ( new_n5511 , n22660 );
nor  g03163 ( new_n5512 , n11011 , new_n5511 );
xnor g03164 ( new_n5513 , n11011 , n22660 );
not  g03165 ( new_n5514 , n1777 );
nor  g03166 ( new_n5515 , new_n5514 , n16029 );
xnor g03167 ( new_n5516 , n1777 , n16029 );
not  g03168 ( new_n5517_1 , n8745 );
nor  g03169 ( new_n5518 , new_n5517_1 , n16476 );
xnor g03170 ( new_n5519 , n8745 , n16476 );
nor  g03171 ( new_n5520 , new_n3947 , n15636 );
nor  g03172 ( new_n5521_1 , n11615 , new_n2441 );
nor  g03173 ( new_n5522 , n20077 , new_n3949 );
nor  g03174 ( new_n5523 , new_n2444_1 , n22433 );
or   g03175 ( new_n5524_1 , n6794 , new_n3952_1 );
nor  g03176 ( new_n5525 , new_n5523 , new_n5524_1 );
nor  g03177 ( new_n5526 , new_n5522 , new_n5525 );
nor  g03178 ( new_n5527 , new_n5521_1 , new_n5526 );
nor  g03179 ( new_n5528 , new_n5520 , new_n5527 );
and  g03180 ( new_n5529 , new_n5519 , new_n5528 );
or   g03181 ( new_n5530 , new_n5518 , new_n5529 );
and  g03182 ( new_n5531 , new_n5516 , new_n5530 );
or   g03183 ( new_n5532_1 , new_n5515 , new_n5531 );
and  g03184 ( new_n5533 , new_n5513 , new_n5532_1 );
or   g03185 ( new_n5534 , new_n5512 , new_n5533 );
and  g03186 ( new_n5535 , new_n5510 , new_n5534 );
or   g03187 ( new_n5536 , new_n5509 , new_n5535 );
and  g03188 ( new_n5537 , new_n5508 , new_n5536 );
or   g03189 ( new_n5538 , new_n5507 , new_n5537 );
and  g03190 ( new_n5539 , new_n5505 , new_n5538 );
or   g03191 ( new_n5540 , new_n5504 , new_n5539 );
and  g03192 ( new_n5541 , new_n5502 , new_n5540 );
nor  g03193 ( new_n5542 , new_n5501 , new_n5541 );
nor  g03194 ( new_n5543 , new_n5504 , new_n5539 );
xnor g03195 ( new_n5544 , new_n5502 , new_n5543 );
nor  g03196 ( new_n5545 , n583 , n22173 );
not  g03197 ( new_n5546 , new_n5545 );
nor  g03198 ( new_n5547 , n2146 , new_n5546 );
not  g03199 ( new_n5548 , new_n5547 );
nor  g03200 ( new_n5549 , n23974 , new_n5548 );
not  g03201 ( new_n5550 , new_n5549 );
nor  g03202 ( new_n5551 , n3909 , new_n5550 );
not  g03203 ( new_n5552 , new_n5551 );
nor  g03204 ( new_n5553 , n20429 , new_n5552 );
not  g03205 ( new_n5554 , new_n5553 );
nor  g03206 ( new_n5555 , n22554 , new_n5554 );
not  g03207 ( new_n5556 , new_n5555 );
nor  g03208 ( new_n5557 , n23913 , new_n5556 );
xnor g03209 ( new_n5558 , n26797 , new_n5557 );
nor  g03210 ( new_n5559 , n10201 , new_n5558 );
not  g03211 ( new_n5560 , n10201 );
xnor g03212 ( new_n5561 , new_n5560 , new_n5558 );
xnor g03213 ( new_n5562 , n23913 , new_n5555 );
nor  g03214 ( new_n5563 , n10593 , new_n5562 );
not  g03215 ( new_n5564_1 , n10593 );
xnor g03216 ( new_n5565 , new_n5564_1 , new_n5562 );
xnor g03217 ( new_n5566 , n22554 , new_n5553 );
nor  g03218 ( new_n5567 , n18290 , new_n5566 );
not  g03219 ( new_n5568 , n18290 );
xnor g03220 ( new_n5569 , new_n5568 , new_n5566 );
xnor g03221 ( new_n5570 , n20429 , new_n5551 );
nor  g03222 ( new_n5571 , n11580 , new_n5570 );
not  g03223 ( new_n5572 , n11580 );
xnor g03224 ( new_n5573 , new_n5572 , new_n5570 );
xnor g03225 ( new_n5574 , n3909 , new_n5549 );
nor  g03226 ( new_n5575 , n15884 , new_n5574 );
not  g03227 ( new_n5576 , n15884 );
xnor g03228 ( new_n5577 , new_n5576 , new_n5574 );
xnor g03229 ( new_n5578 , n23974 , new_n5547 );
nor  g03230 ( new_n5579_1 , n6356 , new_n5578 );
xnor g03231 ( new_n5580 , n2146 , new_n5545 );
nor  g03232 ( new_n5581 , n27104 , new_n5580 );
not  g03233 ( new_n5582 , n27104 );
xnor g03234 ( new_n5583 , new_n5582 , new_n5580 );
not  g03235 ( new_n5584 , n27188 );
xnor g03236 ( new_n5585 , n583 , n22173 );
and  g03237 ( new_n5586 , new_n5584 , new_n5585 );
not  g03238 ( new_n5587 , n583 );
not  g03239 ( new_n5588 , n6611 );
or   g03240 ( new_n5589 , new_n5587 , new_n5588 );
xnor g03241 ( new_n5590 , n27188 , new_n5585 );
and  g03242 ( new_n5591 , new_n5589 , new_n5590 );
or   g03243 ( new_n5592 , new_n5586 , new_n5591 );
and  g03244 ( new_n5593_1 , new_n5583 , new_n5592 );
or   g03245 ( new_n5594 , new_n5581 , new_n5593_1 );
not  g03246 ( new_n5595 , n6356 );
xnor g03247 ( new_n5596 , new_n5595 , new_n5578 );
and  g03248 ( new_n5597 , new_n5594 , new_n5596 );
or   g03249 ( new_n5598 , new_n5579_1 , new_n5597 );
and  g03250 ( new_n5599 , new_n5577 , new_n5598 );
or   g03251 ( new_n5600 , new_n5575 , new_n5599 );
and  g03252 ( new_n5601 , new_n5573 , new_n5600 );
or   g03253 ( new_n5602 , new_n5571 , new_n5601 );
and  g03254 ( new_n5603_1 , new_n5569 , new_n5602 );
or   g03255 ( new_n5604 , new_n5567 , new_n5603_1 );
and  g03256 ( new_n5605_1 , new_n5565 , new_n5604 );
or   g03257 ( new_n5606 , new_n5563 , new_n5605_1 );
and  g03258 ( new_n5607 , new_n5561 , new_n5606 );
nor  g03259 ( new_n5608 , new_n5559 , new_n5607 );
not  g03260 ( new_n5609_1 , new_n5608 );
not  g03261 ( new_n5610 , n12650 );
not  g03262 ( new_n5611 , n26797 );
and  g03263 ( new_n5612 , new_n5611 , new_n5557 );
xnor g03264 ( new_n5613 , n12702 , new_n5612 );
xnor g03265 ( new_n5614 , new_n5610 , new_n5613 );
xnor g03266 ( new_n5615 , new_n5609_1 , new_n5614 );
nor  g03267 ( new_n5616 , new_n5544 , new_n5615 );
xnor g03268 ( new_n5617 , new_n5544 , new_n5615 );
nor  g03269 ( new_n5618 , new_n5507 , new_n5537 );
xnor g03270 ( new_n5619 , new_n5505 , new_n5618 );
not  g03271 ( new_n5620 , new_n5619 );
xor  g03272 ( new_n5621 , new_n5561 , new_n5606 );
and  g03273 ( new_n5622 , new_n5620 , new_n5621 );
xnor g03274 ( new_n5623 , new_n5620 , new_n5621 );
nor  g03275 ( new_n5624 , new_n5509 , new_n5535 );
xnor g03276 ( new_n5625 , new_n5508 , new_n5624 );
not  g03277 ( new_n5626 , new_n5625 );
xor  g03278 ( new_n5627 , new_n5565 , new_n5604 );
and  g03279 ( new_n5628 , new_n5626 , new_n5627 );
xnor g03280 ( new_n5629 , new_n5626 , new_n5627 );
nor  g03281 ( new_n5630 , new_n5512 , new_n5533 );
xnor g03282 ( new_n5631 , new_n5510 , new_n5630 );
not  g03283 ( new_n5632 , new_n5631 );
xor  g03284 ( new_n5633 , new_n5569 , new_n5602 );
and  g03285 ( new_n5634_1 , new_n5632 , new_n5633 );
xnor g03286 ( new_n5635 , new_n5632 , new_n5633 );
nor  g03287 ( new_n5636 , new_n5515 , new_n5531 );
xnor g03288 ( new_n5637 , new_n5513 , new_n5636 );
not  g03289 ( new_n5638 , new_n5637 );
xor  g03290 ( new_n5639 , new_n5573 , new_n5600 );
and  g03291 ( new_n5640 , new_n5638 , new_n5639 );
xnor g03292 ( new_n5641 , new_n5638 , new_n5639 );
nor  g03293 ( new_n5642 , new_n5518 , new_n5529 );
xnor g03294 ( new_n5643_1 , new_n5516 , new_n5642 );
not  g03295 ( new_n5644 , new_n5643_1 );
xor  g03296 ( new_n5645 , new_n5577 , new_n5598 );
and  g03297 ( new_n5646 , new_n5644 , new_n5645 );
xnor g03298 ( new_n5647 , new_n5644 , new_n5645 );
xor  g03299 ( new_n5648 , new_n5519 , new_n5528 );
not  g03300 ( new_n5649 , new_n5648 );
xor  g03301 ( new_n5650 , new_n5594 , new_n5596 );
and  g03302 ( new_n5651 , new_n5649 , new_n5650 );
xnor g03303 ( new_n5652 , new_n5648 , new_n5650 );
xor  g03304 ( new_n5653 , new_n5583 , new_n5592 );
xnor g03305 ( new_n5654 , n11615 , n15636 );
xnor g03306 ( new_n5655 , new_n5526 , new_n5654 );
nor  g03307 ( new_n5656 , new_n5653 , new_n5655 );
xnor g03308 ( new_n5657 , new_n5653 , new_n5655 );
nor  g03309 ( new_n5658 , new_n5587 , new_n5588 );
xnor g03310 ( new_n5659 , new_n5658 , new_n5590 );
xnor g03311 ( new_n5660 , n20077 , n22433 );
xnor g03312 ( new_n5661 , new_n5524_1 , new_n5660 );
nor  g03313 ( new_n5662 , new_n5659 , new_n5661 );
xnor g03314 ( new_n5663 , n6794 , n14090 );
xnor g03315 ( new_n5664 , n583 , n6611 );
nor  g03316 ( new_n5665 , new_n5663 , new_n5664 );
not  g03317 ( new_n5666 , new_n5661 );
xnor g03318 ( new_n5667 , new_n5659 , new_n5666 );
and  g03319 ( new_n5668 , new_n5665 , new_n5667 );
nor  g03320 ( new_n5669 , new_n5662 , new_n5668 );
nor  g03321 ( new_n5670 , new_n5657 , new_n5669 );
nor  g03322 ( new_n5671 , new_n5656 , new_n5670 );
and  g03323 ( new_n5672 , new_n5652 , new_n5671 );
nor  g03324 ( new_n5673 , new_n5651 , new_n5672 );
nor  g03325 ( new_n5674 , new_n5647 , new_n5673 );
nor  g03326 ( new_n5675 , new_n5646 , new_n5674 );
nor  g03327 ( new_n5676 , new_n5641 , new_n5675 );
nor  g03328 ( new_n5677 , new_n5640 , new_n5676 );
nor  g03329 ( new_n5678 , new_n5635 , new_n5677 );
nor  g03330 ( new_n5679 , new_n5634_1 , new_n5678 );
nor  g03331 ( new_n5680_1 , new_n5629 , new_n5679 );
nor  g03332 ( new_n5681 , new_n5628 , new_n5680_1 );
nor  g03333 ( new_n5682 , new_n5623 , new_n5681 );
nor  g03334 ( new_n5683 , new_n5622 , new_n5682 );
nor  g03335 ( new_n5684 , new_n5617 , new_n5683 );
nor  g03336 ( new_n5685 , new_n5616 , new_n5684 );
not  g03337 ( new_n5686 , n12702 );
and  g03338 ( new_n5687_1 , new_n5686 , new_n5612 );
and  g03339 ( new_n5688 , n12650 , new_n5613 );
nor  g03340 ( new_n5689 , n12650 , new_n5613 );
nor  g03341 ( new_n5690 , new_n5609_1 , new_n5689 );
or   g03342 ( new_n5691 , new_n5688 , new_n5690 );
nor  g03343 ( new_n5692 , new_n5687_1 , new_n5691 );
not  g03344 ( new_n5693 , new_n5692 );
and  g03345 ( new_n5694 , new_n5685 , new_n5693 );
and  g03346 ( new_n5695 , new_n5542 , new_n5694 );
or   g03347 ( new_n5696_1 , new_n5685 , new_n5693 );
nor  g03348 ( new_n5697 , new_n5542 , new_n5696_1 );
nor  g03349 ( new_n5698 , new_n5695 , new_n5697 );
not  g03350 ( new_n5699 , new_n5698 );
xnor g03351 ( new_n5700_1 , new_n5499 , new_n5699 );
xnor g03352 ( new_n5701 , new_n5685 , new_n5692 );
xnor g03353 ( new_n5702 , new_n5542 , new_n5701 );
and  g03354 ( new_n5703 , new_n5498 , new_n5702 );
or   g03355 ( new_n5704_1 , new_n5498 , new_n5702 );
xor  g03356 ( new_n5705 , new_n5455 , new_n5496 );
xnor g03357 ( new_n5706 , new_n5617 , new_n5683 );
nor  g03358 ( new_n5707 , new_n5705 , new_n5706 );
xnor g03359 ( new_n5708 , new_n5705 , new_n5706 );
xor  g03360 ( new_n5709 , new_n5458 , new_n5494 );
xnor g03361 ( new_n5710 , new_n5623 , new_n5681 );
nor  g03362 ( new_n5711 , new_n5709 , new_n5710 );
xnor g03363 ( new_n5712 , new_n5709 , new_n5710 );
xor  g03364 ( new_n5713 , new_n5461 , new_n5492 );
xnor g03365 ( new_n5714 , new_n5629 , new_n5679 );
nor  g03366 ( new_n5715 , new_n5713 , new_n5714 );
xnor g03367 ( new_n5716 , new_n5713 , new_n5714 );
xor  g03368 ( new_n5717 , new_n5464 , new_n5490 );
xnor g03369 ( new_n5718 , new_n5635 , new_n5677 );
nor  g03370 ( new_n5719 , new_n5717 , new_n5718 );
xnor g03371 ( new_n5720 , new_n5717 , new_n5718 );
xor  g03372 ( new_n5721 , new_n5467 , new_n5488 );
xnor g03373 ( new_n5722 , new_n5641 , new_n5675 );
nor  g03374 ( new_n5723 , new_n5721 , new_n5722 );
xnor g03375 ( new_n5724 , new_n5721 , new_n5722 );
xor  g03376 ( new_n5725 , new_n5470 , new_n5486 );
xnor g03377 ( new_n5726 , new_n5647 , new_n5673 );
nor  g03378 ( new_n5727 , new_n5725 , new_n5726 );
xnor g03379 ( new_n5728 , new_n5725 , new_n5726 );
xnor g03380 ( new_n5729 , new_n5652 , new_n5671 );
not  g03381 ( new_n5730 , new_n5729 );
xnor g03382 ( new_n5731 , new_n5473 , new_n5484 );
and  g03383 ( new_n5732_1 , new_n5730 , new_n5731 );
xnor g03384 ( new_n5733 , new_n5730 , new_n5731 );
xnor g03385 ( new_n5734 , new_n5657 , new_n5669 );
xnor g03386 ( new_n5735 , n11302 , n12341 );
xnor g03387 ( new_n5736 , new_n5482 , new_n5735 );
and  g03388 ( new_n5737 , new_n5734 , new_n5736 );
xnor g03389 ( new_n5738 , new_n5734 , new_n5736 );
xnor g03390 ( new_n5739 , new_n5663 , new_n5664 );
xnor g03391 ( new_n5740 , n6773 , n12384 );
nor  g03392 ( new_n5741 , new_n5739 , new_n5740 );
xnor g03393 ( new_n5742_1 , n17090 , n20986 );
xnor g03394 ( new_n5743 , new_n5480 , new_n5742_1 );
nor  g03395 ( new_n5744 , new_n5741 , new_n5743 );
xnor g03396 ( new_n5745 , new_n5665 , new_n5667 );
not  g03397 ( new_n5746 , new_n5745 );
xnor g03398 ( new_n5747 , new_n5741 , new_n5743 );
nor  g03399 ( new_n5748 , new_n5746 , new_n5747 );
nor  g03400 ( new_n5749 , new_n5744 , new_n5748 );
nor  g03401 ( new_n5750 , new_n5738 , new_n5749 );
nor  g03402 ( new_n5751 , new_n5737 , new_n5750 );
nor  g03403 ( new_n5752_1 , new_n5733 , new_n5751 );
nor  g03404 ( new_n5753 , new_n5732_1 , new_n5752_1 );
nor  g03405 ( new_n5754 , new_n5728 , new_n5753 );
nor  g03406 ( new_n5755 , new_n5727 , new_n5754 );
nor  g03407 ( new_n5756 , new_n5724 , new_n5755 );
nor  g03408 ( new_n5757 , new_n5723 , new_n5756 );
nor  g03409 ( new_n5758 , new_n5720 , new_n5757 );
nor  g03410 ( new_n5759 , new_n5719 , new_n5758 );
nor  g03411 ( new_n5760 , new_n5716 , new_n5759 );
nor  g03412 ( new_n5761 , new_n5715 , new_n5760 );
nor  g03413 ( new_n5762 , new_n5712 , new_n5761 );
nor  g03414 ( new_n5763 , new_n5711 , new_n5762 );
nor  g03415 ( new_n5764 , new_n5708 , new_n5763 );
nor  g03416 ( new_n5765_1 , new_n5707 , new_n5764 );
and  g03417 ( new_n5766 , new_n5704_1 , new_n5765_1 );
nor  g03418 ( new_n5767 , new_n5703 , new_n5766 );
xnor g03419 ( n457 , new_n5700_1 , new_n5767 );
xnor g03420 ( new_n5769 , n1681 , n24323 );
xnor g03421 ( new_n5770 , new_n2951 , n13781 );
xnor g03422 ( new_n5771 , new_n5769 , new_n5770 );
not  g03423 ( new_n5772 , new_n5771 );
nor  g03424 ( new_n5773 , new_n5663 , new_n5772 );
xnor g03425 ( new_n5774 , new_n5666 , new_n5773 );
not  g03426 ( new_n5775 , new_n5770 );
nor  g03427 ( new_n5776_1 , new_n5769 , new_n5775 );
nor  g03428 ( new_n5777 , new_n4394 , n24323 );
xnor g03429 ( new_n5778 , n25877 , n26443 );
xnor g03430 ( new_n5779 , new_n5777 , new_n5778 );
xnor g03431 ( new_n5780 , new_n5776_1 , new_n5779 );
xnor g03432 ( new_n5781 , new_n2951 , n9399 );
nor  g03433 ( new_n5782_1 , new_n2951 , new_n2383 );
nor  g03434 ( new_n5783 , n11486 , new_n5782_1 );
not  g03435 ( new_n5784 , n11486 );
or   g03436 ( new_n5785 , new_n5784 , new_n2383 );
nor  g03437 ( new_n5786 , new_n2951 , new_n5785 );
nor  g03438 ( new_n5787 , new_n5783 , new_n5786 );
xnor g03439 ( new_n5788 , new_n5781 , new_n5787 );
not  g03440 ( new_n5789 , new_n5788 );
xnor g03441 ( new_n5790 , new_n5780 , new_n5789 );
xnor g03442 ( n463 , new_n5774 , new_n5790 );
xnor g03443 ( new_n5792 , n6775 , n12121 );
xnor g03444 ( new_n5793 , n8920 , new_n5792 );
not  g03445 ( new_n5794 , new_n5793 );
xnor g03446 ( new_n5795 , n5438 , new_n3063 );
xnor g03447 ( n491 , new_n5794 , new_n5795 );
xnor g03448 ( n496 , new_n5733 , new_n5751 );
not  g03449 ( new_n5798 , n12384 );
xnor g03450 ( new_n5799 , new_n5798 , n25926 );
not  g03451 ( new_n5800 , new_n5799 );
xnor g03452 ( new_n5801 , new_n4030 , new_n5800 );
xnor g03453 ( new_n5802 , n16167 , new_n5663 );
not  g03454 ( new_n5803 , new_n5802 );
nor  g03455 ( new_n5804 , new_n5801 , new_n5803 );
not  g03456 ( new_n5805 , n16167 );
or   g03457 ( new_n5806 , new_n5805 , new_n5663 );
not  g03458 ( new_n5807 , n18745 );
xnor g03459 ( new_n5808 , new_n5807 , new_n5666 );
xor  g03460 ( new_n5809 , new_n5806 , new_n5808 );
nor  g03461 ( new_n5810 , new_n5798 , new_n3982 );
xnor g03462 ( new_n5811 , n7657 , n25926 );
xnor g03463 ( new_n5812 , n20986 , new_n5811 );
xnor g03464 ( new_n5813 , new_n5810 , new_n5812 );
not  g03465 ( new_n5814 , new_n5813 );
or   g03466 ( new_n5815 , new_n4030 , new_n5800 );
nor  g03467 ( new_n5816 , n17090 , new_n5815 );
nor  g03468 ( new_n5817 , n6773 , n17090 );
or   g03469 ( new_n5818 , new_n4030 , new_n4111 );
nor  g03470 ( new_n5819 , new_n5799 , new_n5818 );
or   g03471 ( new_n5820 , new_n5817 , new_n5819 );
nor  g03472 ( new_n5821 , new_n5816 , new_n5820 );
xnor g03473 ( new_n5822_1 , new_n5814 , new_n5821 );
xnor g03474 ( new_n5823 , new_n5809 , new_n5822_1 );
xnor g03475 ( n498 , new_n5804 , new_n5823 );
xnor g03476 ( new_n5825 , new_n4237 , n25872 );
nor  g03477 ( new_n5826 , n20259 , n22043 );
or   g03478 ( new_n5827 , new_n5002 , new_n3875 );
xnor g03479 ( new_n5828 , new_n4939_1 , n22043 );
and  g03480 ( new_n5829 , new_n5827 , new_n5828 );
or   g03481 ( new_n5830 , new_n5826 , new_n5829 );
xor  g03482 ( new_n5831 , new_n5825 , new_n5830 );
xnor g03483 ( new_n5832 , new_n4880 , new_n5831 );
nor  g03484 ( new_n5833_1 , new_n5002 , new_n3875 );
xnor g03485 ( new_n5834_1 , new_n5833_1 , new_n5828 );
nor  g03486 ( new_n5835 , new_n4872 , new_n5834_1 );
xnor g03487 ( new_n5836 , new_n5002 , n12121 );
or   g03488 ( new_n5837 , new_n4874 , new_n5836 );
not  g03489 ( new_n5838 , new_n5834_1 );
xnor g03490 ( new_n5839 , new_n4872 , new_n5838 );
and  g03491 ( new_n5840_1 , new_n5837 , new_n5839 );
nor  g03492 ( new_n5841_1 , new_n5835 , new_n5840_1 );
xnor g03493 ( new_n5842_1 , new_n5832 , new_n5841_1 );
xnor g03494 ( new_n5843 , new_n3792 , new_n5842_1 );
xor  g03495 ( new_n5844 , new_n5837 , new_n5839 );
nor  g03496 ( new_n5845 , new_n3759 , new_n5844 );
not  g03497 ( new_n5846 , new_n3796 );
and  g03498 ( new_n5847 , new_n5846 , new_n5844 );
xnor g03499 ( new_n5848 , new_n4874 , new_n5836 );
and  g03500 ( new_n5849 , new_n3799 , new_n5848 );
nor  g03501 ( new_n5850_1 , new_n5847 , new_n5849 );
nor  g03502 ( new_n5851 , new_n5845 , new_n5850_1 );
xor  g03503 ( n521 , new_n5843 , new_n5851 );
not  g03504 ( new_n5853 , new_n5739 );
xnor g03505 ( n548 , new_n5853 , new_n5740 );
xor  g03506 ( n554 , new_n4289 , new_n4308 );
nor  g03507 ( new_n5856 , n15743 , n20658 );
not  g03508 ( new_n5857 , new_n5856 );
nor  g03509 ( new_n5858 , n7524 , new_n5857 );
not  g03510 ( new_n5859 , new_n5858 );
nor  g03511 ( new_n5860 , n4957 , new_n5859 );
not  g03512 ( new_n5861 , new_n5860 );
nor  g03513 ( new_n5862 , n9003 , new_n5861 );
not  g03514 ( new_n5863 , new_n5862 );
nor  g03515 ( new_n5864 , n3161 , new_n5863 );
not  g03516 ( new_n5865 , new_n5864 );
nor  g03517 ( new_n5866 , n25749 , new_n5865 );
not  g03518 ( new_n5867 , new_n5866 );
nor  g03519 ( new_n5868 , n20409 , new_n5867 );
not  g03520 ( new_n5869 , new_n5868 );
nor  g03521 ( new_n5870 , n647 , new_n5869 );
xnor g03522 ( new_n5871 , n2979 , new_n5870 );
not  g03523 ( new_n5872 , n6456 );
xnor g03524 ( new_n5873 , new_n5872 , n9259 );
nor  g03525 ( new_n5874 , n4085 , n21489 );
not  g03526 ( new_n5875 , n4085 );
xnor g03527 ( new_n5876 , new_n5875 , n21489 );
nor  g03528 ( new_n5877 , n20213 , n26725 );
xnor g03529 ( new_n5878 , new_n4844 , n26725 );
nor  g03530 ( new_n5879 , n11980 , n13912 );
not  g03531 ( new_n5880 , n11980 );
xnor g03532 ( new_n5881 , new_n5880 , n13912 );
nor  g03533 ( new_n5882_1 , n3253 , n7670 );
not  g03534 ( new_n5883 , n3253 );
xnor g03535 ( new_n5884 , new_n5883 , n7670 );
nor  g03536 ( new_n5885 , n7759 , n9598 );
not  g03537 ( new_n5886 , n7759 );
xnor g03538 ( new_n5887 , new_n5886 , n9598 );
nor  g03539 ( new_n5888 , n12562 , n22290 );
not  g03540 ( new_n5889 , n12562 );
xnor g03541 ( new_n5890 , new_n5889 , n22290 );
nor  g03542 ( new_n5891 , n7949 , n11273 );
not  g03543 ( new_n5892 , n7949 );
xnor g03544 ( new_n5893 , new_n5892 , n11273 );
nor  g03545 ( new_n5894 , n24374 , n25565 );
not  g03546 ( new_n5895 , n14575 );
nor  g03547 ( new_n5896 , new_n5895 , new_n3635 );
xnor g03548 ( new_n5897 , n24374 , n25565 );
nor  g03549 ( new_n5898 , new_n5896 , new_n5897 );
or   g03550 ( new_n5899 , new_n5894 , new_n5898 );
and  g03551 ( new_n5900 , new_n5893 , new_n5899 );
or   g03552 ( new_n5901 , new_n5891 , new_n5900 );
and  g03553 ( new_n5902 , new_n5890 , new_n5901 );
or   g03554 ( new_n5903_1 , new_n5888 , new_n5902 );
and  g03555 ( new_n5904_1 , new_n5887 , new_n5903_1 );
or   g03556 ( new_n5905 , new_n5885 , new_n5904_1 );
and  g03557 ( new_n5906 , new_n5884 , new_n5905 );
or   g03558 ( new_n5907 , new_n5882_1 , new_n5906 );
and  g03559 ( new_n5908 , new_n5881 , new_n5907 );
or   g03560 ( new_n5909 , new_n5879 , new_n5908 );
and  g03561 ( new_n5910 , new_n5878 , new_n5909 );
or   g03562 ( new_n5911_1 , new_n5877 , new_n5910 );
and  g03563 ( new_n5912 , new_n5876 , new_n5911_1 );
nor  g03564 ( new_n5913 , new_n5874 , new_n5912 );
xnor g03565 ( new_n5914 , new_n5873 , new_n5913 );
not  g03566 ( new_n5915 , new_n5914 );
xnor g03567 ( new_n5916 , new_n5871 , new_n5915 );
xnor g03568 ( new_n5917 , n647 , new_n5868 );
nor  g03569 ( new_n5918 , new_n5877 , new_n5910 );
xnor g03570 ( new_n5919 , new_n5876 , new_n5918 );
and  g03571 ( new_n5920 , new_n5917 , new_n5919 );
not  g03572 ( new_n5921 , new_n5919 );
xnor g03573 ( new_n5922 , new_n5917 , new_n5921 );
xnor g03574 ( new_n5923 , n20409 , new_n5866 );
nor  g03575 ( new_n5924 , new_n5879 , new_n5908 );
xnor g03576 ( new_n5925 , new_n5878 , new_n5924 );
nor  g03577 ( new_n5926 , new_n5923 , new_n5925 );
xnor g03578 ( new_n5927 , new_n5923 , new_n5925 );
xnor g03579 ( new_n5928 , n25749 , new_n5864 );
nor  g03580 ( new_n5929 , new_n5882_1 , new_n5906 );
xnor g03581 ( new_n5930 , new_n5881 , new_n5929 );
nor  g03582 ( new_n5931 , new_n5928 , new_n5930 );
xnor g03583 ( new_n5932 , new_n5928 , new_n5930 );
xnor g03584 ( new_n5933 , n3161 , new_n5862 );
nor  g03585 ( new_n5934 , new_n5885 , new_n5904_1 );
xnor g03586 ( new_n5935 , new_n5884 , new_n5934 );
nor  g03587 ( new_n5936_1 , new_n5933 , new_n5935 );
xnor g03588 ( new_n5937 , new_n5933 , new_n5935 );
xnor g03589 ( new_n5938 , n9003 , new_n5860 );
nor  g03590 ( new_n5939 , new_n5888 , new_n5902 );
xnor g03591 ( new_n5940 , new_n5887 , new_n5939 );
nor  g03592 ( new_n5941 , new_n5938 , new_n5940 );
xnor g03593 ( new_n5942 , new_n5938 , new_n5940 );
xnor g03594 ( new_n5943_1 , n4957 , new_n5858 );
nor  g03595 ( new_n5944 , new_n5891 , new_n5900 );
xnor g03596 ( new_n5945 , new_n5890 , new_n5944 );
nor  g03597 ( new_n5946 , new_n5943_1 , new_n5945 );
not  g03598 ( new_n5947 , new_n5945 );
xnor g03599 ( new_n5948 , new_n5943_1 , new_n5947 );
xnor g03600 ( new_n5949 , n7524 , new_n5856 );
not  g03601 ( new_n5950 , new_n5949 );
nor  g03602 ( new_n5951 , new_n5894 , new_n5898 );
xnor g03603 ( new_n5952 , new_n5893 , new_n5951 );
not  g03604 ( new_n5953 , new_n5952 );
nor  g03605 ( new_n5954 , new_n5950 , new_n5953 );
xnor g03606 ( new_n5955 , new_n5949 , new_n5953 );
xnor g03607 ( new_n5956 , n14575 , n21993 );
nor  g03608 ( new_n5957 , n20658 , new_n5956 );
and  g03609 ( new_n5958 , new_n3794_1 , new_n5957 );
xnor g03610 ( new_n5959 , new_n5896 , new_n5897 );
xnor g03611 ( new_n5960 , new_n3794_1 , n20658 );
not  g03612 ( new_n5961 , new_n5960 );
nor  g03613 ( new_n5962 , new_n5957 , new_n5961 );
nor  g03614 ( new_n5963 , new_n5958 , new_n5962 );
and  g03615 ( new_n5964_1 , new_n5959 , new_n5963 );
nor  g03616 ( new_n5965 , new_n5958 , new_n5964_1 );
and  g03617 ( new_n5966 , new_n5955 , new_n5965 );
nor  g03618 ( new_n5967 , new_n5954 , new_n5966 );
and  g03619 ( new_n5968 , new_n5948 , new_n5967 );
nor  g03620 ( new_n5969 , new_n5946 , new_n5968 );
nor  g03621 ( new_n5970 , new_n5942 , new_n5969 );
nor  g03622 ( new_n5971 , new_n5941 , new_n5970 );
nor  g03623 ( new_n5972 , new_n5937 , new_n5971 );
nor  g03624 ( new_n5973 , new_n5936_1 , new_n5972 );
nor  g03625 ( new_n5974 , new_n5932 , new_n5973 );
nor  g03626 ( new_n5975 , new_n5931 , new_n5974 );
nor  g03627 ( new_n5976 , new_n5927 , new_n5975 );
nor  g03628 ( new_n5977 , new_n5926 , new_n5976 );
and  g03629 ( new_n5978 , new_n5922 , new_n5977 );
or   g03630 ( new_n5979 , new_n5920 , new_n5978 );
xor  g03631 ( new_n5980_1 , new_n5916 , new_n5979 );
not  g03632 ( new_n5981 , n8526 );
not  g03633 ( new_n5982 , n3582 );
xnor g03634 ( new_n5983 , new_n5982 , n21784 );
nor  g03635 ( new_n5984 , n2145 , n5521 );
not  g03636 ( new_n5985 , n2145 );
xnor g03637 ( new_n5986 , new_n5985 , n5521 );
nor  g03638 ( new_n5987 , n5031 , n11926 );
not  g03639 ( new_n5988 , n5031 );
xnor g03640 ( new_n5989 , new_n5988 , n11926 );
nor  g03641 ( new_n5990 , n4325 , n11044 );
not  g03642 ( new_n5991 , n4325 );
xnor g03643 ( new_n5992 , new_n5991 , n11044 );
nor  g03644 ( new_n5993 , n2421 , n5337 );
not  g03645 ( new_n5994 , n2421 );
xnor g03646 ( new_n5995 , new_n5994 , n5337 );
nor  g03647 ( new_n5996 , n626 , n987 );
xnor g03648 ( new_n5997 , new_n4223 , n987 );
nor  g03649 ( new_n5998 , n1204 , n20478 );
xnor g03650 ( new_n5999 , new_n4233 , n20478 );
nor  g03651 ( new_n6000 , n19618 , n26882 );
xnor g03652 ( new_n6001 , new_n4237 , n26882 );
nor  g03653 ( new_n6002 , n22043 , n22619 );
not  g03654 ( new_n6003 , n6775 );
nor  g03655 ( new_n6004 , new_n6003 , new_n3875 );
xnor g03656 ( new_n6005 , n22043 , n22619 );
nor  g03657 ( new_n6006 , new_n6004 , new_n6005 );
or   g03658 ( new_n6007 , new_n6002 , new_n6006 );
and  g03659 ( new_n6008 , new_n6001 , new_n6007 );
or   g03660 ( new_n6009 , new_n6000 , new_n6008 );
and  g03661 ( new_n6010 , new_n5999 , new_n6009 );
or   g03662 ( new_n6011 , new_n5998 , new_n6010 );
and  g03663 ( new_n6012_1 , new_n5997 , new_n6011 );
or   g03664 ( new_n6013 , new_n5996 , new_n6012_1 );
and  g03665 ( new_n6014 , new_n5995 , new_n6013 );
or   g03666 ( new_n6015 , new_n5993 , new_n6014 );
and  g03667 ( new_n6016 , new_n5992 , new_n6015 );
or   g03668 ( new_n6017 , new_n5990 , new_n6016 );
and  g03669 ( new_n6018 , new_n5989 , new_n6017 );
or   g03670 ( new_n6019 , new_n5987 , new_n6018 );
and  g03671 ( new_n6020 , new_n5986 , new_n6019 );
nor  g03672 ( new_n6021 , new_n5984 , new_n6020 );
xnor g03673 ( new_n6022_1 , new_n5983 , new_n6021 );
not  g03674 ( new_n6023 , new_n6022_1 );
xnor g03675 ( new_n6024 , new_n5981 , new_n6023 );
not  g03676 ( new_n6025 , n2816 );
nor  g03677 ( new_n6026 , new_n5987 , new_n6018 );
xnor g03678 ( new_n6027 , new_n5986 , new_n6026 );
nor  g03679 ( new_n6028 , new_n6025 , new_n6027 );
not  g03680 ( new_n6029 , new_n6027 );
xnor g03681 ( new_n6030 , new_n6025 , new_n6029 );
not  g03682 ( new_n6031_1 , n20359 );
nor  g03683 ( new_n6032 , new_n5990 , new_n6016 );
xnor g03684 ( new_n6033 , new_n5989 , new_n6032 );
nor  g03685 ( new_n6034 , new_n6031_1 , new_n6033 );
not  g03686 ( new_n6035 , new_n6033 );
xnor g03687 ( new_n6036 , new_n6031_1 , new_n6035 );
not  g03688 ( new_n6037 , n4409 );
nor  g03689 ( new_n6038 , new_n5993 , new_n6014 );
xnor g03690 ( new_n6039 , new_n5992 , new_n6038 );
nor  g03691 ( new_n6040 , new_n6037 , new_n6039 );
not  g03692 ( new_n6041 , new_n6039 );
xnor g03693 ( new_n6042 , new_n6037 , new_n6041 );
not  g03694 ( new_n6043 , n3570 );
nor  g03695 ( new_n6044_1 , new_n5996 , new_n6012_1 );
xnor g03696 ( new_n6045 , new_n5995 , new_n6044_1 );
nor  g03697 ( new_n6046_1 , new_n6043 , new_n6045 );
not  g03698 ( new_n6047 , new_n6045 );
xnor g03699 ( new_n6048 , new_n6043 , new_n6047 );
not  g03700 ( new_n6049 , n13668 );
nor  g03701 ( new_n6050 , new_n5998 , new_n6010 );
xnor g03702 ( new_n6051 , new_n5997 , new_n6050 );
nor  g03703 ( new_n6052 , new_n6049 , new_n6051 );
not  g03704 ( new_n6053 , new_n6051 );
xnor g03705 ( new_n6054 , new_n6049 , new_n6053 );
not  g03706 ( new_n6055 , n21276 );
nor  g03707 ( new_n6056 , new_n6000 , new_n6008 );
xnor g03708 ( new_n6057 , new_n5999 , new_n6056 );
nor  g03709 ( new_n6058 , new_n6055 , new_n6057 );
not  g03710 ( new_n6059 , new_n6057 );
xnor g03711 ( new_n6060 , new_n6055 , new_n6059 );
not  g03712 ( new_n6061 , n26748 );
nor  g03713 ( new_n6062 , new_n6002 , new_n6006 );
xnor g03714 ( new_n6063 , new_n6001 , new_n6062 );
nor  g03715 ( new_n6064 , new_n6061 , new_n6063 );
xnor g03716 ( new_n6065 , new_n6004 , new_n6005 );
nor  g03717 ( new_n6066 , n10057 , new_n6065 );
or   g03718 ( new_n6067 , new_n4242 , new_n5792 );
not  g03719 ( new_n6068 , n10057 );
xnor g03720 ( new_n6069 , new_n6068 , new_n6065 );
and  g03721 ( new_n6070 , new_n6067 , new_n6069 );
nor  g03722 ( new_n6071 , new_n6066 , new_n6070 );
not  g03723 ( new_n6072 , new_n6063 );
xnor g03724 ( new_n6073 , new_n6061 , new_n6072 );
and  g03725 ( new_n6074 , new_n6071 , new_n6073 );
or   g03726 ( new_n6075 , new_n6064 , new_n6074 );
and  g03727 ( new_n6076 , new_n6060 , new_n6075 );
or   g03728 ( new_n6077 , new_n6058 , new_n6076 );
and  g03729 ( new_n6078 , new_n6054 , new_n6077 );
or   g03730 ( new_n6079 , new_n6052 , new_n6078 );
and  g03731 ( new_n6080 , new_n6048 , new_n6079 );
or   g03732 ( new_n6081 , new_n6046_1 , new_n6080 );
and  g03733 ( new_n6082 , new_n6042 , new_n6081 );
or   g03734 ( new_n6083 , new_n6040 , new_n6082 );
and  g03735 ( new_n6084_1 , new_n6036 , new_n6083 );
or   g03736 ( new_n6085 , new_n6034 , new_n6084_1 );
and  g03737 ( new_n6086 , new_n6030 , new_n6085 );
nor  g03738 ( new_n6087 , new_n6028 , new_n6086 );
xnor g03739 ( new_n6088 , new_n6024 , new_n6087 );
xnor g03740 ( new_n6089 , new_n5980_1 , new_n6088 );
nor  g03741 ( new_n6090 , new_n6034 , new_n6084_1 );
xnor g03742 ( new_n6091 , new_n6030 , new_n6090 );
xor  g03743 ( new_n6092 , new_n5922 , new_n5977 );
nor  g03744 ( new_n6093 , new_n6091 , new_n6092 );
xnor g03745 ( new_n6094 , new_n6091 , new_n6092 );
xnor g03746 ( new_n6095 , new_n5927 , new_n5975 );
nor  g03747 ( new_n6096 , new_n6040 , new_n6082 );
xnor g03748 ( new_n6097 , new_n6036 , new_n6096 );
nor  g03749 ( new_n6098 , new_n6095 , new_n6097 );
xnor g03750 ( new_n6099 , new_n6095 , new_n6097 );
xnor g03751 ( new_n6100 , new_n5932 , new_n5973 );
nor  g03752 ( new_n6101 , new_n6046_1 , new_n6080 );
xnor g03753 ( new_n6102 , new_n6042 , new_n6101 );
nor  g03754 ( new_n6103 , new_n6100 , new_n6102 );
xnor g03755 ( new_n6104_1 , new_n6100 , new_n6102 );
xnor g03756 ( new_n6105_1 , new_n5937 , new_n5971 );
nor  g03757 ( new_n6106 , new_n6052 , new_n6078 );
xnor g03758 ( new_n6107 , new_n6048 , new_n6106 );
nor  g03759 ( new_n6108 , new_n6105_1 , new_n6107 );
xnor g03760 ( new_n6109 , new_n6105_1 , new_n6107 );
xnor g03761 ( new_n6110 , new_n5942 , new_n5969 );
nor  g03762 ( new_n6111 , new_n6058 , new_n6076 );
xnor g03763 ( new_n6112 , new_n6054 , new_n6111 );
nor  g03764 ( new_n6113 , new_n6110 , new_n6112 );
xnor g03765 ( new_n6114 , new_n6110 , new_n6112 );
xnor g03766 ( new_n6115 , new_n5948 , new_n5967 );
xor  g03767 ( new_n6116 , new_n6060 , new_n6075 );
nor  g03768 ( new_n6117 , new_n6115 , new_n6116 );
xnor g03769 ( new_n6118 , new_n6115 , new_n6116 );
xnor g03770 ( new_n6119 , new_n5955 , new_n5965 );
not  g03771 ( new_n6120 , new_n6119 );
xnor g03772 ( new_n6121 , new_n6071 , new_n6073 );
not  g03773 ( new_n6122 , new_n6121 );
nor  g03774 ( new_n6123 , new_n6120 , new_n6122 );
xnor g03775 ( new_n6124 , new_n6120 , new_n6121 );
nor  g03776 ( new_n6125 , new_n4242 , new_n5792 );
xnor g03777 ( new_n6126 , new_n6125 , new_n6069 );
not  g03778 ( new_n6127 , new_n5959 );
xnor g03779 ( new_n6128 , new_n6127 , new_n5963 );
nor  g03780 ( new_n6129 , new_n6126 , new_n6128 );
xnor g03781 ( new_n6130 , new_n3798 , new_n5956 );
nor  g03782 ( new_n6131 , new_n5794 , new_n6130 );
not  g03783 ( new_n6132 , new_n6126 );
xnor g03784 ( new_n6133 , new_n6132 , new_n6128 );
and  g03785 ( new_n6134 , new_n6131 , new_n6133 );
nor  g03786 ( new_n6135 , new_n6129 , new_n6134 );
and  g03787 ( new_n6136 , new_n6124 , new_n6135 );
nor  g03788 ( new_n6137 , new_n6123 , new_n6136 );
nor  g03789 ( new_n6138 , new_n6118 , new_n6137 );
nor  g03790 ( new_n6139 , new_n6117 , new_n6138 );
nor  g03791 ( new_n6140 , new_n6114 , new_n6139 );
nor  g03792 ( new_n6141 , new_n6113 , new_n6140 );
nor  g03793 ( new_n6142 , new_n6109 , new_n6141 );
nor  g03794 ( new_n6143 , new_n6108 , new_n6142 );
nor  g03795 ( new_n6144 , new_n6104_1 , new_n6143 );
nor  g03796 ( new_n6145 , new_n6103 , new_n6144 );
nor  g03797 ( new_n6146 , new_n6099 , new_n6145 );
nor  g03798 ( new_n6147 , new_n6098 , new_n6146 );
nor  g03799 ( new_n6148 , new_n6094 , new_n6147 );
nor  g03800 ( new_n6149 , new_n6093 , new_n6148 );
xnor g03801 ( n567 , new_n6089 , new_n6149 );
nor  g03802 ( new_n6151 , n1831 , n10250 );
not  g03803 ( new_n6152 , n1831 );
xnor g03804 ( new_n6153 , new_n6152 , n10250 );
nor  g03805 ( new_n6154 , n7674 , n13137 );
not  g03806 ( new_n6155 , n7674 );
xnor g03807 ( new_n6156 , new_n6155 , n13137 );
nor  g03808 ( new_n6157 , n6397 , n18452 );
not  g03809 ( new_n6158 , n6397 );
xnor g03810 ( new_n6159 , new_n6158 , n18452 );
nor  g03811 ( new_n6160_1 , n19196 , n21317 );
not  g03812 ( new_n6161 , n19196 );
xnor g03813 ( new_n6162 , new_n6161 , n21317 );
nor  g03814 ( new_n6163 , n12398 , n23586 );
not  g03815 ( new_n6164 , n12398 );
xnor g03816 ( new_n6165 , new_n6164 , n23586 );
nor  g03817 ( new_n6166 , n19789 , n21226 );
not  g03818 ( new_n6167 , n19789 );
xnor g03819 ( new_n6168 , new_n6167 , n21226 );
nor  g03820 ( new_n6169 , n4426 , n20169 );
not  g03821 ( new_n6170 , n4426 );
xnor g03822 ( new_n6171_1 , new_n6170 , n20169 );
nor  g03823 ( new_n6172 , n8285 , n20036 );
not  g03824 ( new_n6173 , n8285 );
xnor g03825 ( new_n6174 , new_n6173 , n20036 );
nor  g03826 ( new_n6175 , n6729 , n11192 );
not  g03827 ( new_n6176 , n9380 );
or   g03828 ( new_n6177 , new_n6176 , new_n2548 );
not  g03829 ( new_n6178 , n6729 );
xnor g03830 ( new_n6179 , new_n6178 , n11192 );
and  g03831 ( new_n6180 , new_n6177 , new_n6179 );
or   g03832 ( new_n6181 , new_n6175 , new_n6180 );
and  g03833 ( new_n6182 , new_n6174 , new_n6181 );
or   g03834 ( new_n6183_1 , new_n6172 , new_n6182 );
and  g03835 ( new_n6184 , new_n6171_1 , new_n6183_1 );
or   g03836 ( new_n6185 , new_n6169 , new_n6184 );
and  g03837 ( new_n6186 , new_n6168 , new_n6185 );
or   g03838 ( new_n6187 , new_n6166 , new_n6186 );
and  g03839 ( new_n6188 , new_n6165 , new_n6187 );
or   g03840 ( new_n6189_1 , new_n6163 , new_n6188 );
and  g03841 ( new_n6190 , new_n6162 , new_n6189_1 );
or   g03842 ( new_n6191 , new_n6160_1 , new_n6190 );
and  g03843 ( new_n6192 , new_n6159 , new_n6191 );
or   g03844 ( new_n6193 , new_n6157 , new_n6192 );
and  g03845 ( new_n6194 , new_n6156 , new_n6193 );
or   g03846 ( new_n6195 , new_n6154 , new_n6194 );
and  g03847 ( new_n6196 , new_n6153 , new_n6195 );
nor  g03848 ( new_n6197 , new_n6151 , new_n6196 );
not  g03849 ( new_n6198 , n8614 );
not  g03850 ( new_n6199 , new_n4011 );
nor  g03851 ( new_n6200 , n25694 , new_n6199 );
not  g03852 ( new_n6201 , new_n6200 );
nor  g03853 ( new_n6202 , n13110 , new_n6201 );
not  g03854 ( new_n6203 , new_n6202 );
nor  g03855 ( new_n6204_1 , n1752 , new_n6203 );
not  g03856 ( new_n6205 , new_n6204_1 );
nor  g03857 ( new_n6206 , n1288 , new_n6205 );
xnor g03858 ( new_n6207 , n3320 , new_n6206 );
not  g03859 ( new_n6208 , new_n6207 );
nor  g03860 ( new_n6209 , new_n6198 , new_n6208 );
not  g03861 ( new_n6210 , new_n6206 );
nor  g03862 ( new_n6211 , n3320 , new_n6210 );
or   g03863 ( new_n6212 , n8614 , new_n6207 );
xnor g03864 ( new_n6213 , n1288 , new_n6204_1 );
nor  g03865 ( new_n6214 , n15182 , new_n6213 );
not  g03866 ( new_n6215 , n15182 );
not  g03867 ( new_n6216 , new_n6213 );
xnor g03868 ( new_n6217 , new_n6215 , new_n6216 );
xnor g03869 ( new_n6218_1 , n1752 , new_n6202 );
nor  g03870 ( new_n6219 , n27037 , new_n6218_1 );
not  g03871 ( new_n6220 , new_n6218_1 );
xnor g03872 ( new_n6221 , n27037 , new_n6220 );
not  g03873 ( new_n6222 , n8964 );
xnor g03874 ( new_n6223_1 , n13110 , new_n6200 );
not  g03875 ( new_n6224 , new_n6223_1 );
nor  g03876 ( new_n6225 , new_n6222 , new_n6224 );
xnor g03877 ( new_n6226 , n8964 , new_n6224 );
not  g03878 ( new_n6227 , n20151 );
nor  g03879 ( new_n6228 , new_n6227 , new_n4013 );
or   g03880 ( new_n6229 , new_n4018 , new_n4041 );
and  g03881 ( new_n6230 , new_n4014_1 , new_n6229 );
or   g03882 ( new_n6231 , new_n6228 , new_n6230 );
and  g03883 ( new_n6232 , new_n6226 , new_n6231 );
nor  g03884 ( new_n6233_1 , new_n6225 , new_n6232 );
and  g03885 ( new_n6234 , new_n6221 , new_n6233_1 );
nor  g03886 ( new_n6235 , new_n6219 , new_n6234 );
nor  g03887 ( new_n6236 , new_n6217 , new_n6235 );
nor  g03888 ( new_n6237 , new_n6214 , new_n6236 );
and  g03889 ( new_n6238 , new_n6212 , new_n6237 );
or   g03890 ( new_n6239 , new_n6211 , new_n6238 );
nor  g03891 ( new_n6240 , new_n6209 , new_n6239 );
nor  g03892 ( new_n6241 , new_n6197 , new_n6240 );
not  g03893 ( new_n6242 , new_n6197 );
xnor g03894 ( new_n6243 , new_n6242 , new_n6240 );
xor  g03895 ( new_n6244 , new_n6153 , new_n6195 );
xnor g03896 ( new_n6245_1 , n8614 , new_n6208 );
xnor g03897 ( new_n6246 , new_n6237 , new_n6245_1 );
nor  g03898 ( new_n6247 , new_n6244 , new_n6246 );
xnor g03899 ( new_n6248_1 , new_n6217 , new_n6235 );
nor  g03900 ( new_n6249 , new_n6157 , new_n6192 );
xnor g03901 ( new_n6250 , new_n6156 , new_n6249 );
not  g03902 ( new_n6251 , new_n6250 );
nor  g03903 ( new_n6252 , new_n6248_1 , new_n6251 );
xnor g03904 ( new_n6253 , new_n6248_1 , new_n6250 );
xnor g03905 ( new_n6254 , new_n6221 , new_n6233_1 );
nor  g03906 ( new_n6255 , new_n6160_1 , new_n6190 );
xnor g03907 ( new_n6256_1 , new_n6159 , new_n6255 );
not  g03908 ( new_n6257 , new_n6256_1 );
nor  g03909 ( new_n6258 , new_n6254 , new_n6257 );
not  g03910 ( new_n6259 , new_n6254 );
xnor g03911 ( new_n6260 , new_n6259 , new_n6257 );
nor  g03912 ( new_n6261 , new_n6163 , new_n6188 );
xnor g03913 ( new_n6262 , new_n6162 , new_n6261 );
nor  g03914 ( new_n6263 , new_n6228 , new_n6230 );
xnor g03915 ( new_n6264 , new_n6226 , new_n6263 );
not  g03916 ( new_n6265 , new_n6264 );
nor  g03917 ( new_n6266 , new_n6262 , new_n6265 );
nor  g03918 ( new_n6267 , new_n6166 , new_n6186 );
xnor g03919 ( new_n6268 , new_n6165 , new_n6267 );
not  g03920 ( new_n6269 , new_n6268 );
nor  g03921 ( new_n6270 , new_n4043 , new_n6269 );
xnor g03922 ( new_n6271_1 , new_n4044 , new_n6269 );
nor  g03923 ( new_n6272 , new_n6169 , new_n6184 );
xnor g03924 ( new_n6273 , new_n6168 , new_n6272 );
not  g03925 ( new_n6274 , new_n6273 );
nor  g03926 ( new_n6275 , new_n6172 , new_n6182 );
xnor g03927 ( new_n6276_1 , new_n6171_1 , new_n6275 );
not  g03928 ( new_n6277 , new_n6276_1 );
nor  g03929 ( new_n6278 , new_n4052 , new_n6277 );
nor  g03930 ( new_n6279 , new_n6175 , new_n6180 );
xnor g03931 ( new_n6280 , new_n6174 , new_n6279 );
nor  g03932 ( new_n6281 , new_n4057 , new_n6280 );
not  g03933 ( new_n6282 , new_n6280 );
xnor g03934 ( new_n6283 , new_n4058 , new_n6282 );
nor  g03935 ( new_n6284 , new_n6176 , new_n2548 );
xnor g03936 ( new_n6285 , new_n6284 , new_n6179 );
nor  g03937 ( new_n6286 , new_n4064 , new_n6285 );
xnor g03938 ( new_n6287 , new_n6176 , n21687 );
not  g03939 ( new_n6288 , new_n6287 );
nor  g03940 ( new_n6289 , new_n2549 , new_n6288 );
xnor g03941 ( new_n6290 , new_n4067 , new_n6285 );
and  g03942 ( new_n6291 , new_n6289 , new_n6290 );
nor  g03943 ( new_n6292 , new_n6286 , new_n6291 );
nor  g03944 ( new_n6293 , new_n6283 , new_n6292 );
nor  g03945 ( new_n6294 , new_n6281 , new_n6293 );
xnor g03946 ( new_n6295 , new_n4052 , new_n6276_1 );
and  g03947 ( new_n6296 , new_n6294 , new_n6295 );
nor  g03948 ( new_n6297 , new_n6278 , new_n6296 );
nor  g03949 ( new_n6298 , new_n6274 , new_n6297 );
xnor g03950 ( new_n6299 , new_n6273 , new_n6297 );
and  g03951 ( new_n6300 , new_n4049 , new_n6299 );
or   g03952 ( new_n6301 , new_n6298 , new_n6300 );
and  g03953 ( new_n6302 , new_n6271_1 , new_n6301 );
nor  g03954 ( new_n6303 , new_n6270 , new_n6302 );
not  g03955 ( new_n6304 , new_n6262 );
xnor g03956 ( new_n6305 , new_n6304 , new_n6265 );
and  g03957 ( new_n6306 , new_n6303 , new_n6305 );
nor  g03958 ( new_n6307 , new_n6266 , new_n6306 );
and  g03959 ( new_n6308_1 , new_n6260 , new_n6307 );
or   g03960 ( new_n6309 , new_n6258 , new_n6308_1 );
and  g03961 ( new_n6310 , new_n6253 , new_n6309 );
nor  g03962 ( new_n6311_1 , new_n6252 , new_n6310 );
not  g03963 ( new_n6312 , new_n6246 );
xnor g03964 ( new_n6313 , new_n6244 , new_n6312 );
and  g03965 ( new_n6314 , new_n6311_1 , new_n6313 );
nor  g03966 ( new_n6315 , new_n6247 , new_n6314 );
and  g03967 ( new_n6316 , new_n6243 , new_n6315 );
nor  g03968 ( new_n6317 , new_n6241 , new_n6316 );
xnor g03969 ( new_n6318 , new_n6243 , new_n6315 );
nor  g03970 ( new_n6319 , n6105 , n15766 );
not  g03971 ( new_n6320 , n15766 );
xnor g03972 ( new_n6321 , n6105 , new_n6320 );
nor  g03973 ( new_n6322 , n3795 , n25629 );
not  g03974 ( new_n6323_1 , n3795 );
xnor g03975 ( new_n6324 , new_n6323_1 , n25629 );
nor  g03976 ( new_n6325 , n7692 , n25464 );
not  g03977 ( new_n6326 , n7692 );
xnor g03978 ( new_n6327 , new_n6326 , n25464 );
nor  g03979 ( new_n6328 , n4590 , n23039 );
not  g03980 ( new_n6329 , n23039 );
xnor g03981 ( new_n6330_1 , n4590 , new_n6329 );
nor  g03982 ( new_n6331 , n13677 , n26752 );
xnor g03983 ( new_n6332 , n13677 , n26752 );
nor  g03984 ( new_n6333 , n6513 , n18926 );
not  g03985 ( new_n6334 , n6513 );
xnor g03986 ( new_n6335 , new_n6334 , n18926 );
not  g03987 ( new_n6336 , n3918 );
nor  g03988 ( new_n6337 , new_n6336 , new_n3967 );
or   g03989 ( new_n6338 , n3918 , n5451 );
nor  g03990 ( new_n6339_1 , n919 , n5330 );
or   g03991 ( new_n6340 , new_n4145 , new_n4149 );
and  g03992 ( new_n6341 , new_n4144 , new_n6340 );
nor  g03993 ( new_n6342 , new_n6339_1 , new_n6341 );
and  g03994 ( new_n6343 , new_n6338 , new_n6342 );
nor  g03995 ( new_n6344 , new_n6337 , new_n6343 );
and  g03996 ( new_n6345 , new_n6335 , new_n6344 );
nor  g03997 ( new_n6346 , new_n6333 , new_n6345 );
nor  g03998 ( new_n6347 , new_n6332 , new_n6346 );
or   g03999 ( new_n6348 , new_n6331 , new_n6347 );
and  g04000 ( new_n6349 , new_n6330_1 , new_n6348 );
or   g04001 ( new_n6350 , new_n6328 , new_n6349 );
and  g04002 ( new_n6351 , new_n6327 , new_n6350 );
or   g04003 ( new_n6352 , new_n6325 , new_n6351 );
and  g04004 ( new_n6353 , new_n6324 , new_n6352 );
or   g04005 ( new_n6354_1 , new_n6322 , new_n6353 );
and  g04006 ( new_n6355 , new_n6321 , new_n6354_1 );
nor  g04007 ( new_n6356_1 , new_n6319 , new_n6355 );
not  g04008 ( new_n6357 , new_n6356_1 );
nor  g04009 ( new_n6358 , new_n6318 , new_n6357 );
xnor g04010 ( new_n6359 , new_n6318 , new_n6357 );
nor  g04011 ( new_n6360 , new_n6322 , new_n6353 );
xnor g04012 ( new_n6361 , new_n6321 , new_n6360 );
not  g04013 ( new_n6362 , new_n6361 );
xnor g04014 ( new_n6363 , new_n6311_1 , new_n6313 );
and  g04015 ( new_n6364 , new_n6362 , new_n6363 );
xnor g04016 ( new_n6365 , new_n6362 , new_n6363 );
xor  g04017 ( new_n6366 , new_n6253 , new_n6309 );
xor  g04018 ( new_n6367 , new_n6324 , new_n6352 );
not  g04019 ( new_n6368 , new_n6367 );
and  g04020 ( new_n6369_1 , new_n6366 , new_n6368 );
xnor g04021 ( new_n6370 , new_n6366 , new_n6368 );
xnor g04022 ( new_n6371 , new_n6260 , new_n6307 );
nor  g04023 ( new_n6372 , new_n6328 , new_n6349 );
xnor g04024 ( new_n6373 , new_n6327 , new_n6372 );
nor  g04025 ( new_n6374 , new_n6371 , new_n6373 );
xnor g04026 ( new_n6375_1 , new_n6371 , new_n6373 );
xor  g04027 ( new_n6376 , new_n6330_1 , new_n6348 );
not  g04028 ( new_n6377 , new_n6376 );
xnor g04029 ( new_n6378 , new_n6303 , new_n6305 );
and  g04030 ( new_n6379_1 , new_n6377 , new_n6378 );
xnor g04031 ( new_n6380 , new_n6377 , new_n6378 );
xor  g04032 ( new_n6381_1 , new_n6271_1 , new_n6301 );
xnor g04033 ( new_n6382 , new_n6332 , new_n6346 );
and  g04034 ( new_n6383_1 , new_n6381_1 , new_n6382 );
xnor g04035 ( new_n6384 , new_n6381_1 , new_n6382 );
xnor g04036 ( new_n6385_1 , new_n4049 , new_n6299 );
xor  g04037 ( new_n6386 , new_n6335 , new_n6344 );
nor  g04038 ( new_n6387 , new_n6385_1 , new_n6386 );
xnor g04039 ( new_n6388 , new_n6385_1 , new_n6386 );
xnor g04040 ( new_n6389 , new_n6294 , new_n6295 );
xnor g04041 ( new_n6390 , new_n6336 , n5451 );
xnor g04042 ( new_n6391 , new_n6342 , new_n6390 );
nor  g04043 ( new_n6392 , new_n6389 , new_n6391 );
xnor g04044 ( new_n6393 , new_n6389 , new_n6391 );
not  g04045 ( new_n6394 , new_n4151_1 );
xnor g04046 ( new_n6395 , new_n6283 , new_n6292 );
and  g04047 ( new_n6396 , new_n6394 , new_n6395 );
xnor g04048 ( new_n6397_1 , new_n6394 , new_n6395 );
xnor g04049 ( new_n6398 , new_n6289 , new_n6290 );
not  g04050 ( new_n6399 , new_n6398 );
nor  g04051 ( new_n6400 , new_n4155 , new_n6399 );
xnor g04052 ( new_n6401 , new_n2549 , new_n6287 );
nor  g04053 ( new_n6402 , new_n4157 , new_n6401 );
xnor g04054 ( new_n6403 , new_n4160 , new_n6399 );
and  g04055 ( new_n6404 , new_n6402 , new_n6403 );
nor  g04056 ( new_n6405 , new_n6400 , new_n6404 );
nor  g04057 ( new_n6406 , new_n6397_1 , new_n6405 );
nor  g04058 ( new_n6407_1 , new_n6396 , new_n6406 );
nor  g04059 ( new_n6408 , new_n6393 , new_n6407_1 );
nor  g04060 ( new_n6409 , new_n6392 , new_n6408 );
nor  g04061 ( new_n6410 , new_n6388 , new_n6409 );
nor  g04062 ( new_n6411 , new_n6387 , new_n6410 );
nor  g04063 ( new_n6412 , new_n6384 , new_n6411 );
nor  g04064 ( new_n6413 , new_n6383_1 , new_n6412 );
nor  g04065 ( new_n6414 , new_n6380 , new_n6413 );
nor  g04066 ( new_n6415 , new_n6379_1 , new_n6414 );
nor  g04067 ( new_n6416 , new_n6375_1 , new_n6415 );
nor  g04068 ( new_n6417 , new_n6374 , new_n6416 );
nor  g04069 ( new_n6418 , new_n6370 , new_n6417 );
nor  g04070 ( new_n6419 , new_n6369_1 , new_n6418 );
nor  g04071 ( new_n6420 , new_n6365 , new_n6419 );
nor  g04072 ( new_n6421 , new_n6364 , new_n6420 );
nor  g04073 ( new_n6422 , new_n6359 , new_n6421 );
nor  g04074 ( new_n6423 , new_n6358 , new_n6422 );
nor  g04075 ( n588 , new_n6317 , new_n6423 );
xnor g04076 ( new_n6425 , n18584 , n19803 );
not  g04077 ( new_n6426 , n12626 );
nor  g04078 ( new_n6427_1 , n4272 , new_n6426 );
and  g04079 ( new_n6428 , new_n4661 , new_n4684 );
nor  g04080 ( new_n6429 , new_n6427_1 , new_n6428 );
xnor g04081 ( new_n6430 , new_n6425 , new_n6429 );
not  g04082 ( new_n6431_1 , new_n6430 );
xnor g04083 ( new_n6432 , n7773 , n16911 );
not  g04084 ( new_n6433 , n376 );
nor  g04085 ( new_n6434 , new_n6433 , n7721 );
xnor g04086 ( new_n6435 , n376 , n7721 );
not  g04087 ( new_n6436 , n5517 );
nor  g04088 ( new_n6437_1 , new_n6436 , n21981 );
xnor g04089 ( new_n6438 , n5517 , n21981 );
not  g04090 ( new_n6439 , n12113 );
nor  g04091 ( new_n6440 , new_n6439 , n12917 );
xnor g04092 ( new_n6441 , n12113 , n12917 );
not  g04093 ( new_n6442 , n10614 );
and  g04094 ( new_n6443 , new_n6442 , n21898 );
nor  g04095 ( new_n6444 , new_n6442 , n21898 );
not  g04096 ( new_n6445 , n11266 );
and  g04097 ( new_n6446 , n9926 , new_n6445 );
nor  g04098 ( new_n6447 , n9926 , new_n6445 );
not  g04099 ( new_n6448 , n22072 );
nor  g04100 ( new_n6449 , n2646 , new_n6448 );
not  g04101 ( new_n6450 , new_n6449 );
nor  g04102 ( new_n6451 , new_n6447 , new_n6450 );
nor  g04103 ( new_n6452 , new_n6446 , new_n6451 );
nor  g04104 ( new_n6453 , new_n6444 , new_n6452 );
nor  g04105 ( new_n6454 , new_n6443 , new_n6453 );
and  g04106 ( new_n6455 , new_n6441 , new_n6454 );
or   g04107 ( new_n6456_1 , new_n6440 , new_n6455 );
and  g04108 ( new_n6457_1 , new_n6438 , new_n6456_1 );
or   g04109 ( new_n6458 , new_n6437_1 , new_n6457_1 );
and  g04110 ( new_n6459 , new_n6435 , new_n6458 );
or   g04111 ( new_n6460 , new_n6434 , new_n6459 );
xor  g04112 ( new_n6461 , new_n6432 , new_n6460 );
nor  g04113 ( new_n6462 , n4939 , n15652 );
not  g04114 ( new_n6463 , new_n6462 );
nor  g04115 ( new_n6464 , n5605 , new_n6463 );
not  g04116 ( new_n6465_1 , new_n6464 );
nor  g04117 ( new_n6466 , n2985 , new_n6465_1 );
not  g04118 ( new_n6467 , new_n6466 );
nor  g04119 ( new_n6468 , n14576 , new_n6467 );
not  g04120 ( new_n6469 , new_n6468 );
nor  g04121 ( new_n6470_1 , n1269 , new_n6469 );
xnor g04122 ( new_n6471 , n16818 , new_n6470_1 );
not  g04123 ( new_n6472 , new_n6471 );
xnor g04124 ( new_n6473 , n1742 , new_n6472 );
xnor g04125 ( new_n6474 , n1269 , new_n6468 );
nor  g04126 ( new_n6475 , n4858 , new_n6474 );
not  g04127 ( new_n6476_1 , new_n6474 );
xnor g04128 ( new_n6477 , n4858 , new_n6476_1 );
xnor g04129 ( new_n6478 , n14576 , new_n6466 );
nor  g04130 ( new_n6479 , n8244 , new_n6478 );
not  g04131 ( new_n6480 , new_n6478 );
xnor g04132 ( new_n6481 , n8244 , new_n6480 );
xnor g04133 ( new_n6482 , n2985 , new_n6464 );
nor  g04134 ( new_n6483 , n9493 , new_n6482 );
xnor g04135 ( new_n6484 , n5605 , new_n6462 );
nor  g04136 ( new_n6485_1 , n15167 , new_n6484 );
not  g04137 ( new_n6486 , new_n6484 );
xnor g04138 ( new_n6487 , n15167 , new_n6486 );
xnor g04139 ( new_n6488 , n4939 , n15652 );
not  g04140 ( new_n6489 , new_n6488 );
nor  g04141 ( new_n6490 , n21095 , new_n6489 );
not  g04142 ( new_n6491 , n4939 );
not  g04143 ( new_n6492 , n8656 );
or   g04144 ( new_n6493 , new_n6491 , new_n6492 );
xnor g04145 ( new_n6494 , n21095 , new_n6488 );
and  g04146 ( new_n6495 , new_n6493 , new_n6494 );
or   g04147 ( new_n6496 , new_n6490 , new_n6495 );
and  g04148 ( new_n6497 , new_n6487 , new_n6496 );
or   g04149 ( new_n6498 , new_n6485_1 , new_n6497 );
not  g04150 ( new_n6499 , new_n6482 );
xnor g04151 ( new_n6500 , n9493 , new_n6499 );
and  g04152 ( new_n6501 , new_n6498 , new_n6500 );
or   g04153 ( new_n6502_1 , new_n6483 , new_n6501 );
and  g04154 ( new_n6503 , new_n6481 , new_n6502_1 );
or   g04155 ( new_n6504 , new_n6479 , new_n6503 );
and  g04156 ( new_n6505 , new_n6477 , new_n6504 );
nor  g04157 ( new_n6506_1 , new_n6475 , new_n6505 );
xnor g04158 ( new_n6507 , new_n6473 , new_n6506_1 );
not  g04159 ( new_n6508 , new_n6507 );
xnor g04160 ( new_n6509 , new_n6461 , new_n6508 );
xor  g04161 ( new_n6510 , new_n6435 , new_n6458 );
not  g04162 ( new_n6511 , new_n6510 );
nor  g04163 ( new_n6512 , new_n6479 , new_n6503 );
xnor g04164 ( new_n6513_1 , new_n6477 , new_n6512 );
nor  g04165 ( new_n6514_1 , new_n6511 , new_n6513_1 );
xnor g04166 ( new_n6515 , new_n6510 , new_n6513_1 );
xnor g04167 ( new_n6516 , new_n6438 , new_n6456_1 );
nor  g04168 ( new_n6517 , new_n6483 , new_n6501 );
xnor g04169 ( new_n6518 , new_n6481 , new_n6517 );
and  g04170 ( new_n6519 , new_n6516 , new_n6518 );
xor  g04171 ( new_n6520 , new_n6438 , new_n6456_1 );
xnor g04172 ( new_n6521 , new_n6520 , new_n6518 );
xnor g04173 ( new_n6522 , new_n6441 , new_n6454 );
nor  g04174 ( new_n6523 , new_n6485_1 , new_n6497 );
xnor g04175 ( new_n6524 , new_n6523 , new_n6500 );
nor  g04176 ( new_n6525 , new_n6522 , new_n6524 );
xor  g04177 ( new_n6526 , new_n6487 , new_n6496 );
xnor g04178 ( new_n6527 , n10614 , n21898 );
xnor g04179 ( new_n6528 , new_n6452 , new_n6527 );
and  g04180 ( new_n6529 , new_n6526 , new_n6528 );
xnor g04181 ( new_n6530 , new_n6526 , new_n6528 );
xnor g04182 ( new_n6531 , n4939 , n8656 );
xnor g04183 ( new_n6532 , n2646 , n22072 );
nor  g04184 ( new_n6533 , new_n6531 , new_n6532 );
xnor g04185 ( new_n6534 , n9926 , n11266 );
xnor g04186 ( new_n6535 , new_n6450 , new_n6534 );
not  g04187 ( new_n6536 , new_n6535 );
nor  g04188 ( new_n6537 , new_n6533 , new_n6536 );
xor  g04189 ( new_n6538 , new_n6493 , new_n6494 );
xnor g04190 ( new_n6539 , new_n6533 , new_n6535 );
and  g04191 ( new_n6540 , new_n6538 , new_n6539 );
nor  g04192 ( new_n6541 , new_n6537 , new_n6540 );
nor  g04193 ( new_n6542_1 , new_n6530 , new_n6541 );
nor  g04194 ( new_n6543 , new_n6529 , new_n6542_1 );
xor  g04195 ( new_n6544 , new_n6522 , new_n6524 );
and  g04196 ( new_n6545 , new_n6543 , new_n6544 );
nor  g04197 ( new_n6546 , new_n6525 , new_n6545 );
and  g04198 ( new_n6547 , new_n6521 , new_n6546 );
nor  g04199 ( new_n6548 , new_n6519 , new_n6547 );
and  g04200 ( new_n6549 , new_n6515 , new_n6548 );
nor  g04201 ( new_n6550 , new_n6514_1 , new_n6549 );
xnor g04202 ( new_n6551 , new_n6509 , new_n6550 );
not  g04203 ( new_n6552 , new_n6551 );
xnor g04204 ( new_n6553 , new_n6431_1 , new_n6552 );
xor  g04205 ( new_n6554 , new_n6515 , new_n6548 );
nor  g04206 ( new_n6555 , new_n4685 , new_n6554 );
xnor g04207 ( new_n6556_1 , new_n4685 , new_n6554 );
xnor g04208 ( new_n6557 , new_n6521 , new_n6546 );
nor  g04209 ( new_n6558_1 , new_n4688 , new_n6557 );
xnor g04210 ( new_n6559 , new_n4688 , new_n6557 );
xnor g04211 ( new_n6560_1 , new_n6543 , new_n6544 );
not  g04212 ( new_n6561 , new_n6560_1 );
nor  g04213 ( new_n6562 , new_n4694 , new_n6561 );
xnor g04214 ( new_n6563 , new_n4694 , new_n6561 );
xnor g04215 ( new_n6564 , new_n6530 , new_n6541 );
nor  g04216 ( new_n6565 , new_n4702 , new_n6564 );
not  g04217 ( new_n6566 , new_n6564 );
xnor g04218 ( new_n6567_1 , new_n4701 , new_n6566 );
xnor g04219 ( new_n6568 , new_n6531 , new_n6532 );
or   g04220 ( new_n6569 , new_n4711 , new_n6568 );
and  g04221 ( new_n6570 , new_n4708 , new_n6569 );
xnor g04222 ( new_n6571 , new_n6538 , new_n6539 );
not  g04223 ( new_n6572 , new_n6571 );
xor  g04224 ( new_n6573 , new_n4708 , new_n6569 );
and  g04225 ( new_n6574 , new_n6572 , new_n6573 );
nor  g04226 ( new_n6575 , new_n6570 , new_n6574 );
nor  g04227 ( new_n6576_1 , new_n6567_1 , new_n6575 );
nor  g04228 ( new_n6577 , new_n6565 , new_n6576_1 );
nor  g04229 ( new_n6578 , new_n6563 , new_n6577 );
nor  g04230 ( new_n6579 , new_n6562 , new_n6578 );
nor  g04231 ( new_n6580 , new_n6559 , new_n6579 );
nor  g04232 ( new_n6581 , new_n6558_1 , new_n6580 );
nor  g04233 ( new_n6582 , new_n6556_1 , new_n6581 );
nor  g04234 ( new_n6583 , new_n6555 , new_n6582 );
xor  g04235 ( n597 , new_n6553 , new_n6583 );
not  g04236 ( new_n6585 , n9646 );
xnor g04237 ( new_n6586 , new_n6585 , n25926 );
xnor g04238 ( new_n6587_1 , n14230 , new_n6586 );
xnor g04239 ( n637 , new_n5802 , new_n6587_1 );
not  g04240 ( new_n6589 , n7421 );
not  g04241 ( new_n6590_1 , n10611 );
xnor g04242 ( new_n6591 , new_n6590_1 , n25797 );
nor  g04243 ( new_n6592 , n2783 , n15967 );
not  g04244 ( new_n6593 , n2783 );
xnor g04245 ( new_n6594 , new_n6593 , n15967 );
nor  g04246 ( new_n6595 , n13319 , n15490 );
not  g04247 ( new_n6596_1 , n18 );
nor  g04248 ( new_n6597 , new_n6596_1 , new_n3756 );
xnor g04249 ( new_n6598 , n13319 , n15490 );
nor  g04250 ( new_n6599 , new_n6597 , new_n6598 );
or   g04251 ( new_n6600 , new_n6595 , new_n6599 );
and  g04252 ( new_n6601 , new_n6594 , new_n6600 );
nor  g04253 ( new_n6602 , new_n6592 , new_n6601 );
xnor g04254 ( new_n6603 , new_n6591 , new_n6602 );
not  g04255 ( new_n6604 , new_n6603 );
xnor g04256 ( new_n6605 , new_n6589 , new_n6604 );
not  g04257 ( new_n6606 , n19680 );
nor  g04258 ( new_n6607 , new_n6595 , new_n6599 );
xnor g04259 ( new_n6608 , new_n6594 , new_n6607 );
nor  g04260 ( new_n6609 , new_n6606 , new_n6608 );
not  g04261 ( new_n6610 , new_n6608 );
xnor g04262 ( new_n6611_1 , new_n6606 , new_n6610 );
xnor g04263 ( new_n6612_1 , new_n6597 , new_n6598 );
nor  g04264 ( new_n6613 , n2809 , new_n6612_1 );
xnor g04265 ( new_n6614 , n18 , n25435 );
or   g04266 ( new_n6615 , new_n4818 , new_n6614 );
not  g04267 ( new_n6616 , n2809 );
xnor g04268 ( new_n6617 , new_n6616 , new_n6612_1 );
and  g04269 ( new_n6618 , new_n6615 , new_n6617 );
nor  g04270 ( new_n6619 , new_n6613 , new_n6618 );
and  g04271 ( new_n6620 , new_n6611_1 , new_n6619 );
or   g04272 ( new_n6621 , new_n6609 , new_n6620 );
xor  g04273 ( new_n6622 , new_n6605 , new_n6621 );
not  g04274 ( new_n6623 , new_n6622 );
xnor g04275 ( new_n6624 , n11056 , n18157 );
nor  g04276 ( new_n6625 , n12161 , n15271 );
xnor g04277 ( new_n6626 , n12161 , n15271 );
nor  g04278 ( new_n6627 , n5026 , n25877 );
not  g04279 ( new_n6628_1 , n8581 );
not  g04280 ( new_n6629 , n24323 );
nor  g04281 ( new_n6630_1 , new_n6628_1 , new_n6629 );
xnor g04282 ( new_n6631_1 , n5026 , n25877 );
nor  g04283 ( new_n6632 , new_n6630_1 , new_n6631_1 );
nor  g04284 ( new_n6633 , new_n6627 , new_n6632 );
nor  g04285 ( new_n6634_1 , new_n6626 , new_n6633 );
nor  g04286 ( new_n6635 , new_n6625 , new_n6634_1 );
xnor g04287 ( new_n6636 , new_n6624 , new_n6635 );
xnor g04288 ( new_n6637 , n20250 , new_n6636 );
xnor g04289 ( new_n6638 , new_n6626 , new_n6633 );
nor  g04290 ( new_n6639 , n5822 , new_n6638 );
xnor g04291 ( new_n6640 , new_n6630_1 , new_n6631_1 );
nor  g04292 ( new_n6641 , n26443 , new_n6640 );
xnor g04293 ( new_n6642 , n8581 , n24323 );
or   g04294 ( new_n6643 , new_n4394 , new_n6642 );
not  g04295 ( new_n6644 , n26443 );
xnor g04296 ( new_n6645 , new_n6644 , new_n6640 );
and  g04297 ( new_n6646 , new_n6643 , new_n6645 );
or   g04298 ( new_n6647 , new_n6641 , new_n6646 );
xnor g04299 ( new_n6648 , new_n4384 , new_n6638 );
and  g04300 ( new_n6649 , new_n6647 , new_n6648 );
nor  g04301 ( new_n6650 , new_n6639 , new_n6649 );
xnor g04302 ( new_n6651 , new_n6637 , new_n6650 );
not  g04303 ( new_n6652_1 , new_n6651 );
xnor g04304 ( new_n6653 , new_n6623 , new_n6652_1 );
xnor g04305 ( new_n6654 , new_n6611_1 , new_n6619 );
xnor g04306 ( new_n6655_1 , new_n6647 , new_n6648 );
and  g04307 ( new_n6656 , new_n6654 , new_n6655_1 );
xor  g04308 ( new_n6657 , new_n6647 , new_n6648 );
xnor g04309 ( new_n6658 , new_n6654 , new_n6657 );
nor  g04310 ( new_n6659_1 , new_n4818 , new_n6614 );
xnor g04311 ( new_n6660 , new_n6659_1 , new_n6617 );
nor  g04312 ( new_n6661 , new_n4394 , new_n6642 );
xnor g04313 ( new_n6662 , new_n6661 , new_n6645 );
not  g04314 ( new_n6663 , new_n6662 );
nor  g04315 ( new_n6664 , new_n6660 , new_n6663 );
xnor g04316 ( new_n6665 , new_n4818 , new_n6614 );
xnor g04317 ( new_n6666 , n1681 , new_n6642 );
nor  g04318 ( new_n6667 , new_n6665 , new_n6666 );
not  g04319 ( new_n6668 , new_n6660 );
xnor g04320 ( new_n6669_1 , new_n6668 , new_n6663 );
and  g04321 ( new_n6670 , new_n6667 , new_n6669_1 );
nor  g04322 ( new_n6671_1 , new_n6664 , new_n6670 );
and  g04323 ( new_n6672 , new_n6658 , new_n6671_1 );
nor  g04324 ( new_n6673_1 , new_n6656 , new_n6672 );
xnor g04325 ( n646 , new_n6653 , new_n6673_1 );
nor  g04326 ( new_n6675 , n2387 , n19494 );
not  g04327 ( new_n6676 , new_n6675 );
nor  g04328 ( new_n6677 , n16223 , new_n6676 );
not  g04329 ( new_n6678 , new_n6677 );
nor  g04330 ( new_n6679 , n26913 , new_n6678 );
xnor g04331 ( new_n6680 , n21832 , new_n6679 );
xnor g04332 ( new_n6681 , new_n5468 , new_n2466 );
nor  g04333 ( new_n6682 , new_n5471 , new_n2470 );
xnor g04334 ( new_n6683 , new_n5471 , new_n2470 );
nor  g04335 ( new_n6684_1 , new_n5475 , new_n2473 );
xnor g04336 ( new_n6685 , n12341 , new_n2475 );
nor  g04337 ( new_n6686 , n12384 , new_n2478 );
and  g04338 ( new_n6687 , new_n5478 , new_n6686 );
xor  g04339 ( new_n6688 , new_n2449 , new_n2480 );
xnor g04340 ( new_n6689 , new_n5478 , new_n6686 );
nor  g04341 ( new_n6690 , new_n6688 , new_n6689 );
or   g04342 ( new_n6691_1 , new_n6687 , new_n6690 );
nor  g04343 ( new_n6692 , new_n6685 , new_n6691_1 );
nor  g04344 ( new_n6693 , new_n6684_1 , new_n6692 );
nor  g04345 ( new_n6694 , new_n6683 , new_n6693 );
nor  g04346 ( new_n6695 , new_n6682 , new_n6694 );
xor  g04347 ( new_n6696 , new_n6681 , new_n6695 );
xnor g04348 ( new_n6697 , new_n6680 , new_n6696 );
xnor g04349 ( new_n6698 , n26913 , new_n6677 );
xor  g04350 ( new_n6699 , new_n6683 , new_n6693 );
and  g04351 ( new_n6700 , new_n6698 , new_n6699 );
xnor g04352 ( new_n6701 , new_n6698 , new_n6699 );
xnor g04353 ( new_n6702 , new_n5798 , new_n2478 );
nor  g04354 ( new_n6703 , new_n3116 , new_n6702 );
and  g04355 ( new_n6704 , new_n2365 , new_n6703 );
xnor g04356 ( new_n6705 , new_n2481 , new_n6689 );
xnor g04357 ( new_n6706_1 , new_n3116 , n19494 );
nor  g04358 ( new_n6707_1 , new_n6703 , new_n6706_1 );
or   g04359 ( new_n6708 , new_n6704 , new_n6707_1 );
nor  g04360 ( new_n6709 , new_n6705 , new_n6708 );
nor  g04361 ( new_n6710 , new_n6704 , new_n6709 );
xnor g04362 ( new_n6711 , n16223 , new_n6675 );
not  g04363 ( new_n6712 , new_n6711 );
nor  g04364 ( new_n6713 , new_n6710 , new_n6712 );
xnor g04365 ( new_n6714 , new_n6685 , new_n6691_1 );
not  g04366 ( new_n6715 , new_n6714 );
xnor g04367 ( new_n6716 , new_n6710 , new_n6711 );
and  g04368 ( new_n6717 , new_n6715 , new_n6716 );
nor  g04369 ( new_n6718 , new_n6713 , new_n6717 );
nor  g04370 ( new_n6719 , new_n6701 , new_n6718 );
nor  g04371 ( new_n6720 , new_n6700 , new_n6719 );
xor  g04372 ( new_n6721 , new_n6697 , new_n6720 );
xnor g04373 ( new_n6722 , new_n3354 , new_n6721 );
xor  g04374 ( new_n6723 , new_n6701 , new_n6718 );
nor  g04375 ( new_n6724 , new_n3358 , new_n6723 );
xnor g04376 ( new_n6725 , new_n6714 , new_n6716 );
and  g04377 ( new_n6726 , new_n3364 , new_n6725 );
xnor g04378 ( new_n6727 , new_n3363 , new_n6725 );
xnor g04379 ( new_n6728 , n2387 , new_n6702 );
and  g04380 ( new_n6729_1 , new_n3367 , new_n6728 );
nor  g04381 ( new_n6730 , new_n3370 , new_n6729_1 );
not  g04382 ( new_n6731 , new_n6705 );
xnor g04383 ( new_n6732 , new_n6731 , new_n6708 );
not  g04384 ( new_n6733 , new_n6732 );
and  g04385 ( new_n6734 , new_n3308 , new_n6729_1 );
nor  g04386 ( new_n6735 , new_n6730 , new_n6734 );
and  g04387 ( new_n6736_1 , new_n6733 , new_n6735 );
nor  g04388 ( new_n6737 , new_n6730 , new_n6736_1 );
and  g04389 ( new_n6738 , new_n6727 , new_n6737 );
or   g04390 ( new_n6739 , new_n6726 , new_n6738 );
xnor g04391 ( new_n6740 , new_n3358 , new_n6723 );
nor  g04392 ( new_n6741 , new_n6739 , new_n6740 );
nor  g04393 ( new_n6742 , new_n6724 , new_n6741 );
xnor g04394 ( n696 , new_n6722 , new_n6742 );
not  g04395 ( new_n6744 , n23697 );
xnor g04396 ( new_n6745 , new_n6744 , n25475 );
not  g04397 ( new_n6746 , new_n6745 );
nor  g04398 ( new_n6747 , n2289 , n23849 );
not  g04399 ( new_n6748 , n2289 );
xnor g04400 ( new_n6749 , new_n6748 , n23849 );
not  g04401 ( new_n6750 , new_n6749 );
nor  g04402 ( new_n6751 , n1112 , n12446 );
not  g04403 ( new_n6752 , n1112 );
xnor g04404 ( new_n6753 , new_n6752 , n12446 );
not  g04405 ( new_n6754 , new_n6753 );
nor  g04406 ( new_n6755 , n11011 , n20179 );
not  g04407 ( new_n6756 , n20179 );
xnor g04408 ( new_n6757 , n11011 , new_n6756 );
not  g04409 ( new_n6758 , new_n6757 );
nor  g04410 ( new_n6759 , n16029 , n19228 );
xnor g04411 ( new_n6760 , new_n3939 , n19228 );
not  g04412 ( new_n6761 , new_n6760 );
nor  g04413 ( new_n6762 , n15539 , n16476 );
not  g04414 ( new_n6763 , n15539 );
xnor g04415 ( new_n6764 , new_n6763 , n16476 );
not  g04416 ( new_n6765 , new_n6764 );
nor  g04417 ( new_n6766 , n8052 , n11615 );
not  g04418 ( new_n6767 , n8052 );
xnor g04419 ( new_n6768 , new_n6767 , n11615 );
not  g04420 ( new_n6769 , new_n6768 );
nor  g04421 ( new_n6770 , n10158 , n22433 );
not  g04422 ( new_n6771 , n18962 );
nor  g04423 ( new_n6772 , new_n3952_1 , new_n6771 );
xnor g04424 ( new_n6773_1 , n10158 , n22433 );
nor  g04425 ( new_n6774 , new_n6772 , new_n6773_1 );
nor  g04426 ( new_n6775_1 , new_n6770 , new_n6774 );
nor  g04427 ( new_n6776 , new_n6769 , new_n6775_1 );
nor  g04428 ( new_n6777 , new_n6766 , new_n6776 );
nor  g04429 ( new_n6778 , new_n6765 , new_n6777 );
nor  g04430 ( new_n6779 , new_n6762 , new_n6778 );
nor  g04431 ( new_n6780 , new_n6761 , new_n6779 );
nor  g04432 ( new_n6781 , new_n6759 , new_n6780 );
nor  g04433 ( new_n6782 , new_n6758 , new_n6781 );
nor  g04434 ( new_n6783 , new_n6755 , new_n6782 );
nor  g04435 ( new_n6784 , new_n6754 , new_n6783 );
nor  g04436 ( new_n6785_1 , new_n6751 , new_n6784 );
nor  g04437 ( new_n6786 , new_n6750 , new_n6785_1 );
nor  g04438 ( new_n6787 , new_n6747 , new_n6786 );
xnor g04439 ( new_n6788 , new_n6746 , new_n6787 );
not  g04440 ( new_n6789 , new_n6788 );
xnor g04441 ( new_n6790_1 , new_n5503 , new_n6789 );
xnor g04442 ( new_n6791_1 , new_n6750 , new_n6785_1 );
and  g04443 ( new_n6792 , n9655 , new_n6791_1 );
xnor g04444 ( new_n6793 , n9655 , new_n6791_1 );
xnor g04445 ( new_n6794_1 , new_n6754 , new_n6783 );
and  g04446 ( new_n6795 , n13490 , new_n6794_1 );
xnor g04447 ( new_n6796 , n13490 , new_n6794_1 );
xnor g04448 ( new_n6797 , new_n6758 , new_n6781 );
not  g04449 ( new_n6798 , new_n6797 );
nor  g04450 ( new_n6799 , new_n5511 , new_n6798 );
xnor g04451 ( new_n6800 , new_n6761 , new_n6779 );
nor  g04452 ( new_n6801 , n1777 , new_n6800 );
not  g04453 ( new_n6802_1 , new_n6800 );
xnor g04454 ( new_n6803 , new_n5514 , new_n6802_1 );
xnor g04455 ( new_n6804 , new_n6765 , new_n6777 );
nor  g04456 ( new_n6805 , n8745 , new_n6804 );
not  g04457 ( new_n6806 , new_n6804 );
xnor g04458 ( new_n6807 , new_n5517_1 , new_n6806 );
xnor g04459 ( new_n6808 , new_n6769 , new_n6775_1 );
not  g04460 ( new_n6809 , new_n6808 );
nor  g04461 ( new_n6810 , new_n2441 , new_n6809 );
xnor g04462 ( new_n6811 , n15636 , new_n6809 );
xnor g04463 ( new_n6812 , n14090 , n18962 );
nor  g04464 ( new_n6813 , new_n2447 , new_n6812 );
nor  g04465 ( new_n6814_1 , n20077 , new_n6813 );
xor  g04466 ( new_n6815 , new_n6772 , new_n6773_1 );
xnor g04467 ( new_n6816 , new_n2444_1 , new_n6813 );
and  g04468 ( new_n6817 , new_n6815 , new_n6816 );
nor  g04469 ( new_n6818 , new_n6814_1 , new_n6817 );
and  g04470 ( new_n6819 , new_n6811 , new_n6818 );
nor  g04471 ( new_n6820 , new_n6810 , new_n6819 );
not  g04472 ( new_n6821 , new_n6820 );
nor  g04473 ( new_n6822 , new_n6807 , new_n6821 );
nor  g04474 ( new_n6823 , new_n6805 , new_n6822 );
nor  g04475 ( new_n6824 , new_n6803 , new_n6823 );
or   g04476 ( new_n6825 , new_n6801 , new_n6824 );
xnor g04477 ( new_n6826_1 , new_n5511 , new_n6798 );
nor  g04478 ( new_n6827 , new_n6825 , new_n6826_1 );
nor  g04479 ( new_n6828 , new_n6799 , new_n6827 );
nor  g04480 ( new_n6829 , new_n6796 , new_n6828 );
nor  g04481 ( new_n6830 , new_n6795 , new_n6829 );
nor  g04482 ( new_n6831 , new_n6793 , new_n6830 );
nor  g04483 ( new_n6832 , new_n6792 , new_n6831 );
xnor g04484 ( new_n6833 , new_n6790_1 , new_n6832 );
xnor g04485 ( new_n6834 , new_n6215 , n21915 );
nor  g04486 ( new_n6835_1 , n13775 , n27037 );
not  g04487 ( new_n6836 , n13775 );
xnor g04488 ( new_n6837 , new_n6836 , n27037 );
nor  g04489 ( new_n6838 , n1293 , n8964 );
not  g04490 ( new_n6839 , n1293 );
xnor g04491 ( new_n6840 , new_n6839 , n8964 );
nor  g04492 ( new_n6841 , n19042 , n20151 );
not  g04493 ( new_n6842 , n19042 );
xnor g04494 ( new_n6843 , new_n6842 , n20151 );
nor  g04495 ( new_n6844 , n7693 , n19472 );
xnor g04496 ( new_n6845 , new_n4015 , n19472 );
not  g04497 ( new_n6846 , n25370 );
nor  g04498 ( new_n6847 , new_n4021 , new_n6846 );
or   g04499 ( new_n6848 , n10405 , n25370 );
nor  g04500 ( new_n6849 , n11302 , n24786 );
or   g04501 ( new_n6850 , new_n4108 , new_n4113 );
and  g04502 ( new_n6851 , new_n4107 , new_n6850 );
nor  g04503 ( new_n6852 , new_n6849 , new_n6851 );
and  g04504 ( new_n6853_1 , new_n6848 , new_n6852 );
nor  g04505 ( new_n6854 , new_n6847 , new_n6853_1 );
and  g04506 ( new_n6855 , new_n6845 , new_n6854 );
or   g04507 ( new_n6856 , new_n6844 , new_n6855 );
and  g04508 ( new_n6857 , new_n6843 , new_n6856 );
or   g04509 ( new_n6858 , new_n6841 , new_n6857 );
and  g04510 ( new_n6859 , new_n6840 , new_n6858 );
or   g04511 ( new_n6860 , new_n6838 , new_n6859 );
and  g04512 ( new_n6861_1 , new_n6837 , new_n6860 );
nor  g04513 ( new_n6862_1 , new_n6835_1 , new_n6861_1 );
xnor g04514 ( new_n6863_1 , new_n6834 , new_n6862_1 );
not  g04515 ( new_n6864 , new_n6863_1 );
xnor g04516 ( new_n6865 , new_n5456 , new_n6864 );
nor  g04517 ( new_n6866 , new_n6838 , new_n6859 );
xnor g04518 ( new_n6867_1 , new_n6837 , new_n6866 );
nor  g04519 ( new_n6868 , new_n5459 , new_n6867_1 );
not  g04520 ( new_n6869 , new_n6867_1 );
xnor g04521 ( new_n6870 , new_n5459 , new_n6869 );
nor  g04522 ( new_n6871 , new_n6841 , new_n6857 );
xnor g04523 ( new_n6872 , new_n6840 , new_n6871 );
nor  g04524 ( new_n6873 , new_n5462 , new_n6872 );
not  g04525 ( new_n6874 , new_n6872 );
xnor g04526 ( new_n6875 , new_n5462 , new_n6874 );
nor  g04527 ( new_n6876 , new_n6844 , new_n6855 );
xnor g04528 ( new_n6877 , new_n6843 , new_n6876 );
nor  g04529 ( new_n6878 , new_n5465 , new_n6877 );
not  g04530 ( new_n6879 , new_n6877 );
xnor g04531 ( new_n6880 , new_n5465 , new_n6879 );
xnor g04532 ( new_n6881 , new_n6845 , new_n6854 );
not  g04533 ( new_n6882 , new_n6881 );
nor  g04534 ( new_n6883 , new_n5468 , new_n6882 );
xnor g04535 ( new_n6884 , n7566 , new_n6882 );
xnor g04536 ( new_n6885 , new_n4021 , n25370 );
xnor g04537 ( new_n6886 , new_n6852 , new_n6885 );
nor  g04538 ( new_n6887 , new_n5471 , new_n6886 );
not  g04539 ( new_n6888 , new_n6886 );
xnor g04540 ( new_n6889 , new_n5471 , new_n6888 );
nor  g04541 ( new_n6890 , new_n5475 , new_n4115 );
nor  g04542 ( new_n6891 , n20986 , new_n4138 );
or   g04543 ( new_n6892 , new_n5798 , new_n4135 );
xnor g04544 ( new_n6893 , new_n5478 , new_n4138 );
and  g04545 ( new_n6894 , new_n6892 , new_n6893 );
nor  g04546 ( new_n6895 , new_n6891 , new_n6894 );
xnor g04547 ( new_n6896 , new_n5475 , new_n4116 );
and  g04548 ( new_n6897 , new_n6895 , new_n6896 );
or   g04549 ( new_n6898 , new_n6890 , new_n6897 );
and  g04550 ( new_n6899 , new_n6889 , new_n6898 );
or   g04551 ( new_n6900 , new_n6887 , new_n6899 );
and  g04552 ( new_n6901 , new_n6884 , new_n6900 );
or   g04553 ( new_n6902 , new_n6883 , new_n6901 );
and  g04554 ( new_n6903 , new_n6880 , new_n6902 );
or   g04555 ( new_n6904 , new_n6878 , new_n6903 );
and  g04556 ( new_n6905 , new_n6875 , new_n6904 );
or   g04557 ( new_n6906 , new_n6873 , new_n6905 );
and  g04558 ( new_n6907 , new_n6870 , new_n6906 );
or   g04559 ( new_n6908 , new_n6868 , new_n6907 );
xor  g04560 ( new_n6909 , new_n6865 , new_n6908 );
xnor g04561 ( new_n6910 , new_n6833 , new_n6909 );
xor  g04562 ( new_n6911 , new_n6870 , new_n6906 );
not  g04563 ( new_n6912 , new_n6911 );
xor  g04564 ( new_n6913 , new_n6793 , new_n6830 );
and  g04565 ( new_n6914 , new_n6912 , new_n6913 );
xnor g04566 ( new_n6915 , new_n6912 , new_n6913 );
xor  g04567 ( new_n6916 , new_n6875 , new_n6904 );
not  g04568 ( new_n6917 , new_n6916 );
xor  g04569 ( new_n6918 , new_n6796 , new_n6828 );
and  g04570 ( new_n6919 , new_n6917 , new_n6918 );
xnor g04571 ( new_n6920 , new_n6917 , new_n6918 );
xor  g04572 ( new_n6921 , new_n6880 , new_n6902 );
not  g04573 ( new_n6922 , new_n6921 );
xor  g04574 ( new_n6923 , new_n6825 , new_n6826_1 );
and  g04575 ( new_n6924 , new_n6922 , new_n6923 );
xnor g04576 ( new_n6925 , new_n6922 , new_n6923 );
xnor g04577 ( new_n6926 , new_n6803 , new_n6823 );
not  g04578 ( new_n6927 , new_n6926 );
xor  g04579 ( new_n6928 , new_n6884 , new_n6900 );
nor  g04580 ( new_n6929 , new_n6927 , new_n6928 );
xnor g04581 ( new_n6930 , new_n6927 , new_n6928 );
xnor g04582 ( new_n6931 , new_n6807 , new_n6820 );
xor  g04583 ( new_n6932 , new_n6889 , new_n6898 );
nor  g04584 ( new_n6933 , new_n6931 , new_n6932 );
xnor g04585 ( new_n6934 , new_n6931 , new_n6932 );
xnor g04586 ( new_n6935 , new_n6895 , new_n6896 );
xnor g04587 ( new_n6936 , new_n6811 , new_n6818 );
not  g04588 ( new_n6937 , new_n6936 );
and  g04589 ( new_n6938 , new_n6935 , new_n6937 );
xnor g04590 ( new_n6939 , new_n6935 , new_n6937 );
nor  g04591 ( new_n6940 , new_n5798 , new_n4135 );
xnor g04592 ( new_n6941 , new_n6940 , new_n6893 );
xnor g04593 ( new_n6942 , new_n6772 , new_n6773_1 );
xnor g04594 ( new_n6943 , new_n6942 , new_n6816 );
not  g04595 ( new_n6944 , new_n6943 );
and  g04596 ( new_n6945 , new_n6941 , new_n6944 );
xnor g04597 ( new_n6946 , n6794 , new_n6812 );
not  g04598 ( new_n6947 , new_n6946 );
xnor g04599 ( new_n6948 , n12384 , new_n4135 );
nor  g04600 ( new_n6949 , new_n6947 , new_n6948 );
xnor g04601 ( new_n6950 , new_n6941 , new_n6943 );
and  g04602 ( new_n6951 , new_n6949 , new_n6950 );
nor  g04603 ( new_n6952 , new_n6945 , new_n6951 );
nor  g04604 ( new_n6953 , new_n6939 , new_n6952 );
nor  g04605 ( new_n6954 , new_n6938 , new_n6953 );
nor  g04606 ( new_n6955 , new_n6934 , new_n6954 );
nor  g04607 ( new_n6956 , new_n6933 , new_n6955 );
nor  g04608 ( new_n6957 , new_n6930 , new_n6956 );
nor  g04609 ( new_n6958 , new_n6929 , new_n6957 );
nor  g04610 ( new_n6959 , new_n6925 , new_n6958 );
nor  g04611 ( new_n6960 , new_n6924 , new_n6959 );
nor  g04612 ( new_n6961 , new_n6920 , new_n6960 );
nor  g04613 ( new_n6962 , new_n6919 , new_n6961 );
nor  g04614 ( new_n6963 , new_n6915 , new_n6962 );
nor  g04615 ( new_n6964 , new_n6914 , new_n6963 );
xnor g04616 ( n723 , new_n6910 , new_n6964 );
xnor g04617 ( new_n6966 , n2272 , n26986 );
not  g04618 ( new_n6967_1 , n25331 );
nor  g04619 ( new_n6968 , n21287 , new_n6967_1 );
xnor g04620 ( new_n6969 , n21287 , n25331 );
not  g04621 ( new_n6970 , n18483 );
nor  g04622 ( new_n6971_1 , n4256 , new_n6970 );
xnor g04623 ( new_n6972 , n4256 , n18483 );
not  g04624 ( new_n6973 , n21934 );
nor  g04625 ( new_n6974 , new_n6973 , n22332 );
xnor g04626 ( new_n6975_1 , n21934 , n22332 );
not  g04627 ( new_n6976 , n18901 );
nor  g04628 ( new_n6977 , new_n6976 , n18907 );
xnor g04629 ( new_n6978 , n18901 , n18907 );
not  g04630 ( new_n6979 , n4376 );
nor  g04631 ( new_n6980 , n2731 , new_n6979 );
xnor g04632 ( new_n6981 , n2731 , n4376 );
not  g04633 ( new_n6982 , n14570 );
nor  g04634 ( new_n6983_1 , new_n6982 , n19911 );
xnor g04635 ( new_n6984 , n14570 , n19911 );
nor  g04636 ( new_n6985_1 , new_n2389 , n23775 );
not  g04637 ( new_n6986 , n23775 );
nor  g04638 ( new_n6987 , n13708 , new_n6986 );
nor  g04639 ( new_n6988 , n8259 , new_n3826 );
not  g04640 ( new_n6989 , n8259 );
nor  g04641 ( new_n6990 , new_n6989 , n18409 );
nor  g04642 ( new_n6991 , new_n2381 , n11479 );
not  g04643 ( new_n6992 , new_n6991 );
nor  g04644 ( new_n6993 , new_n6990 , new_n6992 );
nor  g04645 ( new_n6994 , new_n6988 , new_n6993 );
nor  g04646 ( new_n6995 , new_n6987 , new_n6994 );
nor  g04647 ( new_n6996 , new_n6985_1 , new_n6995 );
and  g04648 ( new_n6997 , new_n6984 , new_n6996 );
or   g04649 ( new_n6998_1 , new_n6983_1 , new_n6997 );
and  g04650 ( new_n6999 , new_n6981 , new_n6998_1 );
or   g04651 ( new_n7000 , new_n6980 , new_n6999 );
and  g04652 ( new_n7001 , new_n6978 , new_n7000 );
or   g04653 ( new_n7002 , new_n6977 , new_n7001 );
and  g04654 ( new_n7003 , new_n6975_1 , new_n7002 );
or   g04655 ( new_n7004 , new_n6974 , new_n7003 );
and  g04656 ( new_n7005 , new_n6972 , new_n7004 );
or   g04657 ( new_n7006 , new_n6971_1 , new_n7005 );
and  g04658 ( new_n7007 , new_n6969 , new_n7006 );
or   g04659 ( new_n7008 , new_n6968 , new_n7007 );
xor  g04660 ( new_n7009 , new_n6966 , new_n7008 );
xnor g04661 ( new_n7010 , n468 , n1255 );
nor  g04662 ( new_n7011 , n5400 , n9512 );
xnor g04663 ( new_n7012 , n5400 , n9512 );
nor  g04664 ( new_n7013 , n16608 , n23923 );
xnor g04665 ( new_n7014 , n16608 , n23923 );
nor  g04666 ( new_n7015 , n329 , n21735 );
xnor g04667 ( new_n7016 , n329 , n21735 );
nor  g04668 ( new_n7017 , n24085 , n24170 );
xnor g04669 ( new_n7018 , n24085 , n24170 );
nor  g04670 ( new_n7019 , n2409 , n14071 );
xnor g04671 ( new_n7020 , n2409 , n14071 );
nor  g04672 ( new_n7021 , n1738 , n8869 );
xnor g04673 ( new_n7022 , n1738 , n8869 );
nor  g04674 ( new_n7023 , n10372 , n12152 );
not  g04675 ( new_n7024 , n7428 );
not  g04676 ( new_n7025 , n19107 );
nor  g04677 ( new_n7026_1 , new_n7024 , new_n7025 );
xnor g04678 ( new_n7027 , n10372 , n12152 );
nor  g04679 ( new_n7028 , new_n7026_1 , new_n7027 );
nor  g04680 ( new_n7029 , new_n7023 , new_n7028 );
nor  g04681 ( new_n7030 , new_n7022 , new_n7029 );
nor  g04682 ( new_n7031 , new_n7021 , new_n7030 );
nor  g04683 ( new_n7032_1 , new_n7020 , new_n7031 );
nor  g04684 ( new_n7033 , new_n7019 , new_n7032_1 );
nor  g04685 ( new_n7034 , new_n7018 , new_n7033 );
nor  g04686 ( new_n7035 , new_n7017 , new_n7034 );
nor  g04687 ( new_n7036 , new_n7016 , new_n7035 );
nor  g04688 ( new_n7037 , new_n7015 , new_n7036 );
nor  g04689 ( new_n7038_1 , new_n7014 , new_n7037 );
nor  g04690 ( new_n7039 , new_n7013 , new_n7038_1 );
nor  g04691 ( new_n7040 , new_n7012 , new_n7039 );
nor  g04692 ( new_n7041 , new_n7011 , new_n7040 );
xnor g04693 ( new_n7042 , new_n7010 , new_n7041 );
not  g04694 ( new_n7043 , n12861 );
xnor g04695 ( new_n7044 , new_n7043 , n14130 );
nor  g04696 ( new_n7045 , n13333 , n16482 );
not  g04697 ( new_n7046 , n13333 );
xnor g04698 ( new_n7047 , new_n7046 , n16482 );
nor  g04699 ( new_n7048 , n2210 , n9942 );
not  g04700 ( new_n7049 , n2210 );
xnor g04701 ( new_n7050 , new_n7049 , n9942 );
nor  g04702 ( new_n7051 , n20604 , n25643 );
or   g04703 ( new_n7052 , new_n5127 , new_n5129 );
and  g04704 ( new_n7053 , new_n5126 , new_n7052 );
or   g04705 ( new_n7054 , new_n7051 , new_n7053 );
and  g04706 ( new_n7055 , new_n7050 , new_n7054 );
or   g04707 ( new_n7056 , new_n7048 , new_n7055 );
and  g04708 ( new_n7057_1 , new_n7047 , new_n7056 );
nor  g04709 ( new_n7058 , new_n7045 , new_n7057_1 );
xnor g04710 ( new_n7059 , new_n7044 , new_n7058 );
nor  g04711 ( new_n7060 , new_n7042 , new_n7059 );
xnor g04712 ( new_n7061 , new_n7042 , new_n7059 );
xnor g04713 ( new_n7062 , new_n7012 , new_n7039 );
nor  g04714 ( new_n7063 , new_n7048 , new_n7055 );
xnor g04715 ( new_n7064 , new_n7047 , new_n7063 );
nor  g04716 ( new_n7065 , new_n7062 , new_n7064 );
xnor g04717 ( new_n7066 , new_n7062 , new_n7064 );
nor  g04718 ( new_n7067 , new_n7051 , new_n7053 );
xnor g04719 ( new_n7068 , new_n7050 , new_n7067 );
xnor g04720 ( new_n7069 , new_n7014 , new_n7037 );
nor  g04721 ( new_n7070 , new_n7068 , new_n7069 );
xnor g04722 ( new_n7071 , new_n7068 , new_n7069 );
xnor g04723 ( new_n7072 , new_n7016 , new_n7035 );
nor  g04724 ( new_n7073 , new_n5131_1 , new_n7072 );
xnor g04725 ( new_n7074 , new_n5131_1 , new_n7072 );
xnor g04726 ( new_n7075 , new_n7018 , new_n7033 );
nor  g04727 ( new_n7076 , new_n5122 , new_n7075 );
xnor g04728 ( new_n7077 , new_n5122 , new_n7075 );
xnor g04729 ( new_n7078 , new_n7020 , new_n7031 );
nor  g04730 ( new_n7079_1 , new_n5112 , new_n7078 );
xnor g04731 ( new_n7080 , new_n5113 , new_n7078 );
xnor g04732 ( new_n7081 , new_n7022 , new_n7029 );
nor  g04733 ( new_n7082 , new_n5102 , new_n7081 );
xnor g04734 ( new_n7083 , new_n5102 , new_n7081 );
xnor g04735 ( new_n7084 , new_n7026_1 , new_n7027 );
nor  g04736 ( new_n7085 , new_n5093 , new_n7084 );
xnor g04737 ( new_n7086 , new_n7024 , n19107 );
nor  g04738 ( new_n7087 , new_n5143 , new_n7086 );
xnor g04739 ( new_n7088 , new_n5094 , new_n7084 );
and  g04740 ( new_n7089 , new_n7087 , new_n7088 );
nor  g04741 ( new_n7090 , new_n7085 , new_n7089 );
nor  g04742 ( new_n7091 , new_n7083 , new_n7090 );
or   g04743 ( new_n7092 , new_n7082 , new_n7091 );
and  g04744 ( new_n7093 , new_n7080 , new_n7092 );
nor  g04745 ( new_n7094 , new_n7079_1 , new_n7093 );
nor  g04746 ( new_n7095 , new_n7077 , new_n7094 );
nor  g04747 ( new_n7096 , new_n7076 , new_n7095 );
nor  g04748 ( new_n7097 , new_n7074 , new_n7096 );
nor  g04749 ( new_n7098 , new_n7073 , new_n7097 );
nor  g04750 ( new_n7099_1 , new_n7071 , new_n7098 );
nor  g04751 ( new_n7100 , new_n7070 , new_n7099_1 );
nor  g04752 ( new_n7101 , new_n7066 , new_n7100 );
nor  g04753 ( new_n7102 , new_n7065 , new_n7101 );
nor  g04754 ( new_n7103 , new_n7061 , new_n7102 );
nor  g04755 ( new_n7104 , new_n7060 , new_n7103 );
xnor g04756 ( new_n7105 , n22253 , n22442 );
nor  g04757 ( new_n7106 , n468 , n1255 );
nor  g04758 ( new_n7107 , new_n7010 , new_n7041 );
nor  g04759 ( new_n7108 , new_n7106 , new_n7107 );
xnor g04760 ( new_n7109 , new_n7105 , new_n7108 );
not  g04761 ( new_n7110 , n8305 );
xnor g04762 ( new_n7111 , new_n7110 , n8856 );
nor  g04763 ( new_n7112 , n12861 , n14130 );
or   g04764 ( new_n7113 , new_n7045 , new_n7057_1 );
and  g04765 ( new_n7114 , new_n7044 , new_n7113 );
nor  g04766 ( new_n7115 , new_n7112 , new_n7114 );
xnor g04767 ( new_n7116 , new_n7111 , new_n7115 );
xnor g04768 ( new_n7117 , new_n7109 , new_n7116 );
xnor g04769 ( new_n7118 , new_n7104 , new_n7117 );
nor  g04770 ( new_n7119 , new_n7009 , new_n7118 );
xnor g04771 ( new_n7120 , new_n7009 , new_n7118 );
xor  g04772 ( new_n7121 , new_n6969 , new_n7006 );
xnor g04773 ( new_n7122 , new_n7061 , new_n7102 );
nor  g04774 ( new_n7123 , new_n7121 , new_n7122 );
xnor g04775 ( new_n7124 , new_n7121 , new_n7122 );
xor  g04776 ( new_n7125 , new_n6972 , new_n7004 );
xnor g04777 ( new_n7126 , new_n7066 , new_n7100 );
nor  g04778 ( new_n7127 , new_n7125 , new_n7126 );
xnor g04779 ( new_n7128 , new_n7125 , new_n7126 );
xor  g04780 ( new_n7129 , new_n6975_1 , new_n7002 );
xnor g04781 ( new_n7130 , new_n7071 , new_n7098 );
nor  g04782 ( new_n7131 , new_n7129 , new_n7130 );
xnor g04783 ( new_n7132 , new_n7129 , new_n7130 );
xor  g04784 ( new_n7133 , new_n6978 , new_n7000 );
xnor g04785 ( new_n7134 , new_n7074 , new_n7096 );
nor  g04786 ( new_n7135 , new_n7133 , new_n7134 );
xnor g04787 ( new_n7136 , new_n7133 , new_n7134 );
xor  g04788 ( new_n7137 , new_n6981 , new_n6998_1 );
xnor g04789 ( new_n7138 , new_n7077 , new_n7094 );
nor  g04790 ( new_n7139_1 , new_n7137 , new_n7138 );
xnor g04791 ( new_n7140 , new_n7137 , new_n7138 );
xor  g04792 ( new_n7141 , new_n7080 , new_n7092 );
xnor g04793 ( new_n7142 , new_n6984 , new_n6996 );
and  g04794 ( new_n7143 , new_n7141 , new_n7142 );
xnor g04795 ( new_n7144 , new_n7083 , new_n7090 );
not  g04796 ( new_n7145 , new_n7144 );
xnor g04797 ( new_n7146 , n13708 , n23775 );
xnor g04798 ( new_n7147 , new_n6994 , new_n7146 );
and  g04799 ( new_n7148 , new_n7145 , new_n7147 );
xnor g04800 ( new_n7149_1 , new_n7144 , new_n7147 );
xnor g04801 ( new_n7150 , new_n5090 , new_n7086 );
xnor g04802 ( new_n7151 , n5704 , n11479 );
nor  g04803 ( new_n7152 , new_n7150 , new_n7151 );
xnor g04804 ( new_n7153 , n8259 , n18409 );
xnor g04805 ( new_n7154 , new_n6992 , new_n7153 );
not  g04806 ( new_n7155 , new_n7154 );
and  g04807 ( new_n7156 , new_n7152 , new_n7155 );
xnor g04808 ( new_n7157 , new_n7087 , new_n7088 );
not  g04809 ( new_n7158 , new_n7157 );
xnor g04810 ( new_n7159 , new_n7152 , new_n7155 );
nor  g04811 ( new_n7160 , new_n7158 , new_n7159 );
nor  g04812 ( new_n7161 , new_n7156 , new_n7160 );
and  g04813 ( new_n7162 , new_n7149_1 , new_n7161 );
nor  g04814 ( new_n7163 , new_n7148 , new_n7162 );
xnor g04815 ( new_n7164 , new_n7141 , new_n7142 );
nor  g04816 ( new_n7165 , new_n7163 , new_n7164 );
nor  g04817 ( new_n7166 , new_n7143 , new_n7165 );
nor  g04818 ( new_n7167 , new_n7140 , new_n7166 );
nor  g04819 ( new_n7168 , new_n7139_1 , new_n7167 );
nor  g04820 ( new_n7169 , new_n7136 , new_n7168 );
nor  g04821 ( new_n7170 , new_n7135 , new_n7169 );
nor  g04822 ( new_n7171 , new_n7132 , new_n7170 );
nor  g04823 ( new_n7172 , new_n7131 , new_n7171 );
nor  g04824 ( new_n7173 , new_n7128 , new_n7172 );
nor  g04825 ( new_n7174 , new_n7127 , new_n7173 );
nor  g04826 ( new_n7175 , new_n7124 , new_n7174 );
nor  g04827 ( new_n7176 , new_n7123 , new_n7175 );
nor  g04828 ( new_n7177 , new_n7120 , new_n7176 );
nor  g04829 ( new_n7178 , new_n7119 , new_n7177 );
not  g04830 ( new_n7179 , n2272 );
nor  g04831 ( new_n7180 , new_n7179 , n26986 );
and  g04832 ( new_n7181 , new_n6966 , new_n7008 );
nor  g04833 ( new_n7182 , new_n7180 , new_n7181 );
nor  g04834 ( new_n7183 , n22253 , n22442 );
nor  g04835 ( new_n7184 , new_n7105 , new_n7108 );
nor  g04836 ( new_n7185 , new_n7183 , new_n7184 );
nor  g04837 ( new_n7186 , n8305 , n8856 );
or   g04838 ( new_n7187 , new_n7112 , new_n7114 );
and  g04839 ( new_n7188 , new_n7111 , new_n7187 );
nor  g04840 ( new_n7189 , new_n7186 , new_n7188 );
xnor g04841 ( new_n7190_1 , new_n7185 , new_n7189 );
nor  g04842 ( new_n7191 , new_n7109 , new_n7116 );
nor  g04843 ( new_n7192 , new_n7104 , new_n7117 );
nor  g04844 ( new_n7193 , new_n7191 , new_n7192 );
xnor g04845 ( new_n7194 , new_n7190_1 , new_n7193 );
not  g04846 ( new_n7195 , new_n7194 );
xnor g04847 ( new_n7196 , new_n7182 , new_n7195 );
xnor g04848 ( n735 , new_n7178 , new_n7196 );
xnor g04849 ( new_n7198 , n14230 , n21138 );
xnor g04850 ( new_n7199 , n19234 , new_n6812 );
not  g04851 ( new_n7200 , new_n7199 );
xnor g04852 ( new_n7201 , n26167 , new_n7200 );
xnor g04853 ( n779 , new_n7198 , new_n7201 );
nor  g04854 ( new_n7203 , new_n5981 , n17458 );
xnor g04855 ( new_n7204 , n8526 , n17458 );
nor  g04856 ( new_n7205 , n1222 , new_n6025 );
xnor g04857 ( new_n7206 , n1222 , n2816 );
nor  g04858 ( new_n7207 , new_n6031_1 , n25240 );
xnor g04859 ( new_n7208 , n20359 , n25240 );
nor  g04860 ( new_n7209 , new_n6037 , n10125 );
xnor g04861 ( new_n7210 , n4409 , n10125 );
nor  g04862 ( new_n7211 , new_n6043 , n8067 );
xnor g04863 ( new_n7212 , n3570 , n8067 );
nor  g04864 ( new_n7213 , new_n6049 , n20923 );
xnor g04865 ( new_n7214 , n13668 , n20923 );
nor  g04866 ( new_n7215 , n18157 , new_n6055 );
xnor g04867 ( new_n7216 , n18157 , n21276 );
not  g04868 ( new_n7217 , n12161 );
nor  g04869 ( new_n7218 , new_n7217 , n26748 );
nor  g04870 ( new_n7219 , n12161 , new_n6061 );
not  g04871 ( new_n7220 , n5026 );
nor  g04872 ( new_n7221 , new_n7220 , n10057 );
nor  g04873 ( new_n7222 , n5026 , new_n6068 );
or   g04874 ( new_n7223 , new_n6628_1 , n8920 );
nor  g04875 ( new_n7224 , new_n7222 , new_n7223 );
nor  g04876 ( new_n7225 , new_n7221 , new_n7224 );
nor  g04877 ( new_n7226 , new_n7219 , new_n7225 );
nor  g04878 ( new_n7227 , new_n7218 , new_n7226 );
and  g04879 ( new_n7228 , new_n7216 , new_n7227 );
or   g04880 ( new_n7229_1 , new_n7215 , new_n7228 );
and  g04881 ( new_n7230_1 , new_n7214 , new_n7229_1 );
or   g04882 ( new_n7231 , new_n7213 , new_n7230_1 );
and  g04883 ( new_n7232 , new_n7212 , new_n7231 );
or   g04884 ( new_n7233_1 , new_n7211 , new_n7232 );
and  g04885 ( new_n7234 , new_n7210 , new_n7233_1 );
or   g04886 ( new_n7235 , new_n7209 , new_n7234 );
and  g04887 ( new_n7236_1 , new_n7208 , new_n7235 );
or   g04888 ( new_n7237 , new_n7207 , new_n7236_1 );
and  g04889 ( new_n7238 , new_n7206 , new_n7237 );
or   g04890 ( new_n7239 , new_n7205 , new_n7238 );
and  g04891 ( new_n7240 , new_n7204 , new_n7239 );
nor  g04892 ( new_n7241 , new_n7203 , new_n7240 );
not  g04893 ( new_n7242 , new_n7241 );
not  g04894 ( new_n7243 , n26986 );
nor  g04895 ( new_n7244 , n19282 , new_n7243 );
xnor g04896 ( new_n7245 , n19282 , n26986 );
and  g04897 ( new_n7246 , new_n2926 , n21287 );
xnor g04898 ( new_n7247 , n12657 , n21287 );
not  g04899 ( new_n7248 , n4256 );
nor  g04900 ( new_n7249 , new_n7248 , n17077 );
xnor g04901 ( new_n7250 , n4256 , n17077 );
not  g04902 ( new_n7251 , n26510 );
and  g04903 ( new_n7252 , n22332 , new_n7251 );
and  g04904 ( new_n7253_1 , new_n3814 , new_n3839 );
or   g04905 ( new_n7254 , new_n7252 , new_n7253_1 );
and  g04906 ( new_n7255 , new_n7250 , new_n7254 );
or   g04907 ( new_n7256_1 , new_n7249 , new_n7255 );
and  g04908 ( new_n7257 , new_n7247 , new_n7256_1 );
or   g04909 ( new_n7258 , new_n7246 , new_n7257 );
and  g04910 ( new_n7259 , new_n7245 , new_n7258 );
nor  g04911 ( new_n7260 , new_n7244 , new_n7259 );
xnor g04912 ( new_n7261 , new_n7242 , new_n7260 );
nor  g04913 ( new_n7262 , new_n7205 , new_n7238 );
xnor g04914 ( new_n7263 , new_n7204 , new_n7262 );
xor  g04915 ( new_n7264 , new_n7245 , new_n7258 );
and  g04916 ( new_n7265 , new_n7263 , new_n7264 );
not  g04917 ( new_n7266 , new_n7263 );
xnor g04918 ( new_n7267 , new_n7266 , new_n7264 );
nor  g04919 ( new_n7268_1 , new_n7207 , new_n7236_1 );
xnor g04920 ( new_n7269 , new_n7206 , new_n7268_1 );
xor  g04921 ( new_n7270 , new_n7247 , new_n7256_1 );
nor  g04922 ( new_n7271 , new_n7269 , new_n7270 );
xnor g04923 ( new_n7272 , new_n7269 , new_n7270 );
nor  g04924 ( new_n7273 , new_n7209 , new_n7234 );
xnor g04925 ( new_n7274 , new_n7208 , new_n7273 );
xor  g04926 ( new_n7275 , new_n7250 , new_n7254 );
nor  g04927 ( new_n7276 , new_n7274 , new_n7275 );
xnor g04928 ( new_n7277_1 , new_n7274 , new_n7275 );
xor  g04929 ( new_n7278 , new_n7210 , new_n7233_1 );
nor  g04930 ( new_n7279 , new_n3840 , new_n7278 );
xnor g04931 ( new_n7280_1 , new_n3840 , new_n7278 );
nor  g04932 ( new_n7281 , new_n7213 , new_n7230_1 );
xnor g04933 ( new_n7282 , new_n7212 , new_n7281 );
nor  g04934 ( new_n7283 , new_n3852 , new_n7282 );
xnor g04935 ( new_n7284 , new_n3852 , new_n7282 );
xor  g04936 ( new_n7285 , new_n7214 , new_n7229_1 );
nor  g04937 ( new_n7286 , new_n3856 , new_n7285 );
xnor g04938 ( new_n7287 , new_n3856 , new_n7285 );
xor  g04939 ( new_n7288 , new_n7216 , new_n7227 );
nor  g04940 ( new_n7289 , new_n3862 , new_n7288 );
not  g04941 ( new_n7290 , new_n7288 );
xnor g04942 ( new_n7291 , new_n3862 , new_n7290 );
xnor g04943 ( new_n7292 , n12161 , n26748 );
xor  g04944 ( new_n7293 , new_n7225 , new_n7292 );
nor  g04945 ( new_n7294 , new_n3868 , new_n7293 );
not  g04946 ( new_n7295 , new_n7293 );
xnor g04947 ( new_n7296 , new_n3868 , new_n7295 );
xnor g04948 ( new_n7297 , n5026 , n10057 );
xnor g04949 ( new_n7298_1 , new_n7223 , new_n7297 );
nor  g04950 ( new_n7299 , new_n3873 , new_n7298_1 );
xnor g04951 ( new_n7300 , n8581 , n8920 );
nor  g04952 ( new_n7301 , new_n3876 , new_n7300 );
not  g04953 ( new_n7302 , new_n7298_1 );
xnor g04954 ( new_n7303 , new_n3873 , new_n7302 );
and  g04955 ( new_n7304 , new_n7301 , new_n7303 );
nor  g04956 ( new_n7305_1 , new_n7299 , new_n7304 );
and  g04957 ( new_n7306 , new_n7296 , new_n7305_1 );
or   g04958 ( new_n7307 , new_n7294 , new_n7306 );
and  g04959 ( new_n7308_1 , new_n7291 , new_n7307 );
nor  g04960 ( new_n7309 , new_n7289 , new_n7308_1 );
nor  g04961 ( new_n7310 , new_n7287 , new_n7309 );
nor  g04962 ( new_n7311 , new_n7286 , new_n7310 );
nor  g04963 ( new_n7312 , new_n7284 , new_n7311 );
nor  g04964 ( new_n7313_1 , new_n7283 , new_n7312 );
nor  g04965 ( new_n7314 , new_n7280_1 , new_n7313_1 );
nor  g04966 ( new_n7315 , new_n7279 , new_n7314 );
nor  g04967 ( new_n7316 , new_n7277_1 , new_n7315 );
nor  g04968 ( new_n7317 , new_n7276 , new_n7316 );
nor  g04969 ( new_n7318 , new_n7272 , new_n7317 );
nor  g04970 ( new_n7319 , new_n7271 , new_n7318 );
and  g04971 ( new_n7320 , new_n7267 , new_n7319 );
nor  g04972 ( new_n7321 , new_n7265 , new_n7320 );
xnor g04973 ( new_n7322 , new_n7261 , new_n7321 );
not  g04974 ( new_n7323 , new_n7322 );
nor  g04975 ( new_n7324 , new_n4798 , n11898 );
xnor g04976 ( new_n7325 , n2979 , n11898 );
nor  g04977 ( new_n7326 , new_n4801 , n19941 );
xnor g04978 ( new_n7327 , n647 , n19941 );
not  g04979 ( new_n7328 , n20409 );
nor  g04980 ( new_n7329 , n1099 , new_n7328 );
xnor g04981 ( new_n7330_1 , n1099 , n20409 );
nor  g04982 ( new_n7331 , n2113 , new_n3725_1 );
xnor g04983 ( new_n7332 , n2113 , n25749 );
nor  g04984 ( new_n7333 , new_n3774 , n21134 );
xnor g04985 ( new_n7334 , n3161 , n21134 );
nor  g04986 ( new_n7335_1 , n6369 , new_n3778 );
xnor g04987 ( new_n7336 , n6369 , n9003 );
nor  g04988 ( new_n7337 , new_n3784 , n25797 );
xnor g04989 ( new_n7338 , n4957 , n25797 );
nor  g04990 ( new_n7339_1 , n7524 , new_n4178 );
nor  g04991 ( new_n7340 , new_n3788 , n15967 );
nor  g04992 ( new_n7341 , new_n3752 , n15743 );
or   g04993 ( new_n7342 , n13319 , new_n3794_1 );
nor  g04994 ( new_n7343 , n20658 , new_n3756 );
and  g04995 ( new_n7344 , new_n7342 , new_n7343 );
nor  g04996 ( new_n7345 , new_n7341 , new_n7344 );
nor  g04997 ( new_n7346_1 , new_n7340 , new_n7345 );
nor  g04998 ( new_n7347 , new_n7339_1 , new_n7346_1 );
and  g04999 ( new_n7348 , new_n7338 , new_n7347 );
or   g05000 ( new_n7349_1 , new_n7337 , new_n7348 );
and  g05001 ( new_n7350 , new_n7336 , new_n7349_1 );
or   g05002 ( new_n7351 , new_n7335_1 , new_n7350 );
and  g05003 ( new_n7352 , new_n7334 , new_n7351 );
or   g05004 ( new_n7353 , new_n7333 , new_n7352 );
and  g05005 ( new_n7354 , new_n7332 , new_n7353 );
or   g05006 ( new_n7355 , new_n7331 , new_n7354 );
and  g05007 ( new_n7356 , new_n7330_1 , new_n7355 );
or   g05008 ( new_n7357 , new_n7329 , new_n7356 );
and  g05009 ( new_n7358 , new_n7327 , new_n7357 );
or   g05010 ( new_n7359 , new_n7326 , new_n7358 );
and  g05011 ( new_n7360 , new_n7325 , new_n7359 );
nor  g05012 ( new_n7361 , new_n7324 , new_n7360 );
not  g05013 ( new_n7362 , new_n7361 );
xnor g05014 ( new_n7363_1 , new_n7323 , new_n7362 );
xor  g05015 ( new_n7364 , new_n7325 , new_n7359 );
xor  g05016 ( new_n7365 , new_n7267 , new_n7319 );
nor  g05017 ( new_n7366 , new_n7364 , new_n7365 );
xnor g05018 ( new_n7367 , new_n7364 , new_n7365 );
xor  g05019 ( new_n7368 , new_n7327 , new_n7357 );
xnor g05020 ( new_n7369 , new_n7272 , new_n7317 );
nor  g05021 ( new_n7370 , new_n7368 , new_n7369 );
xnor g05022 ( new_n7371 , new_n7368 , new_n7369 );
xor  g05023 ( new_n7372 , new_n7330_1 , new_n7355 );
xnor g05024 ( new_n7373 , new_n7277_1 , new_n7315 );
nor  g05025 ( new_n7374 , new_n7372 , new_n7373 );
xnor g05026 ( new_n7375 , new_n7372 , new_n7373 );
xor  g05027 ( new_n7376 , new_n7332 , new_n7353 );
xnor g05028 ( new_n7377_1 , new_n7280_1 , new_n7313_1 );
nor  g05029 ( new_n7378 , new_n7376 , new_n7377_1 );
xnor g05030 ( new_n7379 , new_n7376 , new_n7377_1 );
xor  g05031 ( new_n7380 , new_n7334 , new_n7351 );
xnor g05032 ( new_n7381 , new_n7284 , new_n7311 );
nor  g05033 ( new_n7382 , new_n7380 , new_n7381 );
xnor g05034 ( new_n7383 , new_n7380 , new_n7381 );
xor  g05035 ( new_n7384 , new_n7336 , new_n7349_1 );
xnor g05036 ( new_n7385 , new_n7287 , new_n7309 );
nor  g05037 ( new_n7386 , new_n7384 , new_n7385 );
xnor g05038 ( new_n7387 , new_n7384 , new_n7385 );
nor  g05039 ( new_n7388 , new_n7294 , new_n7306 );
xnor g05040 ( new_n7389 , new_n7291 , new_n7388 );
xnor g05041 ( new_n7390_1 , new_n7338 , new_n7347 );
and  g05042 ( new_n7391 , new_n7389 , new_n7390_1 );
xnor g05043 ( new_n7392 , new_n7296 , new_n7305_1 );
not  g05044 ( new_n7393 , new_n7392 );
xnor g05045 ( new_n7394 , n7524 , n15967 );
xnor g05046 ( new_n7395 , new_n7345 , new_n7394 );
and  g05047 ( new_n7396 , new_n7393 , new_n7395 );
xnor g05048 ( new_n7397 , new_n7393 , new_n7395 );
xnor g05049 ( new_n7398 , n20658 , n25435 );
not  g05050 ( new_n7399 , new_n7300 );
xnor g05051 ( new_n7400 , new_n3876 , new_n7399 );
not  g05052 ( new_n7401 , new_n7400 );
nor  g05053 ( new_n7402 , new_n7398 , new_n7401 );
xnor g05054 ( new_n7403_1 , n13319 , n15743 );
xnor g05055 ( new_n7404 , new_n7343 , new_n7403_1 );
nor  g05056 ( new_n7405 , new_n7402 , new_n7404 );
xnor g05057 ( new_n7406 , new_n7301 , new_n7303 );
not  g05058 ( new_n7407 , new_n7406 );
xnor g05059 ( new_n7408_1 , new_n7402 , new_n7404 );
nor  g05060 ( new_n7409 , new_n7407 , new_n7408_1 );
nor  g05061 ( new_n7410 , new_n7405 , new_n7409 );
nor  g05062 ( new_n7411 , new_n7397 , new_n7410 );
nor  g05063 ( new_n7412 , new_n7396 , new_n7411 );
xnor g05064 ( new_n7413 , new_n7389 , new_n7390_1 );
nor  g05065 ( new_n7414 , new_n7412 , new_n7413 );
nor  g05066 ( new_n7415 , new_n7391 , new_n7414 );
nor  g05067 ( new_n7416 , new_n7387 , new_n7415 );
nor  g05068 ( new_n7417 , new_n7386 , new_n7416 );
nor  g05069 ( new_n7418 , new_n7383 , new_n7417 );
nor  g05070 ( new_n7419 , new_n7382 , new_n7418 );
nor  g05071 ( new_n7420 , new_n7379 , new_n7419 );
nor  g05072 ( new_n7421_1 , new_n7378 , new_n7420 );
nor  g05073 ( new_n7422 , new_n7375 , new_n7421_1 );
nor  g05074 ( new_n7423 , new_n7374 , new_n7422 );
nor  g05075 ( new_n7424 , new_n7371 , new_n7423 );
nor  g05076 ( new_n7425 , new_n7370 , new_n7424 );
nor  g05077 ( new_n7426 , new_n7367 , new_n7425 );
nor  g05078 ( new_n7427 , new_n7366 , new_n7426 );
xnor g05079 ( n809 , new_n7363_1 , new_n7427 );
not  g05080 ( new_n7429 , n2978 );
nor  g05081 ( new_n7430 , new_n7429 , n19282 );
xnor g05082 ( new_n7431 , n2978 , n19282 );
nor  g05083 ( new_n7432_1 , n12657 , new_n6744 );
xnor g05084 ( new_n7433 , n12657 , n23697 );
nor  g05085 ( new_n7434 , new_n6748 , n17077 );
xnor g05086 ( new_n7435 , n2289 , n17077 );
nor  g05087 ( new_n7436 , new_n6752 , n26510 );
xnor g05088 ( new_n7437_1 , n1112 , n26510 );
nor  g05089 ( new_n7438 , new_n6756 , n23068 );
xnor g05090 ( new_n7439 , n20179 , n23068 );
not  g05091 ( new_n7440 , n19228 );
nor  g05092 ( new_n7441 , new_n7440 , n19514 );
xnor g05093 ( new_n7442 , n19228 , n19514 );
nor  g05094 ( new_n7443 , n10053 , new_n6763 );
xnor g05095 ( new_n7444 , n10053 , n15539 );
nor  g05096 ( new_n7445 , n8052 , new_n2947 );
nor  g05097 ( new_n7446 , new_n6767 , n8399 );
nor  g05098 ( new_n7447 , new_n3824 , n10158 );
not  g05099 ( new_n7448 , n10158 );
nor  g05100 ( new_n7449 , n9507 , new_n7448 );
nor  g05101 ( new_n7450 , n18962 , new_n2952 );
not  g05102 ( new_n7451 , new_n7450 );
nor  g05103 ( new_n7452 , new_n7449 , new_n7451 );
nor  g05104 ( new_n7453 , new_n7447 , new_n7452 );
nor  g05105 ( new_n7454 , new_n7446 , new_n7453 );
nor  g05106 ( new_n7455 , new_n7445 , new_n7454 );
and  g05107 ( new_n7456 , new_n7444 , new_n7455 );
or   g05108 ( new_n7457 , new_n7443 , new_n7456 );
and  g05109 ( new_n7458 , new_n7442 , new_n7457 );
or   g05110 ( new_n7459 , new_n7441 , new_n7458 );
and  g05111 ( new_n7460_1 , new_n7439 , new_n7459 );
or   g05112 ( new_n7461 , new_n7438 , new_n7460_1 );
and  g05113 ( new_n7462 , new_n7437_1 , new_n7461 );
or   g05114 ( new_n7463 , new_n7436 , new_n7462 );
and  g05115 ( new_n7464 , new_n7435 , new_n7463 );
or   g05116 ( new_n7465 , new_n7434 , new_n7464 );
and  g05117 ( new_n7466 , new_n7433 , new_n7465 );
or   g05118 ( new_n7467 , new_n7432_1 , new_n7466 );
and  g05119 ( new_n7468 , new_n7431 , new_n7467 );
nor  g05120 ( new_n7469 , new_n7430 , new_n7468 );
nor  g05121 ( new_n7470 , n22626 , n26986 );
not  g05122 ( new_n7471 , new_n2424 );
nor  g05123 ( new_n7472 , new_n7471 , new_n2431 );
not  g05124 ( new_n7473 , new_n7472 );
xnor g05125 ( new_n7474 , n1654 , n4256 );
nor  g05126 ( new_n7475_1 , n13783 , n22332 );
or   g05127 ( new_n7476 , new_n2427 , new_n2428 );
and  g05128 ( new_n7477_1 , new_n2426 , new_n7476 );
nor  g05129 ( new_n7478 , new_n7475_1 , new_n7477_1 );
xnor g05130 ( new_n7479 , new_n7474 , new_n7478 );
nor  g05131 ( new_n7480 , new_n7473 , new_n7479 );
not  g05132 ( new_n7481 , new_n7480 );
not  g05133 ( new_n7482 , n14440 );
xnor g05134 ( new_n7483 , new_n7482 , n21287 );
nor  g05135 ( new_n7484 , n1654 , n4256 );
nor  g05136 ( new_n7485 , new_n7474 , new_n7478 );
nor  g05137 ( new_n7486 , new_n7484 , new_n7485 );
xnor g05138 ( new_n7487 , new_n7483 , new_n7486 );
not  g05139 ( new_n7488 , new_n7487 );
nor  g05140 ( new_n7489 , new_n7481 , new_n7488 );
xnor g05141 ( new_n7490 , n22626 , n26986 );
nor  g05142 ( new_n7491 , n14440 , n21287 );
or   g05143 ( new_n7492 , new_n7484 , new_n7485 );
and  g05144 ( new_n7493 , new_n7483 , new_n7492 );
nor  g05145 ( new_n7494 , new_n7491 , new_n7493 );
xor  g05146 ( new_n7495 , new_n7490 , new_n7494 );
and  g05147 ( new_n7496 , new_n7489 , new_n7495 );
and  g05148 ( new_n7497 , new_n7470 , new_n7496 );
nor  g05149 ( new_n7498 , new_n7490 , new_n7494 );
nor  g05150 ( new_n7499 , new_n7470 , new_n7498 );
not  g05151 ( new_n7500 , new_n7499 );
nor  g05152 ( new_n7501 , new_n7496 , new_n7500 );
nor  g05153 ( new_n7502 , new_n7497 , new_n7501 );
nor  g05154 ( new_n7503 , n3425 , n13494 );
xnor g05155 ( new_n7504 , new_n3217 , n13494 );
not  g05156 ( new_n7505 , new_n7504 );
nor  g05157 ( new_n7506 , n9967 , n25345 );
xnor g05158 ( new_n7507_1 , new_n3198 , n25345 );
not  g05159 ( new_n7508 , n20946 );
nor  g05160 ( new_n7509 , new_n5506 , new_n7508 );
or   g05161 ( new_n7510 , n9655 , n20946 );
nor  g05162 ( new_n7511 , n7751 , n13490 );
nor  g05163 ( new_n7512 , new_n2433 , new_n2459 );
nor  g05164 ( new_n7513 , new_n7511 , new_n7512 );
and  g05165 ( new_n7514_1 , new_n7510 , new_n7513 );
nor  g05166 ( new_n7515 , new_n7509 , new_n7514_1 );
and  g05167 ( new_n7516 , new_n7507_1 , new_n7515 );
nor  g05168 ( new_n7517 , new_n7506 , new_n7516 );
nor  g05169 ( new_n7518 , new_n7505 , new_n7517 );
nor  g05170 ( new_n7519 , new_n7503 , new_n7518 );
and  g05171 ( new_n7520 , new_n7502 , new_n7519 );
or   g05172 ( new_n7521 , new_n7502 , new_n7519 );
xnor g05173 ( new_n7522 , new_n7490 , new_n7494 );
xnor g05174 ( new_n7523 , new_n7489 , new_n7522 );
xnor g05175 ( new_n7524_1 , new_n7505 , new_n7517 );
nor  g05176 ( new_n7525 , new_n7523 , new_n7524_1 );
xnor g05177 ( new_n7526 , new_n7523 , new_n7524_1 );
xnor g05178 ( new_n7527 , new_n7480 , new_n7488 );
xnor g05179 ( new_n7528 , new_n7507_1 , new_n7515 );
nor  g05180 ( new_n7529 , new_n7527 , new_n7528 );
xnor g05181 ( new_n7530 , new_n7527 , new_n7528 );
xnor g05182 ( new_n7531 , new_n7472 , new_n7479 );
xnor g05183 ( new_n7532 , n9655 , n20946 );
xnor g05184 ( new_n7533 , new_n7513 , new_n7532 );
nor  g05185 ( new_n7534 , new_n7531 , new_n7533 );
xnor g05186 ( new_n7535 , new_n7531 , new_n7533 );
nor  g05187 ( new_n7536 , new_n2432 , new_n2460 );
nor  g05188 ( new_n7537 , new_n2461 , new_n2500 );
nor  g05189 ( new_n7538 , new_n7536 , new_n7537 );
nor  g05190 ( new_n7539 , new_n7535 , new_n7538 );
nor  g05191 ( new_n7540 , new_n7534 , new_n7539 );
nor  g05192 ( new_n7541 , new_n7530 , new_n7540 );
nor  g05193 ( new_n7542 , new_n7529 , new_n7541 );
nor  g05194 ( new_n7543 , new_n7526 , new_n7542 );
nor  g05195 ( new_n7544 , new_n7525 , new_n7543 );
and  g05196 ( new_n7545 , new_n7521 , new_n7544 );
or   g05197 ( new_n7546 , new_n7497 , new_n7545 );
nor  g05198 ( new_n7547 , new_n7520 , new_n7546 );
xnor g05199 ( new_n7548 , new_n7469 , new_n7547 );
xnor g05200 ( new_n7549 , new_n7502 , new_n7519 );
xnor g05201 ( new_n7550 , new_n7544 , new_n7549 );
nor  g05202 ( new_n7551 , new_n7469 , new_n7550 );
xnor g05203 ( new_n7552 , new_n7469 , new_n7550 );
xor  g05204 ( new_n7553 , new_n7431 , new_n7467 );
xnor g05205 ( new_n7554 , new_n7526 , new_n7542 );
nor  g05206 ( new_n7555 , new_n7553 , new_n7554 );
xnor g05207 ( new_n7556 , new_n7553 , new_n7554 );
xor  g05208 ( new_n7557 , new_n7433 , new_n7465 );
xnor g05209 ( new_n7558_1 , new_n7530 , new_n7540 );
nor  g05210 ( new_n7559 , new_n7557 , new_n7558_1 );
xnor g05211 ( new_n7560 , new_n7557 , new_n7558_1 );
xor  g05212 ( new_n7561 , new_n7435 , new_n7463 );
xnor g05213 ( new_n7562 , new_n7535 , new_n7538 );
nor  g05214 ( new_n7563 , new_n7561 , new_n7562 );
xnor g05215 ( new_n7564 , new_n7561 , new_n7562 );
xor  g05216 ( new_n7565 , new_n7437_1 , new_n7461 );
nor  g05217 ( new_n7566_1 , new_n2501 , new_n7565 );
xnor g05218 ( new_n7567 , new_n2501 , new_n7565 );
xor  g05219 ( new_n7568 , new_n7439 , new_n7459 );
nor  g05220 ( new_n7569_1 , new_n2504 , new_n7568 );
xnor g05221 ( new_n7570 , new_n2504 , new_n7568 );
xor  g05222 ( new_n7571 , new_n7442 , new_n7457 );
nor  g05223 ( new_n7572_1 , new_n2508 , new_n7571 );
xnor g05224 ( new_n7573 , new_n2508 , new_n7571 );
xnor g05225 ( new_n7574 , new_n7444 , new_n7455 );
and  g05226 ( new_n7575_1 , new_n2513_1 , new_n7574 );
xnor g05227 ( new_n7576 , new_n2513_1 , new_n7574 );
xnor g05228 ( new_n7577 , n8052 , n8399 );
xnor g05229 ( new_n7578 , new_n7453 , new_n7577 );
and  g05230 ( new_n7579 , new_n2516 , new_n7578 );
xnor g05231 ( new_n7580 , new_n2516 , new_n7578 );
xnor g05232 ( new_n7581 , n18962 , n26979 );
or   g05233 ( new_n7582 , new_n2523 , new_n7581 );
xnor g05234 ( new_n7583 , n9507 , n10158 );
xnor g05235 ( new_n7584 , new_n7451 , new_n7583 );
and  g05236 ( new_n7585_1 , new_n7582 , new_n7584 );
xor  g05237 ( new_n7586 , new_n7582 , new_n7584 );
and  g05238 ( new_n7587 , new_n2529 , new_n7586 );
nor  g05239 ( new_n7588_1 , new_n7585_1 , new_n7587 );
nor  g05240 ( new_n7589 , new_n7580 , new_n7588_1 );
nor  g05241 ( new_n7590 , new_n7579 , new_n7589 );
nor  g05242 ( new_n7591 , new_n7576 , new_n7590 );
nor  g05243 ( new_n7592 , new_n7575_1 , new_n7591 );
nor  g05244 ( new_n7593_1 , new_n7573 , new_n7592 );
nor  g05245 ( new_n7594 , new_n7572_1 , new_n7593_1 );
nor  g05246 ( new_n7595 , new_n7570 , new_n7594 );
nor  g05247 ( new_n7596 , new_n7569_1 , new_n7595 );
nor  g05248 ( new_n7597 , new_n7567 , new_n7596 );
nor  g05249 ( new_n7598_1 , new_n7566_1 , new_n7597 );
nor  g05250 ( new_n7599 , new_n7564 , new_n7598_1 );
nor  g05251 ( new_n7600 , new_n7563 , new_n7599 );
nor  g05252 ( new_n7601 , new_n7560 , new_n7600 );
nor  g05253 ( new_n7602 , new_n7559 , new_n7601 );
nor  g05254 ( new_n7603 , new_n7556 , new_n7602 );
nor  g05255 ( new_n7604 , new_n7555 , new_n7603 );
nor  g05256 ( new_n7605 , new_n7552 , new_n7604 );
nor  g05257 ( new_n7606 , new_n7551 , new_n7605 );
xnor g05258 ( n819 , new_n7548 , new_n7606 );
not  g05259 ( new_n7608 , n8856 );
nor  g05260 ( new_n7609 , new_n7608 , n22626 );
xnor g05261 ( new_n7610_1 , n8856 , n22626 );
nor  g05262 ( new_n7611 , new_n3405 , n14440 );
xnor g05263 ( new_n7612 , n14130 , n14440 );
not  g05264 ( new_n7613 , n1654 );
and  g05265 ( new_n7614 , new_n7613 , n16482 );
xnor g05266 ( new_n7615 , n1654 , n16482 );
and  g05267 ( new_n7616_1 , n9942 , new_n2425 );
xnor g05268 ( new_n7617 , n9942 , n13783 );
not  g05269 ( new_n7618 , n26660 );
and  g05270 ( new_n7619 , n25643 , new_n7618 );
xnor g05271 ( new_n7620 , n25643 , n26660 );
nor  g05272 ( new_n7621 , n3018 , new_n5116 );
xnor g05273 ( new_n7622 , n3018 , n9557 );
nor  g05274 ( new_n7623 , new_n5106 , n3480 );
xnor g05275 ( new_n7624 , n3136 , n3480 );
not  g05276 ( new_n7625 , n16722 );
nor  g05277 ( new_n7626 , n6385 , new_n7625 );
nor  g05278 ( new_n7627 , new_n2359 , n16722 );
nor  g05279 ( new_n7628 , new_n5784 , n20138 );
nor  g05280 ( new_n7629 , n11486 , new_n2363_1 );
nor  g05281 ( new_n7630_1 , n9251 , new_n2383 );
not  g05282 ( new_n7631 , new_n7630_1 );
nor  g05283 ( new_n7632 , new_n7629 , new_n7631 );
nor  g05284 ( new_n7633 , new_n7628 , new_n7632 );
nor  g05285 ( new_n7634 , new_n7627 , new_n7633 );
nor  g05286 ( new_n7635 , new_n7626 , new_n7634 );
and  g05287 ( new_n7636 , new_n7624 , new_n7635 );
or   g05288 ( new_n7637 , new_n7623 , new_n7636 );
and  g05289 ( new_n7638 , new_n7622 , new_n7637 );
or   g05290 ( new_n7639 , new_n7621 , new_n7638 );
and  g05291 ( new_n7640 , new_n7620 , new_n7639 );
or   g05292 ( new_n7641 , new_n7619 , new_n7640 );
and  g05293 ( new_n7642 , new_n7617 , new_n7641 );
or   g05294 ( new_n7643_1 , new_n7616_1 , new_n7642 );
and  g05295 ( new_n7644 , new_n7615 , new_n7643_1 );
or   g05296 ( new_n7645 , new_n7614 , new_n7644 );
and  g05297 ( new_n7646 , new_n7612 , new_n7645 );
or   g05298 ( new_n7647_1 , new_n7611 , new_n7646 );
and  g05299 ( new_n7648 , new_n7610_1 , new_n7647_1 );
nor  g05300 ( new_n7649 , new_n7609 , new_n7648 );
not  g05301 ( new_n7650 , new_n7649 );
nor  g05302 ( new_n7651 , new_n5982 , n25120 );
xnor g05303 ( new_n7652 , n3582 , n25120 );
nor  g05304 ( new_n7653 , new_n5985 , n8363 );
xnor g05305 ( new_n7654 , n2145 , n8363 );
nor  g05306 ( new_n7655 , new_n5988 , n14680 );
xnor g05307 ( new_n7656 , n5031 , n14680 );
not  g05308 ( new_n7657_1 , n11044 );
nor  g05309 ( new_n7658 , new_n7657_1 , n17250 );
xnor g05310 ( new_n7659 , n11044 , n17250 );
nor  g05311 ( new_n7660 , new_n5994 , n23160 );
xnor g05312 ( new_n7661 , n2421 , n23160 );
not  g05313 ( new_n7662 , n987 );
nor  g05314 ( new_n7663 , new_n7662 , n16524 );
xnor g05315 ( new_n7664 , n987 , n16524 );
not  g05316 ( new_n7665 , n20478 );
nor  g05317 ( new_n7666 , n11056 , new_n7665 );
xnor g05318 ( new_n7667 , n11056 , n20478 );
not  g05319 ( new_n7668 , n15271 );
nor  g05320 ( new_n7669 , new_n7668 , n26882 );
not  g05321 ( new_n7670_1 , n26882 );
nor  g05322 ( new_n7671 , n15271 , new_n7670_1 );
not  g05323 ( new_n7672 , n22619 );
and  g05324 ( new_n7673 , new_n7672 , n25877 );
nor  g05325 ( new_n7674_1 , new_n7672 , n25877 );
nor  g05326 ( new_n7675 , n6775 , new_n6629 );
not  g05327 ( new_n7676 , new_n7675 );
nor  g05328 ( new_n7677 , new_n7674_1 , new_n7676 );
nor  g05329 ( new_n7678_1 , new_n7673 , new_n7677 );
nor  g05330 ( new_n7679_1 , new_n7671 , new_n7678_1 );
nor  g05331 ( new_n7680 , new_n7669 , new_n7679_1 );
and  g05332 ( new_n7681 , new_n7667 , new_n7680 );
or   g05333 ( new_n7682 , new_n7666 , new_n7681 );
and  g05334 ( new_n7683 , new_n7664 , new_n7682 );
or   g05335 ( new_n7684 , new_n7663 , new_n7683 );
and  g05336 ( new_n7685 , new_n7661 , new_n7684 );
or   g05337 ( new_n7686_1 , new_n7660 , new_n7685 );
and  g05338 ( new_n7687 , new_n7659 , new_n7686_1 );
or   g05339 ( new_n7688 , new_n7658 , new_n7687 );
and  g05340 ( new_n7689 , new_n7656 , new_n7688 );
or   g05341 ( new_n7690 , new_n7655 , new_n7689 );
and  g05342 ( new_n7691 , new_n7654 , new_n7690 );
or   g05343 ( new_n7692_1 , new_n7653 , new_n7691 );
and  g05344 ( new_n7693_1 , new_n7652 , new_n7692_1 );
nor  g05345 ( new_n7694 , new_n7651 , new_n7693_1 );
not  g05346 ( new_n7695 , new_n7694 );
xnor g05347 ( new_n7696 , new_n7650 , new_n7695 );
nor  g05348 ( new_n7697 , new_n7653 , new_n7691 );
xnor g05349 ( new_n7698_1 , new_n7652 , new_n7697 );
nor  g05350 ( new_n7699 , new_n7611 , new_n7646 );
xnor g05351 ( new_n7700 , new_n7610_1 , new_n7699 );
nor  g05352 ( new_n7701 , new_n7698_1 , new_n7700 );
not  g05353 ( new_n7702 , new_n7698_1 );
not  g05354 ( new_n7703 , new_n7700 );
xnor g05355 ( new_n7704 , new_n7702 , new_n7703 );
xor  g05356 ( new_n7705 , new_n7654 , new_n7690 );
xor  g05357 ( new_n7706 , new_n7612 , new_n7645 );
nor  g05358 ( new_n7707 , new_n7705 , new_n7706 );
xnor g05359 ( new_n7708_1 , new_n7705 , new_n7706 );
nor  g05360 ( new_n7709 , new_n7658 , new_n7687 );
xnor g05361 ( new_n7710 , new_n7656 , new_n7709 );
nor  g05362 ( new_n7711 , new_n7616_1 , new_n7642 );
xnor g05363 ( new_n7712 , new_n7615 , new_n7711 );
nor  g05364 ( new_n7713 , new_n7710 , new_n7712 );
not  g05365 ( new_n7714 , new_n7710 );
not  g05366 ( new_n7715 , new_n7712 );
xnor g05367 ( new_n7716 , new_n7714 , new_n7715 );
xor  g05368 ( new_n7717 , new_n7659 , new_n7686_1 );
xor  g05369 ( new_n7718 , new_n7617 , new_n7641 );
nor  g05370 ( new_n7719 , new_n7717 , new_n7718 );
xnor g05371 ( new_n7720 , new_n7717 , new_n7718 );
xor  g05372 ( new_n7721_1 , new_n7661 , new_n7684 );
xor  g05373 ( new_n7722 , new_n7620 , new_n7639 );
nor  g05374 ( new_n7723 , new_n7721_1 , new_n7722 );
xnor g05375 ( new_n7724 , new_n7721_1 , new_n7722 );
xor  g05376 ( new_n7725 , new_n7664 , new_n7682 );
xor  g05377 ( new_n7726 , new_n7622 , new_n7637 );
nor  g05378 ( new_n7727 , new_n7725 , new_n7726 );
xnor g05379 ( new_n7728 , new_n7725 , new_n7726 );
xnor g05380 ( new_n7729 , new_n7667 , new_n7680 );
not  g05381 ( new_n7730 , new_n7729 );
xor  g05382 ( new_n7731_1 , new_n7624 , new_n7635 );
nor  g05383 ( new_n7732 , new_n7730 , new_n7731_1 );
xnor g05384 ( new_n7733 , new_n7730 , new_n7731_1 );
xnor g05385 ( new_n7734 , n15271 , n26882 );
xnor g05386 ( new_n7735 , new_n7678_1 , new_n7734 );
xnor g05387 ( new_n7736 , n6385 , n16722 );
xnor g05388 ( new_n7737 , new_n7633 , new_n7736 );
and  g05389 ( new_n7738 , new_n7735 , new_n7737 );
not  g05390 ( new_n7739 , new_n7735 );
xnor g05391 ( new_n7740 , new_n7739 , new_n7737 );
xnor g05392 ( new_n7741 , n22619 , n25877 );
xnor g05393 ( new_n7742 , new_n7676 , new_n7741 );
not  g05394 ( new_n7743 , new_n7742 );
xnor g05395 ( new_n7744 , n11486 , n20138 );
xnor g05396 ( new_n7745 , new_n7631 , new_n7744 );
not  g05397 ( new_n7746 , new_n7745 );
nor  g05398 ( new_n7747 , new_n7743 , new_n7746 );
xnor g05399 ( new_n7748 , n6775 , n24323 );
xnor g05400 ( new_n7749 , n9251 , n13781 );
or   g05401 ( new_n7750 , new_n7748 , new_n7749 );
xnor g05402 ( new_n7751_1 , new_n7743 , new_n7745 );
and  g05403 ( new_n7752 , new_n7750 , new_n7751_1 );
or   g05404 ( new_n7753 , new_n7747 , new_n7752 );
and  g05405 ( new_n7754 , new_n7740 , new_n7753 );
nor  g05406 ( new_n7755 , new_n7738 , new_n7754 );
nor  g05407 ( new_n7756 , new_n7733 , new_n7755 );
nor  g05408 ( new_n7757 , new_n7732 , new_n7756 );
nor  g05409 ( new_n7758 , new_n7728 , new_n7757 );
nor  g05410 ( new_n7759_1 , new_n7727 , new_n7758 );
nor  g05411 ( new_n7760 , new_n7724 , new_n7759_1 );
nor  g05412 ( new_n7761 , new_n7723 , new_n7760 );
nor  g05413 ( new_n7762 , new_n7720 , new_n7761 );
nor  g05414 ( new_n7763 , new_n7719 , new_n7762 );
nor  g05415 ( new_n7764 , new_n7716 , new_n7763 );
nor  g05416 ( new_n7765 , new_n7713 , new_n7764 );
nor  g05417 ( new_n7766 , new_n7708_1 , new_n7765 );
nor  g05418 ( new_n7767 , new_n7707 , new_n7766 );
nor  g05419 ( new_n7768 , new_n7704 , new_n7767 );
nor  g05420 ( new_n7769_1 , new_n7701 , new_n7768 );
xnor g05421 ( new_n7770 , new_n7696 , new_n7769_1 );
not  g05422 ( new_n7771 , new_n7770 );
not  g05423 ( new_n7772 , n9554 );
not  g05424 ( new_n7773_1 , n26408 );
nor  g05425 ( new_n7774 , n2809 , n15508 );
not  g05426 ( new_n7775 , new_n7774 );
nor  g05427 ( new_n7776 , n19680 , new_n7775 );
not  g05428 ( new_n7777 , new_n7776 );
nor  g05429 ( new_n7778 , n7421 , new_n7777 );
not  g05430 ( new_n7779 , new_n7778 );
nor  g05431 ( new_n7780_1 , n13453 , new_n7779 );
not  g05432 ( new_n7781 , new_n7780_1 );
nor  g05433 ( new_n7782 , n11630 , new_n7781 );
not  g05434 ( new_n7783 , new_n7782 );
nor  g05435 ( new_n7784 , n7377 , new_n7783 );
not  g05436 ( new_n7785 , new_n7784 );
nor  g05437 ( new_n7786 , n18227 , new_n7785 );
and  g05438 ( new_n7787 , new_n7773_1 , new_n7786 );
and  g05439 ( new_n7788_1 , new_n7772 , new_n7787 );
xnor g05440 ( new_n7789 , n9554 , new_n7787 );
nor  g05441 ( new_n7790 , n9259 , new_n7789 );
xnor g05442 ( new_n7791 , n26408 , new_n7786 );
nor  g05443 ( new_n7792 , n21489 , new_n7791 );
xnor g05444 ( new_n7793 , new_n3583 , new_n7791 );
xnor g05445 ( new_n7794_1 , n18227 , new_n7784 );
nor  g05446 ( new_n7795 , n20213 , new_n7794_1 );
xnor g05447 ( new_n7796 , new_n4844 , new_n7794_1 );
xnor g05448 ( new_n7797 , n7377 , new_n7782 );
nor  g05449 ( new_n7798 , n13912 , new_n7797 );
xnor g05450 ( new_n7799 , new_n4848 , new_n7797 );
xnor g05451 ( new_n7800 , n11630 , new_n7780_1 );
nor  g05452 ( new_n7801 , n7670 , new_n7800 );
xnor g05453 ( new_n7802 , new_n4853 , new_n7800 );
xnor g05454 ( new_n7803 , n13453 , new_n7778 );
nor  g05455 ( new_n7804 , n9598 , new_n7803 );
xnor g05456 ( new_n7805 , new_n4857 , new_n7803 );
xnor g05457 ( new_n7806 , n7421 , new_n7776 );
nor  g05458 ( new_n7807 , n22290 , new_n7806 );
xnor g05459 ( new_n7808 , n19680 , new_n7774 );
nor  g05460 ( new_n7809 , n11273 , new_n7808 );
xnor g05461 ( new_n7810 , new_n4867 , new_n7808 );
xnor g05462 ( new_n7811_1 , new_n6616 , n15508 );
nor  g05463 ( new_n7812 , n25565 , new_n7811_1 );
nor  g05464 ( new_n7813 , new_n4818 , new_n3635 );
xnor g05465 ( new_n7814 , n25565 , new_n7811_1 );
nor  g05466 ( new_n7815 , new_n7813 , new_n7814 );
or   g05467 ( new_n7816 , new_n7812 , new_n7815 );
and  g05468 ( new_n7817 , new_n7810 , new_n7816 );
or   g05469 ( new_n7818 , new_n7809 , new_n7817 );
xnor g05470 ( new_n7819 , new_n4863 , new_n7806 );
and  g05471 ( new_n7820 , new_n7818 , new_n7819 );
or   g05472 ( new_n7821 , new_n7807 , new_n7820 );
and  g05473 ( new_n7822 , new_n7805 , new_n7821 );
or   g05474 ( new_n7823 , new_n7804 , new_n7822 );
and  g05475 ( new_n7824 , new_n7802 , new_n7823 );
or   g05476 ( new_n7825 , new_n7801 , new_n7824 );
and  g05477 ( new_n7826 , new_n7799 , new_n7825 );
or   g05478 ( new_n7827 , new_n7798 , new_n7826 );
and  g05479 ( new_n7828 , new_n7796 , new_n7827 );
or   g05480 ( new_n7829 , new_n7795 , new_n7828 );
and  g05481 ( new_n7830_1 , new_n7793 , new_n7829 );
nor  g05482 ( new_n7831 , new_n7792 , new_n7830_1 );
and  g05483 ( new_n7832 , n9259 , new_n7789 );
nor  g05484 ( new_n7833 , new_n7831 , new_n7832 );
nor  g05485 ( new_n7834_1 , new_n7790 , new_n7833 );
nor  g05486 ( new_n7835 , new_n7788_1 , new_n7834_1 );
xnor g05487 ( new_n7836 , new_n7771 , new_n7835 );
xnor g05488 ( new_n7837 , new_n7704 , new_n7767 );
xnor g05489 ( new_n7838 , new_n4797 , new_n7789 );
xnor g05490 ( new_n7839 , new_n7831 , new_n7838 );
not  g05491 ( new_n7840 , new_n7839 );
nor  g05492 ( new_n7841_1 , new_n7837 , new_n7840 );
not  g05493 ( new_n7842 , new_n7837 );
xnor g05494 ( new_n7843 , new_n7842 , new_n7840 );
xnor g05495 ( new_n7844 , new_n7708_1 , new_n7765 );
not  g05496 ( new_n7845 , new_n7844 );
nor  g05497 ( new_n7846 , new_n7795 , new_n7828 );
xnor g05498 ( new_n7847 , new_n7793 , new_n7846 );
nor  g05499 ( new_n7848 , new_n7845 , new_n7847 );
not  g05500 ( new_n7849 , new_n7847 );
xnor g05501 ( new_n7850 , new_n7845 , new_n7849 );
xnor g05502 ( new_n7851 , new_n7716 , new_n7763 );
not  g05503 ( new_n7852 , new_n7851 );
nor  g05504 ( new_n7853 , new_n7798 , new_n7826 );
xnor g05505 ( new_n7854 , new_n7796 , new_n7853 );
nor  g05506 ( new_n7855 , new_n7852 , new_n7854 );
not  g05507 ( new_n7856 , new_n7854 );
xnor g05508 ( new_n7857 , new_n7852 , new_n7856 );
xnor g05509 ( new_n7858 , new_n7720 , new_n7761 );
nor  g05510 ( new_n7859 , new_n7801 , new_n7824 );
xnor g05511 ( new_n7860 , new_n7799 , new_n7859 );
not  g05512 ( new_n7861 , new_n7860 );
nor  g05513 ( new_n7862 , new_n7858 , new_n7861 );
and  g05514 ( new_n7863 , new_n7858 , new_n7861 );
xnor g05515 ( new_n7864 , new_n7724 , new_n7759_1 );
not  g05516 ( new_n7865 , new_n7864 );
xor  g05517 ( new_n7866 , new_n7802 , new_n7823 );
and  g05518 ( new_n7867 , new_n7865 , new_n7866 );
xnor g05519 ( new_n7868 , new_n7865 , new_n7866 );
xor  g05520 ( new_n7869 , new_n7805 , new_n7821 );
not  g05521 ( new_n7870 , new_n7869 );
xnor g05522 ( new_n7871 , new_n7728 , new_n7757 );
nor  g05523 ( new_n7872 , new_n7870 , new_n7871 );
xnor g05524 ( new_n7873 , new_n7870 , new_n7871 );
xnor g05525 ( new_n7874 , new_n7733 , new_n7755 );
nor  g05526 ( new_n7875 , new_n7809 , new_n7817 );
xnor g05527 ( new_n7876_1 , new_n7875 , new_n7819 );
not  g05528 ( new_n7877 , new_n7876_1 );
nor  g05529 ( new_n7878 , new_n7874 , new_n7877 );
not  g05530 ( new_n7879 , new_n7874 );
or   g05531 ( new_n7880 , new_n7879 , new_n7876_1 );
nor  g05532 ( new_n7881 , new_n7747 , new_n7752 );
xnor g05533 ( new_n7882 , new_n7740 , new_n7881 );
xor  g05534 ( new_n7883 , new_n7750 , new_n7751_1 );
not  g05535 ( new_n7884_1 , new_n7883 );
xnor g05536 ( new_n7885 , new_n7813 , new_n7814 );
nor  g05537 ( new_n7886 , new_n7884_1 , new_n7885 );
xnor g05538 ( new_n7887 , n15508 , n21993 );
not  g05539 ( new_n7888 , new_n7748 );
xnor g05540 ( new_n7889 , new_n7888 , new_n7749 );
not  g05541 ( new_n7890 , new_n7889 );
nor  g05542 ( new_n7891 , new_n7887 , new_n7890 );
xnor g05543 ( new_n7892 , new_n7884_1 , new_n7885 );
nor  g05544 ( new_n7893 , new_n7891 , new_n7892 );
nor  g05545 ( new_n7894 , new_n7886 , new_n7893 );
not  g05546 ( new_n7895 , new_n7894 );
nor  g05547 ( new_n7896 , new_n7882 , new_n7895 );
nor  g05548 ( new_n7897 , new_n7812 , new_n7815 );
xnor g05549 ( new_n7898 , new_n7810 , new_n7897 );
not  g05550 ( new_n7899 , new_n7898 );
xnor g05551 ( new_n7900 , new_n7882 , new_n7894 );
and  g05552 ( new_n7901 , new_n7899 , new_n7900 );
nor  g05553 ( new_n7902 , new_n7896 , new_n7901 );
and  g05554 ( new_n7903 , new_n7880 , new_n7902 );
nor  g05555 ( new_n7904 , new_n7878 , new_n7903 );
nor  g05556 ( new_n7905 , new_n7873 , new_n7904 );
nor  g05557 ( new_n7906 , new_n7872 , new_n7905 );
nor  g05558 ( new_n7907 , new_n7868 , new_n7906 );
nor  g05559 ( new_n7908 , new_n7867 , new_n7907 );
nor  g05560 ( new_n7909 , new_n7863 , new_n7908 );
nor  g05561 ( new_n7910 , new_n7862 , new_n7909 );
and  g05562 ( new_n7911 , new_n7857 , new_n7910 );
or   g05563 ( new_n7912 , new_n7855 , new_n7911 );
and  g05564 ( new_n7913 , new_n7850 , new_n7912 );
nor  g05565 ( new_n7914 , new_n7848 , new_n7913 );
and  g05566 ( new_n7915 , new_n7843 , new_n7914 );
nor  g05567 ( new_n7916 , new_n7841_1 , new_n7915 );
xor  g05568 ( n829 , new_n7836 , new_n7916 );
not  g05569 ( new_n7918 , n14826 );
xnor g05570 ( new_n7919 , new_n7918 , n23272 );
nor  g05571 ( new_n7920 , n11481 , n23493 );
xnor g05572 ( new_n7921 , new_n4361 , n23493 );
nor  g05573 ( new_n7922 , n10275 , n16439 );
not  g05574 ( new_n7923 , n10275 );
xnor g05575 ( new_n7924 , new_n7923 , n16439 );
nor  g05576 ( new_n7925 , n15146 , n15241 );
not  g05577 ( new_n7926 , n15146 );
xnor g05578 ( new_n7927 , new_n7926 , n15241 );
nor  g05579 ( new_n7928 , n7678 , n11579 );
xnor g05580 ( new_n7929 , new_n4373 , n11579 );
nor  g05581 ( new_n7930 , n21 , n3785 );
not  g05582 ( new_n7931 , n21 );
xnor g05583 ( new_n7932 , new_n7931 , n3785 );
nor  g05584 ( new_n7933 , n1682 , n20250 );
not  g05585 ( new_n7934 , n1682 );
xnor g05586 ( new_n7935 , new_n7934 , n20250 );
nor  g05587 ( new_n7936 , n5822 , n7963 );
xnor g05588 ( new_n7937_1 , new_n4384 , n7963 );
nor  g05589 ( new_n7938 , n10017 , n26443 );
not  g05590 ( new_n7939 , n3618 );
or   g05591 ( new_n7940 , new_n4394 , new_n7939 );
not  g05592 ( new_n7941 , n10017 );
xnor g05593 ( new_n7942 , new_n7941 , n26443 );
and  g05594 ( new_n7943_1 , new_n7940 , new_n7942 );
or   g05595 ( new_n7944 , new_n7938 , new_n7943_1 );
and  g05596 ( new_n7945 , new_n7937_1 , new_n7944 );
or   g05597 ( new_n7946 , new_n7936 , new_n7945 );
and  g05598 ( new_n7947 , new_n7935 , new_n7946 );
or   g05599 ( new_n7948 , new_n7933 , new_n7947 );
and  g05600 ( new_n7949_1 , new_n7932 , new_n7948 );
or   g05601 ( new_n7950_1 , new_n7930 , new_n7949_1 );
and  g05602 ( new_n7951 , new_n7929 , new_n7950_1 );
or   g05603 ( new_n7952 , new_n7928 , new_n7951 );
and  g05604 ( new_n7953 , new_n7927 , new_n7952 );
or   g05605 ( new_n7954 , new_n7925 , new_n7953 );
and  g05606 ( new_n7955 , new_n7924 , new_n7954 );
or   g05607 ( new_n7956 , new_n7922 , new_n7955 );
and  g05608 ( new_n7957 , new_n7921 , new_n7956 );
nor  g05609 ( new_n7958 , new_n7920 , new_n7957 );
xnor g05610 ( new_n7959_1 , new_n7919 , new_n7958 );
nor  g05611 ( new_n7960 , n22764 , new_n7959_1 );
not  g05612 ( new_n7961 , new_n7959_1 );
xnor g05613 ( new_n7962 , n22764 , new_n7961 );
nor  g05614 ( new_n7963_1 , new_n7922 , new_n7955 );
xnor g05615 ( new_n7964 , new_n7921 , new_n7963_1 );
nor  g05616 ( new_n7965 , n26264 , new_n7964 );
not  g05617 ( new_n7966 , new_n7964 );
xnor g05618 ( new_n7967 , n26264 , new_n7966 );
nor  g05619 ( new_n7968_1 , new_n7925 , new_n7953 );
xnor g05620 ( new_n7969 , new_n7924 , new_n7968_1 );
nor  g05621 ( new_n7970 , n7841 , new_n7969 );
not  g05622 ( new_n7971 , new_n7969 );
xnor g05623 ( new_n7972 , n7841 , new_n7971 );
nor  g05624 ( new_n7973 , new_n7928 , new_n7951 );
xnor g05625 ( new_n7974 , new_n7927 , new_n7973 );
nor  g05626 ( new_n7975 , n16812 , new_n7974 );
not  g05627 ( new_n7976 , new_n7974 );
xnor g05628 ( new_n7977 , n16812 , new_n7976 );
nor  g05629 ( new_n7978 , new_n7930 , new_n7949_1 );
xnor g05630 ( new_n7979 , new_n7929 , new_n7978 );
nor  g05631 ( new_n7980 , n25068 , new_n7979 );
not  g05632 ( new_n7981 , new_n7979 );
xnor g05633 ( new_n7982 , n25068 , new_n7981 );
nor  g05634 ( new_n7983 , new_n7933 , new_n7947 );
xnor g05635 ( new_n7984 , new_n7932 , new_n7983 );
nor  g05636 ( new_n7985 , n2331 , new_n7984 );
not  g05637 ( new_n7986 , new_n7984 );
xnor g05638 ( new_n7987 , n2331 , new_n7986 );
nor  g05639 ( new_n7988 , new_n7936 , new_n7945 );
xnor g05640 ( new_n7989 , new_n7935 , new_n7988 );
nor  g05641 ( new_n7990 , n22631 , new_n7989 );
not  g05642 ( new_n7991 , new_n7989 );
xnor g05643 ( new_n7992_1 , n22631 , new_n7991 );
not  g05644 ( new_n7993 , n16743 );
xor  g05645 ( new_n7994 , new_n7937_1 , new_n7944 );
not  g05646 ( new_n7995 , new_n7994 );
nor  g05647 ( new_n7996 , new_n7993 , new_n7995 );
xnor g05648 ( new_n7997 , n16743 , new_n7995 );
not  g05649 ( new_n7998 , n15258 );
nor  g05650 ( new_n7999_1 , n4588 , new_n2543 );
and  g05651 ( new_n8000 , new_n7998 , new_n7999_1 );
nor  g05652 ( new_n8001 , new_n4394 , new_n7939 );
xnor g05653 ( new_n8002 , new_n8001 , new_n7942 );
not  g05654 ( new_n8003 , new_n8002 );
xnor g05655 ( new_n8004 , n15258 , new_n7999_1 );
and  g05656 ( new_n8005 , new_n8003 , new_n8004 );
nor  g05657 ( new_n8006_1 , new_n8000 , new_n8005 );
and  g05658 ( new_n8007 , new_n7997 , new_n8006_1 );
nor  g05659 ( new_n8008 , new_n7996 , new_n8007 );
and  g05660 ( new_n8009 , new_n7992_1 , new_n8008 );
or   g05661 ( new_n8010 , new_n7990 , new_n8009 );
and  g05662 ( new_n8011 , new_n7987 , new_n8010 );
or   g05663 ( new_n8012 , new_n7985 , new_n8011 );
and  g05664 ( new_n8013 , new_n7982 , new_n8012 );
or   g05665 ( new_n8014 , new_n7980 , new_n8013 );
and  g05666 ( new_n8015 , new_n7977 , new_n8014 );
or   g05667 ( new_n8016 , new_n7975 , new_n8015 );
and  g05668 ( new_n8017 , new_n7972 , new_n8016 );
or   g05669 ( new_n8018 , new_n7970 , new_n8017 );
and  g05670 ( new_n8019 , new_n7967 , new_n8018 );
or   g05671 ( new_n8020 , new_n7965 , new_n8019 );
and  g05672 ( new_n8021 , new_n7962 , new_n8020 );
nor  g05673 ( new_n8022 , new_n7960 , new_n8021 );
nor  g05674 ( new_n8023 , n14826 , n23272 );
or   g05675 ( new_n8024 , new_n7920 , new_n7957 );
and  g05676 ( new_n8025 , new_n7919 , new_n8024 );
nor  g05677 ( new_n8026 , new_n8023 , new_n8025 );
not  g05678 ( new_n8027_1 , new_n8026 );
and  g05679 ( new_n8028 , new_n8022 , new_n8027_1 );
nor  g05680 ( new_n8029 , new_n5686 , n18105 );
xnor g05681 ( new_n8030 , n12702 , n18105 );
nor  g05682 ( new_n8031_1 , n24196 , new_n5611 );
xnor g05683 ( new_n8032 , n24196 , n26797 );
not  g05684 ( new_n8033 , n23913 );
nor  g05685 ( new_n8034 , n16376 , new_n8033 );
xnor g05686 ( new_n8035 , n16376 , n23913 );
not  g05687 ( new_n8036 , n22554 );
nor  g05688 ( new_n8037 , new_n8036 , n25381 );
xnor g05689 ( new_n8038 , n22554 , n25381 );
not  g05690 ( new_n8039 , n20429 );
nor  g05691 ( new_n8040 , n12587 , new_n8039 );
xnor g05692 ( new_n8041 , n12587 , n20429 );
not  g05693 ( new_n8042_1 , n3909 );
nor  g05694 ( new_n8043 , n268 , new_n8042_1 );
xnor g05695 ( new_n8044 , n268 , n3909 );
not  g05696 ( new_n8045 , n23974 );
nor  g05697 ( new_n8046 , new_n8045 , n24879 );
xnor g05698 ( new_n8047 , n23974 , n24879 );
not  g05699 ( new_n8048 , n6785 );
nor  g05700 ( new_n8049 , n2146 , new_n8048 );
not  g05701 ( new_n8050 , n2146 );
nor  g05702 ( new_n8051 , new_n8050 , n6785 );
not  g05703 ( new_n8052_1 , n24032 );
nor  g05704 ( new_n8053 , n22173 , new_n8052_1 );
nor  g05705 ( new_n8054 , n583 , new_n4507 );
not  g05706 ( new_n8055 , n22173 );
or   g05707 ( new_n8056 , new_n8055 , n24032 );
and  g05708 ( new_n8057 , new_n8054 , new_n8056 );
nor  g05709 ( new_n8058 , new_n8053 , new_n8057 );
nor  g05710 ( new_n8059 , new_n8051 , new_n8058 );
nor  g05711 ( new_n8060 , new_n8049 , new_n8059 );
and  g05712 ( new_n8061 , new_n8047 , new_n8060 );
or   g05713 ( new_n8062 , new_n8046 , new_n8061 );
and  g05714 ( new_n8063 , new_n8044 , new_n8062 );
or   g05715 ( new_n8064 , new_n8043 , new_n8063 );
and  g05716 ( new_n8065 , new_n8041 , new_n8064 );
or   g05717 ( new_n8066 , new_n8040 , new_n8065 );
and  g05718 ( new_n8067_1 , new_n8038 , new_n8066 );
or   g05719 ( new_n8068 , new_n8037 , new_n8067_1 );
and  g05720 ( new_n8069 , new_n8035 , new_n8068 );
or   g05721 ( new_n8070 , new_n8034 , new_n8069 );
and  g05722 ( new_n8071 , new_n8032 , new_n8070 );
or   g05723 ( new_n8072 , new_n8031_1 , new_n8071 );
and  g05724 ( new_n8073 , new_n8030 , new_n8072 );
nor  g05725 ( new_n8074 , new_n8029 , new_n8073 );
not  g05726 ( new_n8075 , new_n8074 );
nor  g05727 ( new_n8076 , new_n8031_1 , new_n8071 );
xnor g05728 ( new_n8077 , new_n8030 , new_n8076 );
nor  g05729 ( new_n8078 , n1536 , new_n8077 );
not  g05730 ( new_n8079 , new_n8077 );
xnor g05731 ( new_n8080 , n1536 , new_n8079 );
xor  g05732 ( new_n8081 , new_n8032 , new_n8070 );
nor  g05733 ( new_n8082 , n19454 , new_n8081 );
xnor g05734 ( new_n8083 , n19454 , new_n8081 );
xor  g05735 ( new_n8084 , new_n8035 , new_n8068 );
nor  g05736 ( new_n8085 , n9445 , new_n8084 );
xnor g05737 ( new_n8086 , n9445 , new_n8084 );
xor  g05738 ( new_n8087 , new_n8038 , new_n8066 );
nor  g05739 ( new_n8088 , n1279 , new_n8087 );
xnor g05740 ( new_n8089 , n1279 , new_n8087 );
nor  g05741 ( new_n8090 , new_n8043 , new_n8063 );
xnor g05742 ( new_n8091 , new_n8041 , new_n8090 );
nor  g05743 ( new_n8092 , n8324 , new_n8091 );
not  g05744 ( new_n8093 , new_n8091 );
xnor g05745 ( new_n8094 , n8324 , new_n8093 );
xor  g05746 ( new_n8095_1 , new_n8044 , new_n8062 );
nor  g05747 ( new_n8096 , n12546 , new_n8095_1 );
xnor g05748 ( new_n8097 , n12546 , new_n8095_1 );
xnor g05749 ( new_n8098 , new_n8047 , new_n8060 );
not  g05750 ( new_n8099 , new_n8098 );
nor  g05751 ( new_n8100 , n21078 , new_n8099 );
xnor g05752 ( new_n8101 , n21078 , new_n8098 );
xnor g05753 ( new_n8102 , n2146 , n6785 );
xnor g05754 ( new_n8103_1 , new_n8058 , new_n8102 );
not  g05755 ( new_n8104 , new_n8103_1 );
and  g05756 ( new_n8105 , n24485 , new_n8104 );
or   g05757 ( new_n8106 , n24485 , new_n8104 );
xnor g05758 ( new_n8107 , n22173 , n24032 );
xnor g05759 ( new_n8108 , new_n8054 , new_n8107 );
nor  g05760 ( new_n8109_1 , n2420 , new_n8108 );
not  g05761 ( new_n8110 , n22201 );
or   g05762 ( new_n8111 , new_n8110 , new_n2545 );
not  g05763 ( new_n8112 , n2420 );
xnor g05764 ( new_n8113 , new_n8112 , new_n8108 );
and  g05765 ( new_n8114 , new_n8111 , new_n8113 );
nor  g05766 ( new_n8115 , new_n8109_1 , new_n8114 );
and  g05767 ( new_n8116 , new_n8106 , new_n8115 );
nor  g05768 ( new_n8117 , new_n8105 , new_n8116 );
and  g05769 ( new_n8118 , new_n8101 , new_n8117 );
nor  g05770 ( new_n8119 , new_n8100 , new_n8118 );
nor  g05771 ( new_n8120 , new_n8097 , new_n8119 );
or   g05772 ( new_n8121 , new_n8096 , new_n8120 );
and  g05773 ( new_n8122 , new_n8094 , new_n8121 );
nor  g05774 ( new_n8123 , new_n8092 , new_n8122 );
nor  g05775 ( new_n8124 , new_n8089 , new_n8123 );
nor  g05776 ( new_n8125 , new_n8088 , new_n8124 );
nor  g05777 ( new_n8126 , new_n8086 , new_n8125 );
nor  g05778 ( new_n8127_1 , new_n8085 , new_n8126 );
nor  g05779 ( new_n8128 , new_n8083 , new_n8127_1 );
or   g05780 ( new_n8129 , new_n8082 , new_n8128 );
and  g05781 ( new_n8130_1 , new_n8080 , new_n8129 );
nor  g05782 ( new_n8131 , new_n8078 , new_n8130_1 );
not  g05783 ( new_n8132 , new_n8131 );
nor  g05784 ( new_n8133 , new_n8075 , new_n8132 );
xnor g05785 ( new_n8134 , new_n8022 , new_n8026 );
xnor g05786 ( new_n8135_1 , new_n8074 , new_n8132 );
nor  g05787 ( new_n8136 , new_n8134 , new_n8135_1 );
xnor g05788 ( new_n8137 , new_n8134 , new_n8135_1 );
nor  g05789 ( new_n8138 , new_n7965 , new_n8019 );
xnor g05790 ( new_n8139_1 , new_n7962 , new_n8138 );
xor  g05791 ( new_n8140 , new_n8080 , new_n8129 );
and  g05792 ( new_n8141 , new_n8139_1 , new_n8140 );
xnor g05793 ( new_n8142 , new_n8139_1 , new_n8140 );
xor  g05794 ( new_n8143 , new_n7967 , new_n8018 );
not  g05795 ( new_n8144 , new_n8143 );
xnor g05796 ( new_n8145 , new_n8083 , new_n8127_1 );
nor  g05797 ( new_n8146 , new_n8144 , new_n8145 );
xnor g05798 ( new_n8147 , new_n8144 , new_n8145 );
xor  g05799 ( new_n8148_1 , new_n7972 , new_n8016 );
not  g05800 ( new_n8149_1 , new_n8148_1 );
xnor g05801 ( new_n8150 , new_n8086 , new_n8125 );
nor  g05802 ( new_n8151 , new_n8149_1 , new_n8150 );
xnor g05803 ( new_n8152 , new_n8149_1 , new_n8150 );
xor  g05804 ( new_n8153 , new_n7977 , new_n8014 );
not  g05805 ( new_n8154 , new_n8153 );
xnor g05806 ( new_n8155 , new_n8089 , new_n8123 );
nor  g05807 ( new_n8156 , new_n8154 , new_n8155 );
xnor g05808 ( new_n8157 , new_n8154 , new_n8155 );
nor  g05809 ( new_n8158 , new_n7985 , new_n8011 );
xnor g05810 ( new_n8159_1 , new_n7982 , new_n8158 );
xor  g05811 ( new_n8160 , new_n8094 , new_n8121 );
and  g05812 ( new_n8161 , new_n8159_1 , new_n8160 );
xnor g05813 ( new_n8162 , new_n8159_1 , new_n8160 );
xor  g05814 ( new_n8163 , new_n7987 , new_n8010 );
not  g05815 ( new_n8164 , new_n8163 );
xnor g05816 ( new_n8165 , new_n8097 , new_n8119 );
nor  g05817 ( new_n8166 , new_n8164 , new_n8165 );
xnor g05818 ( new_n8167 , new_n8164 , new_n8165 );
xnor g05819 ( new_n8168 , new_n7992_1 , new_n8008 );
xnor g05820 ( new_n8169 , new_n8101 , new_n8117 );
nor  g05821 ( new_n8170 , new_n8168 , new_n8169 );
xnor g05822 ( new_n8171 , new_n8168 , new_n8169 );
xnor g05823 ( new_n8172 , new_n7997 , new_n8006_1 );
not  g05824 ( new_n8173 , new_n8172 );
xnor g05825 ( new_n8174 , n24485 , new_n8104 );
xnor g05826 ( new_n8175 , new_n8115 , new_n8174 );
nor  g05827 ( new_n8176 , new_n8173 , new_n8175 );
xnor g05828 ( new_n8177 , new_n8172 , new_n8175 );
xor  g05829 ( new_n8178 , new_n8111 , new_n8113 );
xnor g05830 ( new_n8179_1 , new_n8002 , new_n8004 );
nor  g05831 ( new_n8180 , new_n8178 , new_n8179_1 );
not  g05832 ( new_n8181 , new_n2544 );
and  g05833 ( new_n8182 , new_n8181 , new_n2546 );
not  g05834 ( new_n8183 , new_n8179_1 );
xnor g05835 ( new_n8184 , new_n8178 , new_n8183 );
and  g05836 ( new_n8185 , new_n8182 , new_n8184 );
nor  g05837 ( new_n8186 , new_n8180 , new_n8185 );
and  g05838 ( new_n8187 , new_n8177 , new_n8186 );
nor  g05839 ( new_n8188 , new_n8176 , new_n8187 );
nor  g05840 ( new_n8189 , new_n8171 , new_n8188 );
nor  g05841 ( new_n8190 , new_n8170 , new_n8189 );
nor  g05842 ( new_n8191 , new_n8167 , new_n8190 );
nor  g05843 ( new_n8192 , new_n8166 , new_n8191 );
nor  g05844 ( new_n8193 , new_n8162 , new_n8192 );
nor  g05845 ( new_n8194_1 , new_n8161 , new_n8193 );
nor  g05846 ( new_n8195 , new_n8157 , new_n8194_1 );
nor  g05847 ( new_n8196 , new_n8156 , new_n8195 );
nor  g05848 ( new_n8197 , new_n8152 , new_n8196 );
nor  g05849 ( new_n8198 , new_n8151 , new_n8197 );
nor  g05850 ( new_n8199 , new_n8147 , new_n8198 );
nor  g05851 ( new_n8200 , new_n8146 , new_n8199 );
nor  g05852 ( new_n8201 , new_n8142 , new_n8200 );
nor  g05853 ( new_n8202 , new_n8141 , new_n8201 );
nor  g05854 ( new_n8203 , new_n8137 , new_n8202 );
nor  g05855 ( new_n8204 , new_n8136 , new_n8203 );
xor  g05856 ( new_n8205 , new_n8133 , new_n8204 );
xnor g05857 ( n849 , new_n8028 , new_n8205 );
xnor g05858 ( n858 , new_n2529 , new_n2530 );
nor  g05859 ( new_n8208 , n9246 , n16994 );
not  g05860 ( new_n8209 , new_n8208 );
nor  g05861 ( new_n8210 , n10096 , new_n8209 );
not  g05862 ( new_n8211 , new_n8210 );
nor  g05863 ( new_n8212 , n14790 , new_n8211 );
not  g05864 ( new_n8213 , new_n8212 );
nor  g05865 ( new_n8214 , n17251 , new_n8213 );
not  g05866 ( new_n8215_1 , new_n8214 );
nor  g05867 ( new_n8216 , n21674 , new_n8215_1 );
not  g05868 ( new_n8217 , new_n8216 );
nor  g05869 ( new_n8218 , n24638 , new_n8217 );
not  g05870 ( new_n8219 , new_n8218 );
nor  g05871 ( new_n8220 , n18444 , new_n8219 );
not  g05872 ( new_n8221 , new_n8220 );
nor  g05873 ( new_n8222 , n14899 , new_n8221 );
xnor g05874 ( new_n8223 , n3506 , new_n8222 );
xnor g05875 ( new_n8224 , n1314 , new_n8223 );
xnor g05876 ( new_n8225 , n14899 , new_n8220 );
and  g05877 ( new_n8226 , n3306 , new_n8225 );
or   g05878 ( new_n8227 , n3306 , new_n8225 );
xnor g05879 ( new_n8228 , n18444 , new_n8218 );
nor  g05880 ( new_n8229 , n22335 , new_n8228 );
not  g05881 ( new_n8230 , n22335 );
xnor g05882 ( new_n8231 , new_n8230 , new_n8228 );
xnor g05883 ( new_n8232 , n24638 , new_n8216 );
nor  g05884 ( new_n8233 , n24048 , new_n8232 );
not  g05885 ( new_n8234 , n24048 );
xnor g05886 ( new_n8235 , new_n8234 , new_n8232 );
xnor g05887 ( new_n8236 , n21674 , new_n8214 );
nor  g05888 ( new_n8237 , n1525 , new_n8236 );
not  g05889 ( new_n8238 , n1525 );
xnor g05890 ( new_n8239 , new_n8238 , new_n8236 );
xnor g05891 ( new_n8240 , n17251 , new_n8212 );
nor  g05892 ( new_n8241 , n16988 , new_n8240 );
xnor g05893 ( new_n8242 , new_n4638 , new_n8240 );
xnor g05894 ( new_n8243 , n14790 , new_n8210 );
nor  g05895 ( new_n8244_1 , n21779 , new_n8243 );
xnor g05896 ( new_n8245 , n10096 , new_n8208 );
nor  g05897 ( new_n8246 , n5376 , new_n8245 );
xnor g05898 ( new_n8247 , new_n4645 , new_n8245 );
xnor g05899 ( new_n8248 , n9246 , n16994 );
and  g05900 ( new_n8249 , new_n4648 , new_n8248 );
and  g05901 ( new_n8250 , n9246 , n23120 );
xnor g05902 ( new_n8251 , new_n4648 , new_n8248 );
nor  g05903 ( new_n8252 , new_n8250 , new_n8251 );
or   g05904 ( new_n8253 , new_n8249 , new_n8252 );
and  g05905 ( new_n8254 , new_n8247 , new_n8253 );
or   g05906 ( new_n8255_1 , new_n8246 , new_n8254 );
xnor g05907 ( new_n8256_1 , new_n4641 , new_n8243 );
and  g05908 ( new_n8257 , new_n8255_1 , new_n8256_1 );
or   g05909 ( new_n8258 , new_n8244_1 , new_n8257 );
and  g05910 ( new_n8259_1 , new_n8242 , new_n8258 );
or   g05911 ( new_n8260 , new_n8241 , new_n8259_1 );
and  g05912 ( new_n8261 , new_n8239 , new_n8260 );
or   g05913 ( new_n8262 , new_n8237 , new_n8261 );
and  g05914 ( new_n8263 , new_n8235 , new_n8262 );
or   g05915 ( new_n8264 , new_n8233 , new_n8263 );
and  g05916 ( new_n8265 , new_n8231 , new_n8264 );
nor  g05917 ( new_n8266 , new_n8229 , new_n8265 );
and  g05918 ( new_n8267_1 , new_n8227 , new_n8266 );
nor  g05919 ( new_n8268 , new_n8226 , new_n8267_1 );
xnor g05920 ( new_n8269 , new_n8224 , new_n8268 );
nor  g05921 ( new_n8270 , n22442 , new_n8269 );
not  g05922 ( new_n8271 , n22442 );
xnor g05923 ( new_n8272 , new_n8271 , new_n8269 );
not  g05924 ( new_n8273 , n468 );
xnor g05925 ( new_n8274 , n3306 , new_n8225 );
xnor g05926 ( new_n8275 , new_n8266 , new_n8274 );
nor  g05927 ( new_n8276_1 , new_n8273 , new_n8275 );
xnor g05928 ( new_n8277 , n468 , new_n8275 );
xor  g05929 ( new_n8278 , new_n8231 , new_n8264 );
nor  g05930 ( new_n8279 , n5400 , new_n8278 );
not  g05931 ( new_n8280 , n5400 );
xnor g05932 ( new_n8281 , new_n8280 , new_n8278 );
xor  g05933 ( new_n8282 , new_n8235 , new_n8262 );
nor  g05934 ( new_n8283 , n23923 , new_n8282 );
not  g05935 ( new_n8284 , n23923 );
xnor g05936 ( new_n8285_1 , new_n8284 , new_n8282 );
xor  g05937 ( new_n8286 , new_n8239 , new_n8260 );
and  g05938 ( new_n8287 , n329 , new_n8286 );
or   g05939 ( new_n8288_1 , n329 , new_n8286 );
xor  g05940 ( new_n8289 , new_n8255_1 , new_n8256_1 );
nor  g05941 ( new_n8290 , n2409 , new_n8289 );
xnor g05942 ( new_n8291 , n2409 , new_n8289 );
xor  g05943 ( new_n8292 , new_n8247 , new_n8253 );
nor  g05944 ( new_n8293 , n8869 , new_n8292 );
xor  g05945 ( new_n8294 , new_n8250 , new_n8251 );
nor  g05946 ( new_n8295 , n10372 , new_n8294 );
xnor g05947 ( new_n8296 , new_n3562 , n23120 );
nor  g05948 ( new_n8297 , new_n7024 , new_n8296 );
xnor g05949 ( new_n8298 , n10372 , new_n8294 );
nor  g05950 ( new_n8299 , new_n8297 , new_n8298 );
nor  g05951 ( new_n8300 , new_n8295 , new_n8299 );
xnor g05952 ( new_n8301 , n8869 , new_n8292 );
nor  g05953 ( new_n8302 , new_n8300 , new_n8301 );
nor  g05954 ( new_n8303 , new_n8293 , new_n8302 );
nor  g05955 ( new_n8304 , new_n8291 , new_n8303 );
nor  g05956 ( new_n8305_1 , new_n8290 , new_n8304 );
nor  g05957 ( new_n8306_1 , n24170 , new_n8305_1 );
xor  g05958 ( new_n8307 , new_n8242 , new_n8258 );
xnor g05959 ( new_n8308 , n24170 , new_n8305_1 );
nor  g05960 ( new_n8309_1 , new_n8307 , new_n8308 );
nor  g05961 ( new_n8310 , new_n8306_1 , new_n8309_1 );
and  g05962 ( new_n8311 , new_n8288_1 , new_n8310 );
nor  g05963 ( new_n8312 , new_n8287 , new_n8311 );
and  g05964 ( new_n8313 , new_n8285_1 , new_n8312 );
or   g05965 ( new_n8314 , new_n8283 , new_n8313 );
and  g05966 ( new_n8315 , new_n8281 , new_n8314 );
nor  g05967 ( new_n8316 , new_n8279 , new_n8315 );
and  g05968 ( new_n8317 , new_n8277 , new_n8316 );
nor  g05969 ( new_n8318 , new_n8276_1 , new_n8317 );
and  g05970 ( new_n8319 , new_n8272 , new_n8318 );
nor  g05971 ( new_n8320_1 , new_n8270 , new_n8319 );
nor  g05972 ( new_n8321_1 , n1314 , new_n8223 );
nor  g05973 ( new_n8322 , new_n8321_1 , new_n8268 );
not  g05974 ( new_n8323 , n3506 );
and  g05975 ( new_n8324_1 , new_n8323 , new_n8222 );
and  g05976 ( new_n8325 , n1314 , new_n8223 );
or   g05977 ( new_n8326 , new_n8324_1 , new_n8325 );
nor  g05978 ( new_n8327 , new_n8322 , new_n8326 );
xor  g05979 ( new_n8328 , new_n8320_1 , new_n8327 );
not  g05980 ( new_n8329 , new_n8328 );
nor  g05981 ( new_n8330 , n26180 , new_n3472 );
nor  g05982 ( new_n8331 , new_n3473 , new_n3534 );
nor  g05983 ( new_n8332 , new_n8330 , new_n8331 );
not  g05984 ( new_n8333 , new_n8332 );
and  g05985 ( new_n8334 , new_n7608 , new_n3419 );
nor  g05986 ( new_n8335 , n25494 , new_n3420 );
and  g05987 ( new_n8336 , n25494 , new_n3420 );
nor  g05988 ( new_n8337 , new_n8336 , new_n3471 );
nor  g05989 ( new_n8338 , new_n8335 , new_n8337 );
nor  g05990 ( new_n8339_1 , new_n8334 , new_n8338 );
xnor g05991 ( new_n8340 , new_n8333 , new_n8339_1 );
xnor g05992 ( new_n8341 , new_n8329 , new_n8340 );
xor  g05993 ( new_n8342 , new_n8272 , new_n8318 );
nor  g05994 ( new_n8343 , new_n3535 , new_n8342 );
xnor g05995 ( new_n8344 , new_n3535 , new_n8342 );
xor  g05996 ( new_n8345 , new_n8277 , new_n8316 );
and  g05997 ( new_n8346 , new_n3665_1 , new_n8345 );
xnor g05998 ( new_n8347 , new_n3665_1 , new_n8345 );
xor  g05999 ( new_n8348 , new_n8281 , new_n8314 );
nor  g06000 ( new_n8349 , new_n3671 , new_n8348 );
xnor g06001 ( new_n8350 , new_n3671 , new_n8348 );
xor  g06002 ( new_n8351 , new_n8285_1 , new_n8312 );
nor  g06003 ( new_n8352 , new_n3676 , new_n8351 );
not  g06004 ( new_n8353 , n329 );
xnor g06005 ( new_n8354 , new_n8353 , new_n8286 );
xnor g06006 ( new_n8355 , new_n8310 , new_n8354 );
nor  g06007 ( new_n8356 , new_n3681 , new_n8355 );
xnor g06008 ( new_n8357 , new_n3681 , new_n8355 );
xor  g06009 ( new_n8358 , new_n8307 , new_n8308 );
nor  g06010 ( new_n8359 , new_n3686 , new_n8358 );
xor  g06011 ( new_n8360 , new_n8291 , new_n8303 );
nor  g06012 ( new_n8361 , new_n3690 , new_n8360 );
xnor g06013 ( new_n8362 , new_n3690 , new_n8360 );
xor  g06014 ( new_n8363_1 , new_n8300 , new_n8301 );
nor  g06015 ( new_n8364 , new_n3696 , new_n8363_1 );
xor  g06016 ( new_n8365 , new_n8297 , new_n8298 );
nor  g06017 ( new_n8366 , new_n3702 , new_n8365 );
not  g06018 ( new_n8367 , new_n3704 );
xnor g06019 ( new_n8368 , n7428 , new_n8296 );
nor  g06020 ( new_n8369 , new_n8367 , new_n8368 );
xnor g06021 ( new_n8370 , new_n3702 , new_n8365 );
nor  g06022 ( new_n8371 , new_n8369 , new_n8370 );
nor  g06023 ( new_n8372 , new_n8366 , new_n8371 );
xnor g06024 ( new_n8373 , new_n3696 , new_n8363_1 );
nor  g06025 ( new_n8374 , new_n8372 , new_n8373 );
nor  g06026 ( new_n8375 , new_n8364 , new_n8374 );
nor  g06027 ( new_n8376_1 , new_n8362 , new_n8375 );
nor  g06028 ( new_n8377 , new_n8361 , new_n8376_1 );
xnor g06029 ( new_n8378 , new_n3686 , new_n8358 );
nor  g06030 ( new_n8379 , new_n8377 , new_n8378 );
nor  g06031 ( new_n8380 , new_n8359 , new_n8379 );
nor  g06032 ( new_n8381_1 , new_n8357 , new_n8380 );
nor  g06033 ( new_n8382 , new_n8356 , new_n8381_1 );
xnor g06034 ( new_n8383 , new_n3676 , new_n8351 );
nor  g06035 ( new_n8384 , new_n8382 , new_n8383 );
nor  g06036 ( new_n8385 , new_n8352 , new_n8384 );
nor  g06037 ( new_n8386 , new_n8350 , new_n8385 );
nor  g06038 ( new_n8387 , new_n8349 , new_n8386 );
nor  g06039 ( new_n8388 , new_n8347 , new_n8387 );
nor  g06040 ( new_n8389 , new_n8346 , new_n8388 );
nor  g06041 ( new_n8390 , new_n8344 , new_n8389 );
or   g06042 ( new_n8391 , new_n8343 , new_n8390 );
xnor g06043 ( n873 , new_n8341 , new_n8391 );
xnor g06044 ( new_n8393 , n2731 , n4812 );
not  g06045 ( new_n8394 , n24278 );
nor  g06046 ( new_n8395 , n19911 , new_n8394 );
xnor g06047 ( new_n8396 , n19911 , n24278 );
nor  g06048 ( new_n8397 , new_n2389 , n24618 );
not  g06049 ( new_n8398 , n24618 );
nor  g06050 ( new_n8399_1 , n13708 , new_n8398 );
nor  g06051 ( new_n8400 , n3952 , new_n3826 );
nor  g06052 ( new_n8401 , new_n2443 , n18409 );
nor  g06053 ( new_n8402 , new_n2381 , n12315 );
not  g06054 ( new_n8403 , new_n8402 );
nor  g06055 ( new_n8404 , new_n8401 , new_n8403 );
nor  g06056 ( new_n8405_1 , new_n8400 , new_n8404 );
nor  g06057 ( new_n8406 , new_n8399_1 , new_n8405_1 );
nor  g06058 ( new_n8407 , new_n8397 , new_n8406 );
and  g06059 ( new_n8408_1 , new_n8396 , new_n8407 );
or   g06060 ( new_n8409 , new_n8395 , new_n8408_1 );
xor  g06061 ( new_n8410 , new_n8393 , new_n8409 );
xor  g06062 ( new_n8411 , new_n5187 , new_n8410 );
xnor g06063 ( new_n8412 , new_n8396 , new_n8407 );
and  g06064 ( new_n8413 , new_n5191 , new_n8412 );
xnor g06065 ( new_n8414 , n13708 , n24618 );
xnor g06066 ( new_n8415 , new_n8405_1 , new_n8414 );
nor  g06067 ( new_n8416 , new_n5195 , new_n8415 );
xnor g06068 ( new_n8417_1 , new_n5195 , new_n8415 );
xnor g06069 ( new_n8418 , n5704 , n12315 );
nor  g06070 ( new_n8419 , new_n5202 , new_n8418 );
and  g06071 ( new_n8420 , new_n5207 , new_n8419 );
xnor g06072 ( new_n8421 , new_n5207 , new_n8419 );
xnor g06073 ( new_n8422 , n3952 , n18409 );
xnor g06074 ( new_n8423 , new_n8403 , new_n8422 );
nor  g06075 ( new_n8424 , new_n8421 , new_n8423 );
nor  g06076 ( new_n8425 , new_n8420 , new_n8424 );
nor  g06077 ( new_n8426 , new_n8417_1 , new_n8425 );
nor  g06078 ( new_n8427 , new_n8416 , new_n8426 );
xnor g06079 ( new_n8428 , new_n5190 , new_n8412 );
and  g06080 ( new_n8429 , new_n8427 , new_n8428 );
nor  g06081 ( new_n8430 , new_n8413 , new_n8429 );
xor  g06082 ( n879 , new_n8411 , new_n8430 );
not  g06083 ( new_n8432_1 , n18157 );
xnor g06084 ( new_n8433 , new_n8432_1 , new_n7991 );
nor  g06085 ( new_n8434 , n12161 , new_n7995 );
nor  g06086 ( new_n8435 , new_n7220 , new_n8002 );
nor  g06087 ( new_n8436 , new_n6628_1 , new_n2543 );
xnor g06088 ( new_n8437 , new_n7220 , new_n8003 );
and  g06089 ( new_n8438 , new_n8436 , new_n8437 );
nor  g06090 ( new_n8439_1 , new_n8435 , new_n8438 );
xnor g06091 ( new_n8440 , new_n7217 , new_n7995 );
and  g06092 ( new_n8441 , new_n8439_1 , new_n8440 );
nor  g06093 ( new_n8442 , new_n8434 , new_n8441 );
xnor g06094 ( new_n8443 , new_n8433 , new_n8442 );
xnor g06095 ( new_n8444 , new_n8439_1 , new_n8440 );
not  g06096 ( new_n8445 , n14684 );
xnor g06097 ( new_n8446 , new_n8445 , new_n6610 );
nor  g06098 ( new_n8447 , n6631 , new_n6612_1 );
or   g06099 ( new_n8448 , new_n4183 , new_n6614 );
xnor g06100 ( new_n8449 , new_n4180 , new_n6612_1 );
and  g06101 ( new_n8450 , new_n8448 , new_n8449 );
or   g06102 ( new_n8451 , new_n8447 , new_n8450 );
xor  g06103 ( new_n8452 , new_n8446 , new_n8451 );
nor  g06104 ( new_n8453_1 , new_n8444 , new_n8452 );
xnor g06105 ( new_n8454 , new_n8444 , new_n8452 );
xor  g06106 ( new_n8455 , new_n8448 , new_n8449 );
xor  g06107 ( new_n8456 , new_n8436 , new_n8437 );
nor  g06108 ( new_n8457 , new_n8455 , new_n8456 );
xnor g06109 ( new_n8458 , n24732 , new_n6614 );
not  g06110 ( new_n8459 , new_n8458 );
xnor g06111 ( new_n8460 , n8581 , new_n2543 );
nor  g06112 ( new_n8461 , new_n8459 , new_n8460 );
xnor g06113 ( new_n8462 , new_n8455 , new_n8456 );
not  g06114 ( new_n8463 , new_n8462 );
and  g06115 ( new_n8464 , new_n8461 , new_n8463 );
nor  g06116 ( new_n8465 , new_n8457 , new_n8464 );
nor  g06117 ( new_n8466 , new_n8454 , new_n8465 );
nor  g06118 ( new_n8467 , new_n8453_1 , new_n8466 );
xnor g06119 ( new_n8468 , new_n8443 , new_n8467 );
not  g06120 ( new_n8469 , n17035 );
xnor g06121 ( new_n8470 , new_n8469 , new_n6604 );
nor  g06122 ( new_n8471 , n14684 , new_n6610 );
and  g06123 ( new_n8472 , new_n8446 , new_n8451 );
nor  g06124 ( new_n8473 , new_n8471 , new_n8472 );
xnor g06125 ( new_n8474 , new_n8470 , new_n8473 );
xor  g06126 ( n887 , new_n8468 , new_n8474 );
xnor g06127 ( new_n8476 , new_n4917 , new_n6041 );
nor  g06128 ( new_n8477 , new_n4922 , new_n6045 );
xnor g06129 ( new_n8478 , new_n4922 , new_n6047 );
nor  g06130 ( new_n8479 , new_n4927 , new_n6051 );
xnor g06131 ( new_n8480_1 , new_n4927 , new_n6053 );
nor  g06132 ( new_n8481 , new_n4932 , new_n6057 );
xnor g06133 ( new_n8482 , new_n4932 , new_n6059 );
not  g06134 ( new_n8483 , n25872 );
nor  g06135 ( new_n8484 , new_n8483 , new_n6063 );
nor  g06136 ( new_n8485 , n20259 , new_n6065 );
or   g06137 ( new_n8486 , new_n5002 , new_n5792 );
xnor g06138 ( new_n8487 , new_n4939_1 , new_n6065 );
and  g06139 ( new_n8488 , new_n8486 , new_n8487 );
nor  g06140 ( new_n8489_1 , new_n8485 , new_n8488 );
xnor g06141 ( new_n8490 , new_n8483 , new_n6072 );
and  g06142 ( new_n8491 , new_n8489_1 , new_n8490 );
or   g06143 ( new_n8492 , new_n8484 , new_n8491 );
and  g06144 ( new_n8493 , new_n8482 , new_n8492 );
or   g06145 ( new_n8494 , new_n8481 , new_n8493 );
and  g06146 ( new_n8495 , new_n8480_1 , new_n8494 );
or   g06147 ( new_n8496 , new_n8479 , new_n8495 );
and  g06148 ( new_n8497 , new_n8478 , new_n8496 );
nor  g06149 ( new_n8498 , new_n8477 , new_n8497 );
xnor g06150 ( new_n8499 , new_n8476 , new_n8498 );
not  g06151 ( new_n8500 , new_n8499 );
not  g06152 ( new_n8501 , n25119 );
xnor g06153 ( new_n8502 , new_n8501 , new_n2980 );
not  g06154 ( new_n8503 , n1163 );
nor  g06155 ( new_n8504 , new_n8503 , new_n2985_1 );
nor  g06156 ( new_n8505_1 , n18537 , new_n2990 );
not  g06157 ( new_n8506 , n18537 );
xnor g06158 ( new_n8507 , new_n8506 , new_n2990 );
nor  g06159 ( new_n8508 , n7057 , new_n2996 );
xor  g06160 ( new_n8509 , n7057 , new_n2996 );
not  g06161 ( new_n8510_1 , n8381 );
nor  g06162 ( new_n8511 , new_n8510_1 , new_n3002 );
xnor g06163 ( new_n8512 , n8381 , new_n3002 );
nor  g06164 ( new_n8513 , new_n5080 , new_n3063 );
nor  g06165 ( new_n8514 , n20235 , new_n8513 );
xnor g06166 ( new_n8515 , new_n5040 , new_n8513 );
and  g06167 ( new_n8516 , new_n3008 , new_n8515 );
nor  g06168 ( new_n8517 , new_n8514 , new_n8516 );
and  g06169 ( new_n8518 , new_n8512 , new_n8517 );
nor  g06170 ( new_n8519_1 , new_n8511 , new_n8518 );
and  g06171 ( new_n8520 , new_n8509 , new_n8519_1 );
or   g06172 ( new_n8521 , new_n8508 , new_n8520 );
and  g06173 ( new_n8522 , new_n8507 , new_n8521 );
nor  g06174 ( new_n8523 , new_n8505_1 , new_n8522 );
xnor g06175 ( new_n8524 , new_n8503 , new_n2986 );
and  g06176 ( new_n8525 , new_n8523 , new_n8524 );
nor  g06177 ( new_n8526_1 , new_n8504 , new_n8525 );
xnor g06178 ( new_n8527 , new_n8502 , new_n8526_1 );
xnor g06179 ( new_n8528 , new_n8500 , new_n8527 );
nor  g06180 ( new_n8529 , new_n8479 , new_n8495 );
xnor g06181 ( new_n8530 , new_n8478 , new_n8529 );
not  g06182 ( new_n8531 , new_n8530 );
xor  g06183 ( new_n8532 , new_n8523 , new_n8524 );
nor  g06184 ( new_n8533 , new_n8531 , new_n8532 );
xnor g06185 ( new_n8534 , new_n8531 , new_n8532 );
xor  g06186 ( new_n8535_1 , new_n8507 , new_n8521 );
nor  g06187 ( new_n8536 , new_n8481 , new_n8493 );
xnor g06188 ( new_n8537 , new_n8480_1 , new_n8536 );
and  g06189 ( new_n8538 , new_n8535_1 , new_n8537 );
xnor g06190 ( new_n8539 , new_n8535_1 , new_n8537 );
xnor g06191 ( new_n8540 , new_n8509 , new_n8519_1 );
nor  g06192 ( new_n8541 , new_n8484 , new_n8491 );
xnor g06193 ( new_n8542 , new_n8482 , new_n8541 );
not  g06194 ( new_n8543 , new_n8542 );
nor  g06195 ( new_n8544 , new_n8540 , new_n8543 );
xnor g06196 ( new_n8545 , new_n8540 , new_n8543 );
xnor g06197 ( new_n8546 , new_n8512 , new_n8517 );
xnor g06198 ( new_n8547 , new_n8489_1 , new_n8490 );
not  g06199 ( new_n8548 , new_n8547 );
and  g06200 ( new_n8549 , new_n8546 , new_n8548 );
xnor g06201 ( new_n8550_1 , new_n8546 , new_n8548 );
nor  g06202 ( new_n8551 , new_n5002 , new_n5792 );
xnor g06203 ( new_n8552 , new_n8551 , new_n8487 );
not  g06204 ( new_n8553 , new_n8552 );
xnor g06205 ( new_n8554 , new_n3009 , new_n8515 );
and  g06206 ( new_n8555 , new_n8553 , new_n8554 );
xnor g06207 ( new_n8556 , n3925 , new_n5792 );
not  g06208 ( new_n8557 , new_n8556 );
xnor g06209 ( new_n8558 , n12495 , new_n3063 );
nor  g06210 ( new_n8559 , new_n8557 , new_n8558 );
xnor g06211 ( new_n8560 , new_n8552 , new_n8554 );
and  g06212 ( new_n8561 , new_n8559 , new_n8560 );
nor  g06213 ( new_n8562 , new_n8555 , new_n8561 );
nor  g06214 ( new_n8563_1 , new_n8550_1 , new_n8562 );
nor  g06215 ( new_n8564 , new_n8549 , new_n8563_1 );
nor  g06216 ( new_n8565 , new_n8545 , new_n8564 );
nor  g06217 ( new_n8566 , new_n8544 , new_n8565 );
nor  g06218 ( new_n8567 , new_n8539 , new_n8566 );
nor  g06219 ( new_n8568 , new_n8538 , new_n8567 );
nor  g06220 ( new_n8569 , new_n8534 , new_n8568 );
nor  g06221 ( new_n8570 , new_n8533 , new_n8569 );
xnor g06222 ( n904 , new_n8528 , new_n8570 );
not  g06223 ( new_n8572 , n19472 );
nor  g06224 ( new_n8573 , n10158 , n18962 );
not  g06225 ( new_n8574 , new_n8573 );
nor  g06226 ( new_n8575 , n8052 , new_n8574 );
not  g06227 ( new_n8576 , new_n8575 );
nor  g06228 ( new_n8577 , n15539 , new_n8576 );
xnor g06229 ( new_n8578 , n19228 , new_n8577 );
xnor g06230 ( new_n8579 , n21471 , new_n8578 );
xnor g06231 ( new_n8580 , n15539 , new_n8575 );
and  g06232 ( new_n8581_1 , n18737 , new_n8580 );
xnor g06233 ( new_n8582 , n18737 , new_n8580 );
xnor g06234 ( new_n8583 , n8052 , new_n8573 );
not  g06235 ( new_n8584 , new_n8583 );
nor  g06236 ( new_n8585 , new_n3301_1 , new_n8584 );
xnor g06237 ( new_n8586 , n14603 , new_n8584 );
xnor g06238 ( new_n8587 , n10158 , n18962 );
not  g06239 ( new_n8588 , new_n8587 );
nor  g06240 ( new_n8589 , n20794 , new_n8588 );
nor  g06241 ( new_n8590 , new_n6771 , new_n3305 );
xnor g06242 ( new_n8591 , n20794 , new_n8587 );
not  g06243 ( new_n8592 , new_n8591 );
nor  g06244 ( new_n8593 , new_n8590 , new_n8592 );
nor  g06245 ( new_n8594_1 , new_n8589 , new_n8593 );
and  g06246 ( new_n8595 , new_n8586 , new_n8594_1 );
nor  g06247 ( new_n8596 , new_n8585 , new_n8595 );
nor  g06248 ( new_n8597 , new_n8582 , new_n8596 );
nor  g06249 ( new_n8598 , new_n8581_1 , new_n8597 );
xnor g06250 ( new_n8599 , new_n8579 , new_n8598 );
not  g06251 ( new_n8600 , new_n8599 );
xnor g06252 ( new_n8601 , new_n8572 , new_n8600 );
xnor g06253 ( new_n8602 , new_n8582 , new_n8596 );
not  g06254 ( new_n8603 , new_n8602 );
nor  g06255 ( new_n8604 , n25370 , new_n8603 );
not  g06256 ( new_n8605 , n24786 );
xnor g06257 ( new_n8606 , new_n8586 , new_n8594_1 );
nor  g06258 ( new_n8607 , new_n8605 , new_n8606 );
not  g06259 ( new_n8608_1 , new_n8606 );
xnor g06260 ( new_n8609 , new_n8605 , new_n8608_1 );
xnor g06261 ( new_n8610 , n18962 , n23333 );
nor  g06262 ( new_n8611 , new_n4109 , new_n8610 );
and  g06263 ( new_n8612 , new_n8591 , new_n8611 );
xnor g06264 ( new_n8613 , new_n8590 , new_n8592 );
nor  g06265 ( new_n8614_1 , new_n8611 , new_n8613 );
nor  g06266 ( new_n8615 , new_n8612 , new_n8614_1 );
and  g06267 ( new_n8616 , n27120 , new_n8615 );
or   g06268 ( new_n8617 , new_n8612 , new_n8616 );
and  g06269 ( new_n8618 , new_n8609 , new_n8617 );
nor  g06270 ( new_n8619 , new_n8607 , new_n8618 );
xnor g06271 ( new_n8620_1 , new_n6846 , new_n8603 );
and  g06272 ( new_n8621 , new_n8619 , new_n8620_1 );
nor  g06273 ( new_n8622 , new_n8604 , new_n8621 );
xor  g06274 ( new_n8623 , new_n8601 , new_n8622 );
xnor g06275 ( new_n8624 , new_n6696 , new_n8623 );
xnor g06276 ( new_n8625 , new_n8619 , new_n8620_1 );
nor  g06277 ( new_n8626 , new_n6699 , new_n8625 );
xnor g06278 ( new_n8627 , new_n6699 , new_n8625 );
not  g06279 ( new_n8628 , n27120 );
xnor g06280 ( new_n8629 , new_n8628 , new_n8615 );
nor  g06281 ( new_n8630 , new_n6731 , new_n8629 );
xnor g06282 ( new_n8631 , n23065 , new_n8610 );
not  g06283 ( new_n8632 , new_n8631 );
nor  g06284 ( new_n8633 , new_n6702 , new_n8632 );
xnor g06285 ( new_n8634 , new_n6731 , new_n8629 );
nor  g06286 ( new_n8635 , new_n8633 , new_n8634 );
nor  g06287 ( new_n8636 , new_n8630 , new_n8635 );
nor  g06288 ( new_n8637_1 , new_n6715 , new_n8636 );
xor  g06289 ( new_n8638_1 , new_n8609 , new_n8617 );
xnor g06290 ( new_n8639 , new_n6715 , new_n8636 );
nor  g06291 ( new_n8640 , new_n8638_1 , new_n8639 );
nor  g06292 ( new_n8641 , new_n8637_1 , new_n8640 );
nor  g06293 ( new_n8642 , new_n8627 , new_n8641 );
nor  g06294 ( new_n8643 , new_n8626 , new_n8642 );
xnor g06295 ( n948 , new_n8624 , new_n8643 );
xnor g06296 ( new_n8645 , n10250 , n25972 );
not  g06297 ( new_n8646 , n21915 );
nor  g06298 ( new_n8647 , n7674 , new_n8646 );
xnor g06299 ( new_n8648 , n7674 , n21915 );
nor  g06300 ( new_n8649 , n6397 , new_n6836 );
xnor g06301 ( new_n8650 , n6397 , n13775 );
nor  g06302 ( new_n8651 , new_n6839 , n19196 );
xnor g06303 ( new_n8652 , n1293 , n19196 );
nor  g06304 ( new_n8653 , new_n6842 , n23586 );
xnor g06305 ( new_n8654 , n19042 , n23586 );
nor  g06306 ( new_n8655 , new_n8572 , n21226 );
xnor g06307 ( new_n8656_1 , n19472 , n21226 );
nor  g06308 ( new_n8657 , n4426 , new_n6846 );
xnor g06309 ( new_n8658 , n4426 , n25370 );
not  g06310 ( new_n8659 , n20036 );
nor  g06311 ( new_n8660 , new_n8659 , n24786 );
nor  g06312 ( new_n8661 , n20036 , new_n8605 );
nor  g06313 ( new_n8662_1 , new_n4120 , n27120 );
or   g06314 ( new_n8663 , n11192 , new_n8628 );
nor  g06315 ( new_n8664 , new_n6176 , n23065 );
and  g06316 ( new_n8665 , new_n8663 , new_n8664 );
nor  g06317 ( new_n8666 , new_n8662_1 , new_n8665 );
nor  g06318 ( new_n8667 , new_n8661 , new_n8666 );
nor  g06319 ( new_n8668 , new_n8660 , new_n8667 );
and  g06320 ( new_n8669 , new_n8658 , new_n8668 );
or   g06321 ( new_n8670 , new_n8657 , new_n8669 );
and  g06322 ( new_n8671 , new_n8656_1 , new_n8670 );
or   g06323 ( new_n8672 , new_n8655 , new_n8671 );
and  g06324 ( new_n8673 , new_n8654 , new_n8672 );
or   g06325 ( new_n8674 , new_n8653 , new_n8673 );
and  g06326 ( new_n8675 , new_n8652 , new_n8674 );
or   g06327 ( new_n8676 , new_n8651 , new_n8675 );
and  g06328 ( new_n8677 , new_n8650 , new_n8676 );
or   g06329 ( new_n8678_1 , new_n8649 , new_n8677 );
and  g06330 ( new_n8679 , new_n8648 , new_n8678_1 );
or   g06331 ( new_n8680 , new_n8647 , new_n8679 );
xor  g06332 ( new_n8681 , new_n8645 , new_n8680 );
xnor g06333 ( new_n8682 , n2978 , n20040 );
nor  g06334 ( new_n8683 , n19531 , new_n6744 );
xnor g06335 ( new_n8684 , n19531 , n23697 );
nor  g06336 ( new_n8685 , new_n6748 , n18345 );
xnor g06337 ( new_n8686 , n2289 , n18345 );
nor  g06338 ( new_n8687_1 , new_n6752 , n13190 );
xnor g06339 ( new_n8688 , n1112 , n13190 );
nor  g06340 ( new_n8689 , n3460 , new_n6756 );
xnor g06341 ( new_n8690 , n3460 , n20179 );
nor  g06342 ( new_n8691 , n5226 , new_n7440 );
xnor g06343 ( new_n8692 , n5226 , n19228 );
nor  g06344 ( new_n8693 , new_n6763 , n17664 );
xnor g06345 ( new_n8694_1 , n15539 , n17664 );
nor  g06346 ( new_n8695 , n8052 , new_n2578_1 );
nor  g06347 ( new_n8696 , new_n6767 , n23369 );
not  g06348 ( new_n8697 , n1136 );
nor  g06349 ( new_n8698 , new_n8697 , n10158 );
nor  g06350 ( new_n8699 , n1136 , new_n7448 );
nor  g06351 ( new_n8700 , n18962 , new_n2582_1 );
not  g06352 ( new_n8701 , new_n8700 );
nor  g06353 ( new_n8702 , new_n8699 , new_n8701 );
nor  g06354 ( new_n8703 , new_n8698 , new_n8702 );
nor  g06355 ( new_n8704 , new_n8696 , new_n8703 );
nor  g06356 ( new_n8705 , new_n8695 , new_n8704 );
and  g06357 ( new_n8706 , new_n8694_1 , new_n8705 );
or   g06358 ( new_n8707 , new_n8693 , new_n8706 );
and  g06359 ( new_n8708 , new_n8692 , new_n8707 );
or   g06360 ( new_n8709 , new_n8691 , new_n8708 );
and  g06361 ( new_n8710 , new_n8690 , new_n8709 );
or   g06362 ( new_n8711 , new_n8689 , new_n8710 );
and  g06363 ( new_n8712 , new_n8688 , new_n8711 );
or   g06364 ( new_n8713 , new_n8687_1 , new_n8712 );
and  g06365 ( new_n8714 , new_n8686 , new_n8713 );
or   g06366 ( new_n8715 , new_n8685 , new_n8714 );
and  g06367 ( new_n8716_1 , new_n8684 , new_n8715 );
nor  g06368 ( new_n8717 , new_n8683 , new_n8716_1 );
xnor g06369 ( new_n8718 , new_n8682 , new_n8717 );
not  g06370 ( new_n8719 , n12507 );
nor  g06371 ( new_n8720 , n4588 , n15258 );
not  g06372 ( new_n8721_1 , new_n8720 );
nor  g06373 ( new_n8722 , n16743 , new_n8721_1 );
not  g06374 ( new_n8723 , new_n8722 );
nor  g06375 ( new_n8724 , n22631 , new_n8723 );
not  g06376 ( new_n8725 , new_n8724 );
nor  g06377 ( new_n8726 , n2331 , new_n8725 );
not  g06378 ( new_n8727 , new_n8726 );
nor  g06379 ( new_n8728 , n25068 , new_n8727 );
not  g06380 ( new_n8729 , new_n8728 );
nor  g06381 ( new_n8730 , n16812 , new_n8729 );
not  g06382 ( new_n8731 , new_n8730 );
nor  g06383 ( new_n8732 , n7841 , new_n8731 );
not  g06384 ( new_n8733 , new_n8732 );
nor  g06385 ( new_n8734 , n26264 , new_n8733 );
xnor g06386 ( new_n8735 , n22764 , new_n8734 );
xnor g06387 ( new_n8736 , new_n8719 , new_n8735 );
xnor g06388 ( new_n8737 , n26264 , new_n8732 );
and  g06389 ( new_n8738 , n15077 , new_n8737 );
nor  g06390 ( new_n8739 , n15077 , new_n8737 );
xnor g06391 ( new_n8740 , n7841 , new_n8730 );
and  g06392 ( new_n8741 , n3710 , new_n8740 );
or   g06393 ( new_n8742 , n3710 , new_n8740 );
xnor g06394 ( new_n8743 , n16812 , new_n8728 );
nor  g06395 ( new_n8744_1 , n26318 , new_n8743 );
not  g06396 ( new_n8745_1 , n26318 );
xnor g06397 ( new_n8746 , new_n8745_1 , new_n8743 );
xnor g06398 ( new_n8747 , n25068 , new_n8726 );
nor  g06399 ( new_n8748 , n26054 , new_n8747 );
not  g06400 ( new_n8749 , n26054 );
xnor g06401 ( new_n8750 , new_n8749 , new_n8747 );
xnor g06402 ( new_n8751 , n2331 , new_n8724 );
nor  g06403 ( new_n8752 , n19081 , new_n8751 );
not  g06404 ( new_n8753 , n19081 );
xnor g06405 ( new_n8754 , new_n8753 , new_n8751 );
xnor g06406 ( new_n8755 , n22631 , new_n8722 );
nor  g06407 ( new_n8756 , n8309 , new_n8755 );
xnor g06408 ( new_n8757 , n16743 , new_n8720 );
nor  g06409 ( new_n8758 , n19144 , new_n8757 );
not  g06410 ( new_n8759 , n19144 );
xnor g06411 ( new_n8760 , new_n8759 , new_n8757 );
xnor g06412 ( new_n8761 , new_n2542 , n15258 );
nor  g06413 ( new_n8762 , n12593 , new_n8761 );
not  g06414 ( new_n8763 , n13714 );
or   g06415 ( new_n8764 , new_n2542 , new_n8763 );
not  g06416 ( new_n8765 , new_n8761 );
xnor g06417 ( new_n8766 , n12593 , new_n8765 );
and  g06418 ( new_n8767 , new_n8764 , new_n8766 );
or   g06419 ( new_n8768 , new_n8762 , new_n8767 );
and  g06420 ( new_n8769 , new_n8760 , new_n8768 );
or   g06421 ( new_n8770 , new_n8758 , new_n8769 );
not  g06422 ( new_n8771 , n8309 );
xnor g06423 ( new_n8772 , new_n8771 , new_n8755 );
and  g06424 ( new_n8773 , new_n8770 , new_n8772 );
or   g06425 ( new_n8774 , new_n8756 , new_n8773 );
and  g06426 ( new_n8775 , new_n8754 , new_n8774 );
or   g06427 ( new_n8776 , new_n8752 , new_n8775 );
and  g06428 ( new_n8777 , new_n8750 , new_n8776 );
or   g06429 ( new_n8778 , new_n8748 , new_n8777 );
and  g06430 ( new_n8779 , new_n8746 , new_n8778 );
nor  g06431 ( new_n8780 , new_n8744_1 , new_n8779 );
and  g06432 ( new_n8781 , new_n8742 , new_n8780 );
nor  g06433 ( new_n8782_1 , new_n8741 , new_n8781 );
nor  g06434 ( new_n8783 , new_n8739 , new_n8782_1 );
nor  g06435 ( new_n8784 , new_n8738 , new_n8783 );
xnor g06436 ( new_n8785 , new_n8736 , new_n8784 );
xnor g06437 ( new_n8786 , new_n8718 , new_n8785 );
nor  g06438 ( new_n8787 , new_n8685 , new_n8714 );
xnor g06439 ( new_n8788 , new_n8684 , new_n8787 );
not  g06440 ( new_n8789 , n15077 );
xnor g06441 ( new_n8790 , new_n8789 , new_n8737 );
xnor g06442 ( new_n8791 , new_n8782_1 , new_n8790 );
and  g06443 ( new_n8792 , new_n8788 , new_n8791 );
not  g06444 ( new_n8793 , new_n8788 );
xnor g06445 ( new_n8794 , new_n8793 , new_n8791 );
xor  g06446 ( new_n8795 , new_n8686 , new_n8713 );
xnor g06447 ( new_n8796 , n3710 , new_n8740 );
xnor g06448 ( new_n8797 , new_n8780 , new_n8796 );
nor  g06449 ( new_n8798 , new_n8795 , new_n8797 );
xnor g06450 ( new_n8799 , new_n8795 , new_n8797 );
nor  g06451 ( new_n8800 , new_n8689 , new_n8710 );
xnor g06452 ( new_n8801 , new_n8688 , new_n8800 );
not  g06453 ( new_n8802 , new_n8801 );
xor  g06454 ( new_n8803_1 , new_n8746 , new_n8778 );
and  g06455 ( new_n8804 , new_n8802 , new_n8803_1 );
xnor g06456 ( new_n8805 , new_n8802 , new_n8803_1 );
nor  g06457 ( new_n8806_1 , new_n8691 , new_n8708 );
xnor g06458 ( new_n8807 , new_n8690 , new_n8806_1 );
not  g06459 ( new_n8808 , new_n8807 );
xor  g06460 ( new_n8809_1 , new_n8750 , new_n8776 );
and  g06461 ( new_n8810 , new_n8808 , new_n8809_1 );
xnor g06462 ( new_n8811 , new_n8808 , new_n8809_1 );
nor  g06463 ( new_n8812 , new_n8693 , new_n8706 );
xnor g06464 ( new_n8813 , new_n8692 , new_n8812 );
not  g06465 ( new_n8814 , new_n8813 );
xor  g06466 ( new_n8815 , new_n8754 , new_n8774 );
and  g06467 ( new_n8816 , new_n8814 , new_n8815 );
xnor g06468 ( new_n8817 , new_n8814 , new_n8815 );
xnor g06469 ( new_n8818 , new_n8694_1 , new_n8705 );
xor  g06470 ( new_n8819 , new_n8770 , new_n8772 );
and  g06471 ( new_n8820 , new_n8818 , new_n8819 );
not  g06472 ( new_n8821_1 , new_n8818 );
xnor g06473 ( new_n8822 , new_n8821_1 , new_n8819 );
xor  g06474 ( new_n8823 , new_n8760 , new_n8768 );
xnor g06475 ( new_n8824_1 , n8052 , n23369 );
xnor g06476 ( new_n8825 , new_n8703 , new_n8824_1 );
nor  g06477 ( new_n8826 , new_n8823 , new_n8825 );
xnor g06478 ( new_n8827_1 , new_n8823 , new_n8825 );
xor  g06479 ( new_n8828 , new_n8764 , new_n8766 );
xnor g06480 ( new_n8829 , n1136 , n10158 );
xnor g06481 ( new_n8830 , new_n8701 , new_n8829 );
nor  g06482 ( new_n8831 , new_n8828 , new_n8830 );
xnor g06483 ( new_n8832 , n18962 , n19234 );
xnor g06484 ( new_n8833 , n4588 , n13714 );
nor  g06485 ( new_n8834 , new_n8832 , new_n8833 );
not  g06486 ( new_n8835 , new_n8830 );
xnor g06487 ( new_n8836 , new_n8828 , new_n8835 );
and  g06488 ( new_n8837 , new_n8834 , new_n8836 );
nor  g06489 ( new_n8838 , new_n8831 , new_n8837 );
nor  g06490 ( new_n8839 , new_n8827_1 , new_n8838 );
nor  g06491 ( new_n8840 , new_n8826 , new_n8839 );
and  g06492 ( new_n8841 , new_n8822 , new_n8840 );
nor  g06493 ( new_n8842 , new_n8820 , new_n8841 );
nor  g06494 ( new_n8843 , new_n8817 , new_n8842 );
nor  g06495 ( new_n8844 , new_n8816 , new_n8843 );
nor  g06496 ( new_n8845 , new_n8811 , new_n8844 );
nor  g06497 ( new_n8846 , new_n8810 , new_n8845 );
nor  g06498 ( new_n8847 , new_n8805 , new_n8846 );
nor  g06499 ( new_n8848 , new_n8804 , new_n8847 );
nor  g06500 ( new_n8849_1 , new_n8799 , new_n8848 );
nor  g06501 ( new_n8850 , new_n8798 , new_n8849_1 );
and  g06502 ( new_n8851 , new_n8794 , new_n8850 );
nor  g06503 ( new_n8852 , new_n8792 , new_n8851 );
xnor g06504 ( new_n8853 , new_n8786 , new_n8852 );
xnor g06505 ( new_n8854 , new_n8681 , new_n8853 );
xor  g06506 ( new_n8855 , new_n8648 , new_n8678_1 );
xor  g06507 ( new_n8856_1 , new_n8794 , new_n8850 );
nor  g06508 ( new_n8857 , new_n8855 , new_n8856_1 );
xnor g06509 ( new_n8858 , new_n8855 , new_n8856_1 );
xor  g06510 ( new_n8859 , new_n8650 , new_n8676 );
xnor g06511 ( new_n8860 , new_n8799 , new_n8848 );
nor  g06512 ( new_n8861_1 , new_n8859 , new_n8860 );
xnor g06513 ( new_n8862_1 , new_n8859 , new_n8860 );
xor  g06514 ( new_n8863 , new_n8652 , new_n8674 );
xnor g06515 ( new_n8864 , new_n8805 , new_n8846 );
nor  g06516 ( new_n8865 , new_n8863 , new_n8864 );
xnor g06517 ( new_n8866 , new_n8863 , new_n8864 );
xor  g06518 ( new_n8867 , new_n8654 , new_n8672 );
xnor g06519 ( new_n8868 , new_n8811 , new_n8844 );
nor  g06520 ( new_n8869_1 , new_n8867 , new_n8868 );
xnor g06521 ( new_n8870 , new_n8867 , new_n8868 );
xor  g06522 ( new_n8871 , new_n8656_1 , new_n8670 );
xnor g06523 ( new_n8872 , new_n8817 , new_n8842 );
nor  g06524 ( new_n8873 , new_n8871 , new_n8872 );
xnor g06525 ( new_n8874 , new_n8871 , new_n8872 );
xnor g06526 ( new_n8875 , new_n8822 , new_n8840 );
not  g06527 ( new_n8876 , new_n8875 );
xnor g06528 ( new_n8877 , new_n8658 , new_n8668 );
and  g06529 ( new_n8878 , new_n8876 , new_n8877 );
xnor g06530 ( new_n8879 , new_n8876 , new_n8877 );
xnor g06531 ( new_n8880 , new_n8827_1 , new_n8838 );
xnor g06532 ( new_n8881 , n20036 , n24786 );
xnor g06533 ( new_n8882 , new_n8666 , new_n8881 );
and  g06534 ( new_n8883 , new_n8880 , new_n8882 );
xnor g06535 ( new_n8884_1 , new_n8880 , new_n8882 );
xnor g06536 ( new_n8885 , n9380 , n23065 );
xnor g06537 ( new_n8886 , new_n8832 , new_n8833 );
nor  g06538 ( new_n8887 , new_n8885 , new_n8886 );
xnor g06539 ( new_n8888 , n11192 , n27120 );
xnor g06540 ( new_n8889 , new_n8664 , new_n8888 );
nor  g06541 ( new_n8890 , new_n8887 , new_n8889 );
xnor g06542 ( new_n8891 , new_n8834 , new_n8836 );
not  g06543 ( new_n8892 , new_n8891 );
xnor g06544 ( new_n8893 , new_n8887 , new_n8889 );
nor  g06545 ( new_n8894 , new_n8892 , new_n8893 );
nor  g06546 ( new_n8895 , new_n8890 , new_n8894 );
nor  g06547 ( new_n8896 , new_n8884_1 , new_n8895 );
nor  g06548 ( new_n8897 , new_n8883 , new_n8896 );
nor  g06549 ( new_n8898 , new_n8879 , new_n8897 );
nor  g06550 ( new_n8899 , new_n8878 , new_n8898 );
nor  g06551 ( new_n8900 , new_n8874 , new_n8899 );
nor  g06552 ( new_n8901 , new_n8873 , new_n8900 );
nor  g06553 ( new_n8902 , new_n8870 , new_n8901 );
nor  g06554 ( new_n8903 , new_n8869_1 , new_n8902 );
nor  g06555 ( new_n8904 , new_n8866 , new_n8903 );
nor  g06556 ( new_n8905 , new_n8865 , new_n8904 );
nor  g06557 ( new_n8906 , new_n8862_1 , new_n8905 );
nor  g06558 ( new_n8907 , new_n8861_1 , new_n8906 );
nor  g06559 ( new_n8908 , new_n8858 , new_n8907 );
nor  g06560 ( new_n8909_1 , new_n8857 , new_n8908 );
xor  g06561 ( n957 , new_n8854 , new_n8909_1 );
xnor g06562 ( new_n8911_1 , n20385 , new_n8832 );
xnor g06563 ( new_n8912 , new_n4122 , n26167 );
xnor g06564 ( new_n8913 , n21138 , new_n8912 );
xnor g06565 ( n980 , new_n8911_1 , new_n8913 );
nor  g06566 ( new_n8915 , new_n4357 , new_n7702 );
xnor g06567 ( new_n8916 , new_n4357 , new_n7698_1 );
nor  g06568 ( new_n8917 , new_n4359 , new_n7705 );
xnor g06569 ( new_n8918 , new_n4359 , new_n7705 );
nor  g06570 ( new_n8919 , new_n4363 , new_n7710 );
xnor g06571 ( new_n8920_1 , new_n4363 , new_n7710 );
nor  g06572 ( new_n8921 , new_n4367 , new_n7717 );
xnor g06573 ( new_n8922 , new_n4367 , new_n7717 );
nor  g06574 ( new_n8923 , new_n4371 , new_n7721_1 );
xnor g06575 ( new_n8924 , new_n4371 , new_n7721_1 );
nor  g06576 ( new_n8925 , new_n4375 , new_n7725 );
xnor g06577 ( new_n8926 , new_n4375 , new_n7725 );
nor  g06578 ( new_n8927 , new_n4380 , new_n7730 );
xnor g06579 ( new_n8928 , new_n4380 , new_n7730 );
nor  g06580 ( new_n8929 , new_n4388 , new_n7739 );
xnor g06581 ( new_n8930 , new_n4388 , new_n7735 );
nor  g06582 ( new_n8931 , new_n4391 , new_n7742 );
nor  g06583 ( new_n8932 , new_n4395 , new_n7748 );
xnor g06584 ( new_n8933 , new_n4392 , new_n7742 );
and  g06585 ( new_n8934 , new_n8932 , new_n8933 );
nor  g06586 ( new_n8935 , new_n8931 , new_n8934 );
and  g06587 ( new_n8936 , new_n8930 , new_n8935 );
nor  g06588 ( new_n8937 , new_n8929 , new_n8936 );
nor  g06589 ( new_n8938 , new_n8928 , new_n8937 );
nor  g06590 ( new_n8939 , new_n8927 , new_n8938 );
nor  g06591 ( new_n8940 , new_n8926 , new_n8939 );
nor  g06592 ( new_n8941 , new_n8925 , new_n8940 );
nor  g06593 ( new_n8942 , new_n8924 , new_n8941 );
nor  g06594 ( new_n8943_1 , new_n8923 , new_n8942 );
nor  g06595 ( new_n8944 , new_n8922 , new_n8943_1 );
nor  g06596 ( new_n8945 , new_n8921 , new_n8944 );
nor  g06597 ( new_n8946 , new_n8920_1 , new_n8945 );
nor  g06598 ( new_n8947 , new_n8919 , new_n8946 );
nor  g06599 ( new_n8948 , new_n8918 , new_n8947 );
nor  g06600 ( new_n8949 , new_n8917 , new_n8948 );
and  g06601 ( new_n8950 , new_n8916 , new_n8949 );
or   g06602 ( new_n8951 , new_n8915 , new_n8950 );
xnor g06603 ( new_n8952 , new_n4353 , new_n7695 );
xor  g06604 ( new_n8953 , new_n8951 , new_n8952 );
not  g06605 ( new_n8954 , n16544 );
nor  g06606 ( new_n8955 , n12650 , new_n8954 );
xnor g06607 ( new_n8956 , n12650 , n16544 );
nor  g06608 ( new_n8957 , new_n2887_1 , n10201 );
xnor g06609 ( new_n8958 , n6814 , n10201 );
not  g06610 ( new_n8959 , n19701 );
nor  g06611 ( new_n8960 , n10593 , new_n8959 );
xnor g06612 ( new_n8961 , n10593 , n19701 );
not  g06613 ( new_n8962 , n23529 );
nor  g06614 ( new_n8963 , n18290 , new_n8962 );
xnor g06615 ( new_n8964_1 , n18290 , n23529 );
not  g06616 ( new_n8965 , n24620 );
nor  g06617 ( new_n8966 , n11580 , new_n8965 );
xnor g06618 ( new_n8967 , n11580 , n24620 );
not  g06619 ( new_n8968 , n5211 );
nor  g06620 ( new_n8969 , new_n8968 , n15884 );
xnor g06621 ( new_n8970 , n5211 , n15884 );
not  g06622 ( new_n8971_1 , n12956 );
nor  g06623 ( new_n8972 , n6356 , new_n8971_1 );
xnor g06624 ( new_n8973 , n6356 , n12956 );
nor  g06625 ( new_n8974 , n18295 , new_n5582 );
nor  g06626 ( new_n8975 , new_n2903 , n27104 );
nor  g06627 ( new_n8976 , n6502 , new_n5584 );
or   g06628 ( new_n8977 , new_n5033 , n27188 );
nor  g06629 ( new_n8978 , new_n5588 , n15780 );
and  g06630 ( new_n8979 , new_n8977 , new_n8978 );
nor  g06631 ( new_n8980 , new_n8976 , new_n8979 );
nor  g06632 ( new_n8981 , new_n8975 , new_n8980 );
nor  g06633 ( new_n8982_1 , new_n8974 , new_n8981 );
and  g06634 ( new_n8983 , new_n8973 , new_n8982_1 );
or   g06635 ( new_n8984 , new_n8972 , new_n8983 );
and  g06636 ( new_n8985 , new_n8970 , new_n8984 );
or   g06637 ( new_n8986 , new_n8969 , new_n8985 );
and  g06638 ( new_n8987 , new_n8967 , new_n8986 );
or   g06639 ( new_n8988 , new_n8966 , new_n8987 );
and  g06640 ( new_n8989 , new_n8964_1 , new_n8988 );
or   g06641 ( new_n8990 , new_n8963 , new_n8989 );
and  g06642 ( new_n8991 , new_n8961 , new_n8990 );
or   g06643 ( new_n8992 , new_n8960 , new_n8991 );
and  g06644 ( new_n8993_1 , new_n8958 , new_n8992 );
or   g06645 ( new_n8994 , new_n8957 , new_n8993_1 );
and  g06646 ( new_n8995 , new_n8956 , new_n8994 );
nor  g06647 ( new_n8996 , new_n8955 , new_n8995 );
xnor g06648 ( new_n8997 , new_n8953 , new_n8996 );
xor  g06649 ( new_n8998 , new_n8956 , new_n8994 );
xor  g06650 ( new_n8999 , new_n8916 , new_n8949 );
nor  g06651 ( new_n9000 , new_n8998 , new_n8999 );
xnor g06652 ( new_n9001 , new_n8998 , new_n8999 );
xor  g06653 ( new_n9002 , new_n8958 , new_n8992 );
xnor g06654 ( new_n9003_1 , new_n8918 , new_n8947 );
nor  g06655 ( new_n9004 , new_n9002 , new_n9003_1 );
xnor g06656 ( new_n9005 , new_n9002 , new_n9003_1 );
xor  g06657 ( new_n9006 , new_n8961 , new_n8990 );
xnor g06658 ( new_n9007 , new_n8920_1 , new_n8945 );
nor  g06659 ( new_n9008 , new_n9006 , new_n9007 );
xnor g06660 ( new_n9009 , new_n9006 , new_n9007 );
xor  g06661 ( new_n9010 , new_n8964_1 , new_n8988 );
xnor g06662 ( new_n9011 , new_n8922 , new_n8943_1 );
nor  g06663 ( new_n9012_1 , new_n9010 , new_n9011 );
xnor g06664 ( new_n9013 , new_n9010 , new_n9011 );
xor  g06665 ( new_n9014 , new_n8967 , new_n8986 );
xnor g06666 ( new_n9015 , new_n8924 , new_n8941 );
nor  g06667 ( new_n9016 , new_n9014 , new_n9015 );
xnor g06668 ( new_n9017 , new_n9014 , new_n9015 );
xor  g06669 ( new_n9018 , new_n8970 , new_n8984 );
xnor g06670 ( new_n9019 , new_n8926 , new_n8939 );
nor  g06671 ( new_n9020 , new_n9018 , new_n9019 );
xnor g06672 ( new_n9021 , new_n9018 , new_n9019 );
xnor g06673 ( new_n9022 , new_n8928 , new_n8937 );
not  g06674 ( new_n9023 , new_n9022 );
xnor g06675 ( new_n9024 , new_n8973 , new_n8982_1 );
and  g06676 ( new_n9025 , new_n9023 , new_n9024 );
xnor g06677 ( new_n9026 , new_n8930 , new_n8935 );
not  g06678 ( new_n9027 , new_n9026 );
xnor g06679 ( new_n9028 , n18295 , n27104 );
xnor g06680 ( new_n9029 , new_n8980 , new_n9028 );
and  g06681 ( new_n9030 , new_n9027 , new_n9029 );
xnor g06682 ( new_n9031 , new_n9027 , new_n9029 );
xnor g06683 ( new_n9032_1 , n6611 , n15780 );
xnor g06684 ( new_n9033 , new_n4395 , new_n7888 );
not  g06685 ( new_n9034 , new_n9033 );
nor  g06686 ( new_n9035 , new_n9032_1 , new_n9034 );
xnor g06687 ( new_n9036 , n6502 , n27188 );
xnor g06688 ( new_n9037 , new_n8978 , new_n9036 );
nor  g06689 ( new_n9038 , new_n9035 , new_n9037 );
xor  g06690 ( new_n9039 , new_n8932 , new_n8933 );
xnor g06691 ( new_n9040 , new_n9035 , new_n9037 );
nor  g06692 ( new_n9041 , new_n9039 , new_n9040 );
nor  g06693 ( new_n9042_1 , new_n9038 , new_n9041 );
nor  g06694 ( new_n9043 , new_n9031 , new_n9042_1 );
nor  g06695 ( new_n9044 , new_n9030 , new_n9043 );
xnor g06696 ( new_n9045 , new_n9023 , new_n9024 );
nor  g06697 ( new_n9046_1 , new_n9044 , new_n9045 );
nor  g06698 ( new_n9047_1 , new_n9025 , new_n9046_1 );
nor  g06699 ( new_n9048 , new_n9021 , new_n9047_1 );
nor  g06700 ( new_n9049 , new_n9020 , new_n9048 );
nor  g06701 ( new_n9050 , new_n9017 , new_n9049 );
nor  g06702 ( new_n9051 , new_n9016 , new_n9050 );
nor  g06703 ( new_n9052 , new_n9013 , new_n9051 );
nor  g06704 ( new_n9053 , new_n9012_1 , new_n9052 );
nor  g06705 ( new_n9054 , new_n9009 , new_n9053 );
nor  g06706 ( new_n9055 , new_n9008 , new_n9054 );
nor  g06707 ( new_n9056 , new_n9005 , new_n9055 );
nor  g06708 ( new_n9057 , new_n9004 , new_n9056 );
nor  g06709 ( new_n9058 , new_n9001 , new_n9057 );
nor  g06710 ( new_n9059 , new_n9000 , new_n9058 );
xnor g06711 ( n982 , new_n8997 , new_n9059 );
not  g06712 ( new_n9061 , new_n4544 );
not  g06713 ( new_n9062 , n3279 );
nor  g06714 ( new_n9063 , n7339 , n26808 );
not  g06715 ( new_n9064 , new_n9063 );
nor  g06716 ( new_n9065 , n1667 , new_n9064 );
not  g06717 ( new_n9066 , new_n9065 );
nor  g06718 ( new_n9067 , n2680 , new_n9066 );
not  g06719 ( new_n9068 , new_n9067 );
nor  g06720 ( new_n9069 , n2547 , new_n9068 );
not  g06721 ( new_n9070 , new_n9069 );
nor  g06722 ( new_n9071 , n2999 , new_n9070 );
not  g06723 ( new_n9072 , new_n9071 );
nor  g06724 ( new_n9073 , n14702 , new_n9072 );
not  g06725 ( new_n9074 , new_n9073 );
nor  g06726 ( new_n9075 , n13914 , new_n9074 );
and  g06727 ( new_n9076 , new_n9062 , new_n9075 );
xnor g06728 ( new_n9077 , n4306 , new_n9076 );
xnor g06729 ( new_n9078 , n18105 , n23166 );
not  g06730 ( new_n9079 , n10577 );
nor  g06731 ( new_n9080 , new_n9079 , n24196 );
xnor g06732 ( new_n9081 , n10577 , n24196 );
not  g06733 ( new_n9082 , n6381 );
nor  g06734 ( new_n9083 , new_n9082 , n16376 );
xnor g06735 ( new_n9084 , n6381 , n16376 );
not  g06736 ( new_n9085 , n14345 );
nor  g06737 ( new_n9086 , new_n9085 , n25381 );
xnor g06738 ( new_n9087 , n14345 , n25381 );
not  g06739 ( new_n9088 , n11356 );
nor  g06740 ( new_n9089 , new_n9088 , n12587 );
xnor g06741 ( new_n9090_1 , n11356 , n12587 );
not  g06742 ( new_n9091 , n3164 );
nor  g06743 ( new_n9092 , n268 , new_n9091 );
xnor g06744 ( new_n9093 , n268 , n3164 );
nor  g06745 ( new_n9094 , new_n6590_1 , n24879 );
xnor g06746 ( new_n9095 , n10611 , n24879 );
nor  g06747 ( new_n9096 , n2783 , new_n8048 );
nor  g06748 ( new_n9097 , new_n6593 , n6785 );
nor  g06749 ( new_n9098 , n15490 , new_n8052_1 );
not  g06750 ( new_n9099 , n15490 );
nor  g06751 ( new_n9100 , new_n9099 , n24032 );
nor  g06752 ( new_n9101 , n18 , new_n4507 );
not  g06753 ( new_n9102 , new_n9101 );
nor  g06754 ( new_n9103 , new_n9100 , new_n9102 );
nor  g06755 ( new_n9104_1 , new_n9098 , new_n9103 );
nor  g06756 ( new_n9105 , new_n9097 , new_n9104_1 );
nor  g06757 ( new_n9106 , new_n9096 , new_n9105 );
and  g06758 ( new_n9107 , new_n9095 , new_n9106 );
or   g06759 ( new_n9108 , new_n9094 , new_n9107 );
and  g06760 ( new_n9109 , new_n9093 , new_n9108 );
or   g06761 ( new_n9110 , new_n9092 , new_n9109 );
and  g06762 ( new_n9111 , new_n9090_1 , new_n9110 );
or   g06763 ( new_n9112 , new_n9089 , new_n9111 );
and  g06764 ( new_n9113 , new_n9087 , new_n9112 );
or   g06765 ( new_n9114 , new_n9086 , new_n9113 );
and  g06766 ( new_n9115 , new_n9084 , new_n9114 );
or   g06767 ( new_n9116 , new_n9083 , new_n9115 );
and  g06768 ( new_n9117 , new_n9081 , new_n9116 );
nor  g06769 ( new_n9118 , new_n9080 , new_n9117 );
xnor g06770 ( new_n9119 , new_n9078 , new_n9118 );
xor  g06771 ( new_n9120 , new_n9077 , new_n9119 );
xnor g06772 ( new_n9121 , n3279 , new_n9075 );
nor  g06773 ( new_n9122 , new_n9083 , new_n9115 );
xnor g06774 ( new_n9123 , new_n9081 , new_n9122 );
and  g06775 ( new_n9124 , new_n9121 , new_n9123 );
xor  g06776 ( new_n9125 , new_n9121 , new_n9123 );
xnor g06777 ( new_n9126 , n13914 , new_n9073 );
xor  g06778 ( new_n9127 , new_n9084 , new_n9114 );
nor  g06779 ( new_n9128 , new_n9126 , new_n9127 );
xnor g06780 ( new_n9129_1 , new_n9126 , new_n9127 );
xnor g06781 ( new_n9130 , n14702 , new_n9071 );
xor  g06782 ( new_n9131 , new_n9087 , new_n9112 );
nor  g06783 ( new_n9132 , new_n9130 , new_n9131 );
xnor g06784 ( new_n9133 , new_n9130 , new_n9131 );
xnor g06785 ( new_n9134 , n2999 , new_n9069 );
xor  g06786 ( new_n9135 , new_n9090_1 , new_n9110 );
nor  g06787 ( new_n9136 , new_n9134 , new_n9135 );
xnor g06788 ( new_n9137 , n2547 , new_n9067 );
xor  g06789 ( new_n9138 , new_n9093 , new_n9108 );
nor  g06790 ( new_n9139 , new_n9137 , new_n9138 );
xnor g06791 ( new_n9140 , new_n9137 , new_n9138 );
xnor g06792 ( new_n9141 , n2680 , new_n9065 );
xnor g06793 ( new_n9142 , new_n9095 , new_n9106 );
not  g06794 ( new_n9143 , new_n9142 );
nor  g06795 ( new_n9144 , new_n9141 , new_n9143 );
xnor g06796 ( new_n9145 , n1667 , new_n9063 );
xnor g06797 ( new_n9146_1 , n2783 , n6785 );
xnor g06798 ( new_n9147 , new_n9104_1 , new_n9146_1 );
not  g06799 ( new_n9148 , new_n9147 );
nor  g06800 ( new_n9149 , new_n9145 , new_n9148 );
xnor g06801 ( new_n9150 , new_n9145 , new_n9147 );
xnor g06802 ( new_n9151 , n7339 , n26808 );
xnor g06803 ( new_n9152 , n15490 , n24032 );
xnor g06804 ( new_n9153 , new_n9102 , new_n9152 );
nor  g06805 ( new_n9154 , new_n9151 , new_n9153 );
not  g06806 ( new_n9155 , n26808 );
xnor g06807 ( new_n9156 , n18 , n22843 );
nor  g06808 ( new_n9157 , new_n9155 , new_n9156 );
not  g06809 ( new_n9158 , new_n9153 );
xnor g06810 ( new_n9159 , new_n9151 , new_n9158 );
and  g06811 ( new_n9160 , new_n9157 , new_n9159 );
nor  g06812 ( new_n9161 , new_n9154 , new_n9160 );
and  g06813 ( new_n9162 , new_n9150 , new_n9161 );
or   g06814 ( new_n9163 , new_n9149 , new_n9162 );
xnor g06815 ( new_n9164_1 , new_n9141 , new_n9142 );
and  g06816 ( new_n9165 , new_n9163 , new_n9164_1 );
nor  g06817 ( new_n9166_1 , new_n9144 , new_n9165 );
nor  g06818 ( new_n9167 , new_n9140 , new_n9166_1 );
nor  g06819 ( new_n9168 , new_n9139 , new_n9167 );
xnor g06820 ( new_n9169 , new_n9134 , new_n9135 );
nor  g06821 ( new_n9170 , new_n9168 , new_n9169 );
nor  g06822 ( new_n9171 , new_n9136 , new_n9170 );
nor  g06823 ( new_n9172_1 , new_n9133 , new_n9171 );
nor  g06824 ( new_n9173 , new_n9132 , new_n9172_1 );
nor  g06825 ( new_n9174 , new_n9129_1 , new_n9173 );
nor  g06826 ( new_n9175 , new_n9128 , new_n9174 );
and  g06827 ( new_n9176 , new_n9125 , new_n9175 );
or   g06828 ( new_n9177 , new_n9124 , new_n9176 );
xor  g06829 ( new_n9178 , new_n9120 , new_n9177 );
xnor g06830 ( new_n9179 , new_n9061 , new_n9178 );
xor  g06831 ( new_n9180 , new_n9125 , new_n9175 );
nor  g06832 ( new_n9181 , new_n4549 , new_n9180 );
xnor g06833 ( new_n9182_1 , new_n4549 , new_n9180 );
xnor g06834 ( new_n9183 , new_n9129_1 , new_n9173 );
nor  g06835 ( new_n9184 , new_n4554 , new_n9183 );
xnor g06836 ( new_n9185 , new_n4554 , new_n9183 );
xnor g06837 ( new_n9186 , new_n9133 , new_n9171 );
nor  g06838 ( new_n9187 , new_n4559 , new_n9186 );
xnor g06839 ( new_n9188 , new_n4559 , new_n9186 );
xnor g06840 ( new_n9189 , new_n9168 , new_n9169 );
nor  g06841 ( new_n9190 , new_n4564 , new_n9189 );
xnor g06842 ( new_n9191_1 , new_n4564 , new_n9189 );
xnor g06843 ( new_n9192 , new_n9140 , new_n9166_1 );
nor  g06844 ( new_n9193 , new_n4568 , new_n9192 );
xnor g06845 ( new_n9194 , new_n4568 , new_n9192 );
xor  g06846 ( new_n9195 , new_n9163 , new_n9164_1 );
and  g06847 ( new_n9196 , new_n4575 , new_n9195 );
xnor g06848 ( new_n9197 , new_n4573 , new_n9195 );
xor  g06849 ( new_n9198 , new_n9150 , new_n9161 );
nor  g06850 ( new_n9199 , new_n4579 , new_n9198 );
xnor g06851 ( new_n9200 , new_n4591 , new_n9198 );
xnor g06852 ( new_n9201 , new_n9157 , new_n9159 );
nor  g06853 ( new_n9202 , new_n4581 , new_n9201 );
xnor g06854 ( new_n9203 , n26808 , new_n9156 );
and  g06855 ( new_n9204 , new_n4585 , new_n9203 );
xor  g06856 ( new_n9205 , new_n4581 , new_n9201 );
and  g06857 ( new_n9206 , new_n9204 , new_n9205 );
or   g06858 ( new_n9207 , new_n9202 , new_n9206 );
and  g06859 ( new_n9208 , new_n9200 , new_n9207 );
nor  g06860 ( new_n9209 , new_n9199 , new_n9208 );
and  g06861 ( new_n9210 , new_n9197 , new_n9209 );
nor  g06862 ( new_n9211 , new_n9196 , new_n9210 );
nor  g06863 ( new_n9212 , new_n9194 , new_n9211 );
nor  g06864 ( new_n9213 , new_n9193 , new_n9212 );
nor  g06865 ( new_n9214 , new_n9191_1 , new_n9213 );
nor  g06866 ( new_n9215 , new_n9190 , new_n9214 );
nor  g06867 ( new_n9216 , new_n9188 , new_n9215 );
nor  g06868 ( new_n9217_1 , new_n9187 , new_n9216 );
nor  g06869 ( new_n9218 , new_n9185 , new_n9217_1 );
nor  g06870 ( new_n9219 , new_n9184 , new_n9218 );
nor  g06871 ( new_n9220_1 , new_n9182_1 , new_n9219 );
nor  g06872 ( new_n9221 , new_n9181 , new_n9220_1 );
xnor g06873 ( n984 , new_n9179 , new_n9221 );
xnor g06874 ( n1005 , new_n9188 , new_n9215 );
xnor g06875 ( n1016 , new_n3344 , new_n3387 );
xnor g06876 ( n1020 , new_n4086 , new_n4100_1 );
xnor g06877 ( new_n9226 , new_n2853_1 , n18290 );
nor  g06878 ( new_n9227 , n2035 , n11580 );
xnor g06879 ( new_n9228 , n2035 , n11580 );
nor  g06880 ( new_n9229 , n5213 , n15884 );
xnor g06881 ( new_n9230 , new_n2859 , n15884 );
nor  g06882 ( new_n9231 , n4665 , n6356 );
xnor g06883 ( new_n9232 , new_n2862 , n6356 );
nor  g06884 ( new_n9233 , n19005 , n27104 );
xnor g06885 ( new_n9234 , new_n2866 , n27104 );
nor  g06886 ( new_n9235 , n4326 , n27188 );
or   g06887 ( new_n9236 , new_n5287 , new_n5588 );
xnor g06888 ( new_n9237 , new_n2869 , n27188 );
and  g06889 ( new_n9238 , new_n9236 , new_n9237 );
or   g06890 ( new_n9239 , new_n9235 , new_n9238 );
and  g06891 ( new_n9240 , new_n9234 , new_n9239 );
or   g06892 ( new_n9241 , new_n9233 , new_n9240 );
and  g06893 ( new_n9242 , new_n9232 , new_n9241 );
or   g06894 ( new_n9243 , new_n9231 , new_n9242 );
and  g06895 ( new_n9244 , new_n9230 , new_n9243 );
nor  g06896 ( new_n9245 , new_n9229 , new_n9244 );
nor  g06897 ( new_n9246_1 , new_n9228 , new_n9245 );
or   g06898 ( new_n9247 , new_n9227 , new_n9246_1 );
xor  g06899 ( new_n9248 , new_n9226 , new_n9247 );
not  g06900 ( new_n9249 , new_n9248 );
xnor g06901 ( new_n9250 , new_n8962 , new_n9249 );
xnor g06902 ( new_n9251_1 , new_n9228 , new_n9245 );
nor  g06903 ( new_n9252 , n24620 , new_n9251_1 );
xnor g06904 ( new_n9253 , new_n8965 , new_n9251_1 );
nor  g06905 ( new_n9254 , new_n9231 , new_n9242 );
xnor g06906 ( new_n9255 , new_n9230 , new_n9254 );
not  g06907 ( new_n9256 , new_n9255 );
nor  g06908 ( new_n9257 , n5211 , new_n9256 );
xnor g06909 ( new_n9258 , new_n8968 , new_n9256 );
nor  g06910 ( new_n9259_1 , new_n9233 , new_n9240 );
xnor g06911 ( new_n9260 , new_n9232 , new_n9259_1 );
not  g06912 ( new_n9261_1 , new_n9260 );
nor  g06913 ( new_n9262 , n12956 , new_n9261_1 );
xnor g06914 ( new_n9263 , new_n8971_1 , new_n9261_1 );
nor  g06915 ( new_n9264 , new_n9235 , new_n9238 );
xnor g06916 ( new_n9265 , new_n9234 , new_n9264 );
not  g06917 ( new_n9266 , new_n9265 );
nor  g06918 ( new_n9267 , n18295 , new_n9266 );
nor  g06919 ( new_n9268 , new_n5287 , new_n5588 );
xnor g06920 ( new_n9269 , new_n9268 , new_n9237 );
nor  g06921 ( new_n9270 , new_n5033 , new_n9269 );
xnor g06922 ( new_n9271 , new_n5287 , n6611 );
not  g06923 ( new_n9272 , new_n9271 );
nor  g06924 ( new_n9273 , new_n2907 , new_n9272 );
not  g06925 ( new_n9274 , new_n9269 );
xnor g06926 ( new_n9275 , new_n5033 , new_n9274 );
and  g06927 ( new_n9276 , new_n9273 , new_n9275 );
nor  g06928 ( new_n9277 , new_n9270 , new_n9276 );
xnor g06929 ( new_n9278 , new_n2903 , new_n9266 );
and  g06930 ( new_n9279 , new_n9277 , new_n9278 );
or   g06931 ( new_n9280 , new_n9267 , new_n9279 );
and  g06932 ( new_n9281 , new_n9263 , new_n9280 );
or   g06933 ( new_n9282 , new_n9262 , new_n9281 );
and  g06934 ( new_n9283 , new_n9258 , new_n9282 );
or   g06935 ( new_n9284 , new_n9257 , new_n9283 );
and  g06936 ( new_n9285 , new_n9253 , new_n9284 );
or   g06937 ( new_n9286 , new_n9252 , new_n9285 );
xor  g06938 ( new_n9287_1 , new_n9250 , new_n9286 );
xnor g06939 ( new_n9288 , new_n6037 , n17250 );
nor  g06940 ( new_n9289 , n3570 , n23160 );
xnor g06941 ( new_n9290 , new_n6043 , n23160 );
nor  g06942 ( new_n9291 , n13668 , n16524 );
xnor g06943 ( new_n9292 , new_n6049 , n16524 );
nor  g06944 ( new_n9293 , n11056 , n21276 );
not  g06945 ( new_n9294 , n11056 );
xnor g06946 ( new_n9295 , new_n9294 , n21276 );
nor  g06947 ( new_n9296 , n15271 , n26748 );
xnor g06948 ( new_n9297 , new_n7668 , n26748 );
nor  g06949 ( new_n9298 , n10057 , n25877 );
nor  g06950 ( new_n9299 , new_n4242 , new_n6629 );
xnor g06951 ( new_n9300 , n10057 , n25877 );
nor  g06952 ( new_n9301 , new_n9299 , new_n9300 );
or   g06953 ( new_n9302 , new_n9298 , new_n9301 );
and  g06954 ( new_n9303 , new_n9297 , new_n9302 );
or   g06955 ( new_n9304 , new_n9296 , new_n9303 );
and  g06956 ( new_n9305 , new_n9295 , new_n9304 );
or   g06957 ( new_n9306 , new_n9293 , new_n9305 );
and  g06958 ( new_n9307 , new_n9292 , new_n9306 );
or   g06959 ( new_n9308_1 , new_n9291 , new_n9307 );
and  g06960 ( new_n9309 , new_n9290 , new_n9308_1 );
nor  g06961 ( new_n9310 , new_n9289 , new_n9309 );
xnor g06962 ( new_n9311 , new_n9288 , new_n9310 );
not  g06963 ( new_n9312 , new_n9311 );
xnor g06964 ( new_n9313 , n11044 , new_n9312 );
nor  g06965 ( new_n9314 , new_n9291 , new_n9307 );
xnor g06966 ( new_n9315 , new_n9290 , new_n9314 );
nor  g06967 ( new_n9316 , new_n5994 , new_n9315 );
not  g06968 ( new_n9317 , new_n9315 );
xnor g06969 ( new_n9318_1 , n2421 , new_n9317 );
nor  g06970 ( new_n9319 , new_n9293 , new_n9305 );
xnor g06971 ( new_n9320 , new_n9292 , new_n9319 );
nor  g06972 ( new_n9321 , new_n7662 , new_n9320 );
not  g06973 ( new_n9322 , new_n9320 );
xnor g06974 ( new_n9323_1 , n987 , new_n9322 );
nor  g06975 ( new_n9324 , new_n9296 , new_n9303 );
xnor g06976 ( new_n9325 , new_n9295 , new_n9324 );
nor  g06977 ( new_n9326 , new_n7665 , new_n9325 );
not  g06978 ( new_n9327 , new_n9325 );
xnor g06979 ( new_n9328 , n20478 , new_n9327 );
nor  g06980 ( new_n9329 , new_n9298 , new_n9301 );
xnor g06981 ( new_n9330 , new_n9297 , new_n9329 );
nor  g06982 ( new_n9331 , new_n7670_1 , new_n9330 );
xnor g06983 ( new_n9332 , new_n9299 , new_n9300 );
nor  g06984 ( new_n9333 , n22619 , new_n9332 );
xnor g06985 ( new_n9334 , new_n4242 , n24323 );
not  g06986 ( new_n9335 , new_n9334 );
nor  g06987 ( new_n9336 , new_n6003 , new_n9335 );
xnor g06988 ( new_n9337 , n22619 , new_n9332 );
nor  g06989 ( new_n9338 , new_n9336 , new_n9337 );
or   g06990 ( new_n9339 , new_n9333 , new_n9338 );
not  g06991 ( new_n9340 , new_n9330 );
xnor g06992 ( new_n9341 , n26882 , new_n9340 );
nor  g06993 ( new_n9342 , new_n9339 , new_n9341 );
nor  g06994 ( new_n9343 , new_n9331 , new_n9342 );
nor  g06995 ( new_n9344_1 , new_n9328 , new_n9343 );
nor  g06996 ( new_n9345 , new_n9326 , new_n9344_1 );
nor  g06997 ( new_n9346 , new_n9323_1 , new_n9345 );
nor  g06998 ( new_n9347 , new_n9321 , new_n9346 );
nor  g06999 ( new_n9348 , new_n9318_1 , new_n9347 );
nor  g07000 ( new_n9349 , new_n9316 , new_n9348 );
xnor g07001 ( new_n9350 , new_n9313 , new_n9349 );
not  g07002 ( new_n9351 , new_n9350 );
xnor g07003 ( new_n9352 , new_n9287_1 , new_n9351 );
xor  g07004 ( new_n9353 , new_n9253 , new_n9284 );
xnor g07005 ( new_n9354 , new_n9318_1 , new_n9347 );
not  g07006 ( new_n9355 , new_n9354 );
and  g07007 ( new_n9356 , new_n9353 , new_n9355 );
xnor g07008 ( new_n9357 , new_n9353 , new_n9355 );
xor  g07009 ( new_n9358 , new_n9258 , new_n9282 );
xnor g07010 ( new_n9359 , new_n9323_1 , new_n9345 );
not  g07011 ( new_n9360 , new_n9359 );
and  g07012 ( new_n9361 , new_n9358 , new_n9360 );
xnor g07013 ( new_n9362 , new_n9358 , new_n9360 );
xor  g07014 ( new_n9363 , new_n9263 , new_n9280 );
xnor g07015 ( new_n9364_1 , new_n9328 , new_n9343 );
not  g07016 ( new_n9365 , new_n9364_1 );
and  g07017 ( new_n9366 , new_n9363 , new_n9365 );
xnor g07018 ( new_n9367 , new_n9363 , new_n9365 );
xnor g07019 ( new_n9368 , new_n9277 , new_n9278 );
not  g07020 ( new_n9369 , new_n9368 );
xor  g07021 ( new_n9370 , new_n9339 , new_n9341 );
and  g07022 ( new_n9371_1 , new_n9369 , new_n9370 );
xnor g07023 ( new_n9372_1 , new_n9369 , new_n9370 );
xor  g07024 ( new_n9373 , new_n9336 , new_n9337 );
xor  g07025 ( new_n9374 , new_n9273 , new_n9275 );
nor  g07026 ( new_n9375 , new_n9373 , new_n9374 );
xnor g07027 ( new_n9376 , n6775 , new_n9335 );
not  g07028 ( new_n9377 , new_n9376 );
xnor g07029 ( new_n9378 , n15780 , new_n9272 );
nor  g07030 ( new_n9379 , new_n9377 , new_n9378 );
not  g07031 ( new_n9380_1 , new_n9373 );
xnor g07032 ( new_n9381 , new_n9380_1 , new_n9374 );
and  g07033 ( new_n9382_1 , new_n9379 , new_n9381 );
nor  g07034 ( new_n9383 , new_n9375 , new_n9382_1 );
nor  g07035 ( new_n9384 , new_n9372_1 , new_n9383 );
nor  g07036 ( new_n9385 , new_n9371_1 , new_n9384 );
nor  g07037 ( new_n9386 , new_n9367 , new_n9385 );
nor  g07038 ( new_n9387 , new_n9366 , new_n9386 );
nor  g07039 ( new_n9388 , new_n9362 , new_n9387 );
nor  g07040 ( new_n9389 , new_n9361 , new_n9388 );
nor  g07041 ( new_n9390 , new_n9357 , new_n9389 );
nor  g07042 ( new_n9391 , new_n9356 , new_n9390 );
xnor g07043 ( n1044 , new_n9352 , new_n9391 );
nor  g07044 ( new_n9393 , n6775 , n22619 );
not  g07045 ( new_n9394 , new_n9393 );
nor  g07046 ( new_n9395 , n26882 , new_n9394 );
xnor g07047 ( new_n9396_1 , n20478 , new_n9395 );
xnor g07048 ( new_n9397 , new_n4932 , new_n9396_1 );
xnor g07049 ( new_n9398 , n26882 , new_n9393 );
and  g07050 ( new_n9399_1 , n25872 , new_n9398 );
xnor g07051 ( new_n9400 , new_n8483 , new_n9398 );
xnor g07052 ( new_n9401 , n6775 , n22619 );
nor  g07053 ( new_n9402 , new_n4939_1 , new_n9401 );
nor  g07054 ( new_n9403_1 , new_n5002 , new_n6003 );
xnor g07055 ( new_n9404 , n20259 , new_n9401 );
and  g07056 ( new_n9405 , new_n9403_1 , new_n9404 );
or   g07057 ( new_n9406 , new_n9402 , new_n9405 );
and  g07058 ( new_n9407 , new_n9400 , new_n9406 );
nor  g07059 ( new_n9408 , new_n9399_1 , new_n9407 );
xnor g07060 ( new_n9409 , new_n9397 , new_n9408 );
nor  g07061 ( new_n9410 , n2088 , n9399 );
not  g07062 ( new_n9411 , new_n9410 );
nor  g07063 ( new_n9412 , n16396 , new_n9411 );
xnor g07064 ( new_n9413 , n25074 , new_n9412 );
xnor g07065 ( new_n9414 , new_n2398 , new_n9413 );
xnor g07066 ( new_n9415 , n16396 , new_n9410 );
and  g07067 ( new_n9416 , n16722 , new_n9415 );
xnor g07068 ( new_n9417 , new_n7625 , new_n9415 );
not  g07069 ( new_n9418 , new_n5781 );
and  g07070 ( new_n9419_1 , new_n9418 , new_n5787 );
nor  g07071 ( new_n9420 , new_n5783 , new_n9419_1 );
and  g07072 ( new_n9421 , new_n9417 , new_n9420 );
nor  g07073 ( new_n9422 , new_n9416 , new_n9421 );
xnor g07074 ( new_n9423_1 , new_n9414 , new_n9422 );
xnor g07075 ( new_n9424 , new_n9409 , new_n9423_1 );
xnor g07076 ( new_n9425 , new_n9417 , new_n9420 );
nor  g07077 ( new_n9426 , new_n9402 , new_n9405 );
xnor g07078 ( new_n9427 , new_n9400 , new_n9426 );
not  g07079 ( new_n9428 , new_n9427 );
nor  g07080 ( new_n9429 , new_n9425 , new_n9428 );
xnor g07081 ( new_n9430_1 , new_n9425 , new_n9428 );
xnor g07082 ( new_n9431 , new_n9403_1 , new_n9404 );
nor  g07083 ( new_n9432 , new_n5788 , new_n9431 );
xnor g07084 ( new_n9433 , new_n5002 , n6775 );
not  g07085 ( new_n9434 , new_n9433 );
nor  g07086 ( new_n9435_1 , new_n5775 , new_n9434 );
xnor g07087 ( new_n9436 , new_n5789 , new_n9431 );
and  g07088 ( new_n9437 , new_n9435_1 , new_n9436 );
nor  g07089 ( new_n9438 , new_n9432 , new_n9437 );
nor  g07090 ( new_n9439 , new_n9430_1 , new_n9438 );
nor  g07091 ( new_n9440 , new_n9429 , new_n9439 );
xor  g07092 ( new_n9441 , new_n9424 , new_n9440 );
xnor g07093 ( new_n9442 , n7057 , n12956 );
nor  g07094 ( new_n9443 , n8381 , new_n2903 );
nor  g07095 ( new_n9444 , new_n8510_1 , n18295 );
nor  g07096 ( new_n9445_1 , new_n5033 , n20235 );
or   g07097 ( new_n9446 , n6502 , new_n5040 );
nor  g07098 ( new_n9447 , n12495 , new_n2907 );
and  g07099 ( new_n9448 , new_n9446 , new_n9447 );
nor  g07100 ( new_n9449 , new_n9445_1 , new_n9448 );
nor  g07101 ( new_n9450 , new_n9444 , new_n9449 );
or   g07102 ( new_n9451_1 , new_n9443 , new_n9450 );
xnor g07103 ( new_n9452 , new_n9442 , new_n9451_1 );
xor  g07104 ( new_n9453 , new_n9441 , new_n9452 );
xor  g07105 ( new_n9454 , new_n9430_1 , new_n9438 );
not  g07106 ( new_n9455 , new_n9454 );
xnor g07107 ( new_n9456 , n8381 , n18295 );
xnor g07108 ( new_n9457 , new_n9449 , new_n9456 );
and  g07109 ( new_n9458_1 , new_n9455 , new_n9457 );
xnor g07110 ( new_n9459_1 , new_n9455 , new_n9457 );
xnor g07111 ( new_n9460_1 , n12495 , n15780 );
xnor g07112 ( new_n9461 , new_n5775 , new_n9433 );
not  g07113 ( new_n9462 , new_n9461 );
nor  g07114 ( new_n9463 , new_n9460_1 , new_n9462 );
xnor g07115 ( new_n9464 , n6502 , n20235 );
xnor g07116 ( new_n9465 , new_n9447 , new_n9464 );
nor  g07117 ( new_n9466 , new_n9463 , new_n9465 );
xnor g07118 ( new_n9467 , new_n9435_1 , new_n9436 );
not  g07119 ( new_n9468 , new_n9467 );
xnor g07120 ( new_n9469 , new_n9463 , new_n9465 );
nor  g07121 ( new_n9470 , new_n9468 , new_n9469 );
nor  g07122 ( new_n9471 , new_n9466 , new_n9470 );
nor  g07123 ( new_n9472 , new_n9459_1 , new_n9471 );
nor  g07124 ( new_n9473 , new_n9458_1 , new_n9472 );
xor  g07125 ( n1060 , new_n9453 , new_n9473 );
xnor g07126 ( n1069 , new_n3348 , new_n3385 );
not  g07127 ( new_n9476 , n3959 );
xnor g07128 ( new_n9477 , new_n9476 , n9832 );
nor  g07129 ( new_n9478 , n1558 , n11566 );
not  g07130 ( new_n9479 , n1558 );
xnor g07131 ( new_n9480 , new_n9479 , n11566 );
nor  g07132 ( new_n9481 , n21749 , n26744 );
xnor g07133 ( new_n9482 , n21749 , n26744 );
nor  g07134 ( new_n9483 , n7769 , n26625 );
not  g07135 ( new_n9484 , n14230 );
not  g07136 ( new_n9485 , n21138 );
or   g07137 ( new_n9486 , new_n9484 , new_n9485 );
not  g07138 ( new_n9487 , n7769 );
xnor g07139 ( new_n9488 , new_n9487 , n26625 );
and  g07140 ( new_n9489 , new_n9486 , new_n9488 );
nor  g07141 ( new_n9490 , new_n9483 , new_n9489 );
nor  g07142 ( new_n9491 , new_n9482 , new_n9490 );
or   g07143 ( new_n9492 , new_n9481 , new_n9491 );
and  g07144 ( new_n9493_1 , new_n9480 , new_n9492 );
nor  g07145 ( new_n9494 , new_n9478 , new_n9493_1 );
xnor g07146 ( new_n9495 , new_n9477 , new_n9494 );
nor  g07147 ( new_n9496 , n22591 , n26167 );
not  g07148 ( new_n9497 , new_n9496 );
nor  g07149 ( new_n9498 , n17095 , new_n9497 );
not  g07150 ( new_n9499 , new_n9498 );
nor  g07151 ( new_n9500 , n15378 , new_n9499 );
xnor g07152 ( new_n9501 , n19575 , new_n9500 );
not  g07153 ( new_n9502 , n5226 );
xnor g07154 ( new_n9503 , new_n9502 , new_n6802_1 );
nor  g07155 ( new_n9504 , new_n2574 , new_n6806 );
xnor g07156 ( new_n9505 , new_n2574 , new_n6806 );
nor  g07157 ( new_n9506 , new_n2578_1 , new_n6809 );
xnor g07158 ( new_n9507_1 , new_n2578_1 , new_n6809 );
nor  g07159 ( new_n9508_1 , n1136 , new_n6942 );
nor  g07160 ( new_n9509 , new_n2582_1 , new_n6812 );
xnor g07161 ( new_n9510 , n1136 , new_n6942 );
nor  g07162 ( new_n9511 , new_n9509 , new_n9510 );
or   g07163 ( new_n9512_1 , new_n9508_1 , new_n9511 );
nor  g07164 ( new_n9513 , new_n9507_1 , new_n9512_1 );
nor  g07165 ( new_n9514 , new_n9506 , new_n9513 );
nor  g07166 ( new_n9515 , new_n9505 , new_n9514 );
nor  g07167 ( new_n9516 , new_n9504 , new_n9515 );
xor  g07168 ( new_n9517 , new_n9503 , new_n9516 );
not  g07169 ( new_n9518 , new_n9517 );
xnor g07170 ( new_n9519 , new_n9501 , new_n9518 );
xor  g07171 ( new_n9520 , new_n9505 , new_n9514 );
xnor g07172 ( new_n9521 , n15378 , new_n9498 );
nor  g07173 ( new_n9522 , new_n9520 , new_n9521 );
xnor g07174 ( new_n9523 , new_n9520 , new_n9521 );
nor  g07175 ( new_n9524 , new_n9508_1 , new_n9511 );
xnor g07176 ( new_n9525 , new_n9507_1 , new_n9524 );
xnor g07177 ( new_n9526 , n17095 , new_n9496 );
nor  g07178 ( new_n9527 , new_n9525 , new_n9526 );
not  g07179 ( new_n9528 , new_n9525 );
xnor g07180 ( new_n9529 , new_n9528 , new_n9526 );
xnor g07181 ( new_n9530 , new_n9509 , new_n9510 );
not  g07182 ( new_n9531 , n22591 );
not  g07183 ( new_n9532 , n26167 );
nor  g07184 ( new_n9533 , new_n9532 , new_n7199 );
xnor g07185 ( new_n9534 , new_n9531 , new_n9533 );
and  g07186 ( new_n9535 , new_n9530 , new_n9534 );
or   g07187 ( new_n9536 , new_n9532 , new_n7200 );
nor  g07188 ( new_n9537 , n22591 , new_n9536 );
nor  g07189 ( new_n9538 , new_n9535 , new_n9537 );
and  g07190 ( new_n9539 , new_n9529 , new_n9538 );
nor  g07191 ( new_n9540 , new_n9527 , new_n9539 );
nor  g07192 ( new_n9541 , new_n9523 , new_n9540 );
or   g07193 ( new_n9542 , new_n9522 , new_n9541 );
xor  g07194 ( new_n9543 , new_n9519 , new_n9542 );
xnor g07195 ( new_n9544 , new_n9495 , new_n9543 );
xnor g07196 ( new_n9545 , new_n9523 , new_n9540 );
xor  g07197 ( new_n9546 , new_n9480 , new_n9492 );
nor  g07198 ( new_n9547 , new_n9545 , new_n9546 );
xnor g07199 ( new_n9548 , new_n9545 , new_n9546 );
not  g07200 ( new_n9549 , new_n9548 );
xor  g07201 ( new_n9550 , new_n9529 , new_n9538 );
xnor g07202 ( new_n9551 , new_n9482 , new_n9490 );
nor  g07203 ( new_n9552_1 , new_n9550 , new_n9551 );
xor  g07204 ( new_n9553 , new_n9550 , new_n9551 );
not  g07205 ( new_n9554_1 , new_n9530 );
xnor g07206 ( new_n9555 , new_n9554_1 , new_n9534 );
nor  g07207 ( new_n9556_1 , new_n9484 , new_n9485 );
xnor g07208 ( new_n9557_1 , new_n9556_1 , new_n9488 );
nor  g07209 ( new_n9558_1 , new_n9555 , new_n9557_1 );
nor  g07210 ( new_n9559 , new_n7198 , new_n7201 );
not  g07211 ( new_n9560 , new_n9557_1 );
xnor g07212 ( new_n9561 , new_n9555 , new_n9560 );
and  g07213 ( new_n9562 , new_n9559 , new_n9561 );
nor  g07214 ( new_n9563 , new_n9558_1 , new_n9562 );
and  g07215 ( new_n9564 , new_n9553 , new_n9563 );
nor  g07216 ( new_n9565 , new_n9552_1 , new_n9564 );
and  g07217 ( new_n9566 , new_n9549 , new_n9565 );
nor  g07218 ( new_n9567 , new_n9547 , new_n9566 );
xor  g07219 ( n1111 , new_n9544 , new_n9567 );
xnor g07220 ( new_n9569 , new_n4431 , new_n2607 );
nor  g07221 ( new_n9570 , new_n4435 , new_n2611 );
xnor g07222 ( new_n9571 , new_n4435 , new_n2611 );
nor  g07223 ( new_n9572 , new_n4442 , new_n2647 );
nor  g07224 ( new_n9573 , n11011 , new_n2615 );
xnor g07225 ( new_n9574 , n11011 , new_n2615 );
nor  g07226 ( new_n9575 , n16029 , new_n2618 );
xnor g07227 ( new_n9576 , new_n3939 , new_n2618 );
nor  g07228 ( new_n9577 , new_n3943 , new_n2623 );
xnor g07229 ( new_n9578 , new_n3943 , new_n2623 );
nor  g07230 ( new_n9579 , new_n3947 , new_n2636 );
nor  g07231 ( new_n9580 , n22433 , new_n2627 );
nor  g07232 ( new_n9581 , new_n3952_1 , new_n2630 );
xnor g07233 ( new_n9582 , n22433 , new_n2627 );
nor  g07234 ( new_n9583 , new_n9581 , new_n9582 );
nor  g07235 ( new_n9584 , new_n9580 , new_n9583 );
xnor g07236 ( new_n9585 , n11615 , new_n2636 );
and  g07237 ( new_n9586 , new_n9584 , new_n9585 );
nor  g07238 ( new_n9587 , new_n9579 , new_n9586 );
nor  g07239 ( new_n9588 , new_n9578 , new_n9587 );
nor  g07240 ( new_n9589 , new_n9577 , new_n9588 );
and  g07241 ( new_n9590 , new_n9576 , new_n9589 );
nor  g07242 ( new_n9591 , new_n9575 , new_n9590 );
nor  g07243 ( new_n9592 , new_n9574 , new_n9591 );
or   g07244 ( new_n9593 , new_n9573 , new_n9592 );
xnor g07245 ( new_n9594 , new_n4442 , new_n2647 );
nor  g07246 ( new_n9595 , new_n9593 , new_n9594 );
nor  g07247 ( new_n9596 , new_n9572 , new_n9595 );
nor  g07248 ( new_n9597 , new_n9571 , new_n9596 );
nor  g07249 ( new_n9598_1 , new_n9570 , new_n9597 );
xor  g07250 ( new_n9599 , new_n9569 , new_n9598_1 );
not  g07251 ( new_n9600 , new_n9599 );
not  g07252 ( new_n9601 , new_n9412 );
nor  g07253 ( new_n9602 , n25074 , new_n9601 );
not  g07254 ( new_n9603 , new_n9602 );
nor  g07255 ( new_n9604 , n8006 , new_n9603 );
not  g07256 ( new_n9605 , new_n9604 );
nor  g07257 ( new_n9606 , n20929 , new_n9605 );
not  g07258 ( new_n9607 , new_n9606 );
nor  g07259 ( new_n9608 , n10710 , new_n9607 );
not  g07260 ( new_n9609 , new_n9608 );
nor  g07261 ( new_n9610 , n11841 , new_n9609 );
xnor g07262 ( new_n9611 , n27089 , new_n9610 );
xnor g07263 ( new_n9612 , new_n2725 , new_n9611 );
xnor g07264 ( new_n9613 , n11841 , new_n9608 );
and  g07265 ( new_n9614 , new_n2729 , new_n9613 );
not  g07266 ( new_n9615 , new_n2729 );
xnor g07267 ( new_n9616_1 , new_n9615 , new_n9613 );
xnor g07268 ( new_n9617 , n10710 , new_n9606 );
nor  g07269 ( new_n9618 , new_n2733 , new_n9617 );
xnor g07270 ( new_n9619 , new_n2733 , new_n9617 );
xnor g07271 ( new_n9620 , n20929 , new_n9604 );
nor  g07272 ( new_n9621 , new_n2738 , new_n9620 );
xnor g07273 ( new_n9622_1 , new_n2740 , new_n9620 );
xnor g07274 ( new_n9623 , n8006 , new_n9602 );
nor  g07275 ( new_n9624 , new_n2744 , new_n9623 );
nor  g07276 ( new_n9625 , new_n2748 , new_n9413 );
not  g07277 ( new_n9626_1 , new_n2748 );
xnor g07278 ( new_n9627 , new_n9626_1 , new_n9413 );
nor  g07279 ( new_n9628 , new_n2753 , new_n9415 );
not  g07280 ( new_n9629 , new_n2753 );
xnor g07281 ( new_n9630 , new_n9629 , new_n9415 );
nor  g07282 ( new_n9631 , new_n2759 , new_n5781 );
nor  g07283 ( new_n9632 , n2088 , new_n2761_1 );
xnor g07284 ( new_n9633_1 , new_n2763 , new_n5781 );
and  g07285 ( new_n9634 , new_n9632 , new_n9633_1 );
or   g07286 ( new_n9635_1 , new_n9631 , new_n9634 );
and  g07287 ( new_n9636 , new_n9630 , new_n9635_1 );
or   g07288 ( new_n9637 , new_n9628 , new_n9636 );
and  g07289 ( new_n9638 , new_n9627 , new_n9637 );
or   g07290 ( new_n9639 , new_n9625 , new_n9638 );
xnor g07291 ( new_n9640 , new_n2771 , new_n9623 );
and  g07292 ( new_n9641 , new_n9639 , new_n9640 );
or   g07293 ( new_n9642 , new_n9624 , new_n9641 );
and  g07294 ( new_n9643 , new_n9622_1 , new_n9642 );
nor  g07295 ( new_n9644 , new_n9621 , new_n9643 );
nor  g07296 ( new_n9645 , new_n9619 , new_n9644 );
nor  g07297 ( new_n9646_1 , new_n9618 , new_n9645 );
and  g07298 ( new_n9647 , new_n9616_1 , new_n9646_1 );
or   g07299 ( new_n9648_1 , new_n9614 , new_n9647 );
xor  g07300 ( new_n9649 , new_n9612 , new_n9648_1 );
xnor g07301 ( new_n9650 , new_n9600 , new_n9649 );
xor  g07302 ( new_n9651 , new_n9571 , new_n9596 );
not  g07303 ( new_n9652 , new_n9651 );
xnor g07304 ( new_n9653 , new_n9616_1 , new_n9646_1 );
nor  g07305 ( new_n9654 , new_n9652 , new_n9653 );
xnor g07306 ( new_n9655_1 , new_n9651 , new_n9653 );
nor  g07307 ( new_n9656 , new_n9573 , new_n9592 );
xnor g07308 ( new_n9657 , new_n9656 , new_n9594 );
xnor g07309 ( new_n9658 , new_n9619 , new_n9644 );
nor  g07310 ( new_n9659 , new_n9657 , new_n9658 );
not  g07311 ( new_n9660 , new_n9657 );
xnor g07312 ( new_n9661 , new_n9660 , new_n9658 );
xnor g07313 ( new_n9662 , new_n9574 , new_n9591 );
not  g07314 ( new_n9663 , new_n9662 );
xor  g07315 ( new_n9664 , new_n9622_1 , new_n9642 );
nor  g07316 ( new_n9665 , new_n9663 , new_n9664 );
xnor g07317 ( new_n9666 , new_n9662 , new_n9664 );
xnor g07318 ( new_n9667 , new_n9576 , new_n9589 );
not  g07319 ( new_n9668 , new_n9667 );
xor  g07320 ( new_n9669 , new_n9639 , new_n9640 );
nor  g07321 ( new_n9670 , new_n9668 , new_n9669 );
xnor g07322 ( new_n9671 , new_n9667 , new_n9669 );
xor  g07323 ( new_n9672 , new_n9627 , new_n9637 );
xnor g07324 ( new_n9673 , new_n9578 , new_n9587 );
nor  g07325 ( new_n9674 , new_n9672 , new_n9673 );
not  g07326 ( new_n9675 , new_n9673 );
xnor g07327 ( new_n9676 , new_n9672 , new_n9675 );
xor  g07328 ( new_n9677 , new_n9630 , new_n9635_1 );
xnor g07329 ( new_n9678 , new_n9584 , new_n9585 );
nor  g07330 ( new_n9679 , new_n9677 , new_n9678 );
not  g07331 ( new_n9680 , new_n9678 );
xnor g07332 ( new_n9681 , new_n9677 , new_n9680 );
xnor g07333 ( new_n9682 , new_n9632 , new_n9633_1 );
xnor g07334 ( new_n9683 , new_n9581 , new_n9582 );
nor  g07335 ( new_n9684 , new_n9682 , new_n9683 );
xnor g07336 ( new_n9685 , n14090 , new_n2630 );
not  g07337 ( new_n9686 , new_n9685 );
xnor g07338 ( new_n9687 , new_n2951 , new_n2761_1 );
nor  g07339 ( new_n9688 , new_n9686 , new_n9687 );
xnor g07340 ( new_n9689_1 , new_n9682 , new_n9683 );
nor  g07341 ( new_n9690 , new_n9688 , new_n9689_1 );
nor  g07342 ( new_n9691 , new_n9684 , new_n9690 );
and  g07343 ( new_n9692 , new_n9681 , new_n9691 );
or   g07344 ( new_n9693 , new_n9679 , new_n9692 );
and  g07345 ( new_n9694 , new_n9676 , new_n9693 );
or   g07346 ( new_n9695_1 , new_n9674 , new_n9694 );
and  g07347 ( new_n9696 , new_n9671 , new_n9695_1 );
or   g07348 ( new_n9697 , new_n9670 , new_n9696 );
and  g07349 ( new_n9698 , new_n9666 , new_n9697 );
nor  g07350 ( new_n9699_1 , new_n9665 , new_n9698 );
and  g07351 ( new_n9700 , new_n9661 , new_n9699_1 );
nor  g07352 ( new_n9701 , new_n9659 , new_n9700 );
and  g07353 ( new_n9702 , new_n9655_1 , new_n9701 );
nor  g07354 ( new_n9703 , new_n9654 , new_n9702 );
xnor g07355 ( n1119 , new_n9650 , new_n9703 );
xnor g07356 ( new_n9705 , new_n7879 , new_n7877 );
xnor g07357 ( n1120 , new_n7902 , new_n9705 );
xnor g07358 ( new_n9707 , n3925 , n9246 );
xnor g07359 ( new_n9708 , new_n7749 , new_n9707 );
not  g07360 ( new_n9709 , new_n9708 );
xnor g07361 ( new_n9710 , n7428 , n12495 );
xnor g07362 ( n1196 , new_n9709 , new_n9710 );
xnor g07363 ( new_n9712 , n15636 , n16223 );
nor  g07364 ( new_n9713 , n19494 , new_n2444_1 );
or   g07365 ( new_n9714 , new_n2365 , n20077 );
nor  g07366 ( new_n9715 , n2387 , new_n2447 );
and  g07367 ( new_n9716 , new_n9714 , new_n9715 );
or   g07368 ( new_n9717 , new_n9713 , new_n9716 );
xor  g07369 ( new_n9718 , new_n9712 , new_n9717 );
xnor g07370 ( new_n9719 , new_n7882 , new_n9718 );
xnor g07371 ( new_n9720 , n2387 , n6794 );
nor  g07372 ( new_n9721 , new_n7890 , new_n9720 );
xnor g07373 ( new_n9722 , n19494 , n20077 );
xnor g07374 ( new_n9723 , new_n9715 , new_n9722 );
nor  g07375 ( new_n9724 , new_n9721 , new_n9723 );
xnor g07376 ( new_n9725 , new_n9721 , new_n9723 );
nor  g07377 ( new_n9726_1 , new_n7884_1 , new_n9725 );
nor  g07378 ( new_n9727 , new_n9724 , new_n9726_1 );
xnor g07379 ( n1237 , new_n9719 , new_n9727 );
xnor g07380 ( new_n9729 , new_n5498 , new_n5702 );
xnor g07381 ( n1239 , new_n5765_1 , new_n9729 );
xnor g07382 ( new_n9731 , n1536 , n22764 );
nor  g07383 ( new_n9732 , n19454 , n26264 );
xnor g07384 ( new_n9733 , n19454 , n26264 );
nor  g07385 ( new_n9734 , n7841 , n9445 );
xnor g07386 ( new_n9735 , n7841 , n9445 );
nor  g07387 ( new_n9736 , n1279 , n16812 );
xnor g07388 ( new_n9737 , n1279 , n16812 );
nor  g07389 ( new_n9738 , n8324 , n25068 );
xnor g07390 ( new_n9739 , n8324 , n25068 );
nor  g07391 ( new_n9740 , n2331 , n12546 );
xnor g07392 ( new_n9741 , n2331 , n12546 );
nor  g07393 ( new_n9742 , n21078 , n22631 );
xnor g07394 ( new_n9743 , n21078 , n22631 );
nor  g07395 ( new_n9744 , n16743 , n24485 );
xnor g07396 ( new_n9745 , n16743 , n24485 );
nor  g07397 ( new_n9746 , n2420 , n15258 );
nor  g07398 ( new_n9747 , new_n2542 , new_n8110 );
xnor g07399 ( new_n9748 , n2420 , n15258 );
nor  g07400 ( new_n9749 , new_n9747 , new_n9748 );
nor  g07401 ( new_n9750 , new_n9746 , new_n9749 );
nor  g07402 ( new_n9751 , new_n9745 , new_n9750 );
nor  g07403 ( new_n9752 , new_n9744 , new_n9751 );
nor  g07404 ( new_n9753_1 , new_n9743 , new_n9752 );
nor  g07405 ( new_n9754 , new_n9742 , new_n9753_1 );
nor  g07406 ( new_n9755 , new_n9741 , new_n9754 );
nor  g07407 ( new_n9756 , new_n9740 , new_n9755 );
nor  g07408 ( new_n9757 , new_n9739 , new_n9756 );
nor  g07409 ( new_n9758 , new_n9738 , new_n9757 );
nor  g07410 ( new_n9759 , new_n9737 , new_n9758 );
nor  g07411 ( new_n9760 , new_n9736 , new_n9759 );
nor  g07412 ( new_n9761_1 , new_n9735 , new_n9760 );
nor  g07413 ( new_n9762 , new_n9734 , new_n9761_1 );
nor  g07414 ( new_n9763_1 , new_n9733 , new_n9762 );
nor  g07415 ( new_n9764 , new_n9732 , new_n9763_1 );
xnor g07416 ( new_n9765 , new_n9731 , new_n9764 );
nor  g07417 ( new_n9766 , n2416 , new_n9765 );
xnor g07418 ( new_n9767_1 , n2416 , new_n9765 );
xnor g07419 ( new_n9768 , new_n9733 , new_n9762 );
nor  g07420 ( new_n9769 , n21905 , new_n9768 );
xnor g07421 ( new_n9770 , n21905 , new_n9768 );
xnor g07422 ( new_n9771_1 , new_n9735 , new_n9760 );
nor  g07423 ( new_n9772 , n22918 , new_n9771_1 );
xnor g07424 ( new_n9773 , n22918 , new_n9771_1 );
xnor g07425 ( new_n9774 , new_n9737 , new_n9758 );
nor  g07426 ( new_n9775 , n25923 , new_n9774 );
xnor g07427 ( new_n9776 , n25923 , new_n9774 );
xnor g07428 ( new_n9777 , new_n9739 , new_n9756 );
nor  g07429 ( new_n9778_1 , n6790 , new_n9777 );
xnor g07430 ( new_n9779 , n6790 , new_n9777 );
xnor g07431 ( new_n9780 , new_n9741 , new_n9754 );
nor  g07432 ( new_n9781 , n22879 , new_n9780 );
xnor g07433 ( new_n9782 , n22879 , new_n9780 );
xnor g07434 ( new_n9783_1 , new_n9743 , new_n9752 );
nor  g07435 ( new_n9784 , n2117 , new_n9783_1 );
xnor g07436 ( new_n9785 , n2117 , new_n9783_1 );
xnor g07437 ( new_n9786 , new_n9745 , new_n9750 );
nor  g07438 ( new_n9787 , n5882 , new_n9786 );
xnor g07439 ( new_n9788 , new_n9747 , new_n9748 );
nor  g07440 ( new_n9789 , n11775 , new_n9788 );
not  g07441 ( new_n9790 , n27134 );
xnor g07442 ( new_n9791 , n4588 , n22201 );
or   g07443 ( new_n9792 , new_n9790 , new_n9791 );
not  g07444 ( new_n9793 , n11775 );
xnor g07445 ( new_n9794 , new_n9793 , new_n9788 );
and  g07446 ( new_n9795 , new_n9792 , new_n9794 );
nor  g07447 ( new_n9796 , new_n9789 , new_n9795 );
xnor g07448 ( new_n9797 , n5882 , new_n9786 );
nor  g07449 ( new_n9798 , new_n9796 , new_n9797 );
nor  g07450 ( new_n9799 , new_n9787 , new_n9798 );
nor  g07451 ( new_n9800 , new_n9785 , new_n9799 );
nor  g07452 ( new_n9801 , new_n9784 , new_n9800 );
nor  g07453 ( new_n9802 , new_n9782 , new_n9801 );
nor  g07454 ( new_n9803_1 , new_n9781 , new_n9802 );
nor  g07455 ( new_n9804 , new_n9779 , new_n9803_1 );
nor  g07456 ( new_n9805 , new_n9778_1 , new_n9804 );
nor  g07457 ( new_n9806 , new_n9776 , new_n9805 );
nor  g07458 ( new_n9807 , new_n9775 , new_n9806 );
nor  g07459 ( new_n9808 , new_n9773 , new_n9807 );
nor  g07460 ( new_n9809 , new_n9772 , new_n9808 );
nor  g07461 ( new_n9810 , new_n9770 , new_n9809 );
nor  g07462 ( new_n9811 , new_n9769 , new_n9810 );
nor  g07463 ( new_n9812 , new_n9767_1 , new_n9811 );
nor  g07464 ( new_n9813 , new_n9766 , new_n9812 );
nor  g07465 ( new_n9814 , n1536 , n22764 );
nor  g07466 ( new_n9815 , new_n9731 , new_n9764 );
nor  g07467 ( new_n9816 , new_n9814 , new_n9815 );
and  g07468 ( new_n9817 , new_n9813 , new_n9816 );
nor  g07469 ( new_n9818 , n8405 , n23493 );
nor  g07470 ( new_n9819 , n10275 , n22359 );
nor  g07471 ( new_n9820 , n5532 , n15146 );
nor  g07472 ( new_n9821 , n3962 , n11579 );
nor  g07473 ( new_n9822 , n21 , n23513 );
xnor g07474 ( new_n9823 , n21 , n23513 );
nor  g07475 ( new_n9824 , n1682 , n6427 );
and  g07476 ( new_n9825 , n1682 , n6427 );
nor  g07477 ( new_n9826 , n6590 , n7963 );
nor  g07478 ( new_n9827 , n10017 , n20349 );
not  g07479 ( new_n9828 , n15936 );
nor  g07480 ( new_n9829 , new_n7939 , new_n9828 );
not  g07481 ( new_n9830 , n20349 );
nor  g07482 ( new_n9831 , new_n7941 , new_n9830 );
nor  g07483 ( new_n9832_1 , new_n9829 , new_n9831 );
nor  g07484 ( new_n9833_1 , new_n9827 , new_n9832_1 );
not  g07485 ( new_n9834 , n6590 );
not  g07486 ( new_n9835 , n7963 );
nor  g07487 ( new_n9836 , new_n9834 , new_n9835 );
nor  g07488 ( new_n9837 , new_n9833_1 , new_n9836 );
nor  g07489 ( new_n9838_1 , new_n9826 , new_n9837 );
nor  g07490 ( new_n9839 , new_n9825 , new_n9838_1 );
nor  g07491 ( new_n9840 , new_n9824 , new_n9839 );
nor  g07492 ( new_n9841 , new_n9823 , new_n9840 );
nor  g07493 ( new_n9842 , new_n9822 , new_n9841 );
xnor g07494 ( new_n9843 , n3962 , n11579 );
nor  g07495 ( new_n9844 , new_n9842 , new_n9843 );
nor  g07496 ( new_n9845 , new_n9821 , new_n9844 );
xnor g07497 ( new_n9846 , n5532 , n15146 );
nor  g07498 ( new_n9847 , new_n9845 , new_n9846 );
nor  g07499 ( new_n9848 , new_n9820 , new_n9847 );
xnor g07500 ( new_n9849 , n10275 , n22359 );
nor  g07501 ( new_n9850 , new_n9848 , new_n9849 );
nor  g07502 ( new_n9851 , new_n9819 , new_n9850 );
xnor g07503 ( new_n9852 , n8405 , n23493 );
nor  g07504 ( new_n9853 , new_n9851 , new_n9852 );
nor  g07505 ( new_n9854 , new_n9818 , new_n9853 );
xnor g07506 ( new_n9855 , n13549 , n14826 );
xnor g07507 ( new_n9856 , new_n9854 , new_n9855 );
nor  g07508 ( new_n9857 , n18105 , new_n9856 );
xnor g07509 ( new_n9858 , n18105 , new_n9856 );
xnor g07510 ( new_n9859 , new_n9851 , new_n9852 );
nor  g07511 ( new_n9860 , n24196 , new_n9859 );
xnor g07512 ( new_n9861 , n24196 , new_n9859 );
xnor g07513 ( new_n9862 , new_n9848 , new_n9849 );
nor  g07514 ( new_n9863 , n16376 , new_n9862 );
xnor g07515 ( new_n9864 , n16376 , new_n9862 );
xnor g07516 ( new_n9865 , new_n9845 , new_n9846 );
nor  g07517 ( new_n9866 , n25381 , new_n9865 );
xnor g07518 ( new_n9867_1 , n25381 , new_n9865 );
xnor g07519 ( new_n9868 , new_n9842 , new_n9843 );
nor  g07520 ( new_n9869 , n12587 , new_n9868 );
xnor g07521 ( new_n9870 , n12587 , new_n9868 );
xnor g07522 ( new_n9871 , new_n9823 , new_n9840 );
nor  g07523 ( new_n9872_1 , n268 , new_n9871 );
xnor g07524 ( new_n9873 , n268 , new_n9871 );
xnor g07525 ( new_n9874 , new_n7934 , n6427 );
not  g07526 ( new_n9875 , new_n9874 );
xnor g07527 ( new_n9876 , new_n9838_1 , new_n9875 );
nor  g07528 ( new_n9877 , n24879 , new_n9876 );
xnor g07529 ( new_n9878 , n24879 , new_n9876 );
xnor g07530 ( new_n9879 , n6590 , n7963 );
xnor g07531 ( new_n9880 , new_n9833_1 , new_n9879 );
nor  g07532 ( new_n9881 , n6785 , new_n9880 );
xnor g07533 ( new_n9882 , n10017 , n20349 );
xnor g07534 ( new_n9883 , new_n9829 , new_n9882 );
nor  g07535 ( new_n9884 , n24032 , new_n9883 );
xnor g07536 ( new_n9885 , n3618 , n15936 );
or   g07537 ( new_n9886 , new_n4507 , new_n9885 );
xnor g07538 ( new_n9887 , new_n8052_1 , new_n9883 );
and  g07539 ( new_n9888 , new_n9886 , new_n9887 );
nor  g07540 ( new_n9889 , new_n9884 , new_n9888 );
xnor g07541 ( new_n9890_1 , n6785 , new_n9880 );
nor  g07542 ( new_n9891 , new_n9889 , new_n9890_1 );
nor  g07543 ( new_n9892 , new_n9881 , new_n9891 );
nor  g07544 ( new_n9893 , new_n9878 , new_n9892 );
nor  g07545 ( new_n9894 , new_n9877 , new_n9893 );
nor  g07546 ( new_n9895 , new_n9873 , new_n9894 );
nor  g07547 ( new_n9896 , new_n9872_1 , new_n9895 );
nor  g07548 ( new_n9897 , new_n9870 , new_n9896 );
nor  g07549 ( new_n9898 , new_n9869 , new_n9897 );
nor  g07550 ( new_n9899 , new_n9867_1 , new_n9898 );
nor  g07551 ( new_n9900 , new_n9866 , new_n9899 );
nor  g07552 ( new_n9901 , new_n9864 , new_n9900 );
nor  g07553 ( new_n9902 , new_n9863 , new_n9901 );
nor  g07554 ( new_n9903 , new_n9861 , new_n9902 );
nor  g07555 ( new_n9904 , new_n9860 , new_n9903 );
nor  g07556 ( new_n9905 , new_n9858 , new_n9904 );
nor  g07557 ( new_n9906 , new_n9857 , new_n9905 );
nor  g07558 ( new_n9907 , new_n9854 , new_n9855 );
nor  g07559 ( new_n9908 , n13549 , n14826 );
nor  g07560 ( new_n9909 , new_n9907 , new_n9908 );
nand g07561 ( new_n9910 , new_n9906 , new_n9909 );
xnor g07562 ( new_n9911 , new_n9817 , new_n9910 );
xnor g07563 ( new_n9912 , new_n9813 , new_n9816 );
xnor g07564 ( new_n9913 , new_n9906 , new_n9909 );
not  g07565 ( new_n9914 , new_n9913 );
and  g07566 ( new_n9915 , new_n9912 , new_n9914 );
xnor g07567 ( new_n9916 , new_n9912 , new_n9914 );
xnor g07568 ( new_n9917_1 , new_n9767_1 , new_n9811 );
xnor g07569 ( new_n9918 , new_n9858 , new_n9904 );
not  g07570 ( new_n9919_1 , new_n9918 );
nor  g07571 ( new_n9920 , new_n9917_1 , new_n9919_1 );
xnor g07572 ( new_n9921 , new_n9917_1 , new_n9919_1 );
xnor g07573 ( new_n9922 , new_n9770 , new_n9809 );
xnor g07574 ( new_n9923 , new_n9861 , new_n9902 );
not  g07575 ( new_n9924 , new_n9923 );
nor  g07576 ( new_n9925 , new_n9922 , new_n9924 );
xnor g07577 ( new_n9926_1 , new_n9922 , new_n9924 );
xnor g07578 ( new_n9927 , new_n9773 , new_n9807 );
xnor g07579 ( new_n9928 , new_n9864 , new_n9900 );
not  g07580 ( new_n9929 , new_n9928 );
nor  g07581 ( new_n9930 , new_n9927 , new_n9929 );
xnor g07582 ( new_n9931 , new_n9927 , new_n9929 );
xnor g07583 ( new_n9932 , new_n9776 , new_n9805 );
xnor g07584 ( new_n9933 , new_n9867_1 , new_n9898 );
not  g07585 ( new_n9934_1 , new_n9933 );
nor  g07586 ( new_n9935 , new_n9932 , new_n9934_1 );
xnor g07587 ( new_n9936 , new_n9932 , new_n9934_1 );
xnor g07588 ( new_n9937 , new_n9779 , new_n9803_1 );
xnor g07589 ( new_n9938_1 , new_n9870 , new_n9896 );
not  g07590 ( new_n9939 , new_n9938_1 );
nor  g07591 ( new_n9940 , new_n9937 , new_n9939 );
xnor g07592 ( new_n9941 , new_n9937 , new_n9939 );
xnor g07593 ( new_n9942_1 , new_n9782 , new_n9801 );
xor  g07594 ( new_n9943 , new_n9873 , new_n9894 );
nor  g07595 ( new_n9944 , new_n9942_1 , new_n9943 );
xnor g07596 ( new_n9945 , new_n9942_1 , new_n9943 );
xnor g07597 ( new_n9946_1 , new_n9785 , new_n9799 );
xnor g07598 ( new_n9947 , new_n9878 , new_n9892 );
not  g07599 ( new_n9948 , new_n9947 );
nor  g07600 ( new_n9949 , new_n9946_1 , new_n9948 );
xnor g07601 ( new_n9950 , new_n9946_1 , new_n9948 );
xnor g07602 ( new_n9951 , new_n9796 , new_n9797 );
xnor g07603 ( new_n9952 , new_n9889 , new_n9890_1 );
not  g07604 ( new_n9953 , new_n9952 );
nor  g07605 ( new_n9954 , new_n9951 , new_n9953 );
xnor g07606 ( new_n9955 , new_n9951 , new_n9953 );
xor  g07607 ( new_n9956 , new_n9792 , new_n9794 );
not  g07608 ( new_n9957 , new_n9956 );
nor  g07609 ( new_n9958 , new_n4507 , new_n9885 );
xnor g07610 ( new_n9959 , new_n9958 , new_n9887 );
nor  g07611 ( new_n9960 , new_n9957 , new_n9959 );
xnor g07612 ( new_n9961 , n27134 , new_n9791 );
xnor g07613 ( new_n9962 , n22843 , new_n9885 );
not  g07614 ( new_n9963 , new_n9962 );
nor  g07615 ( new_n9964 , new_n9961 , new_n9963 );
not  g07616 ( new_n9965 , new_n9959 );
xnor g07617 ( new_n9966 , new_n9957 , new_n9965 );
and  g07618 ( new_n9967_1 , new_n9964 , new_n9966 );
nor  g07619 ( new_n9968_1 , new_n9960 , new_n9967_1 );
nor  g07620 ( new_n9969 , new_n9955 , new_n9968_1 );
nor  g07621 ( new_n9970 , new_n9954 , new_n9969 );
nor  g07622 ( new_n9971 , new_n9950 , new_n9970 );
nor  g07623 ( new_n9972 , new_n9949 , new_n9971 );
nor  g07624 ( new_n9973 , new_n9945 , new_n9972 );
nor  g07625 ( new_n9974 , new_n9944 , new_n9973 );
nor  g07626 ( new_n9975 , new_n9941 , new_n9974 );
nor  g07627 ( new_n9976 , new_n9940 , new_n9975 );
nor  g07628 ( new_n9977 , new_n9936 , new_n9976 );
nor  g07629 ( new_n9978 , new_n9935 , new_n9977 );
nor  g07630 ( new_n9979 , new_n9931 , new_n9978 );
nor  g07631 ( new_n9980 , new_n9930 , new_n9979 );
nor  g07632 ( new_n9981 , new_n9926_1 , new_n9980 );
nor  g07633 ( new_n9982 , new_n9925 , new_n9981 );
nor  g07634 ( new_n9983 , new_n9921 , new_n9982 );
nor  g07635 ( new_n9984 , new_n9920 , new_n9983 );
nor  g07636 ( new_n9985 , new_n9916 , new_n9984 );
nor  g07637 ( new_n9986 , new_n9915 , new_n9985 );
xnor g07638 ( n1302 , new_n9911 , new_n9986 );
nor  g07639 ( new_n9988 , new_n8719 , n13951 );
xnor g07640 ( new_n9989 , n12507 , n13951 );
nor  g07641 ( new_n9990 , new_n8789 , n22793 );
xnor g07642 ( new_n9991 , n15077 , n22793 );
not  g07643 ( new_n9992 , n3710 );
nor  g07644 ( new_n9993 , new_n9992 , n8439 );
xnor g07645 ( new_n9994 , n3710 , n8439 );
nor  g07646 ( new_n9995 , n25523 , new_n8745_1 );
xnor g07647 ( new_n9996 , n25523 , n26318 );
nor  g07648 ( new_n9997 , n5579 , new_n8749 );
xnor g07649 ( new_n9998 , n5579 , n26054 );
nor  g07650 ( new_n9999 , new_n8753 , n23430 );
xnor g07651 ( new_n10000 , n19081 , n23430 );
nor  g07652 ( new_n10001 , new_n8771 , n10411 );
xnor g07653 ( new_n10002 , n8309 , n10411 );
not  g07654 ( new_n10003 , n16971 );
nor  g07655 ( new_n10004 , new_n10003 , n19144 );
nor  g07656 ( new_n10005 , n16971 , new_n8759 );
nor  g07657 ( new_n10006 , new_n2756 , n12593 );
not  g07658 ( new_n10007 , n12593 );
nor  g07659 ( new_n10008 , n11503 , new_n10007 );
nor  g07660 ( new_n10009_1 , n13714 , new_n2828 );
not  g07661 ( new_n10010_1 , new_n10009_1 );
nor  g07662 ( new_n10011 , new_n10008 , new_n10010_1 );
nor  g07663 ( new_n10012 , new_n10006 , new_n10011 );
nor  g07664 ( new_n10013 , new_n10005 , new_n10012 );
nor  g07665 ( new_n10014 , new_n10004 , new_n10013 );
and  g07666 ( new_n10015 , new_n10002 , new_n10014 );
or   g07667 ( new_n10016 , new_n10001 , new_n10015 );
and  g07668 ( new_n10017_1 , new_n10000 , new_n10016 );
or   g07669 ( new_n10018_1 , new_n9999 , new_n10017_1 );
and  g07670 ( new_n10019_1 , new_n9998 , new_n10018_1 );
or   g07671 ( new_n10020 , new_n9997 , new_n10019_1 );
and  g07672 ( new_n10021_1 , new_n9996 , new_n10020 );
or   g07673 ( new_n10022 , new_n9995 , new_n10021_1 );
and  g07674 ( new_n10023 , new_n9994 , new_n10022 );
or   g07675 ( new_n10024 , new_n9993 , new_n10023 );
and  g07676 ( new_n10025 , new_n9991 , new_n10024 );
or   g07677 ( new_n10026 , new_n9990 , new_n10025 );
and  g07678 ( new_n10027 , new_n9989 , new_n10026 );
nor  g07679 ( new_n10028 , new_n9988 , new_n10027 );
nor  g07680 ( new_n10029 , n11220 , n12650 );
not  g07681 ( new_n10030 , n11220 );
xnor g07682 ( new_n10031 , new_n10030 , n12650 );
nor  g07683 ( new_n10032 , n10201 , n22379 );
xnor g07684 ( new_n10033 , new_n5560 , n22379 );
nor  g07685 ( new_n10034 , n1662 , n10593 );
xnor g07686 ( new_n10035 , new_n2850 , n10593 );
nor  g07687 ( new_n10036 , n12875 , n18290 );
and  g07688 ( new_n10037 , new_n9226 , new_n9247 );
or   g07689 ( new_n10038 , new_n10036 , new_n10037 );
and  g07690 ( new_n10039 , new_n10035 , new_n10038 );
or   g07691 ( new_n10040 , new_n10034 , new_n10039 );
and  g07692 ( new_n10041 , new_n10033 , new_n10040 );
or   g07693 ( new_n10042 , new_n10032 , new_n10041 );
and  g07694 ( new_n10043 , new_n10031 , new_n10042 );
nor  g07695 ( new_n10044 , new_n10029 , new_n10043 );
not  g07696 ( new_n10045 , new_n10044 );
nor  g07697 ( new_n10046 , n2944 , n22270 );
or   g07698 ( new_n10047 , new_n2676 , new_n2717 );
and  g07699 ( new_n10048 , new_n2675 , new_n10047 );
nor  g07700 ( new_n10049 , new_n10046 , new_n10048 );
not  g07701 ( new_n10050 , new_n10049 );
xnor g07702 ( new_n10051 , new_n10045 , new_n10050 );
not  g07703 ( new_n10052 , new_n2719 );
nor  g07704 ( new_n10053_1 , new_n10032 , new_n10041 );
xnor g07705 ( new_n10054 , new_n10031 , new_n10053_1 );
nor  g07706 ( new_n10055_1 , new_n10052 , new_n10054 );
nor  g07707 ( new_n10056 , new_n10034 , new_n10039 );
xnor g07708 ( new_n10057_1 , new_n10033 , new_n10056 );
not  g07709 ( new_n10058 , new_n10057_1 );
nor  g07710 ( new_n10059 , new_n2723 , new_n10058 );
xnor g07711 ( new_n10060 , new_n2725 , new_n10057_1 );
nor  g07712 ( new_n10061 , new_n10036 , new_n10037 );
xnor g07713 ( new_n10062 , new_n10035 , new_n10061 );
not  g07714 ( new_n10063 , new_n10062 );
nor  g07715 ( new_n10064 , new_n2729 , new_n10063 );
xnor g07716 ( new_n10065 , new_n9615 , new_n10062 );
nor  g07717 ( new_n10066 , new_n2733 , new_n9249 );
nor  g07718 ( new_n10067 , new_n2738 , new_n9251_1 );
xnor g07719 ( new_n10068 , new_n2740 , new_n9251_1 );
nor  g07720 ( new_n10069 , new_n2771 , new_n9255 );
nor  g07721 ( new_n10070 , new_n2748 , new_n9261_1 );
xnor g07722 ( new_n10071 , new_n9626_1 , new_n9261_1 );
nor  g07723 ( new_n10072 , new_n2753 , new_n9266 );
xnor g07724 ( new_n10073 , new_n9629 , new_n9266 );
nor  g07725 ( new_n10074 , new_n2759 , new_n9274 );
nor  g07726 ( new_n10075 , new_n2761_1 , new_n9271 );
xnor g07727 ( new_n10076 , new_n2763 , new_n9274 );
and  g07728 ( new_n10077 , new_n10075 , new_n10076 );
or   g07729 ( new_n10078 , new_n10074 , new_n10077 );
and  g07730 ( new_n10079 , new_n10073 , new_n10078 );
or   g07731 ( new_n10080 , new_n10072 , new_n10079 );
and  g07732 ( new_n10081 , new_n10071 , new_n10080 );
nor  g07733 ( new_n10082 , new_n10070 , new_n10081 );
xnor g07734 ( new_n10083 , new_n2771 , new_n9256 );
and  g07735 ( new_n10084 , new_n10082 , new_n10083 );
nor  g07736 ( new_n10085 , new_n10069 , new_n10084 );
and  g07737 ( new_n10086 , new_n10068 , new_n10085 );
nor  g07738 ( new_n10087 , new_n10067 , new_n10086 );
xnor g07739 ( new_n10088 , new_n2733 , new_n9249 );
nor  g07740 ( new_n10089 , new_n10087 , new_n10088 );
nor  g07741 ( new_n10090 , new_n10066 , new_n10089 );
nor  g07742 ( new_n10091 , new_n10065 , new_n10090 );
nor  g07743 ( new_n10092 , new_n10064 , new_n10091 );
nor  g07744 ( new_n10093 , new_n10060 , new_n10092 );
nor  g07745 ( new_n10094 , new_n10059 , new_n10093 );
not  g07746 ( new_n10095 , new_n10054 );
xnor g07747 ( new_n10096_1 , new_n10052 , new_n10095 );
and  g07748 ( new_n10097 , new_n10094 , new_n10096_1 );
or   g07749 ( new_n10098 , new_n10055_1 , new_n10097 );
xor  g07750 ( new_n10099 , new_n10051 , new_n10098 );
xnor g07751 ( new_n10100 , new_n10028 , new_n10099 );
xor  g07752 ( new_n10101_1 , new_n9989 , new_n10026 );
xor  g07753 ( new_n10102 , new_n10094 , new_n10096_1 );
nor  g07754 ( new_n10103 , new_n10101_1 , new_n10102 );
xnor g07755 ( new_n10104 , new_n10101_1 , new_n10102 );
xor  g07756 ( new_n10105 , new_n9991 , new_n10024 );
xnor g07757 ( new_n10106 , new_n10060 , new_n10092 );
nor  g07758 ( new_n10107 , new_n10105 , new_n10106 );
xnor g07759 ( new_n10108 , new_n10105 , new_n10106 );
xor  g07760 ( new_n10109 , new_n9994 , new_n10022 );
xnor g07761 ( new_n10110 , new_n10065 , new_n10090 );
nor  g07762 ( new_n10111_1 , new_n10109 , new_n10110 );
xnor g07763 ( new_n10112 , new_n10109 , new_n10110 );
xor  g07764 ( new_n10113 , new_n9996 , new_n10020 );
xnor g07765 ( new_n10114 , new_n10087 , new_n10088 );
nor  g07766 ( new_n10115 , new_n10113 , new_n10114 );
xnor g07767 ( new_n10116 , new_n10113 , new_n10114 );
xor  g07768 ( new_n10117_1 , new_n9998 , new_n10018_1 );
xnor g07769 ( new_n10118 , new_n10068 , new_n10085 );
nor  g07770 ( new_n10119 , new_n10117_1 , new_n10118 );
xor  g07771 ( new_n10120 , new_n10000 , new_n10016 );
xor  g07772 ( new_n10121 , new_n10082 , new_n10083 );
nor  g07773 ( new_n10122 , new_n10120 , new_n10121 );
xnor g07774 ( new_n10123 , new_n10120 , new_n10121 );
xor  g07775 ( new_n10124 , new_n10071 , new_n10080 );
xnor g07776 ( new_n10125_1 , new_n10002 , new_n10014 );
and  g07777 ( new_n10126 , new_n10124 , new_n10125_1 );
nor  g07778 ( new_n10127 , new_n10074 , new_n10077 );
xnor g07779 ( new_n10128 , new_n10073 , new_n10127 );
xnor g07780 ( new_n10129 , n16971 , n19144 );
xnor g07781 ( new_n10130 , new_n10012 , new_n10129 );
and  g07782 ( new_n10131 , new_n10128 , new_n10130 );
not  g07783 ( new_n10132 , new_n10128 );
xnor g07784 ( new_n10133 , new_n10132 , new_n10130 );
xnor g07785 ( new_n10134 , new_n2761_1 , new_n9272 );
xnor g07786 ( new_n10135 , n13714 , n18151 );
nor  g07787 ( new_n10136 , new_n10134 , new_n10135 );
xnor g07788 ( new_n10137 , n11503 , n12593 );
xnor g07789 ( new_n10138 , new_n10010_1 , new_n10137 );
not  g07790 ( new_n10139 , new_n10138 );
and  g07791 ( new_n10140 , new_n10136 , new_n10139 );
xnor g07792 ( new_n10141 , new_n10075 , new_n10076 );
not  g07793 ( new_n10142 , new_n10141 );
xnor g07794 ( new_n10143 , new_n10136 , new_n10139 );
nor  g07795 ( new_n10144 , new_n10142 , new_n10143 );
nor  g07796 ( new_n10145 , new_n10140 , new_n10144 );
and  g07797 ( new_n10146 , new_n10133 , new_n10145 );
nor  g07798 ( new_n10147 , new_n10131 , new_n10146 );
xnor g07799 ( new_n10148 , new_n10124 , new_n10125_1 );
nor  g07800 ( new_n10149 , new_n10147 , new_n10148 );
nor  g07801 ( new_n10150 , new_n10126 , new_n10149 );
nor  g07802 ( new_n10151 , new_n10123 , new_n10150 );
nor  g07803 ( new_n10152 , new_n10122 , new_n10151 );
xnor g07804 ( new_n10153 , new_n10117_1 , new_n10118 );
nor  g07805 ( new_n10154 , new_n10152 , new_n10153 );
nor  g07806 ( new_n10155 , new_n10119 , new_n10154 );
nor  g07807 ( new_n10156 , new_n10116 , new_n10155 );
nor  g07808 ( new_n10157 , new_n10115 , new_n10156 );
nor  g07809 ( new_n10158_1 , new_n10112 , new_n10157 );
nor  g07810 ( new_n10159 , new_n10111_1 , new_n10158_1 );
nor  g07811 ( new_n10160 , new_n10108 , new_n10159 );
nor  g07812 ( new_n10161 , new_n10107 , new_n10160 );
nor  g07813 ( new_n10162 , new_n10104 , new_n10161 );
nor  g07814 ( new_n10163 , new_n10103 , new_n10162 );
xnor g07815 ( n1332 , new_n10100 , new_n10163 );
not  g07816 ( new_n10165_1 , new_n5542 );
nor  g07817 ( new_n10166 , n14692 , new_n5544 );
not  g07818 ( new_n10167 , new_n5544 );
xnor g07819 ( new_n10168 , n14692 , new_n10167 );
nor  g07820 ( new_n10169 , n4100 , new_n5619 );
not  g07821 ( new_n10170 , n4100 );
xnor g07822 ( new_n10171 , new_n10170 , new_n5620 );
nor  g07823 ( new_n10172 , n21957 , new_n5625 );
not  g07824 ( new_n10173 , n21957 );
xnor g07825 ( new_n10174 , new_n10173 , new_n5626 );
nor  g07826 ( new_n10175 , n15761 , new_n5631 );
not  g07827 ( new_n10176 , n15761 );
xnor g07828 ( new_n10177 , new_n10176 , new_n5632 );
nor  g07829 ( new_n10178 , n11201 , new_n5637 );
not  g07830 ( new_n10179 , n11201 );
xnor g07831 ( new_n10180 , new_n10179 , new_n5638 );
nor  g07832 ( new_n10181 , n18690 , new_n5643_1 );
not  g07833 ( new_n10182 , n18690 );
xnor g07834 ( new_n10183 , new_n10182 , new_n5644 );
nor  g07835 ( new_n10184 , n12153 , new_n5648 );
xnor g07836 ( new_n10185 , n12153 , new_n5649 );
not  g07837 ( new_n10186 , n13044 );
nor  g07838 ( new_n10187 , new_n10186 , new_n5655 );
nand g07839 ( new_n10188 , new_n10186 , new_n5655 );
nor  g07840 ( new_n10189 , n18745 , new_n5666 );
and  g07841 ( new_n10190 , new_n5806 , new_n5808 );
nor  g07842 ( new_n10191 , new_n10189 , new_n10190 );
and  g07843 ( new_n10192 , new_n10188 , new_n10191 );
nor  g07844 ( new_n10193 , new_n10187 , new_n10192 );
and  g07845 ( new_n10194 , new_n10185 , new_n10193 );
nor  g07846 ( new_n10195 , new_n10184 , new_n10194 );
nor  g07847 ( new_n10196 , new_n10183 , new_n10195 );
nor  g07848 ( new_n10197 , new_n10181 , new_n10196 );
nor  g07849 ( new_n10198 , new_n10180 , new_n10197 );
nor  g07850 ( new_n10199 , new_n10178 , new_n10198 );
nor  g07851 ( new_n10200 , new_n10177 , new_n10199 );
nor  g07852 ( new_n10201_1 , new_n10175 , new_n10200 );
nor  g07853 ( new_n10202 , new_n10174 , new_n10201_1 );
nor  g07854 ( new_n10203 , new_n10172 , new_n10202 );
nor  g07855 ( new_n10204 , new_n10171 , new_n10203 );
or   g07856 ( new_n10205 , new_n10169 , new_n10204 );
and  g07857 ( new_n10206 , new_n10168 , new_n10205 );
nor  g07858 ( new_n10207 , new_n10166 , new_n10206 );
not  g07859 ( new_n10208 , new_n10207 );
nor  g07860 ( new_n10209 , new_n10165_1 , new_n10208 );
not  g07861 ( new_n10210 , new_n10209 );
not  g07862 ( new_n10211 , new_n5817 );
nor  g07863 ( new_n10212 , n11302 , new_n10211 );
not  g07864 ( new_n10213 , new_n10212 );
nor  g07865 ( new_n10214 , n10405 , new_n10213 );
not  g07866 ( new_n10215 , new_n10214 );
nor  g07867 ( new_n10216 , n7693 , new_n10215 );
not  g07868 ( new_n10217 , new_n10216 );
nor  g07869 ( new_n10218 , n20151 , new_n10217 );
not  g07870 ( new_n10219 , new_n10218 );
nor  g07871 ( new_n10220 , n8964 , new_n10219 );
not  g07872 ( new_n10221 , new_n10220 );
nor  g07873 ( new_n10222 , n27037 , new_n10221 );
and  g07874 ( new_n10223 , new_n6215 , new_n10222 );
and  g07875 ( new_n10224 , new_n6198 , new_n10223 );
nor  g07876 ( new_n10225 , n7657 , n25926 );
not  g07877 ( new_n10226 , new_n10225 );
nor  g07878 ( new_n10227 , n5330 , new_n10226 );
not  g07879 ( new_n10228 , new_n10227 );
nor  g07880 ( new_n10229 , n5451 , new_n10228 );
not  g07881 ( new_n10230 , new_n10229 );
nor  g07882 ( new_n10231 , n18926 , new_n10230 );
not  g07883 ( new_n10232 , new_n10231 );
nor  g07884 ( new_n10233 , n13677 , new_n10232 );
not  g07885 ( new_n10234 , new_n10233 );
nor  g07886 ( new_n10235 , n23039 , new_n10234 );
not  g07887 ( new_n10236_1 , new_n10235 );
nor  g07888 ( new_n10237 , n7692 , new_n10236_1 );
not  g07889 ( new_n10238 , new_n10237 );
nor  g07890 ( new_n10239_1 , n25629 , new_n10238 );
and  g07891 ( new_n10240 , new_n6320 , new_n10239_1 );
xnor g07892 ( new_n10241 , n15766 , new_n10239_1 );
nor  g07893 ( new_n10242 , n23895 , new_n10241 );
xnor g07894 ( new_n10243 , n25629 , new_n10237 );
nor  g07895 ( new_n10244_1 , n17351 , new_n10243 );
xnor g07896 ( new_n10245 , new_n5456 , new_n10243 );
xnor g07897 ( new_n10246 , n7692 , new_n10235 );
nor  g07898 ( new_n10247 , n11736 , new_n10246 );
xnor g07899 ( new_n10248 , new_n5459 , new_n10246 );
xnor g07900 ( new_n10249 , n23039 , new_n10233 );
nor  g07901 ( new_n10250_1 , n23200 , new_n10249 );
xnor g07902 ( new_n10251 , new_n5462 , new_n10249 );
xnor g07903 ( new_n10252 , n13677 , new_n10231 );
nor  g07904 ( new_n10253 , n17959 , new_n10252 );
xnor g07905 ( new_n10254 , n18926 , new_n10229 );
nor  g07906 ( new_n10255 , n7566 , new_n10254 );
xnor g07907 ( new_n10256 , new_n5468 , new_n10254 );
xnor g07908 ( new_n10257 , n5451 , new_n10227 );
and  g07909 ( new_n10258 , n7731 , new_n10257 );
nor  g07910 ( new_n10259 , n7731 , new_n10257 );
xnor g07911 ( new_n10260 , n5330 , new_n10225 );
and  g07912 ( new_n10261_1 , n12341 , new_n10260 );
xnor g07913 ( new_n10262_1 , new_n5475 , new_n10260 );
nor  g07914 ( new_n10263 , new_n5478 , new_n5811 );
and  g07915 ( new_n10264 , new_n5810 , new_n5812 );
or   g07916 ( new_n10265 , new_n10263 , new_n10264 );
and  g07917 ( new_n10266 , new_n10262_1 , new_n10265 );
nor  g07918 ( new_n10267 , new_n10261_1 , new_n10266 );
nor  g07919 ( new_n10268 , new_n10259 , new_n10267 );
nor  g07920 ( new_n10269 , new_n10258 , new_n10268 );
and  g07921 ( new_n10270 , new_n10256 , new_n10269 );
or   g07922 ( new_n10271 , new_n10255 , new_n10270 );
xnor g07923 ( new_n10272 , new_n5465 , new_n10252 );
and  g07924 ( new_n10273 , new_n10271 , new_n10272 );
or   g07925 ( new_n10274 , new_n10253 , new_n10273 );
and  g07926 ( new_n10275_1 , new_n10251 , new_n10274 );
or   g07927 ( new_n10276 , new_n10250_1 , new_n10275_1 );
and  g07928 ( new_n10277 , new_n10248 , new_n10276 );
or   g07929 ( new_n10278 , new_n10247 , new_n10277 );
and  g07930 ( new_n10279 , new_n10245 , new_n10278 );
nor  g07931 ( new_n10280 , new_n10244_1 , new_n10279 );
not  g07932 ( new_n10281 , new_n10241 );
nor  g07933 ( new_n10282 , new_n5453 , new_n10281 );
nor  g07934 ( new_n10283 , new_n10280 , new_n10282 );
nor  g07935 ( new_n10284 , new_n10242 , new_n10283 );
nor  g07936 ( new_n10285 , new_n10240 , new_n10284 );
nor  g07937 ( new_n10286 , new_n10224 , new_n10285 );
xnor g07938 ( new_n10287_1 , n8614 , new_n10223 );
not  g07939 ( new_n10288 , new_n10287_1 );
xnor g07940 ( new_n10289 , n23895 , new_n10281 );
xnor g07941 ( new_n10290 , new_n10280 , new_n10289 );
nor  g07942 ( new_n10291 , new_n10288 , new_n10290 );
xnor g07943 ( new_n10292 , n15182 , new_n10222 );
nor  g07944 ( new_n10293 , new_n10247 , new_n10277 );
xnor g07945 ( new_n10294 , new_n10245 , new_n10293 );
not  g07946 ( new_n10295_1 , new_n10294 );
nor  g07947 ( new_n10296 , new_n10292 , new_n10295_1 );
xnor g07948 ( new_n10297 , new_n10292 , new_n10294 );
xnor g07949 ( new_n10298 , n27037 , new_n10220 );
xor  g07950 ( new_n10299 , new_n10248 , new_n10276 );
not  g07951 ( new_n10300 , new_n10299 );
nor  g07952 ( new_n10301 , new_n10298 , new_n10300 );
xnor g07953 ( new_n10302 , new_n10298 , new_n10300 );
xnor g07954 ( new_n10303 , n8964 , new_n10218 );
xor  g07955 ( new_n10304 , new_n10251 , new_n10274 );
not  g07956 ( new_n10305 , new_n10304 );
nor  g07957 ( new_n10306 , new_n10303 , new_n10305 );
xnor g07958 ( new_n10307 , new_n10303 , new_n10304 );
xnor g07959 ( new_n10308 , n20151 , new_n10216 );
xor  g07960 ( new_n10309 , new_n10271 , new_n10272 );
not  g07961 ( new_n10310 , new_n10309 );
nor  g07962 ( new_n10311 , new_n10308 , new_n10310 );
xnor g07963 ( new_n10312 , new_n10308 , new_n10310 );
xnor g07964 ( new_n10313 , n7693 , new_n10214 );
xnor g07965 ( new_n10314 , new_n10256 , new_n10269 );
nor  g07966 ( new_n10315 , new_n10313 , new_n10314 );
xor  g07967 ( new_n10316 , new_n10313 , new_n10314 );
xnor g07968 ( new_n10317 , n10405 , new_n10212 );
xnor g07969 ( new_n10318 , new_n5471 , new_n10257 );
xnor g07970 ( new_n10319 , new_n10267 , new_n10318 );
nor  g07971 ( new_n10320 , new_n10317 , new_n10319 );
xnor g07972 ( new_n10321_1 , new_n10317 , new_n10319 );
xor  g07973 ( new_n10322 , new_n10262_1 , new_n10265 );
xnor g07974 ( new_n10323 , n11302 , new_n5817 );
nor  g07975 ( new_n10324 , new_n10322 , new_n10323 );
xnor g07976 ( new_n10325 , new_n10322 , new_n10323 );
and  g07977 ( new_n10326_1 , new_n5813 , new_n5821 );
nor  g07978 ( new_n10327_1 , new_n5820 , new_n10326_1 );
nor  g07979 ( new_n10328 , new_n10325 , new_n10327_1 );
nor  g07980 ( new_n10329 , new_n10324 , new_n10328 );
nor  g07981 ( new_n10330_1 , new_n10321_1 , new_n10329 );
or   g07982 ( new_n10331 , new_n10320 , new_n10330_1 );
and  g07983 ( new_n10332 , new_n10316 , new_n10331 );
nor  g07984 ( new_n10333 , new_n10315 , new_n10332 );
nor  g07985 ( new_n10334 , new_n10312 , new_n10333 );
or   g07986 ( new_n10335 , new_n10311 , new_n10334 );
and  g07987 ( new_n10336 , new_n10307 , new_n10335 );
nor  g07988 ( new_n10337 , new_n10306 , new_n10336 );
nor  g07989 ( new_n10338 , new_n10302 , new_n10337 );
or   g07990 ( new_n10339 , new_n10301 , new_n10338 );
and  g07991 ( new_n10340_1 , new_n10297 , new_n10339 );
nor  g07992 ( new_n10341 , new_n10296 , new_n10340_1 );
not  g07993 ( new_n10342 , new_n10290 );
xnor g07994 ( new_n10343 , new_n10288 , new_n10342 );
and  g07995 ( new_n10344 , new_n10341 , new_n10343 );
nor  g07996 ( new_n10345_1 , new_n10291 , new_n10344 );
and  g07997 ( new_n10346 , new_n10286 , new_n10345_1 );
xnor g07998 ( new_n10347 , new_n10210 , new_n10346 );
xnor g07999 ( new_n10348 , new_n5542 , new_n10208 );
xnor g08000 ( new_n10349 , new_n10224 , new_n10285 );
xnor g08001 ( new_n10350 , new_n10345_1 , new_n10349 );
nor  g08002 ( new_n10351 , new_n10348 , new_n10350 );
not  g08003 ( new_n10352 , new_n10348 );
xnor g08004 ( new_n10353 , new_n10352 , new_n10350 );
xor  g08005 ( new_n10354 , new_n10168 , new_n10205 );
xnor g08006 ( new_n10355 , new_n10341 , new_n10343 );
nor  g08007 ( new_n10356_1 , new_n10354 , new_n10355 );
xor  g08008 ( new_n10357 , new_n10354 , new_n10355 );
xnor g08009 ( new_n10358 , new_n10297 , new_n10339 );
xnor g08010 ( new_n10359 , new_n10171 , new_n10203 );
and  g08011 ( new_n10360 , new_n10358 , new_n10359 );
xnor g08012 ( new_n10361 , new_n10302 , new_n10337 );
xnor g08013 ( new_n10362 , new_n10174 , new_n10201_1 );
nor  g08014 ( new_n10363 , new_n10361 , new_n10362 );
xnor g08015 ( new_n10364 , new_n10361 , new_n10362 );
not  g08016 ( new_n10365 , new_n10364 );
xnor g08017 ( new_n10366 , new_n10307 , new_n10335 );
xnor g08018 ( new_n10367 , new_n10177 , new_n10199 );
and  g08019 ( new_n10368 , new_n10366 , new_n10367 );
xnor g08020 ( new_n10369 , new_n10312 , new_n10333 );
xnor g08021 ( new_n10370 , new_n10180 , new_n10197 );
nor  g08022 ( new_n10371 , new_n10369 , new_n10370 );
xnor g08023 ( new_n10372_1 , new_n10369 , new_n10370 );
not  g08024 ( new_n10373 , new_n10372_1 );
xnor g08025 ( new_n10374 , new_n10316 , new_n10331 );
xnor g08026 ( new_n10375 , new_n10183 , new_n10195 );
and  g08027 ( new_n10376 , new_n10374 , new_n10375 );
xor  g08028 ( new_n10377 , new_n10374 , new_n10375 );
xnor g08029 ( new_n10378 , new_n10321_1 , new_n10329 );
xnor g08030 ( new_n10379 , new_n10185 , new_n10193 );
nor  g08031 ( new_n10380 , new_n10378 , new_n10379 );
xnor g08032 ( new_n10381 , new_n10378 , new_n10379 );
xnor g08033 ( new_n10382 , new_n10325 , new_n10327_1 );
xnor g08034 ( new_n10383 , new_n10186 , new_n5655 );
xnor g08035 ( new_n10384 , new_n10191 , new_n10383 );
nor  g08036 ( new_n10385_1 , new_n10382 , new_n10384 );
and  g08037 ( new_n10386 , new_n5809 , new_n5822_1 );
nor  g08038 ( new_n10387_1 , new_n5804 , new_n5823 );
nor  g08039 ( new_n10388_1 , new_n10386 , new_n10387_1 );
xnor g08040 ( new_n10389 , new_n10382 , new_n10384 );
nor  g08041 ( new_n10390_1 , new_n10388_1 , new_n10389 );
nor  g08042 ( new_n10391 , new_n10385_1 , new_n10390_1 );
nor  g08043 ( new_n10392 , new_n10381 , new_n10391 );
nor  g08044 ( new_n10393 , new_n10380 , new_n10392 );
and  g08045 ( new_n10394 , new_n10377 , new_n10393 );
nor  g08046 ( new_n10395 , new_n10376 , new_n10394 );
and  g08047 ( new_n10396 , new_n10373 , new_n10395 );
nor  g08048 ( new_n10397 , new_n10371 , new_n10396 );
xor  g08049 ( new_n10398 , new_n10366 , new_n10367 );
and  g08050 ( new_n10399 , new_n10397 , new_n10398 );
nor  g08051 ( new_n10400 , new_n10368 , new_n10399 );
and  g08052 ( new_n10401 , new_n10365 , new_n10400 );
nor  g08053 ( new_n10402 , new_n10363 , new_n10401 );
xor  g08054 ( new_n10403 , new_n10358 , new_n10359 );
and  g08055 ( new_n10404_1 , new_n10402 , new_n10403 );
or   g08056 ( new_n10405_1 , new_n10360 , new_n10404_1 );
and  g08057 ( new_n10406 , new_n10357 , new_n10405_1 );
nor  g08058 ( new_n10407 , new_n10356_1 , new_n10406 );
and  g08059 ( new_n10408 , new_n10353 , new_n10407 );
nor  g08060 ( new_n10409_1 , new_n10351 , new_n10408 );
not  g08061 ( new_n10410 , new_n10409_1 );
xnor g08062 ( n1357 , new_n10347 , new_n10410 );
xnor g08063 ( new_n10412 , n25240 , new_n7971 );
nor  g08064 ( new_n10413 , n10125 , new_n7976 );
not  g08065 ( new_n10414 , n10125 );
xnor g08066 ( new_n10415 , new_n10414 , new_n7976 );
nor  g08067 ( new_n10416 , n8067 , new_n7981 );
xnor g08068 ( new_n10417 , n8067 , new_n7981 );
nor  g08069 ( new_n10418 , n20923 , new_n7986 );
xnor g08070 ( new_n10419 , n20923 , new_n7986 );
nor  g08071 ( new_n10420_1 , n18157 , new_n7991 );
or   g08072 ( new_n10421 , new_n8434 , new_n8441 );
and  g08073 ( new_n10422 , new_n8433 , new_n10421 );
nor  g08074 ( new_n10423 , new_n10420_1 , new_n10422 );
nor  g08075 ( new_n10424 , new_n10419 , new_n10423 );
nor  g08076 ( new_n10425 , new_n10418 , new_n10424 );
nor  g08077 ( new_n10426 , new_n10417 , new_n10425 );
or   g08078 ( new_n10427 , new_n10416 , new_n10426 );
and  g08079 ( new_n10428 , new_n10415 , new_n10427 );
nor  g08080 ( new_n10429 , new_n10413 , new_n10428 );
xnor g08081 ( new_n10430 , new_n10412 , new_n10429 );
not  g08082 ( new_n10431 , n5077 );
xnor g08083 ( new_n10432_1 , n1099 , n6381 );
nor  g08084 ( new_n10433 , n2113 , n14345 );
not  g08085 ( new_n10434 , n2113 );
xnor g08086 ( new_n10435 , new_n10434 , n14345 );
nor  g08087 ( new_n10436 , n11356 , n21134 );
xnor g08088 ( new_n10437 , new_n9088 , n21134 );
nor  g08089 ( new_n10438 , new_n9091 , new_n4165_1 );
or   g08090 ( new_n10439 , n3164 , n6369 );
nor  g08091 ( new_n10440 , n10611 , n25797 );
or   g08092 ( new_n10441 , new_n6592 , new_n6601 );
and  g08093 ( new_n10442 , new_n6591 , new_n10441 );
nor  g08094 ( new_n10443 , new_n10440 , new_n10442 );
and  g08095 ( new_n10444 , new_n10439 , new_n10443 );
nor  g08096 ( new_n10445 , new_n10438 , new_n10444 );
and  g08097 ( new_n10446 , new_n10437 , new_n10445 );
or   g08098 ( new_n10447 , new_n10436 , new_n10446 );
and  g08099 ( new_n10448 , new_n10435 , new_n10447 );
nor  g08100 ( new_n10449 , new_n10433 , new_n10448 );
xnor g08101 ( new_n10450 , new_n10432_1 , new_n10449 );
xnor g08102 ( new_n10451 , new_n10431 , new_n10450 );
not  g08103 ( new_n10452 , n15546 );
nor  g08104 ( new_n10453 , new_n10436 , new_n10446 );
xnor g08105 ( new_n10454 , new_n10435 , new_n10453 );
nor  g08106 ( new_n10455 , new_n10452 , new_n10454 );
not  g08107 ( new_n10456 , new_n10454 );
xnor g08108 ( new_n10457 , new_n10452 , new_n10456 );
xnor g08109 ( new_n10458 , new_n10437 , new_n10445 );
nor  g08110 ( new_n10459 , n26452 , new_n10458 );
not  g08111 ( new_n10460 , n19905 );
xnor g08112 ( new_n10461 , new_n9091 , n6369 );
xnor g08113 ( new_n10462 , new_n10443 , new_n10461 );
nor  g08114 ( new_n10463 , new_n10460 , new_n10462 );
not  g08115 ( new_n10464 , new_n10462 );
xnor g08116 ( new_n10465 , new_n10460 , new_n10464 );
nor  g08117 ( new_n10466 , new_n8469 , new_n6603 );
and  g08118 ( new_n10467 , new_n8470 , new_n8473 );
or   g08119 ( new_n10468 , new_n10466 , new_n10467 );
and  g08120 ( new_n10469 , new_n10465 , new_n10468 );
nor  g08121 ( new_n10470 , new_n10463 , new_n10469 );
not  g08122 ( new_n10471 , new_n10458 );
xnor g08123 ( new_n10472 , n26452 , new_n10471 );
and  g08124 ( new_n10473 , new_n10470 , new_n10472 );
nor  g08125 ( new_n10474 , new_n10459 , new_n10473 );
and  g08126 ( new_n10475 , new_n10457 , new_n10474 );
nor  g08127 ( new_n10476 , new_n10455 , new_n10475 );
xor  g08128 ( new_n10477 , new_n10451 , new_n10476 );
xnor g08129 ( new_n10478 , new_n10430 , new_n10477 );
xor  g08130 ( new_n10479 , new_n10415 , new_n10427 );
xnor g08131 ( new_n10480 , new_n10457 , new_n10474 );
not  g08132 ( new_n10481 , new_n10480 );
and  g08133 ( new_n10482 , new_n10479 , new_n10481 );
xnor g08134 ( new_n10483 , new_n10479 , new_n10481 );
xnor g08135 ( new_n10484_1 , new_n10417 , new_n10425 );
xor  g08136 ( new_n10485 , new_n10470 , new_n10472 );
nor  g08137 ( new_n10486 , new_n10484_1 , new_n10485 );
xnor g08138 ( new_n10487 , new_n10484_1 , new_n10485 );
xnor g08139 ( new_n10488 , new_n10419 , new_n10423 );
nor  g08140 ( new_n10489_1 , new_n10466 , new_n10467 );
xnor g08141 ( new_n10490 , new_n10465 , new_n10489_1 );
not  g08142 ( new_n10491 , new_n10490 );
nor  g08143 ( new_n10492 , new_n10488 , new_n10491 );
xnor g08144 ( new_n10493 , new_n10488 , new_n10490 );
not  g08145 ( new_n10494 , new_n8467 );
nor  g08146 ( new_n10495 , new_n8443 , new_n10494 );
and  g08147 ( new_n10496 , new_n8468 , new_n8474 );
nor  g08148 ( new_n10497 , new_n10495 , new_n10496 );
and  g08149 ( new_n10498 , new_n10493 , new_n10497 );
nor  g08150 ( new_n10499 , new_n10492 , new_n10498 );
nor  g08151 ( new_n10500 , new_n10487 , new_n10499 );
nor  g08152 ( new_n10501 , new_n10486 , new_n10500 );
nor  g08153 ( new_n10502 , new_n10483 , new_n10501 );
nor  g08154 ( new_n10503 , new_n10482 , new_n10502 );
xnor g08155 ( n1371 , new_n10478 , new_n10503 );
xnor g08156 ( new_n10505 , n15241 , n17250 );
not  g08157 ( new_n10506 , n23160 );
nor  g08158 ( new_n10507 , n7678 , new_n10506 );
and  g08159 ( new_n10508 , new_n4377 , n16524 );
xnor g08160 ( new_n10509 , n3785 , n16524 );
nor  g08161 ( new_n10510 , n11056 , new_n4382 );
nor  g08162 ( new_n10511 , new_n4384 , n15271 );
xnor g08163 ( new_n10512 , n5822 , n15271 );
nor  g08164 ( new_n10513 , n25877 , new_n6644 );
and  g08165 ( new_n10514_1 , new_n5777 , new_n5778 );
or   g08166 ( new_n10515 , new_n10513 , new_n10514_1 );
and  g08167 ( new_n10516 , new_n10512 , new_n10515 );
or   g08168 ( new_n10517 , new_n10511 , new_n10516 );
xnor g08169 ( new_n10518 , n11056 , n20250 );
and  g08170 ( new_n10519 , new_n10517 , new_n10518 );
nor  g08171 ( new_n10520 , new_n10510 , new_n10519 );
and  g08172 ( new_n10521 , new_n10509 , new_n10520 );
or   g08173 ( new_n10522 , new_n10508 , new_n10521 );
xnor g08174 ( new_n10523 , n7678 , n23160 );
and  g08175 ( new_n10524 , new_n10522 , new_n10523 );
or   g08176 ( new_n10525_1 , new_n10507 , new_n10524 );
xor  g08177 ( new_n10526 , new_n10505 , new_n10525_1 );
xnor g08178 ( new_n10527 , new_n2425 , new_n9617 );
not  g08179 ( new_n10528 , new_n10527 );
nor  g08180 ( new_n10529 , n26660 , new_n9620 );
xnor g08181 ( new_n10530 , new_n7618 , new_n9620 );
and  g08182 ( new_n10531 , n3018 , new_n9623 );
nor  g08183 ( new_n10532 , n3018 , new_n9623 );
and  g08184 ( new_n10533 , n3480 , new_n9413 );
not  g08185 ( new_n10534 , new_n9414 );
nor  g08186 ( new_n10535 , new_n10534 , new_n9422 );
nor  g08187 ( new_n10536 , new_n10533 , new_n10535 );
nor  g08188 ( new_n10537 , new_n10532 , new_n10536 );
nor  g08189 ( new_n10538 , new_n10531 , new_n10537 );
and  g08190 ( new_n10539 , new_n10530 , new_n10538 );
nor  g08191 ( new_n10540_1 , new_n10529 , new_n10539 );
xnor g08192 ( new_n10541 , new_n10528 , new_n10540_1 );
xnor g08193 ( new_n10542 , new_n10526 , new_n10541 );
xnor g08194 ( new_n10543 , new_n10530 , new_n10538 );
xor  g08195 ( new_n10544 , new_n10522 , new_n10523 );
and  g08196 ( new_n10545 , new_n10543 , new_n10544 );
not  g08197 ( new_n10546 , new_n10543 );
xnor g08198 ( new_n10547 , new_n10546 , new_n10544 );
xnor g08199 ( new_n10548 , new_n10509 , new_n10520 );
not  g08200 ( new_n10549 , new_n10548 );
not  g08201 ( new_n10550 , n3018 );
xnor g08202 ( new_n10551 , new_n10550 , new_n9623 );
xnor g08203 ( new_n10552 , new_n10536 , new_n10551 );
nor  g08204 ( new_n10553 , new_n10549 , new_n10552 );
not  g08205 ( new_n10554 , new_n10552 );
xnor g08206 ( new_n10555 , new_n10548 , new_n10554 );
nor  g08207 ( new_n10556 , new_n10511 , new_n10516 );
xnor g08208 ( new_n10557 , new_n10556 , new_n10518 );
not  g08209 ( new_n10558 , new_n10557 );
nor  g08210 ( new_n10559 , new_n9423_1 , new_n10558 );
xnor g08211 ( new_n10560 , new_n9423_1 , new_n10557 );
xor  g08212 ( new_n10561_1 , new_n10512 , new_n10515 );
nor  g08213 ( new_n10562 , new_n9425 , new_n10561_1 );
xnor g08214 ( new_n10563 , new_n9425 , new_n10561_1 );
and  g08215 ( new_n10564_1 , new_n5776_1 , new_n5779 );
nor  g08216 ( new_n10565 , new_n5780 , new_n5788 );
nor  g08217 ( new_n10566 , new_n10564_1 , new_n10565 );
nor  g08218 ( new_n10567 , new_n10563 , new_n10566 );
nor  g08219 ( new_n10568 , new_n10562 , new_n10567 );
and  g08220 ( new_n10569 , new_n10560 , new_n10568 );
nor  g08221 ( new_n10570 , new_n10559 , new_n10569 );
nor  g08222 ( new_n10571 , new_n10555 , new_n10570 );
nor  g08223 ( new_n10572 , new_n10553 , new_n10571 );
and  g08224 ( new_n10573 , new_n10547 , new_n10572 );
nor  g08225 ( new_n10574 , new_n10545 , new_n10573 );
xnor g08226 ( new_n10575 , new_n10542 , new_n10574 );
not  g08227 ( new_n10576 , new_n10575 );
xnor g08228 ( new_n10577_1 , new_n5632 , new_n10576 );
xor  g08229 ( new_n10578 , new_n10547 , new_n10572 );
nor  g08230 ( new_n10579 , new_n5637 , new_n10578 );
xnor g08231 ( new_n10580 , new_n5637 , new_n10578 );
not  g08232 ( new_n10581 , new_n10580 );
xor  g08233 ( new_n10582 , new_n10555 , new_n10570 );
nor  g08234 ( new_n10583 , new_n5644 , new_n10582 );
xnor g08235 ( new_n10584 , new_n10560 , new_n10568 );
nor  g08236 ( new_n10585 , new_n5648 , new_n10584 );
xnor g08237 ( new_n10586 , new_n5648 , new_n10584 );
not  g08238 ( new_n10587 , new_n10586 );
xor  g08239 ( new_n10588_1 , new_n10563 , new_n10566 );
not  g08240 ( new_n10589 , new_n10588_1 );
nor  g08241 ( new_n10590 , new_n5655 , new_n10589 );
and  g08242 ( new_n10591 , new_n5666 , new_n5773 );
not  g08243 ( new_n10592 , new_n5790 );
nor  g08244 ( new_n10593_1 , new_n5774 , new_n10592 );
nor  g08245 ( new_n10594 , new_n10591 , new_n10593_1 );
xnor g08246 ( new_n10595_1 , new_n5655 , new_n10589 );
nor  g08247 ( new_n10596 , new_n10594 , new_n10595_1 );
nor  g08248 ( new_n10597 , new_n10590 , new_n10596 );
and  g08249 ( new_n10598 , new_n10587 , new_n10597 );
nor  g08250 ( new_n10599 , new_n10585 , new_n10598 );
not  g08251 ( new_n10600 , new_n10582 );
xnor g08252 ( new_n10601 , new_n5644 , new_n10600 );
and  g08253 ( new_n10602 , new_n10599 , new_n10601 );
nor  g08254 ( new_n10603 , new_n10583 , new_n10602 );
and  g08255 ( new_n10604 , new_n10581 , new_n10603 );
nor  g08256 ( new_n10605 , new_n10579 , new_n10604 );
xor  g08257 ( n1385 , new_n10577_1 , new_n10605 );
xnor g08258 ( new_n10607 , n24732 , n26808 );
not  g08259 ( new_n10608 , new_n10607 );
nor  g08260 ( new_n10609 , new_n4183 , new_n9155 );
xnor g08261 ( new_n10610 , n6631 , n7339 );
xnor g08262 ( new_n10611_1 , new_n10609 , new_n10610 );
nor  g08263 ( new_n10612 , new_n10608 , new_n10611_1 );
not  g08264 ( new_n10613 , new_n10612 );
not  g08265 ( new_n10614_1 , n1667 );
xnor g08266 ( new_n10615 , new_n10614_1 , n14684 );
nor  g08267 ( new_n10616 , n6631 , n7339 );
nor  g08268 ( new_n10617_1 , new_n10609 , new_n10610 );
nor  g08269 ( new_n10618 , new_n10616 , new_n10617_1 );
xnor g08270 ( new_n10619 , new_n10615 , new_n10618 );
not  g08271 ( new_n10620 , new_n10619 );
nor  g08272 ( new_n10621 , new_n10613 , new_n10620 );
not  g08273 ( new_n10622 , new_n10621 );
not  g08274 ( new_n10623 , n2680 );
xnor g08275 ( new_n10624 , new_n10623 , n17035 );
nor  g08276 ( new_n10625 , n1667 , n14684 );
or   g08277 ( new_n10626 , new_n10616 , new_n10617_1 );
and  g08278 ( new_n10627 , new_n10615 , new_n10626 );
nor  g08279 ( new_n10628_1 , new_n10625 , new_n10627 );
xnor g08280 ( new_n10629 , new_n10624 , new_n10628_1 );
not  g08281 ( new_n10630 , new_n10629 );
nor  g08282 ( new_n10631 , new_n10622 , new_n10630 );
not  g08283 ( new_n10632 , new_n10631 );
not  g08284 ( new_n10633 , n2547 );
xnor g08285 ( new_n10634 , new_n10633 , n19905 );
nor  g08286 ( new_n10635 , n2680 , n17035 );
or   g08287 ( new_n10636 , new_n10625 , new_n10627 );
and  g08288 ( new_n10637 , new_n10624 , new_n10636 );
nor  g08289 ( new_n10638 , new_n10635 , new_n10637 );
xnor g08290 ( new_n10639 , new_n10634 , new_n10638 );
not  g08291 ( new_n10640 , new_n10639 );
nor  g08292 ( new_n10641 , new_n10632 , new_n10640 );
not  g08293 ( new_n10642 , new_n10641 );
not  g08294 ( new_n10643 , n2999 );
xnor g08295 ( new_n10644 , new_n10643 , n26452 );
nor  g08296 ( new_n10645 , n2547 , n19905 );
not  g08297 ( new_n10646 , new_n10634 );
nor  g08298 ( new_n10647_1 , new_n10646 , new_n10638 );
nor  g08299 ( new_n10648 , new_n10645 , new_n10647_1 );
xnor g08300 ( new_n10649 , new_n10644 , new_n10648 );
not  g08301 ( new_n10650_1 , new_n10649 );
nor  g08302 ( new_n10651 , new_n10642 , new_n10650_1 );
not  g08303 ( new_n10652 , new_n10651 );
xnor g08304 ( new_n10653_1 , n14702 , new_n10452 );
nor  g08305 ( new_n10654 , n2999 , n26452 );
not  g08306 ( new_n10655 , new_n10644 );
nor  g08307 ( new_n10656 , new_n10655 , new_n10648 );
nor  g08308 ( new_n10657 , new_n10654 , new_n10656 );
xnor g08309 ( new_n10658 , new_n10653_1 , new_n10657 );
not  g08310 ( new_n10659 , new_n10658 );
nor  g08311 ( new_n10660 , new_n10652 , new_n10659 );
not  g08312 ( new_n10661 , new_n10660 );
xnor g08313 ( new_n10662 , new_n10431 , n13914 );
nor  g08314 ( new_n10663 , n14702 , n15546 );
not  g08315 ( new_n10664 , new_n10653_1 );
nor  g08316 ( new_n10665 , new_n10664 , new_n10657 );
nor  g08317 ( new_n10666 , new_n10663 , new_n10665 );
xnor g08318 ( new_n10667 , new_n10662 , new_n10666 );
not  g08319 ( new_n10668 , new_n10667 );
nor  g08320 ( new_n10669 , new_n10661 , new_n10668 );
not  g08321 ( new_n10670 , new_n10669 );
xnor g08322 ( new_n10671 , new_n9062 , n18035 );
nor  g08323 ( new_n10672 , n5077 , n13914 );
not  g08324 ( new_n10673 , new_n10662 );
nor  g08325 ( new_n10674 , new_n10673 , new_n10666 );
nor  g08326 ( new_n10675 , new_n10672 , new_n10674 );
xnor g08327 ( new_n10676 , new_n10671 , new_n10675 );
not  g08328 ( new_n10677 , new_n10676 );
nor  g08329 ( new_n10678 , new_n10670 , new_n10677 );
not  g08330 ( new_n10679 , n4306 );
xnor g08331 ( new_n10680 , new_n10679 , n8827 );
nor  g08332 ( new_n10681 , n3279 , n18035 );
not  g08333 ( new_n10682 , new_n10671 );
nor  g08334 ( new_n10683 , new_n10682 , new_n10675 );
nor  g08335 ( new_n10684 , new_n10681 , new_n10683 );
xnor g08336 ( new_n10685 , new_n10680 , new_n10684 );
xor  g08337 ( new_n10686 , new_n10678 , new_n10685 );
xnor g08338 ( new_n10687 , new_n7959_1 , new_n10686 );
xnor g08339 ( new_n10688 , new_n10669 , new_n10677 );
nor  g08340 ( new_n10689 , new_n7966 , new_n10688 );
xnor g08341 ( new_n10690 , new_n7964 , new_n10688 );
xnor g08342 ( new_n10691 , new_n10660 , new_n10668 );
nor  g08343 ( new_n10692_1 , new_n7971 , new_n10691 );
xnor g08344 ( new_n10693 , new_n7969 , new_n10691 );
xnor g08345 ( new_n10694_1 , new_n10651 , new_n10659 );
nor  g08346 ( new_n10695 , new_n7976 , new_n10694_1 );
xnor g08347 ( new_n10696 , new_n7974 , new_n10694_1 );
xnor g08348 ( new_n10697 , new_n10641 , new_n10650_1 );
nor  g08349 ( new_n10698 , new_n7981 , new_n10697 );
xnor g08350 ( new_n10699 , new_n7979 , new_n10697 );
xnor g08351 ( new_n10700 , new_n10631 , new_n10640 );
nor  g08352 ( new_n10701_1 , new_n7986 , new_n10700 );
xnor g08353 ( new_n10702 , new_n7984 , new_n10700 );
xnor g08354 ( new_n10703 , new_n10621 , new_n10630 );
nor  g08355 ( new_n10704 , new_n7991 , new_n10703 );
xnor g08356 ( new_n10705 , new_n7991 , new_n10703 );
xnor g08357 ( new_n10706 , new_n10612 , new_n10620 );
nor  g08358 ( new_n10707 , new_n7995 , new_n10706 );
xnor g08359 ( new_n10708 , new_n7995 , new_n10706 );
nor  g08360 ( new_n10709 , new_n2543 , new_n10607 );
nor  g08361 ( new_n10710_1 , new_n8003 , new_n10709 );
nor  g08362 ( new_n10711 , new_n10607 , new_n10610 );
or   g08363 ( new_n10712_1 , new_n10612 , new_n10711 );
and  g08364 ( new_n10713 , new_n7942 , new_n10709 );
nor  g08365 ( new_n10714 , new_n10710_1 , new_n10713 );
and  g08366 ( new_n10715 , new_n10712_1 , new_n10714 );
nor  g08367 ( new_n10716 , new_n10710_1 , new_n10715 );
nor  g08368 ( new_n10717 , new_n10708 , new_n10716 );
nor  g08369 ( new_n10718 , new_n10707 , new_n10717 );
nor  g08370 ( new_n10719 , new_n10705 , new_n10718 );
or   g08371 ( new_n10720 , new_n10704 , new_n10719 );
and  g08372 ( new_n10721 , new_n10702 , new_n10720 );
or   g08373 ( new_n10722 , new_n10701_1 , new_n10721 );
and  g08374 ( new_n10723 , new_n10699 , new_n10722 );
or   g08375 ( new_n10724 , new_n10698 , new_n10723 );
and  g08376 ( new_n10725 , new_n10696 , new_n10724 );
or   g08377 ( new_n10726 , new_n10695 , new_n10725 );
and  g08378 ( new_n10727 , new_n10693 , new_n10726 );
or   g08379 ( new_n10728 , new_n10692_1 , new_n10727 );
and  g08380 ( new_n10729 , new_n10690 , new_n10728 );
or   g08381 ( new_n10730 , new_n10689 , new_n10729 );
xor  g08382 ( new_n10731 , new_n10687 , new_n10730 );
xnor g08383 ( new_n10732 , new_n9119 , new_n10731 );
xor  g08384 ( new_n10733 , new_n10690 , new_n10728 );
and  g08385 ( new_n10734 , new_n9123 , new_n10733 );
xnor g08386 ( new_n10735 , new_n9123 , new_n10733 );
xor  g08387 ( new_n10736 , new_n10693 , new_n10726 );
and  g08388 ( new_n10737 , new_n9127 , new_n10736 );
xnor g08389 ( new_n10738 , new_n9127 , new_n10736 );
xor  g08390 ( new_n10739_1 , new_n10696 , new_n10724 );
and  g08391 ( new_n10740 , new_n9131 , new_n10739_1 );
xnor g08392 ( new_n10741 , new_n9131 , new_n10739_1 );
xor  g08393 ( new_n10742 , new_n10699 , new_n10722 );
and  g08394 ( new_n10743 , new_n9135 , new_n10742 );
xnor g08395 ( new_n10744 , new_n9135 , new_n10742 );
xor  g08396 ( new_n10745 , new_n10702 , new_n10720 );
and  g08397 ( new_n10746 , new_n9138 , new_n10745 );
xnor g08398 ( new_n10747 , new_n9138 , new_n10745 );
xnor g08399 ( new_n10748 , new_n10705 , new_n10718 );
nor  g08400 ( new_n10749 , new_n9142 , new_n10748 );
xnor g08401 ( new_n10750 , new_n10708 , new_n10716 );
nor  g08402 ( new_n10751 , new_n9147 , new_n10750 );
xnor g08403 ( new_n10752 , new_n9147 , new_n10750 );
xnor g08404 ( new_n10753 , new_n2543 , new_n10608 );
nor  g08405 ( new_n10754 , new_n9156 , new_n10753 );
and  g08406 ( new_n10755 , new_n9158 , new_n10754 );
xnor g08407 ( new_n10756_1 , new_n9153 , new_n10754 );
xnor g08408 ( new_n10757 , new_n10712_1 , new_n10714 );
not  g08409 ( new_n10758 , new_n10757 );
and  g08410 ( new_n10759 , new_n10756_1 , new_n10758 );
nor  g08411 ( new_n10760 , new_n10755 , new_n10759 );
nor  g08412 ( new_n10761 , new_n10752 , new_n10760 );
nor  g08413 ( new_n10762 , new_n10751 , new_n10761 );
xnor g08414 ( new_n10763_1 , new_n9142 , new_n10748 );
nor  g08415 ( new_n10764 , new_n10762 , new_n10763_1 );
nor  g08416 ( new_n10765 , new_n10749 , new_n10764 );
nor  g08417 ( new_n10766 , new_n10747 , new_n10765 );
nor  g08418 ( new_n10767 , new_n10746 , new_n10766 );
nor  g08419 ( new_n10768 , new_n10744 , new_n10767 );
nor  g08420 ( new_n10769 , new_n10743 , new_n10768 );
nor  g08421 ( new_n10770 , new_n10741 , new_n10769 );
nor  g08422 ( new_n10771 , new_n10740 , new_n10770 );
nor  g08423 ( new_n10772 , new_n10738 , new_n10771 );
nor  g08424 ( new_n10773 , new_n10737 , new_n10772 );
nor  g08425 ( new_n10774 , new_n10735 , new_n10773 );
nor  g08426 ( new_n10775_1 , new_n10734 , new_n10774 );
xnor g08427 ( n1498 , new_n10732 , new_n10775_1 );
not  g08428 ( new_n10777 , new_n5956 );
xnor g08429 ( new_n10778 , n9090 , n20658 );
xnor g08430 ( new_n10779 , new_n10777 , new_n10778 );
xnor g08431 ( n1501 , new_n5004 , new_n10779 );
nor  g08432 ( new_n10781 , n11473 , n15506 );
not  g08433 ( new_n10782 , new_n10781 );
nor  g08434 ( new_n10783 , n5131 , new_n10782 );
not  g08435 ( new_n10784 , new_n10783 );
nor  g08436 ( new_n10785 , n21538 , new_n10784 );
not  g08437 ( new_n10786 , new_n10785 );
nor  g08438 ( new_n10787 , n25094 , new_n10786 );
not  g08439 ( new_n10788 , new_n10787 );
nor  g08440 ( new_n10789 , n1611 , new_n10788 );
xnor g08441 ( new_n10790 , n752 , new_n10789 );
xnor g08442 ( new_n10791 , new_n9660 , new_n10790 );
xnor g08443 ( new_n10792_1 , n1611 , new_n10787 );
nor  g08444 ( new_n10793 , new_n9662 , new_n10792_1 );
xnor g08445 ( new_n10794 , new_n9662 , new_n10792_1 );
xnor g08446 ( new_n10795 , n25094 , new_n10785 );
nor  g08447 ( new_n10796 , new_n9667 , new_n10795 );
xnor g08448 ( new_n10797 , new_n9667 , new_n10795 );
xnor g08449 ( new_n10798 , n21538 , new_n10783 );
and  g08450 ( new_n10799 , new_n9675 , new_n10798 );
xnor g08451 ( new_n10800 , n5131 , new_n10781 );
nor  g08452 ( new_n10801 , new_n9680 , new_n10800 );
xnor g08453 ( new_n10802 , new_n9680 , new_n10800 );
not  g08454 ( new_n10803 , n15506 );
nor  g08455 ( new_n10804 , new_n10803 , new_n9686 );
xnor g08456 ( new_n10805 , n11473 , n15506 );
not  g08457 ( new_n10806 , new_n10805 );
nor  g08458 ( new_n10807 , new_n10804 , new_n10806 );
not  g08459 ( new_n10808 , new_n9683 );
not  g08460 ( new_n10809 , n11473 );
and  g08461 ( new_n10810 , new_n10809 , new_n10804 );
nor  g08462 ( new_n10811 , new_n10807 , new_n10810 );
and  g08463 ( new_n10812 , new_n10808 , new_n10811 );
nor  g08464 ( new_n10813 , new_n10807 , new_n10812 );
nor  g08465 ( new_n10814 , new_n10802 , new_n10813 );
nor  g08466 ( new_n10815 , new_n10801 , new_n10814 );
xnor g08467 ( new_n10816 , new_n9673 , new_n10798 );
and  g08468 ( new_n10817_1 , new_n10815 , new_n10816 );
or   g08469 ( new_n10818 , new_n10799 , new_n10817_1 );
nor  g08470 ( new_n10819 , new_n10797 , new_n10818 );
nor  g08471 ( new_n10820 , new_n10796 , new_n10819 );
nor  g08472 ( new_n10821 , new_n10794 , new_n10820 );
nor  g08473 ( new_n10822 , new_n10793 , new_n10821 );
xor  g08474 ( new_n10823 , new_n10791 , new_n10822 );
not  g08475 ( new_n10824 , n20470 );
xnor g08476 ( new_n10825 , n3366 , new_n10824 );
and  g08477 ( new_n10826 , n21222 , n26565 );
or   g08478 ( new_n10827 , n21222 , n26565 );
nor  g08479 ( new_n10828 , n3959 , n9832 );
or   g08480 ( new_n10829 , new_n9478 , new_n9493_1 );
and  g08481 ( new_n10830 , new_n9477 , new_n10829 );
nor  g08482 ( new_n10831 , new_n10828 , new_n10830 );
and  g08483 ( new_n10832 , new_n10827 , new_n10831 );
nor  g08484 ( new_n10833 , new_n10826 , new_n10832 );
xor  g08485 ( new_n10834_1 , new_n10825 , new_n10833 );
xnor g08486 ( new_n10835 , new_n10823 , new_n10834_1 );
xor  g08487 ( new_n10836 , new_n10794 , new_n10820 );
not  g08488 ( new_n10837 , n21222 );
xnor g08489 ( new_n10838 , new_n10837 , n26565 );
xnor g08490 ( new_n10839 , new_n10831 , new_n10838 );
not  g08491 ( new_n10840 , new_n10839 );
and  g08492 ( new_n10841 , new_n10836 , new_n10840 );
xnor g08493 ( new_n10842 , new_n10836 , new_n10840 );
not  g08494 ( new_n10843 , new_n9495 );
xor  g08495 ( new_n10844 , new_n10797 , new_n10818 );
and  g08496 ( new_n10845 , new_n10843 , new_n10844 );
xnor g08497 ( new_n10846 , new_n10843 , new_n10844 );
xnor g08498 ( new_n10847 , new_n10815 , new_n10816 );
not  g08499 ( new_n10848 , new_n10847 );
nor  g08500 ( new_n10849 , new_n9546 , new_n10848 );
xnor g08501 ( new_n10850 , new_n9546 , new_n10848 );
xor  g08502 ( new_n10851_1 , new_n10802 , new_n10813 );
nor  g08503 ( new_n10852 , new_n9551 , new_n10851_1 );
xnor g08504 ( new_n10853 , new_n10808 , new_n10811 );
nor  g08505 ( new_n10854 , new_n9557_1 , new_n10853 );
xnor g08506 ( new_n10855 , n15506 , new_n9686 );
nor  g08507 ( new_n10856 , new_n7198 , new_n10855 );
xnor g08508 ( new_n10857 , new_n9560 , new_n10853 );
and  g08509 ( new_n10858 , new_n10856 , new_n10857 );
nor  g08510 ( new_n10859 , new_n10854 , new_n10858 );
xor  g08511 ( new_n10860 , new_n9551 , new_n10851_1 );
and  g08512 ( new_n10861 , new_n10859 , new_n10860 );
or   g08513 ( new_n10862 , new_n10852 , new_n10861 );
nor  g08514 ( new_n10863 , new_n10850 , new_n10862 );
nor  g08515 ( new_n10864 , new_n10849 , new_n10863 );
nor  g08516 ( new_n10865 , new_n10846 , new_n10864 );
nor  g08517 ( new_n10866 , new_n10845 , new_n10865 );
nor  g08518 ( new_n10867 , new_n10842 , new_n10866 );
nor  g08519 ( new_n10868 , new_n10841 , new_n10867 );
xnor g08520 ( n1518 , new_n10835 , new_n10868 );
not  g08521 ( new_n10870 , n17458 );
nor  g08522 ( new_n10871 , n14826 , new_n10870 );
xnor g08523 ( new_n10872 , n14826 , n17458 );
not  g08524 ( new_n10873 , n1222 );
nor  g08525 ( new_n10874_1 , new_n10873 , n23493 );
xnor g08526 ( new_n10875 , n1222 , n23493 );
not  g08527 ( new_n10876 , n25240 );
nor  g08528 ( new_n10877 , n10275 , new_n10876 );
xnor g08529 ( new_n10878 , n10275 , n25240 );
nor  g08530 ( new_n10879 , new_n10414 , n15146 );
xnor g08531 ( new_n10880 , n10125 , n15146 );
not  g08532 ( new_n10881 , n8067 );
nor  g08533 ( new_n10882 , new_n10881 , n11579 );
xnor g08534 ( new_n10883 , n8067 , n11579 );
not  g08535 ( new_n10884 , n20923 );
nor  g08536 ( new_n10885 , n21 , new_n10884 );
xnor g08537 ( new_n10886 , n21 , n20923 );
nor  g08538 ( new_n10887 , n1682 , new_n8432_1 );
xnor g08539 ( new_n10888 , n1682 , n18157 );
nor  g08540 ( new_n10889 , new_n9835 , n12161 );
nor  g08541 ( new_n10890 , n7963 , new_n7217 );
nor  g08542 ( new_n10891 , n5026 , new_n7941 );
nor  g08543 ( new_n10892 , new_n7220 , n10017 );
nor  g08544 ( new_n10893 , new_n7939 , n8581 );
not  g08545 ( new_n10894 , new_n10893 );
nor  g08546 ( new_n10895 , new_n10892 , new_n10894 );
nor  g08547 ( new_n10896 , new_n10891 , new_n10895 );
nor  g08548 ( new_n10897 , new_n10890 , new_n10896 );
nor  g08549 ( new_n10898 , new_n10889 , new_n10897 );
and  g08550 ( new_n10899 , new_n10888 , new_n10898 );
or   g08551 ( new_n10900 , new_n10887 , new_n10899 );
and  g08552 ( new_n10901 , new_n10886 , new_n10900 );
or   g08553 ( new_n10902 , new_n10885 , new_n10901 );
and  g08554 ( new_n10903 , new_n10883 , new_n10902 );
or   g08555 ( new_n10904 , new_n10882 , new_n10903 );
and  g08556 ( new_n10905 , new_n10880 , new_n10904 );
or   g08557 ( new_n10906 , new_n10879 , new_n10905 );
and  g08558 ( new_n10907 , new_n10878 , new_n10906 );
or   g08559 ( new_n10908 , new_n10877 , new_n10907 );
and  g08560 ( new_n10909 , new_n10875 , new_n10908 );
or   g08561 ( new_n10910 , new_n10874_1 , new_n10909 );
and  g08562 ( new_n10911 , new_n10872 , new_n10910 );
nor  g08563 ( new_n10912 , new_n10871 , new_n10911 );
not  g08564 ( new_n10913 , new_n4200 );
nor  g08565 ( new_n10914 , n3468 , new_n10913 );
not  g08566 ( new_n10915 , new_n10914 );
nor  g08567 ( new_n10916 , n12821 , new_n10915 );
not  g08568 ( new_n10917 , new_n10916 );
nor  g08569 ( new_n10918 , n22492 , new_n10917 );
not  g08570 ( new_n10919 , new_n10918 );
nor  g08571 ( new_n10920 , n7330 , new_n10919 );
not  g08572 ( new_n10921 , new_n10920 );
nor  g08573 ( new_n10922 , n767 , new_n10921 );
xnor g08574 ( new_n10923 , n2944 , new_n10922 );
and  g08575 ( new_n10924_1 , n19282 , new_n10923 );
and  g08576 ( new_n10925 , new_n2674 , new_n10922 );
xnor g08577 ( new_n10926 , n767 , new_n10920 );
nor  g08578 ( new_n10927 , n12657 , new_n10926 );
xnor g08579 ( new_n10928 , new_n2926 , new_n10926 );
xnor g08580 ( new_n10929 , n7330 , new_n10918 );
and  g08581 ( new_n10930 , n17077 , new_n10929 );
xnor g08582 ( new_n10931 , n17077 , new_n10929 );
xnor g08583 ( new_n10932 , n22492 , new_n10916 );
not  g08584 ( new_n10933 , new_n10932 );
nor  g08585 ( new_n10934 , new_n7251 , new_n10933 );
xnor g08586 ( new_n10935 , n26510 , new_n10933 );
xnor g08587 ( new_n10936 , n12821 , new_n10914 );
not  g08588 ( new_n10937 , new_n10936 );
nor  g08589 ( new_n10938 , new_n3815 , new_n10937 );
nor  g08590 ( new_n10939 , n23068 , new_n10936 );
and  g08591 ( new_n10940 , n19514 , new_n4201 );
or   g08592 ( new_n10941 , new_n4205_1 , new_n4219 );
and  g08593 ( new_n10942 , new_n4203 , new_n10941 );
nor  g08594 ( new_n10943_1 , new_n10940 , new_n10942 );
nor  g08595 ( new_n10944 , new_n10939 , new_n10943_1 );
or   g08596 ( new_n10945 , new_n10938 , new_n10944 );
and  g08597 ( new_n10946 , new_n10935 , new_n10945 );
nor  g08598 ( new_n10947 , new_n10934 , new_n10946 );
nor  g08599 ( new_n10948 , new_n10931 , new_n10947 );
nor  g08600 ( new_n10949 , new_n10930 , new_n10948 );
and  g08601 ( new_n10950 , new_n10928 , new_n10949 );
nor  g08602 ( new_n10951 , new_n10927 , new_n10950 );
or   g08603 ( new_n10952 , n19282 , new_n10923 );
and  g08604 ( new_n10953 , new_n10951 , new_n10952 );
or   g08605 ( new_n10954 , new_n10925 , new_n10953 );
nor  g08606 ( new_n10955 , new_n10924_1 , new_n10954 );
nor  g08607 ( new_n10956 , new_n10912 , new_n10955 );
xor  g08608 ( new_n10957 , new_n10872 , new_n10910 );
not  g08609 ( new_n10958 , n19282 );
xnor g08610 ( new_n10959 , new_n10958 , new_n10923 );
xnor g08611 ( new_n10960 , new_n10951 , new_n10959 );
not  g08612 ( new_n10961_1 , new_n10960 );
nor  g08613 ( new_n10962 , new_n10957 , new_n10961_1 );
xnor g08614 ( new_n10963 , new_n10957 , new_n10961_1 );
xor  g08615 ( new_n10964 , new_n10875 , new_n10908 );
xnor g08616 ( new_n10965 , new_n10928 , new_n10949 );
nor  g08617 ( new_n10966 , new_n10964 , new_n10965 );
xnor g08618 ( new_n10967 , new_n10964 , new_n10965 );
xor  g08619 ( new_n10968 , new_n10878 , new_n10906 );
xnor g08620 ( new_n10969 , new_n10931 , new_n10947 );
not  g08621 ( new_n10970 , new_n10969 );
nor  g08622 ( new_n10971 , new_n10968 , new_n10970 );
xnor g08623 ( new_n10972 , new_n10968 , new_n10970 );
xor  g08624 ( new_n10973 , new_n10880 , new_n10904 );
xor  g08625 ( new_n10974 , new_n10935 , new_n10945 );
nor  g08626 ( new_n10975 , new_n10973 , new_n10974 );
xnor g08627 ( new_n10976 , new_n10973 , new_n10974 );
xor  g08628 ( new_n10977 , new_n10883 , new_n10902 );
xnor g08629 ( new_n10978 , n23068 , new_n10937 );
xnor g08630 ( new_n10979 , new_n10943_1 , new_n10978 );
nor  g08631 ( new_n10980 , new_n10977 , new_n10979 );
xnor g08632 ( new_n10981 , new_n10977 , new_n10979 );
xor  g08633 ( new_n10982 , new_n10886 , new_n10900 );
nor  g08634 ( new_n10983 , new_n4221_1 , new_n10982 );
xnor g08635 ( new_n10984 , new_n10888 , new_n10898 );
not  g08636 ( new_n10985 , new_n10984 );
nor  g08637 ( new_n10986 , new_n4254 , new_n10985 );
xnor g08638 ( new_n10987 , new_n4255 , new_n10984 );
xnor g08639 ( new_n10988 , n7963 , n12161 );
xnor g08640 ( new_n10989 , new_n10896 , new_n10988 );
and  g08641 ( new_n10990 , new_n4290 , new_n10989 );
xnor g08642 ( new_n10991 , new_n4290 , new_n10989 );
xnor g08643 ( new_n10992 , n3618 , n8581 );
nor  g08644 ( new_n10993 , new_n4268 , new_n10992 );
xnor g08645 ( new_n10994 , n5026 , n10017 );
xnor g08646 ( new_n10995 , new_n10894 , new_n10994 );
not  g08647 ( new_n10996 , new_n10995 );
nor  g08648 ( new_n10997 , new_n10993 , new_n10996 );
xnor g08649 ( new_n10998 , new_n10993 , new_n10995 );
and  g08650 ( new_n10999 , new_n4262 , new_n10998 );
nor  g08651 ( new_n11000 , new_n10997 , new_n10999 );
nor  g08652 ( new_n11001 , new_n10991 , new_n11000 );
nor  g08653 ( new_n11002 , new_n10990 , new_n11001 );
nor  g08654 ( new_n11003 , new_n10987 , new_n11002 );
nor  g08655 ( new_n11004 , new_n10986 , new_n11003 );
xnor g08656 ( new_n11005_1 , new_n4221_1 , new_n10982 );
nor  g08657 ( new_n11006 , new_n11004 , new_n11005_1 );
nor  g08658 ( new_n11007 , new_n10983 , new_n11006 );
nor  g08659 ( new_n11008 , new_n10981 , new_n11007 );
nor  g08660 ( new_n11009 , new_n10980 , new_n11008 );
nor  g08661 ( new_n11010 , new_n10976 , new_n11009 );
nor  g08662 ( new_n11011_1 , new_n10975 , new_n11010 );
nor  g08663 ( new_n11012 , new_n10972 , new_n11011_1 );
nor  g08664 ( new_n11013 , new_n10971 , new_n11012 );
nor  g08665 ( new_n11014 , new_n10967 , new_n11013 );
nor  g08666 ( new_n11015 , new_n10966 , new_n11014 );
nor  g08667 ( new_n11016 , new_n10963 , new_n11015 );
nor  g08668 ( new_n11017 , new_n10962 , new_n11016 );
not  g08669 ( new_n11018 , new_n10912 );
xnor g08670 ( new_n11019 , new_n11018 , new_n10955 );
and  g08671 ( new_n11020 , new_n11017 , new_n11019 );
nor  g08672 ( new_n11021 , new_n10956 , new_n11020 );
nor  g08673 ( new_n11022 , new_n7429 , n20040 );
or   g08674 ( new_n11023_1 , new_n8683 , new_n8716_1 );
and  g08675 ( new_n11024 , new_n8682 , new_n11023_1 );
nor  g08676 ( new_n11025_1 , new_n11022 , new_n11024 );
not  g08677 ( new_n11026 , new_n11025_1 );
xnor g08678 ( new_n11027 , new_n11021 , new_n11026 );
xor  g08679 ( new_n11028 , new_n11017 , new_n11019 );
nor  g08680 ( new_n11029 , new_n11025_1 , new_n11028 );
xnor g08681 ( new_n11030 , new_n10963 , new_n11015 );
nor  g08682 ( new_n11031 , new_n8718 , new_n11030 );
not  g08683 ( new_n11032 , new_n8718 );
not  g08684 ( new_n11033 , new_n11030 );
xnor g08685 ( new_n11034 , new_n11032 , new_n11033 );
xnor g08686 ( new_n11035 , new_n10967 , new_n11013 );
nor  g08687 ( new_n11036 , new_n8788 , new_n11035 );
not  g08688 ( new_n11037 , new_n11035 );
xnor g08689 ( new_n11038 , new_n8793 , new_n11037 );
xnor g08690 ( new_n11039 , new_n10972 , new_n11011_1 );
nor  g08691 ( new_n11040 , new_n8795 , new_n11039 );
xnor g08692 ( new_n11041 , new_n8795 , new_n11039 );
xnor g08693 ( new_n11042 , new_n10976 , new_n11009 );
nor  g08694 ( new_n11043 , new_n8801 , new_n11042 );
not  g08695 ( new_n11044_1 , new_n11042 );
xnor g08696 ( new_n11045 , new_n8802 , new_n11044_1 );
xnor g08697 ( new_n11046 , new_n10981 , new_n11007 );
nor  g08698 ( new_n11047 , new_n8807 , new_n11046 );
not  g08699 ( new_n11048 , new_n11046 );
xnor g08700 ( new_n11049 , new_n8807 , new_n11048 );
xnor g08701 ( new_n11050 , new_n11004 , new_n11005_1 );
not  g08702 ( new_n11051 , new_n11050 );
nor  g08703 ( new_n11052 , new_n8814 , new_n11051 );
xnor g08704 ( new_n11053 , new_n10987 , new_n11002 );
nor  g08705 ( new_n11054 , new_n8821_1 , new_n11053 );
not  g08706 ( new_n11055 , new_n11053 );
xnor g08707 ( new_n11056_1 , new_n8818 , new_n11055 );
not  g08708 ( new_n11057 , new_n8825 );
xnor g08709 ( new_n11058 , new_n10991 , new_n11000 );
nor  g08710 ( new_n11059 , new_n11057 , new_n11058 );
xnor g08711 ( new_n11060 , new_n4267 , new_n10992 );
not  g08712 ( new_n11061 , new_n11060 );
nor  g08713 ( new_n11062 , new_n8832 , new_n11061 );
and  g08714 ( new_n11063_1 , new_n8835 , new_n11062 );
xnor g08715 ( new_n11064 , new_n4270 , new_n10998 );
xnor g08716 ( new_n11065 , new_n8830 , new_n11062 );
not  g08717 ( new_n11066 , new_n11065 );
nor  g08718 ( new_n11067 , new_n11064 , new_n11066 );
nor  g08719 ( new_n11068 , new_n11063_1 , new_n11067 );
not  g08720 ( new_n11069 , new_n11058 );
xnor g08721 ( new_n11070 , new_n11057 , new_n11069 );
and  g08722 ( new_n11071 , new_n11068 , new_n11070 );
nor  g08723 ( new_n11072 , new_n11059 , new_n11071 );
nor  g08724 ( new_n11073 , new_n11056_1 , new_n11072 );
nor  g08725 ( new_n11074 , new_n11054 , new_n11073 );
xnor g08726 ( new_n11075 , new_n8813 , new_n11051 );
and  g08727 ( new_n11076 , new_n11074 , new_n11075 );
nor  g08728 ( new_n11077 , new_n11052 , new_n11076 );
and  g08729 ( new_n11078_1 , new_n11049 , new_n11077 );
nor  g08730 ( new_n11079 , new_n11047 , new_n11078_1 );
nor  g08731 ( new_n11080_1 , new_n11045 , new_n11079 );
nor  g08732 ( new_n11081 , new_n11043 , new_n11080_1 );
nor  g08733 ( new_n11082 , new_n11041 , new_n11081 );
nor  g08734 ( new_n11083 , new_n11040 , new_n11082 );
nor  g08735 ( new_n11084 , new_n11038 , new_n11083 );
nor  g08736 ( new_n11085 , new_n11036 , new_n11084 );
nor  g08737 ( new_n11086 , new_n11034 , new_n11085 );
nor  g08738 ( new_n11087 , new_n11031 , new_n11086 );
xnor g08739 ( new_n11088 , new_n11025_1 , new_n11028 );
nor  g08740 ( new_n11089 , new_n11087 , new_n11088 );
nor  g08741 ( new_n11090 , new_n11029 , new_n11089 );
xor  g08742 ( n1527 , new_n11027 , new_n11090 );
xnor g08743 ( new_n11092 , n23463 , n25345 );
nor  g08744 ( new_n11093 , n9655 , new_n3095 );
xnor g08745 ( new_n11094_1 , n9655 , n13074 );
nor  g08746 ( new_n11095 , new_n3099 , n13490 );
xnor g08747 ( new_n11096 , n10739 , n13490 );
nor  g08748 ( new_n11097 , new_n2350 , n22660 );
xnor g08749 ( new_n11098 , n21753 , n22660 );
nor  g08750 ( new_n11099 , n1777 , new_n2353 );
xnor g08751 ( new_n11100 , n1777 , n21832 );
nor  g08752 ( new_n11101_1 , n8745 , new_n2356 );
nor  g08753 ( new_n11102 , new_n2441 , n16223 );
and  g08754 ( new_n11103_1 , new_n9712 , new_n9717 );
nor  g08755 ( new_n11104 , new_n11102 , new_n11103_1 );
xnor g08756 ( new_n11105 , n8745 , n26913 );
and  g08757 ( new_n11106 , new_n11104 , new_n11105 );
or   g08758 ( new_n11107 , new_n11101_1 , new_n11106 );
and  g08759 ( new_n11108 , new_n11100 , new_n11107 );
or   g08760 ( new_n11109 , new_n11099 , new_n11108 );
and  g08761 ( new_n11110 , new_n11098 , new_n11109 );
or   g08762 ( new_n11111 , new_n11097 , new_n11110 );
and  g08763 ( new_n11112 , new_n11096 , new_n11111 );
or   g08764 ( new_n11113 , new_n11095 , new_n11112 );
and  g08765 ( new_n11114 , new_n11094_1 , new_n11113 );
or   g08766 ( new_n11115 , new_n11093 , new_n11114 );
xor  g08767 ( new_n11116 , new_n11092 , new_n11115 );
xnor g08768 ( new_n11117 , new_n7845 , new_n11116 );
xor  g08769 ( new_n11118 , new_n11094_1 , new_n11113 );
nor  g08770 ( new_n11119 , new_n7851 , new_n11118 );
xnor g08771 ( new_n11120_1 , new_n7851 , new_n11118 );
xor  g08772 ( new_n11121_1 , new_n11096 , new_n11111 );
nor  g08773 ( new_n11122 , new_n7858 , new_n11121_1 );
xnor g08774 ( new_n11123 , new_n7858 , new_n11121_1 );
xor  g08775 ( new_n11124 , new_n11098 , new_n11109 );
nor  g08776 ( new_n11125 , new_n7864 , new_n11124 );
xnor g08777 ( new_n11126 , new_n7864 , new_n11124 );
xor  g08778 ( new_n11127_1 , new_n11100 , new_n11107 );
nor  g08779 ( new_n11128 , new_n7871 , new_n11127_1 );
xnor g08780 ( new_n11129 , new_n7871 , new_n11127_1 );
xnor g08781 ( new_n11130 , new_n11104 , new_n11105 );
and  g08782 ( new_n11131 , new_n7879 , new_n11130 );
and  g08783 ( new_n11132_1 , new_n7882 , new_n9718 );
nor  g08784 ( new_n11133 , new_n9719 , new_n9727 );
nor  g08785 ( new_n11134_1 , new_n11132_1 , new_n11133 );
xnor g08786 ( new_n11135 , new_n7879 , new_n11130 );
nor  g08787 ( new_n11136 , new_n11134_1 , new_n11135 );
nor  g08788 ( new_n11137 , new_n11131 , new_n11136 );
nor  g08789 ( new_n11138_1 , new_n11129 , new_n11137 );
nor  g08790 ( new_n11139 , new_n11128 , new_n11138_1 );
nor  g08791 ( new_n11140 , new_n11126 , new_n11139 );
nor  g08792 ( new_n11141 , new_n11125 , new_n11140 );
nor  g08793 ( new_n11142 , new_n11123 , new_n11141 );
nor  g08794 ( new_n11143 , new_n11122 , new_n11142 );
nor  g08795 ( new_n11144 , new_n11120_1 , new_n11143 );
nor  g08796 ( new_n11145 , new_n11119 , new_n11144 );
xor  g08797 ( n1580 , new_n11117 , new_n11145 );
xnor g08798 ( new_n11147 , n12315 , n18962 );
nor  g08799 ( new_n11148 , new_n7401 , new_n11147 );
nor  g08800 ( new_n11149 , n12315 , new_n6771 );
xnor g08801 ( new_n11150 , n3952 , n10158 );
xnor g08802 ( new_n11151 , new_n11149 , new_n11150 );
xnor g08803 ( new_n11152 , new_n11148 , new_n11151 );
xnor g08804 ( n1586 , new_n7407 , new_n11152 );
xnor g08805 ( new_n11154 , n1483 , n19539 );
not  g08806 ( new_n11155 , n8194 );
nor  g08807 ( new_n11156 , new_n11155 , n24093 );
xnor g08808 ( new_n11157 , n8194 , n24093 );
not  g08809 ( new_n11158 , n23657 );
nor  g08810 ( new_n11159 , n23035 , new_n11158 );
xnor g08811 ( new_n11160 , n23035 , n23657 );
not  g08812 ( new_n11161 , n16911 );
nor  g08813 ( new_n11162 , n7773 , new_n11161 );
and  g08814 ( new_n11163 , new_n6432 , new_n6460 );
or   g08815 ( new_n11164 , new_n11162 , new_n11163 );
and  g08816 ( new_n11165 , new_n11160 , new_n11164 );
or   g08817 ( new_n11166 , new_n11159 , new_n11165 );
and  g08818 ( new_n11167 , new_n11157 , new_n11166 );
or   g08819 ( new_n11168 , new_n11156 , new_n11167 );
xor  g08820 ( new_n11169 , new_n11154 , new_n11168 );
xnor g08821 ( new_n11170 , n1314 , n25494 );
and  g08822 ( new_n11171 , n3306 , new_n3424 );
xnor g08823 ( new_n11172 , n3306 , n10117 );
nor  g08824 ( new_n11173 , n13460 , new_n8230 );
xnor g08825 ( new_n11174 , n13460 , n22335 );
nor  g08826 ( new_n11175 , n6104 , new_n8234 );
nor  g08827 ( new_n11176 , new_n8238 , n4119 );
and  g08828 ( new_n11177 , new_n4637 , new_n4659 );
or   g08829 ( new_n11178 , new_n11176 , new_n11177 );
xnor g08830 ( new_n11179 , n6104 , n24048 );
and  g08831 ( new_n11180 , new_n11178 , new_n11179 );
or   g08832 ( new_n11181 , new_n11175 , new_n11180 );
and  g08833 ( new_n11182_1 , new_n11174 , new_n11181 );
or   g08834 ( new_n11183 , new_n11173 , new_n11182_1 );
and  g08835 ( new_n11184_1 , new_n11172 , new_n11183 );
or   g08836 ( new_n11185 , new_n11171 , new_n11184_1 );
xor  g08837 ( new_n11186 , new_n11170 , new_n11185 );
xnor g08838 ( new_n11187 , n23717 , n25296 );
not  g08839 ( new_n11188 , n7788 );
nor  g08840 ( new_n11189 , new_n11188 , n20013 );
xnor g08841 ( new_n11190 , n7788 , n20013 );
not  g08842 ( new_n11191 , n5443 );
nor  g08843 ( new_n11192_1 , n1320 , new_n11191 );
xnor g08844 ( new_n11193 , n1320 , n5443 );
not  g08845 ( new_n11194 , n18584 );
nor  g08846 ( new_n11195 , new_n11194 , n19803 );
or   g08847 ( new_n11196 , new_n6427_1 , new_n6428 );
and  g08848 ( new_n11197 , new_n6425 , new_n11196 );
or   g08849 ( new_n11198 , new_n11195 , new_n11197 );
and  g08850 ( new_n11199 , new_n11193 , new_n11198 );
or   g08851 ( new_n11200 , new_n11192_1 , new_n11199 );
and  g08852 ( new_n11201_1 , new_n11190 , new_n11200 );
or   g08853 ( new_n11202 , new_n11189 , new_n11201_1 );
xor  g08854 ( new_n11203 , new_n11187 , new_n11202 );
xnor g08855 ( new_n11204 , new_n11186 , new_n11203 );
xor  g08856 ( new_n11205 , new_n11172 , new_n11183 );
xor  g08857 ( new_n11206 , new_n11190 , new_n11200 );
and  g08858 ( new_n11207 , new_n11205 , new_n11206 );
xor  g08859 ( new_n11208 , new_n11205 , new_n11206 );
xor  g08860 ( new_n11209 , new_n11174 , new_n11181 );
xor  g08861 ( new_n11210 , new_n11193 , new_n11198 );
nor  g08862 ( new_n11211 , new_n11209 , new_n11210 );
xnor g08863 ( new_n11212 , new_n11209 , new_n11210 );
not  g08864 ( new_n11213 , new_n11212 );
xor  g08865 ( new_n11214 , new_n11178 , new_n11179 );
and  g08866 ( new_n11215 , new_n6430 , new_n11214 );
xnor g08867 ( new_n11216 , new_n6430 , new_n11214 );
and  g08868 ( new_n11217 , new_n4660 , new_n4685 );
nor  g08869 ( new_n11218 , new_n4686 , new_n4722_1 );
nor  g08870 ( new_n11219 , new_n11217 , new_n11218 );
nor  g08871 ( new_n11220_1 , new_n11216 , new_n11219 );
nor  g08872 ( new_n11221 , new_n11215 , new_n11220_1 );
and  g08873 ( new_n11222 , new_n11213 , new_n11221 );
nor  g08874 ( new_n11223_1 , new_n11211 , new_n11222 );
and  g08875 ( new_n11224 , new_n11208 , new_n11223_1 );
nor  g08876 ( new_n11225 , new_n11207 , new_n11224 );
xnor g08877 ( new_n11226 , new_n11204 , new_n11225 );
xnor g08878 ( new_n11227 , new_n11169 , new_n11226 );
xor  g08879 ( new_n11228 , new_n11157 , new_n11166 );
xor  g08880 ( new_n11229 , new_n11208 , new_n11223_1 );
nor  g08881 ( new_n11230 , new_n11228 , new_n11229 );
xnor g08882 ( new_n11231 , new_n11228 , new_n11229 );
xor  g08883 ( new_n11232 , new_n11160 , new_n11164 );
xnor g08884 ( new_n11233 , new_n11213 , new_n11221 );
nor  g08885 ( new_n11234_1 , new_n11232 , new_n11233 );
xnor g08886 ( new_n11235 , new_n11232 , new_n11233 );
xnor g08887 ( new_n11236 , new_n11216 , new_n11219 );
not  g08888 ( new_n11237 , new_n11236 );
nor  g08889 ( new_n11238 , new_n6461 , new_n11237 );
xnor g08890 ( new_n11239 , new_n6461 , new_n11237 );
not  g08891 ( new_n11240 , new_n4723 );
nor  g08892 ( new_n11241 , new_n11240 , new_n6510 );
nor  g08893 ( new_n11242 , new_n4726 , new_n6520 );
xnor g08894 ( new_n11243 , new_n4726 , new_n6520 );
and  g08895 ( new_n11244 , new_n4730 , new_n6522 );
and  g08896 ( new_n11245_1 , new_n4734 , new_n6528 );
xnor g08897 ( new_n11246 , new_n4734 , new_n6528 );
nor  g08898 ( new_n11247 , new_n4740 , new_n6532 );
nor  g08899 ( new_n11248 , new_n6536 , new_n11247 );
xnor g08900 ( new_n11249 , new_n6535 , new_n11247 );
and  g08901 ( new_n11250 , new_n4745_1 , new_n11249 );
nor  g08902 ( new_n11251 , new_n11248 , new_n11250 );
nor  g08903 ( new_n11252 , new_n11246 , new_n11251 );
nor  g08904 ( new_n11253 , new_n11245_1 , new_n11252 );
xnor g08905 ( new_n11254 , new_n4730 , new_n6522 );
nor  g08906 ( new_n11255 , new_n11253 , new_n11254 );
nor  g08907 ( new_n11256 , new_n11244 , new_n11255 );
nor  g08908 ( new_n11257 , new_n11243 , new_n11256 );
nor  g08909 ( new_n11258 , new_n11242 , new_n11257 );
xnor g08910 ( new_n11259 , new_n11240 , new_n6510 );
nor  g08911 ( new_n11260 , new_n11258 , new_n11259 );
nor  g08912 ( new_n11261_1 , new_n11241 , new_n11260 );
nor  g08913 ( new_n11262 , new_n11239 , new_n11261_1 );
nor  g08914 ( new_n11263 , new_n11238 , new_n11262 );
nor  g08915 ( new_n11264 , new_n11235 , new_n11263 );
nor  g08916 ( new_n11265 , new_n11234_1 , new_n11264 );
nor  g08917 ( new_n11266_1 , new_n11231 , new_n11265 );
nor  g08918 ( new_n11267 , new_n11230 , new_n11266_1 );
xor  g08919 ( n1590 , new_n11227 , new_n11267 );
xnor g08920 ( n1602 , new_n7576 , new_n7590 );
xor  g08921 ( n1634 , new_n2790 , new_n2845 );
xnor g08922 ( n1636 , new_n11231 , new_n11265 );
nor  g08923 ( new_n11272 , n4514 , n10514 );
not  g08924 ( new_n11273_1 , n4514 );
xnor g08925 ( new_n11274 , new_n11273_1 , n10514 );
nor  g08926 ( new_n11275_1 , n3984 , n18649 );
not  g08927 ( new_n11276 , n18649 );
xnor g08928 ( new_n11277 , n3984 , new_n11276 );
and  g08929 ( new_n11278 , n6218 , n19652 );
or   g08930 ( new_n11279 , n6218 , n19652 );
nor  g08931 ( new_n11280 , n3366 , n20470 );
and  g08932 ( new_n11281 , new_n10825 , new_n10833 );
nor  g08933 ( new_n11282 , new_n11280 , new_n11281 );
and  g08934 ( new_n11283 , new_n11279 , new_n11282 );
nor  g08935 ( new_n11284 , new_n11278 , new_n11283 );
and  g08936 ( new_n11285 , new_n11277 , new_n11284 );
or   g08937 ( new_n11286 , new_n11275_1 , new_n11285 );
and  g08938 ( new_n11287 , new_n11274 , new_n11286 );
nor  g08939 ( new_n11288 , new_n11272 , new_n11287 );
not  g08940 ( new_n11289 , n20040 );
xnor g08941 ( new_n11290_1 , new_n7429 , n18880 );
not  g08942 ( new_n11291 , new_n11290_1 );
nor  g08943 ( new_n11292 , n23697 , n25475 );
nor  g08944 ( new_n11293 , new_n6746 , new_n6787 );
nor  g08945 ( new_n11294 , new_n11292 , new_n11293 );
xnor g08946 ( new_n11295 , new_n11291 , new_n11294 );
not  g08947 ( new_n11296 , new_n11295 );
nor  g08948 ( new_n11297 , new_n11289 , new_n11296 );
xnor g08949 ( new_n11298 , new_n11289 , new_n11296 );
nor  g08950 ( new_n11299 , new_n2558 , new_n6789 );
xnor g08951 ( new_n11300 , new_n2558 , new_n6789 );
nor  g08952 ( new_n11301 , n18345 , new_n6791_1 );
xnor g08953 ( new_n11302_1 , n18345 , new_n6791_1 );
nor  g08954 ( new_n11303 , n13190 , new_n6794_1 );
xnor g08955 ( new_n11304 , new_n2566 , new_n6794_1 );
not  g08956 ( new_n11305 , n3460 );
nor  g08957 ( new_n11306 , new_n11305 , new_n6798 );
nor  g08958 ( new_n11307 , new_n9502 , new_n6802_1 );
nor  g08959 ( new_n11308 , new_n9503 , new_n9516 );
nor  g08960 ( new_n11309 , new_n11307 , new_n11308 );
xnor g08961 ( new_n11310 , new_n11305 , new_n6798 );
nor  g08962 ( new_n11311 , new_n11309 , new_n11310 );
nor  g08963 ( new_n11312 , new_n11306 , new_n11311 );
and  g08964 ( new_n11313_1 , new_n11304 , new_n11312 );
nor  g08965 ( new_n11314 , new_n11303 , new_n11313_1 );
nor  g08966 ( new_n11315 , new_n11302_1 , new_n11314 );
or   g08967 ( new_n11316 , new_n11301 , new_n11315 );
nor  g08968 ( new_n11317 , new_n11300 , new_n11316 );
nor  g08969 ( new_n11318 , new_n11299 , new_n11317 );
nor  g08970 ( new_n11319 , new_n11298 , new_n11318 );
nor  g08971 ( new_n11320 , new_n11297 , new_n11319 );
nor  g08972 ( new_n11321 , n2978 , n18880 );
nor  g08973 ( new_n11322 , new_n11291 , new_n11294 );
nor  g08974 ( new_n11323 , new_n11321 , new_n11322 );
xnor g08975 ( new_n11324 , new_n11320 , new_n11323 );
not  g08976 ( new_n11325_1 , n7569 );
not  g08977 ( new_n11326_1 , n17037 );
not  g08978 ( new_n11327 , new_n9500 );
nor  g08979 ( new_n11328 , n19575 , new_n11327 );
not  g08980 ( new_n11329 , new_n11328 );
nor  g08981 ( new_n11330_1 , n26512 , new_n11329 );
not  g08982 ( new_n11331 , new_n11330_1 );
nor  g08983 ( new_n11332 , n26191 , new_n11331 );
not  g08984 ( new_n11333 , new_n11332 );
nor  g08985 ( new_n11334 , n5386 , new_n11333 );
and  g08986 ( new_n11335 , new_n11326_1 , new_n11334 );
and  g08987 ( new_n11336 , new_n11325_1 , new_n11335 );
xnor g08988 ( new_n11337 , new_n11324 , new_n11336 );
xnor g08989 ( new_n11338 , new_n11298 , new_n11318 );
not  g08990 ( new_n11339 , new_n11338 );
xnor g08991 ( new_n11340 , n7569 , new_n11335 );
nor  g08992 ( new_n11341 , new_n11339 , new_n11340 );
xnor g08993 ( new_n11342 , new_n11339 , new_n11340 );
nor  g08994 ( new_n11343 , new_n11301 , new_n11315 );
xnor g08995 ( new_n11344 , new_n11300 , new_n11343 );
xnor g08996 ( new_n11345 , n17037 , new_n11334 );
nor  g08997 ( new_n11346 , new_n11344 , new_n11345 );
xnor g08998 ( new_n11347_1 , new_n11344 , new_n11345 );
xnor g08999 ( new_n11348_1 , new_n11302_1 , new_n11314 );
xnor g09000 ( new_n11349 , n5386 , new_n11332 );
nor  g09001 ( new_n11350 , new_n11348_1 , new_n11349 );
xnor g09002 ( new_n11351 , new_n11348_1 , new_n11349 );
xnor g09003 ( new_n11352_1 , new_n11304 , new_n11312 );
xnor g09004 ( new_n11353 , n26191 , new_n11330_1 );
nor  g09005 ( new_n11354 , new_n11352_1 , new_n11353 );
xnor g09006 ( new_n11355 , n26512 , new_n11328 );
not  g09007 ( new_n11356_1 , new_n11355 );
xor  g09008 ( new_n11357 , new_n11309 , new_n11310 );
not  g09009 ( new_n11358 , new_n11357 );
nor  g09010 ( new_n11359 , new_n11356_1 , new_n11358 );
xnor g09011 ( new_n11360 , new_n11356_1 , new_n11358 );
nor  g09012 ( new_n11361 , new_n9501 , new_n9517 );
and  g09013 ( new_n11362 , new_n9519 , new_n9542 );
or   g09014 ( new_n11363 , new_n11361 , new_n11362 );
nor  g09015 ( new_n11364 , new_n11360 , new_n11363 );
nor  g09016 ( new_n11365 , new_n11359 , new_n11364 );
not  g09017 ( new_n11366 , new_n11352_1 );
xnor g09018 ( new_n11367 , new_n11366 , new_n11353 );
and  g09019 ( new_n11368 , new_n11365 , new_n11367 );
nor  g09020 ( new_n11369 , new_n11354 , new_n11368 );
nor  g09021 ( new_n11370 , new_n11351 , new_n11369 );
nor  g09022 ( new_n11371 , new_n11350 , new_n11370 );
nor  g09023 ( new_n11372 , new_n11347_1 , new_n11371 );
nor  g09024 ( new_n11373 , new_n11346 , new_n11372 );
nor  g09025 ( new_n11374 , new_n11342 , new_n11373 );
nor  g09026 ( new_n11375_1 , new_n11341 , new_n11374 );
xnor g09027 ( new_n11376 , new_n11337 , new_n11375_1 );
xnor g09028 ( new_n11377 , new_n11288 , new_n11376 );
xor  g09029 ( new_n11378 , new_n11342 , new_n11373 );
xor  g09030 ( new_n11379_1 , new_n11274 , new_n11286 );
not  g09031 ( new_n11380 , new_n11379_1 );
and  g09032 ( new_n11381 , new_n11378 , new_n11380 );
xnor g09033 ( new_n11382 , new_n11378 , new_n11380 );
xnor g09034 ( new_n11383 , new_n11347_1 , new_n11371 );
xnor g09035 ( new_n11384 , new_n11277 , new_n11284 );
not  g09036 ( new_n11385 , new_n11384 );
nor  g09037 ( new_n11386_1 , new_n11383 , new_n11385 );
xnor g09038 ( new_n11387 , new_n11383 , new_n11385 );
xor  g09039 ( new_n11388 , new_n11351 , new_n11369 );
not  g09040 ( new_n11389 , n6218 );
xnor g09041 ( new_n11390 , new_n11389 , n19652 );
xnor g09042 ( new_n11391_1 , new_n11282 , new_n11390 );
not  g09043 ( new_n11392 , new_n11391_1 );
and  g09044 ( new_n11393 , new_n11388 , new_n11392 );
xnor g09045 ( new_n11394 , new_n11388 , new_n11392 );
xnor g09046 ( new_n11395 , new_n11365 , new_n11367 );
nor  g09047 ( new_n11396 , new_n10834_1 , new_n11395 );
xnor g09048 ( new_n11397 , new_n10834_1 , new_n11395 );
xor  g09049 ( new_n11398_1 , new_n11360 , new_n11363 );
and  g09050 ( new_n11399 , new_n10839 , new_n11398_1 );
nor  g09051 ( new_n11400 , new_n10839 , new_n11398_1 );
nor  g09052 ( new_n11401 , new_n10843 , new_n9543 );
and  g09053 ( new_n11402 , new_n9544 , new_n9567 );
nor  g09054 ( new_n11403_1 , new_n11401 , new_n11402 );
nor  g09055 ( new_n11404 , new_n11400 , new_n11403_1 );
or   g09056 ( new_n11405 , new_n11399 , new_n11404 );
nor  g09057 ( new_n11406 , new_n11397 , new_n11405 );
nor  g09058 ( new_n11407 , new_n11396 , new_n11406 );
nor  g09059 ( new_n11408 , new_n11394 , new_n11407 );
nor  g09060 ( new_n11409 , new_n11393 , new_n11408 );
nor  g09061 ( new_n11410 , new_n11387 , new_n11409 );
nor  g09062 ( new_n11411 , new_n11386_1 , new_n11410 );
nor  g09063 ( new_n11412 , new_n11382 , new_n11411 );
nor  g09064 ( new_n11413 , new_n11381 , new_n11412 );
xnor g09065 ( n1684 , new_n11377 , new_n11413 );
xnor g09066 ( new_n11415 , n3984 , new_n6216 );
nor  g09067 ( new_n11416 , n19652 , new_n6218_1 );
xnor g09068 ( new_n11417 , n19652 , new_n6220 );
nor  g09069 ( new_n11418 , n3366 , new_n6223_1 );
xnor g09070 ( new_n11419_1 , n3366 , new_n6224 );
nor  g09071 ( new_n11420 , n26565 , new_n4012 );
xnor g09072 ( new_n11421 , n26565 , new_n4013 );
nor  g09073 ( new_n11422 , n3959 , new_n4016 );
xnor g09074 ( new_n11423 , n3959 , new_n4017 );
nor  g09075 ( new_n11424_1 , n11566 , new_n4019 );
xor  g09076 ( new_n11425 , n11566 , new_n4019 );
nor  g09077 ( new_n11426 , n26744 , new_n4023 );
xnor g09078 ( new_n11427 , n26744 , new_n4025 );
nor  g09079 ( new_n11428 , n26625 , new_n4028 );
or   g09080 ( new_n11429 , new_n9484 , new_n4031 );
xnor g09081 ( new_n11430 , n26625 , new_n4027 );
and  g09082 ( new_n11431 , new_n11429 , new_n11430 );
or   g09083 ( new_n11432 , new_n11428 , new_n11431 );
and  g09084 ( new_n11433 , new_n11427 , new_n11432 );
or   g09085 ( new_n11434 , new_n11426 , new_n11433 );
and  g09086 ( new_n11435 , new_n11425 , new_n11434 );
or   g09087 ( new_n11436 , new_n11424_1 , new_n11435 );
and  g09088 ( new_n11437 , new_n11423 , new_n11436 );
or   g09089 ( new_n11438 , new_n11422 , new_n11437 );
and  g09090 ( new_n11439_1 , new_n11421 , new_n11438 );
or   g09091 ( new_n11440 , new_n11420 , new_n11439_1 );
and  g09092 ( new_n11441 , new_n11419_1 , new_n11440 );
or   g09093 ( new_n11442 , new_n11418 , new_n11441 );
and  g09094 ( new_n11443 , new_n11417 , new_n11442 );
or   g09095 ( new_n11444 , new_n11416 , new_n11443 );
xor  g09096 ( new_n11445 , new_n11415 , new_n11444 );
nor  g09097 ( new_n11446 , n13026 , new_n11445 );
xor  g09098 ( new_n11447 , n13026 , new_n11445 );
xor  g09099 ( new_n11448 , new_n11417 , new_n11442 );
nor  g09100 ( new_n11449 , n2175 , new_n11448 );
xor  g09101 ( new_n11450 , n2175 , new_n11448 );
xor  g09102 ( new_n11451 , new_n11419_1 , new_n11440 );
nor  g09103 ( new_n11452 , n752 , new_n11451 );
xnor g09104 ( new_n11453 , n752 , new_n11451 );
xor  g09105 ( new_n11454 , new_n11421 , new_n11438 );
nor  g09106 ( new_n11455_1 , n1611 , new_n11454 );
xor  g09107 ( new_n11456 , new_n11423 , new_n11436 );
nor  g09108 ( new_n11457 , n25094 , new_n11456 );
xnor g09109 ( new_n11458 , n25094 , new_n11456 );
xor  g09110 ( new_n11459 , new_n11425 , new_n11434 );
nor  g09111 ( new_n11460 , n21538 , new_n11459 );
xnor g09112 ( new_n11461 , n21538 , new_n11459 );
xor  g09113 ( new_n11462_1 , new_n11427 , new_n11432 );
nor  g09114 ( new_n11463 , n5131 , new_n11462_1 );
xor  g09115 ( new_n11464 , new_n11429 , new_n11430 );
nor  g09116 ( new_n11465 , n11473 , new_n11464 );
xnor g09117 ( new_n11466 , new_n9484 , n19922 );
or   g09118 ( new_n11467 , new_n10803 , new_n11466 );
xnor g09119 ( new_n11468 , new_n10809 , new_n11464 );
and  g09120 ( new_n11469 , new_n11467 , new_n11468 );
nor  g09121 ( new_n11470_1 , new_n11465 , new_n11469 );
xnor g09122 ( new_n11471 , n5131 , new_n11462_1 );
nor  g09123 ( new_n11472_1 , new_n11470_1 , new_n11471 );
nor  g09124 ( new_n11473_1 , new_n11463 , new_n11472_1 );
nor  g09125 ( new_n11474 , new_n11461 , new_n11473_1 );
nor  g09126 ( new_n11475 , new_n11460 , new_n11474 );
nor  g09127 ( new_n11476 , new_n11458 , new_n11475 );
nor  g09128 ( new_n11477 , new_n11457 , new_n11476 );
xnor g09129 ( new_n11478 , n1611 , new_n11454 );
nor  g09130 ( new_n11479_1 , new_n11477 , new_n11478 );
nor  g09131 ( new_n11480 , new_n11455_1 , new_n11479_1 );
nor  g09132 ( new_n11481_1 , new_n11453 , new_n11480 );
or   g09133 ( new_n11482 , new_n11452 , new_n11481_1 );
and  g09134 ( new_n11483 , new_n11450 , new_n11482 );
or   g09135 ( new_n11484 , new_n11449 , new_n11483 );
and  g09136 ( new_n11485 , new_n11447 , new_n11484 );
nor  g09137 ( new_n11486_1 , new_n11446 , new_n11485 );
and  g09138 ( new_n11487 , n23912 , new_n11486_1 );
xnor g09139 ( new_n11488 , n23912 , new_n11486_1 );
nor  g09140 ( new_n11489 , n3984 , new_n6213 );
and  g09141 ( new_n11490 , new_n11415 , new_n11444 );
nor  g09142 ( new_n11491 , new_n11489 , new_n11490 );
not  g09143 ( new_n11492 , new_n11491 );
xnor g09144 ( new_n11493 , n4514 , new_n6208 );
xnor g09145 ( new_n11494 , new_n11492 , new_n11493 );
nor  g09146 ( new_n11495 , new_n11488 , new_n11494 );
nor  g09147 ( new_n11496_1 , new_n11487 , new_n11495 );
nor  g09148 ( new_n11497 , new_n11273_1 , new_n6208 );
nor  g09149 ( new_n11498 , n4514 , new_n6207 );
nor  g09150 ( new_n11499 , new_n11492 , new_n11498 );
or   g09151 ( new_n11500 , new_n6211 , new_n11499 );
or   g09152 ( new_n11501 , new_n11497 , new_n11500 );
and  g09153 ( new_n11502 , new_n11496_1 , new_n11501 );
nor  g09154 ( new_n11503_1 , n15766 , new_n4477 );
xnor g09155 ( new_n11504 , new_n6320 , new_n4477 );
nor  g09156 ( new_n11505 , n25629 , new_n4482 );
xnor g09157 ( new_n11506_1 , n25629 , new_n4481 );
nor  g09158 ( new_n11507 , n7692 , new_n4488 );
xnor g09159 ( new_n11508 , new_n6326 , new_n4488 );
nor  g09160 ( new_n11509 , n23039 , new_n4493 );
xnor g09161 ( new_n11510 , n23039 , new_n4493 );
nor  g09162 ( new_n11511 , n13677 , new_n3963 );
nor  g09163 ( new_n11512 , new_n3964 , new_n3995 );
nor  g09164 ( new_n11513 , new_n11511 , new_n11512 );
nor  g09165 ( new_n11514 , new_n11510 , new_n11513 );
or   g09166 ( new_n11515_1 , new_n11509 , new_n11514 );
and  g09167 ( new_n11516 , new_n11508 , new_n11515_1 );
or   g09168 ( new_n11517 , new_n11507 , new_n11516 );
and  g09169 ( new_n11518 , new_n11506_1 , new_n11517 );
or   g09170 ( new_n11519 , new_n11505 , new_n11518 );
and  g09171 ( new_n11520 , new_n11504 , new_n11519 );
nor  g09172 ( new_n11521 , new_n11503_1 , new_n11520 );
not  g09173 ( new_n11522 , new_n11521 );
nor  g09174 ( new_n11523 , new_n4538 , new_n11522 );
not  g09175 ( new_n11524 , new_n11523 );
xnor g09176 ( new_n11525 , new_n4453 , new_n11522 );
xor  g09177 ( new_n11526 , new_n11496_1 , new_n11501 );
nor  g09178 ( new_n11527 , new_n11525 , new_n11526 );
xnor g09179 ( new_n11528 , new_n11525 , new_n11526 );
xor  g09180 ( new_n11529 , new_n11504 , new_n11519 );
not  g09181 ( new_n11530 , new_n11529 );
xnor g09182 ( new_n11531 , new_n11488 , new_n11494 );
nor  g09183 ( new_n11532 , new_n11530 , new_n11531 );
xor  g09184 ( new_n11533 , new_n11506_1 , new_n11517 );
not  g09185 ( new_n11534 , new_n11533 );
xor  g09186 ( new_n11535 , new_n11447 , new_n11484 );
nor  g09187 ( new_n11536 , new_n11534 , new_n11535 );
xnor g09188 ( new_n11537 , new_n11534 , new_n11535 );
xor  g09189 ( new_n11538_1 , new_n11508 , new_n11515_1 );
not  g09190 ( new_n11539 , new_n11538_1 );
xor  g09191 ( new_n11540 , new_n11450 , new_n11482 );
nor  g09192 ( new_n11541 , new_n11539 , new_n11540 );
xnor g09193 ( new_n11542 , new_n11539 , new_n11540 );
xnor g09194 ( new_n11543 , new_n11510 , new_n11513 );
xor  g09195 ( new_n11544 , new_n11453 , new_n11480 );
nor  g09196 ( new_n11545 , new_n11543 , new_n11544 );
xnor g09197 ( new_n11546 , new_n11543 , new_n11544 );
xor  g09198 ( new_n11547 , new_n11477 , new_n11478 );
nor  g09199 ( new_n11548_1 , new_n3996 , new_n11547 );
xnor g09200 ( new_n11549 , new_n3996 , new_n11547 );
not  g09201 ( new_n11550 , new_n4080 );
xor  g09202 ( new_n11551 , new_n11458 , new_n11475 );
nor  g09203 ( new_n11552 , new_n11550 , new_n11551 );
xor  g09204 ( new_n11553 , new_n11461 , new_n11473_1 );
nor  g09205 ( new_n11554 , new_n4084 , new_n11553 );
xnor g09206 ( new_n11555 , new_n4084 , new_n11553 );
xor  g09207 ( new_n11556 , new_n11470_1 , new_n11471 );
nor  g09208 ( new_n11557 , new_n4087 , new_n11556 );
xor  g09209 ( new_n11558 , new_n11467 , new_n11468 );
nor  g09210 ( new_n11559 , new_n4092 , new_n11558 );
xnor g09211 ( new_n11560 , n15506 , new_n11466 );
nor  g09212 ( new_n11561 , new_n4094 , new_n11560 );
xnor g09213 ( new_n11562 , new_n4092 , new_n11558 );
nor  g09214 ( new_n11563 , new_n11561 , new_n11562 );
nor  g09215 ( new_n11564_1 , new_n11559 , new_n11563 );
xnor g09216 ( new_n11565 , new_n4087 , new_n11556 );
nor  g09217 ( new_n11566_1 , new_n11564_1 , new_n11565 );
nor  g09218 ( new_n11567 , new_n11557 , new_n11566_1 );
nor  g09219 ( new_n11568 , new_n11555 , new_n11567 );
nor  g09220 ( new_n11569 , new_n11554 , new_n11568 );
xnor g09221 ( new_n11570 , new_n11550 , new_n11551 );
nor  g09222 ( new_n11571 , new_n11569 , new_n11570 );
nor  g09223 ( new_n11572 , new_n11552 , new_n11571 );
nor  g09224 ( new_n11573 , new_n11549 , new_n11572 );
nor  g09225 ( new_n11574 , new_n11548_1 , new_n11573 );
nor  g09226 ( new_n11575 , new_n11546 , new_n11574 );
nor  g09227 ( new_n11576 , new_n11545 , new_n11575 );
nor  g09228 ( new_n11577 , new_n11542 , new_n11576 );
nor  g09229 ( new_n11578 , new_n11541 , new_n11577 );
nor  g09230 ( new_n11579_1 , new_n11537 , new_n11578 );
nor  g09231 ( new_n11580_1 , new_n11536 , new_n11579_1 );
xnor g09232 ( new_n11581 , new_n11530 , new_n11531 );
nor  g09233 ( new_n11582 , new_n11580_1 , new_n11581 );
nor  g09234 ( new_n11583 , new_n11532 , new_n11582 );
nor  g09235 ( new_n11584 , new_n11528 , new_n11583 );
nor  g09236 ( new_n11585 , new_n11527 , new_n11584 );
xnor g09237 ( new_n11586 , new_n11524 , new_n11585 );
xnor g09238 ( n1701 , new_n11502 , new_n11586 );
xnor g09239 ( n1703 , new_n3894 , new_n3924 );
xnor g09240 ( n1721 , new_n4551 , new_n4604 );
nor  g09241 ( new_n11590 , new_n4353 , new_n7694 );
and  g09242 ( new_n11591_1 , new_n8951 , new_n8952 );
nor  g09243 ( new_n11592 , new_n11590 , new_n11591_1 );
not  g09244 ( new_n11593 , new_n11592 );
and  g09245 ( new_n11594 , new_n8996 , new_n11593 );
nor  g09246 ( new_n11595 , new_n8953 , new_n8996 );
nor  g09247 ( new_n11596 , new_n8997 , new_n9059 );
nor  g09248 ( new_n11597 , new_n11595 , new_n11596 );
nor  g09249 ( new_n11598 , new_n11594 , new_n11597 );
nor  g09250 ( new_n11599 , new_n8996 , new_n11593 );
nor  g09251 ( new_n11600 , new_n11596 , new_n11599 );
nor  g09252 ( n1760 , new_n11598 , new_n11600 );
xnor g09253 ( n1791 , new_n4090 , new_n4098 );
xnor g09254 ( new_n11603 , n16502 , n23333 );
xnor g09255 ( n1808 , new_n11603 , new_n3368 );
nor  g09256 ( new_n11605 , new_n7650 , new_n7695 );
nor  g09257 ( new_n11606 , new_n7696 , new_n7769_1 );
nor  g09258 ( new_n11607_1 , new_n11605 , new_n11606 );
nor  g09259 ( new_n11608 , new_n3087 , n13494 );
xnor g09260 ( new_n11609 , n4319 , n13494 );
not  g09261 ( new_n11610 , n23463 );
nor  g09262 ( new_n11611 , new_n11610 , n25345 );
and  g09263 ( new_n11612 , new_n11092 , new_n11115 );
or   g09264 ( new_n11613 , new_n11611 , new_n11612 );
and  g09265 ( new_n11614 , new_n11609 , new_n11613 );
nor  g09266 ( new_n11615_1 , new_n11608 , new_n11614 );
and  g09267 ( new_n11616 , new_n11607_1 , new_n11615_1 );
nor  g09268 ( new_n11617 , new_n7770 , new_n11615_1 );
xnor g09269 ( new_n11618 , new_n7771 , new_n11615_1 );
xor  g09270 ( new_n11619 , new_n11609 , new_n11613 );
and  g09271 ( new_n11620 , new_n7837 , new_n11619 );
xnor g09272 ( new_n11621 , new_n7842 , new_n11619 );
and  g09273 ( new_n11622 , new_n7844 , new_n11116 );
and  g09274 ( new_n11623 , new_n11117 , new_n11145 );
or   g09275 ( new_n11624 , new_n11622 , new_n11623 );
and  g09276 ( new_n11625 , new_n11621 , new_n11624 );
nor  g09277 ( new_n11626 , new_n11620 , new_n11625 );
and  g09278 ( new_n11627 , new_n11618 , new_n11626 );
nor  g09279 ( new_n11628 , new_n11617 , new_n11627 );
nor  g09280 ( new_n11629 , new_n11616 , new_n11628 );
nor  g09281 ( new_n11630_1 , new_n11607_1 , new_n11615_1 );
nor  g09282 ( new_n11631 , new_n11627 , new_n11630_1 );
nor  g09283 ( n1821 , new_n11629 , new_n11631 );
xnor g09284 ( n1832 , new_n6947 , new_n6948 );
xnor g09285 ( new_n11634 , new_n7179 , n9934 );
nor  g09286 ( new_n11635 , n18496 , n25331 );
not  g09287 ( new_n11636 , n18496 );
xnor g09288 ( new_n11637 , new_n11636 , n25331 );
nor  g09289 ( new_n11638 , n18483 , n26224 );
xnor g09290 ( new_n11639 , n18483 , n26224 );
nor  g09291 ( new_n11640 , n19327 , n21934 );
xnor g09292 ( new_n11641 , n19327 , n21934 );
nor  g09293 ( new_n11642 , n18901 , n22597 );
xnor g09294 ( new_n11643 , n18901 , n22597 );
nor  g09295 ( new_n11644 , n4376 , n26107 );
xnor g09296 ( new_n11645 , n4376 , n26107 );
nor  g09297 ( new_n11646 , n342 , n14570 );
xnor g09298 ( new_n11647_1 , n342 , n14570 );
nor  g09299 ( new_n11648 , n23775 , n26553 );
xnor g09300 ( new_n11649 , n23775 , n26553 );
nor  g09301 ( new_n11650 , n4964 , n8259 );
not  g09302 ( new_n11651 , n11479 );
or   g09303 ( new_n11652 , new_n3755_1 , new_n11651 );
xnor g09304 ( new_n11653 , new_n4776 , n8259 );
and  g09305 ( new_n11654 , new_n11652 , new_n11653 );
nor  g09306 ( new_n11655 , new_n11650 , new_n11654 );
nor  g09307 ( new_n11656 , new_n11649 , new_n11655 );
nor  g09308 ( new_n11657 , new_n11648 , new_n11656 );
nor  g09309 ( new_n11658 , new_n11647_1 , new_n11657 );
nor  g09310 ( new_n11659 , new_n11646 , new_n11658 );
nor  g09311 ( new_n11660 , new_n11645 , new_n11659 );
nor  g09312 ( new_n11661 , new_n11644 , new_n11660 );
nor  g09313 ( new_n11662 , new_n11643 , new_n11661 );
nor  g09314 ( new_n11663 , new_n11642 , new_n11662 );
nor  g09315 ( new_n11664 , new_n11641 , new_n11663 );
nor  g09316 ( new_n11665 , new_n11640 , new_n11664 );
nor  g09317 ( new_n11666 , new_n11639 , new_n11665 );
or   g09318 ( new_n11667_1 , new_n11638 , new_n11666 );
and  g09319 ( new_n11668 , new_n11637 , new_n11667_1 );
or   g09320 ( new_n11669 , new_n11635 , new_n11668 );
xor  g09321 ( new_n11670 , new_n11634 , new_n11669 );
xnor g09322 ( new_n11671 , n2160 , new_n11670 );
xor  g09323 ( new_n11672 , new_n11637 , new_n11667_1 );
nor  g09324 ( new_n11673 , n10763 , new_n11672 );
not  g09325 ( new_n11674_1 , n10763 );
xnor g09326 ( new_n11675 , new_n11674_1 , new_n11672 );
xnor g09327 ( new_n11676 , new_n11639 , new_n11665 );
nor  g09328 ( new_n11677 , new_n2890 , new_n11676 );
xnor g09329 ( new_n11678 , new_n2890 , new_n11676 );
xnor g09330 ( new_n11679 , new_n11641 , new_n11663 );
nor  g09331 ( new_n11680 , new_n2893 , new_n11679 );
xnor g09332 ( new_n11681 , new_n2893 , new_n11679 );
xnor g09333 ( new_n11682_1 , new_n11643 , new_n11661 );
nor  g09334 ( new_n11683 , new_n2896 , new_n11682_1 );
xnor g09335 ( new_n11684 , new_n2896 , new_n11682_1 );
not  g09336 ( new_n11685 , n12811 );
xnor g09337 ( new_n11686 , new_n11645 , new_n11659 );
nor  g09338 ( new_n11687 , new_n11685 , new_n11686 );
xnor g09339 ( new_n11688 , new_n11685 , new_n11686 );
not  g09340 ( new_n11689 , n1118 );
xnor g09341 ( new_n11690 , new_n11647_1 , new_n11657 );
nor  g09342 ( new_n11691 , new_n11689 , new_n11690 );
xnor g09343 ( new_n11692 , new_n11689 , new_n11690 );
not  g09344 ( new_n11693 , n25974 );
xnor g09345 ( new_n11694 , new_n11649 , new_n11655 );
nor  g09346 ( new_n11695 , new_n11693 , new_n11694 );
xnor g09347 ( new_n11696 , n25974 , new_n11694 );
xnor g09348 ( new_n11697 , new_n3755_1 , n11479 );
nor  g09349 ( new_n11698 , new_n2906 , new_n11697 );
nor  g09350 ( new_n11699 , n1630 , new_n11698 );
xor  g09351 ( new_n11700 , new_n11652 , new_n11653 );
xnor g09352 ( new_n11701 , new_n2909 , new_n11698 );
not  g09353 ( new_n11702 , new_n11701 );
nor  g09354 ( new_n11703 , new_n11700 , new_n11702 );
nor  g09355 ( new_n11704 , new_n11699 , new_n11703 );
and  g09356 ( new_n11705 , new_n11696 , new_n11704 );
nor  g09357 ( new_n11706 , new_n11695 , new_n11705 );
nor  g09358 ( new_n11707 , new_n11692 , new_n11706 );
nor  g09359 ( new_n11708 , new_n11691 , new_n11707 );
nor  g09360 ( new_n11709 , new_n11688 , new_n11708 );
nor  g09361 ( new_n11710_1 , new_n11687 , new_n11709 );
nor  g09362 ( new_n11711 , new_n11684 , new_n11710_1 );
nor  g09363 ( new_n11712_1 , new_n11683 , new_n11711 );
nor  g09364 ( new_n11713 , new_n11681 , new_n11712_1 );
nor  g09365 ( new_n11714 , new_n11680 , new_n11713 );
nor  g09366 ( new_n11715 , new_n11678 , new_n11714 );
nor  g09367 ( new_n11716 , new_n11677 , new_n11715 );
and  g09368 ( new_n11717 , new_n11675 , new_n11716 );
nor  g09369 ( new_n11718 , new_n11673 , new_n11717 );
xnor g09370 ( new_n11719 , new_n11671 , new_n11718 );
not  g09371 ( new_n11720 , new_n3849 );
nor  g09372 ( new_n11721 , n4325 , new_n11720 );
not  g09373 ( new_n11722 , new_n11721 );
nor  g09374 ( new_n11723 , n11926 , new_n11722 );
not  g09375 ( new_n11724_1 , new_n11723 );
nor  g09376 ( new_n11725 , n5521 , new_n11724_1 );
xnor g09377 ( new_n11726 , n21784 , new_n11725 );
xnor g09378 ( new_n11727 , new_n7264 , new_n11726 );
xnor g09379 ( new_n11728 , n5521 , new_n11723 );
nor  g09380 ( new_n11729 , new_n7270 , new_n11728 );
xnor g09381 ( new_n11730 , new_n7270 , new_n11728 );
xnor g09382 ( new_n11731 , n11926 , new_n11721 );
nor  g09383 ( new_n11732 , new_n7275 , new_n11731 );
xnor g09384 ( new_n11733 , new_n7275 , new_n11731 );
nor  g09385 ( new_n11734 , new_n3840 , new_n3850_1 );
nor  g09386 ( new_n11735 , new_n3851 , new_n3888 );
nor  g09387 ( new_n11736_1 , new_n11734 , new_n11735 );
nor  g09388 ( new_n11737 , new_n11733 , new_n11736_1 );
nor  g09389 ( new_n11738 , new_n11732 , new_n11737 );
nor  g09390 ( new_n11739 , new_n11730 , new_n11738 );
nor  g09391 ( new_n11740 , new_n11729 , new_n11739 );
xnor g09392 ( new_n11741_1 , new_n11727 , new_n11740 );
not  g09393 ( new_n11742 , new_n11741_1 );
xnor g09394 ( new_n11743 , new_n11719 , new_n11742 );
xnor g09395 ( new_n11744 , new_n11675 , new_n11716 );
xnor g09396 ( new_n11745 , new_n11730 , new_n11738 );
not  g09397 ( new_n11746 , new_n11745 );
and  g09398 ( new_n11747 , new_n11744 , new_n11746 );
xnor g09399 ( new_n11748 , new_n11744 , new_n11746 );
xnor g09400 ( new_n11749_1 , new_n11678 , new_n11714 );
xnor g09401 ( new_n11750 , new_n11733 , new_n11736_1 );
nor  g09402 ( new_n11751 , new_n11749_1 , new_n11750 );
xnor g09403 ( new_n11752 , new_n11749_1 , new_n11750 );
xnor g09404 ( new_n11753 , new_n11681 , new_n11712_1 );
nor  g09405 ( new_n11754 , new_n3889 , new_n11753 );
xnor g09406 ( new_n11755 , new_n3889 , new_n11753 );
xnor g09407 ( new_n11756 , new_n11684 , new_n11710_1 );
nor  g09408 ( new_n11757 , new_n3891_1 , new_n11756 );
xnor g09409 ( new_n11758 , new_n3891_1 , new_n11756 );
xnor g09410 ( new_n11759 , new_n11688 , new_n11708 );
nor  g09411 ( new_n11760 , new_n3895 , new_n11759 );
xnor g09412 ( new_n11761 , new_n3895 , new_n11759 );
xnor g09413 ( new_n11762 , new_n11692 , new_n11706 );
nor  g09414 ( new_n11763 , new_n3900 , new_n11762 );
xnor g09415 ( new_n11764 , new_n3900 , new_n11762 );
xnor g09416 ( new_n11765 , new_n11696 , new_n11704 );
nor  g09417 ( new_n11766 , new_n3904 , new_n11765 );
xnor g09418 ( new_n11767 , new_n3904 , new_n11765 );
not  g09419 ( new_n11768 , new_n11767 );
xnor g09420 ( new_n11769 , n1451 , new_n11697 );
nor  g09421 ( new_n11770_1 , new_n3914 , new_n11769 );
xnor g09422 ( new_n11771_1 , new_n11700 , new_n11701 );
and  g09423 ( new_n11772 , new_n11770_1 , new_n11771_1 );
xnor g09424 ( new_n11773 , new_n11770_1 , new_n11771_1 );
nor  g09425 ( new_n11774 , new_n3908 , new_n11773 );
nor  g09426 ( new_n11775_1 , new_n11772 , new_n11774 );
and  g09427 ( new_n11776 , new_n11768 , new_n11775_1 );
nor  g09428 ( new_n11777 , new_n11766 , new_n11776 );
nor  g09429 ( new_n11778 , new_n11764 , new_n11777 );
nor  g09430 ( new_n11779 , new_n11763 , new_n11778 );
nor  g09431 ( new_n11780 , new_n11761 , new_n11779 );
nor  g09432 ( new_n11781 , new_n11760 , new_n11780 );
nor  g09433 ( new_n11782 , new_n11758 , new_n11781 );
nor  g09434 ( new_n11783 , new_n11757 , new_n11782 );
nor  g09435 ( new_n11784 , new_n11755 , new_n11783 );
nor  g09436 ( new_n11785 , new_n11754 , new_n11784 );
nor  g09437 ( new_n11786 , new_n11752 , new_n11785 );
nor  g09438 ( new_n11787 , new_n11751 , new_n11786 );
nor  g09439 ( new_n11788 , new_n11748 , new_n11787 );
nor  g09440 ( new_n11789 , new_n11747 , new_n11788 );
xnor g09441 ( n1859 , new_n11743 , new_n11789 );
xnor g09442 ( n1860 , new_n5189 , new_n5215 );
not  g09443 ( new_n11792 , new_n11323 );
nor  g09444 ( new_n11793 , new_n11320 , new_n11792 );
not  g09445 ( new_n11794 , new_n11793 );
not  g09446 ( new_n11795 , n10250 );
nor  g09447 ( new_n11796 , n15182 , n21915 );
or   g09448 ( new_n11797 , new_n6835_1 , new_n6861_1 );
and  g09449 ( new_n11798 , new_n6834 , new_n11797 );
nor  g09450 ( new_n11799 , new_n11796 , new_n11798 );
not  g09451 ( new_n11800 , new_n11799 );
xnor g09452 ( new_n11801 , new_n6198 , n25972 );
xnor g09453 ( new_n11802 , new_n11800 , new_n11801 );
not  g09454 ( new_n11803 , new_n11802 );
nor  g09455 ( new_n11804 , new_n11795 , new_n11803 );
xnor g09456 ( new_n11805 , new_n11795 , new_n11802 );
nor  g09457 ( new_n11806 , new_n6155 , new_n6863_1 );
xnor g09458 ( new_n11807 , new_n6155 , new_n6864 );
nor  g09459 ( new_n11808 , new_n6158 , new_n6867_1 );
xnor g09460 ( new_n11809 , new_n6158 , new_n6869 );
nor  g09461 ( new_n11810 , new_n6161 , new_n6872 );
xnor g09462 ( new_n11811 , new_n6161 , new_n6874 );
not  g09463 ( new_n11812 , n23586 );
nor  g09464 ( new_n11813 , new_n11812 , new_n6877 );
nor  g09465 ( new_n11814 , n21226 , new_n6881 );
xnor g09466 ( new_n11815 , n21226 , new_n6882 );
nor  g09467 ( new_n11816 , new_n6170 , new_n6886 );
xnor g09468 ( new_n11817 , new_n6170 , new_n6888 );
nor  g09469 ( new_n11818_1 , n20036 , new_n4116 );
nor  g09470 ( new_n11819 , new_n4120 , new_n4130 );
nor  g09471 ( new_n11820 , new_n6176 , new_n4135 );
xnor g09472 ( new_n11821 , new_n4120 , new_n4138 );
and  g09473 ( new_n11822 , new_n11820 , new_n11821 );
nor  g09474 ( new_n11823 , new_n11819 , new_n11822 );
xnor g09475 ( new_n11824 , new_n8659 , new_n4116 );
and  g09476 ( new_n11825 , new_n11823 , new_n11824 );
nor  g09477 ( new_n11826 , new_n11818_1 , new_n11825 );
and  g09478 ( new_n11827 , new_n11817 , new_n11826 );
nor  g09479 ( new_n11828 , new_n11816 , new_n11827 );
and  g09480 ( new_n11829 , new_n11815 , new_n11828 );
nor  g09481 ( new_n11830 , new_n11814 , new_n11829 );
xnor g09482 ( new_n11831 , new_n11812 , new_n6879 );
and  g09483 ( new_n11832 , new_n11830 , new_n11831 );
or   g09484 ( new_n11833 , new_n11813 , new_n11832 );
and  g09485 ( new_n11834 , new_n11811 , new_n11833 );
or   g09486 ( new_n11835 , new_n11810 , new_n11834 );
and  g09487 ( new_n11836 , new_n11809 , new_n11835 );
or   g09488 ( new_n11837_1 , new_n11808 , new_n11836 );
and  g09489 ( new_n11838 , new_n11807 , new_n11837_1 );
or   g09490 ( new_n11839 , new_n11806 , new_n11838 );
and  g09491 ( new_n11840 , new_n11805 , new_n11839 );
nor  g09492 ( new_n11841_1 , new_n11804 , new_n11840 );
not  g09493 ( new_n11842_1 , n25972 );
nor  g09494 ( new_n11843_1 , new_n6198 , new_n11842_1 );
nor  g09495 ( new_n11844 , n8614 , n25972 );
nor  g09496 ( new_n11845 , new_n11800 , new_n11844 );
nor  g09497 ( new_n11846 , new_n11843_1 , new_n11845 );
nor  g09498 ( new_n11847 , new_n11841_1 , new_n11846 );
nor  g09499 ( new_n11848 , new_n11794 , new_n11847 );
xnor g09500 ( new_n11849 , new_n11794 , new_n11847 );
not  g09501 ( new_n11850 , new_n11324 );
not  g09502 ( new_n11851 , new_n11846 );
xnor g09503 ( new_n11852 , new_n11841_1 , new_n11851 );
nor  g09504 ( new_n11853 , new_n11850 , new_n11852 );
xnor g09505 ( new_n11854 , new_n11850 , new_n11852 );
xor  g09506 ( new_n11855 , new_n11805 , new_n11839 );
nor  g09507 ( new_n11856 , new_n11338 , new_n11855 );
xnor g09508 ( new_n11857 , new_n11338 , new_n11855 );
not  g09509 ( new_n11858 , new_n11344 );
xor  g09510 ( new_n11859 , new_n11807 , new_n11837_1 );
nor  g09511 ( new_n11860 , new_n11858 , new_n11859 );
xnor g09512 ( new_n11861 , new_n11858 , new_n11859 );
not  g09513 ( new_n11862 , new_n11348_1 );
xor  g09514 ( new_n11863 , new_n11809 , new_n11835 );
nor  g09515 ( new_n11864 , new_n11862 , new_n11863 );
xnor g09516 ( new_n11865 , new_n11862 , new_n11863 );
xor  g09517 ( new_n11866 , new_n11811 , new_n11833 );
nor  g09518 ( new_n11867 , new_n11366 , new_n11866 );
xnor g09519 ( new_n11868 , new_n11366 , new_n11866 );
xor  g09520 ( new_n11869 , new_n11830 , new_n11831 );
nor  g09521 ( new_n11870 , new_n11358 , new_n11869 );
xnor g09522 ( new_n11871 , new_n11358 , new_n11869 );
xnor g09523 ( new_n11872 , new_n11815 , new_n11828 );
nor  g09524 ( new_n11873 , new_n9518 , new_n11872 );
xnor g09525 ( new_n11874 , new_n9518 , new_n11872 );
not  g09526 ( new_n11875 , new_n9520 );
xor  g09527 ( new_n11876 , new_n11817 , new_n11826 );
nor  g09528 ( new_n11877 , new_n11875 , new_n11876 );
xnor g09529 ( new_n11878 , new_n11875 , new_n11876 );
xnor g09530 ( new_n11879 , new_n11823 , new_n11824 );
nor  g09531 ( new_n11880 , new_n9528 , new_n11879 );
xnor g09532 ( new_n11881 , new_n9528 , new_n11879 );
xor  g09533 ( new_n11882 , new_n11820 , new_n11821 );
nor  g09534 ( new_n11883 , new_n9554_1 , new_n11882 );
xnor g09535 ( new_n11884 , n9380 , new_n4135 );
nor  g09536 ( new_n11885 , new_n7200 , new_n11884 );
xnor g09537 ( new_n11886 , new_n9530 , new_n11882 );
and  g09538 ( new_n11887 , new_n11885 , new_n11886 );
nor  g09539 ( new_n11888 , new_n11883 , new_n11887 );
nor  g09540 ( new_n11889 , new_n11881 , new_n11888 );
nor  g09541 ( new_n11890 , new_n11880 , new_n11889 );
nor  g09542 ( new_n11891 , new_n11878 , new_n11890 );
nor  g09543 ( new_n11892 , new_n11877 , new_n11891 );
nor  g09544 ( new_n11893 , new_n11874 , new_n11892 );
nor  g09545 ( new_n11894 , new_n11873 , new_n11893 );
nor  g09546 ( new_n11895 , new_n11871 , new_n11894 );
nor  g09547 ( new_n11896 , new_n11870 , new_n11895 );
nor  g09548 ( new_n11897 , new_n11868 , new_n11896 );
nor  g09549 ( new_n11898_1 , new_n11867 , new_n11897 );
nor  g09550 ( new_n11899 , new_n11865 , new_n11898_1 );
nor  g09551 ( new_n11900 , new_n11864 , new_n11899 );
nor  g09552 ( new_n11901 , new_n11861 , new_n11900 );
nor  g09553 ( new_n11902 , new_n11860 , new_n11901 );
nor  g09554 ( new_n11903 , new_n11857 , new_n11902 );
nor  g09555 ( new_n11904 , new_n11856 , new_n11903 );
nor  g09556 ( new_n11905_1 , new_n11854 , new_n11904 );
nor  g09557 ( new_n11906 , new_n11853 , new_n11905_1 );
nor  g09558 ( new_n11907 , new_n11849 , new_n11906 );
or   g09559 ( n1861 , new_n11848 , new_n11907 );
nor  g09560 ( new_n11909 , n12593 , n13714 );
not  g09561 ( new_n11910 , new_n11909 );
nor  g09562 ( new_n11911 , n19144 , new_n11910 );
not  g09563 ( new_n11912 , new_n11911 );
nor  g09564 ( new_n11913 , n8309 , new_n11912 );
not  g09565 ( new_n11914 , new_n11913 );
nor  g09566 ( new_n11915 , n19081 , new_n11914 );
not  g09567 ( new_n11916 , new_n11915 );
nor  g09568 ( new_n11917 , n26054 , new_n11916 );
xnor g09569 ( new_n11918 , n26318 , new_n11917 );
xnor g09570 ( new_n11919 , new_n5348 , new_n11918 );
xnor g09571 ( new_n11920 , n26054 , new_n11915 );
nor  g09572 ( new_n11921 , new_n5391 , new_n11920 );
xnor g09573 ( new_n11922 , n19081 , new_n11913 );
nor  g09574 ( new_n11923 , new_n5388 , new_n11922 );
xnor g09575 ( new_n11924 , new_n5388 , new_n11922 );
xnor g09576 ( new_n11925 , n8309 , new_n11911 );
nor  g09577 ( new_n11926_1 , new_n5358 , new_n11925 );
xnor g09578 ( new_n11927 , n19144 , new_n11909 );
nor  g09579 ( new_n11928 , new_n5376_1 , new_n11927 );
xnor g09580 ( new_n11929 , new_n5362 , new_n11927 );
nor  g09581 ( new_n11930 , new_n8763 , new_n5368 );
xnor g09582 ( new_n11931 , n12593 , new_n11930 );
nor  g09583 ( new_n11932 , new_n5365 , new_n11931 );
or   g09584 ( new_n11933 , new_n8763 , new_n5369 );
nor  g09585 ( new_n11934 , n12593 , new_n11933 );
nor  g09586 ( new_n11935 , new_n11932 , new_n11934 );
and  g09587 ( new_n11936 , new_n11929 , new_n11935 );
nor  g09588 ( new_n11937 , new_n11928 , new_n11936 );
xnor g09589 ( new_n11938 , new_n5358 , new_n11925 );
nor  g09590 ( new_n11939 , new_n11937 , new_n11938 );
nor  g09591 ( new_n11940 , new_n11926_1 , new_n11939 );
nor  g09592 ( new_n11941 , new_n11924 , new_n11940 );
nor  g09593 ( new_n11942 , new_n11923 , new_n11941 );
xnor g09594 ( new_n11943 , new_n5391 , new_n11920 );
nor  g09595 ( new_n11944 , new_n11942 , new_n11943 );
nor  g09596 ( new_n11945 , new_n11921 , new_n11944 );
xnor g09597 ( new_n11946 , new_n11919 , new_n11945 );
not  g09598 ( new_n11947 , new_n8577 );
nor  g09599 ( new_n11948 , n19228 , new_n11947 );
not  g09600 ( new_n11949 , new_n11948 );
nor  g09601 ( new_n11950 , n20179 , new_n11949 );
xnor g09602 ( new_n11951 , n1112 , new_n11950 );
xnor g09603 ( new_n11952 , new_n7278 , new_n11951 );
not  g09604 ( new_n11953 , new_n7282 );
xnor g09605 ( new_n11954 , n20179 , new_n11948 );
not  g09606 ( new_n11955 , new_n11954 );
nor  g09607 ( new_n11956 , new_n11953 , new_n11955 );
xnor g09608 ( new_n11957 , new_n11953 , new_n11955 );
nor  g09609 ( new_n11958 , new_n7285 , new_n8578 );
xnor g09610 ( new_n11959 , new_n7285 , new_n8578 );
nor  g09611 ( new_n11960 , new_n7288 , new_n8580 );
xnor g09612 ( new_n11961 , new_n7288 , new_n8580 );
nor  g09613 ( new_n11962 , new_n7295 , new_n8584 );
or   g09614 ( new_n11963 , new_n7293 , new_n8583 );
nor  g09615 ( new_n11964 , new_n7302 , new_n8588 );
nor  g09616 ( new_n11965_1 , new_n6771 , new_n7300 );
xnor g09617 ( new_n11966 , new_n7302 , new_n8588 );
nor  g09618 ( new_n11967 , new_n11965_1 , new_n11966 );
nor  g09619 ( new_n11968 , new_n11964 , new_n11967 );
and  g09620 ( new_n11969 , new_n11963 , new_n11968 );
or   g09621 ( new_n11970 , new_n11962 , new_n11969 );
nor  g09622 ( new_n11971 , new_n11961 , new_n11970 );
nor  g09623 ( new_n11972 , new_n11960 , new_n11971 );
nor  g09624 ( new_n11973 , new_n11959 , new_n11972 );
or   g09625 ( new_n11974 , new_n11958 , new_n11973 );
nor  g09626 ( new_n11975 , new_n11957 , new_n11974 );
nor  g09627 ( new_n11976 , new_n11956 , new_n11975 );
xor  g09628 ( new_n11977 , new_n11952 , new_n11976 );
xnor g09629 ( new_n11978 , new_n11946 , new_n11977 );
xnor g09630 ( new_n11979 , new_n11957 , new_n11974 );
xnor g09631 ( new_n11980_1 , new_n11942 , new_n11943 );
not  g09632 ( new_n11981 , new_n11980_1 );
and  g09633 ( new_n11982 , new_n11979 , new_n11981 );
xnor g09634 ( new_n11983 , new_n11979 , new_n11981 );
xnor g09635 ( new_n11984 , new_n11924 , new_n11940 );
xnor g09636 ( new_n11985 , new_n11959 , new_n11972 );
nor  g09637 ( new_n11986 , new_n11984 , new_n11985 );
xnor g09638 ( new_n11987 , new_n11984 , new_n11985 );
xnor g09639 ( new_n11988 , new_n11937 , new_n11938 );
xnor g09640 ( new_n11989 , new_n11961 , new_n11970 );
nor  g09641 ( new_n11990 , new_n11988 , new_n11989 );
xnor g09642 ( new_n11991 , new_n11988 , new_n11989 );
xnor g09643 ( new_n11992 , new_n11929 , new_n11935 );
xnor g09644 ( new_n11993 , new_n7295 , new_n8584 );
xnor g09645 ( new_n11994 , new_n11968 , new_n11993 );
nor  g09646 ( new_n11995 , new_n11992 , new_n11994 );
xnor g09647 ( new_n11996 , new_n11992 , new_n11994 );
xnor g09648 ( new_n11997 , new_n11965_1 , new_n11966 );
xnor g09649 ( new_n11998 , new_n5372 , new_n11931 );
nor  g09650 ( new_n11999 , new_n11997 , new_n11998 );
xnor g09651 ( new_n12000_1 , n18962 , new_n7300 );
not  g09652 ( new_n12001 , new_n12000_1 );
xnor g09653 ( new_n12002 , new_n8763 , new_n5369 );
nor  g09654 ( new_n12003_1 , new_n12001 , new_n12002 );
xnor g09655 ( new_n12004 , new_n11997 , new_n11998 );
nor  g09656 ( new_n12005 , new_n12003_1 , new_n12004 );
nor  g09657 ( new_n12006 , new_n11999 , new_n12005 );
nor  g09658 ( new_n12007 , new_n11996 , new_n12006 );
nor  g09659 ( new_n12008 , new_n11995 , new_n12007 );
nor  g09660 ( new_n12009 , new_n11991 , new_n12008 );
nor  g09661 ( new_n12010 , new_n11990 , new_n12009 );
nor  g09662 ( new_n12011_1 , new_n11987 , new_n12010 );
nor  g09663 ( new_n12012 , new_n11986 , new_n12011_1 );
nor  g09664 ( new_n12013 , new_n11983 , new_n12012 );
nor  g09665 ( new_n12014 , new_n11982 , new_n12013 );
xnor g09666 ( n1891 , new_n11978 , new_n12014 );
xnor g09667 ( new_n12016 , n1949 , n20169 );
and  g09668 ( new_n12017 , new_n6173 , n9323 );
nor  g09669 ( new_n12018 , new_n6173 , n9323 );
and  g09670 ( new_n12019 , new_n6178 , n10792 );
or   g09671 ( new_n12020 , new_n6178 , n10792 );
nor  g09672 ( new_n12021 , new_n4031 , n21687 );
and  g09673 ( new_n12022 , new_n12020 , new_n12021 );
nor  g09674 ( new_n12023 , new_n12019 , new_n12022 );
nor  g09675 ( new_n12024 , new_n12018 , new_n12023 );
or   g09676 ( new_n12025 , new_n12017 , new_n12024 );
xor  g09677 ( new_n12026 , new_n12016 , new_n12025 );
xnor g09678 ( new_n12027 , new_n6560_1 , new_n12026 );
xnor g09679 ( new_n12028 , n8285 , n9323 );
xnor g09680 ( new_n12029 , new_n12023 , new_n12028 );
and  g09681 ( new_n12030 , new_n6566 , new_n12029 );
xnor g09682 ( new_n12031 , new_n6566 , new_n12029 );
xnor g09683 ( new_n12032 , n19922 , n21687 );
nor  g09684 ( new_n12033 , new_n6568 , new_n12032 );
xnor g09685 ( new_n12034 , n6729 , n10792 );
xnor g09686 ( new_n12035 , new_n12021 , new_n12034 );
nor  g09687 ( new_n12036 , new_n12033 , new_n12035 );
xnor g09688 ( new_n12037 , new_n12033 , new_n12035 );
nor  g09689 ( new_n12038 , new_n6571 , new_n12037 );
nor  g09690 ( new_n12039 , new_n12036 , new_n12038 );
nor  g09691 ( new_n12040 , new_n12031 , new_n12039 );
nor  g09692 ( new_n12041 , new_n12030 , new_n12040 );
xnor g09693 ( n1925 , new_n12027 , new_n12041 );
xnor g09694 ( n1942 , new_n7570 , new_n7594 );
xnor g09695 ( n1972 , new_n6365 , new_n6419 );
and  g09696 ( new_n12045 , new_n8718 , new_n8785 );
nor  g09697 ( new_n12046 , new_n8786 , new_n8852 );
nor  g09698 ( new_n12047 , new_n12045 , new_n12046 );
not  g09699 ( new_n12048 , n22764 );
and  g09700 ( new_n12049 , new_n12048 , new_n8734 );
and  g09701 ( new_n12050 , n12507 , new_n8735 );
nor  g09702 ( new_n12051 , n12507 , new_n8735 );
nor  g09703 ( new_n12052 , new_n12051 , new_n8784 );
or   g09704 ( new_n12053 , new_n12050 , new_n12052 );
nor  g09705 ( new_n12054 , new_n12049 , new_n12053 );
and  g09706 ( new_n12055 , new_n11026 , new_n12054 );
and  g09707 ( new_n12056 , new_n12047 , new_n12055 );
or   g09708 ( new_n12057 , new_n11026 , new_n12054 );
nor  g09709 ( new_n12058 , new_n12047 , new_n12057 );
nor  g09710 ( new_n12059 , new_n12056 , new_n12058 );
and  g09711 ( new_n12060 , new_n11018 , new_n12059 );
xnor g09712 ( new_n12061 , new_n10912 , new_n12059 );
xnor g09713 ( new_n12062 , new_n11025_1 , new_n12054 );
xnor g09714 ( new_n12063 , new_n12047 , new_n12062 );
not  g09715 ( new_n12064 , new_n12063 );
nor  g09716 ( new_n12065 , new_n10912 , new_n12064 );
xnor g09717 ( new_n12066 , new_n10912 , new_n12064 );
not  g09718 ( new_n12067 , new_n8853 );
nor  g09719 ( new_n12068 , new_n12067 , new_n10957 );
nor  g09720 ( new_n12069 , new_n8856_1 , new_n10964 );
xnor g09721 ( new_n12070 , new_n8856_1 , new_n10964 );
nor  g09722 ( new_n12071 , new_n8860 , new_n10968 );
xnor g09723 ( new_n12072_1 , new_n8860 , new_n10968 );
nor  g09724 ( new_n12073 , new_n8864 , new_n10973 );
xnor g09725 ( new_n12074 , new_n8864 , new_n10973 );
nor  g09726 ( new_n12075 , new_n8868 , new_n10977 );
xnor g09727 ( new_n12076 , new_n8868 , new_n10977 );
nor  g09728 ( new_n12077 , new_n8872 , new_n10982 );
xnor g09729 ( new_n12078 , new_n8872 , new_n10982 );
nor  g09730 ( new_n12079 , new_n8875 , new_n10985 );
xnor g09731 ( new_n12080 , new_n8876 , new_n10984 );
and  g09732 ( new_n12081 , new_n8880 , new_n10989 );
xnor g09733 ( new_n12082 , new_n8880 , new_n10989 );
nor  g09734 ( new_n12083 , new_n8886 , new_n10992 );
nor  g09735 ( new_n12084 , new_n10996 , new_n12083 );
xnor g09736 ( new_n12085 , new_n10995 , new_n12083 );
and  g09737 ( new_n12086 , new_n8891 , new_n12085 );
nor  g09738 ( new_n12087 , new_n12084 , new_n12086 );
nor  g09739 ( new_n12088 , new_n12082 , new_n12087 );
nor  g09740 ( new_n12089 , new_n12081 , new_n12088 );
nor  g09741 ( new_n12090 , new_n12080 , new_n12089 );
nor  g09742 ( new_n12091 , new_n12079 , new_n12090 );
nor  g09743 ( new_n12092 , new_n12078 , new_n12091 );
nor  g09744 ( new_n12093 , new_n12077 , new_n12092 );
nor  g09745 ( new_n12094 , new_n12076 , new_n12093 );
nor  g09746 ( new_n12095 , new_n12075 , new_n12094 );
nor  g09747 ( new_n12096 , new_n12074 , new_n12095 );
nor  g09748 ( new_n12097 , new_n12073 , new_n12096 );
nor  g09749 ( new_n12098 , new_n12072_1 , new_n12097 );
nor  g09750 ( new_n12099 , new_n12071 , new_n12098 );
nor  g09751 ( new_n12100 , new_n12070 , new_n12099 );
nor  g09752 ( new_n12101 , new_n12069 , new_n12100 );
xnor g09753 ( new_n12102 , new_n12067 , new_n10957 );
nor  g09754 ( new_n12103 , new_n12101 , new_n12102 );
nor  g09755 ( new_n12104 , new_n12068 , new_n12103 );
nor  g09756 ( new_n12105 , new_n12066 , new_n12104 );
nor  g09757 ( new_n12106 , new_n12065 , new_n12105 );
and  g09758 ( new_n12107 , new_n12061 , new_n12106 );
nor  g09759 ( n1981 , new_n12060 , new_n12107 );
xnor g09760 ( n2004 , new_n12101 , new_n12102 );
not  g09761 ( new_n12110 , n5140 );
nor  g09762 ( new_n12111 , new_n12110 , n6105 );
xnor g09763 ( new_n12112 , n5140 , n6105 );
not  g09764 ( new_n12113_1 , n6204 );
nor  g09765 ( new_n12114 , n3795 , new_n12113_1 );
xnor g09766 ( new_n12115 , n3795 , n6204 );
not  g09767 ( new_n12116 , n3349 );
nor  g09768 ( new_n12117 , new_n12116 , n25464 );
xnor g09769 ( new_n12118 , n3349 , n25464 );
not  g09770 ( new_n12119 , n1742 );
nor  g09771 ( new_n12120 , new_n12119 , n4590 );
xnor g09772 ( new_n12121_1 , n1742 , n4590 );
not  g09773 ( new_n12122 , n4858 );
nor  g09774 ( new_n12123 , new_n12122 , n26752 );
xnor g09775 ( new_n12124 , n4858 , n26752 );
not  g09776 ( new_n12125 , n8244 );
nor  g09777 ( new_n12126 , n6513 , new_n12125 );
xnor g09778 ( new_n12127 , n6513 , n8244 );
not  g09779 ( new_n12128 , n9493 );
nor  g09780 ( new_n12129 , n3918 , new_n12128 );
xnor g09781 ( new_n12130 , n3918 , n9493 );
nor  g09782 ( new_n12131_1 , new_n4143 , n15167 );
not  g09783 ( new_n12132 , n15167 );
nor  g09784 ( new_n12133 , n919 , new_n12132 );
not  g09785 ( new_n12134 , n21095 );
and  g09786 ( new_n12135 , new_n12134 , n25316 );
nor  g09787 ( new_n12136 , new_n12134 , n25316 );
nor  g09788 ( new_n12137 , n8656 , new_n4146_1 );
not  g09789 ( new_n12138 , new_n12137 );
nor  g09790 ( new_n12139 , new_n12136 , new_n12138 );
nor  g09791 ( new_n12140 , new_n12135 , new_n12139 );
nor  g09792 ( new_n12141 , new_n12133 , new_n12140 );
nor  g09793 ( new_n12142 , new_n12131_1 , new_n12141 );
and  g09794 ( new_n12143 , new_n12130 , new_n12142 );
or   g09795 ( new_n12144 , new_n12129 , new_n12143 );
and  g09796 ( new_n12145 , new_n12127 , new_n12144 );
or   g09797 ( new_n12146_1 , new_n12126 , new_n12145 );
and  g09798 ( new_n12147 , new_n12124 , new_n12146_1 );
or   g09799 ( new_n12148 , new_n12123 , new_n12147 );
and  g09800 ( new_n12149 , new_n12121_1 , new_n12148 );
or   g09801 ( new_n12150 , new_n12120 , new_n12149 );
and  g09802 ( new_n12151 , new_n12118 , new_n12150 );
or   g09803 ( new_n12152_1 , new_n12117 , new_n12151 );
and  g09804 ( new_n12153_1 , new_n12115 , new_n12152_1 );
or   g09805 ( new_n12154 , new_n12114 , new_n12153_1 );
and  g09806 ( new_n12155 , new_n12112 , new_n12154 );
nor  g09807 ( new_n12156 , new_n12111 , new_n12155 );
nor  g09808 ( new_n12157_1 , n10018 , new_n6208 );
not  g09809 ( new_n12158_1 , n10018 );
nor  g09810 ( new_n12159 , new_n12158_1 , new_n6207 );
nor  g09811 ( new_n12160 , n2184 , new_n6216 );
xnor g09812 ( new_n12161_1 , n2184 , new_n6213 );
nor  g09813 ( new_n12162 , n3541 , new_n6220 );
xnor g09814 ( new_n12163 , n3541 , new_n6218_1 );
nor  g09815 ( new_n12164 , n16818 , new_n6224 );
xnor g09816 ( new_n12165 , n16818 , new_n6223_1 );
nor  g09817 ( new_n12166 , n1269 , new_n4013 );
xnor g09818 ( new_n12167 , n1269 , new_n4012 );
nor  g09819 ( new_n12168 , n14576 , new_n4017 );
xnor g09820 ( new_n12169 , n14576 , new_n4016 );
not  g09821 ( new_n12170 , n2985 );
nor  g09822 ( new_n12171 , new_n12170 , new_n4019 );
xnor g09823 ( new_n12172 , n2985 , new_n4019 );
nor  g09824 ( new_n12173 , n5605 , new_n4025 );
and  g09825 ( new_n12174 , n15652 , new_n4027 );
nor  g09826 ( new_n12175 , new_n6491 , n19922 );
xnor g09827 ( new_n12176 , n15652 , new_n4028 );
and  g09828 ( new_n12177 , new_n12175 , new_n12176 );
nor  g09829 ( new_n12178 , new_n12174 , new_n12177 );
xnor g09830 ( new_n12179_1 , n5605 , new_n4023 );
and  g09831 ( new_n12180 , new_n12178 , new_n12179_1 );
nor  g09832 ( new_n12181 , new_n12173 , new_n12180 );
and  g09833 ( new_n12182 , new_n12172 , new_n12181 );
nor  g09834 ( new_n12183 , new_n12171 , new_n12182 );
and  g09835 ( new_n12184 , new_n12169 , new_n12183 );
or   g09836 ( new_n12185 , new_n12168 , new_n12184 );
and  g09837 ( new_n12186 , new_n12167 , new_n12185 );
or   g09838 ( new_n12187 , new_n12166 , new_n12186 );
and  g09839 ( new_n12188 , new_n12165 , new_n12187 );
or   g09840 ( new_n12189 , new_n12164 , new_n12188 );
and  g09841 ( new_n12190 , new_n12163 , new_n12189 );
or   g09842 ( new_n12191 , new_n12162 , new_n12190 );
and  g09843 ( new_n12192_1 , new_n12161_1 , new_n12191 );
nor  g09844 ( new_n12193 , new_n12160 , new_n12192_1 );
nor  g09845 ( new_n12194 , new_n12159 , new_n12193 );
xor  g09846 ( new_n12195 , new_n6211 , new_n12194 );
nor  g09847 ( new_n12196 , new_n12157_1 , new_n12195 );
xnor g09848 ( new_n12197 , new_n6242 , new_n12196 );
xnor g09849 ( new_n12198 , new_n12158_1 , new_n6208 );
xnor g09850 ( new_n12199 , new_n12193 , new_n12198 );
not  g09851 ( new_n12200 , new_n12199 );
and  g09852 ( new_n12201 , new_n6244 , new_n12200 );
xnor g09853 ( new_n12202 , new_n6244 , new_n12200 );
xor  g09854 ( new_n12203 , new_n12161_1 , new_n12191 );
nor  g09855 ( new_n12204 , new_n6251 , new_n12203 );
xnor g09856 ( new_n12205 , new_n6251 , new_n12203 );
xor  g09857 ( new_n12206 , new_n12163 , new_n12189 );
nor  g09858 ( new_n12207 , new_n6257 , new_n12206 );
xnor g09859 ( new_n12208 , new_n6257 , new_n12206 );
xor  g09860 ( new_n12209_1 , new_n12165 , new_n12187 );
nor  g09861 ( new_n12210 , new_n6304 , new_n12209_1 );
xor  g09862 ( new_n12211 , new_n12167 , new_n12185 );
nor  g09863 ( new_n12212 , new_n6269 , new_n12211 );
xnor g09864 ( new_n12213 , new_n6269 , new_n12211 );
xor  g09865 ( new_n12214 , new_n12169 , new_n12183 );
nor  g09866 ( new_n12215 , new_n6274 , new_n12214 );
xnor g09867 ( new_n12216 , new_n6274 , new_n12214 );
xnor g09868 ( new_n12217 , new_n12172 , new_n12181 );
nor  g09869 ( new_n12218 , new_n6277 , new_n12217 );
xnor g09870 ( new_n12219 , new_n12178 , new_n12179_1 );
nor  g09871 ( new_n12220 , new_n6280 , new_n12219 );
xnor g09872 ( new_n12221 , new_n6280 , new_n12219 );
xor  g09873 ( new_n12222 , new_n12175 , new_n12176 );
nor  g09874 ( new_n12223_1 , new_n6285 , new_n12222 );
xnor g09875 ( new_n12224 , n4939 , n19922 );
nor  g09876 ( new_n12225_1 , new_n6288 , new_n12224 );
not  g09877 ( new_n12226 , new_n6285 );
xnor g09878 ( new_n12227 , new_n12226 , new_n12222 );
and  g09879 ( new_n12228_1 , new_n12225_1 , new_n12227 );
nor  g09880 ( new_n12229 , new_n12223_1 , new_n12228_1 );
nor  g09881 ( new_n12230 , new_n12221 , new_n12229 );
nor  g09882 ( new_n12231 , new_n12220 , new_n12230 );
xnor g09883 ( new_n12232 , new_n6276_1 , new_n12217 );
and  g09884 ( new_n12233 , new_n12231 , new_n12232 );
nor  g09885 ( new_n12234 , new_n12218 , new_n12233 );
nor  g09886 ( new_n12235_1 , new_n12216 , new_n12234 );
nor  g09887 ( new_n12236 , new_n12215 , new_n12235_1 );
nor  g09888 ( new_n12237 , new_n12213 , new_n12236 );
nor  g09889 ( new_n12238 , new_n12212 , new_n12237 );
xnor g09890 ( new_n12239 , new_n6304 , new_n12209_1 );
nor  g09891 ( new_n12240 , new_n12238 , new_n12239 );
nor  g09892 ( new_n12241 , new_n12210 , new_n12240 );
nor  g09893 ( new_n12242 , new_n12208 , new_n12241 );
nor  g09894 ( new_n12243 , new_n12207 , new_n12242 );
nor  g09895 ( new_n12244 , new_n12205 , new_n12243 );
nor  g09896 ( new_n12245 , new_n12204 , new_n12244 );
nor  g09897 ( new_n12246 , new_n12202 , new_n12245 );
nor  g09898 ( new_n12247 , new_n12201 , new_n12246 );
xnor g09899 ( new_n12248 , new_n12197 , new_n12247 );
nor  g09900 ( new_n12249 , new_n12156 , new_n12248 );
xnor g09901 ( new_n12250 , new_n12156 , new_n12248 );
xor  g09902 ( new_n12251 , new_n12112 , new_n12154 );
xnor g09903 ( new_n12252 , new_n12202 , new_n12245 );
nor  g09904 ( new_n12253 , new_n12251 , new_n12252 );
xnor g09905 ( new_n12254 , new_n12251 , new_n12252 );
xor  g09906 ( new_n12255 , new_n12115 , new_n12152_1 );
xnor g09907 ( new_n12256 , new_n12205 , new_n12243 );
nor  g09908 ( new_n12257 , new_n12255 , new_n12256 );
xnor g09909 ( new_n12258 , new_n12255 , new_n12256 );
xor  g09910 ( new_n12259 , new_n12118 , new_n12150 );
xnor g09911 ( new_n12260 , new_n12208 , new_n12241 );
nor  g09912 ( new_n12261 , new_n12259 , new_n12260 );
xnor g09913 ( new_n12262 , new_n12259 , new_n12260 );
xor  g09914 ( new_n12263 , new_n12121_1 , new_n12148 );
xnor g09915 ( new_n12264 , new_n12238 , new_n12239 );
nor  g09916 ( new_n12265 , new_n12263 , new_n12264 );
xnor g09917 ( new_n12266 , new_n12263 , new_n12264 );
xor  g09918 ( new_n12267 , new_n12124 , new_n12146_1 );
xnor g09919 ( new_n12268 , new_n12213 , new_n12236 );
nor  g09920 ( new_n12269 , new_n12267 , new_n12268 );
xnor g09921 ( new_n12270 , new_n12267 , new_n12268 );
xor  g09922 ( new_n12271 , new_n12127 , new_n12144 );
xnor g09923 ( new_n12272 , new_n12216 , new_n12234 );
nor  g09924 ( new_n12273 , new_n12271 , new_n12272 );
xnor g09925 ( new_n12274 , new_n12271 , new_n12272 );
xnor g09926 ( new_n12275 , new_n12130 , new_n12142 );
xnor g09927 ( new_n12276 , new_n12231 , new_n12232 );
not  g09928 ( new_n12277 , new_n12276 );
and  g09929 ( new_n12278 , new_n12275 , new_n12277 );
xnor g09930 ( new_n12279 , new_n12275 , new_n12277 );
xnor g09931 ( new_n12280 , new_n12221 , new_n12229 );
xnor g09932 ( new_n12281 , n919 , n15167 );
xnor g09933 ( new_n12282 , new_n12140 , new_n12281 );
and  g09934 ( new_n12283 , new_n12280 , new_n12282 );
xnor g09935 ( new_n12284 , new_n12280 , new_n12282 );
xnor g09936 ( new_n12285 , new_n6287 , new_n12224 );
not  g09937 ( new_n12286 , new_n12285 );
xnor g09938 ( new_n12287 , n8656 , n20385 );
nor  g09939 ( new_n12288 , new_n12286 , new_n12287 );
xnor g09940 ( new_n12289 , n21095 , n25316 );
xnor g09941 ( new_n12290 , new_n12138 , new_n12289 );
not  g09942 ( new_n12291 , new_n12290 );
nor  g09943 ( new_n12292 , new_n12288 , new_n12291 );
xnor g09944 ( new_n12293 , new_n12225_1 , new_n12227 );
xnor g09945 ( new_n12294 , new_n12288 , new_n12290 );
and  g09946 ( new_n12295 , new_n12293 , new_n12294 );
nor  g09947 ( new_n12296 , new_n12292 , new_n12295 );
nor  g09948 ( new_n12297 , new_n12284 , new_n12296 );
nor  g09949 ( new_n12298 , new_n12283 , new_n12297 );
nor  g09950 ( new_n12299 , new_n12279 , new_n12298 );
nor  g09951 ( new_n12300 , new_n12278 , new_n12299 );
nor  g09952 ( new_n12301 , new_n12274 , new_n12300 );
nor  g09953 ( new_n12302_1 , new_n12273 , new_n12301 );
nor  g09954 ( new_n12303 , new_n12270 , new_n12302_1 );
nor  g09955 ( new_n12304_1 , new_n12269 , new_n12303 );
nor  g09956 ( new_n12305 , new_n12266 , new_n12304_1 );
nor  g09957 ( new_n12306 , new_n12265 , new_n12305 );
nor  g09958 ( new_n12307 , new_n12262 , new_n12306 );
nor  g09959 ( new_n12308 , new_n12261 , new_n12307 );
nor  g09960 ( new_n12309 , new_n12258 , new_n12308 );
nor  g09961 ( new_n12310 , new_n12257 , new_n12309 );
nor  g09962 ( new_n12311 , new_n12254 , new_n12310 );
nor  g09963 ( new_n12312 , new_n12253 , new_n12311 );
nor  g09964 ( new_n12313 , new_n12250 , new_n12312 );
nor  g09965 ( new_n12314 , new_n12249 , new_n12313 );
not  g09966 ( new_n12315_1 , new_n12314 );
nor  g09967 ( new_n12316 , new_n6242 , new_n12196 );
and  g09968 ( new_n12317 , new_n6211 , new_n12194 );
nand g09969 ( new_n12318 , new_n6242 , new_n12196 );
and  g09970 ( new_n12319 , new_n12318 , new_n12247 );
or   g09971 ( new_n12320 , new_n12317 , new_n12319 );
nor  g09972 ( new_n12321 , new_n12316 , new_n12320 );
and  g09973 ( n2007 , new_n12315_1 , new_n12321 );
xnor g09974 ( n2061 , new_n8884_1 , new_n8895 );
xnor g09975 ( new_n12324_1 , new_n7122 , new_n11205 );
nor  g09976 ( new_n12325_1 , new_n7126 , new_n11209 );
xnor g09977 ( new_n12326 , new_n7126 , new_n11209 );
nor  g09978 ( new_n12327 , new_n7130 , new_n11214 );
nor  g09979 ( new_n12328 , new_n4660 , new_n7134 );
xnor g09980 ( new_n12329_1 , new_n4660 , new_n7134 );
nor  g09981 ( new_n12330_1 , new_n4687 , new_n7138 );
xnor g09982 ( new_n12331 , new_n4687 , new_n7138 );
and  g09983 ( new_n12332 , new_n4691 , new_n7141 );
nor  g09984 ( new_n12333 , new_n4699 , new_n7144 );
xnor g09985 ( new_n12334 , new_n4699 , new_n7145 );
nor  g09986 ( new_n12335 , new_n4710 , new_n7150 );
and  g09987 ( new_n12336 , new_n4713 , new_n12335 );
xnor g09988 ( new_n12337 , new_n4706 , new_n12335 );
and  g09989 ( new_n12338 , new_n7157 , new_n12337 );
nor  g09990 ( new_n12339 , new_n12336 , new_n12338 );
and  g09991 ( new_n12340 , new_n12334 , new_n12339 );
nor  g09992 ( new_n12341_1 , new_n12333 , new_n12340 );
xnor g09993 ( new_n12342 , new_n4691 , new_n7141 );
nor  g09994 ( new_n12343 , new_n12341_1 , new_n12342 );
nor  g09995 ( new_n12344 , new_n12332 , new_n12343 );
nor  g09996 ( new_n12345 , new_n12331 , new_n12344 );
nor  g09997 ( new_n12346_1 , new_n12330_1 , new_n12345 );
nor  g09998 ( new_n12347 , new_n12329_1 , new_n12346_1 );
nor  g09999 ( new_n12348 , new_n12328 , new_n12347 );
xnor g10000 ( new_n12349_1 , new_n7130 , new_n11214 );
nor  g10001 ( new_n12350 , new_n12348 , new_n12349_1 );
nor  g10002 ( new_n12351 , new_n12327 , new_n12350 );
nor  g10003 ( new_n12352 , new_n12326 , new_n12351 );
nor  g10004 ( new_n12353 , new_n12325_1 , new_n12352 );
xnor g10005 ( n2092 , new_n12324_1 , new_n12353 );
xnor g10006 ( new_n12355 , n10650 , n22253 );
nor  g10007 ( new_n12356 , n1255 , n12900 );
xnor g10008 ( new_n12357 , n1255 , n12900 );
nor  g10009 ( new_n12358 , n9512 , n20411 );
xnor g10010 ( new_n12359 , n9512 , n20411 );
nor  g10011 ( new_n12360 , n16608 , n17069 );
xnor g10012 ( new_n12361 , n16608 , n17069 );
nor  g10013 ( new_n12362 , n15918 , n21735 );
xnor g10014 ( new_n12363 , n15918 , n21735 );
nor  g10015 ( new_n12364_1 , n17784 , n24085 );
xnor g10016 ( new_n12365 , n17784 , n24085 );
nor  g10017 ( new_n12366 , n14071 , n14323 );
xnor g10018 ( new_n12367 , n14071 , n14323 );
nor  g10019 ( new_n12368 , n1738 , n2886 );
xnor g10020 ( new_n12369 , n1738 , n2886 );
nor  g10021 ( new_n12370 , n1040 , n12152 );
not  g10022 ( new_n12371 , n9090 );
or   g10023 ( new_n12372 , new_n12371 , new_n7025 );
not  g10024 ( new_n12373 , n1040 );
xnor g10025 ( new_n12374 , new_n12373 , n12152 );
and  g10026 ( new_n12375 , new_n12372 , new_n12374 );
nor  g10027 ( new_n12376 , new_n12370 , new_n12375 );
nor  g10028 ( new_n12377 , new_n12369 , new_n12376 );
nor  g10029 ( new_n12378 , new_n12368 , new_n12377 );
nor  g10030 ( new_n12379 , new_n12367 , new_n12378 );
nor  g10031 ( new_n12380_1 , new_n12366 , new_n12379 );
nor  g10032 ( new_n12381 , new_n12365 , new_n12380_1 );
nor  g10033 ( new_n12382 , new_n12364_1 , new_n12381 );
nor  g10034 ( new_n12383_1 , new_n12363 , new_n12382 );
nor  g10035 ( new_n12384_1 , new_n12362 , new_n12383_1 );
nor  g10036 ( new_n12385 , new_n12361 , new_n12384_1 );
nor  g10037 ( new_n12386 , new_n12360 , new_n12385 );
nor  g10038 ( new_n12387 , new_n12359 , new_n12386 );
nor  g10039 ( new_n12388 , new_n12358 , new_n12387 );
nor  g10040 ( new_n12389 , new_n12357 , new_n12388 );
nor  g10041 ( new_n12390 , new_n12356 , new_n12389 );
xnor g10042 ( new_n12391 , new_n12355 , new_n12390 );
nor  g10043 ( new_n12392 , new_n7179 , new_n12391 );
xnor g10044 ( new_n12393 , new_n7179 , new_n12391 );
xnor g10045 ( new_n12394 , new_n12357 , new_n12388 );
nor  g10046 ( new_n12395 , new_n6967_1 , new_n12394 );
xnor g10047 ( new_n12396 , new_n6967_1 , new_n12394 );
xnor g10048 ( new_n12397_1 , new_n12359 , new_n12386 );
nor  g10049 ( new_n12398_1 , new_n6970 , new_n12397_1 );
xnor g10050 ( new_n12399 , new_n6970 , new_n12397_1 );
xnor g10051 ( new_n12400 , new_n12361 , new_n12384_1 );
nor  g10052 ( new_n12401 , new_n6973 , new_n12400 );
xnor g10053 ( new_n12402 , new_n6973 , new_n12400 );
xnor g10054 ( new_n12403 , new_n12363 , new_n12382 );
nor  g10055 ( new_n12404 , new_n6976 , new_n12403 );
xnor g10056 ( new_n12405 , new_n6976 , new_n12403 );
xnor g10057 ( new_n12406 , new_n12365 , new_n12380_1 );
nor  g10058 ( new_n12407 , new_n6979 , new_n12406 );
xnor g10059 ( new_n12408_1 , new_n6979 , new_n12406 );
xnor g10060 ( new_n12409 , new_n12367 , new_n12378 );
nor  g10061 ( new_n12410 , new_n6982 , new_n12409 );
xnor g10062 ( new_n12411 , new_n6982 , new_n12409 );
xnor g10063 ( new_n12412 , new_n12369 , new_n12376 );
nor  g10064 ( new_n12413 , new_n6986 , new_n12412 );
xnor g10065 ( new_n12414 , n23775 , new_n12412 );
xnor g10066 ( new_n12415 , new_n12371 , n19107 );
nor  g10067 ( new_n12416 , new_n11651 , new_n12415 );
nor  g10068 ( new_n12417 , n8259 , new_n12416 );
xor  g10069 ( new_n12418 , new_n12372 , new_n12374 );
xnor g10070 ( new_n12419 , new_n6989 , new_n12416 );
not  g10071 ( new_n12420 , new_n12419 );
nor  g10072 ( new_n12421 , new_n12418 , new_n12420 );
nor  g10073 ( new_n12422 , new_n12417 , new_n12421 );
and  g10074 ( new_n12423 , new_n12414 , new_n12422 );
nor  g10075 ( new_n12424 , new_n12413 , new_n12423 );
nor  g10076 ( new_n12425 , new_n12411 , new_n12424 );
nor  g10077 ( new_n12426 , new_n12410 , new_n12425 );
nor  g10078 ( new_n12427 , new_n12408_1 , new_n12426 );
nor  g10079 ( new_n12428 , new_n12407 , new_n12427 );
nor  g10080 ( new_n12429 , new_n12405 , new_n12428 );
nor  g10081 ( new_n12430 , new_n12404 , new_n12429 );
nor  g10082 ( new_n12431 , new_n12402 , new_n12430 );
nor  g10083 ( new_n12432 , new_n12401 , new_n12431 );
nor  g10084 ( new_n12433 , new_n12399 , new_n12432 );
nor  g10085 ( new_n12434 , new_n12398_1 , new_n12433 );
nor  g10086 ( new_n12435 , new_n12396 , new_n12434 );
nor  g10087 ( new_n12436 , new_n12395 , new_n12435 );
nor  g10088 ( new_n12437 , new_n12393 , new_n12436 );
nor  g10089 ( new_n12438 , new_n12392 , new_n12437 );
nor  g10090 ( new_n12439 , n10650 , n22253 );
nor  g10091 ( new_n12440 , new_n12355 , new_n12390 );
nor  g10092 ( new_n12441 , new_n12439 , new_n12440 );
nor  g10093 ( new_n12442 , new_n12438 , new_n12441 );
not  g10094 ( new_n12443 , n9934 );
nor  g10095 ( new_n12444 , n4964 , n7876 );
not  g10096 ( new_n12445 , new_n12444 );
nor  g10097 ( new_n12446_1 , n26553 , new_n12445 );
not  g10098 ( new_n12447 , new_n12446_1 );
nor  g10099 ( new_n12448 , n342 , new_n12447 );
not  g10100 ( new_n12449_1 , new_n12448 );
nor  g10101 ( new_n12450 , n26107 , new_n12449_1 );
not  g10102 ( new_n12451 , new_n12450 );
nor  g10103 ( new_n12452 , n22597 , new_n12451 );
not  g10104 ( new_n12453 , new_n12452 );
nor  g10105 ( new_n12454 , n19327 , new_n12453 );
not  g10106 ( new_n12455 , new_n12454 );
nor  g10107 ( new_n12456 , n26224 , new_n12455 );
and  g10108 ( new_n12457 , new_n11636 , new_n12456 );
and  g10109 ( new_n12458 , new_n12443 , new_n12457 );
xnor g10110 ( new_n12459 , new_n12443 , new_n12457 );
nor  g10111 ( new_n12460 , n5704 , n18409 );
not  g10112 ( new_n12461_1 , new_n12460 );
nor  g10113 ( new_n12462_1 , n13708 , new_n12461_1 );
not  g10114 ( new_n12463 , new_n12462_1 );
nor  g10115 ( new_n12464 , n19911 , new_n12463 );
not  g10116 ( new_n12465 , new_n12464 );
nor  g10117 ( new_n12466 , n2731 , new_n12465 );
not  g10118 ( new_n12467_1 , new_n12466 );
nor  g10119 ( new_n12468 , n18907 , new_n12467_1 );
not  g10120 ( new_n12469_1 , new_n12468 );
nor  g10121 ( new_n12470 , n22332 , new_n12469_1 );
not  g10122 ( new_n12471 , new_n12470 );
nor  g10123 ( new_n12472 , n4256 , new_n12471 );
xnor g10124 ( new_n12473 , n21287 , new_n12472 );
nor  g10125 ( new_n12474 , n12861 , new_n12473 );
xnor g10126 ( new_n12475 , new_n7043 , new_n12473 );
xnor g10127 ( new_n12476 , n4256 , new_n12470 );
nor  g10128 ( new_n12477 , n13333 , new_n12476 );
xnor g10129 ( new_n12478 , new_n7046 , new_n12476 );
xnor g10130 ( new_n12479 , n22332 , new_n12468 );
nor  g10131 ( new_n12480 , n2210 , new_n12479 );
xnor g10132 ( new_n12481 , new_n7049 , new_n12479 );
xnor g10133 ( new_n12482 , n18907 , new_n12466 );
nor  g10134 ( new_n12483 , n20604 , new_n12482 );
xnor g10135 ( new_n12484 , new_n5125 , new_n12482 );
xnor g10136 ( new_n12485 , n2731 , new_n12464 );
nor  g10137 ( new_n12486 , n16158 , new_n12485 );
xnor g10138 ( new_n12487 , new_n4614 , new_n12485 );
xnor g10139 ( new_n12488 , n19911 , new_n12462_1 );
nor  g10140 ( new_n12489 , n5752 , new_n12488 );
xnor g10141 ( new_n12490 , n13708 , new_n12460 );
nor  g10142 ( new_n12491 , n18171 , new_n12490 );
xnor g10143 ( new_n12492 , new_n4620 , new_n12490 );
xnor g10144 ( new_n12493 , n5704 , n18409 );
and  g10145 ( new_n12494 , new_n4623 , new_n12493 );
or   g10146 ( new_n12495_1 , new_n2381 , new_n4626 );
xnor g10147 ( new_n12496 , n25073 , new_n12493 );
and  g10148 ( new_n12497 , new_n12495_1 , new_n12496 );
or   g10149 ( new_n12498 , new_n12494 , new_n12497 );
and  g10150 ( new_n12499 , new_n12492 , new_n12498 );
or   g10151 ( new_n12500 , new_n12491 , new_n12499 );
xnor g10152 ( new_n12501 , new_n4617 , new_n12488 );
and  g10153 ( new_n12502 , new_n12500 , new_n12501 );
or   g10154 ( new_n12503 , new_n12489 , new_n12502 );
and  g10155 ( new_n12504 , new_n12487 , new_n12503 );
or   g10156 ( new_n12505 , new_n12486 , new_n12504 );
and  g10157 ( new_n12506 , new_n12484 , new_n12505 );
or   g10158 ( new_n12507_1 , new_n12483 , new_n12506 );
and  g10159 ( new_n12508 , new_n12481 , new_n12507_1 );
or   g10160 ( new_n12509 , new_n12480 , new_n12508 );
and  g10161 ( new_n12510 , new_n12478 , new_n12509 );
or   g10162 ( new_n12511 , new_n12477 , new_n12510 );
and  g10163 ( new_n12512 , new_n12475 , new_n12511 );
nor  g10164 ( new_n12513 , new_n12474 , new_n12512 );
not  g10165 ( new_n12514 , new_n12472 );
nor  g10166 ( new_n12515_1 , n21287 , new_n12514 );
xnor g10167 ( new_n12516_1 , n26986 , new_n12515_1 );
xnor g10168 ( new_n12517 , new_n7110 , new_n12516_1 );
xnor g10169 ( new_n12518 , new_n12513 , new_n12517 );
nor  g10170 ( new_n12519 , new_n12459 , new_n12518 );
xnor g10171 ( new_n12520 , new_n12459 , new_n12518 );
xnor g10172 ( new_n12521 , new_n11636 , new_n12456 );
nor  g10173 ( new_n12522 , new_n12477 , new_n12510 );
xnor g10174 ( new_n12523 , new_n12475 , new_n12522 );
nor  g10175 ( new_n12524 , new_n12521 , new_n12523 );
xnor g10176 ( new_n12525 , new_n12521 , new_n12523 );
not  g10177 ( new_n12526 , n26224 );
xnor g10178 ( new_n12527 , new_n12526 , new_n12454 );
xor  g10179 ( new_n12528 , new_n12478 , new_n12509 );
nor  g10180 ( new_n12529 , new_n12527 , new_n12528 );
xnor g10181 ( new_n12530 , new_n12527 , new_n12528 );
xnor g10182 ( new_n12531 , new_n3726 , new_n12452 );
nor  g10183 ( new_n12532 , new_n12483 , new_n12506 );
xnor g10184 ( new_n12533 , new_n12481 , new_n12532 );
nor  g10185 ( new_n12534 , new_n12531 , new_n12533 );
xnor g10186 ( new_n12535 , new_n12531 , new_n12533 );
xnor g10187 ( new_n12536 , new_n3740_1 , new_n12450 );
xor  g10188 ( new_n12537 , new_n12484 , new_n12505 );
nor  g10189 ( new_n12538 , new_n12536 , new_n12537 );
xnor g10190 ( new_n12539 , new_n12536 , new_n12537 );
xnor g10191 ( new_n12540_1 , n26107 , new_n12448 );
not  g10192 ( new_n12541 , new_n12540_1 );
nor  g10193 ( new_n12542 , new_n12489 , new_n12502 );
xnor g10194 ( new_n12543 , new_n12487 , new_n12542 );
nor  g10195 ( new_n12544 , new_n12541 , new_n12543 );
not  g10196 ( new_n12545_1 , new_n12543 );
xnor g10197 ( new_n12546_1 , new_n12541 , new_n12545_1 );
xnor g10198 ( new_n12547 , n342 , new_n12446_1 );
xnor g10199 ( new_n12548 , new_n12500 , new_n12501 );
and  g10200 ( new_n12549 , new_n12547 , new_n12548 );
xor  g10201 ( new_n12550 , new_n12500 , new_n12501 );
xnor g10202 ( new_n12551 , new_n12547 , new_n12550 );
nor  g10203 ( new_n12552_1 , new_n12494 , new_n12497 );
xnor g10204 ( new_n12553 , new_n12492 , new_n12552_1 );
not  g10205 ( new_n12554 , new_n12553 );
xnor g10206 ( new_n12555 , n26553 , new_n12444 );
and  g10207 ( new_n12556 , new_n12554 , new_n12555 );
xnor g10208 ( new_n12557 , new_n12553 , new_n12555 );
xnor g10209 ( new_n12558 , n4964 , n7876 );
nor  g10210 ( new_n12559 , new_n2381 , new_n4626 );
xnor g10211 ( new_n12560 , new_n12559 , new_n12496 );
nor  g10212 ( new_n12561 , new_n12558 , new_n12560 );
xnor g10213 ( new_n12562_1 , new_n2381 , n22309 );
not  g10214 ( new_n12563 , new_n12562_1 );
nor  g10215 ( new_n12564 , new_n3755_1 , new_n12563 );
not  g10216 ( new_n12565 , new_n12560 );
xnor g10217 ( new_n12566_1 , new_n12558 , new_n12565 );
and  g10218 ( new_n12567 , new_n12564 , new_n12566_1 );
or   g10219 ( new_n12568 , new_n12561 , new_n12567 );
and  g10220 ( new_n12569_1 , new_n12557 , new_n12568 );
or   g10221 ( new_n12570 , new_n12556 , new_n12569_1 );
and  g10222 ( new_n12571 , new_n12551 , new_n12570 );
or   g10223 ( new_n12572 , new_n12549 , new_n12571 );
and  g10224 ( new_n12573 , new_n12546_1 , new_n12572 );
nor  g10225 ( new_n12574 , new_n12544 , new_n12573 );
nor  g10226 ( new_n12575 , new_n12539 , new_n12574 );
nor  g10227 ( new_n12576 , new_n12538 , new_n12575 );
nor  g10228 ( new_n12577 , new_n12535 , new_n12576 );
nor  g10229 ( new_n12578 , new_n12534 , new_n12577 );
nor  g10230 ( new_n12579 , new_n12530 , new_n12578 );
nor  g10231 ( new_n12580 , new_n12529 , new_n12579 );
nor  g10232 ( new_n12581 , new_n12525 , new_n12580 );
nor  g10233 ( new_n12582 , new_n12524 , new_n12581 );
nor  g10234 ( new_n12583 , new_n12520 , new_n12582 );
or   g10235 ( new_n12584 , new_n12519 , new_n12583 );
nor  g10236 ( new_n12585 , new_n12458 , new_n12584 );
and  g10237 ( new_n12586 , new_n7243 , new_n12515_1 );
nor  g10238 ( new_n12587_1 , n8305 , new_n12516_1 );
and  g10239 ( new_n12588 , n8305 , new_n12516_1 );
nor  g10240 ( new_n12589 , new_n12513 , new_n12588 );
nor  g10241 ( new_n12590 , new_n12587_1 , new_n12589 );
or   g10242 ( new_n12591 , new_n12586 , new_n12590 );
and  g10243 ( new_n12592 , new_n12585 , new_n12591 );
xnor g10244 ( new_n12593_1 , new_n12442 , new_n12592 );
xnor g10245 ( new_n12594 , new_n12438 , new_n12441 );
nor  g10246 ( new_n12595 , new_n12586 , new_n12590 );
xnor g10247 ( new_n12596 , new_n12585 , new_n12595 );
not  g10248 ( new_n12597 , new_n12596 );
nor  g10249 ( new_n12598 , new_n12594 , new_n12597 );
xnor g10250 ( new_n12599 , new_n12594 , new_n12597 );
xnor g10251 ( new_n12600 , new_n12393 , new_n12436 );
xnor g10252 ( new_n12601 , new_n12520 , new_n12582 );
not  g10253 ( new_n12602 , new_n12601 );
nor  g10254 ( new_n12603 , new_n12600 , new_n12602 );
xnor g10255 ( new_n12604 , new_n12600 , new_n12602 );
xnor g10256 ( new_n12605 , new_n12396 , new_n12434 );
xnor g10257 ( new_n12606 , new_n12525 , new_n12580 );
not  g10258 ( new_n12607_1 , new_n12606 );
nor  g10259 ( new_n12608 , new_n12605 , new_n12607_1 );
xnor g10260 ( new_n12609 , new_n12605 , new_n12607_1 );
xnor g10261 ( new_n12610 , new_n12399 , new_n12432 );
xnor g10262 ( new_n12611 , new_n12530 , new_n12578 );
not  g10263 ( new_n12612 , new_n12611 );
nor  g10264 ( new_n12613 , new_n12610 , new_n12612 );
xnor g10265 ( new_n12614 , new_n12610 , new_n12612 );
xnor g10266 ( new_n12615 , new_n12402 , new_n12430 );
xnor g10267 ( new_n12616 , new_n12535 , new_n12576 );
not  g10268 ( new_n12617 , new_n12616 );
nor  g10269 ( new_n12618 , new_n12615 , new_n12617 );
xnor g10270 ( new_n12619 , new_n12615 , new_n12617 );
xnor g10271 ( new_n12620_1 , new_n12405 , new_n12428 );
xnor g10272 ( new_n12621_1 , new_n12539 , new_n12574 );
not  g10273 ( new_n12622 , new_n12621_1 );
nor  g10274 ( new_n12623 , new_n12620_1 , new_n12622 );
xnor g10275 ( new_n12624 , new_n12620_1 , new_n12622 );
xnor g10276 ( new_n12625 , new_n12408_1 , new_n12426 );
xor  g10277 ( new_n12626_1 , new_n12546_1 , new_n12572 );
nor  g10278 ( new_n12627 , new_n12625 , new_n12626_1 );
xnor g10279 ( new_n12628 , new_n12625 , new_n12626_1 );
xnor g10280 ( new_n12629 , new_n12411 , new_n12424 );
xor  g10281 ( new_n12630 , new_n12551 , new_n12570 );
nor  g10282 ( new_n12631 , new_n12629 , new_n12630 );
xnor g10283 ( new_n12632 , new_n12629 , new_n12630 );
xnor g10284 ( new_n12633 , new_n12414 , new_n12422 );
nor  g10285 ( new_n12634 , new_n12561 , new_n12567 );
xnor g10286 ( new_n12635 , new_n12557 , new_n12634 );
nor  g10287 ( new_n12636 , new_n12633 , new_n12635 );
not  g10288 ( new_n12637 , new_n12635 );
xnor g10289 ( new_n12638 , new_n12633 , new_n12637 );
xnor g10290 ( new_n12639 , new_n12564 , new_n12566_1 );
xnor g10291 ( new_n12640 , new_n12418 , new_n12419 );
not  g10292 ( new_n12641 , new_n12640 );
nor  g10293 ( new_n12642 , new_n12639 , new_n12641 );
xnor g10294 ( new_n12643 , n11479 , new_n12415 );
xnor g10295 ( new_n12644 , n7876 , new_n12563 );
not  g10296 ( new_n12645 , new_n12644 );
nor  g10297 ( new_n12646 , new_n12643 , new_n12645 );
xnor g10298 ( new_n12647 , new_n12639 , new_n12640 );
and  g10299 ( new_n12648 , new_n12646 , new_n12647 );
nor  g10300 ( new_n12649 , new_n12642 , new_n12648 );
and  g10301 ( new_n12650_1 , new_n12638 , new_n12649 );
nor  g10302 ( new_n12651 , new_n12636 , new_n12650_1 );
nor  g10303 ( new_n12652 , new_n12632 , new_n12651 );
nor  g10304 ( new_n12653 , new_n12631 , new_n12652 );
nor  g10305 ( new_n12654_1 , new_n12628 , new_n12653 );
nor  g10306 ( new_n12655 , new_n12627 , new_n12654_1 );
nor  g10307 ( new_n12656 , new_n12624 , new_n12655 );
nor  g10308 ( new_n12657_1 , new_n12623 , new_n12656 );
nor  g10309 ( new_n12658 , new_n12619 , new_n12657_1 );
nor  g10310 ( new_n12659 , new_n12618 , new_n12658 );
nor  g10311 ( new_n12660 , new_n12614 , new_n12659 );
nor  g10312 ( new_n12661 , new_n12613 , new_n12660 );
nor  g10313 ( new_n12662 , new_n12609 , new_n12661 );
nor  g10314 ( new_n12663 , new_n12608 , new_n12662 );
nor  g10315 ( new_n12664 , new_n12604 , new_n12663 );
nor  g10316 ( new_n12665_1 , new_n12603 , new_n12664 );
nor  g10317 ( new_n12666 , new_n12599 , new_n12665_1 );
nor  g10318 ( new_n12667 , new_n12598 , new_n12666 );
xnor g10319 ( n2095 , new_n12593_1 , new_n12667 );
xnor g10320 ( n2105 , new_n11258 , new_n11259 );
not  g10321 ( new_n12670_1 , new_n6088 );
not  g10322 ( new_n12671 , n11898 );
xnor g10323 ( new_n12672 , new_n12671 , n23166 );
not  g10324 ( new_n12673 , n19941 );
nor  g10325 ( new_n12674 , new_n9079 , new_n12673 );
or   g10326 ( new_n12675 , n10577 , n19941 );
nor  g10327 ( new_n12676 , n1099 , n6381 );
nor  g10328 ( new_n12677 , new_n10432_1 , new_n10449 );
nor  g10329 ( new_n12678 , new_n12676 , new_n12677 );
and  g10330 ( new_n12679 , new_n12675 , new_n12678 );
nor  g10331 ( new_n12680 , new_n12674 , new_n12679 );
xor  g10332 ( new_n12681 , new_n12672 , new_n12680 );
xnor g10333 ( new_n12682 , n8827 , new_n12681 );
not  g10334 ( new_n12683 , n18035 );
xnor g10335 ( new_n12684 , new_n9079 , n19941 );
xnor g10336 ( new_n12685 , new_n12678 , new_n12684 );
nor  g10337 ( new_n12686 , new_n12683 , new_n12685 );
not  g10338 ( new_n12687 , new_n12685 );
xnor g10339 ( new_n12688 , new_n12683 , new_n12687 );
nor  g10340 ( new_n12689 , n5077 , new_n10450 );
and  g10341 ( new_n12690 , new_n10451 , new_n10476 );
nor  g10342 ( new_n12691 , new_n12689 , new_n12690 );
and  g10343 ( new_n12692 , new_n12688 , new_n12691 );
or   g10344 ( new_n12693 , new_n12686 , new_n12692 );
xor  g10345 ( new_n12694 , new_n12682 , new_n12693 );
xnor g10346 ( new_n12695 , new_n12670_1 , new_n12694 );
xnor g10347 ( new_n12696 , new_n12688 , new_n12691 );
nor  g10348 ( new_n12697 , new_n6091 , new_n12696 );
not  g10349 ( new_n12698 , new_n6091 );
not  g10350 ( new_n12699 , new_n12696 );
xnor g10351 ( new_n12700 , new_n12698 , new_n12699 );
nor  g10352 ( new_n12701 , new_n6097 , new_n10477 );
xnor g10353 ( new_n12702_1 , new_n6097 , new_n10477 );
nor  g10354 ( new_n12703 , new_n6102 , new_n10480 );
not  g10355 ( new_n12704 , new_n6102 );
xnor g10356 ( new_n12705 , new_n12704 , new_n10481 );
nor  g10357 ( new_n12706 , new_n6107 , new_n10485 );
xnor g10358 ( new_n12707_1 , new_n6107 , new_n10485 );
nor  g10359 ( new_n12708 , new_n6112 , new_n10491 );
xnor g10360 ( new_n12709 , new_n6112 , new_n10491 );
nor  g10361 ( new_n12710 , new_n6116 , new_n8474 );
xnor g10362 ( new_n12711 , new_n6116 , new_n8474 );
nor  g10363 ( new_n12712 , new_n6122 , new_n8452 );
xnor g10364 ( new_n12713 , new_n6122 , new_n8452 );
nor  g10365 ( new_n12714 , new_n6132 , new_n8455 );
nor  g10366 ( new_n12715 , new_n5793 , new_n8459 );
xnor g10367 ( new_n12716 , new_n6126 , new_n8455 );
and  g10368 ( new_n12717 , new_n12715 , new_n12716 );
nor  g10369 ( new_n12718 , new_n12714 , new_n12717 );
nor  g10370 ( new_n12719 , new_n12713 , new_n12718 );
nor  g10371 ( new_n12720 , new_n12712 , new_n12719 );
nor  g10372 ( new_n12721 , new_n12711 , new_n12720 );
nor  g10373 ( new_n12722 , new_n12710 , new_n12721 );
nor  g10374 ( new_n12723 , new_n12709 , new_n12722 );
nor  g10375 ( new_n12724 , new_n12708 , new_n12723 );
nor  g10376 ( new_n12725_1 , new_n12707_1 , new_n12724 );
nor  g10377 ( new_n12726 , new_n12706 , new_n12725_1 );
nor  g10378 ( new_n12727_1 , new_n12705 , new_n12726 );
nor  g10379 ( new_n12728 , new_n12703 , new_n12727_1 );
nor  g10380 ( new_n12729 , new_n12702_1 , new_n12728 );
nor  g10381 ( new_n12730 , new_n12701 , new_n12729 );
nor  g10382 ( new_n12731 , new_n12700 , new_n12730 );
nor  g10383 ( new_n12732 , new_n12697 , new_n12731 );
xnor g10384 ( n2122 , new_n12695 , new_n12732 );
xnor g10385 ( n2147 , new_n2809_1 , new_n2837 );
xnor g10386 ( n2209 , new_n10365 , new_n10400 );
xnor g10387 ( n2214 , new_n5663 , new_n5771 );
xnor g10388 ( new_n12737 , new_n4195 , new_n11051 );
nor  g10389 ( new_n12738 , new_n4285 , new_n11053 );
xnor g10390 ( new_n12739 , new_n4285 , new_n11055 );
nor  g10391 ( new_n12740_1 , new_n4293 , new_n11069 );
xnor g10392 ( new_n12741 , new_n4293 , new_n11058 );
and  g10393 ( new_n12742_1 , new_n4299 , new_n11064 );
nor  g10394 ( new_n12743 , new_n4301 , new_n11061 );
xnor g10395 ( new_n12744 , new_n4299 , new_n11064 );
nor  g10396 ( new_n12745 , new_n12743 , new_n12744 );
nor  g10397 ( new_n12746_1 , new_n12742_1 , new_n12745 );
and  g10398 ( new_n12747 , new_n12741 , new_n12746_1 );
nor  g10399 ( new_n12748 , new_n12740_1 , new_n12747 );
and  g10400 ( new_n12749 , new_n12739 , new_n12748 );
nor  g10401 ( new_n12750 , new_n12738 , new_n12749 );
xnor g10402 ( n2238 , new_n12737 , new_n12750 );
xor  g10403 ( n2327 , new_n11074 , new_n11075 );
xnor g10404 ( n2343 , new_n5724 , new_n5755 );
not  g10405 ( new_n12754 , n13453 );
xnor g10406 ( new_n12755 , new_n12754 , new_n10464 );
nor  g10407 ( new_n12756_1 , new_n6589 , new_n6603 );
and  g10408 ( new_n12757 , new_n6605 , new_n6621 );
nor  g10409 ( new_n12758 , new_n12756_1 , new_n12757 );
xnor g10410 ( new_n12759 , new_n12755 , new_n12758 );
xnor g10411 ( new_n12760 , n16524 , n20923 );
nor  g10412 ( new_n12761 , n11056 , n18157 );
nor  g10413 ( new_n12762 , new_n6624 , new_n6635 );
nor  g10414 ( new_n12763 , new_n12761 , new_n12762 );
xnor g10415 ( new_n12764 , new_n12760 , new_n12763 );
xnor g10416 ( new_n12765 , n3785 , new_n12764 );
nor  g10417 ( new_n12766 , n20250 , new_n6636 );
nor  g10418 ( new_n12767 , new_n6637 , new_n6650 );
nor  g10419 ( new_n12768 , new_n12766 , new_n12767 );
xnor g10420 ( new_n12769 , new_n12765 , new_n12768 );
not  g10421 ( new_n12770 , new_n12769 );
xnor g10422 ( new_n12771 , new_n12759 , new_n12770 );
nor  g10423 ( new_n12772 , new_n6623 , new_n6651 );
and  g10424 ( new_n12773 , new_n6653 , new_n6673_1 );
nor  g10425 ( new_n12774 , new_n12772 , new_n12773 );
xnor g10426 ( n2361 , new_n12771 , new_n12774 );
xnor g10427 ( n2363 , new_n8367 , new_n3705 );
xnor g10428 ( n2374 , new_n4566 , new_n4598 );
xnor g10429 ( new_n12778 , n1204 , n7305 );
nor  g10430 ( new_n12779 , n19618 , n25872 );
and  g10431 ( new_n12780 , new_n5825 , new_n5830 );
nor  g10432 ( new_n12781 , new_n12779 , new_n12780 );
xnor g10433 ( new_n12782 , new_n12778 , new_n12781 );
nor  g10434 ( new_n12783_1 , new_n4864 , new_n12782 );
xor  g10435 ( new_n12784 , new_n4864 , new_n12782 );
nor  g10436 ( new_n12785 , new_n4880 , new_n5831 );
nor  g10437 ( new_n12786 , new_n5832 , new_n5841_1 );
nor  g10438 ( new_n12787 , new_n12785 , new_n12786 );
and  g10439 ( new_n12788 , new_n12784 , new_n12787 );
nor  g10440 ( new_n12789 , new_n12783_1 , new_n12788 );
xnor g10441 ( new_n12790 , new_n4223 , n20826 );
nor  g10442 ( new_n12791 , n1204 , n7305 );
nor  g10443 ( new_n12792 , new_n12778 , new_n12781 );
or   g10444 ( new_n12793 , new_n12791 , new_n12792 );
xor  g10445 ( new_n12794 , new_n12790 , new_n12793 );
not  g10446 ( new_n12795 , new_n12794 );
xnor g10447 ( new_n12796 , new_n12789 , new_n12795 );
xnor g10448 ( new_n12797 , new_n4859 , new_n12796 );
xnor g10449 ( new_n12798 , new_n3780 , new_n12797 );
xor  g10450 ( new_n12799 , new_n12784 , new_n12787 );
nor  g10451 ( new_n12800 , new_n3785_1 , new_n12799 );
nor  g10452 ( new_n12801_1 , new_n3790 , new_n5842_1 );
and  g10453 ( new_n12802 , new_n5843 , new_n5851 );
nor  g10454 ( new_n12803 , new_n12801_1 , new_n12802 );
xnor g10455 ( new_n12804 , new_n3785_1 , new_n12799 );
nor  g10456 ( new_n12805 , new_n12803 , new_n12804 );
or   g10457 ( new_n12806 , new_n12800 , new_n12805 );
xor  g10458 ( n2388 , new_n12798 , new_n12806 );
not  g10459 ( new_n12808 , n2160 );
xnor g10460 ( new_n12809 , new_n12808 , n7335 );
nor  g10461 ( new_n12810 , n5696 , n10763 );
and  g10462 ( new_n12811_1 , new_n5305 , new_n5334 );
or   g10463 ( new_n12812_1 , new_n12810 , new_n12811_1 );
xor  g10464 ( new_n12813 , new_n12809 , new_n12812_1 );
xnor g10465 ( new_n12814 , n3425 , n11220 );
nor  g10466 ( new_n12815 , n9967 , n22379 );
nor  g10467 ( new_n12816_1 , new_n5271 , new_n5303 );
nor  g10468 ( new_n12817 , new_n12815 , new_n12816_1 );
xnor g10469 ( new_n12818 , new_n12814 , new_n12817 );
xnor g10470 ( new_n12819 , new_n12813 , new_n12818 );
nor  g10471 ( new_n12820 , new_n5304 , new_n5335 );
nor  g10472 ( new_n12821_1 , new_n5336 , new_n5398 );
nor  g10473 ( new_n12822 , new_n12820 , new_n12821_1 );
xnor g10474 ( new_n12823 , new_n12819 , new_n12822 );
not  g10475 ( new_n12824 , new_n12823 );
not  g10476 ( new_n12825 , new_n5231 );
nor  g10477 ( new_n12826 , n337 , new_n12825 );
xnor g10478 ( new_n12827 , n7593 , new_n12826 );
xnor g10479 ( new_n12828 , new_n3086 , new_n12827 );
nor  g10480 ( new_n12829 , n6485 , new_n5232 );
and  g10481 ( new_n12830 , new_n5233 , new_n5269 );
nor  g10482 ( new_n12831 , new_n12829 , new_n12830 );
xnor g10483 ( new_n12832 , new_n12828 , new_n12831 );
xnor g10484 ( new_n12833 , new_n12824 , new_n12832 );
nor  g10485 ( new_n12834 , new_n5270 , new_n5399_1 );
and  g10486 ( new_n12835 , new_n5401 , new_n5451_1 );
or   g10487 ( new_n12836 , new_n12834 , new_n12835 );
xor  g10488 ( n2440 , new_n12833 , new_n12836 );
xnor g10489 ( n2444 , new_n11394 , new_n11407 );
xnor g10490 ( n2513 , new_n3257 , new_n5083 );
xnor g10491 ( new_n12840 , n14323 , new_n5943_1 );
not  g10492 ( new_n12841 , n2886 );
nor  g10493 ( new_n12842 , new_n12841 , new_n5950 );
xnor g10494 ( new_n12843_1 , n2886 , new_n5950 );
nor  g10495 ( new_n12844 , new_n12373 , new_n5961 );
nor  g10496 ( new_n12845 , new_n12371 , new_n3798 );
xnor g10497 ( new_n12846 , n1040 , new_n5961 );
and  g10498 ( new_n12847 , new_n12845 , new_n12846 );
or   g10499 ( new_n12848 , new_n12844 , new_n12847 );
and  g10500 ( new_n12849 , new_n12843_1 , new_n12848 );
nor  g10501 ( new_n12850 , new_n12842 , new_n12849 );
xnor g10502 ( new_n12851 , new_n12840 , new_n12850 );
xnor g10503 ( new_n12852 , n12562 , new_n12851 );
xor  g10504 ( new_n12853 , new_n12843_1 , new_n12848 );
nor  g10505 ( new_n12854 , n7949 , new_n12853 );
xnor g10506 ( new_n12855 , new_n5892 , new_n12853 );
nor  g10507 ( new_n12856 , new_n5895 , new_n10778 );
nor  g10508 ( new_n12857 , n24374 , new_n12856 );
xnor g10509 ( new_n12858 , new_n12845 , new_n12846 );
xor  g10510 ( new_n12859 , n24374 , new_n12856 );
and  g10511 ( new_n12860 , new_n12858 , new_n12859 );
or   g10512 ( new_n12861_1 , new_n12857 , new_n12860 );
and  g10513 ( new_n12862 , new_n12855 , new_n12861_1 );
nor  g10514 ( new_n12863 , new_n12854 , new_n12862 );
xor  g10515 ( new_n12864_1 , new_n12852 , new_n12863 );
xnor g10516 ( new_n12865_1 , new_n12630 , new_n12864_1 );
xor  g10517 ( new_n12866 , new_n12855 , new_n12861_1 );
and  g10518 ( new_n12867 , new_n12637 , new_n12866 );
xnor g10519 ( new_n12868 , new_n12637 , new_n12866 );
not  g10520 ( new_n12869 , new_n12858 );
xnor g10521 ( new_n12870_1 , new_n12869 , new_n12859 );
and  g10522 ( new_n12871_1 , new_n12639 , new_n12870_1 );
xnor g10523 ( new_n12872 , n14575 , new_n10778 );
and  g10524 ( new_n12873_1 , new_n12644 , new_n12872 );
xnor g10525 ( new_n12874 , new_n12639 , new_n12870_1 );
nor  g10526 ( new_n12875_1 , new_n12873_1 , new_n12874 );
nor  g10527 ( new_n12876 , new_n12871_1 , new_n12875_1 );
nor  g10528 ( new_n12877 , new_n12868 , new_n12876 );
nor  g10529 ( new_n12878 , new_n12867 , new_n12877 );
xnor g10530 ( n2515 , new_n12865_1 , new_n12878 );
xnor g10531 ( n2533 , new_n10741 , new_n10769 );
nor  g10532 ( new_n12881 , new_n3217 , n26986 );
xnor g10533 ( new_n12882 , n3425 , n26986 );
nor  g10534 ( new_n12883 , new_n3198 , n21287 );
xnor g10535 ( new_n12884 , n9967 , n21287 );
nor  g10536 ( new_n12885 , n4256 , new_n7508 );
xnor g10537 ( new_n12886 , n4256 , n20946 );
nor  g10538 ( new_n12887 , new_n5275 , n22332 );
xnor g10539 ( new_n12888 , n7751 , n22332 );
not  g10540 ( new_n12889 , n26823 );
nor  g10541 ( new_n12890 , n18907 , new_n12889 );
xnor g10542 ( new_n12891 , n18907 , n26823 );
nor  g10543 ( new_n12892_1 , n2731 , new_n5280 );
and  g10544 ( new_n12893 , new_n8393 , new_n8409 );
or   g10545 ( new_n12894 , new_n12892_1 , new_n12893 );
and  g10546 ( new_n12895 , new_n12891 , new_n12894 );
or   g10547 ( new_n12896 , new_n12890 , new_n12895 );
and  g10548 ( new_n12897 , new_n12888 , new_n12896 );
or   g10549 ( new_n12898 , new_n12887 , new_n12897 );
and  g10550 ( new_n12899 , new_n12886 , new_n12898 );
or   g10551 ( new_n12900_1 , new_n12885 , new_n12899 );
and  g10552 ( new_n12901 , new_n12884 , new_n12900_1 );
or   g10553 ( new_n12902 , new_n12883 , new_n12901 );
and  g10554 ( new_n12903 , new_n12882 , new_n12902 );
nor  g10555 ( new_n12904_1 , new_n12881 , new_n12903 );
not  g10556 ( new_n12905 , new_n7059 );
not  g10557 ( new_n12906 , new_n7064 );
not  g10558 ( new_n12907 , new_n5124 );
nor  g10559 ( new_n12908 , new_n12907 , new_n5132 );
not  g10560 ( new_n12909 , new_n12908 );
not  g10561 ( new_n12910 , new_n7068 );
nor  g10562 ( new_n12911 , new_n12909 , new_n12910 );
not  g10563 ( new_n12912 , new_n12911 );
nor  g10564 ( new_n12913 , new_n12906 , new_n12912 );
not  g10565 ( new_n12914 , new_n12913 );
nor  g10566 ( new_n12915 , new_n12905 , new_n12914 );
and  g10567 ( new_n12916 , new_n7116 , new_n12915 );
and  g10568 ( new_n12917_1 , new_n7186 , new_n12916 );
not  g10569 ( new_n12918 , new_n7189 );
nor  g10570 ( new_n12919 , new_n12918 , new_n12916 );
nor  g10571 ( new_n12920 , new_n12917_1 , new_n12919 );
nor  g10572 ( new_n12921 , new_n3195 , new_n12920 );
xor  g10573 ( new_n12922 , new_n7116 , new_n12915 );
nor  g10574 ( new_n12923 , new_n3137 , new_n12922 );
xnor g10575 ( new_n12924 , new_n3137 , new_n12922 );
xnor g10576 ( new_n12925 , new_n12905 , new_n12913 );
nor  g10577 ( new_n12926 , new_n3141 , new_n12925 );
xnor g10578 ( new_n12927 , new_n3141 , new_n12925 );
xnor g10579 ( new_n12928 , new_n12906 , new_n12911 );
nor  g10580 ( new_n12929 , new_n3145 , new_n12928 );
xnor g10581 ( new_n12930 , new_n3145 , new_n12928 );
xnor g10582 ( new_n12931 , new_n12908 , new_n12910 );
nor  g10583 ( new_n12932 , new_n3149 , new_n12931 );
xnor g10584 ( new_n12933 , new_n3149 , new_n12931 );
nor  g10585 ( new_n12934 , new_n3153 , new_n5133 );
nor  g10586 ( new_n12935 , new_n5134 , new_n5159 );
nor  g10587 ( new_n12936 , new_n12934 , new_n12935 );
nor  g10588 ( new_n12937 , new_n12933 , new_n12936 );
nor  g10589 ( new_n12938 , new_n12932 , new_n12937 );
nor  g10590 ( new_n12939 , new_n12930 , new_n12938 );
nor  g10591 ( new_n12940 , new_n12929 , new_n12939 );
nor  g10592 ( new_n12941_1 , new_n12927 , new_n12940 );
nor  g10593 ( new_n12942_1 , new_n12926 , new_n12941_1 );
nor  g10594 ( new_n12943 , new_n12924 , new_n12942_1 );
nor  g10595 ( new_n12944 , new_n12923 , new_n12943 );
and  g10596 ( new_n12945 , new_n3195 , new_n12920 );
nor  g10597 ( new_n12946 , new_n12944 , new_n12945 );
nor  g10598 ( new_n12947 , new_n12921 , new_n12946 );
nor  g10599 ( new_n12948 , new_n12917_1 , new_n12947 );
xnor g10600 ( new_n12949 , new_n12904_1 , new_n12948 );
xnor g10601 ( new_n12950 , new_n3196 , new_n12920 );
xnor g10602 ( new_n12951 , new_n12944 , new_n12950 );
not  g10603 ( new_n12952 , new_n12951 );
nor  g10604 ( new_n12953 , new_n12904_1 , new_n12952 );
xnor g10605 ( new_n12954 , new_n12904_1 , new_n12952 );
xor  g10606 ( new_n12955 , new_n12882 , new_n12902 );
xnor g10607 ( new_n12956_1 , new_n12924 , new_n12942_1 );
nor  g10608 ( new_n12957 , new_n12955 , new_n12956_1 );
xnor g10609 ( new_n12958 , new_n12955 , new_n12956_1 );
xor  g10610 ( new_n12959 , new_n12884 , new_n12900_1 );
xnor g10611 ( new_n12960 , new_n12927 , new_n12940 );
nor  g10612 ( new_n12961 , new_n12959 , new_n12960 );
xnor g10613 ( new_n12962 , new_n12959 , new_n12960 );
xor  g10614 ( new_n12963 , new_n12886 , new_n12898 );
xnor g10615 ( new_n12964 , new_n12930 , new_n12938 );
nor  g10616 ( new_n12965 , new_n12963 , new_n12964 );
xnor g10617 ( new_n12966 , new_n12963 , new_n12964 );
xor  g10618 ( new_n12967 , new_n12888 , new_n12896 );
xnor g10619 ( new_n12968 , new_n12933 , new_n12936 );
nor  g10620 ( new_n12969 , new_n12967 , new_n12968 );
not  g10621 ( new_n12970 , new_n12968 );
xnor g10622 ( new_n12971 , new_n12967 , new_n12970 );
xor  g10623 ( new_n12972 , new_n12891 , new_n12894 );
and  g10624 ( new_n12973 , new_n5160 , new_n12972 );
xnor g10625 ( new_n12974 , new_n5161 , new_n12972 );
and  g10626 ( new_n12975 , new_n5187 , new_n8410 );
and  g10627 ( new_n12976 , new_n8411 , new_n8430 );
or   g10628 ( new_n12977 , new_n12975 , new_n12976 );
and  g10629 ( new_n12978_1 , new_n12974 , new_n12977 );
nor  g10630 ( new_n12979 , new_n12973 , new_n12978_1 );
and  g10631 ( new_n12980_1 , new_n12971 , new_n12979 );
nor  g10632 ( new_n12981 , new_n12969 , new_n12980_1 );
nor  g10633 ( new_n12982 , new_n12966 , new_n12981 );
nor  g10634 ( new_n12983 , new_n12965 , new_n12982 );
nor  g10635 ( new_n12984 , new_n12962 , new_n12983 );
nor  g10636 ( new_n12985_1 , new_n12961 , new_n12984 );
nor  g10637 ( new_n12986 , new_n12958 , new_n12985_1 );
nor  g10638 ( new_n12987_1 , new_n12957 , new_n12986 );
nor  g10639 ( new_n12988 , new_n12954 , new_n12987_1 );
nor  g10640 ( new_n12989 , new_n12953 , new_n12988 );
xnor g10641 ( n2535 , new_n12949 , new_n12989 );
nor  g10642 ( new_n12991 , n3925 , n20259 );
not  g10643 ( new_n12992_1 , new_n12991 );
nor  g10644 ( new_n12993 , n25872 , new_n12992_1 );
not  g10645 ( new_n12994 , new_n12993 );
nor  g10646 ( new_n12995 , n7305 , new_n12994 );
not  g10647 ( new_n12996 , new_n12995 );
nor  g10648 ( new_n12997 , n20826 , new_n12996 );
xnor g10649 ( new_n12998 , n22198 , new_n12997 );
xnor g10650 ( new_n12999 , n21674 , new_n12998 );
xnor g10651 ( new_n13000 , n20826 , new_n12995 );
nor  g10652 ( new_n13001 , n17251 , new_n13000 );
xnor g10653 ( new_n13002 , n17251 , new_n13000 );
xnor g10654 ( new_n13003 , n7305 , new_n12993 );
nor  g10655 ( new_n13004 , n14790 , new_n13003 );
xnor g10656 ( new_n13005_1 , n25872 , new_n12991 );
nor  g10657 ( new_n13006 , n10096 , new_n13005_1 );
xnor g10658 ( new_n13007 , new_n3555_1 , new_n13005_1 );
xnor g10659 ( new_n13008 , n3925 , n20259 );
and  g10660 ( new_n13009 , new_n3558 , new_n13008 );
or   g10661 ( new_n13010 , new_n5002 , new_n3562 );
xnor g10662 ( new_n13011 , n16994 , new_n13008 );
and  g10663 ( new_n13012 , new_n13010 , new_n13011 );
or   g10664 ( new_n13013 , new_n13009 , new_n13012 );
and  g10665 ( new_n13014 , new_n13007 , new_n13013 );
nor  g10666 ( new_n13015 , new_n13006 , new_n13014 );
xnor g10667 ( new_n13016 , n14790 , new_n13003 );
nor  g10668 ( new_n13017 , new_n13015 , new_n13016 );
nor  g10669 ( new_n13018 , new_n13004 , new_n13017 );
nor  g10670 ( new_n13019 , new_n13002 , new_n13018 );
nor  g10671 ( new_n13020 , new_n13001 , new_n13019 );
xnor g10672 ( new_n13021 , new_n12999 , new_n13020 );
xnor g10673 ( new_n13022 , new_n7722 , new_n13021 );
xnor g10674 ( new_n13023 , new_n13002 , new_n13018 );
nor  g10675 ( new_n13024 , new_n7726 , new_n13023 );
xnor g10676 ( new_n13025 , new_n7726 , new_n13023 );
xnor g10677 ( new_n13026_1 , new_n13015 , new_n13016 );
nor  g10678 ( new_n13027 , new_n7731_1 , new_n13026_1 );
xor  g10679 ( new_n13028 , new_n7731_1 , new_n13026_1 );
xor  g10680 ( new_n13029 , new_n13007 , new_n13013 );
nor  g10681 ( new_n13030 , new_n7737 , new_n13029 );
xnor g10682 ( new_n13031 , new_n7737 , new_n13029 );
xor  g10683 ( new_n13032 , new_n13010 , new_n13011 );
nor  g10684 ( new_n13033 , new_n7745 , new_n13032 );
nor  g10685 ( new_n13034 , new_n7749 , new_n9707 );
xnor g10686 ( new_n13035 , new_n7746 , new_n13032 );
and  g10687 ( new_n13036 , new_n13034 , new_n13035 );
nor  g10688 ( new_n13037 , new_n13033 , new_n13036 );
nor  g10689 ( new_n13038 , new_n13031 , new_n13037 );
nor  g10690 ( new_n13039 , new_n13030 , new_n13038 );
and  g10691 ( new_n13040 , new_n13028 , new_n13039 );
nor  g10692 ( new_n13041 , new_n13027 , new_n13040 );
nor  g10693 ( new_n13042 , new_n13025 , new_n13041 );
nor  g10694 ( new_n13043_1 , new_n13024 , new_n13042 );
xnor g10695 ( new_n13044_1 , new_n13022 , new_n13043_1 );
xnor g10696 ( new_n13045 , n329 , n1163 );
not  g10697 ( new_n13046 , n24170 );
nor  g10698 ( new_n13047 , n18537 , new_n13046 );
xnor g10699 ( new_n13048_1 , n18537 , n24170 );
not  g10700 ( new_n13049 , n2409 );
nor  g10701 ( new_n13050 , new_n13049 , n7057 );
xnor g10702 ( new_n13051 , n2409 , n7057 );
nor  g10703 ( new_n13052 , new_n8510_1 , n8869 );
and  g10704 ( new_n13053 , new_n8510_1 , n8869 );
nor  g10705 ( new_n13054_1 , n10372 , new_n5040 );
nor  g10706 ( new_n13055 , n7428 , new_n5080 );
nand g10707 ( new_n13056 , n10372 , new_n5040 );
and  g10708 ( new_n13057 , new_n13055 , new_n13056 );
nor  g10709 ( new_n13058 , new_n13054_1 , new_n13057 );
nor  g10710 ( new_n13059 , new_n13053 , new_n13058 );
nor  g10711 ( new_n13060 , new_n13052 , new_n13059 );
and  g10712 ( new_n13061 , new_n13051 , new_n13060 );
or   g10713 ( new_n13062 , new_n13050 , new_n13061 );
and  g10714 ( new_n13063 , new_n13048_1 , new_n13062 );
or   g10715 ( new_n13064 , new_n13047 , new_n13063 );
xor  g10716 ( new_n13065 , new_n13045 , new_n13064 );
xnor g10717 ( new_n13066 , new_n13044_1 , new_n13065 );
xor  g10718 ( new_n13067 , new_n13048_1 , new_n13062 );
xnor g10719 ( new_n13068 , new_n13025 , new_n13041 );
nor  g10720 ( new_n13069 , new_n13067 , new_n13068 );
xnor g10721 ( new_n13070 , new_n13067 , new_n13068 );
xnor g10722 ( new_n13071 , new_n13028 , new_n13039 );
not  g10723 ( new_n13072 , new_n13071 );
xnor g10724 ( new_n13073 , new_n13051 , new_n13060 );
and  g10725 ( new_n13074_1 , new_n13072 , new_n13073 );
xnor g10726 ( new_n13075 , new_n13072 , new_n13073 );
xnor g10727 ( new_n13076 , new_n13031 , new_n13037 );
xnor g10728 ( new_n13077 , n8381 , n8869 );
xnor g10729 ( new_n13078 , new_n13058 , new_n13077 );
and  g10730 ( new_n13079 , new_n13076 , new_n13078 );
xnor g10731 ( new_n13080 , new_n13076 , new_n13078 );
nor  g10732 ( new_n13081 , new_n9708 , new_n9710 );
xnor g10733 ( new_n13082_1 , n10372 , n20235 );
xnor g10734 ( new_n13083 , new_n13055 , new_n13082_1 );
nor  g10735 ( new_n13084 , new_n13081 , new_n13083 );
xnor g10736 ( new_n13085 , new_n13034 , new_n13035 );
not  g10737 ( new_n13086 , new_n13085 );
xnor g10738 ( new_n13087 , new_n13081 , new_n13083 );
nor  g10739 ( new_n13088 , new_n13086 , new_n13087 );
nor  g10740 ( new_n13089 , new_n13084 , new_n13088 );
nor  g10741 ( new_n13090 , new_n13080 , new_n13089 );
nor  g10742 ( new_n13091 , new_n13079 , new_n13090 );
nor  g10743 ( new_n13092 , new_n13075 , new_n13091 );
nor  g10744 ( new_n13093 , new_n13074_1 , new_n13092 );
nor  g10745 ( new_n13094 , new_n13070 , new_n13093 );
nor  g10746 ( new_n13095 , new_n13069 , new_n13094 );
xnor g10747 ( n2537 , new_n13066 , new_n13095 );
not  g10748 ( new_n13097 , new_n2987 );
xnor g10749 ( new_n13098 , new_n13097 , new_n10936 );
nor  g10750 ( new_n13099 , new_n2994 , new_n4202 );
xnor g10751 ( new_n13100 , new_n2994 , new_n4201 );
nor  g10752 ( new_n13101 , new_n2998 , new_n4204_1 );
xnor g10753 ( new_n13102 , new_n3000 , new_n4204_1 );
nor  g10754 ( new_n13103 , new_n3004 , new_n4208 );
xnor g10755 ( new_n13104 , new_n3004 , new_n4207 );
and  g10756 ( new_n13105 , new_n3010_1 , new_n4211 );
nor  g10757 ( new_n13106 , n1152 , new_n3015 );
xnor g10758 ( new_n13107 , new_n3011 , new_n4211 );
and  g10759 ( new_n13108 , new_n13106 , new_n13107 );
nor  g10760 ( new_n13109 , new_n13105 , new_n13108 );
and  g10761 ( new_n13110_1 , new_n13104 , new_n13109 );
nor  g10762 ( new_n13111 , new_n13103 , new_n13110_1 );
and  g10763 ( new_n13112 , new_n13102 , new_n13111 );
nor  g10764 ( new_n13113 , new_n13101 , new_n13112 );
and  g10765 ( new_n13114 , new_n13100 , new_n13113 );
or   g10766 ( new_n13115 , new_n13099 , new_n13114 );
xor  g10767 ( new_n13116_1 , new_n13098 , new_n13115 );
xnor g10768 ( new_n13117 , new_n11357 , new_n13116_1 );
xor  g10769 ( new_n13118 , new_n13100 , new_n13113 );
nor  g10770 ( new_n13119 , new_n9517 , new_n13118 );
xnor g10771 ( new_n13120 , new_n9517 , new_n13118 );
xnor g10772 ( new_n13121 , new_n13102 , new_n13111 );
nor  g10773 ( new_n13122_1 , new_n9520 , new_n13121 );
xnor g10774 ( new_n13123 , new_n11875 , new_n13121 );
xnor g10775 ( new_n13124 , new_n13104 , new_n13109 );
nor  g10776 ( new_n13125 , new_n9528 , new_n13124 );
xnor g10777 ( new_n13126 , new_n9525 , new_n13124 );
xnor g10778 ( new_n13127 , new_n13106 , new_n13107 );
nor  g10779 ( new_n13128 , new_n9530 , new_n13127 );
xnor g10780 ( new_n13129 , new_n2698 , new_n3015 );
nor  g10781 ( new_n13130 , new_n7200 , new_n13129 );
xnor g10782 ( new_n13131 , new_n9530 , new_n13127 );
nor  g10783 ( new_n13132 , new_n13130 , new_n13131 );
nor  g10784 ( new_n13133 , new_n13128 , new_n13132 );
and  g10785 ( new_n13134 , new_n13126 , new_n13133 );
nor  g10786 ( new_n13135 , new_n13125 , new_n13134 );
and  g10787 ( new_n13136 , new_n13123 , new_n13135 );
nor  g10788 ( new_n13137_1 , new_n13122_1 , new_n13136 );
nor  g10789 ( new_n13138 , new_n13120 , new_n13137_1 );
nor  g10790 ( new_n13139 , new_n13119 , new_n13138 );
xnor g10791 ( n2553 , new_n13117 , new_n13139 );
xnor g10792 ( n2555 , new_n11761 , new_n11779 );
xnor g10793 ( new_n13142 , n12892 , new_n10607 );
not  g10794 ( new_n13143 , new_n13142 );
nor  g10795 ( new_n13144_1 , new_n9962 , new_n13143 );
not  g10796 ( new_n13145 , n12892 );
nor  g10797 ( new_n13146 , new_n13145 , new_n10607 );
not  g10798 ( new_n13147 , new_n10611_1 );
xnor g10799 ( new_n13148 , n12209 , new_n13147 );
xnor g10800 ( new_n13149 , new_n13146 , new_n13148 );
not  g10801 ( new_n13150 , new_n13149 );
xnor g10802 ( new_n13151 , new_n9965 , new_n13150 );
xnor g10803 ( n2560 , new_n13144_1 , new_n13151 );
nor  g10804 ( new_n13153 , n10650 , n26180 );
xnor g10805 ( new_n13154 , n10650 , n26180 );
nor  g10806 ( new_n13155 , n12900 , n24004 );
xnor g10807 ( new_n13156 , n12900 , n24004 );
nor  g10808 ( new_n13157 , n12871 , n20411 );
xnor g10809 ( new_n13158 , n12871 , n20411 );
nor  g10810 ( new_n13159 , n17069 , n23304 );
xnor g10811 ( new_n13160 , n17069 , n23304 );
nor  g10812 ( new_n13161 , n15918 , n19361 );
xnor g10813 ( new_n13162 , n15918 , n19361 );
nor  g10814 ( new_n13163 , n1437 , n17784 );
xnor g10815 ( new_n13164 , new_n3497 , n17784 );
nor  g10816 ( new_n13165 , n4722 , n14323 );
xnor g10817 ( new_n13166 , new_n3503 , n14323 );
nor  g10818 ( new_n13167 , n2886 , n14633 );
xnor g10819 ( new_n13168_1 , new_n12841 , n14633 );
nor  g10820 ( new_n13169 , n1040 , n8721 );
or   g10821 ( new_n13170 , new_n12371 , new_n3515 );
xnor g10822 ( new_n13171 , new_n12373 , n8721 );
and  g10823 ( new_n13172 , new_n13170 , new_n13171 );
or   g10824 ( new_n13173 , new_n13169 , new_n13172 );
and  g10825 ( new_n13174 , new_n13168_1 , new_n13173 );
or   g10826 ( new_n13175 , new_n13167 , new_n13174 );
and  g10827 ( new_n13176 , new_n13166 , new_n13175 );
or   g10828 ( new_n13177 , new_n13165 , new_n13176 );
and  g10829 ( new_n13178 , new_n13164 , new_n13177 );
nor  g10830 ( new_n13179 , new_n13163 , new_n13178 );
nor  g10831 ( new_n13180 , new_n13162 , new_n13179 );
nor  g10832 ( new_n13181 , new_n13161 , new_n13180 );
nor  g10833 ( new_n13182 , new_n13160 , new_n13181 );
nor  g10834 ( new_n13183 , new_n13159 , new_n13182 );
nor  g10835 ( new_n13184 , new_n13158 , new_n13183 );
nor  g10836 ( new_n13185 , new_n13157 , new_n13184 );
nor  g10837 ( new_n13186 , new_n13156 , new_n13185 );
nor  g10838 ( new_n13187 , new_n13155 , new_n13186 );
nor  g10839 ( new_n13188 , new_n13154 , new_n13187 );
nor  g10840 ( new_n13189 , new_n13153 , new_n13188 );
nor  g10841 ( new_n13190_1 , n6456 , n9259 );
or   g10842 ( new_n13191 , new_n5874 , new_n5912 );
and  g10843 ( new_n13192 , new_n5873 , new_n13191 );
nor  g10844 ( new_n13193 , new_n13190_1 , new_n13192 );
not  g10845 ( new_n13194 , new_n13193 );
nor  g10846 ( new_n13195 , new_n13189 , new_n13194 );
xnor g10847 ( new_n13196 , new_n13189 , new_n13194 );
xnor g10848 ( new_n13197 , new_n13154 , new_n13187 );
nor  g10849 ( new_n13198_1 , new_n5914 , new_n13197 );
xnor g10850 ( new_n13199_1 , new_n5914 , new_n13197 );
xnor g10851 ( new_n13200 , new_n13156 , new_n13185 );
nor  g10852 ( new_n13201 , new_n5919 , new_n13200 );
xnor g10853 ( new_n13202 , new_n5919 , new_n13200 );
xnor g10854 ( new_n13203 , new_n13158 , new_n13183 );
nor  g10855 ( new_n13204_1 , new_n5925 , new_n13203 );
xnor g10856 ( new_n13205 , new_n5925 , new_n13203 );
xnor g10857 ( new_n13206 , new_n13160 , new_n13181 );
nor  g10858 ( new_n13207 , new_n5930 , new_n13206 );
xnor g10859 ( new_n13208 , new_n5930 , new_n13206 );
xnor g10860 ( new_n13209_1 , new_n13162 , new_n13179 );
nor  g10861 ( new_n13210 , new_n5935 , new_n13209_1 );
not  g10862 ( new_n13211 , new_n5935 );
xnor g10863 ( new_n13212 , new_n13211 , new_n13209_1 );
not  g10864 ( new_n13213 , new_n5940 );
xor  g10865 ( new_n13214 , new_n13164 , new_n13177 );
nor  g10866 ( new_n13215 , new_n13213 , new_n13214 );
xnor g10867 ( new_n13216 , new_n13213 , new_n13214 );
nor  g10868 ( new_n13217 , new_n13167 , new_n13174 );
xnor g10869 ( new_n13218 , new_n13166 , new_n13217 );
nor  g10870 ( new_n13219 , new_n5947 , new_n13218 );
xnor g10871 ( new_n13220 , new_n5945 , new_n13218 );
nor  g10872 ( new_n13221 , new_n13169 , new_n13172 );
xnor g10873 ( new_n13222 , new_n13168_1 , new_n13221 );
nor  g10874 ( new_n13223 , new_n5953 , new_n13222 );
xnor g10875 ( new_n13224 , new_n5952 , new_n13222 );
xnor g10876 ( new_n13225 , new_n12371 , n18578 );
nor  g10877 ( new_n13226 , new_n5956 , new_n13225 );
nor  g10878 ( new_n13227 , new_n5959 , new_n13226 );
xnor g10879 ( new_n13228 , new_n13170 , new_n13171 );
not  g10880 ( new_n13229 , new_n13226 );
nor  g10881 ( new_n13230 , new_n5897 , new_n13229 );
nor  g10882 ( new_n13231 , new_n13227 , new_n13230 );
and  g10883 ( new_n13232 , new_n13228 , new_n13231 );
or   g10884 ( new_n13233 , new_n13227 , new_n13232 );
and  g10885 ( new_n13234 , new_n13224 , new_n13233 );
or   g10886 ( new_n13235 , new_n13223 , new_n13234 );
and  g10887 ( new_n13236 , new_n13220 , new_n13235 );
nor  g10888 ( new_n13237 , new_n13219 , new_n13236 );
nor  g10889 ( new_n13238 , new_n13216 , new_n13237 );
nor  g10890 ( new_n13239 , new_n13215 , new_n13238 );
and  g10891 ( new_n13240 , new_n13212 , new_n13239 );
nor  g10892 ( new_n13241 , new_n13210 , new_n13240 );
nor  g10893 ( new_n13242 , new_n13208 , new_n13241 );
nor  g10894 ( new_n13243 , new_n13207 , new_n13242 );
nor  g10895 ( new_n13244 , new_n13205 , new_n13243 );
nor  g10896 ( new_n13245 , new_n13204_1 , new_n13244 );
nor  g10897 ( new_n13246 , new_n13202 , new_n13245 );
nor  g10898 ( new_n13247 , new_n13201 , new_n13246 );
nor  g10899 ( new_n13248 , new_n13199_1 , new_n13247 );
nor  g10900 ( new_n13249 , new_n13198_1 , new_n13248 );
nor  g10901 ( new_n13250 , new_n13196 , new_n13249 );
nor  g10902 ( new_n13251 , new_n13195 , new_n13250 );
xnor g10903 ( new_n13252 , new_n13196 , new_n13249 );
not  g10904 ( new_n13253 , new_n13252 );
not  g10905 ( new_n13254 , n2743 );
nor  g10906 ( new_n13255 , new_n13254 , n3506 );
and  g10907 ( new_n13256 , new_n3536 , new_n3580 );
nor  g10908 ( new_n13257 , new_n13255 , new_n13256 );
and  g10909 ( new_n13258 , new_n13253 , new_n13257 );
xnor g10910 ( new_n13259 , new_n13253 , new_n13257 );
xnor g10911 ( new_n13260 , new_n13199_1 , new_n13247 );
nor  g10912 ( new_n13261 , new_n3582_1 , new_n13260 );
xnor g10913 ( new_n13262 , new_n3582_1 , new_n13260 );
xnor g10914 ( new_n13263_1 , new_n13202 , new_n13245 );
nor  g10915 ( new_n13264 , new_n3601 , new_n13263_1 );
xnor g10916 ( new_n13265 , new_n3601 , new_n13263_1 );
xnor g10917 ( new_n13266 , new_n13205 , new_n13243 );
nor  g10918 ( new_n13267 , new_n3610 , new_n13266 );
xnor g10919 ( new_n13268 , new_n3610 , new_n13266 );
xnor g10920 ( new_n13269 , new_n13208 , new_n13241 );
not  g10921 ( new_n13270_1 , new_n13269 );
and  g10922 ( new_n13271 , new_n3613 , new_n13270_1 );
xnor g10923 ( new_n13272 , new_n3613 , new_n13270_1 );
xnor g10924 ( new_n13273_1 , new_n13212 , new_n13239 );
not  g10925 ( new_n13274 , new_n13273_1 );
and  g10926 ( new_n13275 , new_n3617_1 , new_n13274 );
xnor g10927 ( new_n13276 , new_n3617_1 , new_n13274 );
xnor g10928 ( new_n13277 , new_n13216 , new_n13237 );
and  g10929 ( new_n13278 , new_n3622 , new_n13277 );
xnor g10930 ( new_n13279 , new_n3622 , new_n13277 );
xor  g10931 ( new_n13280 , new_n13220 , new_n13235 );
nor  g10932 ( new_n13281 , new_n3627 , new_n13280 );
xnor g10933 ( new_n13282 , new_n3627 , new_n13280 );
xor  g10934 ( new_n13283 , new_n13224 , new_n13233 );
nor  g10935 ( new_n13284 , new_n3632 , new_n13283 );
xnor g10936 ( new_n13285_1 , new_n3632 , new_n13283 );
xor  g10937 ( new_n13286 , new_n13228 , new_n13231 );
nor  g10938 ( new_n13287 , new_n3638 , new_n13286 );
xnor g10939 ( new_n13288 , new_n5956 , new_n13225 );
nor  g10940 ( new_n13289 , new_n3641 , new_n13288 );
xnor g10941 ( new_n13290 , new_n3639 , new_n13286 );
and  g10942 ( new_n13291 , new_n13289 , new_n13290 );
nor  g10943 ( new_n13292 , new_n13287 , new_n13291 );
nor  g10944 ( new_n13293 , new_n13285_1 , new_n13292 );
nor  g10945 ( new_n13294 , new_n13284 , new_n13293 );
nor  g10946 ( new_n13295 , new_n13282 , new_n13294 );
nor  g10947 ( new_n13296 , new_n13281 , new_n13295 );
nor  g10948 ( new_n13297 , new_n13279 , new_n13296 );
nor  g10949 ( new_n13298 , new_n13278 , new_n13297 );
nor  g10950 ( new_n13299 , new_n13276 , new_n13298 );
nor  g10951 ( new_n13300 , new_n13275 , new_n13299 );
nor  g10952 ( new_n13301 , new_n13272 , new_n13300 );
nor  g10953 ( new_n13302 , new_n13271 , new_n13301 );
nor  g10954 ( new_n13303 , new_n13268 , new_n13302 );
nor  g10955 ( new_n13304 , new_n13267 , new_n13303 );
nor  g10956 ( new_n13305 , new_n13265 , new_n13304 );
nor  g10957 ( new_n13306 , new_n13264 , new_n13305 );
nor  g10958 ( new_n13307 , new_n13262 , new_n13306 );
nor  g10959 ( new_n13308 , new_n13261 , new_n13307 );
nor  g10960 ( new_n13309 , new_n13259 , new_n13308 );
nor  g10961 ( new_n13310 , new_n13258 , new_n13309 );
xor  g10962 ( n2561 , new_n13251 , new_n13310 );
xor  g10963 ( n2573 , new_n8421 , new_n8423 );
xnor g10964 ( new_n13313 , n10411 , n18558 );
nor  g10965 ( new_n13314 , n7149 , new_n10003 );
nor  g10966 ( new_n13315 , new_n2695 , n16971 );
nor  g10967 ( new_n13316 , new_n2756 , n14148 );
nor  g10968 ( new_n13317 , n11503 , new_n2701 );
nor  g10969 ( new_n13318 , n1152 , new_n2828 );
not  g10970 ( new_n13319_1 , new_n13318 );
nor  g10971 ( new_n13320 , new_n13317 , new_n13319_1 );
nor  g10972 ( new_n13321 , new_n13316 , new_n13320 );
nor  g10973 ( new_n13322 , new_n13315 , new_n13321 );
or   g10974 ( new_n13323 , new_n13314 , new_n13322 );
xor  g10975 ( new_n13324 , new_n13313 , new_n13323 );
nor  g10976 ( new_n13325 , new_n9834 , n7963 );
nor  g10977 ( new_n13326 , n6590 , new_n9835 );
nor  g10978 ( new_n13327 , n10017 , new_n9830 );
or   g10979 ( new_n13328 , new_n7941 , n20349 );
nor  g10980 ( new_n13329 , n3618 , new_n9828 );
and  g10981 ( new_n13330 , new_n13328 , new_n13329 );
nor  g10982 ( new_n13331 , new_n13327 , new_n13330 );
nor  g10983 ( new_n13332 , new_n13326 , new_n13331 );
nor  g10984 ( new_n13333_1 , new_n13325 , new_n13332 );
xnor g10985 ( new_n13334 , new_n9874 , new_n13333_1 );
not  g10986 ( new_n13335 , new_n13334 );
xnor g10987 ( new_n13336 , new_n13324 , new_n13335 );
xnor g10988 ( new_n13337 , n7149 , n16971 );
xnor g10989 ( new_n13338_1 , new_n13321 , new_n13337 );
xnor g10990 ( new_n13339 , new_n9879 , new_n13331 );
nor  g10991 ( new_n13340 , new_n13338_1 , new_n13339 );
not  g10992 ( new_n13341 , new_n13339 );
xnor g10993 ( new_n13342 , new_n13338_1 , new_n13341 );
xnor g10994 ( new_n13343 , n1152 , n18151 );
or   g10995 ( new_n13344 , new_n9885 , new_n13343 );
xnor g10996 ( new_n13345 , n11503 , n14148 );
xnor g10997 ( new_n13346 , new_n13319_1 , new_n13345 );
and  g10998 ( new_n13347 , new_n13344 , new_n13346 );
nor  g10999 ( new_n13348 , new_n9885 , new_n13343 );
xnor g11000 ( new_n13349 , new_n13348 , new_n13346 );
xor  g11001 ( new_n13350 , new_n9882 , new_n13329 );
and  g11002 ( new_n13351 , new_n13349 , new_n13350 );
nor  g11003 ( new_n13352 , new_n13347 , new_n13351 );
and  g11004 ( new_n13353 , new_n13342 , new_n13352 );
nor  g11005 ( new_n13354 , new_n13340 , new_n13353 );
xnor g11006 ( new_n13355 , new_n13336 , new_n13354 );
not  g11007 ( new_n13356 , new_n13355 );
xnor g11008 ( new_n13357 , n17035 , n19515 );
not  g11009 ( new_n13358 , n22588 );
nor  g11010 ( new_n13359 , n14684 , new_n13358 );
nor  g11011 ( new_n13360 , new_n8445 , n22588 );
and  g11012 ( new_n13361 , new_n4180 , n12209 );
nor  g11013 ( new_n13362 , new_n4180 , n12209 );
nor  g11014 ( new_n13363 , new_n13145 , n24732 );
not  g11015 ( new_n13364 , new_n13363 );
nor  g11016 ( new_n13365 , new_n13362 , new_n13364 );
nor  g11017 ( new_n13366 , new_n13361 , new_n13365 );
nor  g11018 ( new_n13367_1 , new_n13360 , new_n13366 );
nor  g11019 ( new_n13368 , new_n13359 , new_n13367_1 );
xnor g11020 ( new_n13369 , new_n13357 , new_n13368 );
not  g11021 ( new_n13370 , new_n13369 );
xnor g11022 ( new_n13371 , new_n13356 , new_n13370 );
xnor g11023 ( new_n13372 , new_n13342 , new_n13352 );
xnor g11024 ( new_n13373 , n14684 , n22588 );
xnor g11025 ( new_n13374 , new_n13366 , new_n13373 );
and  g11026 ( new_n13375 , new_n13372 , new_n13374 );
xnor g11027 ( new_n13376 , n12892 , n24732 );
xnor g11028 ( new_n13377 , new_n9885 , new_n13343 );
nor  g11029 ( new_n13378 , new_n13376 , new_n13377 );
xnor g11030 ( new_n13379 , n6631 , n12209 );
xnor g11031 ( new_n13380 , new_n13364 , new_n13379 );
not  g11032 ( new_n13381 , new_n13380 );
nor  g11033 ( new_n13382 , new_n13378 , new_n13381 );
xnor g11034 ( new_n13383 , new_n13378 , new_n13380 );
xnor g11035 ( new_n13384 , new_n9882 , new_n13329 );
xnor g11036 ( new_n13385 , new_n13349 , new_n13384 );
and  g11037 ( new_n13386 , new_n13383 , new_n13385 );
nor  g11038 ( new_n13387 , new_n13382 , new_n13386 );
xnor g11039 ( new_n13388 , new_n13372 , new_n13374 );
nor  g11040 ( new_n13389 , new_n13387 , new_n13388 );
nor  g11041 ( new_n13390 , new_n13375 , new_n13389 );
xnor g11042 ( n2578 , new_n13371 , new_n13390 );
not  g11043 ( new_n13392 , new_n11607_1 );
nor  g11044 ( new_n13393 , new_n7835 , new_n13392 );
not  g11045 ( new_n13394 , new_n7835 );
xnor g11046 ( new_n13395 , new_n13394 , new_n13392 );
nor  g11047 ( new_n13396 , new_n7771 , new_n13394 );
and  g11048 ( new_n13397 , new_n7836 , new_n7916 );
or   g11049 ( new_n13398 , new_n13396 , new_n13397 );
and  g11050 ( new_n13399 , new_n13395 , new_n13398 );
nor  g11051 ( n2582 , new_n13393 , new_n13399 );
xor  g11052 ( n2602 , new_n4295 , new_n4306_1 );
nor  g11053 ( new_n13402 , n2420 , n22201 );
not  g11054 ( new_n13403 , new_n13402 );
nor  g11055 ( new_n13404 , n24485 , new_n13403 );
not  g11056 ( new_n13405 , new_n13404 );
nor  g11057 ( new_n13406 , n21078 , new_n13405 );
not  g11058 ( new_n13407_1 , new_n13406 );
nor  g11059 ( new_n13408 , n12546 , new_n13407_1 );
xnor g11060 ( new_n13409_1 , n8324 , new_n13408 );
xnor g11061 ( new_n13410 , new_n3963 , new_n13409_1 );
xnor g11062 ( new_n13411 , n12546 , new_n13406 );
nor  g11063 ( new_n13412 , new_n3965 , new_n13411 );
xnor g11064 ( new_n13413 , n21078 , new_n13404 );
nor  g11065 ( new_n13414 , new_n3970 , new_n13413 );
xnor g11066 ( new_n13415 , new_n3968 , new_n13413 );
xnor g11067 ( new_n13416 , n24485 , new_n13402 );
and  g11068 ( new_n13417 , new_n3976 , new_n13416 );
xnor g11069 ( new_n13418 , new_n3974 , new_n13416 );
xnor g11070 ( new_n13419_1 , new_n8112 , n22201 );
nor  g11071 ( new_n13420 , new_n3984_1 , new_n13419_1 );
or   g11072 ( new_n13421 , new_n8110 , new_n2551 );
xnor g11073 ( new_n13422 , new_n3980 , new_n13419_1 );
and  g11074 ( new_n13423 , new_n13421 , new_n13422 );
nor  g11075 ( new_n13424_1 , new_n13420 , new_n13423 );
and  g11076 ( new_n13425 , new_n13418 , new_n13424_1 );
nor  g11077 ( new_n13426 , new_n13417 , new_n13425 );
and  g11078 ( new_n13427 , new_n13415 , new_n13426 );
nor  g11079 ( new_n13428 , new_n13414 , new_n13427 );
xnor g11080 ( new_n13429 , new_n3965 , new_n13411 );
nor  g11081 ( new_n13430 , new_n13428 , new_n13429 );
nor  g11082 ( new_n13431 , new_n13412 , new_n13430 );
xnor g11083 ( new_n13432 , new_n13410 , new_n13431 );
xnor g11084 ( new_n13433 , n7678 , new_n8093 );
nor  g11085 ( new_n13434 , n3785 , new_n8095_1 );
xnor g11086 ( new_n13435 , new_n4377 , new_n8095_1 );
nor  g11087 ( new_n13436 , n20250 , new_n8099 );
xnor g11088 ( new_n13437 , new_n4382 , new_n8099 );
nor  g11089 ( new_n13438 , new_n4384 , new_n8103_1 );
or   g11090 ( new_n13439 , n5822 , new_n8104 );
nor  g11091 ( new_n13440 , n26443 , new_n8108 );
or   g11092 ( new_n13441 , new_n4394 , new_n2545 );
xnor g11093 ( new_n13442 , new_n6644 , new_n8108 );
and  g11094 ( new_n13443 , new_n13441 , new_n13442 );
nor  g11095 ( new_n13444 , new_n13440 , new_n13443 );
and  g11096 ( new_n13445 , new_n13439 , new_n13444 );
nor  g11097 ( new_n13446 , new_n13438 , new_n13445 );
and  g11098 ( new_n13447 , new_n13437 , new_n13446 );
or   g11099 ( new_n13448 , new_n13436 , new_n13447 );
and  g11100 ( new_n13449 , new_n13435 , new_n13448 );
nor  g11101 ( new_n13450 , new_n13434 , new_n13449 );
xor  g11102 ( new_n13451 , new_n13433 , new_n13450 );
xnor g11103 ( new_n13452 , new_n13432 , new_n13451 );
xor  g11104 ( new_n13453_1 , new_n13435 , new_n13448 );
xnor g11105 ( new_n13454 , new_n13428 , new_n13429 );
not  g11106 ( new_n13455 , new_n13454 );
and  g11107 ( new_n13456_1 , new_n13453_1 , new_n13455 );
xnor g11108 ( new_n13457_1 , new_n13453_1 , new_n13455 );
xnor g11109 ( new_n13458 , new_n13415 , new_n13426 );
xnor g11110 ( new_n13459 , new_n13437 , new_n13446 );
nor  g11111 ( new_n13460_1 , new_n13458 , new_n13459 );
xor  g11112 ( new_n13461 , new_n13458 , new_n13459 );
xnor g11113 ( new_n13462 , new_n13418 , new_n13424_1 );
xnor g11114 ( new_n13463 , new_n4384 , new_n8104 );
xnor g11115 ( new_n13464 , new_n13444 , new_n13463 );
nor  g11116 ( new_n13465 , new_n13462 , new_n13464 );
xor  g11117 ( new_n13466 , new_n13421 , new_n13422 );
xor  g11118 ( new_n13467 , new_n13441 , new_n13442 );
and  g11119 ( new_n13468 , new_n13466 , new_n13467 );
xnor g11120 ( new_n13469 , new_n4394 , new_n2545 );
xnor g11121 ( new_n13470 , n22201 , new_n2551 );
not  g11122 ( new_n13471 , new_n13470 );
nor  g11123 ( new_n13472 , new_n13469 , new_n13471 );
xnor g11124 ( new_n13473 , new_n13466 , new_n13467 );
nor  g11125 ( new_n13474 , new_n13472 , new_n13473 );
nor  g11126 ( new_n13475 , new_n13468 , new_n13474 );
xor  g11127 ( new_n13476 , new_n13462 , new_n13464 );
and  g11128 ( new_n13477_1 , new_n13475 , new_n13476 );
nor  g11129 ( new_n13478 , new_n13465 , new_n13477_1 );
and  g11130 ( new_n13479 , new_n13461 , new_n13478 );
nor  g11131 ( new_n13480 , new_n13460_1 , new_n13479 );
nor  g11132 ( new_n13481 , new_n13457_1 , new_n13480 );
nor  g11133 ( new_n13482 , new_n13456_1 , new_n13481 );
xnor g11134 ( n2619 , new_n13452 , new_n13482 );
nor  g11135 ( new_n13484_1 , n12900 , new_n5917 );
xnor g11136 ( new_n13485 , n12900 , new_n5917 );
nor  g11137 ( new_n13486_1 , n20411 , new_n5923 );
xnor g11138 ( new_n13487_1 , n20411 , new_n5923 );
nor  g11139 ( new_n13488 , n17069 , new_n5928 );
xnor g11140 ( new_n13489 , n17069 , new_n5928 );
nor  g11141 ( new_n13490_1 , n15918 , new_n5933 );
nor  g11142 ( new_n13491 , n17784 , new_n5938 );
xnor g11143 ( new_n13492 , n17784 , new_n5938 );
and  g11144 ( new_n13493 , n14323 , new_n5943_1 );
nor  g11145 ( new_n13494_1 , new_n12840 , new_n12850 );
nor  g11146 ( new_n13495 , new_n13493 , new_n13494_1 );
not  g11147 ( new_n13496 , new_n13495 );
nor  g11148 ( new_n13497 , new_n13492 , new_n13496 );
nor  g11149 ( new_n13498 , new_n13491 , new_n13497 );
xnor g11150 ( new_n13499 , n15918 , new_n5933 );
nor  g11151 ( new_n13500_1 , new_n13498 , new_n13499 );
nor  g11152 ( new_n13501_1 , new_n13490_1 , new_n13500_1 );
nor  g11153 ( new_n13502 , new_n13489 , new_n13501_1 );
nor  g11154 ( new_n13503 , new_n13488 , new_n13502 );
nor  g11155 ( new_n13504 , new_n13487_1 , new_n13503 );
nor  g11156 ( new_n13505 , new_n13486_1 , new_n13504 );
nor  g11157 ( new_n13506_1 , new_n13485 , new_n13505 );
nor  g11158 ( new_n13507 , new_n13484_1 , new_n13506_1 );
not  g11159 ( new_n13508 , new_n5871 );
xnor g11160 ( new_n13509 , n10650 , new_n13508 );
xnor g11161 ( new_n13510 , new_n13507 , new_n13509 );
not  g11162 ( new_n13511 , new_n13510 );
nor  g11163 ( new_n13512 , n6456 , new_n13511 );
xnor g11164 ( new_n13513 , new_n5872 , new_n13511 );
xnor g11165 ( new_n13514 , new_n13485 , new_n13505 );
nor  g11166 ( new_n13515 , n4085 , new_n13514 );
not  g11167 ( new_n13516 , new_n13514 );
xnor g11168 ( new_n13517 , n4085 , new_n13516 );
xnor g11169 ( new_n13518 , new_n13487_1 , new_n13503 );
nor  g11170 ( new_n13519 , n26725 , new_n13518 );
not  g11171 ( new_n13520 , new_n13518 );
xnor g11172 ( new_n13521 , n26725 , new_n13520 );
xnor g11173 ( new_n13522 , new_n13489 , new_n13501_1 );
nor  g11174 ( new_n13523 , n11980 , new_n13522 );
not  g11175 ( new_n13524 , new_n13522 );
xnor g11176 ( new_n13525 , n11980 , new_n13524 );
xnor g11177 ( new_n13526 , new_n13498 , new_n13499 );
nor  g11178 ( new_n13527 , n3253 , new_n13526 );
xnor g11179 ( new_n13528 , new_n5883 , new_n13526 );
xnor g11180 ( new_n13529 , new_n13492 , new_n13495 );
nor  g11181 ( new_n13530 , new_n5886 , new_n13529 );
not  g11182 ( new_n13531 , new_n13529 );
xnor g11183 ( new_n13532 , new_n5886 , new_n13531 );
nor  g11184 ( new_n13533 , new_n5889 , new_n12851 );
and  g11185 ( new_n13534 , new_n12852 , new_n12863 );
or   g11186 ( new_n13535 , new_n13533 , new_n13534 );
and  g11187 ( new_n13536 , new_n13532 , new_n13535 );
nor  g11188 ( new_n13537 , new_n13530 , new_n13536 );
and  g11189 ( new_n13538 , new_n13528 , new_n13537 );
or   g11190 ( new_n13539 , new_n13527 , new_n13538 );
and  g11191 ( new_n13540 , new_n13525 , new_n13539 );
or   g11192 ( new_n13541 , new_n13523 , new_n13540 );
and  g11193 ( new_n13542 , new_n13521 , new_n13541 );
or   g11194 ( new_n13543 , new_n13519 , new_n13542 );
and  g11195 ( new_n13544 , new_n13517 , new_n13543 );
or   g11196 ( new_n13545 , new_n13515 , new_n13544 );
and  g11197 ( new_n13546 , new_n13513 , new_n13545 );
nor  g11198 ( new_n13547 , new_n13512 , new_n13546 );
or   g11199 ( new_n13548_1 , n10650 , new_n5871 );
and  g11200 ( new_n13549_1 , new_n13507 , new_n13548_1 );
and  g11201 ( new_n13550 , new_n4798 , new_n5870 );
and  g11202 ( new_n13551_1 , n10650 , new_n5871 );
or   g11203 ( new_n13552 , new_n13550 , new_n13551_1 );
nor  g11204 ( new_n13553 , new_n13549_1 , new_n13552 );
and  g11205 ( new_n13554 , new_n13547 , new_n13553 );
nor  g11206 ( new_n13555 , new_n12592 , new_n13554 );
xnor g11207 ( new_n13556 , new_n12592 , new_n13554 );
xnor g11208 ( new_n13557 , new_n13547 , new_n13553 );
and  g11209 ( new_n13558 , new_n12596 , new_n13557 );
xnor g11210 ( new_n13559 , new_n12596 , new_n13557 );
xor  g11211 ( new_n13560 , new_n13513 , new_n13545 );
and  g11212 ( new_n13561 , new_n12601 , new_n13560 );
xnor g11213 ( new_n13562 , new_n12601 , new_n13560 );
xor  g11214 ( new_n13563 , new_n13517 , new_n13543 );
and  g11215 ( new_n13564 , new_n12606 , new_n13563 );
xnor g11216 ( new_n13565 , new_n12606 , new_n13563 );
xor  g11217 ( new_n13566 , new_n13521 , new_n13541 );
and  g11218 ( new_n13567 , new_n12611 , new_n13566 );
xnor g11219 ( new_n13568 , new_n12611 , new_n13566 );
xor  g11220 ( new_n13569 , new_n13525 , new_n13539 );
and  g11221 ( new_n13570 , new_n12616 , new_n13569 );
xnor g11222 ( new_n13571 , new_n12616 , new_n13569 );
xnor g11223 ( new_n13572 , new_n13528 , new_n13537 );
nor  g11224 ( new_n13573 , new_n12622 , new_n13572 );
xnor g11225 ( new_n13574 , new_n12622 , new_n13572 );
xor  g11226 ( new_n13575 , new_n13532 , new_n13535 );
nor  g11227 ( new_n13576 , new_n12626_1 , new_n13575 );
xnor g11228 ( new_n13577 , new_n12626_1 , new_n13575 );
nor  g11229 ( new_n13578 , new_n12630 , new_n12864_1 );
nor  g11230 ( new_n13579 , new_n12865_1 , new_n12878 );
nor  g11231 ( new_n13580 , new_n13578 , new_n13579 );
nor  g11232 ( new_n13581 , new_n13577 , new_n13580 );
nor  g11233 ( new_n13582 , new_n13576 , new_n13581 );
nor  g11234 ( new_n13583 , new_n13574 , new_n13582 );
nor  g11235 ( new_n13584 , new_n13573 , new_n13583 );
nor  g11236 ( new_n13585 , new_n13571 , new_n13584 );
nor  g11237 ( new_n13586 , new_n13570 , new_n13585 );
nor  g11238 ( new_n13587 , new_n13568 , new_n13586 );
nor  g11239 ( new_n13588 , new_n13567 , new_n13587 );
nor  g11240 ( new_n13589 , new_n13565 , new_n13588 );
nor  g11241 ( new_n13590 , new_n13564 , new_n13589 );
nor  g11242 ( new_n13591 , new_n13562 , new_n13590 );
nor  g11243 ( new_n13592 , new_n13561 , new_n13591 );
nor  g11244 ( new_n13593 , new_n13559 , new_n13592 );
nor  g11245 ( new_n13594 , new_n13558 , new_n13593 );
nor  g11246 ( new_n13595 , new_n13556 , new_n13594 );
nor  g11247 ( n2661 , new_n13555 , new_n13595 );
xnor g11248 ( n2693 , new_n11068 , new_n11070 );
xnor g11249 ( new_n13598 , new_n7288 , new_n13324 );
nor  g11250 ( new_n13599 , new_n7295 , new_n13338_1 );
xnor g11251 ( new_n13600 , new_n7295 , new_n13338_1 );
nor  g11252 ( new_n13601 , new_n7298_1 , new_n13346 );
nor  g11253 ( new_n13602_1 , new_n7300 , new_n13343 );
xnor g11254 ( new_n13603 , new_n7302 , new_n13346 );
and  g11255 ( new_n13604 , new_n13602_1 , new_n13603 );
nor  g11256 ( new_n13605 , new_n13601 , new_n13604 );
nor  g11257 ( new_n13606 , new_n13600 , new_n13605 );
nor  g11258 ( new_n13607 , new_n13599 , new_n13606 );
xnor g11259 ( new_n13608 , new_n13598 , new_n13607 );
not  g11260 ( new_n13609 , new_n13608 );
xnor g11261 ( new_n13610 , n4665 , n8309 );
nor  g11262 ( new_n13611 , n19005 , new_n8759 );
nor  g11263 ( new_n13612 , new_n2866 , n19144 );
nor  g11264 ( new_n13613 , n4326 , new_n10007 );
or   g11265 ( new_n13614 , new_n2869 , n12593 );
nor  g11266 ( new_n13615 , n5438 , new_n8763 );
and  g11267 ( new_n13616 , new_n13614 , new_n13615 );
nor  g11268 ( new_n13617 , new_n13613 , new_n13616 );
nor  g11269 ( new_n13618 , new_n13612 , new_n13617 );
or   g11270 ( new_n13619 , new_n13611 , new_n13618 );
xor  g11271 ( new_n13620 , new_n13610 , new_n13619 );
xnor g11272 ( new_n13621 , new_n13609 , new_n13620 );
xnor g11273 ( new_n13622 , new_n13600 , new_n13605 );
xnor g11274 ( new_n13623 , n19005 , n19144 );
xnor g11275 ( new_n13624 , new_n13617 , new_n13623 );
and  g11276 ( new_n13625 , new_n13622 , new_n13624 );
xnor g11277 ( new_n13626_1 , new_n13622 , new_n13624 );
xnor g11278 ( new_n13627 , n5438 , n13714 );
xnor g11279 ( new_n13628 , new_n7399 , new_n13343 );
not  g11280 ( new_n13629 , new_n13628 );
nor  g11281 ( new_n13630 , new_n13627 , new_n13629 );
xnor g11282 ( new_n13631 , n4326 , n12593 );
xnor g11283 ( new_n13632 , new_n13615 , new_n13631 );
nor  g11284 ( new_n13633 , new_n13630 , new_n13632 );
xnor g11285 ( new_n13634 , new_n13602_1 , new_n13603 );
not  g11286 ( new_n13635 , new_n13634 );
xnor g11287 ( new_n13636 , new_n13630 , new_n13632 );
nor  g11288 ( new_n13637 , new_n13635 , new_n13636 );
nor  g11289 ( new_n13638 , new_n13633 , new_n13637 );
nor  g11290 ( new_n13639 , new_n13626_1 , new_n13638 );
nor  g11291 ( new_n13640 , new_n13625 , new_n13639 );
xnor g11292 ( n2703 , new_n13621 , new_n13640 );
xnor g11293 ( n2706 , new_n12711 , new_n12720 );
nor  g11294 ( new_n13643 , new_n6152 , n3320 );
xnor g11295 ( new_n13644 , n1831 , n3320 );
not  g11296 ( new_n13645 , n13137 );
nor  g11297 ( new_n13646 , n1288 , new_n13645 );
xnor g11298 ( new_n13647 , n1288 , n13137 );
not  g11299 ( new_n13648 , n18452 );
nor  g11300 ( new_n13649 , n1752 , new_n13648 );
xnor g11301 ( new_n13650 , n1752 , n18452 );
not  g11302 ( new_n13651 , n21317 );
nor  g11303 ( new_n13652 , n13110 , new_n13651 );
xnor g11304 ( new_n13653 , n13110 , n21317 );
nor  g11305 ( new_n13654 , new_n6164 , n25694 );
xnor g11306 ( new_n13655 , n12398 , n25694 );
nor  g11307 ( new_n13656 , n15424 , new_n6167 );
xnor g11308 ( new_n13657 , n15424 , n19789 );
not  g11309 ( new_n13658 , n1949 );
nor  g11310 ( new_n13659 , new_n13658 , n20169 );
and  g11311 ( new_n13660 , new_n12016 , new_n12025 );
nor  g11312 ( new_n13661 , new_n13659 , new_n13660 );
and  g11313 ( new_n13662 , new_n13657 , new_n13661 );
or   g11314 ( new_n13663 , new_n13656 , new_n13662 );
and  g11315 ( new_n13664 , new_n13655 , new_n13663 );
or   g11316 ( new_n13665 , new_n13654 , new_n13664 );
and  g11317 ( new_n13666 , new_n13653 , new_n13665 );
or   g11318 ( new_n13667 , new_n13652 , new_n13666 );
and  g11319 ( new_n13668_1 , new_n13650 , new_n13667 );
or   g11320 ( new_n13669 , new_n13649 , new_n13668_1 );
and  g11321 ( new_n13670 , new_n13647 , new_n13669 );
or   g11322 ( new_n13671 , new_n13646 , new_n13670 );
and  g11323 ( new_n13672 , new_n13644 , new_n13671 );
nor  g11324 ( new_n13673 , new_n13643 , new_n13672 );
not  g11325 ( new_n13674 , new_n13673 );
not  g11326 ( new_n13675 , n1483 );
nor  g11327 ( new_n13676 , new_n13675 , n19539 );
and  g11328 ( new_n13677_1 , new_n11154 , new_n11168 );
nor  g11329 ( new_n13678 , new_n13676 , new_n13677_1 );
not  g11330 ( new_n13679 , new_n6470_1 );
nor  g11331 ( new_n13680 , n16818 , new_n13679 );
not  g11332 ( new_n13681 , new_n13680 );
nor  g11333 ( new_n13682 , n3541 , new_n13681 );
xnor g11334 ( new_n13683_1 , n2184 , new_n13682 );
nor  g11335 ( new_n13684 , n6204 , new_n13683_1 );
not  g11336 ( new_n13685 , new_n13683_1 );
xnor g11337 ( new_n13686 , n6204 , new_n13685 );
xnor g11338 ( new_n13687 , n3541 , new_n13680 );
not  g11339 ( new_n13688 , new_n13687 );
nor  g11340 ( new_n13689 , new_n12116 , new_n13688 );
nor  g11341 ( new_n13690 , n3349 , new_n13687 );
nor  g11342 ( new_n13691 , new_n12119 , new_n6472 );
or   g11343 ( new_n13692 , n1742 , new_n6471 );
and  g11344 ( new_n13693 , new_n13692 , new_n6506_1 );
nor  g11345 ( new_n13694 , new_n13691 , new_n13693 );
nor  g11346 ( new_n13695 , new_n13690 , new_n13694 );
nor  g11347 ( new_n13696 , new_n13689 , new_n13695 );
and  g11348 ( new_n13697 , new_n13686 , new_n13696 );
nor  g11349 ( new_n13698 , new_n13684 , new_n13697 );
not  g11350 ( new_n13699 , new_n13682 );
nor  g11351 ( new_n13700 , n2184 , new_n13699 );
xnor g11352 ( new_n13701 , n10018 , new_n13700 );
not  g11353 ( new_n13702 , new_n13701 );
xnor g11354 ( new_n13703 , new_n12110 , new_n13702 );
xnor g11355 ( new_n13704 , new_n13698 , new_n13703 );
nor  g11356 ( new_n13705 , new_n11169 , new_n13704 );
xnor g11357 ( new_n13706 , new_n11169 , new_n13704 );
xnor g11358 ( new_n13707 , new_n13686 , new_n13696 );
nor  g11359 ( new_n13708_1 , new_n11228 , new_n13707 );
xnor g11360 ( new_n13709 , new_n11228 , new_n13707 );
not  g11361 ( new_n13710_1 , new_n13709 );
xnor g11362 ( new_n13711 , n3349 , new_n13688 );
xnor g11363 ( new_n13712 , new_n13694 , new_n13711 );
and  g11364 ( new_n13713 , new_n11232 , new_n13712 );
xnor g11365 ( new_n13714_1 , new_n11232 , new_n13712 );
and  g11366 ( new_n13715 , new_n6461 , new_n6508 );
nor  g11367 ( new_n13716 , new_n6509 , new_n6550 );
nor  g11368 ( new_n13717 , new_n13715 , new_n13716 );
nor  g11369 ( new_n13718 , new_n13714_1 , new_n13717 );
nor  g11370 ( new_n13719_1 , new_n13713 , new_n13718 );
and  g11371 ( new_n13720 , new_n13710_1 , new_n13719_1 );
nor  g11372 ( new_n13721 , new_n13708_1 , new_n13720 );
nor  g11373 ( new_n13722_1 , new_n13706 , new_n13721 );
nor  g11374 ( new_n13723 , new_n13705 , new_n13722_1 );
and  g11375 ( new_n13724 , new_n12158_1 , new_n13700 );
nor  g11376 ( new_n13725 , n5140 , new_n13701 );
nor  g11377 ( new_n13726 , new_n12110 , new_n13702 );
nor  g11378 ( new_n13727 , new_n13698 , new_n13726 );
nor  g11379 ( new_n13728 , new_n13725 , new_n13727 );
nor  g11380 ( new_n13729 , new_n13724 , new_n13728 );
not  g11381 ( new_n13730 , new_n13729 );
and  g11382 ( new_n13731 , new_n13723 , new_n13730 );
and  g11383 ( new_n13732 , new_n13678 , new_n13731 );
or   g11384 ( new_n13733 , new_n13723 , new_n13730 );
nor  g11385 ( new_n13734 , new_n13678 , new_n13733 );
nor  g11386 ( new_n13735 , new_n13732 , new_n13734 );
not  g11387 ( new_n13736 , new_n13735 );
xnor g11388 ( new_n13737 , new_n13674 , new_n13736 );
xnor g11389 ( new_n13738 , new_n13723 , new_n13729 );
xnor g11390 ( new_n13739 , new_n13678 , new_n13738 );
and  g11391 ( new_n13740 , new_n13673 , new_n13739 );
or   g11392 ( new_n13741 , new_n13673 , new_n13739 );
xor  g11393 ( new_n13742 , new_n13644 , new_n13671 );
xnor g11394 ( new_n13743 , new_n13706 , new_n13721 );
nor  g11395 ( new_n13744 , new_n13742 , new_n13743 );
xnor g11396 ( new_n13745 , new_n13742 , new_n13743 );
xor  g11397 ( new_n13746 , new_n13647 , new_n13669 );
xnor g11398 ( new_n13747 , new_n13710_1 , new_n13719_1 );
nor  g11399 ( new_n13748 , new_n13746 , new_n13747 );
xnor g11400 ( new_n13749 , new_n13746 , new_n13747 );
xor  g11401 ( new_n13750 , new_n13650 , new_n13667 );
xnor g11402 ( new_n13751 , new_n13714_1 , new_n13717 );
not  g11403 ( new_n13752 , new_n13751 );
nor  g11404 ( new_n13753 , new_n13750 , new_n13752 );
xnor g11405 ( new_n13754_1 , new_n13750 , new_n13752 );
xor  g11406 ( new_n13755 , new_n13653 , new_n13665 );
nor  g11407 ( new_n13756 , new_n6552 , new_n13755 );
xor  g11408 ( new_n13757 , new_n13655 , new_n13663 );
nor  g11409 ( new_n13758 , new_n6554 , new_n13757 );
xnor g11410 ( new_n13759 , new_n6554 , new_n13757 );
not  g11411 ( new_n13760 , new_n6557 );
xnor g11412 ( new_n13761 , new_n13657 , new_n13661 );
and  g11413 ( new_n13762 , new_n13760 , new_n13761 );
xnor g11414 ( new_n13763 , new_n13760 , new_n13761 );
and  g11415 ( new_n13764_1 , new_n6560_1 , new_n12026 );
nor  g11416 ( new_n13765 , new_n12027 , new_n12041 );
nor  g11417 ( new_n13766 , new_n13764_1 , new_n13765 );
nor  g11418 ( new_n13767 , new_n13763 , new_n13766 );
nor  g11419 ( new_n13768 , new_n13762 , new_n13767 );
nor  g11420 ( new_n13769 , new_n13759 , new_n13768 );
nor  g11421 ( new_n13770 , new_n13758 , new_n13769 );
xnor g11422 ( new_n13771 , new_n6552 , new_n13755 );
nor  g11423 ( new_n13772 , new_n13770 , new_n13771 );
nor  g11424 ( new_n13773 , new_n13756 , new_n13772 );
nor  g11425 ( new_n13774 , new_n13754_1 , new_n13773 );
nor  g11426 ( new_n13775_1 , new_n13753 , new_n13774 );
nor  g11427 ( new_n13776 , new_n13749 , new_n13775_1 );
nor  g11428 ( new_n13777 , new_n13748 , new_n13776 );
nor  g11429 ( new_n13778 , new_n13745 , new_n13777 );
nor  g11430 ( new_n13779 , new_n13744 , new_n13778 );
and  g11431 ( new_n13780 , new_n13741 , new_n13779 );
nor  g11432 ( new_n13781_1 , new_n13740 , new_n13780 );
xnor g11433 ( n2711 , new_n13737 , new_n13781_1 );
xnor g11434 ( new_n13783_1 , n2680 , n10611 );
nor  g11435 ( new_n13784 , new_n10614_1 , n2783 );
nor  g11436 ( new_n13785 , n1667 , new_n6593 );
and  g11437 ( new_n13786 , n7339 , new_n9099 );
or   g11438 ( new_n13787 , n7339 , new_n9099 );
nor  g11439 ( new_n13788 , n18 , new_n9155 );
and  g11440 ( new_n13789 , new_n13787 , new_n13788 );
nor  g11441 ( new_n13790 , new_n13786 , new_n13789 );
nor  g11442 ( new_n13791 , new_n13785 , new_n13790 );
or   g11443 ( new_n13792 , new_n13784 , new_n13791 );
xor  g11444 ( new_n13793 , new_n13783_1 , new_n13792 );
xnor g11445 ( new_n13794 , new_n9023 , new_n13793 );
xnor g11446 ( new_n13795 , n1667 , n2783 );
xnor g11447 ( new_n13796 , new_n13790 , new_n13795 );
and  g11448 ( new_n13797 , new_n9027 , new_n13796 );
xnor g11449 ( new_n13798_1 , new_n9027 , new_n13796 );
xnor g11450 ( new_n13799 , n18 , n26808 );
nor  g11451 ( new_n13800 , new_n9034 , new_n13799 );
xnor g11452 ( new_n13801 , n7339 , n15490 );
xnor g11453 ( new_n13802 , new_n13788 , new_n13801 );
nor  g11454 ( new_n13803 , new_n13800 , new_n13802 );
xnor g11455 ( new_n13804 , new_n13800 , new_n13802 );
nor  g11456 ( new_n13805 , new_n9039 , new_n13804 );
nor  g11457 ( new_n13806 , new_n13803 , new_n13805 );
nor  g11458 ( new_n13807 , new_n13798_1 , new_n13806 );
nor  g11459 ( new_n13808 , new_n13797 , new_n13807 );
xnor g11460 ( n2761 , new_n13794 , new_n13808 );
xnor g11461 ( new_n13810 , n8526 , n25120 );
nor  g11462 ( new_n13811 , n2816 , n8363 );
xnor g11463 ( new_n13812 , new_n6025 , n8363 );
nor  g11464 ( new_n13813 , n14680 , n20359 );
xnor g11465 ( new_n13814 , n14680 , n20359 );
nor  g11466 ( new_n13815 , n4409 , n17250 );
or   g11467 ( new_n13816 , new_n9289 , new_n9309 );
and  g11468 ( new_n13817 , new_n9288 , new_n13816 );
nor  g11469 ( new_n13818 , new_n13815 , new_n13817 );
nor  g11470 ( new_n13819 , new_n13814 , new_n13818 );
or   g11471 ( new_n13820 , new_n13813 , new_n13819 );
and  g11472 ( new_n13821 , new_n13812 , new_n13820 );
nor  g11473 ( new_n13822 , new_n13811 , new_n13821 );
xnor g11474 ( new_n13823 , new_n13810 , new_n13822 );
nor  g11475 ( new_n13824 , n17458 , new_n13823 );
xnor g11476 ( new_n13825 , new_n10870 , new_n13823 );
nor  g11477 ( new_n13826 , new_n13813 , new_n13819 );
xnor g11478 ( new_n13827 , new_n13812 , new_n13826 );
nor  g11479 ( new_n13828 , new_n10873 , new_n13827 );
xnor g11480 ( new_n13829 , new_n13814 , new_n13818 );
nor  g11481 ( new_n13830 , n25240 , new_n13829 );
xnor g11482 ( new_n13831 , new_n10876 , new_n13829 );
nor  g11483 ( new_n13832 , new_n10414 , new_n9311 );
xnor g11484 ( new_n13833 , new_n10414 , new_n9312 );
nor  g11485 ( new_n13834 , new_n10881 , new_n9315 );
xnor g11486 ( new_n13835_1 , new_n10881 , new_n9317 );
nor  g11487 ( new_n13836 , new_n10884 , new_n9320 );
xnor g11488 ( new_n13837 , new_n10884 , new_n9322 );
nor  g11489 ( new_n13838 , new_n8432_1 , new_n9325 );
xnor g11490 ( new_n13839 , new_n8432_1 , new_n9327 );
nor  g11491 ( new_n13840 , new_n7217 , new_n9330 );
nor  g11492 ( new_n13841 , n5026 , new_n9332 );
or   g11493 ( new_n13842 , new_n6628_1 , new_n9335 );
xnor g11494 ( new_n13843 , new_n7220 , new_n9332 );
and  g11495 ( new_n13844 , new_n13842 , new_n13843 );
nor  g11496 ( new_n13845 , new_n13841 , new_n13844 );
xnor g11497 ( new_n13846 , new_n7217 , new_n9340 );
and  g11498 ( new_n13847 , new_n13845 , new_n13846 );
or   g11499 ( new_n13848 , new_n13840 , new_n13847 );
and  g11500 ( new_n13849 , new_n13839 , new_n13848 );
or   g11501 ( new_n13850_1 , new_n13838 , new_n13849 );
and  g11502 ( new_n13851_1 , new_n13837 , new_n13850_1 );
or   g11503 ( new_n13852 , new_n13836 , new_n13851_1 );
and  g11504 ( new_n13853 , new_n13835_1 , new_n13852 );
or   g11505 ( new_n13854 , new_n13834 , new_n13853 );
and  g11506 ( new_n13855 , new_n13833 , new_n13854 );
nor  g11507 ( new_n13856 , new_n13832 , new_n13855 );
and  g11508 ( new_n13857 , new_n13831 , new_n13856 );
nor  g11509 ( new_n13858 , new_n13830 , new_n13857 );
not  g11510 ( new_n13859 , new_n13827 );
xnor g11511 ( new_n13860 , new_n10873 , new_n13859 );
and  g11512 ( new_n13861 , new_n13858 , new_n13860 );
nor  g11513 ( new_n13862 , new_n13828 , new_n13861 );
and  g11514 ( new_n13863 , new_n13825 , new_n13862 );
nor  g11515 ( new_n13864 , new_n13824 , new_n13863 );
not  g11516 ( new_n13865 , new_n13864 );
nor  g11517 ( new_n13866 , n8526 , n25120 );
nor  g11518 ( new_n13867 , new_n13810 , new_n13822 );
nor  g11519 ( new_n13868 , new_n13866 , new_n13867 );
not  g11520 ( new_n13869 , new_n13868 );
nor  g11521 ( new_n13870 , new_n13865 , new_n13869 );
not  g11522 ( new_n13871 , new_n3735 );
nor  g11523 ( new_n13872 , n2113 , new_n13871 );
not  g11524 ( new_n13873 , new_n13872 );
nor  g11525 ( new_n13874 , n1099 , new_n13873 );
not  g11526 ( new_n13875 , new_n13874 );
nor  g11527 ( new_n13876 , n19941 , new_n13875 );
xnor g11528 ( new_n13877 , n11898 , new_n13876 );
nor  g11529 ( new_n13878 , new_n4837 , new_n13877 );
not  g11530 ( new_n13879 , new_n13877 );
xnor g11531 ( new_n13880 , new_n4839 , new_n13879 );
xnor g11532 ( new_n13881 , n19941 , new_n13874 );
nor  g11533 ( new_n13882 , new_n4841 , new_n13881 );
xnor g11534 ( new_n13883 , new_n4841 , new_n13881 );
xnor g11535 ( new_n13884 , n1099 , new_n13872 );
nor  g11536 ( new_n13885 , new_n4845 , new_n13884 );
xnor g11537 ( new_n13886 , new_n4845 , new_n13884 );
nor  g11538 ( new_n13887 , new_n3736 , new_n4850_1 );
xnor g11539 ( new_n13888 , new_n3736 , new_n4850_1 );
nor  g11540 ( new_n13889 , new_n3738 , new_n4854 );
xnor g11541 ( new_n13890 , new_n3738 , new_n4854 );
nor  g11542 ( new_n13891 , new_n3742 , new_n4859 );
xnor g11543 ( new_n13892 , new_n3742 , new_n4859 );
nor  g11544 ( new_n13893 , new_n3746 , new_n4864 );
xnor g11545 ( new_n13894 , new_n3746 , new_n4864 );
nor  g11546 ( new_n13895 , new_n3748 , new_n4869 );
xnor g11547 ( new_n13896 , new_n3748 , new_n4880 );
nor  g11548 ( new_n13897 , n25435 , new_n4874 );
and  g11549 ( new_n13898 , new_n3752 , new_n13897 );
nor  g11550 ( new_n13899 , new_n3758_1 , new_n13897 );
nor  g11551 ( new_n13900 , new_n13898 , new_n13899 );
and  g11552 ( new_n13901 , new_n4872 , new_n13900 );
or   g11553 ( new_n13902 , new_n13898 , new_n13901 );
and  g11554 ( new_n13903 , new_n13896 , new_n13902 );
nor  g11555 ( new_n13904 , new_n13895 , new_n13903 );
nor  g11556 ( new_n13905 , new_n13894 , new_n13904 );
nor  g11557 ( new_n13906 , new_n13893 , new_n13905 );
nor  g11558 ( new_n13907 , new_n13892 , new_n13906 );
nor  g11559 ( new_n13908 , new_n13891 , new_n13907 );
nor  g11560 ( new_n13909 , new_n13890 , new_n13908 );
nor  g11561 ( new_n13910 , new_n13889 , new_n13909 );
nor  g11562 ( new_n13911 , new_n13888 , new_n13910 );
nor  g11563 ( new_n13912_1 , new_n13887 , new_n13911 );
nor  g11564 ( new_n13913 , new_n13886 , new_n13912_1 );
nor  g11565 ( new_n13914_1 , new_n13885 , new_n13913 );
nor  g11566 ( new_n13915 , new_n13883 , new_n13914_1 );
nor  g11567 ( new_n13916 , new_n13882 , new_n13915 );
nor  g11568 ( new_n13917 , new_n13880 , new_n13916 );
nor  g11569 ( new_n13918 , new_n13878 , new_n13917 );
not  g11570 ( new_n13919 , new_n4901 );
and  g11571 ( new_n13920 , new_n12671 , new_n13876 );
and  g11572 ( new_n13921 , new_n13919 , new_n13920 );
and  g11573 ( new_n13922_1 , new_n13918 , new_n13921 );
or   g11574 ( new_n13923_1 , new_n13919 , new_n13920 );
nor  g11575 ( new_n13924 , new_n13918 , new_n13923_1 );
nor  g11576 ( new_n13925 , new_n13922_1 , new_n13924 );
and  g11577 ( new_n13926 , new_n13870 , new_n13925 );
or   g11578 ( new_n13927 , new_n13870 , new_n13925 );
xnor g11579 ( new_n13928 , new_n13865 , new_n13868 );
xnor g11580 ( new_n13929 , new_n4901 , new_n13920 );
xnor g11581 ( new_n13930 , new_n13918 , new_n13929 );
nor  g11582 ( new_n13931 , new_n13928 , new_n13930 );
xnor g11583 ( new_n13932 , new_n13928 , new_n13930 );
xnor g11584 ( new_n13933 , new_n13825 , new_n13862 );
xnor g11585 ( new_n13934 , new_n13880 , new_n13916 );
nor  g11586 ( new_n13935 , new_n13933 , new_n13934 );
xnor g11587 ( new_n13936 , new_n13933 , new_n13934 );
xnor g11588 ( new_n13937 , new_n13883 , new_n13914_1 );
xor  g11589 ( new_n13938 , new_n13858 , new_n13860 );
nor  g11590 ( new_n13939 , new_n13937 , new_n13938 );
xnor g11591 ( new_n13940 , new_n13937 , new_n13938 );
xnor g11592 ( new_n13941 , new_n13831 , new_n13856 );
xnor g11593 ( new_n13942 , new_n13886 , new_n13912_1 );
nor  g11594 ( new_n13943 , new_n13941 , new_n13942 );
xnor g11595 ( new_n13944 , new_n13941 , new_n13942 );
xnor g11596 ( new_n13945 , new_n13888 , new_n13910 );
xor  g11597 ( new_n13946 , new_n13833 , new_n13854 );
nor  g11598 ( new_n13947 , new_n13945 , new_n13946 );
xnor g11599 ( new_n13948 , new_n13945 , new_n13946 );
xnor g11600 ( new_n13949 , new_n13890 , new_n13908 );
xor  g11601 ( new_n13950 , new_n13835_1 , new_n13852 );
nor  g11602 ( new_n13951_1 , new_n13949 , new_n13950 );
xnor g11603 ( new_n13952 , new_n13949 , new_n13950 );
xnor g11604 ( new_n13953 , new_n13892 , new_n13906 );
xor  g11605 ( new_n13954 , new_n13837 , new_n13850_1 );
nor  g11606 ( new_n13955 , new_n13953 , new_n13954 );
xnor g11607 ( new_n13956 , new_n13953 , new_n13954 );
xnor g11608 ( new_n13957 , new_n13894 , new_n13904 );
xor  g11609 ( new_n13958 , new_n13839 , new_n13848 );
nor  g11610 ( new_n13959 , new_n13957 , new_n13958 );
xnor g11611 ( new_n13960 , new_n13957 , new_n13958 );
not  g11612 ( new_n13961 , new_n13960 );
xor  g11613 ( new_n13962 , new_n13896 , new_n13902 );
xnor g11614 ( new_n13963 , new_n13845 , new_n13846 );
nor  g11615 ( new_n13964 , new_n13962 , new_n13963 );
xor  g11616 ( new_n13965 , new_n13962 , new_n13963 );
xor  g11617 ( new_n13966 , new_n13842 , new_n13843 );
xnor g11618 ( new_n13967 , new_n4871 , new_n13900 );
and  g11619 ( new_n13968 , new_n13966 , new_n13967 );
xnor g11620 ( new_n13969 , n8581 , new_n9335 );
xnor g11621 ( new_n13970 , n25435 , new_n4874 );
and  g11622 ( new_n13971 , new_n13969 , new_n13970 );
xnor g11623 ( new_n13972 , new_n13966 , new_n13967 );
nor  g11624 ( new_n13973 , new_n13971 , new_n13972 );
nor  g11625 ( new_n13974 , new_n13968 , new_n13973 );
and  g11626 ( new_n13975 , new_n13965 , new_n13974 );
nor  g11627 ( new_n13976 , new_n13964 , new_n13975 );
and  g11628 ( new_n13977 , new_n13961 , new_n13976 );
nor  g11629 ( new_n13978 , new_n13959 , new_n13977 );
nor  g11630 ( new_n13979 , new_n13956 , new_n13978 );
nor  g11631 ( new_n13980 , new_n13955 , new_n13979 );
nor  g11632 ( new_n13981 , new_n13952 , new_n13980 );
nor  g11633 ( new_n13982 , new_n13951_1 , new_n13981 );
nor  g11634 ( new_n13983 , new_n13948 , new_n13982 );
nor  g11635 ( new_n13984 , new_n13947 , new_n13983 );
nor  g11636 ( new_n13985 , new_n13944 , new_n13984 );
nor  g11637 ( new_n13986 , new_n13943 , new_n13985 );
nor  g11638 ( new_n13987 , new_n13940 , new_n13986 );
nor  g11639 ( new_n13988 , new_n13939 , new_n13987 );
nor  g11640 ( new_n13989 , new_n13936 , new_n13988 );
nor  g11641 ( new_n13990 , new_n13935 , new_n13989 );
nor  g11642 ( new_n13991 , new_n13932 , new_n13990 );
nor  g11643 ( new_n13992 , new_n13931 , new_n13991 );
and  g11644 ( new_n13993 , new_n13927 , new_n13992 );
or   g11645 ( new_n13994 , new_n13922_1 , new_n13993 );
nor  g11646 ( n2774 , new_n13926 , new_n13994 );
not  g11647 ( new_n13996 , new_n9395 );
nor  g11648 ( new_n13997 , n20478 , new_n13996 );
not  g11649 ( new_n13998 , new_n13997 );
nor  g11650 ( new_n13999 , n987 , new_n13998 );
not  g11651 ( new_n14000 , new_n13999 );
nor  g11652 ( new_n14001 , n2421 , new_n14000 );
not  g11653 ( new_n14002 , new_n14001 );
nor  g11654 ( new_n14003 , n11044 , new_n14002 );
not  g11655 ( new_n14004_1 , new_n14003 );
nor  g11656 ( new_n14005 , n5031 , new_n14004_1 );
xnor g11657 ( new_n14006 , n2145 , new_n14005 );
xnor g11658 ( new_n14007 , new_n4909 , new_n14006 );
xnor g11659 ( new_n14008 , n5031 , new_n14003 );
nor  g11660 ( new_n14009 , n2659 , new_n14008 );
xnor g11661 ( new_n14010 , new_n4913_1 , new_n14008 );
xnor g11662 ( new_n14011 , n11044 , new_n14001 );
nor  g11663 ( new_n14012 , n24327 , new_n14011 );
xnor g11664 ( new_n14013 , new_n4917 , new_n14011 );
xnor g11665 ( new_n14014 , n2421 , new_n13999 );
nor  g11666 ( new_n14015 , n22198 , new_n14014 );
xnor g11667 ( new_n14016 , n987 , new_n13997 );
and  g11668 ( new_n14017 , n20826 , new_n14016 );
xnor g11669 ( new_n14018 , new_n4927 , new_n14016 );
and  g11670 ( new_n14019 , n7305 , new_n9396_1 );
or   g11671 ( new_n14020 , new_n9399_1 , new_n9407 );
and  g11672 ( new_n14021 , new_n9397 , new_n14020 );
or   g11673 ( new_n14022 , new_n14019 , new_n14021 );
and  g11674 ( new_n14023 , new_n14018 , new_n14022 );
nor  g11675 ( new_n14024 , new_n14017 , new_n14023 );
xnor g11676 ( new_n14025 , new_n4922 , new_n14014 );
and  g11677 ( new_n14026 , new_n14024 , new_n14025 );
or   g11678 ( new_n14027 , new_n14015 , new_n14026 );
and  g11679 ( new_n14028 , new_n14013 , new_n14027 );
or   g11680 ( new_n14029 , new_n14012 , new_n14028 );
and  g11681 ( new_n14030 , new_n14010 , new_n14029 );
nor  g11682 ( new_n14031 , new_n14009 , new_n14030 );
xnor g11683 ( new_n14032 , new_n14007 , new_n14031 );
xnor g11684 ( new_n14033 , new_n3476 , new_n14032 );
nor  g11685 ( new_n14034 , new_n14012 , new_n14028 );
xnor g11686 ( new_n14035 , new_n14010 , new_n14034 );
nor  g11687 ( new_n14036_1 , new_n3480_1 , new_n14035 );
xor  g11688 ( new_n14037 , new_n14013 , new_n14027 );
not  g11689 ( new_n14038 , new_n14037 );
nor  g11690 ( new_n14039 , new_n3486 , new_n14038 );
xnor g11691 ( new_n14040 , new_n3486 , new_n14038 );
xnor g11692 ( new_n14041 , new_n14024 , new_n14025 );
nor  g11693 ( new_n14042 , new_n3491 , new_n14041 );
not  g11694 ( new_n14043 , new_n14041 );
xnor g11695 ( new_n14044 , new_n3490 , new_n14043 );
nor  g11696 ( new_n14045 , new_n14019 , new_n14021 );
xnor g11697 ( new_n14046 , new_n14018 , new_n14045 );
nor  g11698 ( new_n14047 , new_n3495 , new_n14046 );
not  g11699 ( new_n14048 , new_n14046 );
xnor g11700 ( new_n14049 , new_n3495 , new_n14048 );
not  g11701 ( new_n14050 , new_n9409 );
nor  g11702 ( new_n14051 , new_n3500 , new_n14050 );
xnor g11703 ( new_n14052 , new_n3501 , new_n14050 );
nor  g11704 ( new_n14053 , new_n3507 , new_n9428 );
xnor g11705 ( new_n14054 , new_n3509 , new_n9428 );
nor  g11706 ( new_n14055 , new_n3513 , new_n9431 );
nor  g11707 ( new_n14056 , new_n3516_1 , new_n9434 );
not  g11708 ( new_n14057 , new_n9431 );
xnor g11709 ( new_n14058 , new_n3513 , new_n14057 );
and  g11710 ( new_n14059_1 , new_n14056 , new_n14058 );
or   g11711 ( new_n14060 , new_n14055 , new_n14059_1 );
and  g11712 ( new_n14061 , new_n14054 , new_n14060 );
or   g11713 ( new_n14062 , new_n14053 , new_n14061 );
and  g11714 ( new_n14063 , new_n14052 , new_n14062 );
nor  g11715 ( new_n14064 , new_n14051 , new_n14063 );
and  g11716 ( new_n14065 , new_n14049 , new_n14064 );
nor  g11717 ( new_n14066 , new_n14047 , new_n14065 );
nor  g11718 ( new_n14067 , new_n14044 , new_n14066 );
nor  g11719 ( new_n14068 , new_n14042 , new_n14067 );
nor  g11720 ( new_n14069 , new_n14040 , new_n14068 );
nor  g11721 ( new_n14070 , new_n14039 , new_n14069 );
xnor g11722 ( new_n14071_1 , new_n3481 , new_n14035 );
and  g11723 ( new_n14072 , new_n14070 , new_n14071_1 );
nor  g11724 ( new_n14073 , new_n14036_1 , new_n14072 );
xnor g11725 ( new_n14074 , new_n14033 , new_n14073 );
not  g11726 ( new_n14075 , new_n14074 );
xnor g11727 ( new_n14076 , n7026 , new_n3603 );
nor  g11728 ( new_n14077 , new_n3540 , new_n3611 );
or   g11729 ( new_n14078 , n13719 , new_n3608 );
nor  g11730 ( new_n14079 , n442 , new_n3614 );
xnor g11731 ( new_n14080 , new_n3543 , new_n3614 );
nor  g11732 ( new_n14081_1 , n9172 , new_n3618_1 );
xnor g11733 ( new_n14082 , n9172 , new_n3618_1 );
nor  g11734 ( new_n14083 , n4913 , new_n3621 );
xnor g11735 ( new_n14084 , new_n3549 , new_n3621 );
nor  g11736 ( new_n14085 , n604 , new_n3625 );
nor  g11737 ( new_n14086 , n16824 , new_n3629 );
xnor g11738 ( new_n14087 , n16824 , new_n3630 );
nor  g11739 ( new_n14088 , n16521 , new_n3636 );
nand g11740 ( new_n14089 , n7139 , n21993 );
xnor g11741 ( new_n14090_1 , n16521 , new_n3643 );
and  g11742 ( new_n14091 , new_n14089 , new_n14090_1 );
or   g11743 ( new_n14092 , new_n14088 , new_n14091 );
and  g11744 ( new_n14093 , new_n14087 , new_n14092 );
or   g11745 ( new_n14094 , new_n14086 , new_n14093 );
xnor g11746 ( new_n14095_1 , n604 , new_n3626 );
and  g11747 ( new_n14096 , new_n14094 , new_n14095_1 );
or   g11748 ( new_n14097 , new_n14085 , new_n14096 );
and  g11749 ( new_n14098 , new_n14084 , new_n14097 );
nor  g11750 ( new_n14099 , new_n14083 , new_n14098 );
nor  g11751 ( new_n14100 , new_n14082 , new_n14099 );
or   g11752 ( new_n14101 , new_n14081_1 , new_n14100 );
and  g11753 ( new_n14102 , new_n14080 , new_n14101 );
nor  g11754 ( new_n14103 , new_n14079 , new_n14102 );
and  g11755 ( new_n14104 , new_n14078 , new_n14103 );
nor  g11756 ( new_n14105 , new_n14077 , new_n14104 );
xnor g11757 ( new_n14106 , new_n14076 , new_n14105 );
xnor g11758 ( new_n14107_1 , new_n14075 , new_n14106 );
xnor g11759 ( new_n14108 , new_n14070 , new_n14071_1 );
xnor g11760 ( new_n14109 , n13719 , new_n3611 );
xnor g11761 ( new_n14110 , new_n14103 , new_n14109 );
nor  g11762 ( new_n14111 , new_n14108 , new_n14110 );
not  g11763 ( new_n14112 , new_n14108 );
xnor g11764 ( new_n14113 , new_n14112 , new_n14110 );
xor  g11765 ( new_n14114 , new_n14080 , new_n14101 );
xnor g11766 ( new_n14115 , new_n14040 , new_n14068 );
not  g11767 ( new_n14116 , new_n14115 );
and  g11768 ( new_n14117 , new_n14114 , new_n14116 );
xnor g11769 ( new_n14118 , new_n14114 , new_n14116 );
xnor g11770 ( new_n14119 , new_n14082 , new_n14099 );
xnor g11771 ( new_n14120 , new_n14044 , new_n14066 );
nor  g11772 ( new_n14121_1 , new_n14119 , new_n14120 );
not  g11773 ( new_n14122 , new_n14120 );
xnor g11774 ( new_n14123 , new_n14119 , new_n14122 );
xor  g11775 ( new_n14124 , new_n14084 , new_n14097 );
xor  g11776 ( new_n14125 , new_n14049 , new_n14064 );
nor  g11777 ( new_n14126_1 , new_n14124 , new_n14125 );
xor  g11778 ( new_n14127 , new_n14094 , new_n14095_1 );
nor  g11779 ( new_n14128 , new_n14053 , new_n14061 );
xnor g11780 ( new_n14129 , new_n14052 , new_n14128 );
not  g11781 ( new_n14130_1 , new_n14129 );
nor  g11782 ( new_n14131 , new_n14127 , new_n14130_1 );
xnor g11783 ( new_n14132 , new_n14127 , new_n14129 );
xor  g11784 ( new_n14133 , new_n14087 , new_n14092 );
nor  g11785 ( new_n14134 , new_n14055 , new_n14059_1 );
xnor g11786 ( new_n14135 , new_n14054 , new_n14134 );
not  g11787 ( new_n14136_1 , new_n14135 );
nor  g11788 ( new_n14137 , new_n14133 , new_n14136_1 );
xnor g11789 ( new_n14138 , new_n14133 , new_n14135 );
xnor g11790 ( new_n14139 , new_n14056 , new_n14058 );
not  g11791 ( new_n14140 , new_n14139 );
nor  g11792 ( new_n14141 , new_n14090_1 , new_n14140 );
xor  g11793 ( new_n14142 , new_n14089 , new_n14090_1 );
nor  g11794 ( new_n14143 , new_n14139 , new_n14142 );
xnor g11795 ( new_n14144 , n7139 , n21993 );
xnor g11796 ( new_n14145 , new_n3516_1 , new_n9433 );
not  g11797 ( new_n14146 , new_n14145 );
nor  g11798 ( new_n14147_1 , new_n14144 , new_n14146 );
nor  g11799 ( new_n14148_1 , new_n14143 , new_n14147_1 );
nor  g11800 ( new_n14149 , new_n14141 , new_n14148_1 );
and  g11801 ( new_n14150 , new_n14138 , new_n14149 );
or   g11802 ( new_n14151 , new_n14137 , new_n14150 );
and  g11803 ( new_n14152 , new_n14132 , new_n14151 );
nor  g11804 ( new_n14153 , new_n14131 , new_n14152 );
xnor g11805 ( new_n14154 , new_n14124 , new_n14125 );
nor  g11806 ( new_n14155 , new_n14153 , new_n14154 );
nor  g11807 ( new_n14156 , new_n14126_1 , new_n14155 );
and  g11808 ( new_n14157 , new_n14123 , new_n14156 );
nor  g11809 ( new_n14158 , new_n14121_1 , new_n14157 );
nor  g11810 ( new_n14159 , new_n14118 , new_n14158 );
nor  g11811 ( new_n14160 , new_n14117 , new_n14159 );
and  g11812 ( new_n14161 , new_n14113 , new_n14160 );
nor  g11813 ( new_n14162 , new_n14111 , new_n14161 );
xnor g11814 ( n2779 , new_n14107_1 , new_n14162 );
nor  g11815 ( new_n14164 , n25751 , new_n10243 );
not  g11816 ( new_n14165 , n25751 );
xnor g11817 ( new_n14166 , new_n14165 , new_n10243 );
nor  g11818 ( new_n14167 , n26053 , new_n10246 );
not  g11819 ( new_n14168 , n26053 );
xnor g11820 ( new_n14169 , new_n14168 , new_n10246 );
nor  g11821 ( new_n14170 , n7917 , new_n10249 );
not  g11822 ( new_n14171 , n7917 );
xnor g11823 ( new_n14172 , new_n14171 , new_n10249 );
nor  g11824 ( new_n14173 , n17302 , new_n10252 );
not  g11825 ( new_n14174_1 , n17302 );
xnor g11826 ( new_n14175 , new_n14174_1 , new_n10252 );
nor  g11827 ( new_n14176 , n2013 , new_n10254 );
not  g11828 ( new_n14177 , n2013 );
xnor g11829 ( new_n14178 , new_n14177 , new_n10254 );
nor  g11830 ( new_n14179 , n23755 , new_n10257 );
nor  g11831 ( new_n14180 , n19163 , new_n10260 );
not  g11832 ( new_n14181 , n19163 );
xnor g11833 ( new_n14182 , new_n14181 , new_n10260 );
not  g11834 ( new_n14183 , n22358 );
and  g11835 ( new_n14184 , new_n14183 , new_n5811 );
nor  g11836 ( new_n14185 , new_n6585 , new_n3982 );
xnor g11837 ( new_n14186 , new_n14183 , new_n5811 );
nor  g11838 ( new_n14187 , new_n14185 , new_n14186 );
or   g11839 ( new_n14188 , new_n14184 , new_n14187 );
and  g11840 ( new_n14189 , new_n14182 , new_n14188 );
or   g11841 ( new_n14190_1 , new_n14180 , new_n14189 );
not  g11842 ( new_n14191 , n23755 );
xnor g11843 ( new_n14192 , new_n14191 , new_n10257 );
and  g11844 ( new_n14193 , new_n14190_1 , new_n14192 );
or   g11845 ( new_n14194 , new_n14179 , new_n14193 );
and  g11846 ( new_n14195 , new_n14178 , new_n14194 );
or   g11847 ( new_n14196 , new_n14176 , new_n14195 );
and  g11848 ( new_n14197 , new_n14175 , new_n14196 );
or   g11849 ( new_n14198 , new_n14173 , new_n14197 );
and  g11850 ( new_n14199 , new_n14172 , new_n14198 );
or   g11851 ( new_n14200 , new_n14170 , new_n14199 );
and  g11852 ( new_n14201 , new_n14169 , new_n14200 );
or   g11853 ( new_n14202 , new_n14167 , new_n14201 );
and  g11854 ( new_n14203 , new_n14166 , new_n14202 );
nor  g11855 ( new_n14204 , new_n14164 , new_n14203 );
xnor g11856 ( new_n14205 , n25586 , new_n10281 );
xnor g11857 ( new_n14206 , new_n14204 , new_n14205 );
xnor g11858 ( new_n14207 , n4514 , new_n14206 );
xor  g11859 ( new_n14208 , new_n14166 , new_n14202 );
nor  g11860 ( new_n14209 , n3984 , new_n14208 );
xnor g11861 ( new_n14210 , n3984 , new_n14208 );
xor  g11862 ( new_n14211_1 , new_n14169 , new_n14200 );
nor  g11863 ( new_n14212 , n19652 , new_n14211_1 );
xnor g11864 ( new_n14213 , n19652 , new_n14211_1 );
xor  g11865 ( new_n14214 , new_n14172 , new_n14198 );
nor  g11866 ( new_n14215 , n3366 , new_n14214 );
xor  g11867 ( new_n14216 , new_n14175 , new_n14196 );
nor  g11868 ( new_n14217 , n26565 , new_n14216 );
xnor g11869 ( new_n14218 , n26565 , new_n14216 );
xor  g11870 ( new_n14219 , new_n14178 , new_n14194 );
nor  g11871 ( new_n14220 , n3959 , new_n14219 );
xnor g11872 ( new_n14221 , n3959 , new_n14219 );
xor  g11873 ( new_n14222_1 , new_n14190_1 , new_n14192 );
nor  g11874 ( new_n14223 , n11566 , new_n14222_1 );
xnor g11875 ( new_n14224 , n11566 , new_n14222_1 );
xor  g11876 ( new_n14225 , new_n14182 , new_n14188 );
nor  g11877 ( new_n14226 , n26744 , new_n14225 );
xor  g11878 ( new_n14227 , new_n14185 , new_n14186 );
nor  g11879 ( new_n14228 , n26625 , new_n14227 );
nor  g11880 ( new_n14229 , new_n9484 , new_n6586 );
xnor g11881 ( new_n14230_1 , n26625 , new_n14227 );
nor  g11882 ( new_n14231 , new_n14229 , new_n14230_1 );
nor  g11883 ( new_n14232 , new_n14228 , new_n14231 );
xnor g11884 ( new_n14233 , n26744 , new_n14225 );
nor  g11885 ( new_n14234 , new_n14232 , new_n14233 );
nor  g11886 ( new_n14235 , new_n14226 , new_n14234 );
nor  g11887 ( new_n14236 , new_n14224 , new_n14235 );
nor  g11888 ( new_n14237 , new_n14223 , new_n14236 );
nor  g11889 ( new_n14238 , new_n14221 , new_n14237 );
nor  g11890 ( new_n14239 , new_n14220 , new_n14238 );
nor  g11891 ( new_n14240 , new_n14218 , new_n14239 );
nor  g11892 ( new_n14241 , new_n14217 , new_n14240 );
xnor g11893 ( new_n14242 , n3366 , new_n14214 );
nor  g11894 ( new_n14243 , new_n14241 , new_n14242 );
nor  g11895 ( new_n14244 , new_n14215 , new_n14243 );
nor  g11896 ( new_n14245 , new_n14213 , new_n14244 );
nor  g11897 ( new_n14246 , new_n14212 , new_n14245 );
nor  g11898 ( new_n14247 , new_n14210 , new_n14246 );
nor  g11899 ( new_n14248 , new_n14209 , new_n14247 );
xnor g11900 ( new_n14249 , new_n14207 , new_n14248 );
and  g11901 ( new_n14250 , new_n10354 , new_n14249 );
xnor g11902 ( new_n14251 , new_n10354 , new_n14249 );
xor  g11903 ( new_n14252 , new_n14210 , new_n14246 );
nor  g11904 ( new_n14253 , new_n10359 , new_n14252 );
xnor g11905 ( new_n14254 , new_n10359 , new_n14252 );
xor  g11906 ( new_n14255 , new_n14213 , new_n14244 );
nor  g11907 ( new_n14256 , new_n10362 , new_n14255 );
xnor g11908 ( new_n14257 , new_n10362 , new_n14255 );
xor  g11909 ( new_n14258 , new_n14241 , new_n14242 );
nor  g11910 ( new_n14259 , new_n10367 , new_n14258 );
xnor g11911 ( new_n14260 , new_n10367 , new_n14258 );
xor  g11912 ( new_n14261 , new_n14218 , new_n14239 );
nor  g11913 ( new_n14262 , new_n10370 , new_n14261 );
xnor g11914 ( new_n14263 , new_n10370 , new_n14261 );
xor  g11915 ( new_n14264 , new_n14221 , new_n14237 );
nor  g11916 ( new_n14265 , new_n10375 , new_n14264 );
xnor g11917 ( new_n14266 , new_n10375 , new_n14264 );
xor  g11918 ( new_n14267_1 , new_n14224 , new_n14235 );
nor  g11919 ( new_n14268 , new_n10379 , new_n14267_1 );
xnor g11920 ( new_n14269 , new_n10379 , new_n14267_1 );
xor  g11921 ( new_n14270 , new_n14232 , new_n14233 );
nor  g11922 ( new_n14271_1 , new_n10384 , new_n14270 );
xnor g11923 ( new_n14272 , new_n10384 , new_n14270 );
xnor g11924 ( new_n14273 , new_n14229 , new_n14230_1 );
not  g11925 ( new_n14274 , new_n14273 );
nor  g11926 ( new_n14275_1 , new_n5808 , new_n14274 );
nor  g11927 ( new_n14276 , new_n5803 , new_n6587_1 );
nor  g11928 ( new_n14277_1 , new_n5809 , new_n14273 );
nor  g11929 ( new_n14278 , new_n14276 , new_n14277_1 );
nor  g11930 ( new_n14279 , new_n14275_1 , new_n14278 );
nor  g11931 ( new_n14280 , new_n14272 , new_n14279 );
nor  g11932 ( new_n14281 , new_n14271_1 , new_n14280 );
nor  g11933 ( new_n14282 , new_n14269 , new_n14281 );
nor  g11934 ( new_n14283 , new_n14268 , new_n14282 );
nor  g11935 ( new_n14284 , new_n14266 , new_n14283 );
nor  g11936 ( new_n14285 , new_n14265 , new_n14284 );
nor  g11937 ( new_n14286 , new_n14263 , new_n14285 );
nor  g11938 ( new_n14287 , new_n14262 , new_n14286 );
nor  g11939 ( new_n14288 , new_n14260 , new_n14287 );
nor  g11940 ( new_n14289 , new_n14259 , new_n14288 );
nor  g11941 ( new_n14290 , new_n14257 , new_n14289 );
nor  g11942 ( new_n14291 , new_n14256 , new_n14290 );
nor  g11943 ( new_n14292 , new_n14254 , new_n14291 );
nor  g11944 ( new_n14293 , new_n14253 , new_n14292 );
nor  g11945 ( new_n14294_1 , new_n14251 , new_n14293 );
nor  g11946 ( new_n14295 , new_n14250 , new_n14294_1 );
xnor g11947 ( new_n14296 , new_n10352 , new_n14295 );
and  g11948 ( new_n14297 , n4514 , new_n14206 );
not  g11949 ( new_n14298 , new_n14248 );
nor  g11950 ( new_n14299 , new_n14207 , new_n14298 );
or   g11951 ( new_n14300 , new_n14297 , new_n14299 );
or   g11952 ( new_n14301 , n25586 , new_n10241 );
and  g11953 ( new_n14302 , new_n14204 , new_n14301 );
not  g11954 ( new_n14303 , n25586 );
nor  g11955 ( new_n14304 , new_n14303 , new_n10281 );
or   g11956 ( new_n14305 , new_n10240 , new_n14304 );
nor  g11957 ( new_n14306 , new_n14302 , new_n14305 );
xnor g11958 ( new_n14307 , new_n14300 , new_n14306 );
xnor g11959 ( n2826 , new_n14296 , new_n14307 );
nor  g11960 ( new_n14309 , new_n12110 , new_n6244 );
xnor g11961 ( new_n14310_1 , n5140 , new_n6244 );
nor  g11962 ( new_n14311 , new_n12113_1 , new_n6250 );
xnor g11963 ( new_n14312 , new_n12113_1 , new_n6251 );
nor  g11964 ( new_n14313 , new_n12116 , new_n6256_1 );
xnor g11965 ( new_n14314 , new_n12116 , new_n6257 );
nor  g11966 ( new_n14315 , new_n12119 , new_n6262 );
xnor g11967 ( new_n14316 , new_n12119 , new_n6304 );
nor  g11968 ( new_n14317 , new_n12122 , new_n6268 );
nor  g11969 ( new_n14318 , n8244 , new_n6274 );
xnor g11970 ( new_n14319 , new_n12125 , new_n6274 );
nor  g11971 ( new_n14320 , new_n12128 , new_n6276_1 );
xnor g11972 ( new_n14321 , new_n12128 , new_n6277 );
nor  g11973 ( new_n14322 , n15167 , new_n6282 );
nor  g11974 ( new_n14323_1 , new_n12134 , new_n6285 );
nor  g11975 ( new_n14324 , new_n6492 , new_n6288 );
xnor g11976 ( new_n14325 , new_n12134 , new_n12226 );
and  g11977 ( new_n14326_1 , new_n14324 , new_n14325 );
nor  g11978 ( new_n14327 , new_n14323_1 , new_n14326_1 );
xnor g11979 ( new_n14328 , new_n12132 , new_n6282 );
and  g11980 ( new_n14329 , new_n14327 , new_n14328 );
nor  g11981 ( new_n14330 , new_n14322 , new_n14329 );
and  g11982 ( new_n14331 , new_n14321 , new_n14330 );
nor  g11983 ( new_n14332 , new_n14320 , new_n14331 );
and  g11984 ( new_n14333 , new_n14319 , new_n14332 );
nor  g11985 ( new_n14334 , new_n14318 , new_n14333 );
xnor g11986 ( new_n14335 , new_n12122 , new_n6269 );
and  g11987 ( new_n14336 , new_n14334 , new_n14335 );
or   g11988 ( new_n14337 , new_n14317 , new_n14336 );
and  g11989 ( new_n14338 , new_n14316 , new_n14337 );
or   g11990 ( new_n14339 , new_n14315 , new_n14338 );
and  g11991 ( new_n14340 , new_n14314 , new_n14339 );
or   g11992 ( new_n14341 , new_n14313 , new_n14340 );
and  g11993 ( new_n14342_1 , new_n14312 , new_n14341 );
or   g11994 ( new_n14343 , new_n14311 , new_n14342_1 );
and  g11995 ( new_n14344 , new_n14310_1 , new_n14343 );
nor  g11996 ( new_n14345_1 , new_n14309 , new_n14344 );
nor  g11997 ( new_n14346 , new_n6242 , new_n14345_1 );
not  g11998 ( new_n14347 , n25365 );
nor  g11999 ( new_n14348 , new_n14347 , new_n2603 );
or   g12000 ( new_n14349 , new_n2606 , new_n2653 );
and  g12001 ( new_n14350 , new_n2604 , new_n14349 );
nor  g12002 ( new_n14351 , new_n14348 , new_n14350 );
nor  g12003 ( new_n14352 , n9396 , n20040 );
nor  g12004 ( new_n14353_1 , new_n2556 , new_n2601 );
nor  g12005 ( new_n14354 , new_n14352 , new_n14353_1 );
not  g12006 ( new_n14355 , new_n14354 );
nor  g12007 ( new_n14356 , new_n14351 , new_n14355 );
not  g12008 ( new_n14357 , new_n14356 );
xnor g12009 ( new_n14358 , new_n14346 , new_n14357 );
xnor g12010 ( new_n14359 , new_n6197 , new_n14345_1 );
not  g12011 ( new_n14360 , new_n14359 );
xnor g12012 ( new_n14361 , new_n14351 , new_n14354 );
and  g12013 ( new_n14362 , new_n14360 , new_n14361 );
xnor g12014 ( new_n14363 , new_n14360 , new_n14361 );
xor  g12015 ( new_n14364_1 , new_n14310_1 , new_n14343 );
nor  g12016 ( new_n14365 , new_n2656 , new_n14364_1 );
xnor g12017 ( new_n14366 , new_n2656 , new_n14364_1 );
xor  g12018 ( new_n14367 , new_n14312 , new_n14341 );
nor  g12019 ( new_n14368 , new_n2787 , new_n14367 );
xnor g12020 ( new_n14369 , new_n2787 , new_n14367 );
not  g12021 ( new_n14370 , new_n2792 );
xor  g12022 ( new_n14371 , new_n14314 , new_n14339 );
nor  g12023 ( new_n14372 , new_n14370 , new_n14371 );
xnor g12024 ( new_n14373 , new_n14370 , new_n14371 );
xor  g12025 ( new_n14374 , new_n14316 , new_n14337 );
nor  g12026 ( new_n14375_1 , new_n2796 , new_n14374 );
xnor g12027 ( new_n14376 , new_n2796 , new_n14374 );
xor  g12028 ( new_n14377 , new_n14334 , new_n14335 );
nor  g12029 ( new_n14378 , new_n2802 , new_n14377 );
xnor g12030 ( new_n14379 , new_n2802 , new_n14377 );
xnor g12031 ( new_n14380 , new_n14319 , new_n14332 );
nor  g12032 ( new_n14381 , new_n2806 , new_n14380 );
xnor g12033 ( new_n14382 , new_n2806 , new_n14380 );
xor  g12034 ( new_n14383 , new_n14321 , new_n14330 );
nor  g12035 ( new_n14384 , new_n2814 , new_n14383 );
xnor g12036 ( new_n14385 , new_n2814 , new_n14383 );
xnor g12037 ( new_n14386 , new_n14327 , new_n14328 );
nor  g12038 ( new_n14387 , new_n2817 , new_n14386 );
xnor g12039 ( new_n14388 , new_n2817 , new_n14386 );
xor  g12040 ( new_n14389 , new_n14324 , new_n14325 );
nor  g12041 ( new_n14390 , new_n2823 , new_n14389 );
xnor g12042 ( new_n14391 , n8656 , new_n6288 );
nor  g12043 ( new_n14392 , new_n2827 , new_n14391 );
xnor g12044 ( new_n14393 , new_n2824 , new_n14389 );
and  g12045 ( new_n14394 , new_n14392 , new_n14393 );
nor  g12046 ( new_n14395 , new_n14390 , new_n14394 );
nor  g12047 ( new_n14396 , new_n14388 , new_n14395 );
nor  g12048 ( new_n14397 , new_n14387 , new_n14396 );
nor  g12049 ( new_n14398 , new_n14385 , new_n14397 );
nor  g12050 ( new_n14399 , new_n14384 , new_n14398 );
nor  g12051 ( new_n14400 , new_n14382 , new_n14399 );
nor  g12052 ( new_n14401 , new_n14381 , new_n14400 );
nor  g12053 ( new_n14402 , new_n14379 , new_n14401 );
nor  g12054 ( new_n14403 , new_n14378 , new_n14402 );
nor  g12055 ( new_n14404 , new_n14376 , new_n14403 );
nor  g12056 ( new_n14405 , new_n14375_1 , new_n14404 );
nor  g12057 ( new_n14406 , new_n14373 , new_n14405 );
nor  g12058 ( new_n14407 , new_n14372 , new_n14406 );
nor  g12059 ( new_n14408 , new_n14369 , new_n14407 );
nor  g12060 ( new_n14409 , new_n14368 , new_n14408 );
nor  g12061 ( new_n14410 , new_n14366 , new_n14409 );
nor  g12062 ( new_n14411 , new_n14365 , new_n14410 );
nor  g12063 ( new_n14412_1 , new_n14363 , new_n14411 );
nor  g12064 ( new_n14413 , new_n14362 , new_n14412_1 );
xnor g12065 ( n2853 , new_n14358 , new_n14413 );
xnor g12066 ( new_n14415 , n2035 , n7099 );
nor  g12067 ( new_n14416 , n5213 , new_n11685 );
xnor g12068 ( new_n14417 , n5213 , n12811 );
nor  g12069 ( new_n14418 , new_n11689 , n4665 );
xnor g12070 ( new_n14419 , n1118 , n4665 );
nor  g12071 ( new_n14420 , new_n2866 , n25974 );
nor  g12072 ( new_n14421 , n19005 , new_n11693 );
nor  g12073 ( new_n14422 , n1630 , new_n2869 );
nor  g12074 ( new_n14423 , new_n2909 , n4326 );
nor  g12075 ( new_n14424 , n1451 , new_n5287 );
not  g12076 ( new_n14425 , new_n14424 );
nor  g12077 ( new_n14426 , new_n14423 , new_n14425 );
nor  g12078 ( new_n14427 , new_n14422 , new_n14426 );
nor  g12079 ( new_n14428 , new_n14421 , new_n14427 );
nor  g12080 ( new_n14429 , new_n14420 , new_n14428 );
and  g12081 ( new_n14430 , new_n14419 , new_n14429 );
or   g12082 ( new_n14431 , new_n14418 , new_n14430 );
and  g12083 ( new_n14432 , new_n14417 , new_n14431 );
or   g12084 ( new_n14433 , new_n14416 , new_n14432 );
xor  g12085 ( new_n14434 , new_n14415 , new_n14433 );
not  g12086 ( new_n14435 , n5337 );
not  g12087 ( new_n14436 , new_n4228 );
nor  g12088 ( new_n14437 , n13668 , new_n14436 );
xnor g12089 ( new_n14438 , n3570 , new_n14437 );
xnor g12090 ( new_n14439 , new_n14435 , new_n14438 );
and  g12091 ( new_n14440_1 , n626 , new_n4229 );
or   g12092 ( new_n14441 , new_n4232 , new_n4249 );
and  g12093 ( new_n14442 , new_n4230 , new_n14441 );
nor  g12094 ( new_n14443 , new_n14440_1 , new_n14442 );
xnor g12095 ( new_n14444 , new_n14439 , new_n14443 );
not  g12096 ( new_n14445 , new_n14444 );
xnor g12097 ( new_n14446 , new_n10979 , new_n14445 );
not  g12098 ( new_n14447 , new_n4251 );
nor  g12099 ( new_n14448 , new_n4222 , new_n14447 );
and  g12100 ( new_n14449 , new_n4252 , new_n4282 );
nor  g12101 ( new_n14450 , new_n14448 , new_n14449 );
xnor g12102 ( new_n14451 , new_n14446 , new_n14450 );
not  g12103 ( new_n14452 , new_n14451 );
xnor g12104 ( new_n14453 , new_n14434 , new_n14452 );
xor  g12105 ( new_n14454 , new_n14417 , new_n14431 );
nor  g12106 ( new_n14455 , new_n4283 , new_n14454 );
xnor g12107 ( new_n14456 , new_n14419 , new_n14429 );
and  g12108 ( new_n14457_1 , new_n4287 , new_n14456 );
xnor g12109 ( new_n14458 , new_n4287 , new_n14456 );
xnor g12110 ( new_n14459 , n19005 , n25974 );
xnor g12111 ( new_n14460 , new_n14427 , new_n14459 );
and  g12112 ( new_n14461 , new_n4292 , new_n14460 );
xnor g12113 ( new_n14462 , new_n4291 , new_n14460 );
xnor g12114 ( new_n14463 , n1451 , n5438 );
nor  g12115 ( new_n14464_1 , new_n4303 , new_n14463 );
xnor g12116 ( new_n14465 , n1630 , n4326 );
xnor g12117 ( new_n14466 , new_n14425 , new_n14465 );
not  g12118 ( new_n14467 , new_n14466 );
and  g12119 ( new_n14468 , new_n14464_1 , new_n14467 );
xnor g12120 ( new_n14469 , new_n14464_1 , new_n14467 );
nor  g12121 ( new_n14470 , new_n4296 , new_n14469 );
nor  g12122 ( new_n14471_1 , new_n14468 , new_n14470 );
and  g12123 ( new_n14472 , new_n14462 , new_n14471_1 );
nor  g12124 ( new_n14473 , new_n14461 , new_n14472 );
nor  g12125 ( new_n14474 , new_n14458 , new_n14473 );
nor  g12126 ( new_n14475_1 , new_n14457_1 , new_n14474 );
xnor g12127 ( new_n14476 , new_n4283 , new_n14454 );
nor  g12128 ( new_n14477 , new_n14475_1 , new_n14476 );
nor  g12129 ( new_n14478 , new_n14455 , new_n14477 );
xor  g12130 ( n2860 , new_n14453 , new_n14478 );
xnor g12131 ( n2887 , new_n13568 , new_n13586 );
not  g12132 ( new_n14481 , new_n14437 );
nor  g12133 ( new_n14482 , n3570 , new_n14481 );
not  g12134 ( new_n14483 , new_n14482 );
nor  g12135 ( new_n14484 , n4409 , new_n14483 );
not  g12136 ( new_n14485 , new_n14484 );
nor  g12137 ( new_n14486 , n20359 , new_n14485 );
and  g12138 ( new_n14487 , new_n6025 , new_n14486 );
xnor g12139 ( new_n14488 , n8526 , new_n14487 );
nor  g12140 ( new_n14489 , n21784 , new_n14488 );
xnor g12141 ( new_n14490 , n2816 , new_n14486 );
and  g12142 ( new_n14491 , n5521 , new_n14490 );
or   g12143 ( new_n14492 , n5521 , new_n14490 );
xnor g12144 ( new_n14493 , n20359 , new_n14484 );
nor  g12145 ( new_n14494 , n11926 , new_n14493 );
xnor g12146 ( new_n14495 , n11926 , new_n14493 );
xnor g12147 ( new_n14496 , n4409 , new_n14482 );
and  g12148 ( new_n14497 , n4325 , new_n14496 );
nor  g12149 ( new_n14498 , n4325 , new_n14496 );
and  g12150 ( new_n14499 , n5337 , new_n14438 );
nor  g12151 ( new_n14500 , n5337 , new_n14438 );
nor  g12152 ( new_n14501 , new_n14500 , new_n14443 );
nor  g12153 ( new_n14502 , new_n14499 , new_n14501 );
nor  g12154 ( new_n14503 , new_n14498 , new_n14502 );
or   g12155 ( new_n14504 , new_n14497 , new_n14503 );
nor  g12156 ( new_n14505 , new_n14495 , new_n14504 );
nor  g12157 ( new_n14506 , new_n14494 , new_n14505 );
and  g12158 ( new_n14507 , new_n14492 , new_n14506 );
nor  g12159 ( new_n14508 , new_n14491 , new_n14507 );
nor  g12160 ( new_n14509 , new_n14489 , new_n14508 );
and  g12161 ( new_n14510_1 , new_n5981 , new_n14487 );
and  g12162 ( new_n14511 , n21784 , new_n14488 );
or   g12163 ( new_n14512 , new_n14510_1 , new_n14511 );
nor  g12164 ( new_n14513 , new_n14509 , new_n14512 );
not  g12165 ( new_n14514 , new_n14513 );
xnor g12166 ( new_n14515 , new_n10955 , new_n14514 );
not  g12167 ( new_n14516 , n21784 );
xnor g12168 ( new_n14517 , new_n14516 , new_n14488 );
xnor g12169 ( new_n14518 , new_n14508 , new_n14517 );
and  g12170 ( new_n14519 , new_n10961_1 , new_n14518 );
xnor g12171 ( new_n14520 , new_n10960 , new_n14518 );
xnor g12172 ( new_n14521 , n5521 , new_n14490 );
xnor g12173 ( new_n14522 , new_n14506 , new_n14521 );
nor  g12174 ( new_n14523 , new_n10965 , new_n14522 );
xnor g12175 ( new_n14524 , new_n10965 , new_n14522 );
nor  g12176 ( new_n14525 , new_n14497 , new_n14503 );
xnor g12177 ( new_n14526 , new_n14495 , new_n14525 );
and  g12178 ( new_n14527 , new_n10969 , new_n14526 );
xnor g12179 ( new_n14528 , new_n5991 , new_n14496 );
xnor g12180 ( new_n14529 , new_n14502 , new_n14528 );
and  g12181 ( new_n14530 , new_n10974 , new_n14529 );
xnor g12182 ( new_n14531 , new_n10974 , new_n14529 );
and  g12183 ( new_n14532 , new_n10979 , new_n14444 );
or   g12184 ( new_n14533 , new_n14448 , new_n14449 );
and  g12185 ( new_n14534 , new_n14446 , new_n14533 );
nor  g12186 ( new_n14535 , new_n14532 , new_n14534 );
nor  g12187 ( new_n14536 , new_n14531 , new_n14535 );
nor  g12188 ( new_n14537 , new_n14530 , new_n14536 );
xnor g12189 ( new_n14538 , new_n10970 , new_n14526 );
and  g12190 ( new_n14539 , new_n14537 , new_n14538 );
nor  g12191 ( new_n14540 , new_n14527 , new_n14539 );
nor  g12192 ( new_n14541_1 , new_n14524 , new_n14540 );
nor  g12193 ( new_n14542 , new_n14523 , new_n14541_1 );
and  g12194 ( new_n14543 , new_n14520 , new_n14542 );
nor  g12195 ( new_n14544 , new_n14519 , new_n14543 );
xnor g12196 ( new_n14545 , new_n14515 , new_n14544 );
not  g12197 ( new_n14546_1 , new_n14545 );
not  g12198 ( new_n14547_1 , n8827 );
not  g12199 ( new_n14548 , new_n4170 );
nor  g12200 ( new_n14549 , n19905 , new_n14548 );
not  g12201 ( new_n14550 , new_n14549 );
nor  g12202 ( new_n14551 , n26452 , new_n14550 );
not  g12203 ( new_n14552 , new_n14551 );
nor  g12204 ( new_n14553 , n15546 , new_n14552 );
not  g12205 ( new_n14554 , new_n14553 );
nor  g12206 ( new_n14555 , n5077 , new_n14554 );
and  g12207 ( new_n14556 , new_n12683 , new_n14555 );
and  g12208 ( new_n14557 , new_n14547_1 , new_n14556 );
xnor g12209 ( new_n14558 , n8827 , new_n14556 );
nor  g12210 ( new_n14559 , n11898 , new_n14558 );
xnor g12211 ( new_n14560 , n18035 , new_n14555 );
nor  g12212 ( new_n14561 , n19941 , new_n14560 );
xnor g12213 ( new_n14562 , new_n12673 , new_n14560 );
xnor g12214 ( new_n14563 , n5077 , new_n14553 );
nor  g12215 ( new_n14564 , n1099 , new_n14563 );
xnor g12216 ( new_n14565 , n1099 , new_n14563 );
xnor g12217 ( new_n14566 , n15546 , new_n14551 );
nor  g12218 ( new_n14567 , n2113 , new_n14566 );
xnor g12219 ( new_n14568 , n26452 , new_n14549 );
nor  g12220 ( new_n14569 , n21134 , new_n14568 );
xnor g12221 ( new_n14570_1 , n21134 , new_n14568 );
nor  g12222 ( new_n14571 , n6369 , new_n4171 );
and  g12223 ( new_n14572 , new_n4172_1 , new_n4193 );
nor  g12224 ( new_n14573 , new_n14571 , new_n14572 );
nor  g12225 ( new_n14574 , new_n14570_1 , new_n14573 );
or   g12226 ( new_n14575_1 , new_n14569 , new_n14574 );
xnor g12227 ( new_n14576_1 , new_n10434 , new_n14566 );
and  g12228 ( new_n14577 , new_n14575_1 , new_n14576_1 );
nor  g12229 ( new_n14578 , new_n14567 , new_n14577 );
nor  g12230 ( new_n14579 , new_n14565 , new_n14578 );
or   g12231 ( new_n14580 , new_n14564 , new_n14579 );
and  g12232 ( new_n14581 , new_n14562 , new_n14580 );
nor  g12233 ( new_n14582 , new_n14561 , new_n14581 );
and  g12234 ( new_n14583 , n11898 , new_n14558 );
nor  g12235 ( new_n14584 , new_n14582 , new_n14583 );
nor  g12236 ( new_n14585 , new_n14559 , new_n14584 );
nor  g12237 ( new_n14586 , new_n14557 , new_n14585 );
xnor g12238 ( new_n14587 , new_n14546_1 , new_n14586 );
xnor g12239 ( new_n14588 , new_n14520 , new_n14542 );
not  g12240 ( new_n14589 , new_n14588 );
xnor g12241 ( new_n14590 , new_n12671 , new_n14558 );
xnor g12242 ( new_n14591 , new_n14582 , new_n14590 );
not  g12243 ( new_n14592 , new_n14591 );
nor  g12244 ( new_n14593_1 , new_n14589 , new_n14592 );
xnor g12245 ( new_n14594 , new_n14589 , new_n14592 );
xor  g12246 ( new_n14595 , new_n14562 , new_n14580 );
not  g12247 ( new_n14596 , new_n14595 );
xnor g12248 ( new_n14597 , new_n14524 , new_n14540 );
nor  g12249 ( new_n14598 , new_n14596 , new_n14597 );
xnor g12250 ( new_n14599 , new_n14596 , new_n14597 );
xnor g12251 ( new_n14600 , new_n14565 , new_n14578 );
xnor g12252 ( new_n14601 , new_n14537 , new_n14538 );
nor  g12253 ( new_n14602 , new_n14600 , new_n14601 );
not  g12254 ( new_n14603_1 , new_n14600 );
not  g12255 ( new_n14604 , new_n14601 );
xnor g12256 ( new_n14605 , new_n14603_1 , new_n14604 );
xnor g12257 ( new_n14606 , new_n14531 , new_n14535 );
xor  g12258 ( new_n14607 , new_n14575_1 , new_n14576_1 );
and  g12259 ( new_n14608 , new_n14606 , new_n14607 );
xnor g12260 ( new_n14609 , new_n14606 , new_n14607 );
xnor g12261 ( new_n14610 , new_n14570_1 , new_n14573 );
nor  g12262 ( new_n14611 , new_n14451 , new_n14610 );
not  g12263 ( new_n14612 , new_n14610 );
xnor g12264 ( new_n14613 , new_n14452 , new_n14612 );
nor  g12265 ( new_n14614 , new_n4194 , new_n4283 );
and  g12266 ( new_n14615 , new_n4284 , new_n4310 );
nor  g12267 ( new_n14616 , new_n14614 , new_n14615 );
nor  g12268 ( new_n14617 , new_n14613 , new_n14616 );
nor  g12269 ( new_n14618 , new_n14611 , new_n14617 );
nor  g12270 ( new_n14619 , new_n14609 , new_n14618 );
nor  g12271 ( new_n14620 , new_n14608 , new_n14619 );
nor  g12272 ( new_n14621 , new_n14605 , new_n14620 );
nor  g12273 ( new_n14622 , new_n14602 , new_n14621 );
nor  g12274 ( new_n14623 , new_n14599 , new_n14622 );
nor  g12275 ( new_n14624 , new_n14598 , new_n14623 );
nor  g12276 ( new_n14625 , new_n14594 , new_n14624 );
nor  g12277 ( new_n14626 , new_n14593_1 , new_n14625 );
xor  g12278 ( n2929 , new_n14587 , new_n14626 );
not  g12279 ( new_n14628 , new_n7269 );
xnor g12280 ( new_n14629 , n767 , n22793 );
not  g12281 ( new_n14630 , n7330 );
nor  g12282 ( new_n14631 , new_n14630 , n8439 );
xnor g12283 ( new_n14632 , n7330 , n8439 );
nor  g12284 ( new_n14633_1 , new_n2683 , n25523 );
xnor g12285 ( new_n14634 , n22492 , n25523 );
not  g12286 ( new_n14635 , n12821 );
nor  g12287 ( new_n14636_1 , n5579 , new_n14635 );
xnor g12288 ( new_n14637 , n5579 , n12821 );
nor  g12289 ( new_n14638 , new_n2689 , n23430 );
xnor g12290 ( new_n14639 , n3468 , n23430 );
not  g12291 ( new_n14640 , n10411 );
nor  g12292 ( new_n14641 , new_n14640 , n18558 );
and  g12293 ( new_n14642 , new_n13313 , new_n13323 );
nor  g12294 ( new_n14643 , new_n14641 , new_n14642 );
and  g12295 ( new_n14644 , new_n14639 , new_n14643 );
or   g12296 ( new_n14645 , new_n14638 , new_n14644 );
and  g12297 ( new_n14646 , new_n14637 , new_n14645 );
or   g12298 ( new_n14647 , new_n14636_1 , new_n14646 );
and  g12299 ( new_n14648 , new_n14634 , new_n14647 );
or   g12300 ( new_n14649 , new_n14633_1 , new_n14648 );
and  g12301 ( new_n14650 , new_n14632 , new_n14649 );
nor  g12302 ( new_n14651 , new_n14631 , new_n14650 );
xnor g12303 ( new_n14652 , new_n14629 , new_n14651 );
not  g12304 ( new_n14653 , new_n14652 );
xnor g12305 ( new_n14654 , new_n14628 , new_n14653 );
xor  g12306 ( new_n14655 , new_n14632 , new_n14649 );
and  g12307 ( new_n14656 , new_n7274 , new_n14655 );
not  g12308 ( new_n14657 , new_n7274 );
xnor g12309 ( new_n14658 , new_n14657 , new_n14655 );
xor  g12310 ( new_n14659 , new_n14634 , new_n14647 );
nor  g12311 ( new_n14660 , new_n7278 , new_n14659 );
xnor g12312 ( new_n14661 , new_n7278 , new_n14659 );
xor  g12313 ( new_n14662 , new_n14637 , new_n14645 );
nor  g12314 ( new_n14663 , new_n7282 , new_n14662 );
xnor g12315 ( new_n14664 , new_n11953 , new_n14662 );
xnor g12316 ( new_n14665 , new_n14639 , new_n14643 );
not  g12317 ( new_n14666 , new_n14665 );
and  g12318 ( new_n14667 , new_n7285 , new_n14666 );
xnor g12319 ( new_n14668 , new_n7285 , new_n14665 );
nor  g12320 ( new_n14669 , new_n7290 , new_n13324 );
or   g12321 ( new_n14670 , new_n13599 , new_n13606 );
and  g12322 ( new_n14671 , new_n13598 , new_n14670 );
or   g12323 ( new_n14672 , new_n14669 , new_n14671 );
and  g12324 ( new_n14673 , new_n14668 , new_n14672 );
nor  g12325 ( new_n14674 , new_n14667 , new_n14673 );
and  g12326 ( new_n14675 , new_n14664 , new_n14674 );
nor  g12327 ( new_n14676 , new_n14663 , new_n14675 );
nor  g12328 ( new_n14677 , new_n14661 , new_n14676 );
nor  g12329 ( new_n14678 , new_n14660 , new_n14677 );
and  g12330 ( new_n14679 , new_n14658 , new_n14678 );
nor  g12331 ( new_n14680_1 , new_n14656 , new_n14679 );
xnor g12332 ( new_n14681 , new_n14654 , new_n14680_1 );
not  g12333 ( new_n14682 , new_n14681 );
xnor g12334 ( new_n14683 , n15077 , n22379 );
nor  g12335 ( new_n14684_1 , new_n2850 , n3710 );
xnor g12336 ( new_n14685 , n1662 , n3710 );
nor  g12337 ( new_n14686 , new_n2853_1 , n26318 );
xnor g12338 ( new_n14687 , n12875 , n26318 );
nor  g12339 ( new_n14688 , new_n2856 , n26054 );
xnor g12340 ( new_n14689 , n2035 , n26054 );
nor  g12341 ( new_n14690 , new_n2859 , n19081 );
or   g12342 ( new_n14691 , n5213 , new_n8753 );
nor  g12343 ( new_n14692_1 , n4665 , new_n8771 );
and  g12344 ( new_n14693 , new_n13610 , new_n13619 );
nor  g12345 ( new_n14694 , new_n14692_1 , new_n14693 );
and  g12346 ( new_n14695 , new_n14691 , new_n14694 );
or   g12347 ( new_n14696 , new_n14690 , new_n14695 );
and  g12348 ( new_n14697 , new_n14689 , new_n14696 );
or   g12349 ( new_n14698 , new_n14688 , new_n14697 );
and  g12350 ( new_n14699 , new_n14687 , new_n14698 );
or   g12351 ( new_n14700 , new_n14686 , new_n14699 );
and  g12352 ( new_n14701_1 , new_n14685 , new_n14700 );
or   g12353 ( new_n14702_1 , new_n14684_1 , new_n14701_1 );
xor  g12354 ( new_n14703 , new_n14683 , new_n14702_1 );
xnor g12355 ( new_n14704_1 , new_n14682 , new_n14703 );
xor  g12356 ( new_n14705 , new_n14685 , new_n14700 );
xor  g12357 ( new_n14706 , new_n14658 , new_n14678 );
nor  g12358 ( new_n14707 , new_n14705 , new_n14706 );
xnor g12359 ( new_n14708 , new_n14705 , new_n14706 );
xor  g12360 ( new_n14709 , new_n14687 , new_n14698 );
xnor g12361 ( new_n14710 , new_n14661 , new_n14676 );
nor  g12362 ( new_n14711 , new_n14709 , new_n14710 );
xnor g12363 ( new_n14712 , new_n14709 , new_n14710 );
xor  g12364 ( new_n14713 , new_n14689 , new_n14696 );
xnor g12365 ( new_n14714 , new_n14664 , new_n14674 );
nor  g12366 ( new_n14715 , new_n14713 , new_n14714 );
nor  g12367 ( new_n14716 , new_n14669 , new_n14671 );
xnor g12368 ( new_n14717 , new_n14668 , new_n14716 );
not  g12369 ( new_n14718 , new_n14717 );
xnor g12370 ( new_n14719 , n5213 , n19081 );
xnor g12371 ( new_n14720 , new_n14694 , new_n14719 );
and  g12372 ( new_n14721 , new_n14718 , new_n14720 );
xnor g12373 ( new_n14722 , new_n14718 , new_n14720 );
and  g12374 ( new_n14723 , new_n13609 , new_n13620 );
nor  g12375 ( new_n14724 , new_n13621 , new_n13640 );
nor  g12376 ( new_n14725 , new_n14723 , new_n14724 );
nor  g12377 ( new_n14726 , new_n14722 , new_n14725 );
nor  g12378 ( new_n14727 , new_n14721 , new_n14726 );
xnor g12379 ( new_n14728 , new_n14713 , new_n14714 );
nor  g12380 ( new_n14729 , new_n14727 , new_n14728 );
nor  g12381 ( new_n14730 , new_n14715 , new_n14729 );
nor  g12382 ( new_n14731 , new_n14712 , new_n14730 );
nor  g12383 ( new_n14732 , new_n14711 , new_n14731 );
nor  g12384 ( new_n14733 , new_n14708 , new_n14732 );
nor  g12385 ( new_n14734_1 , new_n14707 , new_n14733 );
xnor g12386 ( n2948 , new_n14704_1 , new_n14734_1 );
xor  g12387 ( n2961 , new_n14132 , new_n14151 );
xnor g12388 ( n2971 , new_n11239 , new_n11261_1 );
xnor g12389 ( n3010 , new_n2515_1 , new_n2534 );
xor  g12390 ( n3017 , new_n6727 , new_n6737 );
xnor g12391 ( new_n14740 , new_n8996 , new_n11592 );
xnor g12392 ( n3020 , new_n11597 , new_n14740 );
xnor g12393 ( n3067 , new_n6114 , new_n6139 );
xnor g12394 ( new_n14743 , new_n2582_1 , n23541 );
xnor g12395 ( new_n14744 , n4588 , n27134 );
xnor g12396 ( new_n14745 , new_n14743 , new_n14744 );
xnor g12397 ( n3076 , new_n9885 , new_n14745 );
nor  g12398 ( new_n14747 , n18 , n15490 );
not  g12399 ( new_n14748 , new_n14747 );
nor  g12400 ( new_n14749 , n2783 , new_n14748 );
xnor g12401 ( new_n14750 , n10611 , new_n14749 );
xnor g12402 ( new_n14751 , new_n6589 , new_n14750 );
xnor g12403 ( new_n14752 , n2783 , new_n14747 );
not  g12404 ( new_n14753 , new_n14752 );
nor  g12405 ( new_n14754 , new_n6606 , new_n14753 );
xnor g12406 ( new_n14755 , n19680 , new_n14753 );
xnor g12407 ( new_n14756 , n18 , n15490 );
and  g12408 ( new_n14757 , new_n6616 , new_n14756 );
or   g12409 ( new_n14758 , new_n6596_1 , new_n4818 );
xnor g12410 ( new_n14759 , n2809 , new_n14756 );
and  g12411 ( new_n14760 , new_n14758 , new_n14759 );
nor  g12412 ( new_n14761 , new_n14757 , new_n14760 );
and  g12413 ( new_n14762 , new_n14755 , new_n14761 );
or   g12414 ( new_n14763_1 , new_n14754 , new_n14762 );
xor  g12415 ( new_n14764 , new_n14751 , new_n14763_1 );
xnor g12416 ( new_n14765 , new_n10584 , new_n14764 );
xnor g12417 ( new_n14766 , new_n14755 , new_n14761 );
nor  g12418 ( new_n14767 , new_n10589 , new_n14766 );
xnor g12419 ( new_n14768 , new_n10588_1 , new_n14766 );
nor  g12420 ( new_n14769 , new_n5790 , new_n14759 );
xor  g12421 ( new_n14770 , new_n14758 , new_n14759 );
nor  g12422 ( new_n14771 , new_n10592 , new_n14770 );
xnor g12423 ( new_n14772_1 , n18 , n15508 );
nor  g12424 ( new_n14773 , new_n5772 , new_n14772_1 );
nor  g12425 ( new_n14774 , new_n14771 , new_n14773 );
nor  g12426 ( new_n14775 , new_n14769 , new_n14774 );
and  g12427 ( new_n14776 , new_n14768 , new_n14775 );
nor  g12428 ( new_n14777 , new_n14767 , new_n14776 );
xor  g12429 ( n3089 , new_n14765 , new_n14777 );
xnor g12430 ( n3125 , new_n5200 , new_n5201 );
xnor g12431 ( new_n14780 , new_n10958 , n21839 );
nor  g12432 ( new_n14781 , n12657 , n27089 );
or   g12433 ( new_n14782 , new_n2928 , new_n2967 );
and  g12434 ( new_n14783 , new_n2927 , new_n14782 );
nor  g12435 ( new_n14784 , new_n14781 , new_n14783 );
xnor g12436 ( new_n14785 , new_n14780 , new_n14784 );
nor  g12437 ( new_n14786 , new_n10923 , new_n14785 );
xnor g12438 ( new_n14787 , new_n10923 , new_n14785 );
nor  g12439 ( new_n14788 , new_n2969 , new_n10926 );
nor  g12440 ( new_n14789 , new_n2973 , new_n10929 );
xnor g12441 ( new_n14790_1 , new_n2974 , new_n10929 );
not  g12442 ( new_n14791 , new_n2981 );
nor  g12443 ( new_n14792 , new_n14791 , new_n10933 );
xnor g12444 ( new_n14793 , new_n14791 , new_n10932 );
nor  g12445 ( new_n14794 , new_n13097 , new_n10937 );
and  g12446 ( new_n14795 , new_n13098 , new_n13115 );
or   g12447 ( new_n14796 , new_n14794 , new_n14795 );
and  g12448 ( new_n14797 , new_n14793 , new_n14796 );
nor  g12449 ( new_n14798 , new_n14792 , new_n14797 );
and  g12450 ( new_n14799 , new_n14790_1 , new_n14798 );
or   g12451 ( new_n14800 , new_n14789 , new_n14799 );
not  g12452 ( new_n14801_1 , new_n2969 );
xnor g12453 ( new_n14802 , new_n14801_1 , new_n10926 );
and  g12454 ( new_n14803 , new_n14800 , new_n14802 );
nor  g12455 ( new_n14804 , new_n14788 , new_n14803 );
nor  g12456 ( new_n14805 , new_n14787 , new_n14804 );
nor  g12457 ( new_n14806 , new_n14786 , new_n14805 );
nor  g12458 ( new_n14807 , n19282 , n21839 );
or   g12459 ( new_n14808 , new_n14781 , new_n14783 );
and  g12460 ( new_n14809 , new_n14780 , new_n14808 );
nor  g12461 ( new_n14810 , new_n14807 , new_n14809 );
not  g12462 ( new_n14811 , new_n14810 );
and  g12463 ( new_n14812 , new_n10925 , new_n14811 );
and  g12464 ( new_n14813 , new_n14806 , new_n14812 );
or   g12465 ( new_n14814 , new_n10925 , new_n14811 );
nor  g12466 ( new_n14815 , new_n14806 , new_n14814 );
nor  g12467 ( new_n14816 , new_n14813 , new_n14815 );
xnor g12468 ( new_n14817 , new_n11794 , new_n14816 );
xnor g12469 ( new_n14818 , new_n10925 , new_n14810 );
xnor g12470 ( new_n14819_1 , new_n14806 , new_n14818 );
nor  g12471 ( new_n14820 , new_n11324 , new_n14819_1 );
xnor g12472 ( new_n14821 , new_n11324 , new_n14819_1 );
xnor g12473 ( new_n14822 , new_n14787 , new_n14804 );
nor  g12474 ( new_n14823 , new_n11339 , new_n14822 );
xnor g12475 ( new_n14824 , new_n11339 , new_n14822 );
xor  g12476 ( new_n14825 , new_n14800 , new_n14802 );
and  g12477 ( new_n14826_1 , new_n11858 , new_n14825 );
xnor g12478 ( new_n14827_1 , new_n11858 , new_n14825 );
xnor g12479 ( new_n14828 , new_n14790_1 , new_n14798 );
nor  g12480 ( new_n14829 , new_n11348_1 , new_n14828 );
xnor g12481 ( new_n14830 , new_n11348_1 , new_n14828 );
xor  g12482 ( new_n14831 , new_n14793 , new_n14796 );
nor  g12483 ( new_n14832 , new_n11352_1 , new_n14831 );
xnor g12484 ( new_n14833 , new_n11352_1 , new_n14831 );
nor  g12485 ( new_n14834 , new_n11357 , new_n13116_1 );
nor  g12486 ( new_n14835 , new_n13117 , new_n13139 );
nor  g12487 ( new_n14836 , new_n14834 , new_n14835 );
nor  g12488 ( new_n14837 , new_n14833 , new_n14836 );
nor  g12489 ( new_n14838 , new_n14832 , new_n14837 );
nor  g12490 ( new_n14839_1 , new_n14830 , new_n14838 );
nor  g12491 ( new_n14840 , new_n14829 , new_n14839_1 );
nor  g12492 ( new_n14841 , new_n14827_1 , new_n14840 );
nor  g12493 ( new_n14842 , new_n14826_1 , new_n14841 );
nor  g12494 ( new_n14843 , new_n14824 , new_n14842 );
nor  g12495 ( new_n14844 , new_n14823 , new_n14843 );
nor  g12496 ( new_n14845 , new_n14821 , new_n14844 );
nor  g12497 ( new_n14846 , new_n14820 , new_n14845 );
not  g12498 ( new_n14847 , new_n14846 );
xnor g12499 ( n3126 , new_n14817 , new_n14847 );
xnor g12500 ( n3208 , new_n11865 , new_n11898_1 );
xnor g12501 ( n3219 , new_n13971 , new_n13972 );
xnor g12502 ( n3235 , new_n14388 , new_n14395 );
xnor g12503 ( n3244 , new_n11126 , new_n11139 );
nor  g12504 ( new_n14853 , n5532 , new_n7926 );
not  g12505 ( new_n14854 , n11579 );
nor  g12506 ( new_n14855 , n3962 , new_n14854 );
nor  g12507 ( new_n14856 , new_n7931 , n23513 );
and  g12508 ( new_n14857 , new_n9875 , new_n13333_1 );
nor  g12509 ( new_n14858 , new_n7934 , n6427 );
or   g12510 ( new_n14859 , new_n14857 , new_n14858 );
and  g12511 ( new_n14860 , new_n9823 , new_n14859 );
or   g12512 ( new_n14861 , new_n14856 , new_n14860 );
and  g12513 ( new_n14862 , new_n9843 , new_n14861 );
or   g12514 ( new_n14863 , new_n14855 , new_n14862 );
and  g12515 ( new_n14864 , new_n9846 , new_n14863 );
or   g12516 ( new_n14865 , new_n14853 , new_n14864 );
xor  g12517 ( new_n14866 , new_n9849 , new_n14865 );
xnor g12518 ( new_n14867 , new_n14655 , new_n14866 );
xor  g12519 ( new_n14868 , new_n9846 , new_n14863 );
nor  g12520 ( new_n14869 , new_n14659 , new_n14868 );
xnor g12521 ( new_n14870 , new_n14659 , new_n14868 );
xor  g12522 ( new_n14871 , new_n9843 , new_n14861 );
nor  g12523 ( new_n14872 , new_n14662 , new_n14871 );
xnor g12524 ( new_n14873 , new_n14662 , new_n14871 );
xor  g12525 ( new_n14874 , new_n9823 , new_n14859 );
nor  g12526 ( new_n14875 , new_n14666 , new_n14874 );
xnor g12527 ( new_n14876 , new_n14665 , new_n14874 );
nor  g12528 ( new_n14877 , new_n13324 , new_n13335 );
nor  g12529 ( new_n14878 , new_n13336 , new_n13354 );
nor  g12530 ( new_n14879 , new_n14877 , new_n14878 );
and  g12531 ( new_n14880 , new_n14876 , new_n14879 );
nor  g12532 ( new_n14881 , new_n14875 , new_n14880 );
nor  g12533 ( new_n14882 , new_n14873 , new_n14881 );
nor  g12534 ( new_n14883 , new_n14872 , new_n14882 );
nor  g12535 ( new_n14884 , new_n14870 , new_n14883 );
nor  g12536 ( new_n14885 , new_n14869 , new_n14884 );
xnor g12537 ( new_n14886 , new_n14867 , new_n14885 );
not  g12538 ( new_n14887 , new_n14886 );
nor  g12539 ( new_n14888 , n16247 , n23541 );
not  g12540 ( new_n14889 , new_n14888 );
nor  g12541 ( new_n14890 , n8638 , new_n14889 );
not  g12542 ( new_n14891_1 , new_n14890 );
nor  g12543 ( new_n14892 , n15979 , new_n14891_1 );
not  g12544 ( new_n14893 , new_n14892 );
nor  g12545 ( new_n14894 , n26483 , new_n14893 );
not  g12546 ( new_n14895 , new_n14894 );
nor  g12547 ( new_n14896 , n24768 , new_n14895 );
not  g12548 ( new_n14897 , new_n14896 );
nor  g12549 ( new_n14898 , n8687 , new_n14897 );
xnor g12550 ( new_n14899_1 , n19270 , new_n14898 );
xnor g12551 ( new_n14900 , new_n2562 , new_n14899_1 );
xnor g12552 ( new_n14901 , n8687 , new_n14896 );
nor  g12553 ( new_n14902 , n13190 , new_n14901 );
xnor g12554 ( new_n14903 , new_n2566 , new_n14901 );
xnor g12555 ( new_n14904 , n24768 , new_n14894 );
nor  g12556 ( new_n14905 , n3460 , new_n14904 );
xnor g12557 ( new_n14906 , new_n11305 , new_n14904 );
xnor g12558 ( new_n14907 , n26483 , new_n14892 );
nor  g12559 ( new_n14908 , n5226 , new_n14907 );
xnor g12560 ( new_n14909 , new_n9502 , new_n14907 );
xnor g12561 ( new_n14910 , n15979 , new_n14890 );
nor  g12562 ( new_n14911 , n17664 , new_n14910 );
xnor g12563 ( new_n14912 , n8638 , new_n14888 );
nor  g12564 ( new_n14913 , n23369 , new_n14912 );
xnor g12565 ( new_n14914 , new_n2578_1 , new_n14912 );
xnor g12566 ( new_n14915 , n16247 , n23541 );
and  g12567 ( new_n14916 , new_n8697 , new_n14915 );
or   g12568 ( new_n14917 , new_n2582_1 , new_n2629 );
xnor g12569 ( new_n14918 , n1136 , new_n14915 );
and  g12570 ( new_n14919 , new_n14917 , new_n14918 );
or   g12571 ( new_n14920 , new_n14916 , new_n14919 );
and  g12572 ( new_n14921 , new_n14914 , new_n14920 );
or   g12573 ( new_n14922 , new_n14913 , new_n14921 );
xnor g12574 ( new_n14923 , new_n2574 , new_n14910 );
and  g12575 ( new_n14924 , new_n14922 , new_n14923 );
or   g12576 ( new_n14925 , new_n14911 , new_n14924 );
and  g12577 ( new_n14926 , new_n14909 , new_n14925 );
or   g12578 ( new_n14927 , new_n14908 , new_n14926 );
and  g12579 ( new_n14928 , new_n14906 , new_n14927 );
or   g12580 ( new_n14929 , new_n14905 , new_n14928 );
and  g12581 ( new_n14930 , new_n14903 , new_n14929 );
nor  g12582 ( new_n14931_1 , new_n14902 , new_n14930 );
xnor g12583 ( new_n14932 , new_n14900 , new_n14931_1 );
xnor g12584 ( new_n14933 , new_n14887 , new_n14932 );
nor  g12585 ( new_n14934 , new_n14905 , new_n14928 );
xnor g12586 ( new_n14935 , new_n14903 , new_n14934 );
not  g12587 ( new_n14936 , new_n14935 );
xnor g12588 ( new_n14937 , new_n14870 , new_n14883 );
nor  g12589 ( new_n14938 , new_n14936 , new_n14937 );
nor  g12590 ( new_n14939 , new_n14908 , new_n14926 );
xnor g12591 ( new_n14940 , new_n14906 , new_n14939 );
not  g12592 ( new_n14941 , new_n14940 );
xnor g12593 ( new_n14942 , new_n14873 , new_n14881 );
nor  g12594 ( new_n14943 , new_n14941 , new_n14942 );
not  g12595 ( new_n14944_1 , new_n14942 );
xnor g12596 ( new_n14945 , new_n14940 , new_n14944_1 );
nor  g12597 ( new_n14946 , new_n14911 , new_n14924 );
xnor g12598 ( new_n14947 , new_n14909 , new_n14946 );
not  g12599 ( new_n14948 , new_n14947 );
xnor g12600 ( new_n14949 , new_n14876 , new_n14879 );
nor  g12601 ( new_n14950 , new_n14948 , new_n14949 );
nor  g12602 ( new_n14951 , new_n14913 , new_n14921 );
xnor g12603 ( new_n14952 , new_n14951 , new_n14923 );
not  g12604 ( new_n14953 , new_n14952 );
nor  g12605 ( new_n14954_1 , new_n13356 , new_n14953 );
xnor g12606 ( new_n14955 , new_n13356 , new_n14952 );
xor  g12607 ( new_n14956 , new_n14914 , new_n14920 );
nor  g12608 ( new_n14957 , new_n13372 , new_n14956 );
xor  g12609 ( new_n14958 , new_n13372 , new_n14956 );
nor  g12610 ( new_n14959 , new_n2582_1 , new_n2629 );
xnor g12611 ( new_n14960 , new_n14959 , new_n14918 );
and  g12612 ( new_n14961 , new_n13385 , new_n14960 );
not  g12613 ( new_n14962 , new_n14743 );
nor  g12614 ( new_n14963 , new_n13377 , new_n14962 );
xnor g12615 ( new_n14964 , new_n13385 , new_n14960 );
nor  g12616 ( new_n14965 , new_n14963 , new_n14964 );
nor  g12617 ( new_n14966 , new_n14961 , new_n14965 );
and  g12618 ( new_n14967 , new_n14958 , new_n14966 );
nor  g12619 ( new_n14968 , new_n14957 , new_n14967 );
and  g12620 ( new_n14969 , new_n14955 , new_n14968 );
nor  g12621 ( new_n14970 , new_n14954_1 , new_n14969 );
not  g12622 ( new_n14971 , new_n14949 );
xnor g12623 ( new_n14972 , new_n14947 , new_n14971 );
nor  g12624 ( new_n14973 , new_n14970 , new_n14972 );
nor  g12625 ( new_n14974 , new_n14950 , new_n14973 );
nor  g12626 ( new_n14975 , new_n14945 , new_n14974 );
nor  g12627 ( new_n14976 , new_n14943 , new_n14975 );
xnor g12628 ( new_n14977_1 , new_n14936 , new_n14937 );
nor  g12629 ( new_n14978 , new_n14976 , new_n14977_1 );
nor  g12630 ( new_n14979 , new_n14938 , new_n14978 );
xnor g12631 ( n3263 , new_n14933 , new_n14979 );
xnor g12632 ( n3289 , new_n12078 , new_n12091 );
xnor g12633 ( new_n14982 , new_n8968 , n21832 );
nor  g12634 ( new_n14983 , new_n8971_1 , new_n2356 );
or   g12635 ( new_n14984 , n12956 , n26913 );
nor  g12636 ( new_n14985 , n16223 , n18295 );
or   g12637 ( new_n14986 , new_n5031_1 , new_n5035 );
and  g12638 ( new_n14987 , new_n5030 , new_n14986 );
nor  g12639 ( new_n14988 , new_n14985 , new_n14987 );
and  g12640 ( new_n14989_1 , new_n14984 , new_n14988 );
nor  g12641 ( new_n14990 , new_n14983 , new_n14989_1 );
xor  g12642 ( new_n14991 , new_n14982 , new_n14990 );
xnor g12643 ( new_n14992 , new_n8506 , new_n14991 );
xnor g12644 ( new_n14993 , new_n8971_1 , n26913 );
xnor g12645 ( new_n14994 , new_n14988 , new_n14993 );
nor  g12646 ( new_n14995 , n7057 , new_n14994 );
not  g12647 ( new_n14996 , new_n14994 );
xnor g12648 ( new_n14997 , n7057 , new_n14996 );
nor  g12649 ( new_n14998 , n8381 , new_n5037 );
or   g12650 ( new_n14999 , new_n5044 , new_n5049 );
and  g12651 ( new_n15000 , new_n5039 , new_n14999 );
or   g12652 ( new_n15001 , new_n14998 , new_n15000 );
and  g12653 ( new_n15002_1 , new_n14997 , new_n15001 );
nor  g12654 ( new_n15003 , new_n14995 , new_n15002_1 );
xnor g12655 ( new_n15004_1 , new_n14992 , new_n15003 );
not  g12656 ( new_n15005 , new_n15004_1 );
xnor g12657 ( new_n15006 , n21649 , new_n14048 );
nor  g12658 ( new_n15007 , n18274 , new_n9409 );
xnor g12659 ( new_n15008 , n18274 , new_n14050 );
nor  g12660 ( new_n15009 , n3828 , new_n9427 );
nor  g12661 ( new_n15010 , n23842 , new_n14057 );
not  g12662 ( new_n15011_1 , n21654 );
or   g12663 ( new_n15012 , new_n15011_1 , new_n9434 );
xnor g12664 ( new_n15013 , new_n5172 , new_n14057 );
and  g12665 ( new_n15014 , new_n15012 , new_n15013 );
or   g12666 ( new_n15015 , new_n15010 , new_n15014 );
xnor g12667 ( new_n15016 , n3828 , new_n9428 );
and  g12668 ( new_n15017 , new_n15015 , new_n15016 );
or   g12669 ( new_n15018 , new_n15009 , new_n15017 );
and  g12670 ( new_n15019_1 , new_n15008 , new_n15018 );
nor  g12671 ( new_n15020 , new_n15007 , new_n15019_1 );
xor  g12672 ( new_n15021 , new_n15006 , new_n15020 );
xnor g12673 ( new_n15022 , new_n15005 , new_n15021 );
nor  g12674 ( new_n15023 , new_n14998 , new_n15000 );
xnor g12675 ( new_n15024 , new_n14997 , new_n15023 );
xor  g12676 ( new_n15025 , new_n15008 , new_n15018 );
and  g12677 ( new_n15026 , new_n15024 , new_n15025 );
xnor g12678 ( new_n15027 , new_n15024 , new_n15025 );
xor  g12679 ( new_n15028 , new_n15015 , new_n15016 );
and  g12680 ( new_n15029 , new_n5051 , new_n15028 );
xor  g12681 ( new_n15030 , new_n15012 , new_n15013 );
and  g12682 ( new_n15031_1 , new_n5077_1 , new_n15030 );
xnor g12683 ( new_n15032 , n21654 , new_n9434 );
not  g12684 ( new_n15033_1 , new_n15032 );
nor  g12685 ( new_n15034 , new_n5081 , new_n15033_1 );
xnor g12686 ( new_n15035 , new_n5077_1 , new_n15030 );
nor  g12687 ( new_n15036 , new_n15034 , new_n15035 );
nor  g12688 ( new_n15037 , new_n15031_1 , new_n15036 );
xnor g12689 ( new_n15038 , new_n5051 , new_n15028 );
nor  g12690 ( new_n15039 , new_n15037 , new_n15038 );
nor  g12691 ( new_n15040 , new_n15029 , new_n15039 );
nor  g12692 ( new_n15041 , new_n15027 , new_n15040 );
nor  g12693 ( new_n15042 , new_n15026 , new_n15041 );
xnor g12694 ( n3301 , new_n15022 , new_n15042 );
xnor g12695 ( new_n15044 , n3030 , new_n10639 );
not  g12696 ( new_n15045 , n19515 );
nor  g12697 ( new_n15046 , new_n15045 , new_n10629 );
xnor g12698 ( new_n15047 , new_n15045 , new_n10630 );
nor  g12699 ( new_n15048 , new_n13358 , new_n10619 );
xnor g12700 ( new_n15049 , new_n13358 , new_n10620 );
nor  g12701 ( new_n15050 , n12209 , new_n10611_1 );
or   g12702 ( new_n15051 , new_n13145 , new_n10607 );
and  g12703 ( new_n15052_1 , new_n15051 , new_n13148 );
nor  g12704 ( new_n15053_1 , new_n15050 , new_n15052_1 );
and  g12705 ( new_n15054 , new_n15049 , new_n15053_1 );
or   g12706 ( new_n15055 , new_n15048 , new_n15054 );
and  g12707 ( new_n15056 , new_n15047 , new_n15055 );
nor  g12708 ( new_n15057 , new_n15046 , new_n15056 );
xnor g12709 ( new_n15058 , new_n15044 , new_n15057 );
not  g12710 ( new_n15059 , new_n15058 );
xnor g12711 ( new_n15060 , new_n9943 , new_n15059 );
nor  g12712 ( new_n15061 , new_n15048 , new_n15054 );
xnor g12713 ( new_n15062 , new_n15047 , new_n15061 );
not  g12714 ( new_n15063 , new_n15062 );
nor  g12715 ( new_n15064 , new_n9947 , new_n15063 );
xnor g12716 ( new_n15065 , new_n9948 , new_n15062 );
xnor g12717 ( new_n15066 , new_n15049 , new_n15053_1 );
nor  g12718 ( new_n15067 , new_n9952 , new_n15066 );
not  g12719 ( new_n15068 , new_n15066 );
xnor g12720 ( new_n15069 , new_n9953 , new_n15068 );
nor  g12721 ( new_n15070 , new_n9965 , new_n13149 );
and  g12722 ( new_n15071 , new_n13144_1 , new_n13151 );
nor  g12723 ( new_n15072 , new_n15070 , new_n15071 );
nor  g12724 ( new_n15073 , new_n15069 , new_n15072 );
nor  g12725 ( new_n15074 , new_n15067 , new_n15073 );
nor  g12726 ( new_n15075 , new_n15065 , new_n15074 );
nor  g12727 ( new_n15076 , new_n15064 , new_n15075 );
xor  g12728 ( n3316 , new_n15060 , new_n15076 );
xnor g12729 ( n3332 , new_n13123 , new_n13135 );
nor  g12730 ( new_n15079 , n17458 , new_n7961 );
xnor g12731 ( new_n15080 , new_n10870 , new_n7961 );
nor  g12732 ( new_n15081 , n1222 , new_n7966 );
xnor g12733 ( new_n15082_1 , new_n10873 , new_n7966 );
nor  g12734 ( new_n15083 , n25240 , new_n7971 );
nor  g12735 ( new_n15084 , new_n10412 , new_n10429 );
or   g12736 ( new_n15085 , new_n15083 , new_n15084 );
and  g12737 ( new_n15086 , new_n15082_1 , new_n15085 );
or   g12738 ( new_n15087 , new_n15081 , new_n15086 );
and  g12739 ( new_n15088 , new_n15080 , new_n15087 );
nor  g12740 ( new_n15089 , new_n15079 , new_n15088 );
and  g12741 ( new_n15090 , new_n8026 , new_n15089 );
nor  g12742 ( new_n15091 , new_n14547_1 , new_n12681 );
and  g12743 ( new_n15092 , new_n12682 , new_n12693 );
nor  g12744 ( new_n15093 , new_n15091 , new_n15092 );
nor  g12745 ( new_n15094_1 , n11898 , n23166 );
and  g12746 ( new_n15095 , new_n12672 , new_n12680 );
or   g12747 ( new_n15096 , new_n15094_1 , new_n15095 );
nor  g12748 ( new_n15097 , new_n15093 , new_n15096 );
not  g12749 ( new_n15098 , new_n15097 );
xnor g12750 ( new_n15099 , new_n15090 , new_n15098 );
xnor g12751 ( new_n15100 , new_n8027_1 , new_n15089 );
xnor g12752 ( new_n15101 , new_n15093 , new_n15096 );
nor  g12753 ( new_n15102 , new_n15100 , new_n15101 );
xnor g12754 ( new_n15103 , new_n15100 , new_n15101 );
not  g12755 ( new_n15104 , new_n15103 );
xor  g12756 ( new_n15105 , new_n15080 , new_n15087 );
nor  g12757 ( new_n15106 , new_n12694 , new_n15105 );
xor  g12758 ( new_n15107 , new_n12694 , new_n15105 );
xor  g12759 ( new_n15108 , new_n15082_1 , new_n15085 );
and  g12760 ( new_n15109 , new_n12699 , new_n15108 );
nor  g12761 ( new_n15110 , new_n10430 , new_n10477 );
nor  g12762 ( new_n15111 , new_n10478 , new_n10503 );
nor  g12763 ( new_n15112 , new_n15110 , new_n15111 );
xnor g12764 ( new_n15113 , new_n12699 , new_n15108 );
nor  g12765 ( new_n15114 , new_n15112 , new_n15113 );
nor  g12766 ( new_n15115 , new_n15109 , new_n15114 );
and  g12767 ( new_n15116 , new_n15107 , new_n15115 );
nor  g12768 ( new_n15117 , new_n15106 , new_n15116 );
and  g12769 ( new_n15118_1 , new_n15104 , new_n15117 );
nor  g12770 ( new_n15119 , new_n15102 , new_n15118_1 );
xnor g12771 ( n3340 , new_n15099 , new_n15119 );
xnor g12772 ( new_n15121 , n5077 , n13851 );
nor  g12773 ( new_n15122 , new_n10452 , n24937 );
xnor g12774 ( new_n15123 , n15546 , n24937 );
not  g12775 ( new_n15124 , n5098 );
and  g12776 ( new_n15125 , new_n15124 , n26452 );
xnor g12777 ( new_n15126 , n5098 , n26452 );
nor  g12778 ( new_n15127 , n3030 , new_n10460 );
xnor g12779 ( new_n15128_1 , n3030 , n19905 );
nor  g12780 ( new_n15129 , n17035 , new_n15045 );
or   g12781 ( new_n15130 , new_n13359 , new_n13367_1 );
and  g12782 ( new_n15131 , new_n13357 , new_n15130 );
nor  g12783 ( new_n15132 , new_n15129 , new_n15131 );
and  g12784 ( new_n15133 , new_n15128_1 , new_n15132 );
or   g12785 ( new_n15134 , new_n15127 , new_n15133 );
and  g12786 ( new_n15135 , new_n15126 , new_n15134 );
or   g12787 ( new_n15136 , new_n15125 , new_n15135 );
and  g12788 ( new_n15137 , new_n15123 , new_n15136 );
or   g12789 ( new_n15138 , new_n15122 , new_n15137 );
xor  g12790 ( new_n15139_1 , new_n15121 , new_n15138 );
xnor g12791 ( new_n15140 , new_n14887 , new_n15139_1 );
xor  g12792 ( new_n15141 , new_n15123 , new_n15136 );
nor  g12793 ( new_n15142 , new_n14937 , new_n15141 );
xnor g12794 ( new_n15143 , new_n14937 , new_n15141 );
xor  g12795 ( new_n15144 , new_n15126 , new_n15134 );
nor  g12796 ( new_n15145_1 , new_n14942 , new_n15144 );
xnor g12797 ( new_n15146_1 , new_n14944_1 , new_n15144 );
xnor g12798 ( new_n15147 , new_n15128_1 , new_n15132 );
nor  g12799 ( new_n15148 , new_n14971 , new_n15147 );
not  g12800 ( new_n15149 , new_n15147 );
xnor g12801 ( new_n15150 , new_n14971 , new_n15149 );
nor  g12802 ( new_n15151 , new_n13356 , new_n13370 );
nor  g12803 ( new_n15152 , new_n13371 , new_n13390 );
nor  g12804 ( new_n15153 , new_n15151 , new_n15152 );
and  g12805 ( new_n15154 , new_n15150 , new_n15153 );
nor  g12806 ( new_n15155 , new_n15148 , new_n15154 );
and  g12807 ( new_n15156 , new_n15146_1 , new_n15155 );
nor  g12808 ( new_n15157 , new_n15145_1 , new_n15156 );
nor  g12809 ( new_n15158 , new_n15143 , new_n15157 );
nor  g12810 ( new_n15159 , new_n15142 , new_n15158 );
xor  g12811 ( n3343 , new_n15140 , new_n15159 );
not  g12812 ( new_n15161 , new_n14898 );
nor  g12813 ( new_n15162 , n19270 , new_n15161 );
not  g12814 ( new_n15163 , new_n15162 );
nor  g12815 ( new_n15164 , n14704 , new_n15163 );
and  g12816 ( new_n15165_1 , new_n14347 , new_n15164 );
xnor g12817 ( new_n15166 , n25365 , new_n15164 );
nor  g12818 ( new_n15167_1 , n20040 , new_n15166 );
xnor g12819 ( new_n15168 , n14704 , new_n15162 );
nor  g12820 ( new_n15169 , n19531 , new_n15168 );
xnor g12821 ( new_n15170 , new_n2558 , new_n15168 );
nor  g12822 ( new_n15171 , n18345 , new_n14899_1 );
or   g12823 ( new_n15172 , new_n14902 , new_n14930 );
and  g12824 ( new_n15173 , new_n14900 , new_n15172 );
or   g12825 ( new_n15174 , new_n15171 , new_n15173 );
and  g12826 ( new_n15175 , new_n15170 , new_n15174 );
nor  g12827 ( new_n15176_1 , new_n15169 , new_n15175 );
and  g12828 ( new_n15177 , n20040 , new_n15166 );
nor  g12829 ( new_n15178 , new_n15176_1 , new_n15177 );
nor  g12830 ( new_n15179 , new_n15167_1 , new_n15178 );
nor  g12831 ( new_n15180_1 , new_n15165_1 , new_n15179 );
xnor g12832 ( new_n15181 , new_n11289 , new_n15166 );
xnor g12833 ( new_n15182_1 , new_n15176_1 , new_n15181 );
nor  g12834 ( new_n15183 , new_n13702 , new_n15182_1 );
not  g12835 ( new_n15184 , new_n15182_1 );
nor  g12836 ( new_n15185 , new_n13701 , new_n15184 );
nor  g12837 ( new_n15186 , new_n15171 , new_n15173 );
xnor g12838 ( new_n15187 , new_n15170 , new_n15186 );
nor  g12839 ( new_n15188 , new_n13685 , new_n15187 );
not  g12840 ( new_n15189 , new_n15187 );
xnor g12841 ( new_n15190 , new_n13685 , new_n15189 );
nor  g12842 ( new_n15191 , new_n13688 , new_n14932 );
not  g12843 ( new_n15192 , new_n14932 );
xnor g12844 ( new_n15193 , new_n13688 , new_n15192 );
nor  g12845 ( new_n15194 , new_n6472 , new_n14935 );
xnor g12846 ( new_n15195 , new_n6472 , new_n14936 );
nor  g12847 ( new_n15196 , new_n6476_1 , new_n14940 );
nor  g12848 ( new_n15197 , new_n6480 , new_n14947 );
xnor g12849 ( new_n15198 , new_n6480 , new_n14948 );
nor  g12850 ( new_n15199 , new_n6482 , new_n14953 );
xnor g12851 ( new_n15200 , new_n6499 , new_n14953 );
nor  g12852 ( new_n15201 , new_n6486 , new_n14956 );
xnor g12853 ( new_n15202 , new_n6484 , new_n14956 );
not  g12854 ( new_n15203 , new_n14960 );
nor  g12855 ( new_n15204 , new_n6489 , new_n15203 );
or   g12856 ( new_n15205_1 , new_n6491 , new_n14962 );
xnor g12857 ( new_n15206 , new_n6488 , new_n15203 );
and  g12858 ( new_n15207 , new_n15205_1 , new_n15206 );
nor  g12859 ( new_n15208 , new_n15204 , new_n15207 );
and  g12860 ( new_n15209 , new_n15202 , new_n15208 );
nor  g12861 ( new_n15210 , new_n15201 , new_n15209 );
and  g12862 ( new_n15211 , new_n15200 , new_n15210 );
nor  g12863 ( new_n15212 , new_n15199 , new_n15211 );
and  g12864 ( new_n15213 , new_n15198 , new_n15212 );
or   g12865 ( new_n15214 , new_n15197 , new_n15213 );
xnor g12866 ( new_n15215 , new_n6476_1 , new_n14941 );
and  g12867 ( new_n15216 , new_n15214 , new_n15215 );
or   g12868 ( new_n15217 , new_n15196 , new_n15216 );
and  g12869 ( new_n15218 , new_n15195 , new_n15217 );
or   g12870 ( new_n15219 , new_n15194 , new_n15218 );
and  g12871 ( new_n15220 , new_n15193 , new_n15219 );
or   g12872 ( new_n15221 , new_n15191 , new_n15220 );
and  g12873 ( new_n15222 , new_n15190 , new_n15221 );
nor  g12874 ( new_n15223 , new_n15188 , new_n15222 );
nor  g12875 ( new_n15224 , new_n15185 , new_n15223 );
or   g12876 ( new_n15225 , new_n13724 , new_n15224 );
or   g12877 ( new_n15226 , new_n15183 , new_n15225 );
xnor g12878 ( new_n15227 , new_n15180_1 , new_n15226 );
and  g12879 ( new_n15228 , new_n11795 , new_n12251 );
xnor g12880 ( new_n15229 , new_n11795 , new_n12251 );
and  g12881 ( new_n15230_1 , new_n6155 , new_n12255 );
xnor g12882 ( new_n15231 , new_n6155 , new_n12255 );
and  g12883 ( new_n15232 , new_n6158 , new_n12259 );
xnor g12884 ( new_n15233 , new_n6158 , new_n12259 );
and  g12885 ( new_n15234 , new_n6161 , new_n12263 );
xnor g12886 ( new_n15235 , new_n6161 , new_n12263 );
and  g12887 ( new_n15236 , new_n11812 , new_n12267 );
xnor g12888 ( new_n15237 , new_n11812 , new_n12267 );
not  g12889 ( new_n15238 , n21226 );
and  g12890 ( new_n15239 , new_n15238 , new_n12271 );
xnor g12891 ( new_n15240 , new_n15238 , new_n12271 );
nor  g12892 ( new_n15241_1 , n4426 , new_n12275 );
xnor g12893 ( new_n15242 , new_n6170 , new_n12275 );
nor  g12894 ( new_n15243 , n20036 , new_n12282 );
xnor g12895 ( new_n15244 , new_n8659 , new_n12282 );
nor  g12896 ( new_n15245 , new_n4120 , new_n12291 );
or   g12897 ( new_n15246 , n9380 , new_n12287 );
xnor g12898 ( new_n15247 , new_n4120 , new_n12290 );
and  g12899 ( new_n15248 , new_n15246 , new_n15247 );
nor  g12900 ( new_n15249 , new_n15245 , new_n15248 );
and  g12901 ( new_n15250 , new_n15244 , new_n15249 );
or   g12902 ( new_n15251 , new_n15243 , new_n15250 );
and  g12903 ( new_n15252 , new_n15242 , new_n15251 );
nor  g12904 ( new_n15253 , new_n15241_1 , new_n15252 );
nor  g12905 ( new_n15254 , new_n15240 , new_n15253 );
nor  g12906 ( new_n15255_1 , new_n15239 , new_n15254 );
nor  g12907 ( new_n15256 , new_n15237 , new_n15255_1 );
nor  g12908 ( new_n15257 , new_n15236 , new_n15256 );
nor  g12909 ( new_n15258_1 , new_n15235 , new_n15257 );
nor  g12910 ( new_n15259 , new_n15234 , new_n15258_1 );
nor  g12911 ( new_n15260 , new_n15233 , new_n15259 );
nor  g12912 ( new_n15261 , new_n15232 , new_n15260 );
nor  g12913 ( new_n15262 , new_n15231 , new_n15261 );
nor  g12914 ( new_n15263 , new_n15230_1 , new_n15262 );
nor  g12915 ( new_n15264 , new_n15229 , new_n15263 );
nor  g12916 ( new_n15265 , new_n15228 , new_n15264 );
xnor g12917 ( new_n15266 , new_n12156 , new_n15265 );
nor  g12918 ( new_n15267 , new_n15227 , new_n15266 );
xnor g12919 ( new_n15268 , new_n15229 , new_n15263 );
xnor g12920 ( new_n15269 , new_n13702 , new_n15184 );
xnor g12921 ( new_n15270 , new_n15223 , new_n15269 );
nor  g12922 ( new_n15271_1 , new_n15268 , new_n15270 );
xnor g12923 ( new_n15272 , new_n15268 , new_n15270 );
xnor g12924 ( new_n15273 , new_n15231 , new_n15261 );
xor  g12925 ( new_n15274 , new_n15190 , new_n15221 );
nor  g12926 ( new_n15275_1 , new_n15273 , new_n15274 );
xnor g12927 ( new_n15276 , new_n15273 , new_n15274 );
xnor g12928 ( new_n15277 , new_n15233 , new_n15259 );
xor  g12929 ( new_n15278 , new_n15193 , new_n15219 );
nor  g12930 ( new_n15279 , new_n15277 , new_n15278 );
xnor g12931 ( new_n15280 , new_n15277 , new_n15278 );
xnor g12932 ( new_n15281 , new_n15235 , new_n15257 );
xor  g12933 ( new_n15282 , new_n15195 , new_n15217 );
nor  g12934 ( new_n15283 , new_n15281 , new_n15282 );
xnor g12935 ( new_n15284 , new_n15281 , new_n15282 );
xnor g12936 ( new_n15285 , new_n15237 , new_n15255_1 );
xor  g12937 ( new_n15286 , new_n15214 , new_n15215 );
nor  g12938 ( new_n15287 , new_n15285 , new_n15286 );
xnor g12939 ( new_n15288 , new_n15285 , new_n15286 );
xnor g12940 ( new_n15289_1 , new_n15240 , new_n15253 );
xnor g12941 ( new_n15290 , new_n15198 , new_n15212 );
not  g12942 ( new_n15291 , new_n15290 );
nor  g12943 ( new_n15292 , new_n15289_1 , new_n15291 );
xnor g12944 ( new_n15293 , new_n15289_1 , new_n15291 );
xor  g12945 ( new_n15294 , new_n15242 , new_n15251 );
xnor g12946 ( new_n15295 , new_n15200 , new_n15210 );
not  g12947 ( new_n15296 , new_n15295 );
and  g12948 ( new_n15297 , new_n15294 , new_n15296 );
xnor g12949 ( new_n15298 , new_n15294 , new_n15296 );
xnor g12950 ( new_n15299 , new_n15244 , new_n15249 );
xnor g12951 ( new_n15300_1 , new_n15202 , new_n15208 );
not  g12952 ( new_n15301 , new_n15300_1 );
nor  g12953 ( new_n15302 , new_n15299 , new_n15301 );
nor  g12954 ( new_n15303 , new_n6491 , new_n14962 );
xnor g12955 ( new_n15304 , new_n15303 , new_n15206 );
not  g12956 ( new_n15305 , new_n15304 );
xor  g12957 ( new_n15306 , new_n15246 , new_n15247 );
and  g12958 ( new_n15307_1 , new_n15305 , new_n15306 );
xnor g12959 ( new_n15308 , n4939 , new_n14962 );
not  g12960 ( new_n15309 , new_n15308 );
xnor g12961 ( new_n15310 , new_n6176 , new_n12287 );
nor  g12962 ( new_n15311 , new_n15309 , new_n15310 );
xnor g12963 ( new_n15312 , new_n15304 , new_n15306 );
and  g12964 ( new_n15313 , new_n15311 , new_n15312 );
nor  g12965 ( new_n15314 , new_n15307_1 , new_n15313 );
xnor g12966 ( new_n15315 , new_n15299 , new_n15300_1 );
and  g12967 ( new_n15316 , new_n15314 , new_n15315 );
nor  g12968 ( new_n15317 , new_n15302 , new_n15316 );
nor  g12969 ( new_n15318 , new_n15298 , new_n15317 );
nor  g12970 ( new_n15319 , new_n15297 , new_n15318 );
nor  g12971 ( new_n15320 , new_n15293 , new_n15319 );
nor  g12972 ( new_n15321 , new_n15292 , new_n15320 );
nor  g12973 ( new_n15322 , new_n15288 , new_n15321 );
nor  g12974 ( new_n15323 , new_n15287 , new_n15322 );
nor  g12975 ( new_n15324 , new_n15284 , new_n15323 );
nor  g12976 ( new_n15325 , new_n15283 , new_n15324 );
nor  g12977 ( new_n15326 , new_n15280 , new_n15325 );
nor  g12978 ( new_n15327_1 , new_n15279 , new_n15326 );
nor  g12979 ( new_n15328 , new_n15276 , new_n15327_1 );
nor  g12980 ( new_n15329 , new_n15275_1 , new_n15328 );
nor  g12981 ( new_n15330 , new_n15272 , new_n15329 );
nor  g12982 ( new_n15331 , new_n15271_1 , new_n15330 );
xnor g12983 ( new_n15332_1 , new_n15227 , new_n15266 );
nor  g12984 ( new_n15333 , new_n15331 , new_n15332_1 );
nor  g12985 ( new_n15334 , new_n15267 , new_n15333 );
nor  g12986 ( new_n15335 , new_n15180_1 , new_n15226 );
or   g12987 ( new_n15336 , new_n12111 , new_n12155 );
and  g12988 ( new_n15337 , new_n15336 , new_n15265 );
xor  g12989 ( new_n15338 , new_n15335 , new_n15337 );
xnor g12990 ( n3390 , new_n15334 , new_n15338 );
xnor g12991 ( n3426 , new_n6572 , new_n6573 );
not  g12992 ( new_n15341 , new_n4740 );
xnor g12993 ( n3451 , new_n4739 , new_n15341 );
xnor g12994 ( n3459 , new_n11991 , new_n12008 );
xnor g12995 ( new_n15344 , new_n5587 , n6773 );
xnor g12996 ( new_n15345_1 , n21687 , new_n15344 );
nor  g12997 ( new_n15346 , new_n13471 , new_n15345_1 );
nor  g12998 ( new_n15347 , new_n2548 , new_n15344 );
nor  g12999 ( new_n15348 , n6729 , new_n15347 );
or   g13000 ( new_n15349 , new_n6178 , new_n2548 );
nor  g13001 ( new_n15350 , new_n15349 , new_n15344 );
nor  g13002 ( new_n15351 , new_n15348 , new_n15350 );
nor  g13003 ( new_n15352 , new_n5587 , new_n4030 );
xnor g13004 ( new_n15353_1 , n17090 , n22173 );
xor  g13005 ( new_n15354 , new_n15352 , new_n15353_1 );
xnor g13006 ( new_n15355 , new_n15351 , new_n15354 );
not  g13007 ( new_n15356 , new_n15355 );
xnor g13008 ( new_n15357 , new_n13466 , new_n15356 );
xnor g13009 ( n3502 , new_n15346 , new_n15357 );
xnor g13010 ( n3516 , new_n10738 , new_n10771 );
nor  g13011 ( new_n15360 , n22274 , n24129 );
not  g13012 ( new_n15361 , new_n15360 );
nor  g13013 ( new_n15362 , n1689 , new_n15361 );
not  g13014 ( new_n15363 , new_n15362 );
nor  g13015 ( new_n15364 , n19608 , new_n15363 );
not  g13016 ( new_n15365 , new_n15364 );
nor  g13017 ( new_n15366_1 , n25126 , new_n15365 );
not  g13018 ( new_n15367 , new_n15366_1 );
nor  g13019 ( new_n15368 , n10712 , new_n15367 );
xnor g13020 ( new_n15369 , n18145 , new_n15368 );
xnor g13021 ( new_n15370 , n15761 , new_n15369 );
xnor g13022 ( new_n15371 , n10712 , new_n15366_1 );
nor  g13023 ( new_n15372 , new_n10179 , new_n15371 );
xnor g13024 ( new_n15373 , n11201 , new_n15371 );
xnor g13025 ( new_n15374 , n25126 , new_n15364 );
nor  g13026 ( new_n15375 , new_n10182 , new_n15374 );
xnor g13027 ( new_n15376 , n18690 , new_n15374 );
xnor g13028 ( new_n15377 , n19608 , new_n15363 );
and  g13029 ( new_n15378_1 , n12153 , new_n15377 );
xnor g13030 ( new_n15379 , n19608 , new_n15362 );
xnor g13031 ( new_n15380 , n12153 , new_n15379 );
xnor g13032 ( new_n15381 , n1689 , new_n15360 );
nor  g13033 ( new_n15382_1 , new_n10186 , new_n15381 );
xnor g13034 ( new_n15383 , n13044 , new_n15381 );
xnor g13035 ( new_n15384 , new_n4118 , n24129 );
nor  g13036 ( new_n15385 , new_n5807 , new_n15384 );
nor  g13037 ( new_n15386 , new_n5805 , n24129 );
xnor g13038 ( new_n15387 , n18745 , new_n15384 );
and  g13039 ( new_n15388 , new_n15386 , new_n15387 );
or   g13040 ( new_n15389 , new_n15385 , new_n15388 );
and  g13041 ( new_n15390 , new_n15383 , new_n15389 );
or   g13042 ( new_n15391 , new_n15382_1 , new_n15390 );
and  g13043 ( new_n15392 , new_n15380 , new_n15391 );
or   g13044 ( new_n15393 , new_n15378_1 , new_n15392 );
and  g13045 ( new_n15394 , new_n15376 , new_n15393 );
or   g13046 ( new_n15395 , new_n15375 , new_n15394 );
and  g13047 ( new_n15396 , new_n15373 , new_n15395 );
or   g13048 ( new_n15397 , new_n15372 , new_n15396 );
xor  g13049 ( new_n15398 , new_n15370 , new_n15397 );
xnor g13050 ( new_n15399 , new_n6874 , new_n15398 );
xor  g13051 ( new_n15400 , new_n15373 , new_n15395 );
and  g13052 ( new_n15401 , new_n6877 , new_n15400 );
xnor g13053 ( new_n15402 , new_n6877 , new_n15400 );
xor  g13054 ( new_n15403 , new_n15376 , new_n15393 );
and  g13055 ( new_n15404 , new_n6882 , new_n15403 );
xnor g13056 ( new_n15405 , new_n6882 , new_n15403 );
xor  g13057 ( new_n15406 , new_n15380 , new_n15391 );
and  g13058 ( new_n15407_1 , new_n6886 , new_n15406 );
xnor g13059 ( new_n15408 , new_n6888 , new_n15406 );
xor  g13060 ( new_n15409 , new_n15383 , new_n15389 );
nor  g13061 ( new_n15410 , new_n4115 , new_n15409 );
xnor g13062 ( new_n15411 , new_n4116 , new_n15409 );
xor  g13063 ( new_n15412 , new_n15386 , new_n15387 );
nor  g13064 ( new_n15413 , new_n4130 , new_n15412 );
xnor g13065 ( new_n15414 , n16167 , n24129 );
nor  g13066 ( new_n15415 , new_n4135 , new_n15414 );
xnor g13067 ( new_n15416 , new_n4138 , new_n15412 );
and  g13068 ( new_n15417 , new_n15415 , new_n15416 );
or   g13069 ( new_n15418 , new_n15413 , new_n15417 );
and  g13070 ( new_n15419 , new_n15411 , new_n15418 );
nor  g13071 ( new_n15420 , new_n15410 , new_n15419 );
and  g13072 ( new_n15421 , new_n15408 , new_n15420 );
nor  g13073 ( new_n15422 , new_n15407_1 , new_n15421 );
nor  g13074 ( new_n15423 , new_n15405 , new_n15422 );
nor  g13075 ( new_n15424_1 , new_n15404 , new_n15423 );
nor  g13076 ( new_n15425 , new_n15402 , new_n15424_1 );
or   g13077 ( new_n15426 , new_n15401 , new_n15425 );
xor  g13078 ( new_n15427 , new_n15399 , new_n15426 );
xnor g13079 ( new_n15428_1 , new_n10305 , new_n15427 );
xnor g13080 ( new_n15429 , new_n15402 , new_n15424_1 );
nor  g13081 ( new_n15430 , new_n10310 , new_n15429 );
xnor g13082 ( new_n15431 , new_n10310 , new_n15429 );
xnor g13083 ( new_n15432 , new_n15405 , new_n15422 );
nor  g13084 ( new_n15433 , new_n10314 , new_n15432 );
xnor g13085 ( new_n15434 , new_n10314 , new_n15432 );
xnor g13086 ( new_n15435_1 , new_n15408 , new_n15420 );
nor  g13087 ( new_n15436 , new_n10319 , new_n15435_1 );
xor  g13088 ( new_n15437 , new_n15411 , new_n15418 );
nor  g13089 ( new_n15438_1 , new_n10322 , new_n15437 );
xnor g13090 ( new_n15439 , new_n10322 , new_n15437 );
xor  g13091 ( new_n15440 , new_n15415 , new_n15416 );
nor  g13092 ( new_n15441 , new_n5814 , new_n15440 );
xnor g13093 ( new_n15442 , new_n4134_1 , new_n15414 );
and  g13094 ( new_n15443 , new_n5799 , new_n15442 );
xnor g13095 ( new_n15444 , new_n5814 , new_n15440 );
nor  g13096 ( new_n15445 , new_n15443 , new_n15444 );
nor  g13097 ( new_n15446 , new_n15441 , new_n15445 );
nor  g13098 ( new_n15447 , new_n15439 , new_n15446 );
nor  g13099 ( new_n15448 , new_n15438_1 , new_n15447 );
xnor g13100 ( new_n15449 , new_n10319 , new_n15435_1 );
nor  g13101 ( new_n15450 , new_n15448 , new_n15449 );
nor  g13102 ( new_n15451 , new_n15436 , new_n15450 );
nor  g13103 ( new_n15452 , new_n15434 , new_n15451 );
nor  g13104 ( new_n15453 , new_n15433 , new_n15452 );
nor  g13105 ( new_n15454 , new_n15431 , new_n15453 );
nor  g13106 ( new_n15455 , new_n15430 , new_n15454 );
xor  g13107 ( n3528 , new_n15428_1 , new_n15455 );
xnor g13108 ( n3555 , new_n9001 , new_n9057 );
nor  g13109 ( new_n15458 , new_n2673 , new_n10052 );
and  g13110 ( new_n15459 , new_n2720 , new_n2782 );
nor  g13111 ( new_n15460 , new_n15458 , new_n15459 );
not  g13112 ( new_n15461 , new_n15460 );
nor  g13113 ( new_n15462 , n13951 , new_n2672 );
and  g13114 ( new_n15463 , new_n15462 , new_n10050 );
and  g13115 ( new_n15464 , new_n15461 , new_n15463 );
or   g13116 ( new_n15465_1 , new_n15462 , new_n10050 );
nor  g13117 ( new_n15466 , new_n15461 , new_n15465_1 );
nor  g13118 ( new_n15467_1 , new_n15464 , new_n15466 );
nor  g13119 ( new_n15468 , new_n14356 , new_n15467_1 );
xnor g13120 ( new_n15469 , new_n14356 , new_n15467_1 );
xnor g13121 ( new_n15470_1 , new_n15462 , new_n10049 );
xnor g13122 ( new_n15471 , new_n15461 , new_n15470_1 );
nor  g13123 ( new_n15472 , new_n14361 , new_n15471 );
xnor g13124 ( new_n15473 , new_n14361 , new_n15471 );
nor  g13125 ( new_n15474 , new_n2655 , new_n2783_1 );
and  g13126 ( new_n15475 , new_n2784 , new_n2847 );
nor  g13127 ( new_n15476 , new_n15474 , new_n15475 );
nor  g13128 ( new_n15477_1 , new_n15473 , new_n15476 );
nor  g13129 ( new_n15478 , new_n15472 , new_n15477_1 );
nor  g13130 ( new_n15479 , new_n15469 , new_n15478 );
nor  g13131 ( new_n15480 , new_n15468 , new_n15479 );
nor  g13132 ( n3561 , new_n15464 , new_n15480 );
xnor g13133 ( new_n15482 , n14680 , n16439 );
and  g13134 ( new_n15483 , new_n4369 , n17250 );
and  g13135 ( new_n15484 , new_n10505 , new_n10525_1 );
or   g13136 ( new_n15485 , new_n15483 , new_n15484 );
xor  g13137 ( new_n15486 , new_n15482 , new_n15485 );
xnor g13138 ( new_n15487 , new_n7613 , new_n9613 );
not  g13139 ( new_n15488 , new_n15487 );
nor  g13140 ( new_n15489 , n13783 , new_n9617 );
nor  g13141 ( new_n15490_1 , new_n10528 , new_n10540_1 );
nor  g13142 ( new_n15491 , new_n15489 , new_n15490_1 );
xnor g13143 ( new_n15492 , new_n15488 , new_n15491 );
xnor g13144 ( new_n15493 , new_n15486 , new_n15492 );
and  g13145 ( new_n15494 , new_n10526 , new_n10541 );
nor  g13146 ( new_n15495 , new_n10542 , new_n10574 );
nor  g13147 ( new_n15496_1 , new_n15494 , new_n15495 );
xnor g13148 ( new_n15497 , new_n15493 , new_n15496_1 );
not  g13149 ( new_n15498 , new_n15497 );
xnor g13150 ( new_n15499 , new_n5625 , new_n15498 );
nor  g13151 ( new_n15500 , new_n5632 , new_n10575 );
and  g13152 ( new_n15501_1 , new_n10577_1 , new_n10605 );
nor  g13153 ( new_n15502 , new_n15500 , new_n15501_1 );
xor  g13154 ( n3563 , new_n15499 , new_n15502 );
xor  g13155 ( n3617 , new_n6131 , new_n6133 );
xnor g13156 ( new_n15505 , n8305 , n22253 );
and  g13157 ( new_n15506_1 , n1255 , new_n7043 );
xnor g13158 ( new_n15507 , n1255 , n12861 );
and  g13159 ( new_n15508_1 , n9512 , new_n7046 );
xnor g13160 ( new_n15509 , n9512 , n13333 );
and  g13161 ( new_n15510 , new_n7049 , n16608 );
and  g13162 ( new_n15511 , new_n5125 , n21735 );
and  g13163 ( new_n15512 , new_n4613 , new_n4635 );
or   g13164 ( new_n15513 , new_n15511 , new_n15512 );
xnor g13165 ( new_n15514 , n2210 , n16608 );
and  g13166 ( new_n15515 , new_n15513 , new_n15514 );
or   g13167 ( new_n15516 , new_n15510 , new_n15515 );
and  g13168 ( new_n15517 , new_n15509 , new_n15516 );
or   g13169 ( new_n15518 , new_n15508_1 , new_n15517 );
and  g13170 ( new_n15519 , new_n15507 , new_n15518 );
or   g13171 ( new_n15520 , new_n15506_1 , new_n15519 );
xor  g13172 ( new_n15521 , new_n15505 , new_n15520 );
xnor g13173 ( new_n15522 , new_n11226 , new_n15521 );
xor  g13174 ( new_n15523 , new_n15507 , new_n15518 );
nor  g13175 ( new_n15524 , new_n11229 , new_n15523 );
xnor g13176 ( new_n15525 , new_n11229 , new_n15523 );
xor  g13177 ( new_n15526 , new_n15509 , new_n15516 );
nor  g13178 ( new_n15527 , new_n11233 , new_n15526 );
xor  g13179 ( new_n15528 , new_n15513 , new_n15514 );
and  g13180 ( new_n15529 , new_n11237 , new_n15528 );
xnor g13181 ( new_n15530 , new_n11236 , new_n15528 );
and  g13182 ( new_n15531 , new_n4636 , new_n11240 );
and  g13183 ( new_n15532 , new_n4724 , new_n4756 );
or   g13184 ( new_n15533 , new_n15531 , new_n15532 );
and  g13185 ( new_n15534 , new_n15530 , new_n15533 );
nor  g13186 ( new_n15535 , new_n15529 , new_n15534 );
xnor g13187 ( new_n15536 , new_n11233 , new_n15526 );
not  g13188 ( new_n15537 , new_n15536 );
and  g13189 ( new_n15538 , new_n15535 , new_n15537 );
nor  g13190 ( new_n15539_1 , new_n15527 , new_n15538 );
nor  g13191 ( new_n15540 , new_n15525 , new_n15539_1 );
nor  g13192 ( new_n15541 , new_n15524 , new_n15540 );
xor  g13193 ( n3642 , new_n15522 , new_n15541 );
xnor g13194 ( new_n15543 , new_n3087 , n16544 );
nor  g13195 ( new_n15544 , n6814 , n23463 );
xnor g13196 ( new_n15545 , new_n2887_1 , n23463 );
nor  g13197 ( new_n15546_1 , n13074 , n19701 );
xnor g13198 ( new_n15547 , new_n3095 , n19701 );
nor  g13199 ( new_n15548 , n10739 , n23529 );
xnor g13200 ( new_n15549 , new_n3099 , n23529 );
nor  g13201 ( new_n15550 , n21753 , n24620 );
xnor g13202 ( new_n15551 , new_n2350 , n24620 );
nor  g13203 ( new_n15552 , n5211 , n21832 );
and  g13204 ( new_n15553 , new_n14982 , new_n14990 );
or   g13205 ( new_n15554 , new_n15552 , new_n15553 );
and  g13206 ( new_n15555_1 , new_n15551 , new_n15554 );
or   g13207 ( new_n15556 , new_n15550 , new_n15555_1 );
and  g13208 ( new_n15557 , new_n15549 , new_n15556 );
or   g13209 ( new_n15558_1 , new_n15548 , new_n15557 );
and  g13210 ( new_n15559_1 , new_n15547 , new_n15558_1 );
or   g13211 ( new_n15560 , new_n15546_1 , new_n15559_1 );
and  g13212 ( new_n15561 , new_n15545 , new_n15560 );
nor  g13213 ( new_n15562 , new_n15544 , new_n15561 );
xnor g13214 ( new_n15563 , new_n15543 , new_n15562 );
not  g13215 ( new_n15564 , new_n15563 );
xnor g13216 ( new_n15565 , n3324 , new_n15564 );
nor  g13217 ( new_n15566 , new_n15546_1 , new_n15559_1 );
xnor g13218 ( new_n15567 , new_n15545 , new_n15566 );
nor  g13219 ( new_n15568 , n17911 , new_n15567 );
not  g13220 ( new_n15569 , new_n15567 );
xnor g13221 ( new_n15570_1 , n17911 , new_n15569 );
nor  g13222 ( new_n15571 , new_n15548 , new_n15557 );
xnor g13223 ( new_n15572 , new_n15547 , new_n15571 );
nor  g13224 ( new_n15573_1 , n21997 , new_n15572 );
not  g13225 ( new_n15574 , new_n15572 );
xnor g13226 ( new_n15575 , n21997 , new_n15574 );
nor  g13227 ( new_n15576 , new_n15550 , new_n15555_1 );
xnor g13228 ( new_n15577 , new_n15549 , new_n15576 );
nor  g13229 ( new_n15578 , n25119 , new_n15577 );
xnor g13230 ( new_n15579 , new_n8501 , new_n15577 );
nor  g13231 ( new_n15580 , new_n15552 , new_n15553 );
xnor g13232 ( new_n15581 , new_n15551 , new_n15580 );
not  g13233 ( new_n15582 , new_n15581 );
nor  g13234 ( new_n15583 , new_n8503 , new_n15582 );
nor  g13235 ( new_n15584 , n18537 , new_n14991 );
or   g13236 ( new_n15585 , new_n14995 , new_n15002_1 );
and  g13237 ( new_n15586 , new_n14992 , new_n15585 );
nor  g13238 ( new_n15587 , new_n15584 , new_n15586 );
xnor g13239 ( new_n15588_1 , n1163 , new_n15582 );
and  g13240 ( new_n15589 , new_n15587 , new_n15588_1 );
nor  g13241 ( new_n15590_1 , new_n15583 , new_n15589 );
and  g13242 ( new_n15591 , new_n15579 , new_n15590_1 );
or   g13243 ( new_n15592 , new_n15578 , new_n15591 );
and  g13244 ( new_n15593 , new_n15575 , new_n15592 );
or   g13245 ( new_n15594 , new_n15573_1 , new_n15593 );
and  g13246 ( new_n15595 , new_n15570_1 , new_n15594 );
nor  g13247 ( new_n15596 , new_n15568 , new_n15595 );
xnor g13248 ( new_n15597 , new_n15565 , new_n15596 );
xnor g13249 ( new_n15598_1 , n16507 , n23250 );
not  g13250 ( new_n15599 , n11455 );
nor  g13251 ( new_n15600 , new_n15599 , n22470 );
xnor g13252 ( new_n15601 , n11455 , n22470 );
not  g13253 ( new_n15602_1 , n3945 );
nor  g13254 ( new_n15603 , new_n15602_1 , n19116 );
xnor g13255 ( new_n15604 , n3945 , n19116 );
not  g13256 ( new_n15605 , n5255 );
nor  g13257 ( new_n15606 , new_n15605 , n6861 );
xnor g13258 ( new_n15607 , n5255 , n6861 );
nor  g13259 ( new_n15608 , n19357 , new_n5163 );
xnor g13260 ( new_n15609 , n19357 , n21649 );
nor  g13261 ( new_n15610 , n2328 , new_n5166 );
not  g13262 ( new_n15611 , n15053 );
nor  g13263 ( new_n15612 , n3828 , new_n15611 );
nor  g13264 ( new_n15613 , new_n5065 , new_n5069 );
nor  g13265 ( new_n15614_1 , new_n15612 , new_n15613 );
xnor g13266 ( new_n15615 , n2328 , n18274 );
and  g13267 ( new_n15616 , new_n15614_1 , new_n15615 );
or   g13268 ( new_n15617 , new_n15610 , new_n15616 );
and  g13269 ( new_n15618 , new_n15609 , new_n15617 );
or   g13270 ( new_n15619 , new_n15608 , new_n15618 );
and  g13271 ( new_n15620 , new_n15607 , new_n15619 );
or   g13272 ( new_n15621 , new_n15606 , new_n15620 );
and  g13273 ( new_n15622 , new_n15604 , new_n15621 );
or   g13274 ( new_n15623 , new_n15603 , new_n15622 );
and  g13275 ( new_n15624 , new_n15601 , new_n15623 );
or   g13276 ( new_n15625 , new_n15600 , new_n15624 );
xor  g13277 ( new_n15626 , new_n15598_1 , new_n15625 );
nor  g13278 ( new_n15627 , n4967 , new_n15626 );
xnor g13279 ( new_n15628 , n4967 , new_n15626 );
xor  g13280 ( new_n15629 , new_n15601 , new_n15623 );
nor  g13281 ( new_n15630 , n15602 , new_n15629 );
xor  g13282 ( new_n15631 , new_n15604 , new_n15621 );
and  g13283 ( new_n15632 , n8694 , new_n15631 );
xor  g13284 ( new_n15633 , new_n15607 , new_n15619 );
nor  g13285 ( new_n15634 , n12380 , new_n15633 );
xnor g13286 ( new_n15635 , n12380 , new_n15633 );
xor  g13287 ( new_n15636_1 , new_n15609 , new_n15617 );
nor  g13288 ( new_n15637 , n8943 , new_n15636_1 );
xnor g13289 ( new_n15638 , n8943 , new_n15636_1 );
not  g13290 ( new_n15639 , new_n15638 );
not  g13291 ( new_n15640 , n8255 );
xnor g13292 ( new_n15641 , new_n15614_1 , new_n15615 );
nor  g13293 ( new_n15642 , new_n15640 , new_n15641 );
xnor g13294 ( new_n15643 , new_n5065 , new_n5069 );
and  g13295 ( new_n15644 , n11184 , new_n15643 );
not  g13296 ( new_n15645 , new_n5071 );
nor  g13297 ( new_n15646 , new_n5063 , new_n15645 );
nor  g13298 ( new_n15647 , new_n15644 , new_n15646 );
xnor g13299 ( new_n15648 , n8255 , new_n15641 );
not  g13300 ( new_n15649 , new_n15648 );
nor  g13301 ( new_n15650 , new_n15647 , new_n15649 );
nor  g13302 ( new_n15651 , new_n15642 , new_n15650 );
and  g13303 ( new_n15652_1 , new_n15639 , new_n15651 );
nor  g13304 ( new_n15653 , new_n15637 , new_n15652_1 );
nor  g13305 ( new_n15654 , new_n15635 , new_n15653 );
nor  g13306 ( new_n15655 , new_n15634 , new_n15654 );
xnor g13307 ( new_n15656 , n8694 , new_n15631 );
not  g13308 ( new_n15657 , new_n15656 );
and  g13309 ( new_n15658 , new_n15655 , new_n15657 );
nor  g13310 ( new_n15659 , new_n15632 , new_n15658 );
not  g13311 ( new_n15660 , n15602 );
xnor g13312 ( new_n15661 , new_n15660 , new_n15629 );
and  g13313 ( new_n15662_1 , new_n15659 , new_n15661 );
nor  g13314 ( new_n15663 , new_n15630 , new_n15662_1 );
nor  g13315 ( new_n15664 , new_n15628 , new_n15663 );
nor  g13316 ( new_n15665 , new_n15627 , new_n15664 );
xnor g13317 ( new_n15666 , n5101 , n6659 );
not  g13318 ( new_n15667 , n23250 );
nor  g13319 ( new_n15668 , n16507 , new_n15667 );
and  g13320 ( new_n15669 , new_n15598_1 , new_n15625 );
or   g13321 ( new_n15670 , new_n15668 , new_n15669 );
xor  g13322 ( new_n15671 , new_n15666 , new_n15670 );
xnor g13323 ( new_n15672 , n13419 , new_n15671 );
xor  g13324 ( new_n15673 , new_n15665 , new_n15672 );
xor  g13325 ( new_n15674 , new_n15597 , new_n15673 );
nor  g13326 ( new_n15675 , new_n15573_1 , new_n15593 );
xnor g13327 ( new_n15676 , new_n15570_1 , new_n15675 );
not  g13328 ( new_n15677 , new_n15676 );
xnor g13329 ( new_n15678 , new_n15628 , new_n15663 );
nor  g13330 ( new_n15679 , new_n15677 , new_n15678 );
xnor g13331 ( new_n15680 , new_n15677 , new_n15678 );
xor  g13332 ( new_n15681 , new_n15575 , new_n15592 );
not  g13333 ( new_n15682 , new_n15661 );
xnor g13334 ( new_n15683 , new_n15659 , new_n15682 );
and  g13335 ( new_n15684 , new_n15681 , new_n15683 );
xnor g13336 ( new_n15685 , new_n15681 , new_n15683 );
xnor g13337 ( new_n15686 , new_n15579 , new_n15590_1 );
xnor g13338 ( new_n15687 , new_n15655 , new_n15656 );
nor  g13339 ( new_n15688 , new_n15686 , new_n15687 );
xnor g13340 ( new_n15689 , new_n15686 , new_n15687 );
xnor g13341 ( new_n15690 , new_n15635 , new_n15653 );
xor  g13342 ( new_n15691 , new_n15587 , new_n15588_1 );
nor  g13343 ( new_n15692 , new_n15690 , new_n15691 );
xnor g13344 ( new_n15693 , new_n15690 , new_n15691 );
xnor g13345 ( new_n15694 , new_n15638 , new_n15651 );
and  g13346 ( new_n15695 , new_n15004_1 , new_n15694 );
xnor g13347 ( new_n15696 , new_n15004_1 , new_n15694 );
not  g13348 ( new_n15697 , new_n15024 );
xnor g13349 ( new_n15698 , new_n15647 , new_n15648 );
nor  g13350 ( new_n15699 , new_n15697 , new_n15698 );
xnor g13351 ( new_n15700 , new_n15697 , new_n15698 );
nor  g13352 ( new_n15701 , new_n5052 , new_n5072 );
nor  g13353 ( new_n15702 , new_n5073 , new_n5088 );
nor  g13354 ( new_n15703 , new_n15701 , new_n15702 );
nor  g13355 ( new_n15704 , new_n15700 , new_n15703 );
nor  g13356 ( new_n15705 , new_n15699 , new_n15704 );
nor  g13357 ( new_n15706 , new_n15696 , new_n15705 );
nor  g13358 ( new_n15707 , new_n15695 , new_n15706 );
nor  g13359 ( new_n15708 , new_n15693 , new_n15707 );
nor  g13360 ( new_n15709 , new_n15692 , new_n15708 );
nor  g13361 ( new_n15710 , new_n15689 , new_n15709 );
nor  g13362 ( new_n15711 , new_n15688 , new_n15710 );
nor  g13363 ( new_n15712 , new_n15685 , new_n15711 );
nor  g13364 ( new_n15713 , new_n15684 , new_n15712 );
nor  g13365 ( new_n15714 , new_n15680 , new_n15713 );
nor  g13366 ( new_n15715 , new_n15679 , new_n15714 );
xor  g13367 ( n3649 , new_n15674 , new_n15715 );
nor  g13368 ( new_n15717 , n14230 , n26625 );
not  g13369 ( new_n15718 , new_n15717 );
nor  g13370 ( new_n15719 , n26744 , new_n15718 );
not  g13371 ( new_n15720 , new_n15719 );
nor  g13372 ( new_n15721 , n11566 , new_n15720 );
not  g13373 ( new_n15722 , new_n15721 );
nor  g13374 ( new_n15723 , n3959 , new_n15722 );
not  g13375 ( new_n15724 , new_n15723 );
nor  g13376 ( new_n15725 , n26565 , new_n15724 );
xnor g13377 ( new_n15726 , n3366 , new_n15725 );
xnor g13378 ( new_n15727 , n26191 , new_n15726 );
xnor g13379 ( new_n15728 , n26565 , new_n15723 );
not  g13380 ( new_n15729 , new_n15728 );
nor  g13381 ( new_n15730 , n26512 , new_n15729 );
xnor g13382 ( new_n15731 , n26512 , new_n15728 );
not  g13383 ( new_n15732 , n19575 );
xnor g13384 ( new_n15733 , n3959 , new_n15721 );
and  g13385 ( new_n15734 , new_n15732 , new_n15733 );
xnor g13386 ( new_n15735 , n19575 , new_n15733 );
not  g13387 ( new_n15736 , n15378 );
xnor g13388 ( new_n15737 , n11566 , new_n15719 );
and  g13389 ( new_n15738 , new_n15736 , new_n15737 );
xnor g13390 ( new_n15739 , n15378 , new_n15737 );
xnor g13391 ( new_n15740 , n26744 , new_n15717 );
not  g13392 ( new_n15741 , new_n15740 );
nor  g13393 ( new_n15742 , n17095 , new_n15741 );
xnor g13394 ( new_n15743_1 , new_n9484 , n26625 );
nor  g13395 ( new_n15744 , new_n9531 , new_n15743_1 );
nor  g13396 ( new_n15745 , n14230 , new_n9532 );
xnor g13397 ( new_n15746 , n22591 , new_n15743_1 );
and  g13398 ( new_n15747 , new_n15745 , new_n15746 );
nor  g13399 ( new_n15748 , new_n15744 , new_n15747 );
xnor g13400 ( new_n15749_1 , n17095 , new_n15740 );
and  g13401 ( new_n15750 , new_n15748 , new_n15749_1 );
or   g13402 ( new_n15751 , new_n15742 , new_n15750 );
and  g13403 ( new_n15752 , new_n15739 , new_n15751 );
or   g13404 ( new_n15753 , new_n15738 , new_n15752 );
and  g13405 ( new_n15754 , new_n15735 , new_n15753 );
or   g13406 ( new_n15755 , new_n15734 , new_n15754 );
and  g13407 ( new_n15756 , new_n15731 , new_n15755 );
or   g13408 ( new_n15757 , new_n15730 , new_n15756 );
xor  g13409 ( new_n15758 , new_n15727 , new_n15757 );
xnor g13410 ( new_n15759 , n7917 , new_n15758 );
xor  g13411 ( new_n15760 , new_n15731 , new_n15755 );
and  g13412 ( new_n15761_1 , new_n14174_1 , new_n15760 );
xnor g13413 ( new_n15762_1 , n17302 , new_n15760 );
xor  g13414 ( new_n15763 , new_n15735 , new_n15753 );
nor  g13415 ( new_n15764 , new_n14177 , new_n15763 );
xnor g13416 ( new_n15765 , new_n14177 , new_n15763 );
xor  g13417 ( new_n15766_1 , new_n15739 , new_n15751 );
nor  g13418 ( new_n15767 , new_n14191 , new_n15766_1 );
xnor g13419 ( new_n15768 , new_n14191 , new_n15766_1 );
xor  g13420 ( new_n15769 , new_n15748 , new_n15749_1 );
nor  g13421 ( new_n15770 , new_n14181 , new_n15769 );
xnor g13422 ( new_n15771 , new_n14181 , new_n15769 );
xnor g13423 ( new_n15772 , new_n15745 , new_n15746 );
nor  g13424 ( new_n15773 , new_n14183 , new_n15772 );
not  g13425 ( new_n15774 , new_n15772 );
or   g13426 ( new_n15775 , n22358 , new_n15774 );
xnor g13427 ( new_n15776 , n14230 , n26167 );
and  g13428 ( new_n15777 , n9646 , new_n15776 );
and  g13429 ( new_n15778 , new_n15775 , new_n15777 );
nor  g13430 ( new_n15779 , new_n15773 , new_n15778 );
nor  g13431 ( new_n15780_1 , new_n15771 , new_n15779 );
nor  g13432 ( new_n15781 , new_n15770 , new_n15780_1 );
nor  g13433 ( new_n15782 , new_n15768 , new_n15781 );
nor  g13434 ( new_n15783 , new_n15767 , new_n15782 );
nor  g13435 ( new_n15784 , new_n15765 , new_n15783 );
nor  g13436 ( new_n15785 , new_n15764 , new_n15784 );
and  g13437 ( new_n15786 , new_n15762_1 , new_n15785 );
or   g13438 ( new_n15787 , new_n15761_1 , new_n15786 );
xor  g13439 ( new_n15788 , new_n15759 , new_n15787 );
xnor g13440 ( new_n15789 , new_n6918 , new_n15788 );
xor  g13441 ( new_n15790 , new_n15762_1 , new_n15785 );
nor  g13442 ( new_n15791 , new_n6923 , new_n15790 );
xnor g13443 ( new_n15792 , new_n6923 , new_n15790 );
xnor g13444 ( new_n15793_1 , new_n15765 , new_n15783 );
nor  g13445 ( new_n15794 , new_n6926 , new_n15793_1 );
xnor g13446 ( new_n15795 , new_n6926 , new_n15793_1 );
not  g13447 ( new_n15796 , new_n6931 );
xnor g13448 ( new_n15797 , new_n15768 , new_n15781 );
nor  g13449 ( new_n15798 , new_n15796 , new_n15797 );
xnor g13450 ( new_n15799 , new_n15796 , new_n15797 );
xnor g13451 ( new_n15800 , new_n15771 , new_n15779 );
nor  g13452 ( new_n15801 , new_n6937 , new_n15800 );
xnor g13453 ( new_n15802 , new_n6936 , new_n15800 );
xnor g13454 ( new_n15803 , n22358 , new_n15774 );
xnor g13455 ( new_n15804 , new_n15777 , new_n15803 );
nor  g13456 ( new_n15805 , new_n6943 , new_n15804 );
xnor g13457 ( new_n15806 , new_n6585 , new_n15776 );
nor  g13458 ( new_n15807 , new_n6947 , new_n15806 );
xnor g13459 ( new_n15808 , new_n6944 , new_n15804 );
and  g13460 ( new_n15809 , new_n15807 , new_n15808 );
nor  g13461 ( new_n15810 , new_n15805 , new_n15809 );
and  g13462 ( new_n15811 , new_n15802 , new_n15810 );
nor  g13463 ( new_n15812_1 , new_n15801 , new_n15811 );
nor  g13464 ( new_n15813 , new_n15799 , new_n15812_1 );
nor  g13465 ( new_n15814 , new_n15798 , new_n15813 );
nor  g13466 ( new_n15815_1 , new_n15795 , new_n15814 );
nor  g13467 ( new_n15816_1 , new_n15794 , new_n15815_1 );
nor  g13468 ( new_n15817 , new_n15792 , new_n15816_1 );
nor  g13469 ( new_n15818 , new_n15791 , new_n15817 );
xnor g13470 ( n3665 , new_n15789 , new_n15818 );
xnor g13471 ( n3679 , new_n5801 , new_n5802 );
nor  g13472 ( new_n15821 , n7139 , n16521 );
not  g13473 ( new_n15822 , new_n15821 );
nor  g13474 ( new_n15823 , n16824 , new_n15822 );
not  g13475 ( new_n15824 , new_n15823 );
nor  g13476 ( new_n15825 , n604 , new_n15824 );
not  g13477 ( new_n15826 , new_n15825 );
nor  g13478 ( new_n15827 , n4913 , new_n15826 );
not  g13479 ( new_n15828 , new_n15827 );
nor  g13480 ( new_n15829 , n9172 , new_n15828 );
not  g13481 ( new_n15830 , new_n15829 );
nor  g13482 ( new_n15831_1 , n442 , new_n15830 );
not  g13483 ( new_n15832 , new_n15831_1 );
nor  g13484 ( new_n15833 , n13719 , new_n15832 );
xnor g13485 ( new_n15834 , n7026 , new_n15833 );
xnor g13486 ( new_n15835 , new_n5921 , new_n15834 );
xnor g13487 ( new_n15836 , n13719 , new_n15831_1 );
and  g13488 ( new_n15837 , new_n5925 , new_n15836 );
not  g13489 ( new_n15838 , new_n5925 );
xnor g13490 ( new_n15839 , new_n15838 , new_n15836 );
xnor g13491 ( new_n15840 , n442 , new_n15829 );
nor  g13492 ( new_n15841 , new_n5930 , new_n15840 );
not  g13493 ( new_n15842 , new_n5930 );
xnor g13494 ( new_n15843 , new_n15842 , new_n15840 );
xnor g13495 ( new_n15844 , n9172 , new_n15827 );
nor  g13496 ( new_n15845 , new_n5935 , new_n15844 );
xnor g13497 ( new_n15846_1 , new_n13211 , new_n15844 );
xnor g13498 ( new_n15847 , n4913 , new_n15825 );
nor  g13499 ( new_n15848 , new_n5940 , new_n15847 );
xnor g13500 ( new_n15849 , new_n13213 , new_n15847 );
xnor g13501 ( new_n15850 , n604 , new_n15823 );
nor  g13502 ( new_n15851 , new_n5945 , new_n15850 );
xnor g13503 ( new_n15852 , new_n5947 , new_n15850 );
xnor g13504 ( new_n15853 , n16824 , new_n15821 );
nor  g13505 ( new_n15854 , new_n5952 , new_n15853 );
xnor g13506 ( new_n15855 , new_n5953 , new_n15853 );
nor  g13507 ( new_n15856 , new_n5956 , new_n15822 );
nor  g13508 ( new_n15857 , n7139 , new_n10777 );
xnor g13509 ( new_n15858 , new_n3560 , new_n15857 );
and  g13510 ( new_n15859_1 , new_n5959 , new_n15858 );
or   g13511 ( new_n15860 , new_n15856 , new_n15859_1 );
and  g13512 ( new_n15861 , new_n15855 , new_n15860 );
or   g13513 ( new_n15862 , new_n15854 , new_n15861 );
and  g13514 ( new_n15863 , new_n15852 , new_n15862 );
or   g13515 ( new_n15864 , new_n15851 , new_n15863 );
and  g13516 ( new_n15865 , new_n15849 , new_n15864 );
or   g13517 ( new_n15866 , new_n15848 , new_n15865 );
and  g13518 ( new_n15867 , new_n15846_1 , new_n15866 );
or   g13519 ( new_n15868 , new_n15845 , new_n15867 );
and  g13520 ( new_n15869_1 , new_n15843 , new_n15868 );
nor  g13521 ( new_n15870 , new_n15841 , new_n15869_1 );
and  g13522 ( new_n15871 , new_n15839 , new_n15870 );
or   g13523 ( new_n15872 , new_n15837 , new_n15871 );
xor  g13524 ( new_n15873 , new_n15835 , new_n15872 );
xnor g13525 ( new_n15874 , new_n4909 , new_n6029 );
nor  g13526 ( new_n15875 , new_n4913_1 , new_n6033 );
xnor g13527 ( new_n15876 , new_n4913_1 , new_n6035 );
nor  g13528 ( new_n15877 , new_n4917 , new_n6039 );
or   g13529 ( new_n15878 , new_n8477 , new_n8497 );
and  g13530 ( new_n15879 , new_n8476 , new_n15878 );
or   g13531 ( new_n15880 , new_n15877 , new_n15879 );
and  g13532 ( new_n15881 , new_n15876 , new_n15880 );
nor  g13533 ( new_n15882 , new_n15875 , new_n15881 );
xnor g13534 ( new_n15883 , new_n15874 , new_n15882 );
xnor g13535 ( new_n15884_1 , new_n15873 , new_n15883 );
xor  g13536 ( new_n15885_1 , new_n15876 , new_n15880 );
xor  g13537 ( new_n15886 , new_n15839 , new_n15870 );
nor  g13538 ( new_n15887 , new_n15885_1 , new_n15886 );
xnor g13539 ( new_n15888 , new_n15885_1 , new_n15886 );
xor  g13540 ( new_n15889_1 , new_n15843 , new_n15868 );
and  g13541 ( new_n15890 , new_n8500 , new_n15889_1 );
xnor g13542 ( new_n15891 , new_n8500 , new_n15889_1 );
xor  g13543 ( new_n15892 , new_n15846_1 , new_n15866 );
and  g13544 ( new_n15893 , new_n8531 , new_n15892 );
xnor g13545 ( new_n15894 , new_n8531 , new_n15892 );
not  g13546 ( new_n15895 , new_n8537 );
xor  g13547 ( new_n15896 , new_n15849 , new_n15864 );
and  g13548 ( new_n15897 , new_n15895 , new_n15896 );
xnor g13549 ( new_n15898 , new_n15895 , new_n15896 );
xor  g13550 ( new_n15899 , new_n15852 , new_n15862 );
and  g13551 ( new_n15900 , new_n8543 , new_n15899 );
xnor g13552 ( new_n15901 , new_n8542 , new_n15899 );
xor  g13553 ( new_n15902 , new_n15855 , new_n15860 );
nor  g13554 ( new_n15903 , new_n8547 , new_n15902 );
xnor g13555 ( new_n15904 , new_n8548 , new_n15902 );
xnor g13556 ( new_n15905 , new_n6127 , new_n15858 );
and  g13557 ( new_n15906 , new_n8552 , new_n15905 );
xnor g13558 ( new_n15907 , n7139 , new_n5956 );
and  g13559 ( new_n15908 , new_n8556 , new_n15907 );
xnor g13560 ( new_n15909 , new_n8552 , new_n15905 );
nor  g13561 ( new_n15910 , new_n15908 , new_n15909 );
nor  g13562 ( new_n15911 , new_n15906 , new_n15910 );
and  g13563 ( new_n15912 , new_n15904 , new_n15911 );
nor  g13564 ( new_n15913 , new_n15903 , new_n15912 );
and  g13565 ( new_n15914 , new_n15901 , new_n15913 );
nor  g13566 ( new_n15915 , new_n15900 , new_n15914 );
nor  g13567 ( new_n15916 , new_n15898 , new_n15915 );
nor  g13568 ( new_n15917_1 , new_n15897 , new_n15916 );
nor  g13569 ( new_n15918_1 , new_n15894 , new_n15917_1 );
nor  g13570 ( new_n15919 , new_n15893 , new_n15918_1 );
nor  g13571 ( new_n15920 , new_n15891 , new_n15919 );
nor  g13572 ( new_n15921 , new_n15890 , new_n15920 );
nor  g13573 ( new_n15922_1 , new_n15888 , new_n15921 );
nor  g13574 ( new_n15923 , new_n15887 , new_n15922_1 );
xnor g13575 ( n3725 , new_n15884_1 , new_n15923 );
nor  g13576 ( new_n15925 , n3425 , n11220 );
nor  g13577 ( new_n15926 , new_n12814 , new_n12817 );
nor  g13578 ( new_n15927 , new_n15925 , new_n15926 );
nor  g13579 ( new_n15928 , n2160 , n7335 );
and  g13580 ( new_n15929 , new_n12809 , new_n12812_1 );
nor  g13581 ( new_n15930 , new_n15928 , new_n15929 );
xnor g13582 ( new_n15931 , new_n15927 , new_n15930 );
nor  g13583 ( new_n15932 , new_n12813 , new_n12818 );
nor  g13584 ( new_n15933 , new_n12819 , new_n12822 );
nor  g13585 ( new_n15934 , new_n15932 , new_n15933 );
not  g13586 ( new_n15935 , new_n15934 );
xnor g13587 ( new_n15936_1 , new_n15931 , new_n15935 );
xnor g13588 ( new_n15937 , new_n14514 , new_n15936_1 );
nor  g13589 ( new_n15938 , new_n12824 , new_n14518 );
xnor g13590 ( new_n15939 , new_n12823 , new_n14518 );
and  g13591 ( new_n15940 , new_n5400_1 , new_n14522 );
xnor g13592 ( new_n15941 , new_n5399_1 , new_n14522 );
nor  g13593 ( new_n15942 , new_n5403_1 , new_n14526 );
not  g13594 ( new_n15943 , new_n5409 );
nor  g13595 ( new_n15944 , new_n15943 , new_n14529 );
xnor g13596 ( new_n15945 , new_n15943 , new_n14529 );
nor  g13597 ( new_n15946 , new_n5413 , new_n14444 );
xnor g13598 ( new_n15947_1 , new_n5414 , new_n14445 );
nor  g13599 ( new_n15948 , new_n4251 , new_n5418 );
nor  g13600 ( new_n15949 , new_n4258 , new_n5421 );
xnor g13601 ( new_n15950 , new_n4257 , new_n5421 );
nor  g13602 ( new_n15951 , new_n4261 , new_n5427 );
xnor g13603 ( new_n15952 , new_n4277 , new_n5427 );
nor  g13604 ( new_n15953 , new_n4264 , new_n5432 );
or   g13605 ( new_n15954 , new_n4244 , new_n5430_1 );
nor  g13606 ( new_n15955 , new_n4266_1 , new_n5436 );
and  g13607 ( new_n15956_1 , new_n15954 , new_n15955 );
or   g13608 ( new_n15957 , new_n15953 , new_n15956_1 );
and  g13609 ( new_n15958_1 , new_n15952 , new_n15957 );
or   g13610 ( new_n15959 , new_n15951 , new_n15958_1 );
and  g13611 ( new_n15960 , new_n15950 , new_n15959 );
nor  g13612 ( new_n15961 , new_n15949 , new_n15960 );
xnor g13613 ( new_n15962 , new_n14447 , new_n5418 );
and  g13614 ( new_n15963 , new_n15961 , new_n15962 );
nor  g13615 ( new_n15964 , new_n15948 , new_n15963 );
nor  g13616 ( new_n15965 , new_n15947_1 , new_n15964 );
nor  g13617 ( new_n15966 , new_n15946 , new_n15965 );
nor  g13618 ( new_n15967_1 , new_n15945 , new_n15966 );
nor  g13619 ( new_n15968 , new_n15944 , new_n15967_1 );
xnor g13620 ( new_n15969 , new_n5404 , new_n14526 );
and  g13621 ( new_n15970 , new_n15968 , new_n15969 );
or   g13622 ( new_n15971 , new_n15942 , new_n15970 );
and  g13623 ( new_n15972 , new_n15941 , new_n15971 );
nor  g13624 ( new_n15973 , new_n15940 , new_n15972 );
and  g13625 ( new_n15974 , new_n15939 , new_n15973 );
nor  g13626 ( new_n15975 , new_n15938 , new_n15974 );
xnor g13627 ( n3733 , new_n15937 , new_n15975 );
xnor g13628 ( new_n15977 , n24937 , new_n10658 );
nor  g13629 ( new_n15978 , new_n15124 , new_n10649 );
xnor g13630 ( new_n15979_1 , new_n15124 , new_n10650_1 );
and  g13631 ( new_n15980 , n3030 , new_n10640 );
or   g13632 ( new_n15981 , new_n15046 , new_n15056 );
and  g13633 ( new_n15982 , new_n15044 , new_n15981 );
or   g13634 ( new_n15983 , new_n15980 , new_n15982 );
and  g13635 ( new_n15984 , new_n15979_1 , new_n15983 );
nor  g13636 ( new_n15985 , new_n15978 , new_n15984 );
xnor g13637 ( new_n15986_1 , new_n15977 , new_n15985 );
not  g13638 ( new_n15987 , new_n15986_1 );
xnor g13639 ( new_n15988 , new_n9934_1 , new_n15987 );
nor  g13640 ( new_n15989 , new_n15980 , new_n15982 );
xnor g13641 ( new_n15990 , new_n15979_1 , new_n15989 );
nor  g13642 ( new_n15991 , new_n9939 , new_n15990 );
not  g13643 ( new_n15992 , new_n15990 );
xnor g13644 ( new_n15993 , new_n9939 , new_n15992 );
nor  g13645 ( new_n15994 , new_n9943 , new_n15058 );
and  g13646 ( new_n15995 , new_n15060 , new_n15076 );
or   g13647 ( new_n15996 , new_n15994 , new_n15995 );
and  g13648 ( new_n15997 , new_n15993 , new_n15996 );
or   g13649 ( new_n15998 , new_n15991 , new_n15997 );
xor  g13650 ( n3755 , new_n15988 , new_n15998 );
xnor g13651 ( n3758 , new_n9017 , new_n9049 );
not  g13652 ( new_n16001 , new_n15368 );
nor  g13653 ( new_n16002 , n18145 , new_n16001 );
not  g13654 ( new_n16003 , new_n16002 );
nor  g13655 ( new_n16004 , n655 , new_n16003 );
not  g13656 ( new_n16005 , new_n16004 );
nor  g13657 ( new_n16006 , n19033 , new_n16005 );
xnor g13658 ( new_n16007 , n2570 , new_n16006 );
xnor g13659 ( new_n16008 , n14692 , new_n16007 );
xnor g13660 ( new_n16009 , n19033 , new_n16004 );
nor  g13661 ( new_n16010 , new_n10170 , new_n16009 );
xnor g13662 ( new_n16011 , n4100 , new_n16009 );
xnor g13663 ( new_n16012 , n655 , new_n16002 );
nor  g13664 ( new_n16013_1 , new_n10173 , new_n16012 );
xnor g13665 ( new_n16014 , n21957 , new_n16012 );
nor  g13666 ( new_n16015 , new_n10176 , new_n15369 );
and  g13667 ( new_n16016 , new_n15370 , new_n15397 );
or   g13668 ( new_n16017 , new_n16015 , new_n16016 );
and  g13669 ( new_n16018 , new_n16014 , new_n16017 );
or   g13670 ( new_n16019 , new_n16013_1 , new_n16018 );
and  g13671 ( new_n16020 , new_n16011 , new_n16019 );
or   g13672 ( new_n16021 , new_n16010 , new_n16020 );
xor  g13673 ( new_n16022 , new_n16008 , new_n16021 );
and  g13674 ( new_n16023 , new_n11803 , new_n16022 );
xnor g13675 ( new_n16024 , new_n11803 , new_n16022 );
xor  g13676 ( new_n16025 , new_n16011 , new_n16019 );
and  g13677 ( new_n16026 , new_n6863_1 , new_n16025 );
xnor g13678 ( new_n16027 , new_n6863_1 , new_n16025 );
xor  g13679 ( new_n16028 , new_n16014 , new_n16017 );
and  g13680 ( new_n16029_1 , new_n6867_1 , new_n16028 );
xnor g13681 ( new_n16030 , new_n6867_1 , new_n16028 );
and  g13682 ( new_n16031 , new_n6872 , new_n15398 );
and  g13683 ( new_n16032 , new_n15399 , new_n15426 );
nor  g13684 ( new_n16033 , new_n16031 , new_n16032 );
nor  g13685 ( new_n16034 , new_n16030 , new_n16033 );
nor  g13686 ( new_n16035 , new_n16029_1 , new_n16034 );
nor  g13687 ( new_n16036 , new_n16027 , new_n16035 );
nor  g13688 ( new_n16037 , new_n16026 , new_n16036 );
nor  g13689 ( new_n16038 , new_n16024 , new_n16037 );
nor  g13690 ( new_n16039 , new_n16023 , new_n16038 );
not  g13691 ( new_n16040 , new_n16006 );
nor  g13692 ( new_n16041 , n2570 , new_n16040 );
xnor g13693 ( new_n16042 , n2570 , new_n16040 );
and  g13694 ( new_n16043 , n14692 , new_n16042 );
and  g13695 ( new_n16044 , new_n16008 , new_n16021 );
nor  g13696 ( new_n16045 , new_n16043 , new_n16044 );
xnor g13697 ( new_n16046 , new_n16041 , new_n16045 );
xnor g13698 ( new_n16047 , new_n11846 , new_n16046 );
xnor g13699 ( new_n16048 , new_n16039 , new_n16047 );
nor  g13700 ( new_n16049 , new_n10285 , new_n16048 );
xnor g13701 ( new_n16050 , new_n10285 , new_n16048 );
xnor g13702 ( new_n16051 , new_n16024 , new_n16037 );
nor  g13703 ( new_n16052 , new_n10342 , new_n16051 );
xnor g13704 ( new_n16053 , new_n10342 , new_n16051 );
xnor g13705 ( new_n16054 , new_n16027 , new_n16035 );
nor  g13706 ( new_n16055 , new_n10295_1 , new_n16054 );
xnor g13707 ( new_n16056 , new_n10295_1 , new_n16054 );
xnor g13708 ( new_n16057 , new_n16030 , new_n16033 );
nor  g13709 ( new_n16058 , new_n10300 , new_n16057 );
xnor g13710 ( new_n16059 , new_n10299 , new_n16057 );
nor  g13711 ( new_n16060_1 , new_n10304 , new_n15427 );
and  g13712 ( new_n16061 , new_n15428_1 , new_n15455 );
nor  g13713 ( new_n16062_1 , new_n16060_1 , new_n16061 );
and  g13714 ( new_n16063 , new_n16059 , new_n16062_1 );
nor  g13715 ( new_n16064 , new_n16058 , new_n16063 );
nor  g13716 ( new_n16065 , new_n16056 , new_n16064 );
nor  g13717 ( new_n16066 , new_n16055 , new_n16065 );
nor  g13718 ( new_n16067 , new_n16053 , new_n16066 );
nor  g13719 ( new_n16068_1 , new_n16052 , new_n16067 );
nor  g13720 ( new_n16069 , new_n16050 , new_n16068_1 );
nor  g13721 ( new_n16070 , new_n16049 , new_n16069 );
not  g13722 ( new_n16071 , new_n16070 );
nor  g13723 ( new_n16072 , new_n11846 , new_n16046 );
and  g13724 ( new_n16073 , new_n16041 , new_n16045 );
nand g13725 ( new_n16074 , new_n11846 , new_n16046 );
and  g13726 ( new_n16075 , new_n16039 , new_n16074 );
or   g13727 ( new_n16076 , new_n16073 , new_n16075 );
nor  g13728 ( new_n16077 , new_n16072 , new_n16076 );
xnor g13729 ( n3760 , new_n16071 , new_n16077 );
xnor g13730 ( n3781 , new_n3898 , new_n3922 );
xnor g13731 ( n3794 , new_n13276 , new_n13298 );
xnor g13732 ( new_n16081 , new_n3755_1 , n9246 );
and  g13733 ( new_n16082 , new_n16081 , new_n10779 );
nor  g13734 ( new_n16083 , new_n5008 , new_n16082 );
and  g13735 ( new_n16084 , new_n4777_1 , new_n16082 );
nor  g13736 ( new_n16085 , new_n16083 , new_n16084 );
nor  g13737 ( new_n16086 , new_n5956 , new_n10778 );
nor  g13738 ( new_n16087 , new_n5897 , new_n5956 );
nor  g13739 ( new_n16088 , new_n10777 , new_n5959 );
nor  g13740 ( new_n16089 , new_n16087 , new_n16088 );
xnor g13741 ( new_n16090 , new_n12869 , new_n16089 );
xnor g13742 ( new_n16091 , new_n16086 , new_n16090 );
xor  g13743 ( n3842 , new_n16085 , new_n16091 );
xnor g13744 ( n3850 , new_n8891 , new_n12085 );
xnor g13745 ( n3869 , new_n4297 , new_n14469 );
xnor g13746 ( new_n16095 , n919 , n21749 );
nor  g13747 ( new_n16096 , n7769 , n25316 );
or   g13748 ( new_n16097 , new_n4146_1 , new_n9485 );
xnor g13749 ( new_n16098_1 , new_n9487 , n25316 );
and  g13750 ( new_n16099 , new_n16097 , new_n16098_1 );
nor  g13751 ( new_n16100 , new_n16096 , new_n16099 );
xnor g13752 ( new_n16101 , new_n16095 , new_n16100 );
xnor g13753 ( new_n16102 , n19584 , new_n16101 );
not  g13754 ( new_n16103 , n15332 );
xnor g13755 ( new_n16104 , new_n4146_1 , n21138 );
nor  g13756 ( new_n16105 , new_n16103 , new_n16104 );
nor  g13757 ( new_n16106 , n5060 , new_n16105 );
xor  g13758 ( new_n16107 , new_n16097 , new_n16098_1 );
xnor g13759 ( new_n16108 , n5060 , new_n16105 );
nor  g13760 ( new_n16109 , new_n16107 , new_n16108 );
nor  g13761 ( new_n16110_1 , new_n16106 , new_n16109 );
xnor g13762 ( new_n16111 , new_n16102 , new_n16110_1 );
xnor g13763 ( new_n16112 , new_n15301 , new_n16111 );
xor  g13764 ( new_n16113 , new_n16107 , new_n16108 );
nor  g13765 ( new_n16114 , new_n15305 , new_n16113 );
xnor g13766 ( new_n16115 , n15332 , new_n16104 );
nor  g13767 ( new_n16116 , new_n15309 , new_n16115 );
xnor g13768 ( new_n16117 , new_n15305 , new_n16113 );
nor  g13769 ( new_n16118 , new_n16116 , new_n16117 );
nor  g13770 ( new_n16119 , new_n16114 , new_n16118 );
xnor g13771 ( n3871 , new_n16112 , new_n16119 );
xor  g13772 ( n3891 , new_n15904 , new_n15911 );
xnor g13773 ( new_n16122 , n2570 , n10250 );
nor  g13774 ( new_n16123 , new_n6155 , n19033 );
xnor g13775 ( new_n16124 , n7674 , n19033 );
nor  g13776 ( new_n16125 , n655 , new_n6158 );
xnor g13777 ( new_n16126 , n655 , n6397 );
nor  g13778 ( new_n16127 , n18145 , new_n6161 );
xnor g13779 ( new_n16128 , n18145 , n19196 );
nor  g13780 ( new_n16129 , n10712 , new_n11812 );
xnor g13781 ( new_n16130 , n10712 , n23586 );
nor  g13782 ( new_n16131 , new_n15238 , n25126 );
xnor g13783 ( new_n16132 , n21226 , n25126 );
nor  g13784 ( new_n16133 , new_n6170 , n19608 );
not  g13785 ( new_n16134 , n1689 );
nor  g13786 ( new_n16135 , new_n16134 , n20036 );
or   g13787 ( new_n16136 , new_n4119_1 , new_n4125 );
and  g13788 ( new_n16137 , new_n4117 , new_n16136 );
nor  g13789 ( new_n16138 , new_n16135 , new_n16137 );
xnor g13790 ( new_n16139 , n4426 , n19608 );
and  g13791 ( new_n16140 , new_n16138 , new_n16139 );
or   g13792 ( new_n16141 , new_n16133 , new_n16140 );
and  g13793 ( new_n16142_1 , new_n16132 , new_n16141 );
or   g13794 ( new_n16143 , new_n16131 , new_n16142_1 );
and  g13795 ( new_n16144 , new_n16130 , new_n16143 );
or   g13796 ( new_n16145 , new_n16129 , new_n16144 );
and  g13797 ( new_n16146 , new_n16128 , new_n16145 );
or   g13798 ( new_n16147 , new_n16127 , new_n16146 );
and  g13799 ( new_n16148 , new_n16126 , new_n16147 );
or   g13800 ( new_n16149 , new_n16125 , new_n16148 );
and  g13801 ( new_n16150 , new_n16124 , new_n16149 );
or   g13802 ( new_n16151 , new_n16123 , new_n16150 );
xor  g13803 ( new_n16152 , new_n16122 , new_n16151 );
xnor g13804 ( new_n16153 , new_n11802 , new_n16152 );
xor  g13805 ( new_n16154 , new_n16124 , new_n16149 );
nor  g13806 ( new_n16155 , new_n6864 , new_n16154 );
xnor g13807 ( new_n16156 , new_n6863_1 , new_n16154 );
xor  g13808 ( new_n16157 , new_n16126 , new_n16147 );
nor  g13809 ( new_n16158_1 , new_n6869 , new_n16157 );
xnor g13810 ( new_n16159 , new_n6867_1 , new_n16157 );
xor  g13811 ( new_n16160 , new_n16128 , new_n16145 );
nor  g13812 ( new_n16161 , new_n6874 , new_n16160 );
xnor g13813 ( new_n16162 , new_n6872 , new_n16160 );
xor  g13814 ( new_n16163 , new_n16130 , new_n16143 );
nor  g13815 ( new_n16164 , new_n6879 , new_n16163 );
xnor g13816 ( new_n16165 , new_n6877 , new_n16163 );
xor  g13817 ( new_n16166 , new_n16132 , new_n16141 );
nor  g13818 ( new_n16167_1 , new_n6881 , new_n16166 );
xnor g13819 ( new_n16168 , new_n6881 , new_n16166 );
xnor g13820 ( new_n16169 , new_n16138 , new_n16139 );
not  g13821 ( new_n16170 , new_n16169 );
nor  g13822 ( new_n16171 , new_n6888 , new_n16170 );
xnor g13823 ( new_n16172 , new_n6888 , new_n16169 );
not  g13824 ( new_n16173 , new_n4127 );
nor  g13825 ( new_n16174 , new_n4116 , new_n16173 );
and  g13826 ( new_n16175 , new_n4128 , new_n4141 );
or   g13827 ( new_n16176 , new_n16174 , new_n16175 );
and  g13828 ( new_n16177 , new_n16172 , new_n16176 );
nor  g13829 ( new_n16178 , new_n16171 , new_n16177 );
nor  g13830 ( new_n16179 , new_n16168 , new_n16178 );
or   g13831 ( new_n16180 , new_n16167_1 , new_n16179 );
and  g13832 ( new_n16181 , new_n16165 , new_n16180 );
or   g13833 ( new_n16182 , new_n16164 , new_n16181 );
and  g13834 ( new_n16183 , new_n16162 , new_n16182 );
or   g13835 ( new_n16184 , new_n16161 , new_n16183 );
and  g13836 ( new_n16185_1 , new_n16159 , new_n16184 );
or   g13837 ( new_n16186 , new_n16158_1 , new_n16185_1 );
and  g13838 ( new_n16187 , new_n16156 , new_n16186 );
nor  g13839 ( new_n16188 , new_n16155 , new_n16187 );
xnor g13840 ( new_n16189 , new_n16153 , new_n16188 );
xnor g13841 ( new_n16190 , new_n6361 , new_n16189 );
xor  g13842 ( new_n16191 , new_n16156 , new_n16186 );
and  g13843 ( new_n16192 , new_n6368 , new_n16191 );
xnor g13844 ( new_n16193 , new_n6368 , new_n16191 );
not  g13845 ( new_n16194 , new_n6373 );
xor  g13846 ( new_n16195 , new_n16159 , new_n16184 );
and  g13847 ( new_n16196_1 , new_n16194 , new_n16195 );
xnor g13848 ( new_n16197 , new_n16194 , new_n16195 );
xor  g13849 ( new_n16198 , new_n16162 , new_n16182 );
and  g13850 ( new_n16199 , new_n6377 , new_n16198 );
xnor g13851 ( new_n16200 , new_n6377 , new_n16198 );
xor  g13852 ( new_n16201 , new_n16165 , new_n16180 );
and  g13853 ( new_n16202 , new_n6382 , new_n16201 );
xnor g13854 ( new_n16203 , new_n6382 , new_n16201 );
xnor g13855 ( new_n16204 , new_n16168 , new_n16178 );
nor  g13856 ( new_n16205 , new_n6386 , new_n16204 );
xnor g13857 ( new_n16206_1 , new_n6386 , new_n16204 );
not  g13858 ( new_n16207 , new_n6391 );
xor  g13859 ( new_n16208 , new_n16172 , new_n16176 );
and  g13860 ( new_n16209 , new_n16207 , new_n16208 );
xnor g13861 ( new_n16210 , new_n16207 , new_n16208 );
nor  g13862 ( new_n16211 , new_n4142 , new_n4151_1 );
nor  g13863 ( new_n16212 , new_n4152_1 , new_n4163 );
nor  g13864 ( new_n16213 , new_n16211 , new_n16212 );
nor  g13865 ( new_n16214 , new_n16210 , new_n16213 );
nor  g13866 ( new_n16215_1 , new_n16209 , new_n16214 );
nor  g13867 ( new_n16216 , new_n16206_1 , new_n16215_1 );
nor  g13868 ( new_n16217_1 , new_n16205 , new_n16216 );
nor  g13869 ( new_n16218_1 , new_n16203 , new_n16217_1 );
nor  g13870 ( new_n16219_1 , new_n16202 , new_n16218_1 );
nor  g13871 ( new_n16220 , new_n16200 , new_n16219_1 );
nor  g13872 ( new_n16221 , new_n16199 , new_n16220 );
nor  g13873 ( new_n16222 , new_n16197 , new_n16221 );
nor  g13874 ( new_n16223_1 , new_n16196_1 , new_n16222 );
nor  g13875 ( new_n16224 , new_n16193 , new_n16223_1 );
nor  g13876 ( new_n16225 , new_n16192 , new_n16224 );
xnor g13877 ( n3932 , new_n16190 , new_n16225 );
xnor g13878 ( n3934 , new_n3915 , new_n3916 );
xnor g13879 ( n3971 , new_n4095 , new_n4096 );
nor  g13880 ( new_n16229 , n5026 , n8581 );
not  g13881 ( new_n16230_1 , new_n16229 );
nor  g13882 ( new_n16231 , n12161 , new_n16230_1 );
not  g13883 ( new_n16232 , new_n16231 );
nor  g13884 ( new_n16233 , n18157 , new_n16232 );
not  g13885 ( new_n16234 , new_n16233 );
nor  g13886 ( new_n16235 , n20923 , new_n16234 );
not  g13887 ( new_n16236 , new_n16235 );
nor  g13888 ( new_n16237 , n8067 , new_n16236 );
not  g13889 ( new_n16238 , new_n16237 );
nor  g13890 ( new_n16239 , n10125 , new_n16238 );
not  g13891 ( new_n16240 , new_n16239 );
nor  g13892 ( new_n16241 , n25240 , new_n16240 );
xnor g13893 ( new_n16242 , n1222 , new_n16241 );
xnor g13894 ( new_n16243_1 , new_n8789 , new_n16242 );
xnor g13895 ( new_n16244 , n25240 , new_n16239 );
nor  g13896 ( new_n16245 , n3710 , new_n16244 );
xnor g13897 ( new_n16246 , new_n9992 , new_n16244 );
xnor g13898 ( new_n16247_1 , n10125 , new_n16237 );
and  g13899 ( new_n16248 , n26318 , new_n16247_1 );
or   g13900 ( new_n16249 , n26318 , new_n16247_1 );
xnor g13901 ( new_n16250 , n8067 , new_n16235 );
nor  g13902 ( new_n16251 , n26054 , new_n16250 );
xnor g13903 ( new_n16252 , new_n8749 , new_n16250 );
xnor g13904 ( new_n16253 , n20923 , new_n16233 );
nor  g13905 ( new_n16254 , n19081 , new_n16253 );
xnor g13906 ( new_n16255 , new_n8753 , new_n16253 );
xnor g13907 ( new_n16256 , n18157 , new_n16231 );
nor  g13908 ( new_n16257 , n8309 , new_n16256 );
xnor g13909 ( new_n16258 , n12161 , new_n16229 );
nor  g13910 ( new_n16259 , n19144 , new_n16258 );
xnor g13911 ( new_n16260 , new_n8759 , new_n16258 );
xnor g13912 ( new_n16261 , new_n7220 , n8581 );
nor  g13913 ( new_n16262 , n12593 , new_n16261 );
or   g13914 ( new_n16263 , new_n6628_1 , new_n8763 );
xnor g13915 ( new_n16264 , new_n10007 , new_n16261 );
and  g13916 ( new_n16265 , new_n16263 , new_n16264 );
or   g13917 ( new_n16266 , new_n16262 , new_n16265 );
and  g13918 ( new_n16267 , new_n16260 , new_n16266 );
or   g13919 ( new_n16268 , new_n16259 , new_n16267 );
xnor g13920 ( new_n16269 , new_n8771 , new_n16256 );
and  g13921 ( new_n16270 , new_n16268 , new_n16269 );
or   g13922 ( new_n16271 , new_n16257 , new_n16270 );
and  g13923 ( new_n16272 , new_n16255 , new_n16271 );
or   g13924 ( new_n16273 , new_n16254 , new_n16272 );
and  g13925 ( new_n16274 , new_n16252 , new_n16273 );
nor  g13926 ( new_n16275_1 , new_n16251 , new_n16274 );
and  g13927 ( new_n16276 , new_n16249 , new_n16275_1 );
nor  g13928 ( new_n16277 , new_n16248 , new_n16276 );
and  g13929 ( new_n16278 , new_n16246 , new_n16277 );
or   g13930 ( new_n16279_1 , new_n16245 , new_n16278 );
xor  g13931 ( new_n16280 , new_n16243_1 , new_n16279_1 );
xnor g13932 ( new_n16281 , n26797 , new_n16280 );
xnor g13933 ( new_n16282 , new_n16246 , new_n16277 );
not  g13934 ( new_n16283 , new_n16282 );
nor  g13935 ( new_n16284 , new_n8033 , new_n16283 );
xnor g13936 ( new_n16285 , n23913 , new_n16283 );
xnor g13937 ( new_n16286 , new_n8745_1 , new_n16247_1 );
xnor g13938 ( new_n16287 , new_n16275_1 , new_n16286 );
nor  g13939 ( new_n16288 , new_n8036 , new_n16287 );
not  g13940 ( new_n16289 , new_n16287 );
xnor g13941 ( new_n16290 , new_n8036 , new_n16289 );
nor  g13942 ( new_n16291 , new_n16254 , new_n16272 );
xnor g13943 ( new_n16292 , new_n16252 , new_n16291 );
nor  g13944 ( new_n16293 , new_n8039 , new_n16292 );
not  g13945 ( new_n16294 , new_n16292 );
xnor g13946 ( new_n16295 , new_n8039 , new_n16294 );
xor  g13947 ( new_n16296 , new_n16255 , new_n16271 );
nor  g13948 ( new_n16297 , new_n8042_1 , new_n16296 );
xnor g13949 ( new_n16298 , n3909 , new_n16296 );
xor  g13950 ( new_n16299 , new_n16268 , new_n16269 );
nor  g13951 ( new_n16300 , new_n8045 , new_n16299 );
xnor g13952 ( new_n16301 , n23974 , new_n16299 );
xor  g13953 ( new_n16302 , new_n16260 , new_n16266 );
nor  g13954 ( new_n16303 , new_n8050 , new_n16302 );
xnor g13955 ( new_n16304 , n2146 , new_n16302 );
xor  g13956 ( new_n16305 , new_n16263 , new_n16264 );
nor  g13957 ( new_n16306 , new_n8055 , new_n16305 );
xnor g13958 ( new_n16307 , n8581 , n13714 );
nor  g13959 ( new_n16308 , new_n5587 , new_n16307 );
xnor g13960 ( new_n16309 , n22173 , new_n16305 );
and  g13961 ( new_n16310 , new_n16308 , new_n16309 );
or   g13962 ( new_n16311 , new_n16306 , new_n16310 );
and  g13963 ( new_n16312 , new_n16304 , new_n16311 );
or   g13964 ( new_n16313 , new_n16303 , new_n16312 );
and  g13965 ( new_n16314 , new_n16301 , new_n16313 );
or   g13966 ( new_n16315 , new_n16300 , new_n16314 );
and  g13967 ( new_n16316 , new_n16298 , new_n16315 );
or   g13968 ( new_n16317 , new_n16297 , new_n16316 );
and  g13969 ( new_n16318 , new_n16295 , new_n16317 );
or   g13970 ( new_n16319 , new_n16293 , new_n16318 );
and  g13971 ( new_n16320 , new_n16290 , new_n16319 );
or   g13972 ( new_n16321 , new_n16288 , new_n16320 );
and  g13973 ( new_n16322_1 , new_n16285 , new_n16321 );
nor  g13974 ( new_n16323 , new_n16284 , new_n16322_1 );
xnor g13975 ( new_n16324 , new_n16281 , new_n16323 );
xnor g13976 ( new_n16325 , new_n8144 , new_n16324 );
xor  g13977 ( new_n16326 , new_n16285 , new_n16321 );
nor  g13978 ( new_n16327_1 , new_n8149_1 , new_n16326 );
xnor g13979 ( new_n16328 , new_n8149_1 , new_n16326 );
xor  g13980 ( new_n16329 , new_n16290 , new_n16319 );
nor  g13981 ( new_n16330 , new_n8154 , new_n16329 );
xnor g13982 ( new_n16331 , new_n8154 , new_n16329 );
not  g13983 ( new_n16332 , new_n8159_1 );
xor  g13984 ( new_n16333 , new_n16295 , new_n16317 );
nor  g13985 ( new_n16334 , new_n16332 , new_n16333 );
xnor g13986 ( new_n16335 , new_n16332 , new_n16333 );
xor  g13987 ( new_n16336 , new_n16298 , new_n16315 );
nor  g13988 ( new_n16337 , new_n8164 , new_n16336 );
xnor g13989 ( new_n16338 , new_n8164 , new_n16336 );
xor  g13990 ( new_n16339 , new_n16301 , new_n16313 );
nor  g13991 ( new_n16340 , new_n8168 , new_n16339 );
xnor g13992 ( new_n16341 , new_n8168 , new_n16339 );
xor  g13993 ( new_n16342 , new_n16304 , new_n16311 );
nor  g13994 ( new_n16343 , new_n8173 , new_n16342 );
xor  g13995 ( new_n16344 , new_n16308 , new_n16309 );
nor  g13996 ( new_n16345 , new_n8183 , new_n16344 );
xnor g13997 ( new_n16346 , n583 , new_n16307 );
and  g13998 ( new_n16347 , new_n8181 , new_n16346 );
xnor g13999 ( new_n16348 , new_n8183 , new_n16344 );
nor  g14000 ( new_n16349 , new_n16347 , new_n16348 );
nor  g14001 ( new_n16350_1 , new_n16345 , new_n16349 );
xnor g14002 ( new_n16351 , new_n8173 , new_n16342 );
nor  g14003 ( new_n16352 , new_n16350_1 , new_n16351 );
nor  g14004 ( new_n16353 , new_n16343 , new_n16352 );
nor  g14005 ( new_n16354 , new_n16341 , new_n16353 );
nor  g14006 ( new_n16355 , new_n16340 , new_n16354 );
nor  g14007 ( new_n16356 , new_n16338 , new_n16355 );
nor  g14008 ( new_n16357 , new_n16337 , new_n16356 );
nor  g14009 ( new_n16358 , new_n16335 , new_n16357 );
nor  g14010 ( new_n16359 , new_n16334 , new_n16358 );
nor  g14011 ( new_n16360 , new_n16331 , new_n16359 );
nor  g14012 ( new_n16361 , new_n16330 , new_n16360 );
nor  g14013 ( new_n16362 , new_n16328 , new_n16361 );
nor  g14014 ( new_n16363 , new_n16327_1 , new_n16362 );
xnor g14015 ( n3983 , new_n16325 , new_n16363 );
not  g14016 ( new_n16365 , new_n6666 );
xnor g14017 ( new_n16366 , n583 , n13714 );
xnor g14018 ( new_n16367_1 , n6611 , new_n16366 );
nor  g14019 ( new_n16368 , new_n16365 , new_n16367_1 );
or   g14020 ( new_n16369 , new_n5588 , new_n16366 );
nor  g14021 ( new_n16370 , new_n5587 , new_n8763 );
xnor g14022 ( new_n16371 , n12593 , n22173 );
xnor g14023 ( new_n16372 , new_n16370 , new_n16371 );
xnor g14024 ( new_n16373 , new_n5584 , new_n16372 );
xor  g14025 ( new_n16374 , new_n16369 , new_n16373 );
xnor g14026 ( new_n16375 , new_n16368 , new_n16374 );
xnor g14027 ( n4000 , new_n6662 , new_n16375 );
xnor g14028 ( new_n16377 , n20179 , n26823 );
nor  g14029 ( new_n16378 , new_n5280 , n19228 );
xnor g14030 ( new_n16379_1 , n4812 , n19228 );
nor  g14031 ( new_n16380 , n15539 , new_n8394 );
xnor g14032 ( new_n16381 , n15539 , n24278 );
nor  g14033 ( new_n16382 , n8052 , new_n8398 );
or   g14034 ( new_n16383 , new_n6767 , n24618 );
nor  g14035 ( new_n16384 , n3952 , new_n7448 );
and  g14036 ( new_n16385 , new_n11149 , new_n11150 );
nor  g14037 ( new_n16386 , new_n16384 , new_n16385 );
and  g14038 ( new_n16387 , new_n16383 , new_n16386 );
or   g14039 ( new_n16388 , new_n16382 , new_n16387 );
and  g14040 ( new_n16389 , new_n16381 , new_n16388 );
or   g14041 ( new_n16390 , new_n16380 , new_n16389 );
and  g14042 ( new_n16391 , new_n16379_1 , new_n16390 );
or   g14043 ( new_n16392 , new_n16378 , new_n16391 );
xor  g14044 ( new_n16393 , new_n16377 , new_n16392 );
xnor g14045 ( new_n16394 , new_n7381 , new_n16393 );
xor  g14046 ( new_n16395 , new_n16379_1 , new_n16390 );
nor  g14047 ( new_n16396_1 , new_n7385 , new_n16395 );
xnor g14048 ( new_n16397 , new_n7385 , new_n16395 );
not  g14049 ( new_n16398_1 , new_n7389 );
xor  g14050 ( new_n16399 , new_n16381 , new_n16388 );
nor  g14051 ( new_n16400 , new_n16398_1 , new_n16399 );
xnor g14052 ( new_n16401 , n8052 , n24618 );
xnor g14053 ( new_n16402 , new_n16386 , new_n16401 );
and  g14054 ( new_n16403 , new_n7393 , new_n16402 );
xnor g14055 ( new_n16404 , new_n7392 , new_n16402 );
and  g14056 ( new_n16405 , new_n11148 , new_n11151 );
nor  g14057 ( new_n16406_1 , new_n7406 , new_n11152 );
nor  g14058 ( new_n16407_1 , new_n16405 , new_n16406_1 );
and  g14059 ( new_n16408 , new_n16404 , new_n16407_1 );
nor  g14060 ( new_n16409 , new_n16403 , new_n16408 );
xnor g14061 ( new_n16410 , new_n16398_1 , new_n16399 );
nor  g14062 ( new_n16411 , new_n16409 , new_n16410 );
nor  g14063 ( new_n16412 , new_n16400 , new_n16411 );
nor  g14064 ( new_n16413 , new_n16397 , new_n16412 );
nor  g14065 ( new_n16414 , new_n16396_1 , new_n16413 );
xnor g14066 ( n4010 , new_n16394 , new_n16414 );
xnor g14067 ( new_n16416 , n2160 , n11220 );
nor  g14068 ( new_n16417 , new_n11674_1 , n22379 );
xnor g14069 ( new_n16418 , n10763 , n22379 );
nor  g14070 ( new_n16419_1 , n1662 , new_n2890 );
xnor g14071 ( new_n16420 , n1662 , n7437 );
nor  g14072 ( new_n16421 , n12875 , new_n2893 );
nor  g14073 ( new_n16422 , n2035 , new_n2896 );
and  g14074 ( new_n16423 , new_n14415 , new_n14433 );
or   g14075 ( new_n16424_1 , new_n16422 , new_n16423 );
xnor g14076 ( new_n16425 , n12875 , n20700 );
and  g14077 ( new_n16426 , new_n16424_1 , new_n16425 );
or   g14078 ( new_n16427 , new_n16421 , new_n16426 );
and  g14079 ( new_n16428_1 , new_n16420 , new_n16427 );
or   g14080 ( new_n16429 , new_n16419_1 , new_n16428_1 );
and  g14081 ( new_n16430 , new_n16418 , new_n16429 );
or   g14082 ( new_n16431 , new_n16417 , new_n16430 );
xor  g14083 ( new_n16432 , new_n16416 , new_n16431 );
xnor g14084 ( new_n16433_1 , new_n14588 , new_n16432 );
xor  g14085 ( new_n16434 , new_n16418 , new_n16429 );
nor  g14086 ( new_n16435 , new_n14597 , new_n16434 );
xnor g14087 ( new_n16436 , new_n14597 , new_n16434 );
xor  g14088 ( new_n16437 , new_n16420 , new_n16427 );
nor  g14089 ( new_n16438 , new_n14601 , new_n16437 );
xor  g14090 ( new_n16439_1 , new_n16424_1 , new_n16425 );
not  g14091 ( new_n16440_1 , new_n16439_1 );
nor  g14092 ( new_n16441 , new_n14606 , new_n16440_1 );
xnor g14093 ( new_n16442 , new_n14606 , new_n16439_1 );
and  g14094 ( new_n16443 , new_n14434 , new_n14451 );
and  g14095 ( new_n16444 , new_n14453 , new_n14478 );
or   g14096 ( new_n16445_1 , new_n16443 , new_n16444 );
and  g14097 ( new_n16446 , new_n16442 , new_n16445_1 );
nor  g14098 ( new_n16447 , new_n16441 , new_n16446 );
xnor g14099 ( new_n16448 , new_n14604 , new_n16437 );
and  g14100 ( new_n16449 , new_n16447 , new_n16448 );
nor  g14101 ( new_n16450 , new_n16438 , new_n16449 );
nor  g14102 ( new_n16451 , new_n16436 , new_n16450 );
nor  g14103 ( new_n16452 , new_n16435 , new_n16451 );
xor  g14104 ( n4014 , new_n16433_1 , new_n16452 );
xnor g14105 ( new_n16454 , new_n11636 , new_n13881 );
nor  g14106 ( new_n16455 , n26224 , new_n13884 );
xnor g14107 ( new_n16456 , new_n12526 , new_n13884 );
nor  g14108 ( new_n16457 , n19327 , new_n3736 );
or   g14109 ( new_n16458 , new_n3739 , new_n3769 );
and  g14110 ( new_n16459 , new_n3737 , new_n16458 );
or   g14111 ( new_n16460_1 , new_n16457 , new_n16459 );
and  g14112 ( new_n16461 , new_n16456 , new_n16460_1 );
nor  g14113 ( new_n16462 , new_n16455 , new_n16461 );
xnor g14114 ( new_n16463 , new_n16454 , new_n16462 );
not  g14115 ( new_n16464 , new_n16463 );
xnor g14116 ( new_n16465 , new_n4801 , new_n16464 );
nor  g14117 ( new_n16466 , new_n16457 , new_n16459 );
xnor g14118 ( new_n16467 , new_n16456 , new_n16466 );
nor  g14119 ( new_n16468 , new_n7328 , new_n16467 );
not  g14120 ( new_n16469 , new_n16467 );
xnor g14121 ( new_n16470 , new_n7328 , new_n16469 );
nor  g14122 ( new_n16471 , new_n3725_1 , new_n3771 );
and  g14123 ( new_n16472 , new_n3773 , new_n3812 );
or   g14124 ( new_n16473 , new_n16471 , new_n16472 );
and  g14125 ( new_n16474 , new_n16470 , new_n16473 );
or   g14126 ( new_n16475 , new_n16468 , new_n16474 );
xor  g14127 ( new_n16476_1 , new_n16465 , new_n16475 );
xnor g14128 ( new_n16477 , new_n11745 , new_n16476_1 );
xor  g14129 ( new_n16478 , new_n16470 , new_n16473 );
nor  g14130 ( new_n16479 , new_n11750 , new_n16478 );
xnor g14131 ( new_n16480 , new_n11750 , new_n16478 );
nor  g14132 ( new_n16481_1 , new_n3813 , new_n3889 );
nor  g14133 ( new_n16482_1 , new_n3890 , new_n3926 );
nor  g14134 ( new_n16483 , new_n16481_1 , new_n16482_1 );
nor  g14135 ( new_n16484 , new_n16480 , new_n16483 );
nor  g14136 ( new_n16485 , new_n16479 , new_n16484 );
xnor g14137 ( n4071 , new_n16477 , new_n16485 );
xnor g14138 ( n4088 , new_n12713 , new_n12718 );
not  g14139 ( new_n16488 , n7593 );
and  g14140 ( new_n16489 , new_n16488 , new_n12826 );
nor  g14141 ( new_n16490 , n5025 , new_n12827 );
and  g14142 ( new_n16491 , n5025 , new_n12827 );
nor  g14143 ( new_n16492 , new_n16491 , new_n12831 );
nor  g14144 ( new_n16493_1 , new_n16490 , new_n16492 );
nor  g14145 ( new_n16494 , new_n16489 , new_n16493_1 );
not  g14146 ( new_n16495 , new_n16494 );
not  g14147 ( new_n16496 , new_n15927 );
nor  g14148 ( new_n16497 , new_n16496 , new_n15930 );
and  g14149 ( new_n16498 , new_n16496 , new_n15930 );
nor  g14150 ( new_n16499 , new_n16498 , new_n15935 );
nor  g14151 ( new_n16500 , new_n16497 , new_n16499 );
not  g14152 ( new_n16501 , new_n16500 );
nor  g14153 ( new_n16502_1 , new_n16495 , new_n16501 );
not  g14154 ( new_n16503 , new_n15936_1 );
nor  g14155 ( new_n16504 , new_n16503 , new_n16494 );
or   g14156 ( new_n16505 , new_n15936_1 , new_n16495 );
nor  g14157 ( new_n16506_1 , new_n12823 , new_n12832 );
and  g14158 ( new_n16507_1 , new_n12833 , new_n12836 );
nor  g14159 ( new_n16508 , new_n16506_1 , new_n16507_1 );
and  g14160 ( new_n16509 , new_n16505 , new_n16508 );
nor  g14161 ( new_n16510 , new_n16504 , new_n16509 );
nor  g14162 ( new_n16511 , new_n16502_1 , new_n16510 );
nor  g14163 ( new_n16512 , new_n16494 , new_n16500 );
nor  g14164 ( new_n16513 , new_n16509 , new_n16512 );
nor  g14165 ( n4089 , new_n16511 , new_n16513 );
not  g14166 ( new_n16515 , new_n11950 );
nor  g14167 ( new_n16516_1 , n1112 , new_n16515 );
xnor g14168 ( new_n16517_1 , n2289 , new_n16516_1 );
not  g14169 ( new_n16518 , new_n16517_1 );
xnor g14170 ( new_n16519 , n3228 , new_n16518 );
nor  g14171 ( new_n16520 , n5302 , new_n11951 );
xnor g14172 ( new_n16521_1 , n5302 , new_n11951 );
and  g14173 ( new_n16522 , n25738 , new_n11954 );
or   g14174 ( new_n16523 , n25738 , new_n11954 );
nor  g14175 ( new_n16524_1 , n21471 , new_n8578 );
not  g14176 ( new_n16525 , new_n8598 );
nor  g14177 ( new_n16526 , new_n8579 , new_n16525 );
nor  g14178 ( new_n16527_1 , new_n16524_1 , new_n16526 );
and  g14179 ( new_n16528 , new_n16523 , new_n16527_1 );
nor  g14180 ( new_n16529 , new_n16522 , new_n16528 );
not  g14181 ( new_n16530 , new_n16529 );
nor  g14182 ( new_n16531 , new_n16521_1 , new_n16530 );
nor  g14183 ( new_n16532 , new_n16520 , new_n16531 );
xnor g14184 ( new_n16533 , new_n16519 , new_n16532 );
not  g14185 ( new_n16534 , new_n16533 );
xnor g14186 ( new_n16535 , n13775 , new_n16534 );
xnor g14187 ( new_n16536 , new_n16521_1 , new_n16529 );
not  g14188 ( new_n16537 , new_n16536 );
nor  g14189 ( new_n16538 , n1293 , new_n16537 );
xnor g14190 ( new_n16539 , new_n6839 , new_n16537 );
xnor g14191 ( new_n16540 , n25738 , new_n11955 );
xnor g14192 ( new_n16541 , new_n16527_1 , new_n16540 );
nor  g14193 ( new_n16542 , new_n6842 , new_n16541 );
nor  g14194 ( new_n16543 , new_n8572 , new_n8599 );
and  g14195 ( new_n16544_1 , new_n8601 , new_n8622 );
or   g14196 ( new_n16545 , new_n16543 , new_n16544_1 );
xnor g14197 ( new_n16546 , n19042 , new_n16541 );
and  g14198 ( new_n16547 , new_n16545 , new_n16546 );
nor  g14199 ( new_n16548 , new_n16542 , new_n16547 );
and  g14200 ( new_n16549 , new_n16539 , new_n16548 );
nor  g14201 ( new_n16550 , new_n16538 , new_n16549 );
xnor g14202 ( new_n16551 , new_n16535 , new_n16550 );
xnor g14203 ( new_n16552 , new_n5459 , new_n7533 );
nor  g14204 ( new_n16553 , new_n5462 , new_n2460 );
xnor g14205 ( new_n16554_1 , new_n5462 , new_n2460 );
nor  g14206 ( new_n16555 , new_n5465 , new_n2463 );
xnor g14207 ( new_n16556 , new_n5465 , new_n2463 );
nor  g14208 ( new_n16557 , new_n5468 , new_n2466 );
nor  g14209 ( new_n16558 , new_n6681 , new_n6695 );
nor  g14210 ( new_n16559 , new_n16557 , new_n16558 );
nor  g14211 ( new_n16560 , new_n16556 , new_n16559 );
nor  g14212 ( new_n16561 , new_n16555 , new_n16560 );
nor  g14213 ( new_n16562 , new_n16554_1 , new_n16561 );
nor  g14214 ( new_n16563 , new_n16553 , new_n16562 );
xor  g14215 ( new_n16564 , new_n16552 , new_n16563 );
xnor g14216 ( new_n16565 , new_n16551 , new_n16564 );
xnor g14217 ( new_n16566 , new_n16539 , new_n16548 );
xor  g14218 ( new_n16567 , new_n16554_1 , new_n16561 );
nor  g14219 ( new_n16568 , new_n16566 , new_n16567 );
xnor g14220 ( new_n16569 , new_n16566 , new_n16567 );
xnor g14221 ( new_n16570 , new_n16556 , new_n16559 );
not  g14222 ( new_n16571 , new_n16570 );
xor  g14223 ( new_n16572 , new_n16545 , new_n16546 );
nor  g14224 ( new_n16573 , new_n16571 , new_n16572 );
nor  g14225 ( new_n16574 , new_n6696 , new_n8623 );
nor  g14226 ( new_n16575 , new_n8624 , new_n8643 );
nor  g14227 ( new_n16576 , new_n16574 , new_n16575 );
xnor g14228 ( new_n16577 , new_n16571 , new_n16572 );
nor  g14229 ( new_n16578 , new_n16576 , new_n16577 );
nor  g14230 ( new_n16579 , new_n16573 , new_n16578 );
nor  g14231 ( new_n16580 , new_n16569 , new_n16579 );
nor  g14232 ( new_n16581 , new_n16568 , new_n16580 );
xnor g14233 ( n4103 , new_n16565 , new_n16581 );
nor  g14234 ( new_n16583_1 , new_n12595 , new_n14513 );
xnor g14235 ( new_n16584_1 , new_n12595 , new_n14514 );
not  g14236 ( new_n16585 , new_n12518 );
nor  g14237 ( new_n16586 , new_n16585 , new_n14518 );
not  g14238 ( new_n16587 , new_n12523 );
nor  g14239 ( new_n16588 , new_n16587 , new_n14522 );
xnor g14240 ( new_n16589_1 , new_n12523 , new_n14522 );
and  g14241 ( new_n16590 , new_n12528 , new_n14526 );
xnor g14242 ( new_n16591 , new_n12528 , new_n14526 );
not  g14243 ( new_n16592 , new_n12533 );
nor  g14244 ( new_n16593 , new_n16592 , new_n14529 );
xnor g14245 ( new_n16594 , new_n12533 , new_n14529 );
and  g14246 ( new_n16595 , new_n12537 , new_n14445 );
nor  g14247 ( new_n16596_1 , new_n4251 , new_n12545_1 );
xnor g14248 ( new_n16597 , new_n14447 , new_n12545_1 );
nor  g14249 ( new_n16598 , new_n4258 , new_n12550 );
xnor g14250 ( new_n16599 , new_n4257 , new_n12550 );
nor  g14251 ( new_n16600 , new_n4277 , new_n12554 );
xnor g14252 ( new_n16601 , new_n4277 , new_n12553 );
not  g14253 ( new_n16602 , new_n4264 );
nor  g14254 ( new_n16603 , new_n16602 , new_n12565 );
or   g14255 ( new_n16604 , new_n4266_1 , new_n12563 );
xnor g14256 ( new_n16605 , new_n16602 , new_n12560 );
and  g14257 ( new_n16606 , new_n16604 , new_n16605 );
or   g14258 ( new_n16607 , new_n16603 , new_n16606 );
and  g14259 ( new_n16608_1 , new_n16601 , new_n16607 );
nor  g14260 ( new_n16609 , new_n16600 , new_n16608_1 );
and  g14261 ( new_n16610 , new_n16599 , new_n16609 );
nor  g14262 ( new_n16611 , new_n16598 , new_n16610 );
and  g14263 ( new_n16612 , new_n16597 , new_n16611 );
nor  g14264 ( new_n16613 , new_n16596_1 , new_n16612 );
xnor g14265 ( new_n16614 , new_n12537 , new_n14445 );
nor  g14266 ( new_n16615 , new_n16613 , new_n16614 );
or   g14267 ( new_n16616 , new_n16595 , new_n16615 );
and  g14268 ( new_n16617_1 , new_n16594 , new_n16616 );
nor  g14269 ( new_n16618 , new_n16593 , new_n16617_1 );
nor  g14270 ( new_n16619 , new_n16591 , new_n16618 );
or   g14271 ( new_n16620 , new_n16590 , new_n16619 );
and  g14272 ( new_n16621 , new_n16589_1 , new_n16620 );
or   g14273 ( new_n16622 , new_n16588 , new_n16621 );
xnor g14274 ( new_n16623 , new_n12518 , new_n14518 );
and  g14275 ( new_n16624 , new_n16622 , new_n16623 );
nor  g14276 ( new_n16625 , new_n16586 , new_n16624 );
and  g14277 ( new_n16626 , new_n16584_1 , new_n16625 );
nor  g14278 ( new_n16627 , new_n16583_1 , new_n16626 );
not  g14279 ( new_n16628 , new_n16627 );
nor  g14280 ( new_n16629 , new_n5872 , new_n13508 );
or   g14281 ( new_n16630_1 , n6456 , new_n5871 );
nor  g14282 ( new_n16631 , n4085 , new_n5917 );
xnor g14283 ( new_n16632 , new_n5875 , new_n5917 );
nor  g14284 ( new_n16633 , n26725 , new_n5923 );
xnor g14285 ( new_n16634 , n26725 , new_n5923 );
nor  g14286 ( new_n16635 , n11980 , new_n5928 );
xnor g14287 ( new_n16636 , new_n5880 , new_n5928 );
nor  g14288 ( new_n16637 , n3253 , new_n5933 );
xnor g14289 ( new_n16638 , new_n5883 , new_n5933 );
nor  g14290 ( new_n16639 , n7759 , new_n5938 );
xnor g14291 ( new_n16640_1 , new_n5886 , new_n5938 );
nor  g14292 ( new_n16641 , n12562 , new_n5943_1 );
nor  g14293 ( new_n16642 , n7949 , new_n5949 );
xnor g14294 ( new_n16643 , n7949 , new_n5950 );
nor  g14295 ( new_n16644 , n24374 , new_n5960 );
or   g14296 ( new_n16645 , new_n5895 , new_n3798 );
xnor g14297 ( new_n16646 , n24374 , new_n5961 );
and  g14298 ( new_n16647 , new_n16645 , new_n16646 );
or   g14299 ( new_n16648 , new_n16644 , new_n16647 );
and  g14300 ( new_n16649 , new_n16643 , new_n16648 );
or   g14301 ( new_n16650 , new_n16642 , new_n16649 );
xnor g14302 ( new_n16651 , new_n5889 , new_n5943_1 );
and  g14303 ( new_n16652 , new_n16650 , new_n16651 );
or   g14304 ( new_n16653 , new_n16641 , new_n16652 );
and  g14305 ( new_n16654 , new_n16640_1 , new_n16653 );
or   g14306 ( new_n16655 , new_n16639 , new_n16654 );
and  g14307 ( new_n16656_1 , new_n16638 , new_n16655 );
or   g14308 ( new_n16657 , new_n16637 , new_n16656_1 );
and  g14309 ( new_n16658 , new_n16636 , new_n16657 );
nor  g14310 ( new_n16659 , new_n16635 , new_n16658 );
nor  g14311 ( new_n16660 , new_n16634 , new_n16659 );
or   g14312 ( new_n16661 , new_n16633 , new_n16660 );
and  g14313 ( new_n16662 , new_n16632 , new_n16661 );
nor  g14314 ( new_n16663 , new_n16631 , new_n16662 );
and  g14315 ( new_n16664 , new_n16630_1 , new_n16663 );
or   g14316 ( new_n16665 , new_n13550 , new_n16664 );
nor  g14317 ( new_n16666 , new_n16629 , new_n16665 );
and  g14318 ( new_n16667 , new_n16628 , new_n16666 );
xor  g14319 ( new_n16668 , new_n16584_1 , new_n16625 );
nor  g14320 ( new_n16669 , new_n16666 , new_n16668 );
xnor g14321 ( new_n16670 , new_n16666 , new_n16668 );
xor  g14322 ( new_n16671 , new_n16622 , new_n16623 );
xnor g14323 ( new_n16672 , n6456 , new_n13508 );
xnor g14324 ( new_n16673 , new_n16663 , new_n16672 );
and  g14325 ( new_n16674_1 , new_n16671 , new_n16673 );
xnor g14326 ( new_n16675 , new_n16671 , new_n16673 );
xor  g14327 ( new_n16676 , new_n16632 , new_n16661 );
xor  g14328 ( new_n16677 , new_n16589_1 , new_n16620 );
and  g14329 ( new_n16678 , new_n16676 , new_n16677 );
xnor g14330 ( new_n16679 , new_n16676 , new_n16677 );
xnor g14331 ( new_n16680 , new_n16634 , new_n16659 );
xnor g14332 ( new_n16681 , new_n16591 , new_n16618 );
nor  g14333 ( new_n16682_1 , new_n16680 , new_n16681 );
xnor g14334 ( new_n16683 , new_n16680 , new_n16681 );
xor  g14335 ( new_n16684_1 , new_n16636 , new_n16657 );
xor  g14336 ( new_n16685 , new_n16594 , new_n16616 );
and  g14337 ( new_n16686 , new_n16684_1 , new_n16685 );
xnor g14338 ( new_n16687 , new_n16684_1 , new_n16685 );
xor  g14339 ( new_n16688_1 , new_n16638 , new_n16655 );
xnor g14340 ( new_n16689 , new_n16613 , new_n16614 );
not  g14341 ( new_n16690 , new_n16689 );
and  g14342 ( new_n16691 , new_n16688_1 , new_n16690 );
xnor g14343 ( new_n16692 , new_n16688_1 , new_n16690 );
xor  g14344 ( new_n16693 , new_n16640_1 , new_n16653 );
xnor g14345 ( new_n16694 , new_n16597 , new_n16611 );
not  g14346 ( new_n16695 , new_n16694 );
and  g14347 ( new_n16696 , new_n16693 , new_n16695 );
xnor g14348 ( new_n16697 , new_n16693 , new_n16695 );
xnor g14349 ( new_n16698 , new_n16599 , new_n16609 );
xor  g14350 ( new_n16699 , new_n16650 , new_n16651 );
and  g14351 ( new_n16700 , new_n16698 , new_n16699 );
not  g14352 ( new_n16701 , new_n16698 );
xnor g14353 ( new_n16702 , new_n16701 , new_n16699 );
xor  g14354 ( new_n16703 , new_n16643 , new_n16648 );
xor  g14355 ( new_n16704 , new_n16601 , new_n16607 );
nor  g14356 ( new_n16705 , new_n16703 , new_n16704 );
xor  g14357 ( new_n16706 , new_n16703 , new_n16704 );
nor  g14358 ( new_n16707 , new_n4266_1 , new_n12563 );
xnor g14359 ( new_n16708 , new_n16707 , new_n16605 );
not  g14360 ( new_n16709 , new_n16708 );
nor  g14361 ( new_n16710 , new_n16646 , new_n16709 );
xor  g14362 ( new_n16711 , new_n16645 , new_n16646 );
nor  g14363 ( new_n16712 , new_n16708 , new_n16711 );
xnor g14364 ( new_n16713 , n14575 , n20658 );
xnor g14365 ( new_n16714 , new_n4266_1 , new_n12562_1 );
not  g14366 ( new_n16715 , new_n16714 );
nor  g14367 ( new_n16716 , new_n16713 , new_n16715 );
nor  g14368 ( new_n16717 , new_n16712 , new_n16716 );
nor  g14369 ( new_n16718 , new_n16710 , new_n16717 );
and  g14370 ( new_n16719 , new_n16706 , new_n16718 );
nor  g14371 ( new_n16720 , new_n16705 , new_n16719 );
and  g14372 ( new_n16721 , new_n16702 , new_n16720 );
nor  g14373 ( new_n16722_1 , new_n16700 , new_n16721 );
nor  g14374 ( new_n16723 , new_n16697 , new_n16722_1 );
nor  g14375 ( new_n16724 , new_n16696 , new_n16723 );
nor  g14376 ( new_n16725 , new_n16692 , new_n16724 );
nor  g14377 ( new_n16726 , new_n16691 , new_n16725 );
nor  g14378 ( new_n16727 , new_n16687 , new_n16726 );
nor  g14379 ( new_n16728 , new_n16686 , new_n16727 );
nor  g14380 ( new_n16729 , new_n16683 , new_n16728 );
nor  g14381 ( new_n16730 , new_n16682_1 , new_n16729 );
nor  g14382 ( new_n16731 , new_n16679 , new_n16730 );
nor  g14383 ( new_n16732 , new_n16678 , new_n16731 );
nor  g14384 ( new_n16733_1 , new_n16675 , new_n16732 );
nor  g14385 ( new_n16734 , new_n16674_1 , new_n16733_1 );
nor  g14386 ( new_n16735 , new_n16670 , new_n16734 );
nor  g14387 ( new_n16736 , new_n16669 , new_n16735 );
nor  g14388 ( new_n16737 , new_n16667 , new_n16736 );
nor  g14389 ( new_n16738 , new_n16628 , new_n16666 );
nor  g14390 ( new_n16739 , new_n16735 , new_n16738 );
nor  g14391 ( n4123 , new_n16737 , new_n16739 );
xnor g14392 ( new_n16741 , new_n7870 , new_n13068 );
nor  g14393 ( new_n16742 , new_n7877 , new_n13071 );
xnor g14394 ( new_n16743_1 , new_n7876_1 , new_n13072 );
not  g14395 ( new_n16744 , new_n13076 );
nor  g14396 ( new_n16745 , new_n7899 , new_n16744 );
xnor g14397 ( new_n16746 , new_n7898 , new_n16744 );
and  g14398 ( new_n16747 , new_n7885 , new_n13086 );
nor  g14399 ( new_n16748 , new_n7887 , new_n9708 );
xnor g14400 ( new_n16749 , new_n7885 , new_n13085 );
and  g14401 ( new_n16750 , new_n16748 , new_n16749 );
nor  g14402 ( new_n16751 , new_n16747 , new_n16750 );
and  g14403 ( new_n16752 , new_n16746 , new_n16751 );
nor  g14404 ( new_n16753 , new_n16745 , new_n16752 );
nor  g14405 ( new_n16754 , new_n16743_1 , new_n16753 );
nor  g14406 ( new_n16755 , new_n16742 , new_n16754 );
xnor g14407 ( n4134 , new_n16741 , new_n16755 );
xnor g14408 ( n4146 , new_n9005 , new_n9055 );
xnor g14409 ( new_n16758 , new_n13958 , new_n15062 );
nor  g14410 ( new_n16759 , new_n13963 , new_n15068 );
xnor g14411 ( new_n16760 , new_n13963 , new_n15066 );
and  g14412 ( new_n16761 , new_n13150 , new_n13966 );
nor  g14413 ( new_n16762 , new_n13143 , new_n13969 );
xnor g14414 ( new_n16763 , new_n13149 , new_n13966 );
and  g14415 ( new_n16764 , new_n16762 , new_n16763 );
nor  g14416 ( new_n16765 , new_n16761 , new_n16764 );
and  g14417 ( new_n16766 , new_n16760 , new_n16765 );
nor  g14418 ( new_n16767 , new_n16759 , new_n16766 );
xnor g14419 ( n4150 , new_n16758 , new_n16767 );
xnor g14420 ( n4151 , new_n12341_1 , new_n12342 );
xnor g14421 ( n4152 , new_n12604 , new_n12663 );
xnor g14422 ( n4153 , new_n6104_1 , new_n6143 );
nor  g14423 ( new_n16772 , n10250 , new_n11842_1 );
and  g14424 ( new_n16773 , new_n8645 , new_n8680 );
nor  g14425 ( new_n16774 , new_n16772 , new_n16773 );
xnor g14426 ( new_n16775 , new_n12059 , new_n16774 );
not  g14427 ( new_n16776 , new_n16774 );
nor  g14428 ( new_n16777 , new_n12063 , new_n16776 );
nor  g14429 ( new_n16778 , new_n12064 , new_n16774 );
and  g14430 ( new_n16779 , new_n8681 , new_n12067 );
and  g14431 ( new_n16780 , new_n8854 , new_n8909_1 );
nor  g14432 ( new_n16781 , new_n16779 , new_n16780 );
nor  g14433 ( new_n16782 , new_n16778 , new_n16781 );
nor  g14434 ( new_n16783 , new_n16777 , new_n16782 );
xnor g14435 ( n4165 , new_n16775 , new_n16783 );
xnor g14436 ( n4172 , new_n11382 , new_n11411 );
xnor g14437 ( n4173 , new_n4745_1 , new_n11249 );
xnor g14438 ( n4176 , new_n6559 , new_n6579 );
xnor g14439 ( n4186 , new_n9039 , new_n9040 );
xnor g14440 ( n4204 , new_n16335 , new_n16357 );
nor  g14441 ( new_n16790 , new_n5500 , new_n11296 );
xnor g14442 ( new_n16791 , new_n5500 , new_n11296 );
nor  g14443 ( new_n16792 , new_n5503 , new_n6789 );
nor  g14444 ( new_n16793 , new_n6790_1 , new_n6832 );
nor  g14445 ( new_n16794 , new_n16792 , new_n16793 );
nor  g14446 ( new_n16795 , new_n16791 , new_n16794 );
nor  g14447 ( new_n16796 , new_n16790 , new_n16795 );
nor  g14448 ( new_n16797 , new_n11792 , new_n16796 );
not  g14449 ( new_n16798_1 , new_n15725 );
nor  g14450 ( new_n16799 , n3366 , new_n16798_1 );
not  g14451 ( new_n16800 , new_n16799 );
nor  g14452 ( new_n16801 , n19652 , new_n16800 );
xnor g14453 ( new_n16802 , n3984 , new_n16801 );
and  g14454 ( new_n16803 , new_n11326_1 , new_n16802 );
xnor g14455 ( new_n16804 , n17037 , new_n16802 );
xnor g14456 ( new_n16805 , n19652 , new_n16800 );
and  g14457 ( new_n16806 , n5386 , new_n16805 );
not  g14458 ( new_n16807 , new_n15726 );
nor  g14459 ( new_n16808 , n26191 , new_n16807 );
and  g14460 ( new_n16809 , new_n15727 , new_n15757 );
nor  g14461 ( new_n16810 , new_n16808 , new_n16809 );
xor  g14462 ( new_n16811 , n5386 , new_n16805 );
and  g14463 ( new_n16812_1 , new_n16810 , new_n16811 );
nor  g14464 ( new_n16813 , new_n16806 , new_n16812_1 );
and  g14465 ( new_n16814 , new_n16804 , new_n16813 );
nor  g14466 ( new_n16815 , new_n16803 , new_n16814 );
not  g14467 ( new_n16816 , new_n16801 );
nor  g14468 ( new_n16817 , n3984 , new_n16816 );
xnor g14469 ( new_n16818_1 , n4514 , new_n16817 );
xnor g14470 ( new_n16819 , n7569 , new_n16818_1 );
xnor g14471 ( new_n16820 , new_n16815 , new_n16819 );
nor  g14472 ( new_n16821 , new_n14303 , new_n16820 );
xnor g14473 ( new_n16822 , new_n14303 , new_n16820 );
xor  g14474 ( new_n16823 , new_n16804 , new_n16813 );
nor  g14475 ( new_n16824_1 , new_n14165 , new_n16823 );
xnor g14476 ( new_n16825 , n25751 , new_n16823 );
xor  g14477 ( new_n16826 , new_n16810 , new_n16811 );
nor  g14478 ( new_n16827 , n26053 , new_n16826 );
xnor g14479 ( new_n16828 , new_n14168 , new_n16826 );
and  g14480 ( new_n16829 , new_n14171 , new_n15758 );
and  g14481 ( new_n16830 , new_n15759 , new_n15787 );
or   g14482 ( new_n16831 , new_n16829 , new_n16830 );
and  g14483 ( new_n16832 , new_n16828 , new_n16831 );
nor  g14484 ( new_n16833 , new_n16827 , new_n16832 );
and  g14485 ( new_n16834_1 , new_n16825 , new_n16833 );
nor  g14486 ( new_n16835 , new_n16824_1 , new_n16834_1 );
nor  g14487 ( new_n16836 , new_n16822 , new_n16835 );
nor  g14488 ( new_n16837_1 , new_n16821 , new_n16836 );
and  g14489 ( new_n16838 , new_n11273_1 , new_n16817 );
nor  g14490 ( new_n16839 , new_n11325_1 , new_n16818_1 );
nor  g14491 ( new_n16840 , new_n16815 , new_n16839 );
and  g14492 ( new_n16841_1 , new_n16838 , new_n16840 );
and  g14493 ( new_n16842 , new_n16837_1 , new_n16841_1 );
and  g14494 ( new_n16843 , new_n11325_1 , new_n16818_1 );
xor  g14495 ( new_n16844 , new_n16838 , new_n16840 );
nor  g14496 ( new_n16845 , new_n16843 , new_n16844 );
not  g14497 ( new_n16846 , new_n16845 );
or   g14498 ( new_n16847 , new_n16837_1 , new_n16846 );
nor  g14499 ( new_n16848 , new_n16841_1 , new_n16847 );
nor  g14500 ( new_n16849 , new_n16842 , new_n16848 );
or   g14501 ( new_n16850 , new_n16797 , new_n16849 );
xnor g14502 ( new_n16851 , new_n16837_1 , new_n16845 );
xnor g14503 ( new_n16852 , new_n11323 , new_n16796 );
not  g14504 ( new_n16853 , new_n16852 );
and  g14505 ( new_n16854 , new_n16851 , new_n16853 );
xnor g14506 ( new_n16855 , new_n16851 , new_n16853 );
xnor g14507 ( new_n16856 , new_n16822 , new_n16835 );
xnor g14508 ( new_n16857 , new_n16791 , new_n16794 );
not  g14509 ( new_n16858 , new_n16857 );
nor  g14510 ( new_n16859 , new_n16856 , new_n16858 );
xnor g14511 ( new_n16860 , new_n16856 , new_n16858 );
not  g14512 ( new_n16861 , new_n6833 );
xnor g14513 ( new_n16862 , new_n16825 , new_n16833 );
nor  g14514 ( new_n16863 , new_n16861 , new_n16862 );
xnor g14515 ( new_n16864 , new_n16861 , new_n16862 );
xor  g14516 ( new_n16865 , new_n16828 , new_n16831 );
nor  g14517 ( new_n16866 , new_n6913 , new_n16865 );
nor  g14518 ( new_n16867 , new_n6918 , new_n15788 );
nor  g14519 ( new_n16868 , new_n15789 , new_n15818 );
nor  g14520 ( new_n16869 , new_n16867 , new_n16868 );
xnor g14521 ( new_n16870 , new_n6913 , new_n16865 );
nor  g14522 ( new_n16871 , new_n16869 , new_n16870 );
nor  g14523 ( new_n16872 , new_n16866 , new_n16871 );
nor  g14524 ( new_n16873 , new_n16864 , new_n16872 );
nor  g14525 ( new_n16874 , new_n16863 , new_n16873 );
nor  g14526 ( new_n16875 , new_n16860 , new_n16874 );
nor  g14527 ( new_n16876 , new_n16859 , new_n16875 );
nor  g14528 ( new_n16877 , new_n16855 , new_n16876 );
nor  g14529 ( new_n16878 , new_n16854 , new_n16877 );
and  g14530 ( new_n16879 , new_n16850 , new_n16878 );
and  g14531 ( new_n16880 , new_n16797 , new_n16849 );
or   g14532 ( new_n16881 , new_n16842 , new_n16880 );
nor  g14533 ( n4205 , new_n16879 , new_n16881 );
not  g14534 ( new_n16883 , new_n12997 );
nor  g14535 ( new_n16884 , n22198 , new_n16883 );
not  g14536 ( new_n16885_1 , new_n16884 );
nor  g14537 ( new_n16886 , n24327 , new_n16885_1 );
xnor g14538 ( new_n16887 , n2659 , new_n16886 );
xnor g14539 ( new_n16888 , n18444 , new_n16887 );
xnor g14540 ( new_n16889 , n24327 , new_n16884 );
nor  g14541 ( new_n16890 , n24638 , new_n16889 );
xnor g14542 ( new_n16891 , n24638 , new_n16889 );
nor  g14543 ( new_n16892 , n21674 , new_n12998 );
nor  g14544 ( new_n16893 , new_n12999 , new_n13020 );
nor  g14545 ( new_n16894 , new_n16892 , new_n16893 );
nor  g14546 ( new_n16895 , new_n16891 , new_n16894 );
nor  g14547 ( new_n16896 , new_n16890 , new_n16895 );
xor  g14548 ( new_n16897 , new_n16888 , new_n16896 );
xnor g14549 ( new_n16898 , new_n7715 , new_n16897 );
xnor g14550 ( new_n16899 , new_n16891 , new_n16894 );
and  g14551 ( new_n16900 , new_n7718 , new_n16899 );
xor  g14552 ( new_n16901 , new_n7718 , new_n16899 );
nor  g14553 ( new_n16902 , new_n7722 , new_n13021 );
nor  g14554 ( new_n16903 , new_n13022 , new_n13043_1 );
nor  g14555 ( new_n16904 , new_n16902 , new_n16903 );
and  g14556 ( new_n16905_1 , new_n16901 , new_n16904 );
nor  g14557 ( new_n16906 , new_n16900 , new_n16905_1 );
xnor g14558 ( new_n16907 , new_n16898 , new_n16906 );
xnor g14559 ( new_n16908 , n5400 , n21997 );
nor  g14560 ( new_n16909 , new_n8284 , n25119 );
xnor g14561 ( new_n16910 , n23923 , n25119 );
nor  g14562 ( new_n16911_1 , new_n8353 , n1163 );
and  g14563 ( new_n16912 , new_n13045 , new_n13064 );
or   g14564 ( new_n16913 , new_n16911_1 , new_n16912 );
and  g14565 ( new_n16914 , new_n16910 , new_n16913 );
or   g14566 ( new_n16915 , new_n16909 , new_n16914 );
xor  g14567 ( new_n16916 , new_n16908 , new_n16915 );
xnor g14568 ( new_n16917 , new_n16907 , new_n16916 );
xor  g14569 ( new_n16918 , new_n16910 , new_n16913 );
xnor g14570 ( new_n16919 , new_n16901 , new_n16904 );
not  g14571 ( new_n16920 , new_n16919 );
and  g14572 ( new_n16921 , new_n16918 , new_n16920 );
xnor g14573 ( new_n16922 , new_n16918 , new_n16919 );
nor  g14574 ( new_n16923 , new_n13044_1 , new_n13065 );
nor  g14575 ( new_n16924 , new_n13066 , new_n13095 );
nor  g14576 ( new_n16925 , new_n16923 , new_n16924 );
and  g14577 ( new_n16926 , new_n16922 , new_n16925 );
or   g14578 ( new_n16927 , new_n16921 , new_n16926 );
xor  g14579 ( n4215 , new_n16917 , new_n16927 );
and  g14580 ( new_n16929 , new_n5985 , new_n14005 );
xnor g14581 ( new_n16930 , n3582 , new_n16929 );
xnor g14582 ( new_n16931 , new_n4907 , new_n16930 );
and  g14583 ( new_n16932 , n2858 , new_n14006 );
or   g14584 ( new_n16933 , n2858 , new_n14006 );
and  g14585 ( new_n16934 , new_n16933 , new_n14031 );
nor  g14586 ( new_n16935 , new_n16932 , new_n16934 );
xnor g14587 ( new_n16936 , new_n16931 , new_n16935 );
not  g14588 ( new_n16937 , new_n9610 );
nor  g14589 ( new_n16938 , n27089 , new_n16937 );
xnor g14590 ( new_n16939 , n21839 , new_n16938 );
not  g14591 ( new_n16940 , new_n16939 );
xnor g14592 ( new_n16941 , n22626 , new_n16940 );
nor  g14593 ( new_n16942 , n14440 , new_n9611 );
xnor g14594 ( new_n16943 , new_n7482 , new_n9611 );
not  g14595 ( new_n16944 , new_n16943 );
nor  g14596 ( new_n16945 , n1654 , new_n9613 );
nor  g14597 ( new_n16946 , new_n15488 , new_n15491 );
nor  g14598 ( new_n16947 , new_n16945 , new_n16946 );
nor  g14599 ( new_n16948 , new_n16944 , new_n16947 );
or   g14600 ( new_n16949 , new_n16942 , new_n16948 );
xnor g14601 ( new_n16950 , new_n16941 , new_n16949 );
xnor g14602 ( new_n16951_1 , new_n16936 , new_n16950 );
xnor g14603 ( new_n16952 , new_n16943 , new_n16947 );
nor  g14604 ( new_n16953 , new_n14032 , new_n16952 );
not  g14605 ( new_n16954_1 , new_n14035 );
nor  g14606 ( new_n16955 , new_n16954_1 , new_n15492 );
xnor g14607 ( new_n16956 , new_n16954_1 , new_n15492 );
nor  g14608 ( new_n16957 , new_n10541 , new_n14038 );
xnor g14609 ( new_n16958 , new_n10541 , new_n14038 );
nor  g14610 ( new_n16959 , new_n10543 , new_n14041 );
xnor g14611 ( new_n16960 , new_n10546 , new_n14043 );
nor  g14612 ( new_n16961 , new_n10554 , new_n14048 );
xnor g14613 ( new_n16962 , new_n10554 , new_n14048 );
and  g14614 ( new_n16963 , new_n9409 , new_n9423_1 );
nor  g14615 ( new_n16964 , new_n9424 , new_n9440 );
nor  g14616 ( new_n16965 , new_n16963 , new_n16964 );
nor  g14617 ( new_n16966 , new_n16962 , new_n16965 );
or   g14618 ( new_n16967 , new_n16961 , new_n16966 );
nor  g14619 ( new_n16968_1 , new_n16960 , new_n16967 );
nor  g14620 ( new_n16969 , new_n16959 , new_n16968_1 );
nor  g14621 ( new_n16970 , new_n16958 , new_n16969 );
nor  g14622 ( new_n16971_1 , new_n16957 , new_n16970 );
nor  g14623 ( new_n16972 , new_n16956 , new_n16971_1 );
nor  g14624 ( new_n16973 , new_n16955 , new_n16972 );
not  g14625 ( new_n16974 , new_n16952 );
xnor g14626 ( new_n16975 , new_n14032 , new_n16974 );
and  g14627 ( new_n16976 , new_n16973 , new_n16975 );
nor  g14628 ( new_n16977 , new_n16953 , new_n16976 );
xnor g14629 ( new_n16978 , new_n16951_1 , new_n16977 );
not  g14630 ( new_n16979 , new_n16978 );
not  g14631 ( new_n16980 , new_n14749 );
nor  g14632 ( new_n16981 , n10611 , new_n16980 );
not  g14633 ( new_n16982 , new_n16981 );
nor  g14634 ( new_n16983 , n3164 , new_n16982 );
not  g14635 ( new_n16984 , new_n16983 );
nor  g14636 ( new_n16985 , n11356 , new_n16984 );
not  g14637 ( new_n16986 , new_n16985 );
nor  g14638 ( new_n16987 , n14345 , new_n16986 );
not  g14639 ( new_n16988_1 , new_n16987 );
nor  g14640 ( new_n16989_1 , n6381 , new_n16988_1 );
not  g14641 ( new_n16990 , new_n16989_1 );
nor  g14642 ( new_n16991 , n10577 , new_n16990 );
xnor g14643 ( new_n16992 , n23166 , new_n16991 );
xnor g14644 ( new_n16993 , new_n7772 , new_n16992 );
xnor g14645 ( new_n16994_1 , n10577 , new_n16989_1 );
nor  g14646 ( new_n16995 , n26408 , new_n16994_1 );
xnor g14647 ( new_n16996 , n26408 , new_n16994_1 );
xnor g14648 ( new_n16997 , n6381 , new_n16987 );
nor  g14649 ( new_n16998 , n18227 , new_n16997 );
xnor g14650 ( new_n16999 , new_n4804_1 , new_n16997 );
xnor g14651 ( new_n17000 , n14345 , new_n16985 );
nor  g14652 ( new_n17001 , n7377 , new_n17000 );
xnor g14653 ( new_n17002 , new_n4807 , new_n17000 );
xnor g14654 ( new_n17003 , n11356 , new_n16983 );
nor  g14655 ( new_n17004 , n11630 , new_n17003 );
xnor g14656 ( new_n17005 , n3164 , new_n16981 );
nor  g14657 ( new_n17006_1 , n13453 , new_n17005 );
xnor g14658 ( new_n17007 , new_n12754 , new_n17005 );
and  g14659 ( new_n17008 , n7421 , new_n14750 );
and  g14660 ( new_n17009 , new_n14751 , new_n14763_1 );
nor  g14661 ( new_n17010 , new_n17008 , new_n17009 );
and  g14662 ( new_n17011 , new_n17007 , new_n17010 );
or   g14663 ( new_n17012 , new_n17006_1 , new_n17011 );
not  g14664 ( new_n17013 , n11630 );
xnor g14665 ( new_n17014 , new_n17013 , new_n17003 );
and  g14666 ( new_n17015 , new_n17012 , new_n17014 );
or   g14667 ( new_n17016 , new_n17004 , new_n17015 );
and  g14668 ( new_n17017 , new_n17002 , new_n17016 );
or   g14669 ( new_n17018 , new_n17001 , new_n17017 );
and  g14670 ( new_n17019 , new_n16999 , new_n17018 );
nor  g14671 ( new_n17020 , new_n16998 , new_n17019 );
nor  g14672 ( new_n17021 , new_n16996 , new_n17020 );
nor  g14673 ( new_n17022 , new_n16995 , new_n17021 );
xnor g14674 ( new_n17023 , new_n16993 , new_n17022 );
not  g14675 ( new_n17024 , new_n17023 );
xnor g14676 ( new_n17025 , new_n16979 , new_n17024 );
xnor g14677 ( new_n17026 , new_n16996 , new_n17020 );
xor  g14678 ( new_n17027 , new_n16973 , new_n16975 );
nor  g14679 ( new_n17028 , new_n17026 , new_n17027 );
xnor g14680 ( new_n17029 , new_n17026 , new_n17027 );
nor  g14681 ( new_n17030 , new_n17001 , new_n17017 );
xnor g14682 ( new_n17031 , new_n16999 , new_n17030 );
not  g14683 ( new_n17032 , new_n17031 );
xor  g14684 ( new_n17033 , new_n16956 , new_n16971_1 );
not  g14685 ( new_n17034 , new_n17033 );
nor  g14686 ( new_n17035_1 , new_n17032 , new_n17034 );
xnor g14687 ( new_n17036 , new_n17032 , new_n17034 );
nor  g14688 ( new_n17037_1 , new_n17004 , new_n17015 );
xnor g14689 ( new_n17038 , new_n17002 , new_n17037_1 );
not  g14690 ( new_n17039 , new_n17038 );
xor  g14691 ( new_n17040 , new_n16958 , new_n16969 );
not  g14692 ( new_n17041 , new_n17040 );
nor  g14693 ( new_n17042 , new_n17039 , new_n17041 );
xnor g14694 ( new_n17043 , new_n17039 , new_n17041 );
nor  g14695 ( new_n17044 , new_n16961 , new_n16966 );
xnor g14696 ( new_n17045 , new_n16960 , new_n17044 );
not  g14697 ( new_n17046 , new_n17045 );
xor  g14698 ( new_n17047 , new_n17012 , new_n17014 );
not  g14699 ( new_n17048 , new_n17047 );
nor  g14700 ( new_n17049 , new_n17046 , new_n17048 );
xnor g14701 ( new_n17050 , new_n17046 , new_n17048 );
xnor g14702 ( new_n17051 , new_n17007 , new_n17010 );
xor  g14703 ( new_n17052 , new_n16962 , new_n16965 );
nor  g14704 ( new_n17053 , new_n17051 , new_n17052 );
not  g14705 ( new_n17054 , new_n17051 );
not  g14706 ( new_n17055 , new_n17052 );
xnor g14707 ( new_n17056 , new_n17054 , new_n17055 );
nor  g14708 ( new_n17057 , new_n9441 , new_n14764 );
xnor g14709 ( new_n17058 , new_n9441 , new_n14764 );
not  g14710 ( new_n17059 , new_n17058 );
nor  g14711 ( new_n17060 , new_n9455 , new_n14766 );
xnor g14712 ( new_n17061 , new_n9455 , new_n14766 );
nor  g14713 ( new_n17062 , new_n9467 , new_n14770 );
nor  g14714 ( new_n17063 , new_n9462 , new_n14772_1 );
xnor g14715 ( new_n17064 , new_n9468 , new_n14770 );
and  g14716 ( new_n17065 , new_n17063 , new_n17064 );
nor  g14717 ( new_n17066 , new_n17062 , new_n17065 );
nor  g14718 ( new_n17067 , new_n17061 , new_n17066 );
nor  g14719 ( new_n17068_1 , new_n17060 , new_n17067 );
and  g14720 ( new_n17069_1 , new_n17059 , new_n17068_1 );
nor  g14721 ( new_n17070_1 , new_n17057 , new_n17069_1 );
nor  g14722 ( new_n17071 , new_n17056 , new_n17070_1 );
nor  g14723 ( new_n17072 , new_n17053 , new_n17071 );
nor  g14724 ( new_n17073 , new_n17050 , new_n17072 );
nor  g14725 ( new_n17074 , new_n17049 , new_n17073 );
nor  g14726 ( new_n17075_1 , new_n17043 , new_n17074 );
nor  g14727 ( new_n17076 , new_n17042 , new_n17075_1 );
nor  g14728 ( new_n17077_1 , new_n17036 , new_n17076 );
nor  g14729 ( new_n17078 , new_n17035_1 , new_n17077_1 );
nor  g14730 ( new_n17079 , new_n17029 , new_n17078 );
or   g14731 ( new_n17080 , new_n17028 , new_n17079 );
xor  g14732 ( n4221 , new_n17025 , new_n17080 );
xnor g14733 ( new_n17082 , new_n4804_1 , new_n10450 );
nor  g14734 ( new_n17083 , new_n4807 , new_n10454 );
xnor g14735 ( new_n17084_1 , new_n4807 , new_n10456 );
nor  g14736 ( new_n17085 , new_n17013 , new_n10471 );
nor  g14737 ( new_n17086 , new_n12754 , new_n10462 );
or   g14738 ( new_n17087 , new_n12756_1 , new_n12757 );
and  g14739 ( new_n17088 , new_n12755 , new_n17087 );
or   g14740 ( new_n17089 , new_n17086 , new_n17088 );
xnor g14741 ( new_n17090_1 , n11630 , new_n10471 );
and  g14742 ( new_n17091 , new_n17089 , new_n17090_1 );
or   g14743 ( new_n17092 , new_n17085 , new_n17091 );
and  g14744 ( new_n17093 , new_n17084_1 , new_n17092 );
nor  g14745 ( new_n17094 , new_n17083 , new_n17093 );
xnor g14746 ( new_n17095_1 , new_n17082 , new_n17094 );
not  g14747 ( new_n17096 , new_n17095_1 );
xnor g14748 ( new_n17097 , new_n15885_1 , new_n17096 );
nor  g14749 ( new_n17098 , new_n17085 , new_n17091 );
xnor g14750 ( new_n17099 , new_n17084_1 , new_n17098 );
not  g14751 ( new_n17100 , new_n17099 );
nor  g14752 ( new_n17101 , new_n8499 , new_n17100 );
xnor g14753 ( new_n17102 , new_n8500 , new_n17099 );
nor  g14754 ( new_n17103 , new_n17086 , new_n17088 );
xnor g14755 ( new_n17104_1 , new_n17103 , new_n17090_1 );
and  g14756 ( new_n17105 , new_n8531 , new_n17104_1 );
xnor g14757 ( new_n17106_1 , new_n8531 , new_n17104_1 );
not  g14758 ( new_n17107 , new_n12759 );
nor  g14759 ( new_n17108 , new_n8537 , new_n17107 );
xnor g14760 ( new_n17109 , new_n15895 , new_n12759 );
nor  g14761 ( new_n17110 , new_n6623 , new_n8542 );
xnor g14762 ( new_n17111 , new_n6623 , new_n8542 );
nor  g14763 ( new_n17112 , new_n6654 , new_n8548 );
xnor g14764 ( new_n17113 , new_n6654 , new_n8548 );
nor  g14765 ( new_n17114 , new_n6660 , new_n8553 );
nor  g14766 ( new_n17115 , new_n6665 , new_n8556 );
xnor g14767 ( new_n17116 , new_n6668 , new_n8553 );
and  g14768 ( new_n17117 , new_n17115 , new_n17116 );
nor  g14769 ( new_n17118 , new_n17114 , new_n17117 );
nor  g14770 ( new_n17119_1 , new_n17113 , new_n17118 );
nor  g14771 ( new_n17120 , new_n17112 , new_n17119_1 );
nor  g14772 ( new_n17121 , new_n17111 , new_n17120 );
nor  g14773 ( new_n17122 , new_n17110 , new_n17121 );
nor  g14774 ( new_n17123 , new_n17109 , new_n17122 );
nor  g14775 ( new_n17124 , new_n17108 , new_n17123 );
nor  g14776 ( new_n17125 , new_n17106_1 , new_n17124 );
nor  g14777 ( new_n17126 , new_n17105 , new_n17125 );
nor  g14778 ( new_n17127 , new_n17102 , new_n17126 );
nor  g14779 ( new_n17128 , new_n17101 , new_n17127 );
xnor g14780 ( n4224 , new_n17097 , new_n17128 );
xor  g14781 ( n4231 , new_n10594 , new_n10595_1 );
xnor g14782 ( new_n17131 , n9934 , new_n13879 );
nor  g14783 ( new_n17132 , n18496 , new_n13881 );
or   g14784 ( new_n17133 , new_n16455 , new_n16461 );
and  g14785 ( new_n17134 , new_n16454 , new_n17133 );
nor  g14786 ( new_n17135 , new_n17132 , new_n17134 );
xnor g14787 ( new_n17136 , new_n17131 , new_n17135 );
not  g14788 ( new_n17137 , new_n17136 );
xnor g14789 ( new_n17138_1 , new_n4798 , new_n17137 );
nor  g14790 ( new_n17139 , new_n4801 , new_n16463 );
and  g14791 ( new_n17140 , new_n16465 , new_n16475 );
or   g14792 ( new_n17141 , new_n17139 , new_n17140 );
xor  g14793 ( new_n17142 , new_n17138_1 , new_n17141 );
xnor g14794 ( new_n17143 , new_n11741_1 , new_n17142 );
nor  g14795 ( new_n17144 , new_n11745 , new_n16476_1 );
nor  g14796 ( new_n17145 , new_n16477 , new_n16485 );
nor  g14797 ( new_n17146 , new_n17144 , new_n17145 );
xnor g14798 ( n4266 , new_n17143 , new_n17146 );
xnor g14799 ( n4340 , new_n6930 , new_n6956 );
xnor g14800 ( new_n17149 , new_n5953 , new_n16088 );
xnor g14801 ( new_n17150 , new_n12853 , new_n17149 );
nor  g14802 ( new_n17151 , new_n12869 , new_n16089 );
nor  g14803 ( new_n17152 , new_n16086 , new_n16090 );
nor  g14804 ( new_n17153 , new_n17151 , new_n17152 );
xor  g14805 ( new_n17154 , new_n17150 , new_n17153 );
xnor g14806 ( new_n17155 , new_n4999 , new_n17154 );
and  g14807 ( new_n17156 , new_n16085 , new_n16091 );
or   g14808 ( new_n17157 , new_n16084 , new_n17156 );
xor  g14809 ( n4374 , new_n17155 , new_n17157 );
xnor g14810 ( n4401 , new_n11034 , new_n11085 );
xor  g14811 ( n4424 , new_n12803 , new_n12804 );
not  g14812 ( new_n17161 , n1881 );
nor  g14813 ( new_n17162 , new_n17161 , new_n10685 );
xnor g14814 ( new_n17163_1 , n1881 , new_n10685 );
nor  g14815 ( new_n17164 , n5834 , new_n10677 );
xnor g14816 ( new_n17165 , n5834 , new_n10676 );
and  g14817 ( new_n17166 , n13851 , new_n10668 );
xnor g14818 ( new_n17167 , n13851 , new_n10667 );
and  g14819 ( new_n17168_1 , n24937 , new_n10659 );
or   g14820 ( new_n17169 , new_n15978 , new_n15984 );
and  g14821 ( new_n17170 , new_n15977 , new_n17169 );
or   g14822 ( new_n17171 , new_n17168_1 , new_n17170 );
and  g14823 ( new_n17172 , new_n17167 , new_n17171 );
nor  g14824 ( new_n17173 , new_n17166 , new_n17172 );
and  g14825 ( new_n17174 , new_n17165 , new_n17173 );
nor  g14826 ( new_n17175 , new_n17164 , new_n17174 );
and  g14827 ( new_n17176 , new_n17163_1 , new_n17175 );
nor  g14828 ( new_n17177 , new_n17162 , new_n17176 );
nor  g14829 ( new_n17178 , n4306 , n8827 );
not  g14830 ( new_n17179 , new_n10680 );
nor  g14831 ( new_n17180 , new_n17179 , new_n10684 );
nor  g14832 ( new_n17181 , new_n17178 , new_n17180 );
xnor g14833 ( new_n17182 , new_n17177 , new_n17181 );
not  g14834 ( new_n17183 , new_n17182 );
xnor g14835 ( new_n17184 , new_n9914 , new_n17183 );
xnor g14836 ( new_n17185 , new_n17163_1 , new_n17175 );
nor  g14837 ( new_n17186 , new_n9918 , new_n17185 );
xnor g14838 ( new_n17187 , new_n9918 , new_n17185 );
xor  g14839 ( new_n17188 , new_n17165 , new_n17173 );
nor  g14840 ( new_n17189 , new_n9923 , new_n17188 );
nor  g14841 ( new_n17190 , new_n17168_1 , new_n17170 );
xnor g14842 ( new_n17191 , new_n17167 , new_n17190 );
nor  g14843 ( new_n17192 , new_n9929 , new_n17191 );
not  g14844 ( new_n17193 , new_n17191 );
xnor g14845 ( new_n17194 , new_n9929 , new_n17193 );
nor  g14846 ( new_n17195 , new_n9934_1 , new_n15986_1 );
and  g14847 ( new_n17196 , new_n15988 , new_n15998 );
or   g14848 ( new_n17197 , new_n17195 , new_n17196 );
and  g14849 ( new_n17198 , new_n17194 , new_n17197 );
nor  g14850 ( new_n17199 , new_n17192 , new_n17198 );
xnor g14851 ( new_n17200 , new_n9924 , new_n17188 );
and  g14852 ( new_n17201 , new_n17199 , new_n17200 );
nor  g14853 ( new_n17202_1 , new_n17189 , new_n17201 );
nor  g14854 ( new_n17203 , new_n17187 , new_n17202_1 );
nor  g14855 ( new_n17204 , new_n17186 , new_n17203 );
xnor g14856 ( n4432 , new_n17184 , new_n17204 );
xnor g14857 ( n4441 , new_n14475_1 , new_n14476 );
nor  g14858 ( new_n17207 , n23065 , n27120 );
not  g14859 ( new_n17208 , new_n17207 );
nor  g14860 ( new_n17209 , n24786 , new_n17208 );
not  g14861 ( new_n17210 , new_n17209 );
nor  g14862 ( new_n17211 , n25370 , new_n17210 );
not  g14863 ( new_n17212 , new_n17211 );
nor  g14864 ( new_n17213 , n19472 , new_n17212 );
not  g14865 ( new_n17214 , new_n17213 );
nor  g14866 ( new_n17215 , n19042 , new_n17214 );
not  g14867 ( new_n17216 , new_n17215 );
nor  g14868 ( new_n17217 , n1293 , new_n17216 );
xnor g14869 ( new_n17218 , n13775 , new_n17217 );
xnor g14870 ( new_n17219_1 , new_n16533 , new_n17218 );
xnor g14871 ( new_n17220 , n1293 , new_n17215 );
nor  g14872 ( new_n17221 , new_n16537 , new_n17220 );
xnor g14873 ( new_n17222 , new_n16537 , new_n17220 );
not  g14874 ( new_n17223 , new_n16541 );
xnor g14875 ( new_n17224 , n19042 , new_n17213 );
nor  g14876 ( new_n17225 , new_n17223 , new_n17224 );
xnor g14877 ( new_n17226 , n19472 , new_n17211 );
nor  g14878 ( new_n17227 , new_n8600 , new_n17226 );
xnor g14879 ( new_n17228 , new_n8599 , new_n17226 );
xnor g14880 ( new_n17229 , n25370 , new_n17209 );
and  g14881 ( new_n17230 , new_n8603 , new_n17229 );
xnor g14882 ( new_n17231 , new_n8602 , new_n17229 );
xnor g14883 ( new_n17232_1 , n24786 , new_n17207 );
nor  g14884 ( new_n17233 , new_n8608_1 , new_n17232_1 );
xnor g14885 ( new_n17234 , new_n8608_1 , new_n17232_1 );
xnor g14886 ( new_n17235 , new_n4109 , n27120 );
nor  g14887 ( new_n17236_1 , new_n8612 , new_n17235 );
nor  g14888 ( new_n17237 , new_n8614_1 , new_n17236_1 );
nor  g14889 ( new_n17238 , new_n17234 , new_n17237 );
nor  g14890 ( new_n17239 , new_n17233 , new_n17238 );
and  g14891 ( new_n17240 , new_n17231 , new_n17239 );
nor  g14892 ( new_n17241 , new_n17230 , new_n17240 );
and  g14893 ( new_n17242 , new_n17228 , new_n17241 );
nor  g14894 ( new_n17243_1 , new_n17227 , new_n17242 );
xnor g14895 ( new_n17244 , new_n17223 , new_n17224 );
nor  g14896 ( new_n17245 , new_n17243_1 , new_n17244 );
nor  g14897 ( new_n17246 , new_n17225 , new_n17245 );
nor  g14898 ( new_n17247 , new_n17222 , new_n17246 );
nor  g14899 ( new_n17248 , new_n17221 , new_n17247 );
xor  g14900 ( new_n17249 , new_n17219_1 , new_n17248 );
not  g14901 ( new_n17250_1 , new_n11917 );
nor  g14902 ( new_n17251_1 , n26318 , new_n17250_1 );
xnor g14903 ( new_n17252 , n3710 , new_n17251_1 );
xnor g14904 ( new_n17253 , new_n5340 , new_n17252 );
nor  g14905 ( new_n17254 , new_n5348 , new_n11918 );
nor  g14906 ( new_n17255 , new_n11919 , new_n11945 );
nor  g14907 ( new_n17256 , new_n17254 , new_n17255 );
xor  g14908 ( new_n17257 , new_n17253 , new_n17256 );
xnor g14909 ( new_n17258 , new_n17249 , new_n17257 );
xnor g14910 ( new_n17259 , new_n17222 , new_n17246 );
nor  g14911 ( new_n17260 , new_n11946 , new_n17259 );
xnor g14912 ( new_n17261 , new_n11946 , new_n17259 );
xnor g14913 ( new_n17262 , new_n17243_1 , new_n17244 );
nor  g14914 ( new_n17263_1 , new_n11980_1 , new_n17262 );
xnor g14915 ( new_n17264 , new_n11981 , new_n17262 );
not  g14916 ( new_n17265 , new_n11984 );
xor  g14917 ( new_n17266 , new_n17228 , new_n17241 );
nor  g14918 ( new_n17267 , new_n17265 , new_n17266 );
xor  g14919 ( new_n17268 , new_n17231 , new_n17239 );
nor  g14920 ( new_n17269 , new_n11988 , new_n17268 );
xnor g14921 ( new_n17270 , new_n11988 , new_n17268 );
xnor g14922 ( new_n17271 , new_n17234 , new_n17237 );
and  g14923 ( new_n17272 , new_n11992 , new_n17271 );
nor  g14924 ( new_n17273 , new_n11992 , new_n17271 );
xor  g14925 ( new_n17274 , new_n8615 , new_n17235 );
nor  g14926 ( new_n17275 , new_n11998 , new_n17274 );
nor  g14927 ( new_n17276 , new_n8632 , new_n12002 );
xnor g14928 ( new_n17277 , new_n11998 , new_n17274 );
nor  g14929 ( new_n17278 , new_n17276 , new_n17277 );
or   g14930 ( new_n17279 , new_n17275 , new_n17278 );
nor  g14931 ( new_n17280 , new_n17273 , new_n17279 );
or   g14932 ( new_n17281 , new_n17272 , new_n17280 );
nor  g14933 ( new_n17282 , new_n17270 , new_n17281 );
or   g14934 ( new_n17283 , new_n17269 , new_n17282 );
xnor g14935 ( new_n17284 , new_n17265 , new_n17266 );
nor  g14936 ( new_n17285_1 , new_n17283 , new_n17284 );
or   g14937 ( new_n17286 , new_n17267 , new_n17285_1 );
not  g14938 ( new_n17287 , new_n17286 );
and  g14939 ( new_n17288 , new_n17264 , new_n17287 );
nor  g14940 ( new_n17289 , new_n17263_1 , new_n17288 );
nor  g14941 ( new_n17290 , new_n17261 , new_n17289 );
nor  g14942 ( new_n17291 , new_n17260 , new_n17290 );
xnor g14943 ( n4451 , new_n17258 , new_n17291 );
xnor g14944 ( new_n17293 , n6659 , n25494 );
nor  g14945 ( new_n17294 , n10117 , new_n15667 );
xnor g14946 ( new_n17295 , n10117 , n23250 );
nor  g14947 ( new_n17296 , new_n15599 , n13460 );
xnor g14948 ( new_n17297 , n11455 , n13460 );
nor  g14949 ( new_n17298 , new_n15602_1 , n6104 );
xnor g14950 ( new_n17299 , n3945 , n6104 );
nor  g14951 ( new_n17300 , n4119 , new_n15605 );
and  g14952 ( new_n17301 , new_n5162 , new_n5183 );
or   g14953 ( new_n17302_1 , new_n17300 , new_n17301 );
and  g14954 ( new_n17303 , new_n17299 , new_n17302_1 );
or   g14955 ( new_n17304 , new_n17298 , new_n17303 );
and  g14956 ( new_n17305 , new_n17297 , new_n17304 );
or   g14957 ( new_n17306 , new_n17296 , new_n17305 );
and  g14958 ( new_n17307 , new_n17295 , new_n17306 );
or   g14959 ( new_n17308 , new_n17294 , new_n17307 );
xor  g14960 ( new_n17309 , new_n17293 , new_n17308 );
xor  g14961 ( new_n17310 , new_n12956_1 , new_n17309 );
xor  g14962 ( new_n17311 , new_n17295 , new_n17306 );
nor  g14963 ( new_n17312 , new_n12960 , new_n17311 );
xnor g14964 ( new_n17313 , new_n12960 , new_n17311 );
xor  g14965 ( new_n17314 , new_n17297 , new_n17304 );
nor  g14966 ( new_n17315 , new_n12964 , new_n17314 );
xnor g14967 ( new_n17316 , new_n12964 , new_n17314 );
not  g14968 ( new_n17317 , new_n17316 );
xor  g14969 ( new_n17318 , new_n17299 , new_n17302_1 );
and  g14970 ( new_n17319 , new_n12968 , new_n17318 );
xnor g14971 ( new_n17320_1 , new_n12970 , new_n17318 );
and  g14972 ( new_n17321 , new_n5160 , new_n5184_1 );
and  g14973 ( new_n17322 , new_n5185 , new_n5217 );
or   g14974 ( new_n17323 , new_n17321 , new_n17322 );
and  g14975 ( new_n17324 , new_n17320_1 , new_n17323 );
nor  g14976 ( new_n17325 , new_n17319 , new_n17324 );
and  g14977 ( new_n17326 , new_n17317 , new_n17325 );
nor  g14978 ( new_n17327 , new_n17315 , new_n17326 );
nor  g14979 ( new_n17328 , new_n17313 , new_n17327 );
nor  g14980 ( new_n17329 , new_n17312 , new_n17328 );
xor  g14981 ( n4476 , new_n17310 , new_n17329 );
not  g14982 ( new_n17331 , new_n11525 );
not  g14983 ( new_n17332 , new_n4003 );
nor  g14984 ( new_n17333 , n12398 , new_n17332 );
not  g14985 ( new_n17334 , new_n17333 );
nor  g14986 ( new_n17335 , n21317 , new_n17334 );
not  g14987 ( new_n17336 , new_n17335 );
nor  g14988 ( new_n17337_1 , n18452 , new_n17336 );
and  g14989 ( new_n17338 , new_n13645 , new_n17337_1 );
and  g14990 ( new_n17339 , new_n6152 , new_n17338 );
xnor g14991 ( new_n17340 , new_n6240 , new_n17339 );
xnor g14992 ( new_n17341 , n1831 , new_n17338 );
nor  g14993 ( new_n17342 , new_n6312 , new_n17341 );
xnor g14994 ( new_n17343 , n13137 , new_n17337_1 );
nor  g14995 ( new_n17344_1 , new_n6248_1 , new_n17343 );
xnor g14996 ( new_n17345 , new_n6248_1 , new_n17343 );
xnor g14997 ( new_n17346 , n18452 , new_n17335 );
nor  g14998 ( new_n17347 , new_n6254 , new_n17346 );
xnor g14999 ( new_n17348 , new_n6259 , new_n17346 );
xnor g15000 ( new_n17349 , n21317 , new_n17333 );
and  g15001 ( new_n17350 , new_n6264 , new_n17349 );
xnor g15002 ( new_n17351_1 , new_n6265 , new_n17349 );
and  g15003 ( new_n17352 , new_n4004 , new_n4043 );
and  g15004 ( new_n17353 , new_n4045 , new_n4076 );
or   g15005 ( new_n17354 , new_n17352 , new_n17353 );
and  g15006 ( new_n17355 , new_n17351_1 , new_n17354 );
nor  g15007 ( new_n17356 , new_n17350 , new_n17355 );
and  g15008 ( new_n17357 , new_n17348 , new_n17356 );
nor  g15009 ( new_n17358 , new_n17347 , new_n17357 );
nor  g15010 ( new_n17359_1 , new_n17345 , new_n17358 );
nor  g15011 ( new_n17360 , new_n17344_1 , new_n17359_1 );
xnor g15012 ( new_n17361 , new_n6312 , new_n17341 );
nor  g15013 ( new_n17362 , new_n17360 , new_n17361 );
nor  g15014 ( new_n17363 , new_n17342 , new_n17362 );
xnor g15015 ( new_n17364 , new_n17340 , new_n17363 );
xnor g15016 ( new_n17365 , new_n17331 , new_n17364 );
xnor g15017 ( new_n17366 , new_n17360 , new_n17361 );
nor  g15018 ( new_n17367 , new_n11530 , new_n17366 );
xnor g15019 ( new_n17368 , new_n11530 , new_n17366 );
xnor g15020 ( new_n17369 , new_n17345 , new_n17358 );
nor  g15021 ( new_n17370 , new_n11534 , new_n17369 );
xnor g15022 ( new_n17371 , new_n11534 , new_n17369 );
xnor g15023 ( new_n17372 , new_n17348 , new_n17356 );
nor  g15024 ( new_n17373 , new_n11539 , new_n17372 );
xnor g15025 ( new_n17374 , new_n11539 , new_n17372 );
xor  g15026 ( new_n17375 , new_n17351_1 , new_n17354 );
nor  g15027 ( new_n17376 , new_n11543 , new_n17375 );
xnor g15028 ( new_n17377 , new_n11543 , new_n17375 );
nor  g15029 ( new_n17378 , new_n3996 , new_n4077 );
nor  g15030 ( new_n17379 , new_n4078 , new_n4104 );
nor  g15031 ( new_n17380 , new_n17378 , new_n17379 );
nor  g15032 ( new_n17381 , new_n17377 , new_n17380 );
nor  g15033 ( new_n17382 , new_n17376 , new_n17381 );
nor  g15034 ( new_n17383 , new_n17374 , new_n17382 );
nor  g15035 ( new_n17384 , new_n17373 , new_n17383 );
nor  g15036 ( new_n17385 , new_n17371 , new_n17384 );
nor  g15037 ( new_n17386 , new_n17370 , new_n17385 );
nor  g15038 ( new_n17387_1 , new_n17368 , new_n17386 );
nor  g15039 ( new_n17388 , new_n17367 , new_n17387_1 );
xnor g15040 ( n4478 , new_n17365 , new_n17388 );
xnor g15041 ( n4529 , new_n12270 , new_n12302_1 );
xnor g15042 ( n4552 , new_n6099 , new_n6145 );
xnor g15043 ( n4595 , new_n6109 , new_n6141 );
xnor g15044 ( n4624 , new_n13948 , new_n13982 );
not  g15045 ( new_n17394 , new_n16886 );
nor  g15046 ( new_n17395 , n2659 , new_n17394 );
xnor g15047 ( new_n17396 , n2858 , new_n17395 );
nor  g15048 ( new_n17397 , n14899 , new_n17396 );
xnor g15049 ( new_n17398 , n14899 , new_n17396 );
nor  g15050 ( new_n17399 , n18444 , new_n16887 );
nor  g15051 ( new_n17400 , new_n16888 , new_n16896 );
nor  g15052 ( new_n17401 , new_n17399 , new_n17400 );
nor  g15053 ( new_n17402 , new_n17398 , new_n17401 );
nor  g15054 ( new_n17403 , new_n17397 , new_n17402 );
and  g15055 ( new_n17404 , new_n4909 , new_n17395 );
xnor g15056 ( new_n17405 , n3740 , new_n17404 );
xnor g15057 ( new_n17406 , new_n8323 , new_n17405 );
xnor g15058 ( new_n17407 , new_n17403 , new_n17406 );
nor  g15059 ( new_n17408 , new_n7703 , new_n17407 );
xnor g15060 ( new_n17409 , new_n7703 , new_n17407 );
xnor g15061 ( new_n17410 , new_n17398 , new_n17401 );
and  g15062 ( new_n17411 , new_n7706 , new_n17410 );
xnor g15063 ( new_n17412 , new_n7706 , new_n17410 );
nor  g15064 ( new_n17413 , new_n7715 , new_n16897 );
nor  g15065 ( new_n17414 , new_n16898 , new_n16906 );
nor  g15066 ( new_n17415 , new_n17413 , new_n17414 );
nor  g15067 ( new_n17416 , new_n17412 , new_n17415 );
nor  g15068 ( new_n17417 , new_n17411 , new_n17416 );
nor  g15069 ( new_n17418 , new_n17409 , new_n17417 );
nor  g15070 ( new_n17419 , new_n17408 , new_n17418 );
and  g15071 ( new_n17420 , new_n4907 , new_n17404 );
and  g15072 ( new_n17421_1 , n3506 , new_n17405 );
or   g15073 ( new_n17422 , n3506 , new_n17405 );
and  g15074 ( new_n17423 , new_n17403 , new_n17422 );
or   g15075 ( new_n17424 , new_n17421_1 , new_n17423 );
nor  g15076 ( new_n17425 , new_n17420 , new_n17424 );
xnor g15077 ( new_n17426 , new_n17419 , new_n17425 );
xnor g15078 ( new_n17427 , new_n7649 , new_n17426 );
not  g15079 ( new_n17428 , new_n17427 );
xnor g15080 ( new_n17429 , new_n13394 , new_n17428 );
xor  g15081 ( new_n17430 , new_n17409 , new_n17417 );
nor  g15082 ( new_n17431 , new_n7840 , new_n17430 );
xnor g15083 ( new_n17432_1 , new_n17412 , new_n17415 );
not  g15084 ( new_n17433 , new_n17432_1 );
nor  g15085 ( new_n17434 , new_n7849 , new_n17433 );
xnor g15086 ( new_n17435 , new_n7849 , new_n17433 );
not  g15087 ( new_n17436_1 , new_n16907 );
nor  g15088 ( new_n17437 , new_n7856 , new_n17436_1 );
xnor g15089 ( new_n17438 , new_n7856 , new_n17436_1 );
nor  g15090 ( new_n17439 , new_n7861 , new_n16920 );
xnor g15091 ( new_n17440_1 , new_n7860 , new_n16920 );
not  g15092 ( new_n17441 , new_n13044_1 );
nor  g15093 ( new_n17442 , new_n7866 , new_n17441 );
nor  g15094 ( new_n17443 , new_n7870 , new_n13068 );
nor  g15095 ( new_n17444 , new_n16741 , new_n16755 );
nor  g15096 ( new_n17445 , new_n17443 , new_n17444 );
xnor g15097 ( new_n17446 , new_n7866 , new_n13044_1 );
and  g15098 ( new_n17447 , new_n17445 , new_n17446 );
nor  g15099 ( new_n17448 , new_n17442 , new_n17447 );
and  g15100 ( new_n17449 , new_n17440_1 , new_n17448 );
nor  g15101 ( new_n17450_1 , new_n17439 , new_n17449 );
nor  g15102 ( new_n17451 , new_n17438 , new_n17450_1 );
nor  g15103 ( new_n17452 , new_n17437 , new_n17451 );
nor  g15104 ( new_n17453 , new_n17435 , new_n17452 );
nor  g15105 ( new_n17454 , new_n17434 , new_n17453 );
xnor g15106 ( new_n17455 , new_n7840 , new_n17430 );
nor  g15107 ( new_n17456 , new_n17454 , new_n17455 );
nor  g15108 ( new_n17457 , new_n17431 , new_n17456 );
xor  g15109 ( n4646 , new_n17429 , new_n17457 );
xnor g15110 ( n4674 , new_n13932 , new_n13990 );
xnor g15111 ( new_n17460 , n3480 , n7057 );
nor  g15112 ( new_n17461_1 , n8381 , new_n7625 );
nor  g15113 ( new_n17462 , new_n8510_1 , n16722 );
nor  g15114 ( new_n17463 , new_n5784 , n20235 );
or   g15115 ( new_n17464 , n11486 , new_n5040 );
nor  g15116 ( new_n17465 , n12495 , new_n2383 );
and  g15117 ( new_n17466_1 , new_n17464 , new_n17465 );
nor  g15118 ( new_n17467 , new_n17463 , new_n17466_1 );
nor  g15119 ( new_n17468 , new_n17462 , new_n17467 );
or   g15120 ( new_n17469 , new_n17461_1 , new_n17468 );
xor  g15121 ( new_n17470 , new_n17460 , new_n17469 );
xnor g15122 ( new_n17471 , new_n3052 , new_n17470 );
xnor g15123 ( new_n17472 , n8381 , n16722 );
xnor g15124 ( new_n17473 , new_n17467 , new_n17472 );
and  g15125 ( new_n17474 , new_n3057 , new_n17473 );
xnor g15126 ( new_n17475 , new_n3057 , new_n17473 );
xnor g15127 ( new_n17476 , n12495 , n13781 );
nor  g15128 ( new_n17477 , new_n3064 , new_n17476 );
nor  g15129 ( new_n17478 , new_n3069 , new_n17477 );
xnor g15130 ( new_n17479 , new_n3069 , new_n17477 );
xnor g15131 ( new_n17480 , n11486 , n20235 );
xnor g15132 ( new_n17481 , new_n17465 , new_n17480 );
nor  g15133 ( new_n17482 , new_n17479 , new_n17481 );
nor  g15134 ( new_n17483 , new_n17478 , new_n17482 );
nor  g15135 ( new_n17484 , new_n17475 , new_n17483 );
nor  g15136 ( new_n17485 , new_n17474 , new_n17484 );
xor  g15137 ( n4693 , new_n17471 , new_n17485 );
xnor g15138 ( n4731 , new_n10587 , new_n10597 );
nor  g15139 ( new_n17488 , new_n5981 , new_n6022_1 );
or   g15140 ( new_n17489 , new_n6028 , new_n6086 );
and  g15141 ( new_n17490 , new_n6024 , new_n17489 );
nor  g15142 ( new_n17491 , new_n17488 , new_n17490 );
nor  g15143 ( new_n17492 , n3582 , n21784 );
or   g15144 ( new_n17493_1 , new_n5984 , new_n6020 );
and  g15145 ( new_n17494 , new_n5983 , new_n17493_1 );
nor  g15146 ( new_n17495 , new_n17492 , new_n17494 );
not  g15147 ( new_n17496 , new_n17495 );
nor  g15148 ( new_n17497 , new_n17491 , new_n17496 );
not  g15149 ( new_n17498 , new_n17497 );
xnor g15150 ( new_n17499 , new_n15097 , new_n17498 );
xnor g15151 ( new_n17500_1 , new_n17491 , new_n17495 );
nor  g15152 ( new_n17501 , new_n15101 , new_n17500_1 );
xnor g15153 ( new_n17502 , new_n15101 , new_n17500_1 );
and  g15154 ( new_n17503 , new_n12670_1 , new_n12694 );
nor  g15155 ( new_n17504 , new_n12695 , new_n12732 );
nor  g15156 ( new_n17505 , new_n17503 , new_n17504 );
nor  g15157 ( new_n17506 , new_n17502 , new_n17505 );
nor  g15158 ( new_n17507 , new_n17501 , new_n17506 );
xnor g15159 ( n4745 , new_n17499 , new_n17507 );
xnor g15160 ( new_n17509 , n6773 , new_n6288 );
xnor g15161 ( n4747 , new_n9686 , new_n17509 );
xnor g15162 ( n4766 , new_n5746 , new_n5747 );
xnor g15163 ( n4770 , new_n13461 , new_n13478 );
xnor g15164 ( n4777 , new_n15308 , new_n16115 );
xnor g15165 ( new_n17514 , n6861 , n17959 );
and  g15166 ( new_n17515 , new_n5468 , n19357 );
xnor g15167 ( new_n17516 , n7566 , n19357 );
and  g15168 ( new_n17517 , n2328 , new_n5471 );
xnor g15169 ( new_n17518 , n2328 , n7731 );
nor  g15170 ( new_n17519 , new_n5475 , n15053 );
nor  g15171 ( new_n17520 , n12341 , new_n15611 );
nor  g15172 ( new_n17521 , new_n5478 , n25471 );
or   g15173 ( new_n17522 , n20986 , new_n5066 );
nor  g15174 ( new_n17523 , new_n5798 , n16502 );
and  g15175 ( new_n17524_1 , new_n17522 , new_n17523 );
nor  g15176 ( new_n17525 , new_n17521 , new_n17524_1 );
nor  g15177 ( new_n17526 , new_n17520 , new_n17525 );
nor  g15178 ( new_n17527 , new_n17519 , new_n17526 );
and  g15179 ( new_n17528 , new_n17518 , new_n17527 );
or   g15180 ( new_n17529_1 , new_n17517 , new_n17528 );
and  g15181 ( new_n17530 , new_n17516 , new_n17529_1 );
or   g15182 ( new_n17531 , new_n17515 , new_n17530 );
xor  g15183 ( new_n17532 , new_n17514 , new_n17531 );
nor  g15184 ( new_n17533 , n6794 , n20077 );
not  g15185 ( new_n17534 , new_n17533 );
nor  g15186 ( new_n17535 , n15636 , new_n17534 );
not  g15187 ( new_n17536 , new_n17535 );
nor  g15188 ( new_n17537 , n8745 , new_n17536 );
not  g15189 ( new_n17538 , new_n17537 );
nor  g15190 ( new_n17539 , n1777 , new_n17538 );
xnor g15191 ( new_n17540 , n22660 , new_n17539 );
xnor g15192 ( new_n17541 , n11580 , new_n17540 );
xnor g15193 ( new_n17542 , n1777 , new_n17537 );
nor  g15194 ( new_n17543 , new_n5576 , new_n17542 );
xnor g15195 ( new_n17544 , n15884 , new_n17542 );
xnor g15196 ( new_n17545 , n8745 , new_n17535 );
nor  g15197 ( new_n17546 , new_n5595 , new_n17545 );
xnor g15198 ( new_n17547 , new_n5595 , new_n17545 );
xnor g15199 ( new_n17548 , n15636 , new_n17533 );
nor  g15200 ( new_n17549 , new_n5582 , new_n17548 );
xnor g15201 ( new_n17550 , n27104 , new_n17548 );
xnor g15202 ( new_n17551 , new_n2447 , n20077 );
nor  g15203 ( new_n17552 , new_n5584 , new_n17551 );
nor  g15204 ( new_n17553 , new_n5588 , n6794 );
xnor g15205 ( new_n17554 , n27188 , new_n17551 );
and  g15206 ( new_n17555 , new_n17553 , new_n17554 );
or   g15207 ( new_n17556 , new_n17552 , new_n17555 );
and  g15208 ( new_n17557_1 , new_n17550 , new_n17556 );
nor  g15209 ( new_n17558 , new_n17549 , new_n17557_1 );
nor  g15210 ( new_n17559 , new_n17547 , new_n17558 );
or   g15211 ( new_n17560 , new_n17546 , new_n17559 );
and  g15212 ( new_n17561 , new_n17544 , new_n17560 );
or   g15213 ( new_n17562 , new_n17543 , new_n17561 );
xor  g15214 ( new_n17563 , new_n17541 , new_n17562 );
xnor g15215 ( new_n17564 , new_n15581 , new_n17563 );
xor  g15216 ( new_n17565 , new_n17544 , new_n17560 );
nor  g15217 ( new_n17566 , new_n14991 , new_n17565 );
xnor g15218 ( new_n17567 , new_n17547 , new_n17558 );
nor  g15219 ( new_n17568 , new_n14996 , new_n17567 );
xnor g15220 ( new_n17569 , new_n14994 , new_n17567 );
xor  g15221 ( new_n17570 , new_n17550 , new_n17556 );
nor  g15222 ( new_n17571 , new_n5037 , new_n17570 );
xnor g15223 ( new_n17572 , new_n5037 , new_n17570 );
xnor g15224 ( new_n17573 , new_n17553 , new_n17554 );
not  g15225 ( new_n17574 , new_n17573 );
nor  g15226 ( new_n17575 , new_n5048 , new_n17574 );
xnor g15227 ( new_n17576 , n6611 , n6794 );
nor  g15228 ( new_n17577 , new_n5042 , new_n17576 );
xnor g15229 ( new_n17578 , new_n5076 , new_n17574 );
and  g15230 ( new_n17579 , new_n17577 , new_n17578 );
nor  g15231 ( new_n17580 , new_n17575 , new_n17579 );
nor  g15232 ( new_n17581 , new_n17572 , new_n17580 );
nor  g15233 ( new_n17582 , new_n17571 , new_n17581 );
and  g15234 ( new_n17583_1 , new_n17569 , new_n17582 );
nor  g15235 ( new_n17584 , new_n17568 , new_n17583_1 );
xor  g15236 ( new_n17585 , new_n14991 , new_n17565 );
and  g15237 ( new_n17586 , new_n17584 , new_n17585 );
nor  g15238 ( new_n17587 , new_n17566 , new_n17586 );
xnor g15239 ( new_n17588 , new_n17564 , new_n17587 );
xnor g15240 ( new_n17589 , new_n17532 , new_n17588 );
xor  g15241 ( new_n17590 , new_n17516 , new_n17529_1 );
xor  g15242 ( new_n17591 , new_n17584 , new_n17585 );
nor  g15243 ( new_n17592_1 , new_n17590 , new_n17591 );
xnor g15244 ( new_n17593 , new_n17590 , new_n17591 );
xnor g15245 ( new_n17594 , new_n17569 , new_n17582 );
not  g15246 ( new_n17595 , new_n17594 );
xnor g15247 ( new_n17596 , new_n17518 , new_n17527 );
and  g15248 ( new_n17597 , new_n17595 , new_n17596 );
xnor g15249 ( new_n17598 , new_n17595 , new_n17596 );
xnor g15250 ( new_n17599 , new_n17572 , new_n17580 );
xnor g15251 ( new_n17600 , n12341 , n15053 );
xnor g15252 ( new_n17601 , new_n17525 , new_n17600 );
and  g15253 ( new_n17602 , new_n17599 , new_n17601 );
xnor g15254 ( new_n17603 , new_n17599 , new_n17601 );
xnor g15255 ( new_n17604 , new_n5041 , new_n17576 );
not  g15256 ( new_n17605 , new_n17604 );
xnor g15257 ( new_n17606 , n12384 , n16502 );
nor  g15258 ( new_n17607 , new_n17605 , new_n17606 );
xnor g15259 ( new_n17608 , n20986 , n25471 );
xnor g15260 ( new_n17609 , new_n17523 , new_n17608 );
nor  g15261 ( new_n17610 , new_n17607 , new_n17609 );
xnor g15262 ( new_n17611 , new_n17577 , new_n17578 );
not  g15263 ( new_n17612 , new_n17611 );
xnor g15264 ( new_n17613 , new_n17607 , new_n17609 );
nor  g15265 ( new_n17614 , new_n17612 , new_n17613 );
nor  g15266 ( new_n17615 , new_n17610 , new_n17614 );
nor  g15267 ( new_n17616 , new_n17603 , new_n17615 );
nor  g15268 ( new_n17617 , new_n17602 , new_n17616 );
nor  g15269 ( new_n17618 , new_n17598 , new_n17617 );
nor  g15270 ( new_n17619 , new_n17597 , new_n17618 );
nor  g15271 ( new_n17620 , new_n17593 , new_n17619 );
nor  g15272 ( new_n17621 , new_n17592_1 , new_n17620 );
xor  g15273 ( n4785 , new_n17589 , new_n17621 );
xnor g15274 ( n4804 , new_n13745 , new_n13777 );
xnor g15275 ( n4810 , new_n15298 , new_n15317 );
not  g15276 ( new_n17625 , n23166 );
nor  g15277 ( new_n17626 , n18105 , new_n17625 );
or   g15278 ( new_n17627 , new_n9080 , new_n9117 );
and  g15279 ( new_n17628 , new_n9078 , new_n17627 );
nor  g15280 ( new_n17629 , new_n17626 , new_n17628 );
nor  g15281 ( new_n17630 , new_n7961 , new_n10686 );
and  g15282 ( new_n17631 , new_n10687 , new_n10730 );
nor  g15283 ( new_n17632 , new_n17630 , new_n17631 );
and  g15284 ( new_n17633 , new_n10678 , new_n10685 );
not  g15285 ( new_n17634 , new_n17181 );
nor  g15286 ( new_n17635 , new_n17633 , new_n17634 );
and  g15287 ( new_n17636 , new_n17178 , new_n17633 );
nor  g15288 ( new_n17637 , new_n17635 , new_n17636 );
xnor g15289 ( new_n17638_1 , new_n8027_1 , new_n17637 );
xnor g15290 ( new_n17639 , new_n17632 , new_n17638_1 );
and  g15291 ( new_n17640 , new_n17629 , new_n17639 );
xnor g15292 ( new_n17641 , new_n17629 , new_n17639 );
and  g15293 ( new_n17642 , new_n9119 , new_n10731 );
nor  g15294 ( new_n17643 , new_n10732 , new_n10775_1 );
nor  g15295 ( new_n17644 , new_n17642 , new_n17643 );
nor  g15296 ( new_n17645 , new_n17641 , new_n17644 );
nor  g15297 ( new_n17646 , new_n17640 , new_n17645 );
or   g15298 ( new_n17647 , new_n8026 , new_n17637 );
and  g15299 ( new_n17648 , new_n17632 , new_n17647 );
and  g15300 ( new_n17649 , new_n8026 , new_n17637 );
or   g15301 ( new_n17650 , new_n17636 , new_n17649 );
or   g15302 ( new_n17651 , new_n17648 , new_n17650 );
nand g15303 ( n4814 , new_n17646 , new_n17651 );
xnor g15304 ( n4850 , new_n15908 , new_n15909 );
xnor g15305 ( n4891 , new_n16687 , new_n16726 );
xnor g15306 ( n4925 , new_n16855 , new_n16876 );
xnor g15307 ( n4947 , new_n15898 , new_n15915 );
xnor g15308 ( n4952 , new_n9377 , new_n9378 );
xnor g15309 ( new_n17658 , n6790 , n25068 );
not  g15310 ( new_n17659 , n2331 );
nor  g15311 ( new_n17660 , new_n17659 , n22879 );
xnor g15312 ( new_n17661 , n2331 , n22879 );
not  g15313 ( new_n17662 , n22631 );
nor  g15314 ( new_n17663 , n2117 , new_n17662 );
xnor g15315 ( new_n17664_1 , n2117 , n22631 );
and  g15316 ( new_n17665 , n5882 , new_n7993 );
nor  g15317 ( new_n17666 , n5882 , new_n7993 );
nor  g15318 ( new_n17667 , new_n9793 , n15258 );
nor  g15319 ( new_n17668 , n4588 , new_n9790 );
not  g15320 ( new_n17669 , new_n17668 );
nor  g15321 ( new_n17670 , n11775 , new_n7998 );
nor  g15322 ( new_n17671 , new_n17669 , new_n17670 );
nor  g15323 ( new_n17672 , new_n17667 , new_n17671 );
nor  g15324 ( new_n17673 , new_n17666 , new_n17672 );
nor  g15325 ( new_n17674 , new_n17665 , new_n17673 );
and  g15326 ( new_n17675 , new_n17664_1 , new_n17674 );
or   g15327 ( new_n17676 , new_n17663 , new_n17675 );
and  g15328 ( new_n17677 , new_n17661 , new_n17676 );
or   g15329 ( new_n17678 , new_n17660 , new_n17677 );
xor  g15330 ( new_n17679 , new_n17658 , new_n17678 );
xnor g15331 ( new_n17680 , new_n14940 , new_n17679 );
xor  g15332 ( new_n17681 , new_n17661 , new_n17676 );
nor  g15333 ( new_n17682 , new_n14948 , new_n17681 );
xnor g15334 ( new_n17683 , new_n14948 , new_n17681 );
xnor g15335 ( new_n17684 , new_n17664_1 , new_n17674 );
and  g15336 ( new_n17685 , new_n14952 , new_n17684 );
xnor g15337 ( new_n17686 , new_n14953 , new_n17684 );
xnor g15338 ( new_n17687_1 , n5882 , n16743 );
xnor g15339 ( new_n17688 , new_n17672 , new_n17687_1 );
nor  g15340 ( new_n17689 , new_n14956 , new_n17688 );
xnor g15341 ( new_n17690 , new_n14956 , new_n17688 );
xnor g15342 ( new_n17691 , n11775 , n15258 );
xnor g15343 ( new_n17692 , new_n17669 , new_n17691 );
nor  g15344 ( new_n17693 , new_n14960 , new_n17692 );
nor  g15345 ( new_n17694 , new_n14962 , new_n14744 );
xnor g15346 ( new_n17695 , new_n15203 , new_n17692 );
and  g15347 ( new_n17696 , new_n17694 , new_n17695 );
nor  g15348 ( new_n17697 , new_n17693 , new_n17696 );
nor  g15349 ( new_n17698 , new_n17690 , new_n17697 );
nor  g15350 ( new_n17699 , new_n17689 , new_n17698 );
and  g15351 ( new_n17700 , new_n17686 , new_n17699 );
nor  g15352 ( new_n17701 , new_n17685 , new_n17700 );
nor  g15353 ( new_n17702 , new_n17683 , new_n17701 );
nor  g15354 ( new_n17703 , new_n17682 , new_n17702 );
xor  g15355 ( new_n17704 , new_n17680 , new_n17703 );
xnor g15356 ( new_n17705 , new_n14871 , new_n17704 );
xnor g15357 ( new_n17706 , new_n17683 , new_n17701 );
nor  g15358 ( new_n17707 , new_n14874 , new_n17706 );
xnor g15359 ( new_n17708 , new_n14874 , new_n17706 );
xnor g15360 ( new_n17709 , new_n17686 , new_n17699 );
nor  g15361 ( new_n17710 , new_n13334 , new_n17709 );
not  g15362 ( new_n17711 , new_n17709 );
xnor g15363 ( new_n17712 , new_n13335 , new_n17711 );
xnor g15364 ( new_n17713 , new_n17690 , new_n17697 );
not  g15365 ( new_n17714 , new_n17713 );
nor  g15366 ( new_n17715 , new_n13341 , new_n17714 );
xnor g15367 ( new_n17716 , new_n13341 , new_n17714 );
not  g15368 ( new_n17717 , new_n14745 );
nor  g15369 ( new_n17718 , new_n9885 , new_n17717 );
nor  g15370 ( new_n17719 , new_n13384 , new_n17718 );
xnor g15371 ( new_n17720 , new_n13384 , new_n17718 );
xor  g15372 ( new_n17721_1 , new_n17694 , new_n17695 );
nor  g15373 ( new_n17722 , new_n17720 , new_n17721_1 );
nor  g15374 ( new_n17723 , new_n17719 , new_n17722 );
nor  g15375 ( new_n17724 , new_n17716 , new_n17723 );
nor  g15376 ( new_n17725 , new_n17715 , new_n17724 );
nor  g15377 ( new_n17726 , new_n17712 , new_n17725 );
nor  g15378 ( new_n17727 , new_n17710 , new_n17726 );
nor  g15379 ( new_n17728 , new_n17708 , new_n17727 );
nor  g15380 ( new_n17729 , new_n17707 , new_n17728 );
xnor g15381 ( n4966 , new_n17705 , new_n17729 );
xnor g15382 ( n4972 , new_n17199 , new_n17200 );
and  g15383 ( new_n17732 , new_n5453 , new_n7524_1 );
xnor g15384 ( new_n17733 , n23895 , new_n7524_1 );
nor  g15385 ( new_n17734 , new_n5456 , new_n7528 );
xnor g15386 ( new_n17735_1 , new_n5456 , new_n7528 );
nor  g15387 ( new_n17736 , new_n5459 , new_n7533 );
nor  g15388 ( new_n17737 , new_n16552 , new_n16563 );
nor  g15389 ( new_n17738_1 , new_n17736 , new_n17737 );
nor  g15390 ( new_n17739 , new_n17735_1 , new_n17738_1 );
nor  g15391 ( new_n17740 , new_n17734 , new_n17739 );
and  g15392 ( new_n17741 , new_n17733 , new_n17740 );
nor  g15393 ( new_n17742 , new_n17732 , new_n17741 );
not  g15394 ( new_n17743 , new_n17742 );
nor  g15395 ( new_n17744 , new_n7519 , new_n17743 );
not  g15396 ( new_n17745 , new_n17744 );
not  g15397 ( new_n17746_1 , new_n16516_1 );
nor  g15398 ( new_n17747 , n2289 , new_n17746_1 );
and  g15399 ( new_n17748 , new_n6744 , new_n17747 );
xnor g15400 ( new_n17749_1 , n2978 , new_n17748 );
xnor g15401 ( new_n17750 , new_n16488 , new_n17749_1 );
xnor g15402 ( new_n17751 , n23697 , new_n17747 );
and  g15403 ( new_n17752 , n337 , new_n17751 );
nor  g15404 ( new_n17753 , n337 , new_n17751 );
and  g15405 ( new_n17754 , n3228 , new_n16517_1 );
or   g15406 ( new_n17755 , n3228 , new_n16517_1 );
and  g15407 ( new_n17756 , new_n17755 , new_n16532 );
nor  g15408 ( new_n17757 , new_n17754 , new_n17756 );
nor  g15409 ( new_n17758 , new_n17753 , new_n17757 );
nor  g15410 ( new_n17759 , new_n17752 , new_n17758 );
xnor g15411 ( new_n17760 , new_n17750 , new_n17759 );
nor  g15412 ( new_n17761 , n25972 , new_n17760 );
xnor g15413 ( new_n17762 , new_n11842_1 , new_n17760 );
xnor g15414 ( new_n17763 , n337 , new_n17751 );
xnor g15415 ( new_n17764 , new_n17757 , new_n17763 );
not  g15416 ( new_n17765 , new_n17764 );
nor  g15417 ( new_n17766 , n21915 , new_n17765 );
nor  g15418 ( new_n17767 , n13775 , new_n16534 );
nor  g15419 ( new_n17768 , new_n16535 , new_n16550 );
or   g15420 ( new_n17769 , new_n17767 , new_n17768 );
xnor g15421 ( new_n17770 , new_n8646 , new_n17765 );
and  g15422 ( new_n17771 , new_n17769 , new_n17770 );
or   g15423 ( new_n17772 , new_n17766 , new_n17771 );
and  g15424 ( new_n17773 , new_n17762 , new_n17772 );
nor  g15425 ( new_n17774 , new_n17761 , new_n17773 );
not  g15426 ( new_n17775 , new_n17774 );
and  g15427 ( new_n17776 , new_n7429 , new_n17748 );
and  g15428 ( new_n17777 , n7593 , new_n17749_1 );
nor  g15429 ( new_n17778 , n7593 , new_n17749_1 );
nor  g15430 ( new_n17779 , new_n17778 , new_n17759 );
or   g15431 ( new_n17780 , new_n17777 , new_n17779 );
nor  g15432 ( new_n17781 , new_n17776 , new_n17780 );
not  g15433 ( new_n17782 , new_n17781 );
nor  g15434 ( new_n17783 , new_n17775 , new_n17782 );
xnor g15435 ( new_n17784_1 , new_n7519 , new_n17742 );
xnor g15436 ( new_n17785 , new_n17775 , new_n17781 );
nor  g15437 ( new_n17786 , new_n17784_1 , new_n17785 );
xnor g15438 ( new_n17787 , new_n17784_1 , new_n17785 );
xnor g15439 ( new_n17788 , new_n17733 , new_n17740 );
not  g15440 ( new_n17789 , new_n17788 );
xor  g15441 ( new_n17790 , new_n17762 , new_n17772 );
nor  g15442 ( new_n17791 , new_n17789 , new_n17790 );
xnor g15443 ( new_n17792 , new_n17788 , new_n17790 );
xnor g15444 ( new_n17793 , new_n17735_1 , new_n17738_1 );
xor  g15445 ( new_n17794 , new_n17769 , new_n17770 );
nor  g15446 ( new_n17795 , new_n17793 , new_n17794 );
nor  g15447 ( new_n17796 , new_n16551 , new_n16564 );
nor  g15448 ( new_n17797 , new_n16565 , new_n16581 );
or   g15449 ( new_n17798 , new_n17796 , new_n17797 );
xnor g15450 ( new_n17799 , new_n17793 , new_n17794 );
nor  g15451 ( new_n17800 , new_n17798 , new_n17799 );
or   g15452 ( new_n17801 , new_n17795 , new_n17800 );
and  g15453 ( new_n17802 , new_n17792 , new_n17801 );
or   g15454 ( new_n17803 , new_n17791 , new_n17802 );
nor  g15455 ( new_n17804 , new_n17787 , new_n17803 );
nor  g15456 ( new_n17805 , new_n17786 , new_n17804 );
xnor g15457 ( new_n17806 , new_n17783 , new_n17805 );
xnor g15458 ( n5011 , new_n17745 , new_n17806 );
nor  g15459 ( new_n17808 , n2944 , new_n10030 );
xnor g15460 ( new_n17809 , n2944 , n11220 );
not  g15461 ( new_n17810 , n22379 );
nor  g15462 ( new_n17811 , n767 , new_n17810 );
and  g15463 ( new_n17812 , new_n2849 , new_n2885 );
or   g15464 ( new_n17813 , new_n17811 , new_n17812 );
and  g15465 ( new_n17814 , new_n17809 , new_n17813 );
nor  g15466 ( new_n17815 , new_n17808 , new_n17814 );
not  g15467 ( new_n17816 , new_n17815 );
nor  g15468 ( new_n17817 , new_n12808 , new_n8954 );
or   g15469 ( new_n17818 , n2160 , n16544 );
nor  g15470 ( new_n17819 , n6814 , n10763 );
and  g15471 ( new_n17820_1 , new_n2888 , new_n2924 );
nor  g15472 ( new_n17821 , new_n17819 , new_n17820_1 );
and  g15473 ( new_n17822 , new_n17818 , new_n17821 );
nor  g15474 ( new_n17823 , new_n17817 , new_n17822 );
nor  g15475 ( new_n17824 , new_n14810 , new_n17823 );
not  g15476 ( new_n17825 , new_n17823 );
xnor g15477 ( new_n17826 , new_n14811 , new_n17825 );
not  g15478 ( new_n17827 , new_n14785 );
xnor g15479 ( new_n17828 , new_n12808 , n16544 );
xnor g15480 ( new_n17829 , new_n17821 , new_n17828 );
nor  g15481 ( new_n17830 , new_n17827 , new_n17829 );
not  g15482 ( new_n17831 , new_n17829 );
xnor g15483 ( new_n17832 , new_n17827 , new_n17831 );
nor  g15484 ( new_n17833 , new_n2925 , new_n14801_1 );
and  g15485 ( new_n17834 , new_n2970 , new_n3031 );
or   g15486 ( new_n17835 , new_n17833 , new_n17834 );
and  g15487 ( new_n17836 , new_n17832 , new_n17835 );
nor  g15488 ( new_n17837 , new_n17830 , new_n17836 );
nor  g15489 ( new_n17838 , new_n17826 , new_n17837 );
nor  g15490 ( new_n17839 , new_n17824 , new_n17838 );
nor  g15491 ( new_n17840 , new_n17816 , new_n17839 );
xnor g15492 ( new_n17841 , new_n17826 , new_n17837 );
not  g15493 ( new_n17842 , new_n17841 );
nor  g15494 ( new_n17843 , new_n17815 , new_n17842 );
nor  g15495 ( new_n17844 , new_n17816 , new_n17841 );
xor  g15496 ( new_n17845 , new_n17809 , new_n17813 );
xor  g15497 ( new_n17846 , new_n17832 , new_n17835 );
nor  g15498 ( new_n17847 , new_n17845 , new_n17846 );
xnor g15499 ( new_n17848 , new_n17845 , new_n17846 );
nor  g15500 ( new_n17849 , new_n2886_1 , new_n3032 );
nor  g15501 ( new_n17850 , new_n3033 , new_n3084 );
nor  g15502 ( new_n17851 , new_n17849 , new_n17850 );
nor  g15503 ( new_n17852 , new_n17848 , new_n17851 );
nor  g15504 ( new_n17853 , new_n17847 , new_n17852 );
nor  g15505 ( new_n17854 , new_n17844 , new_n17853 );
nor  g15506 ( new_n17855_1 , new_n17843 , new_n17854 );
nor  g15507 ( new_n17856 , new_n17840 , new_n17855_1 );
not  g15508 ( new_n17857 , new_n17839 );
nor  g15509 ( new_n17858 , new_n17815 , new_n17857 );
nor  g15510 ( new_n17859 , new_n17854 , new_n17858 );
nor  g15511 ( n5020 , new_n17856 , new_n17859 );
nor  g15512 ( new_n17861 , n11486 , n13781 );
not  g15513 ( new_n17862 , new_n17861 );
nor  g15514 ( new_n17863 , n16722 , new_n17862 );
not  g15515 ( new_n17864 , new_n17863 );
nor  g15516 ( new_n17865 , n3480 , new_n17864 );
xnor g15517 ( new_n17866 , n3018 , new_n17865 );
xnor g15518 ( new_n17867 , new_n2994 , new_n17866 );
xnor g15519 ( new_n17868 , n3480 , new_n17863 );
nor  g15520 ( new_n17869 , new_n2998 , new_n17868 );
xnor g15521 ( new_n17870 , new_n2998 , new_n17868 );
xnor g15522 ( new_n17871 , n16722 , new_n17861 );
nor  g15523 ( new_n17872 , new_n3003 , new_n17871 );
xnor g15524 ( new_n17873 , new_n3003 , new_n17871 );
xnor g15525 ( new_n17874 , new_n5784 , n13781 );
nor  g15526 ( new_n17875 , new_n3011 , new_n17874 );
nor  g15527 ( new_n17876 , n13781 , new_n3015 );
not  g15528 ( new_n17877_1 , new_n17876 );
xnor g15529 ( new_n17878 , new_n3011 , new_n17874 );
nor  g15530 ( new_n17879 , new_n17877_1 , new_n17878 );
nor  g15531 ( new_n17880 , new_n17875 , new_n17879 );
nor  g15532 ( new_n17881 , new_n17873 , new_n17880 );
nor  g15533 ( new_n17882 , new_n17872 , new_n17881 );
nor  g15534 ( new_n17883 , new_n17870 , new_n17882 );
nor  g15535 ( new_n17884 , new_n17869 , new_n17883 );
xor  g15536 ( new_n17885 , new_n17867 , new_n17884 );
xnor g15537 ( new_n17886 , new_n6926 , new_n17885 );
xor  g15538 ( new_n17887 , new_n17870 , new_n17882 );
and  g15539 ( new_n17888 , new_n6931 , new_n17887 );
xnor g15540 ( new_n17889_1 , new_n6931 , new_n17887 );
xor  g15541 ( new_n17890 , new_n17873 , new_n17880 );
and  g15542 ( new_n17891 , new_n6936 , new_n17890 );
xnor g15543 ( new_n17892 , new_n17876 , new_n17878 );
and  g15544 ( new_n17893 , new_n6943 , new_n17892 );
xnor g15545 ( new_n17894 , new_n2383 , new_n3015 );
nor  g15546 ( new_n17895 , new_n6947 , new_n17894 );
xnor g15547 ( new_n17896 , new_n6943 , new_n17892 );
nor  g15548 ( new_n17897 , new_n17895 , new_n17896 );
nor  g15549 ( new_n17898 , new_n17893 , new_n17897 );
xnor g15550 ( new_n17899 , new_n6936 , new_n17890 );
nor  g15551 ( new_n17900 , new_n17898 , new_n17899 );
nor  g15552 ( new_n17901 , new_n17891 , new_n17900 );
nor  g15553 ( new_n17902 , new_n17889_1 , new_n17901 );
nor  g15554 ( new_n17903 , new_n17888 , new_n17902 );
xnor g15555 ( n5024 , new_n17886 , new_n17903 );
xnor g15556 ( n5046 , new_n3684 , new_n3715 );
xnor g15557 ( n5062 , new_n3800 , new_n5848 );
xnor g15558 ( n5064 , new_n12326 , new_n12351 );
xnor g15559 ( new_n17908 , new_n11651 , n12495 );
not  g15560 ( new_n17909 , new_n17908 );
xnor g15561 ( new_n17910 , new_n2477 , new_n17909 );
xnor g15562 ( new_n17911_1 , n7428 , n9251 );
nor  g15563 ( new_n17912_1 , new_n17910 , new_n17911_1 );
nor  g15564 ( new_n17913 , n7428 , new_n2367 );
xnor g15565 ( new_n17914 , n10372 , n20138 );
xnor g15566 ( new_n17915 , new_n17913 , new_n17914 );
xnor g15567 ( new_n17916 , new_n17912_1 , new_n17915 );
nor  g15568 ( new_n17917 , new_n2477 , new_n17908 );
or   g15569 ( new_n17918 , new_n11651 , new_n5080 );
xnor g15570 ( new_n17919 , new_n6989 , n20235 );
xor  g15571 ( new_n17920 , new_n17918 , new_n17919 );
xnor g15572 ( new_n17921 , new_n2386 , new_n17920 );
xnor g15573 ( new_n17922 , new_n17917 , new_n17921 );
not  g15574 ( new_n17923 , new_n17922 );
xnor g15575 ( n5082 , new_n17916 , new_n17923 );
xnor g15576 ( n5120 , new_n13469 , new_n13470 );
xnor g15577 ( n5158 , new_n14609 , new_n14618 );
xnor g15578 ( n5168 , new_n15901 , new_n15913 );
not  g15579 ( new_n17928 , new_n16936 );
xnor g15580 ( new_n17929 , n6659 , new_n17928 );
not  g15581 ( new_n17930 , new_n14032 );
nor  g15582 ( new_n17931_1 , n23250 , new_n17930 );
xnor g15583 ( new_n17932 , new_n15667 , new_n17930 );
nor  g15584 ( new_n17933 , n11455 , new_n16954_1 );
xnor g15585 ( new_n17934 , new_n15599 , new_n16954_1 );
nor  g15586 ( new_n17935 , n3945 , new_n14038 );
xnor g15587 ( new_n17936 , new_n15602_1 , new_n14038 );
nor  g15588 ( new_n17937 , new_n15605 , new_n14043 );
xnor g15589 ( new_n17938 , n5255 , new_n14043 );
nor  g15590 ( new_n17939 , new_n5163 , new_n14048 );
and  g15591 ( new_n17940 , new_n15006 , new_n15020 );
or   g15592 ( new_n17941 , new_n17939 , new_n17940 );
and  g15593 ( new_n17942 , new_n17938 , new_n17941 );
nor  g15594 ( new_n17943 , new_n17937 , new_n17942 );
and  g15595 ( new_n17944 , new_n17936 , new_n17943 );
or   g15596 ( new_n17945 , new_n17935 , new_n17944 );
and  g15597 ( new_n17946 , new_n17934 , new_n17945 );
or   g15598 ( new_n17947 , new_n17933 , new_n17946 );
and  g15599 ( new_n17948_1 , new_n17932 , new_n17947 );
or   g15600 ( new_n17949 , new_n17931_1 , new_n17948_1 );
xor  g15601 ( new_n17950 , new_n17929 , new_n17949 );
xnor g15602 ( new_n17951 , new_n15597 , new_n17950 );
xor  g15603 ( new_n17952 , new_n17932 , new_n17947 );
and  g15604 ( new_n17953 , new_n15676 , new_n17952 );
xnor g15605 ( new_n17954_1 , new_n15676 , new_n17952 );
xor  g15606 ( new_n17955 , new_n17934 , new_n17945 );
and  g15607 ( new_n17956_1 , new_n15681 , new_n17955 );
xnor g15608 ( new_n17957 , new_n15681 , new_n17955 );
xnor g15609 ( new_n17958 , new_n17936 , new_n17943 );
nor  g15610 ( new_n17959_1 , new_n15686 , new_n17958 );
xnor g15611 ( new_n17960 , new_n15686 , new_n17958 );
xor  g15612 ( new_n17961 , new_n17938 , new_n17941 );
nor  g15613 ( new_n17962 , new_n15691 , new_n17961 );
xnor g15614 ( new_n17963_1 , new_n15691 , new_n17961 );
nor  g15615 ( new_n17964 , new_n15005 , new_n15021 );
nor  g15616 ( new_n17965 , new_n15022 , new_n15042 );
nor  g15617 ( new_n17966 , new_n17964 , new_n17965 );
nor  g15618 ( new_n17967 , new_n17963_1 , new_n17966 );
nor  g15619 ( new_n17968_1 , new_n17962 , new_n17967 );
nor  g15620 ( new_n17969 , new_n17960 , new_n17968_1 );
nor  g15621 ( new_n17970 , new_n17959_1 , new_n17969 );
nor  g15622 ( new_n17971 , new_n17957 , new_n17970 );
nor  g15623 ( new_n17972 , new_n17956_1 , new_n17971 );
nor  g15624 ( new_n17973 , new_n17954_1 , new_n17972 );
nor  g15625 ( new_n17974 , new_n17953 , new_n17973 );
xnor g15626 ( n5184 , new_n17951 , new_n17974 );
and  g15627 ( new_n17976_1 , new_n4417 , new_n4533 );
and  g15628 ( new_n17977 , new_n17976_1 , new_n4611 );
or   g15629 ( new_n17978 , new_n4417 , new_n4533 );
nor  g15630 ( new_n17979 , new_n17978 , new_n4611 );
or   g15631 ( n5228 , new_n17977 , new_n17979 );
not  g15632 ( new_n17981 , n1314 );
nor  g15633 ( new_n17982 , new_n17981 , n25494 );
and  g15634 ( new_n17983 , new_n11170 , new_n11185 );
nor  g15635 ( new_n17984 , new_n17982 , new_n17983 );
xnor g15636 ( new_n17985 , new_n7195 , new_n17984 );
nor  g15637 ( new_n17986 , new_n7118 , new_n11186 );
xnor g15638 ( new_n17987 , new_n7118 , new_n11186 );
nor  g15639 ( new_n17988 , new_n7122 , new_n11205 );
nor  g15640 ( new_n17989 , new_n12324_1 , new_n12353 );
nor  g15641 ( new_n17990 , new_n17988 , new_n17989 );
nor  g15642 ( new_n17991 , new_n17987 , new_n17990 );
nor  g15643 ( new_n17992 , new_n17986 , new_n17991 );
xnor g15644 ( n5256 , new_n17985 , new_n17992 );
xor  g15645 ( n5265 , new_n6658 , new_n6671_1 );
xnor g15646 ( n5273 , new_n16683 , new_n16728 );
xnor g15647 ( new_n17996 , n2289 , n20946 );
nor  g15648 ( new_n17997 , n1112 , new_n5275 );
xnor g15649 ( new_n17998_1 , n1112 , n7751 );
nor  g15650 ( new_n17999 , n20179 , new_n12889 );
and  g15651 ( new_n18000 , new_n16377 , new_n16392 );
or   g15652 ( new_n18001 , new_n17999 , new_n18000 );
and  g15653 ( new_n18002 , new_n17998_1 , new_n18001 );
or   g15654 ( new_n18003 , new_n17997 , new_n18002 );
xor  g15655 ( new_n18004 , new_n17996 , new_n18003 );
xnor g15656 ( new_n18005 , new_n7373 , new_n18004 );
xor  g15657 ( new_n18006 , new_n17998_1 , new_n18001 );
nor  g15658 ( new_n18007 , new_n7377_1 , new_n18006 );
xnor g15659 ( new_n18008 , new_n7377_1 , new_n18006 );
nor  g15660 ( new_n18009 , new_n7381 , new_n16393 );
nor  g15661 ( new_n18010 , new_n16394 , new_n16414 );
nor  g15662 ( new_n18011 , new_n18009 , new_n18010 );
nor  g15663 ( new_n18012 , new_n18008 , new_n18011 );
nor  g15664 ( new_n18013 , new_n18007 , new_n18012 );
xnor g15665 ( n5274 , new_n18005 , new_n18013 );
nor  g15666 ( new_n18015 , n20385 , n25316 );
not  g15667 ( new_n18016 , new_n18015 );
nor  g15668 ( new_n18017 , n919 , new_n18016 );
not  g15669 ( new_n18018 , new_n18017 );
nor  g15670 ( new_n18019 , n3918 , new_n18018 );
xnor g15671 ( new_n18020 , n6513 , new_n18019 );
xnor g15672 ( new_n18021 , new_n8814 , new_n18020 );
xnor g15673 ( new_n18022 , n3918 , new_n18017 );
nor  g15674 ( new_n18023 , new_n8821_1 , new_n18022 );
xnor g15675 ( new_n18024 , n919 , new_n18015 );
nor  g15676 ( new_n18025_1 , new_n11057 , new_n18024 );
xnor g15677 ( new_n18026 , new_n8825 , new_n18024 );
xnor g15678 ( new_n18027 , n20385 , n25316 );
nor  g15679 ( new_n18028 , new_n8830 , new_n18027 );
nor  g15680 ( new_n18029 , new_n4146_1 , new_n8832 );
xnor g15681 ( new_n18030 , new_n8835 , new_n18027 );
and  g15682 ( new_n18031 , new_n18029 , new_n18030 );
nor  g15683 ( new_n18032 , new_n18028 , new_n18031 );
and  g15684 ( new_n18033 , new_n18026 , new_n18032 );
nor  g15685 ( new_n18034 , new_n18025_1 , new_n18033 );
xnor g15686 ( new_n18035_1 , new_n8821_1 , new_n18022 );
nor  g15687 ( new_n18036 , new_n18034 , new_n18035_1 );
or   g15688 ( new_n18037 , new_n18023 , new_n18036 );
xor  g15689 ( new_n18038 , new_n18021 , new_n18037 );
not  g15690 ( new_n18039 , new_n18038 );
xnor g15691 ( new_n18040 , n19472 , new_n16166 );
nor  g15692 ( new_n18041 , new_n6846 , new_n16170 );
xnor g15693 ( new_n18042 , n25370 , new_n16170 );
nor  g15694 ( new_n18043_1 , new_n8605 , new_n16173 );
xnor g15695 ( new_n18044 , n24786 , new_n16173 );
and  g15696 ( new_n18045_1 , n27120 , new_n4132 );
or   g15697 ( new_n18046 , n23065 , new_n4136 );
xnor g15698 ( new_n18047 , new_n8628 , new_n4132 );
and  g15699 ( new_n18048 , new_n18046 , new_n18047 );
or   g15700 ( new_n18049 , new_n18045_1 , new_n18048 );
and  g15701 ( new_n18050 , new_n18044 , new_n18049 );
or   g15702 ( new_n18051 , new_n18043_1 , new_n18050 );
and  g15703 ( new_n18052 , new_n18042 , new_n18051 );
or   g15704 ( new_n18053 , new_n18041 , new_n18052 );
xor  g15705 ( new_n18054 , new_n18040 , new_n18053 );
xnor g15706 ( new_n18055 , new_n18039 , new_n18054 );
xor  g15707 ( new_n18056 , new_n18042 , new_n18051 );
xnor g15708 ( new_n18057 , new_n18034 , new_n18035_1 );
nor  g15709 ( new_n18058 , new_n18056 , new_n18057 );
xnor g15710 ( new_n18059_1 , new_n18056 , new_n18057 );
xor  g15711 ( new_n18060 , new_n18044 , new_n18049 );
xnor g15712 ( new_n18061_1 , new_n18026 , new_n18032 );
nor  g15713 ( new_n18062 , new_n18060 , new_n18061_1 );
xnor g15714 ( new_n18063 , new_n18060 , new_n18061_1 );
xnor g15715 ( new_n18064 , new_n18029 , new_n18030 );
not  g15716 ( new_n18065 , new_n18064 );
xor  g15717 ( new_n18066 , new_n18046 , new_n18047 );
nor  g15718 ( new_n18067 , new_n18065 , new_n18066 );
not  g15719 ( new_n18068 , new_n8911_1 );
xnor g15720 ( new_n18069 , new_n4109 , new_n4136 );
nor  g15721 ( new_n18070 , new_n18068 , new_n18069 );
xnor g15722 ( new_n18071_1 , new_n18065 , new_n18066 );
nor  g15723 ( new_n18072 , new_n18070 , new_n18071_1 );
nor  g15724 ( new_n18073 , new_n18067 , new_n18072 );
nor  g15725 ( new_n18074 , new_n18063 , new_n18073 );
nor  g15726 ( new_n18075 , new_n18062 , new_n18074 );
nor  g15727 ( new_n18076 , new_n18059_1 , new_n18075 );
nor  g15728 ( new_n18077 , new_n18058 , new_n18076 );
xnor g15729 ( n5300 , new_n18055 , new_n18077 );
and  g15730 ( new_n18079 , new_n7185 , new_n12918 );
and  g15731 ( new_n18080 , new_n7190_1 , new_n7193 );
nor  g15732 ( new_n18081 , new_n18079 , new_n18080 );
nor  g15733 ( new_n18082 , new_n17984 , new_n18081 );
not  g15734 ( new_n18083 , new_n18081 );
xnor g15735 ( new_n18084 , new_n17984 , new_n18083 );
nor  g15736 ( new_n18085 , new_n7195 , new_n17984 );
nor  g15737 ( new_n18086 , new_n17985 , new_n17992 );
nor  g15738 ( new_n18087 , new_n18085 , new_n18086 );
and  g15739 ( new_n18088 , new_n18084 , new_n18087 );
nor  g15740 ( n5325 , new_n18082 , new_n18088 );
xnor g15741 ( new_n18090 , n17458 , n25120 );
nor  g15742 ( new_n18091 , n1222 , n8363 );
xnor g15743 ( new_n18092 , n1222 , n8363 );
nor  g15744 ( new_n18093 , n14680 , n25240 );
xnor g15745 ( new_n18094 , n14680 , n25240 );
nor  g15746 ( new_n18095 , n10125 , n17250 );
xnor g15747 ( new_n18096 , new_n10414 , n17250 );
nor  g15748 ( new_n18097 , new_n10881 , new_n10506 );
or   g15749 ( new_n18098 , n8067 , n23160 );
nor  g15750 ( new_n18099 , n16524 , n20923 );
nor  g15751 ( new_n18100 , new_n12760 , new_n12763 );
nor  g15752 ( new_n18101 , new_n18099 , new_n18100 );
and  g15753 ( new_n18102 , new_n18098 , new_n18101 );
nor  g15754 ( new_n18103 , new_n18097 , new_n18102 );
and  g15755 ( new_n18104 , new_n18096 , new_n18103 );
nor  g15756 ( new_n18105_1 , new_n18095 , new_n18104 );
nor  g15757 ( new_n18106 , new_n18094 , new_n18105_1 );
nor  g15758 ( new_n18107 , new_n18093 , new_n18106 );
nor  g15759 ( new_n18108 , new_n18092 , new_n18107 );
nor  g15760 ( new_n18109 , new_n18091 , new_n18108 );
xnor g15761 ( new_n18110 , new_n18090 , new_n18109 );
nor  g15762 ( new_n18111 , n23272 , new_n18110 );
xnor g15763 ( new_n18112 , n23272 , new_n18110 );
xnor g15764 ( new_n18113 , new_n18092 , new_n18107 );
nor  g15765 ( new_n18114 , n11481 , new_n18113 );
xnor g15766 ( new_n18115 , n11481 , new_n18113 );
xnor g15767 ( new_n18116 , new_n18094 , new_n18105_1 );
nor  g15768 ( new_n18117 , n16439 , new_n18116 );
xnor g15769 ( new_n18118 , n16439 , new_n18116 );
xnor g15770 ( new_n18119 , new_n18096 , new_n18103 );
nor  g15771 ( new_n18120 , n15241 , new_n18119 );
xnor g15772 ( new_n18121 , n15241 , new_n18119 );
xnor g15773 ( new_n18122 , n8067 , n23160 );
xnor g15774 ( new_n18123 , new_n18101 , new_n18122 );
nor  g15775 ( new_n18124 , n7678 , new_n18123 );
xnor g15776 ( new_n18125 , new_n4373 , new_n18123 );
nor  g15777 ( new_n18126 , n3785 , new_n12764 );
nor  g15778 ( new_n18127 , new_n12765 , new_n12768 );
or   g15779 ( new_n18128 , new_n18126 , new_n18127 );
and  g15780 ( new_n18129 , new_n18125 , new_n18128 );
nor  g15781 ( new_n18130 , new_n18124 , new_n18129 );
nor  g15782 ( new_n18131 , new_n18121 , new_n18130 );
nor  g15783 ( new_n18132 , new_n18120 , new_n18131 );
nor  g15784 ( new_n18133 , new_n18118 , new_n18132 );
nor  g15785 ( new_n18134 , new_n18117 , new_n18133 );
nor  g15786 ( new_n18135 , new_n18115 , new_n18134 );
nor  g15787 ( new_n18136 , new_n18114 , new_n18135 );
nor  g15788 ( new_n18137 , new_n18112 , new_n18136 );
or   g15789 ( new_n18138 , new_n18111 , new_n18137 );
nor  g15790 ( new_n18139 , n17458 , n25120 );
nor  g15791 ( new_n18140 , new_n18090 , new_n18109 );
nor  g15792 ( new_n18141 , new_n18139 , new_n18140 );
not  g15793 ( new_n18142 , new_n18141 );
nor  g15794 ( new_n18143_1 , new_n18138 , new_n18142 );
not  g15795 ( new_n18144 , new_n18143_1 );
xnor g15796 ( new_n18145_1 , n12507 , n12702 );
nor  g15797 ( new_n18146 , n15077 , n26797 );
xnor g15798 ( new_n18147 , n15077 , n26797 );
nor  g15799 ( new_n18148 , n3710 , n23913 );
xnor g15800 ( new_n18149 , n3710 , n23913 );
nor  g15801 ( new_n18150 , n22554 , n26318 );
xnor g15802 ( new_n18151_1 , n22554 , n26318 );
nor  g15803 ( new_n18152_1 , n20429 , n26054 );
xnor g15804 ( new_n18153 , n20429 , n26054 );
nor  g15805 ( new_n18154 , n3909 , n19081 );
xnor g15806 ( new_n18155 , n3909 , n19081 );
nor  g15807 ( new_n18156 , n8309 , n23974 );
xnor g15808 ( new_n18157_1 , new_n8771 , n23974 );
nor  g15809 ( new_n18158 , new_n8050 , new_n8759 );
or   g15810 ( new_n18159 , n2146 , n19144 );
nor  g15811 ( new_n18160 , n12593 , n22173 );
nor  g15812 ( new_n18161 , new_n16370 , new_n16371 );
nor  g15813 ( new_n18162 , new_n18160 , new_n18161 );
and  g15814 ( new_n18163 , new_n18159 , new_n18162 );
nor  g15815 ( new_n18164 , new_n18158 , new_n18163 );
and  g15816 ( new_n18165 , new_n18157_1 , new_n18164 );
nor  g15817 ( new_n18166 , new_n18156 , new_n18165 );
nor  g15818 ( new_n18167 , new_n18155 , new_n18166 );
nor  g15819 ( new_n18168 , new_n18154 , new_n18167 );
nor  g15820 ( new_n18169 , new_n18153 , new_n18168 );
nor  g15821 ( new_n18170 , new_n18152_1 , new_n18169 );
nor  g15822 ( new_n18171_1 , new_n18151_1 , new_n18170 );
nor  g15823 ( new_n18172 , new_n18150 , new_n18171_1 );
nor  g15824 ( new_n18173 , new_n18149 , new_n18172 );
nor  g15825 ( new_n18174 , new_n18148 , new_n18173 );
nor  g15826 ( new_n18175 , new_n18147 , new_n18174 );
nor  g15827 ( new_n18176 , new_n18146 , new_n18175 );
xnor g15828 ( new_n18177 , new_n18145_1 , new_n18176 );
nor  g15829 ( new_n18178 , n12650 , new_n18177 );
xnor g15830 ( new_n18179 , n12650 , new_n18177 );
xnor g15831 ( new_n18180 , new_n18147 , new_n18174 );
nor  g15832 ( new_n18181 , n10201 , new_n18180 );
xnor g15833 ( new_n18182 , n10201 , new_n18180 );
xnor g15834 ( new_n18183 , new_n18149 , new_n18172 );
nor  g15835 ( new_n18184 , n10593 , new_n18183 );
xnor g15836 ( new_n18185 , n10593 , new_n18183 );
xnor g15837 ( new_n18186 , new_n18151_1 , new_n18170 );
nor  g15838 ( new_n18187 , n18290 , new_n18186 );
xnor g15839 ( new_n18188 , new_n18153 , new_n18168 );
nor  g15840 ( new_n18189 , n11580 , new_n18188 );
xnor g15841 ( new_n18190 , n11580 , new_n18188 );
xnor g15842 ( new_n18191 , new_n18155 , new_n18166 );
nor  g15843 ( new_n18192 , n15884 , new_n18191 );
xnor g15844 ( new_n18193_1 , n15884 , new_n18191 );
xnor g15845 ( new_n18194 , new_n18157_1 , new_n18164 );
nor  g15846 ( new_n18195 , n6356 , new_n18194 );
xnor g15847 ( new_n18196 , new_n8050 , n19144 );
xnor g15848 ( new_n18197 , new_n18162 , new_n18196 );
nor  g15849 ( new_n18198 , new_n5582 , new_n18197 );
xnor g15850 ( new_n18199 , n27104 , new_n18197 );
nor  g15851 ( new_n18200 , n27188 , new_n16372 );
and  g15852 ( new_n18201 , new_n16369 , new_n16373 );
nor  g15853 ( new_n18202 , new_n18200 , new_n18201 );
and  g15854 ( new_n18203 , new_n18199 , new_n18202 );
nor  g15855 ( new_n18204 , new_n18198 , new_n18203 );
xnor g15856 ( new_n18205 , new_n5595 , new_n18194 );
and  g15857 ( new_n18206 , new_n18204 , new_n18205 );
nor  g15858 ( new_n18207 , new_n18195 , new_n18206 );
nor  g15859 ( new_n18208 , new_n18193_1 , new_n18207 );
nor  g15860 ( new_n18209 , new_n18192 , new_n18208 );
nor  g15861 ( new_n18210 , new_n18190 , new_n18209 );
nor  g15862 ( new_n18211 , new_n18189 , new_n18210 );
xnor g15863 ( new_n18212 , n18290 , new_n18186 );
nor  g15864 ( new_n18213 , new_n18211 , new_n18212 );
nor  g15865 ( new_n18214 , new_n18187 , new_n18213 );
nor  g15866 ( new_n18215 , new_n18185 , new_n18214 );
nor  g15867 ( new_n18216 , new_n18184 , new_n18215 );
nor  g15868 ( new_n18217 , new_n18182 , new_n18216 );
nor  g15869 ( new_n18218 , new_n18181 , new_n18217 );
nor  g15870 ( new_n18219 , new_n18179 , new_n18218 );
nor  g15871 ( new_n18220 , new_n18178 , new_n18219 );
nor  g15872 ( new_n18221 , n12507 , n12702 );
nor  g15873 ( new_n18222 , new_n18145_1 , new_n18176 );
nor  g15874 ( new_n18223 , new_n18221 , new_n18222 );
and  g15875 ( new_n18224 , new_n18220 , new_n18223 );
xnor g15876 ( new_n18225 , new_n18144 , new_n18224 );
xnor g15877 ( new_n18226 , new_n18138 , new_n18141 );
xnor g15878 ( new_n18227_1 , new_n18220 , new_n18223 );
and  g15879 ( new_n18228 , new_n18226 , new_n18227_1 );
xnor g15880 ( new_n18229 , new_n18226 , new_n18227_1 );
xnor g15881 ( new_n18230 , new_n18112 , new_n18136 );
not  g15882 ( new_n18231 , new_n18230 );
xnor g15883 ( new_n18232_1 , new_n18179 , new_n18218 );
nor  g15884 ( new_n18233 , new_n18231 , new_n18232_1 );
xnor g15885 ( new_n18234 , new_n18231 , new_n18232_1 );
xnor g15886 ( new_n18235 , new_n18115 , new_n18134 );
not  g15887 ( new_n18236 , new_n18235 );
xnor g15888 ( new_n18237 , new_n18182 , new_n18216 );
nor  g15889 ( new_n18238_1 , new_n18236 , new_n18237 );
xnor g15890 ( new_n18239 , new_n18236 , new_n18237 );
xnor g15891 ( new_n18240 , new_n18118 , new_n18132 );
not  g15892 ( new_n18241_1 , new_n18240 );
xnor g15893 ( new_n18242 , new_n18185 , new_n18214 );
nor  g15894 ( new_n18243 , new_n18241_1 , new_n18242 );
xnor g15895 ( new_n18244 , new_n18241_1 , new_n18242 );
xnor g15896 ( new_n18245 , new_n18121 , new_n18130 );
not  g15897 ( new_n18246 , new_n18245 );
xnor g15898 ( new_n18247 , new_n18211 , new_n18212 );
nor  g15899 ( new_n18248 , new_n18246 , new_n18247 );
xnor g15900 ( new_n18249 , new_n18246 , new_n18247 );
xnor g15901 ( new_n18250 , new_n18190 , new_n18209 );
xor  g15902 ( new_n18251 , new_n18125 , new_n18128 );
nor  g15903 ( new_n18252 , new_n18250 , new_n18251 );
xnor g15904 ( new_n18253 , new_n18250 , new_n18251 );
xnor g15905 ( new_n18254_1 , new_n18193_1 , new_n18207 );
nor  g15906 ( new_n18255 , new_n12770 , new_n18254_1 );
xnor g15907 ( new_n18256 , new_n12770 , new_n18254_1 );
xnor g15908 ( new_n18257 , new_n18204 , new_n18205 );
nor  g15909 ( new_n18258 , new_n6652_1 , new_n18257 );
xor  g15910 ( new_n18259 , new_n18199 , new_n18202 );
nor  g15911 ( new_n18260 , new_n6657 , new_n18259 );
xnor g15912 ( new_n18261 , new_n6657 , new_n18259 );
not  g15913 ( new_n18262 , new_n18261 );
nor  g15914 ( new_n18263 , new_n16368 , new_n16374 );
nor  g15915 ( new_n18264 , new_n6663 , new_n16375 );
nor  g15916 ( new_n18265 , new_n18263 , new_n18264 );
and  g15917 ( new_n18266 , new_n18262 , new_n18265 );
nor  g15918 ( new_n18267 , new_n18260 , new_n18266 );
xnor g15919 ( new_n18268 , new_n6652_1 , new_n18257 );
nor  g15920 ( new_n18269 , new_n18267 , new_n18268 );
nor  g15921 ( new_n18270 , new_n18258 , new_n18269 );
nor  g15922 ( new_n18271 , new_n18256 , new_n18270 );
nor  g15923 ( new_n18272 , new_n18255 , new_n18271 );
nor  g15924 ( new_n18273 , new_n18253 , new_n18272 );
nor  g15925 ( new_n18274_1 , new_n18252 , new_n18273 );
nor  g15926 ( new_n18275 , new_n18249 , new_n18274_1 );
nor  g15927 ( new_n18276 , new_n18248 , new_n18275 );
nor  g15928 ( new_n18277 , new_n18244 , new_n18276 );
nor  g15929 ( new_n18278 , new_n18243 , new_n18277 );
nor  g15930 ( new_n18279 , new_n18239 , new_n18278 );
nor  g15931 ( new_n18280 , new_n18238_1 , new_n18279 );
nor  g15932 ( new_n18281 , new_n18234 , new_n18280 );
nor  g15933 ( new_n18282 , new_n18233 , new_n18281 );
nor  g15934 ( new_n18283 , new_n18229 , new_n18282 );
nor  g15935 ( new_n18284 , new_n18228 , new_n18283 );
xnor g15936 ( n5351 , new_n18225 , new_n18284 );
and  g15937 ( n5353 , new_n16071 , new_n16077 );
nor  g15938 ( new_n18287 , n2160 , new_n11670 );
nor  g15939 ( new_n18288_1 , new_n11671 , new_n11718 );
nor  g15940 ( new_n18289 , new_n18287 , new_n18288_1 );
not  g15941 ( new_n18290_1 , new_n18289 );
nor  g15942 ( new_n18291 , n2272 , n9934 );
and  g15943 ( new_n18292 , new_n11634 , new_n11669 );
nor  g15944 ( new_n18293 , new_n18291 , new_n18292 );
nor  g15945 ( new_n18294 , new_n18290_1 , new_n18293 );
and  g15946 ( new_n18295_1 , new_n14516 , new_n11725 );
or   g15947 ( new_n18296 , new_n7260 , new_n18295_1 );
nor  g15948 ( new_n18297 , new_n7264 , new_n11726 );
nor  g15949 ( new_n18298 , new_n11727 , new_n11740 );
nor  g15950 ( new_n18299 , new_n18297 , new_n18298 );
nor  g15951 ( new_n18300 , new_n18296 , new_n18299 );
xnor g15952 ( new_n18301_1 , new_n18294 , new_n18300 );
xnor g15953 ( new_n18302 , new_n18289 , new_n18293 );
not  g15954 ( new_n18303 , new_n7260 );
xnor g15955 ( new_n18304_1 , new_n18303 , new_n18295_1 );
xnor g15956 ( new_n18305 , new_n18299 , new_n18304_1 );
not  g15957 ( new_n18306 , new_n18305 );
and  g15958 ( new_n18307 , new_n18302 , new_n18306 );
xnor g15959 ( new_n18308 , new_n18302 , new_n18306 );
and  g15960 ( new_n18309 , new_n11719 , new_n11742 );
nor  g15961 ( new_n18310_1 , new_n11743 , new_n11789 );
nor  g15962 ( new_n18311_1 , new_n18309 , new_n18310_1 );
nor  g15963 ( new_n18312 , new_n18308 , new_n18311_1 );
nor  g15964 ( new_n18313 , new_n18307 , new_n18312 );
xnor g15965 ( n5399 , new_n18301_1 , new_n18313 );
nor  g15966 ( new_n18315 , new_n4798 , new_n17136 );
and  g15967 ( new_n18316 , new_n17138_1 , new_n17141 );
nor  g15968 ( new_n18317 , new_n18315 , new_n18316 );
nor  g15969 ( new_n18318 , new_n12443 , new_n13879 );
or   g15970 ( new_n18319 , n9934 , new_n13877 );
and  g15971 ( new_n18320 , new_n18319 , new_n17135 );
or   g15972 ( new_n18321 , new_n13920 , new_n18320 );
nor  g15973 ( new_n18322 , new_n18318 , new_n18321 );
not  g15974 ( new_n18323_1 , new_n18322 );
nor  g15975 ( new_n18324 , new_n18317 , new_n18323_1 );
xnor g15976 ( new_n18325 , new_n18300 , new_n18324 );
xnor g15977 ( new_n18326 , new_n18317 , new_n18322 );
nor  g15978 ( new_n18327 , new_n18305 , new_n18326 );
nor  g15979 ( new_n18328 , new_n11741_1 , new_n17142 );
nor  g15980 ( new_n18329 , new_n17143 , new_n17146 );
nor  g15981 ( new_n18330 , new_n18328 , new_n18329 );
xnor g15982 ( new_n18331 , new_n18305 , new_n18326 );
nor  g15983 ( new_n18332_1 , new_n18330 , new_n18331 );
nor  g15984 ( new_n18333 , new_n18327 , new_n18332_1 );
xnor g15985 ( n5403 , new_n18325 , new_n18333 );
xnor g15986 ( n5430 , new_n15288 , new_n15321 );
or   g15987 ( new_n18336 , new_n14300 , new_n14306 );
and  g15988 ( new_n18337 , new_n10348 , new_n14295 );
nor  g15989 ( new_n18338 , new_n10348 , new_n14295 );
nor  g15990 ( new_n18339 , new_n18338 , new_n14307 );
or   g15991 ( new_n18340 , new_n18337 , new_n18339 );
nor  g15992 ( new_n18341 , new_n10209 , new_n18340 );
and  g15993 ( n5439 , new_n18336 , new_n18341 );
xnor g15994 ( n5472 , new_n12076 , new_n12093 );
xnor g15995 ( n5485 , new_n8350 , new_n8385 );
xnor g15996 ( n5524 , new_n17787 , new_n17803 );
not  g15997 ( new_n18346 , new_n16088 );
nor  g15998 ( new_n18347 , new_n5953 , new_n18346 );
not  g15999 ( new_n18348 , new_n18347 );
nor  g16000 ( new_n18349 , new_n5947 , new_n18348 );
not  g16001 ( new_n18350_1 , new_n18349 );
nor  g16002 ( new_n18351 , new_n13213 , new_n18350_1 );
not  g16003 ( new_n18352 , new_n18351 );
nor  g16004 ( new_n18353 , new_n13211 , new_n18352 );
not  g16005 ( new_n18354 , new_n18353 );
nor  g16006 ( new_n18355 , new_n15842 , new_n18354 );
not  g16007 ( new_n18356 , new_n18355 );
nor  g16008 ( new_n18357 , new_n15838 , new_n18356 );
not  g16009 ( new_n18358 , new_n18357 );
nor  g16010 ( new_n18359 , new_n5921 , new_n18358 );
xnor g16011 ( new_n18360 , new_n5915 , new_n18359 );
nor  g16012 ( new_n18361 , new_n13511 , new_n18360 );
xnor g16013 ( new_n18362_1 , new_n13511 , new_n18360 );
xnor g16014 ( new_n18363 , new_n5921 , new_n18357 );
nor  g16015 ( new_n18364 , new_n13514 , new_n18363 );
xnor g16016 ( new_n18365 , new_n13514 , new_n18363 );
xnor g16017 ( new_n18366 , new_n15838 , new_n18355 );
nor  g16018 ( new_n18367 , new_n13518 , new_n18366 );
xnor g16019 ( new_n18368 , new_n13518 , new_n18366 );
xnor g16020 ( new_n18369 , new_n15842 , new_n18353 );
nor  g16021 ( new_n18370 , new_n13522 , new_n18369 );
xnor g16022 ( new_n18371 , new_n13522 , new_n18369 );
xnor g16023 ( new_n18372 , new_n13211 , new_n18351 );
nor  g16024 ( new_n18373 , new_n13526 , new_n18372 );
xnor g16025 ( new_n18374 , new_n13526 , new_n18372 );
xnor g16026 ( new_n18375 , new_n13213 , new_n18349 );
nor  g16027 ( new_n18376 , new_n13531 , new_n18375 );
xnor g16028 ( new_n18377_1 , new_n13531 , new_n18375 );
xnor g16029 ( new_n18378 , new_n5947 , new_n18347 );
nor  g16030 ( new_n18379 , new_n12853 , new_n17149 );
nor  g16031 ( new_n18380 , new_n17150 , new_n17153 );
nor  g16032 ( new_n18381 , new_n18379 , new_n18380 );
nor  g16033 ( new_n18382 , new_n18378 , new_n18381 );
xor  g16034 ( new_n18383 , new_n18378 , new_n18381 );
and  g16035 ( new_n18384 , new_n12851 , new_n18383 );
nor  g16036 ( new_n18385 , new_n18382 , new_n18384 );
nor  g16037 ( new_n18386 , new_n18377_1 , new_n18385 );
nor  g16038 ( new_n18387 , new_n18376 , new_n18386 );
nor  g16039 ( new_n18388 , new_n18374 , new_n18387 );
nor  g16040 ( new_n18389 , new_n18373 , new_n18388 );
nor  g16041 ( new_n18390 , new_n18371 , new_n18389 );
nor  g16042 ( new_n18391 , new_n18370 , new_n18390 );
nor  g16043 ( new_n18392 , new_n18368 , new_n18391 );
nor  g16044 ( new_n18393 , new_n18367 , new_n18392 );
nor  g16045 ( new_n18394 , new_n18365 , new_n18393 );
nor  g16046 ( new_n18395 , new_n18364 , new_n18394 );
nor  g16047 ( new_n18396 , new_n18362_1 , new_n18395 );
nor  g16048 ( new_n18397 , new_n18361 , new_n18396 );
and  g16049 ( new_n18398 , new_n5914 , new_n18359 );
nor  g16050 ( new_n18399 , new_n13194 , new_n18398 );
and  g16051 ( new_n18400 , new_n13190_1 , new_n18398 );
nor  g16052 ( new_n18401 , new_n18399 , new_n18400 );
xnor g16053 ( new_n18402 , new_n13553 , new_n18401 );
xnor g16054 ( new_n18403 , new_n18397 , new_n18402 );
nor  g16055 ( new_n18404 , new_n4796 , new_n18403 );
xnor g16056 ( new_n18405_1 , new_n4796 , new_n18403 );
xnor g16057 ( new_n18406 , new_n18362_1 , new_n18395 );
nor  g16058 ( new_n18407 , new_n4968 , new_n18406 );
xnor g16059 ( new_n18408 , new_n4968 , new_n18406 );
xnor g16060 ( new_n18409_1 , new_n18365 , new_n18393 );
nor  g16061 ( new_n18410 , new_n4972_1 , new_n18409_1 );
xnor g16062 ( new_n18411 , new_n4972_1 , new_n18409_1 );
xnor g16063 ( new_n18412 , new_n18368 , new_n18391 );
nor  g16064 ( new_n18413 , new_n4976 , new_n18412 );
xnor g16065 ( new_n18414_1 , new_n4976 , new_n18412 );
xnor g16066 ( new_n18415 , new_n18371 , new_n18389 );
nor  g16067 ( new_n18416 , new_n4980 , new_n18415 );
xnor g16068 ( new_n18417 , new_n4980 , new_n18415 );
xnor g16069 ( new_n18418_1 , new_n18374 , new_n18387 );
nor  g16070 ( new_n18419 , new_n4984 , new_n18418_1 );
xnor g16071 ( new_n18420 , new_n4984 , new_n18418_1 );
xnor g16072 ( new_n18421 , new_n18377_1 , new_n18385 );
nor  g16073 ( new_n18422 , new_n4988 , new_n18421 );
xnor g16074 ( new_n18423 , new_n4988 , new_n18421 );
xnor g16075 ( new_n18424 , new_n12851 , new_n18383 );
nor  g16076 ( new_n18425 , new_n4992 , new_n18424 );
xnor g16077 ( new_n18426 , new_n4992 , new_n18424 );
not  g16078 ( new_n18427 , new_n18426 );
nor  g16079 ( new_n18428 , new_n4998 , new_n17154 );
and  g16080 ( new_n18429 , new_n17155 , new_n17157 );
nor  g16081 ( new_n18430 , new_n18428 , new_n18429 );
and  g16082 ( new_n18431 , new_n18427 , new_n18430 );
nor  g16083 ( new_n18432 , new_n18425 , new_n18431 );
nor  g16084 ( new_n18433 , new_n18423 , new_n18432 );
nor  g16085 ( new_n18434 , new_n18422 , new_n18433 );
nor  g16086 ( new_n18435 , new_n18420 , new_n18434 );
nor  g16087 ( new_n18436 , new_n18419 , new_n18435 );
nor  g16088 ( new_n18437_1 , new_n18417 , new_n18436 );
nor  g16089 ( new_n18438 , new_n18416 , new_n18437_1 );
nor  g16090 ( new_n18439_1 , new_n18414_1 , new_n18438 );
nor  g16091 ( new_n18440 , new_n18413 , new_n18439_1 );
nor  g16092 ( new_n18441 , new_n18411 , new_n18440 );
nor  g16093 ( new_n18442 , new_n18410 , new_n18441 );
nor  g16094 ( new_n18443 , new_n18408 , new_n18442 );
nor  g16095 ( new_n18444_1 , new_n18407 , new_n18443 );
nor  g16096 ( new_n18445_1 , new_n18405_1 , new_n18444_1 );
or   g16097 ( new_n18446 , new_n18404 , new_n18445_1 );
nor  g16098 ( new_n18447 , new_n13553 , new_n18401 );
and  g16099 ( new_n18448 , new_n13553 , new_n18401 );
nor  g16100 ( new_n18449 , new_n18397 , new_n18448 );
nor  g16101 ( new_n18450 , new_n18447 , new_n18449 );
nor  g16102 ( new_n18451 , new_n18400 , new_n18450 );
xnor g16103 ( n5564 , new_n18446 , new_n18451 );
xnor g16104 ( n5593 , new_n6939 , new_n6952 );
xnor g16105 ( new_n18454 , new_n13941 , new_n17193 );
nor  g16106 ( new_n18455 , new_n13946 , new_n15987 );
xnor g16107 ( new_n18456 , new_n13946 , new_n15987 );
nor  g16108 ( new_n18457 , new_n13950 , new_n15992 );
xnor g16109 ( new_n18458 , new_n13950 , new_n15992 );
nor  g16110 ( new_n18459 , new_n13954 , new_n15059 );
xnor g16111 ( new_n18460 , new_n13954 , new_n15059 );
nor  g16112 ( new_n18461 , new_n13958 , new_n15063 );
and  g16113 ( new_n18462 , new_n16758 , new_n16767 );
nor  g16114 ( new_n18463 , new_n18461 , new_n18462 );
nor  g16115 ( new_n18464 , new_n18460 , new_n18463 );
nor  g16116 ( new_n18465 , new_n18459 , new_n18464 );
nor  g16117 ( new_n18466 , new_n18458 , new_n18465 );
nor  g16118 ( new_n18467_1 , new_n18457 , new_n18466 );
nor  g16119 ( new_n18468 , new_n18456 , new_n18467_1 );
nor  g16120 ( new_n18469 , new_n18455 , new_n18468 );
xnor g16121 ( n5603 , new_n18454 , new_n18469 );
xnor g16122 ( new_n18471 , n14440 , n17911 );
not  g16123 ( new_n18472 , n21997 );
nor  g16124 ( new_n18473 , n1654 , new_n18472 );
xnor g16125 ( new_n18474 , n1654 , n21997 );
nor  g16126 ( new_n18475 , n13783 , new_n8501 );
xnor g16127 ( new_n18476 , n13783 , n25119 );
nor  g16128 ( new_n18477 , new_n8503 , n26660 );
xnor g16129 ( new_n18478 , n1163 , n26660 );
nor  g16130 ( new_n18479 , n3018 , new_n8506 );
or   g16131 ( new_n18480 , new_n10550 , n18537 );
nor  g16132 ( new_n18481 , new_n2398 , n7057 );
and  g16133 ( new_n18482_1 , new_n17460 , new_n17469 );
nor  g16134 ( new_n18483_1 , new_n18481 , new_n18482_1 );
and  g16135 ( new_n18484 , new_n18480 , new_n18483_1 );
or   g16136 ( new_n18485 , new_n18479 , new_n18484 );
and  g16137 ( new_n18486 , new_n18478 , new_n18485 );
or   g16138 ( new_n18487 , new_n18477 , new_n18486 );
and  g16139 ( new_n18488 , new_n18476 , new_n18487 );
or   g16140 ( new_n18489 , new_n18475 , new_n18488 );
and  g16141 ( new_n18490 , new_n18474 , new_n18489 );
or   g16142 ( new_n18491 , new_n18473 , new_n18490 );
xor  g16143 ( new_n18492 , new_n18471 , new_n18491 );
xor  g16144 ( new_n18493 , new_n3032 , new_n18492 );
xor  g16145 ( new_n18494 , new_n18474 , new_n18489 );
nor  g16146 ( new_n18495 , new_n3035 , new_n18494 );
xnor g16147 ( new_n18496_1 , new_n3035 , new_n18494 );
xor  g16148 ( new_n18497 , new_n18476 , new_n18487 );
nor  g16149 ( new_n18498 , new_n3039 , new_n18497 );
xnor g16150 ( new_n18499 , new_n3039 , new_n18497 );
xor  g16151 ( new_n18500 , new_n18478 , new_n18485 );
nor  g16152 ( new_n18501 , new_n3043 , new_n18500 );
xnor g16153 ( new_n18502 , new_n3043 , new_n18500 );
not  g16154 ( new_n18503 , new_n18502 );
xnor g16155 ( new_n18504 , n3018 , n18537 );
xnor g16156 ( new_n18505 , new_n18483_1 , new_n18504 );
nor  g16157 ( new_n18506 , new_n3048 , new_n18505 );
nor  g16158 ( new_n18507 , new_n3053 , new_n17470 );
and  g16159 ( new_n18508 , new_n17471 , new_n17485 );
or   g16160 ( new_n18509_1 , new_n18507 , new_n18508 );
xnor g16161 ( new_n18510 , new_n3049 , new_n18505 );
and  g16162 ( new_n18511 , new_n18509_1 , new_n18510 );
nor  g16163 ( new_n18512 , new_n18506 , new_n18511 );
and  g16164 ( new_n18513_1 , new_n18503 , new_n18512 );
nor  g16165 ( new_n18514 , new_n18501 , new_n18513_1 );
nor  g16166 ( new_n18515_1 , new_n18499 , new_n18514 );
nor  g16167 ( new_n18516 , new_n18498 , new_n18515_1 );
nor  g16168 ( new_n18517 , new_n18496_1 , new_n18516 );
nor  g16169 ( new_n18518 , new_n18495 , new_n18517 );
xor  g16170 ( n5609 , new_n18493 , new_n18518 );
xnor g16171 ( n5634 , new_n13120 , new_n13137_1 );
nor  g16172 ( new_n18521 , n2978 , new_n3217 );
xnor g16173 ( new_n18522 , n2978 , n3425 );
nor  g16174 ( new_n18523 , new_n3198 , n23697 );
xnor g16175 ( new_n18524 , n9967 , n23697 );
nor  g16176 ( new_n18525 , n2289 , new_n7508 );
and  g16177 ( new_n18526 , new_n17996 , new_n18003 );
or   g16178 ( new_n18527 , new_n18525 , new_n18526 );
and  g16179 ( new_n18528 , new_n18524 , new_n18527 );
or   g16180 ( new_n18529 , new_n18523 , new_n18528 );
and  g16181 ( new_n18530 , new_n18522 , new_n18529 );
nor  g16182 ( new_n18531 , new_n18521 , new_n18530 );
nor  g16183 ( new_n18532 , new_n7322 , new_n18531 );
not  g16184 ( new_n18533 , new_n18531 );
nor  g16185 ( new_n18534 , new_n7323 , new_n18533 );
xor  g16186 ( new_n18535 , new_n18522 , new_n18529 );
nor  g16187 ( new_n18536 , new_n7365 , new_n18535 );
xnor g16188 ( new_n18537_1 , new_n7365 , new_n18535 );
xor  g16189 ( new_n18538 , new_n18524 , new_n18527 );
nor  g16190 ( new_n18539 , new_n7369 , new_n18538 );
xnor g16191 ( new_n18540 , new_n7369 , new_n18538 );
nor  g16192 ( new_n18541 , new_n7373 , new_n18004 );
nor  g16193 ( new_n18542 , new_n18005 , new_n18013 );
nor  g16194 ( new_n18543 , new_n18541 , new_n18542 );
nor  g16195 ( new_n18544 , new_n18540 , new_n18543 );
nor  g16196 ( new_n18545 , new_n18539 , new_n18544 );
nor  g16197 ( new_n18546 , new_n18537_1 , new_n18545 );
nor  g16198 ( new_n18547 , new_n18536 , new_n18546 );
nor  g16199 ( new_n18548 , new_n18534 , new_n18547 );
nor  g16200 ( new_n18549 , new_n18532 , new_n18548 );
nor  g16201 ( new_n18550 , new_n7242 , new_n18303 );
and  g16202 ( new_n18551 , new_n7261 , new_n7321 );
nor  g16203 ( new_n18552 , new_n18550 , new_n18551 );
not  g16204 ( new_n18553 , new_n18552 );
xnor g16205 ( new_n18554 , new_n18531 , new_n18553 );
xnor g16206 ( n5643 , new_n18549 , new_n18554 );
xnor g16207 ( new_n18556 , n5834 , n18035 );
nor  g16208 ( new_n18557 , new_n10431 , n13851 );
and  g16209 ( new_n18558_1 , new_n15121 , new_n15138 );
or   g16210 ( new_n18559 , new_n18557 , new_n18558_1 );
xor  g16211 ( new_n18560 , new_n18556 , new_n18559 );
xnor g16212 ( new_n18561 , new_n14681 , new_n18560 );
nor  g16213 ( new_n18562 , new_n14706 , new_n15139_1 );
xnor g16214 ( new_n18563 , new_n14706 , new_n15139_1 );
nor  g16215 ( new_n18564 , new_n14710 , new_n15141 );
xnor g16216 ( new_n18565 , new_n14710 , new_n15141 );
nor  g16217 ( new_n18566 , new_n14714 , new_n15144 );
xnor g16218 ( new_n18567 , new_n14714 , new_n15144 );
nor  g16219 ( new_n18568 , new_n14717 , new_n15149 );
nor  g16220 ( new_n18569 , new_n13370 , new_n13608 );
xnor g16221 ( new_n18570 , new_n13369 , new_n13609 );
and  g16222 ( new_n18571 , new_n13374 , new_n13622 );
xnor g16223 ( new_n18572_1 , new_n13374 , new_n13622 );
nor  g16224 ( new_n18573 , new_n13376 , new_n13629 );
nor  g16225 ( new_n18574_1 , new_n13381 , new_n18573 );
xnor g16226 ( new_n18575 , new_n13380 , new_n18573 );
and  g16227 ( new_n18576_1 , new_n13634 , new_n18575 );
nor  g16228 ( new_n18577 , new_n18574_1 , new_n18576_1 );
nor  g16229 ( new_n18578_1 , new_n18572_1 , new_n18577 );
nor  g16230 ( new_n18579 , new_n18571 , new_n18578_1 );
nor  g16231 ( new_n18580 , new_n18570 , new_n18579 );
nor  g16232 ( new_n18581 , new_n18569 , new_n18580 );
xnor g16233 ( new_n18582_1 , new_n14718 , new_n15147 );
nor  g16234 ( new_n18583_1 , new_n18581 , new_n18582_1 );
nor  g16235 ( new_n18584_1 , new_n18568 , new_n18583_1 );
nor  g16236 ( new_n18585 , new_n18567 , new_n18584_1 );
nor  g16237 ( new_n18586 , new_n18566 , new_n18585 );
nor  g16238 ( new_n18587 , new_n18565 , new_n18586 );
nor  g16239 ( new_n18588 , new_n18564 , new_n18587 );
nor  g16240 ( new_n18589 , new_n18563 , new_n18588 );
nor  g16241 ( new_n18590 , new_n18562 , new_n18589 );
xor  g16242 ( n5680 , new_n18561 , new_n18590 );
xnor g16243 ( n5687 , new_n14392 , new_n14393 );
xnor g16244 ( n5700 , new_n15439 , new_n15446 );
xor  g16245 ( n5732 , new_n10357 , new_n10405_1 );
xnor g16246 ( new_n18595 , n8381 , n23775 );
nor  g16247 ( new_n18596 , n8259 , n20235 );
and  g16248 ( new_n18597 , new_n17918 , new_n17919 );
nor  g16249 ( new_n18598 , new_n18596 , new_n18597 );
xnor g16250 ( new_n18599 , new_n18595 , new_n18598 );
xnor g16251 ( new_n18600 , new_n2395 , new_n18599 );
nor  g16252 ( new_n18601 , new_n2386 , new_n17920 );
nor  g16253 ( new_n18602 , new_n17917 , new_n17921 );
nor  g16254 ( new_n18603 , new_n18601 , new_n18602 );
xnor g16255 ( new_n18604 , new_n18600 , new_n18603 );
xnor g16256 ( new_n18605 , n6385 , n8869 );
nor  g16257 ( new_n18606 , n10372 , new_n2363_1 );
and  g16258 ( new_n18607 , new_n17913 , new_n17914 );
or   g16259 ( new_n18608 , new_n18606 , new_n18607 );
xor  g16260 ( new_n18609 , new_n18605 , new_n18608 );
xnor g16261 ( new_n18610_1 , new_n18604 , new_n18609 );
and  g16262 ( new_n18611 , new_n17912_1 , new_n17915 );
nor  g16263 ( new_n18612 , new_n17916 , new_n17922 );
nor  g16264 ( new_n18613 , new_n18611 , new_n18612 );
xnor g16265 ( n5742 , new_n18610_1 , new_n18613 );
xnor g16266 ( n5765 , new_n13387 , new_n13388 );
xnor g16267 ( n5776 , new_n12266 , new_n12304_1 );
xnor g16268 ( n5782 , new_n2800 , new_n2841 );
xnor g16269 ( new_n18618 , new_n8503 , n18901 );
nor  g16270 ( new_n18619 , n4376 , n18537 );
xnor g16271 ( new_n18620 , n4376 , n18537 );
nor  g16272 ( new_n18621 , n7057 , n14570 );
xnor g16273 ( new_n18622 , n7057 , n14570 );
nor  g16274 ( new_n18623 , n8381 , n23775 );
nor  g16275 ( new_n18624 , new_n18595 , new_n18598 );
nor  g16276 ( new_n18625 , new_n18623 , new_n18624 );
nor  g16277 ( new_n18626 , new_n18622 , new_n18625 );
nor  g16278 ( new_n18627 , new_n18621 , new_n18626 );
nor  g16279 ( new_n18628 , new_n18620 , new_n18627 );
or   g16280 ( new_n18629 , new_n18619 , new_n18628 );
xor  g16281 ( new_n18630 , new_n18618 , new_n18629 );
xor  g16282 ( new_n18631 , new_n2423 , new_n18630 );
xnor g16283 ( new_n18632 , new_n18620 , new_n18627 );
nor  g16284 ( new_n18633 , new_n2414 , new_n18632 );
xnor g16285 ( new_n18634 , new_n18622 , new_n18625 );
nor  g16286 ( new_n18635_1 , new_n2394 , new_n18599 );
and  g16287 ( new_n18636 , new_n18600 , new_n18603 );
nor  g16288 ( new_n18637 , new_n18635_1 , new_n18636 );
nor  g16289 ( new_n18638 , new_n18634 , new_n18637 );
xnor g16290 ( new_n18639 , new_n18634 , new_n18637 );
nor  g16291 ( new_n18640 , new_n2404 , new_n18639 );
or   g16292 ( new_n18641 , new_n18638 , new_n18640 );
xnor g16293 ( new_n18642 , new_n2415 , new_n18632 );
and  g16294 ( new_n18643 , new_n18641 , new_n18642 );
nor  g16295 ( new_n18644 , new_n18633 , new_n18643 );
xor  g16296 ( new_n18645 , new_n18631 , new_n18644 );
xnor g16297 ( new_n18646 , n7099 , n23068 );
nor  g16298 ( new_n18647 , new_n11685 , n19514 );
xnor g16299 ( new_n18648 , n12811 , n19514 );
nor  g16300 ( new_n18649_1 , new_n11689 , n10053 );
xnor g16301 ( new_n18650 , n1118 , n10053 );
nor  g16302 ( new_n18651 , new_n2947 , n25974 );
nor  g16303 ( new_n18652 , n8399 , new_n11693 );
nor  g16304 ( new_n18653_1 , n1630 , new_n3824 );
or   g16305 ( new_n18654 , new_n2909 , n9507 );
nor  g16306 ( new_n18655 , n1451 , new_n2952 );
and  g16307 ( new_n18656 , new_n18654 , new_n18655 );
nor  g16308 ( new_n18657 , new_n18653_1 , new_n18656 );
nor  g16309 ( new_n18658 , new_n18652 , new_n18657 );
nor  g16310 ( new_n18659 , new_n18651 , new_n18658 );
and  g16311 ( new_n18660 , new_n18650 , new_n18659 );
or   g16312 ( new_n18661 , new_n18649_1 , new_n18660 );
and  g16313 ( new_n18662 , new_n18648 , new_n18661 );
or   g16314 ( new_n18663 , new_n18647 , new_n18662 );
xor  g16315 ( new_n18664 , new_n18646 , new_n18663 );
xnor g16316 ( new_n18665 , new_n18645 , new_n18664 );
not  g16317 ( new_n18666 , new_n18665 );
xor  g16318 ( new_n18667 , new_n18648 , new_n18661 );
not  g16319 ( new_n18668 , new_n18667 );
nor  g16320 ( new_n18669 , new_n18638 , new_n18640 );
xnor g16321 ( new_n18670 , new_n18669 , new_n18642 );
nor  g16322 ( new_n18671 , new_n18668 , new_n18670 );
xnor g16323 ( new_n18672 , new_n2405 , new_n18639 );
xnor g16324 ( new_n18673 , new_n18650 , new_n18659 );
and  g16325 ( new_n18674 , new_n18672 , new_n18673 );
xnor g16326 ( new_n18675 , new_n18672 , new_n18673 );
not  g16327 ( new_n18676 , new_n18604 );
xnor g16328 ( new_n18677 , n8399 , n25974 );
xnor g16329 ( new_n18678 , new_n18657 , new_n18677 );
and  g16330 ( new_n18679_1 , new_n18676 , new_n18678 );
xnor g16331 ( new_n18680 , new_n18676 , new_n18678 );
xnor g16332 ( new_n18681 , n1451 , n26979 );
nor  g16333 ( new_n18682 , new_n17910 , new_n18681 );
xnor g16334 ( new_n18683 , n1630 , n9507 );
xnor g16335 ( new_n18684 , new_n18655 , new_n18683 );
nor  g16336 ( new_n18685 , new_n18682 , new_n18684 );
xnor g16337 ( new_n18686 , new_n18682 , new_n18684 );
nor  g16338 ( new_n18687 , new_n17923 , new_n18686 );
nor  g16339 ( new_n18688 , new_n18685 , new_n18687 );
nor  g16340 ( new_n18689 , new_n18680 , new_n18688 );
nor  g16341 ( new_n18690_1 , new_n18679_1 , new_n18689 );
nor  g16342 ( new_n18691 , new_n18675 , new_n18690_1 );
nor  g16343 ( new_n18692 , new_n18674 , new_n18691 );
xnor g16344 ( new_n18693_1 , new_n18667 , new_n18670 );
and  g16345 ( new_n18694 , new_n18692 , new_n18693_1 );
nor  g16346 ( new_n18695 , new_n18671 , new_n18694 );
xnor g16347 ( n5833 , new_n18666 , new_n18695 );
xnor g16348 ( n5840 , new_n12274 , new_n12300 );
xor  g16349 ( n5841 , new_n18509_1 , new_n18510 );
xnor g16350 ( n5850 , new_n12743 , new_n12744 );
xnor g16351 ( n5903 , new_n18570 , new_n18579 );
xnor g16352 ( new_n18701 , n19042 , new_n16163 );
nor  g16353 ( new_n18702 , new_n8572 , new_n16166 );
and  g16354 ( new_n18703 , new_n18040 , new_n18053 );
or   g16355 ( new_n18704 , new_n18702 , new_n18703 );
xor  g16356 ( new_n18705 , new_n18701 , new_n18704 );
not  g16357 ( new_n18706 , new_n18019 );
nor  g16358 ( new_n18707 , n6513 , new_n18706 );
xnor g16359 ( new_n18708_1 , n26752 , new_n18707 );
xnor g16360 ( new_n18709 , new_n8807 , new_n18708_1 );
nor  g16361 ( new_n18710 , new_n8813 , new_n18020 );
and  g16362 ( new_n18711 , new_n18021 , new_n18037 );
nor  g16363 ( new_n18712 , new_n18710 , new_n18711 );
xnor g16364 ( new_n18713 , new_n18709 , new_n18712 );
xnor g16365 ( new_n18714 , new_n18705 , new_n18713 );
nor  g16366 ( new_n18715 , new_n18039 , new_n18054 );
nor  g16367 ( new_n18716 , new_n18055 , new_n18077 );
nor  g16368 ( new_n18717 , new_n18715 , new_n18716 );
xnor g16369 ( n5904 , new_n18714 , new_n18717 );
xnor g16370 ( new_n18719 , n6814 , n27089 );
nor  g16371 ( new_n18720 , n11841 , new_n8959 );
xnor g16372 ( new_n18721_1 , n11841 , n19701 );
nor  g16373 ( new_n18722 , n10710 , new_n8962 );
xnor g16374 ( new_n18723 , n10710 , n23529 );
nor  g16375 ( new_n18724 , n20929 , new_n8965 );
xnor g16376 ( new_n18725_1 , n20929 , n24620 );
nor  g16377 ( new_n18726 , new_n8968 , n8006 );
xnor g16378 ( new_n18727 , n5211 , n8006 );
nor  g16379 ( new_n18728 , new_n8971_1 , n25074 );
xnor g16380 ( new_n18729 , n12956 , n25074 );
nor  g16381 ( new_n18730 , new_n4328 , n18295 );
nor  g16382 ( new_n18731 , n16396 , new_n2903 );
nor  g16383 ( new_n18732 , n6502 , new_n4331 );
nor  g16384 ( new_n18733 , new_n5033 , n9399 );
nor  g16385 ( new_n18734 , new_n2951 , n15780 );
not  g16386 ( new_n18735 , new_n18734 );
nor  g16387 ( new_n18736 , new_n18733 , new_n18735 );
nor  g16388 ( new_n18737_1 , new_n18732 , new_n18736 );
nor  g16389 ( new_n18738 , new_n18731 , new_n18737_1 );
nor  g16390 ( new_n18739 , new_n18730 , new_n18738 );
and  g16391 ( new_n18740 , new_n18729 , new_n18739 );
or   g16392 ( new_n18741 , new_n18728 , new_n18740 );
and  g16393 ( new_n18742 , new_n18727 , new_n18741 );
or   g16394 ( new_n18743 , new_n18726 , new_n18742 );
and  g16395 ( new_n18744 , new_n18725_1 , new_n18743 );
or   g16396 ( new_n18745_1 , new_n18724 , new_n18744 );
and  g16397 ( new_n18746 , new_n18723 , new_n18745_1 );
or   g16398 ( new_n18747 , new_n18722 , new_n18746 );
and  g16399 ( new_n18748 , new_n18721_1 , new_n18747 );
or   g16400 ( new_n18749 , new_n18720 , new_n18748 );
xor  g16401 ( new_n18750 , new_n18719 , new_n18749 );
xnor g16402 ( new_n18751_1 , new_n10106 , new_n18750 );
xor  g16403 ( new_n18752 , new_n18721_1 , new_n18747 );
nor  g16404 ( new_n18753 , new_n10110 , new_n18752 );
xnor g16405 ( new_n18754 , new_n10110 , new_n18752 );
xor  g16406 ( new_n18755 , new_n18723 , new_n18745_1 );
nor  g16407 ( new_n18756 , new_n10114 , new_n18755 );
xnor g16408 ( new_n18757 , new_n10114 , new_n18755 );
xor  g16409 ( new_n18758 , new_n18725_1 , new_n18743 );
nor  g16410 ( new_n18759 , new_n10118 , new_n18758 );
xor  g16411 ( new_n18760 , new_n18727 , new_n18741 );
nor  g16412 ( new_n18761 , new_n10121 , new_n18760 );
xnor g16413 ( new_n18762 , new_n10121 , new_n18760 );
xnor g16414 ( new_n18763 , new_n18729 , new_n18739 );
and  g16415 ( new_n18764 , new_n10124 , new_n18763 );
xnor g16416 ( new_n18765 , n16396 , n18295 );
xnor g16417 ( new_n18766 , new_n18737_1 , new_n18765 );
and  g16418 ( new_n18767 , new_n10128 , new_n18766 );
xnor g16419 ( new_n18768 , new_n10132 , new_n18766 );
xnor g16420 ( new_n18769 , n2088 , n15780 );
nor  g16421 ( new_n18770 , new_n10134 , new_n18769 );
xnor g16422 ( new_n18771 , n6502 , n9399 );
xnor g16423 ( new_n18772 , new_n18735 , new_n18771 );
not  g16424 ( new_n18773 , new_n18772 );
and  g16425 ( new_n18774 , new_n18770 , new_n18773 );
xnor g16426 ( new_n18775 , new_n18770 , new_n18773 );
nor  g16427 ( new_n18776 , new_n10142 , new_n18775 );
nor  g16428 ( new_n18777 , new_n18774 , new_n18776 );
and  g16429 ( new_n18778 , new_n18768 , new_n18777 );
nor  g16430 ( new_n18779 , new_n18767 , new_n18778 );
xnor g16431 ( new_n18780_1 , new_n10124 , new_n18763 );
nor  g16432 ( new_n18781 , new_n18779 , new_n18780_1 );
nor  g16433 ( new_n18782_1 , new_n18764 , new_n18781 );
nor  g16434 ( new_n18783 , new_n18762 , new_n18782_1 );
nor  g16435 ( new_n18784 , new_n18761 , new_n18783 );
xnor g16436 ( new_n18785 , new_n10118 , new_n18758 );
nor  g16437 ( new_n18786 , new_n18784 , new_n18785 );
nor  g16438 ( new_n18787 , new_n18759 , new_n18786 );
nor  g16439 ( new_n18788 , new_n18757 , new_n18787 );
nor  g16440 ( new_n18789 , new_n18756 , new_n18788 );
nor  g16441 ( new_n18790 , new_n18754 , new_n18789 );
nor  g16442 ( new_n18791 , new_n18753 , new_n18790 );
xnor g16443 ( n5911 , new_n18751_1 , new_n18791 );
xnor g16444 ( n5936 , new_n3913 , new_n11769 );
xnor g16445 ( n5943 , new_n9936 , new_n9976 );
xnor g16446 ( n5964 , new_n13952 , new_n13980 );
nor  g16447 ( new_n18796 , n11184 , new_n5070 );
nor  g16448 ( new_n18797 , n23146 , new_n5057 );
or   g16449 ( new_n18798 , n17968 , new_n5082_1 );
nor  g16450 ( new_n18799 , new_n5061 , new_n18798 );
nor  g16451 ( new_n18800 , new_n18797 , new_n18799 );
nor  g16452 ( new_n18801 , new_n5071 , new_n18800 );
nor  g16453 ( new_n18802_1 , new_n18796 , new_n18801 );
and  g16454 ( new_n18803 , new_n15641 , new_n18802_1 );
nor  g16455 ( new_n18804 , new_n15648 , new_n18802_1 );
nor  g16456 ( new_n18805 , new_n15640 , new_n18804 );
nor  g16457 ( new_n18806 , new_n18803 , new_n18805 );
nor  g16458 ( new_n18807 , new_n15636_1 , new_n18806 );
nand g16459 ( new_n18808 , new_n15638 , new_n18806 );
and  g16460 ( new_n18809 , n8943 , new_n18808 );
nor  g16461 ( new_n18810 , new_n18807 , new_n18809 );
nor  g16462 ( new_n18811 , new_n15633 , new_n18810 );
nand g16463 ( new_n18812 , new_n15635 , new_n18810 );
and  g16464 ( new_n18813 , n12380 , new_n18812 );
nor  g16465 ( new_n18814 , new_n18811 , new_n18813 );
nor  g16466 ( new_n18815 , new_n15631 , new_n18814 );
nand g16467 ( new_n18816 , new_n15656 , new_n18814 );
and  g16468 ( new_n18817 , n8694 , new_n18816 );
nor  g16469 ( new_n18818 , new_n18815 , new_n18817 );
nor  g16470 ( new_n18819 , new_n15629 , new_n18818 );
and  g16471 ( new_n18820 , new_n15682 , new_n18818 );
nor  g16472 ( new_n18821 , new_n15660 , new_n18820 );
or   g16473 ( new_n18822 , new_n18819 , new_n18821 );
xor  g16474 ( new_n18823 , new_n15628 , new_n18822 );
xnor g16475 ( new_n18824 , new_n3224 , new_n18823 );
xnor g16476 ( new_n18825 , new_n15661 , new_n18818 );
and  g16477 ( new_n18826 , new_n3228_1 , new_n18825 );
xnor g16478 ( new_n18827 , new_n3228_1 , new_n18825 );
xnor g16479 ( new_n18828 , new_n15657 , new_n18814 );
and  g16480 ( new_n18829 , new_n3233 , new_n18828 );
xnor g16481 ( new_n18830_1 , new_n3233 , new_n18828 );
xor  g16482 ( new_n18831_1 , new_n15635 , new_n18810 );
and  g16483 ( new_n18832 , new_n3238 , new_n18831_1 );
xnor g16484 ( new_n18833 , new_n3238 , new_n18831_1 );
xnor g16485 ( new_n18834 , new_n15639 , new_n18806 );
and  g16486 ( new_n18835 , new_n3243 , new_n18834 );
xnor g16487 ( new_n18836 , new_n3243 , new_n18834 );
xnor g16488 ( new_n18837 , new_n15649 , new_n18802_1 );
and  g16489 ( new_n18838 , new_n3248 , new_n18837 );
xnor g16490 ( new_n18839 , new_n3248 , new_n18837 );
xnor g16491 ( new_n18840 , new_n15645 , new_n18800 );
and  g16492 ( new_n18841 , new_n3253_1 , new_n18840 );
xnor g16493 ( new_n18842 , new_n3253_1 , new_n18840 );
xnor g16494 ( new_n18843_1 , new_n5074 , new_n18798 );
and  g16495 ( new_n18844 , new_n3261 , new_n18843_1 );
nor  g16496 ( new_n18845 , new_n3257 , new_n5084 );
xnor g16497 ( new_n18846 , new_n3261 , new_n18843_1 );
nor  g16498 ( new_n18847 , new_n18845 , new_n18846 );
nor  g16499 ( new_n18848 , new_n18844 , new_n18847 );
nor  g16500 ( new_n18849 , new_n18842 , new_n18848 );
nor  g16501 ( new_n18850 , new_n18841 , new_n18849 );
nor  g16502 ( new_n18851 , new_n18839 , new_n18850 );
nor  g16503 ( new_n18852 , new_n18838 , new_n18851 );
nor  g16504 ( new_n18853 , new_n18836 , new_n18852 );
nor  g16505 ( new_n18854 , new_n18835 , new_n18853 );
nor  g16506 ( new_n18855 , new_n18833 , new_n18854 );
nor  g16507 ( new_n18856 , new_n18832 , new_n18855 );
nor  g16508 ( new_n18857 , new_n18830_1 , new_n18856 );
nor  g16509 ( new_n18858_1 , new_n18829 , new_n18857 );
nor  g16510 ( new_n18859_1 , new_n18827 , new_n18858_1 );
nor  g16511 ( new_n18860 , new_n18826 , new_n18859_1 );
xnor g16512 ( n5980 , new_n18824 , new_n18860 );
xnor g16513 ( n6012 , new_n11120_1 , new_n11143 );
nor  g16514 ( new_n18863 , n16544 , new_n10095 );
xnor g16515 ( new_n18864_1 , n16544 , new_n10095 );
nor  g16516 ( new_n18865_1 , n6814 , new_n10058 );
xnor g16517 ( new_n18866 , n6814 , new_n10058 );
nor  g16518 ( new_n18867 , n19701 , new_n10063 );
xnor g16519 ( new_n18868 , n19701 , new_n10063 );
nor  g16520 ( new_n18869 , n23529 , new_n9249 );
and  g16521 ( new_n18870 , new_n9250 , new_n9286 );
nor  g16522 ( new_n18871 , new_n18869 , new_n18870 );
nor  g16523 ( new_n18872 , new_n18868 , new_n18871 );
nor  g16524 ( new_n18873 , new_n18867 , new_n18872 );
nor  g16525 ( new_n18874 , new_n18866 , new_n18873 );
nor  g16526 ( new_n18875 , new_n18865_1 , new_n18874 );
nor  g16527 ( new_n18876 , new_n18864_1 , new_n18875 );
nor  g16528 ( new_n18877 , new_n18863 , new_n18876 );
and  g16529 ( new_n18878 , new_n10044 , new_n18877 );
nor  g16530 ( new_n18879 , n3582 , new_n13823 );
xnor g16531 ( new_n18880_1 , n3582 , new_n13823 );
nor  g16532 ( new_n18881 , n2145 , new_n13859 );
xnor g16533 ( new_n18882 , n2145 , new_n13859 );
nor  g16534 ( new_n18883 , n5031 , new_n13829 );
xnor g16535 ( new_n18884 , n5031 , new_n13829 );
nor  g16536 ( new_n18885 , new_n7657_1 , new_n9311 );
nor  g16537 ( new_n18886_1 , new_n9313 , new_n9349 );
or   g16538 ( new_n18887_1 , new_n18885 , new_n18886_1 );
nor  g16539 ( new_n18888 , new_n18884 , new_n18887_1 );
nor  g16540 ( new_n18889 , new_n18883 , new_n18888 );
nor  g16541 ( new_n18890 , new_n18882 , new_n18889 );
nor  g16542 ( new_n18891 , new_n18881 , new_n18890 );
nor  g16543 ( new_n18892 , new_n18880_1 , new_n18891 );
nor  g16544 ( new_n18893 , new_n18879 , new_n18892 );
not  g16545 ( new_n18894 , new_n18893 );
nor  g16546 ( new_n18895 , new_n13869 , new_n18894 );
not  g16547 ( new_n18896 , new_n18895 );
xnor g16548 ( new_n18897 , new_n18878 , new_n18896 );
xnor g16549 ( new_n18898 , new_n10045 , new_n18877 );
xnor g16550 ( new_n18899 , new_n13868 , new_n18894 );
not  g16551 ( new_n18900 , new_n18899 );
nor  g16552 ( new_n18901_1 , new_n18898 , new_n18900 );
xnor g16553 ( new_n18902 , new_n18898 , new_n18900 );
xnor g16554 ( new_n18903 , new_n18864_1 , new_n18875 );
xor  g16555 ( new_n18904 , new_n18880_1 , new_n18891 );
nor  g16556 ( new_n18905 , new_n18903 , new_n18904 );
xnor g16557 ( new_n18906 , new_n18903 , new_n18904 );
xnor g16558 ( new_n18907_1 , new_n18866 , new_n18873 );
xor  g16559 ( new_n18908 , new_n18882 , new_n18889 );
nor  g16560 ( new_n18909 , new_n18907_1 , new_n18908 );
xnor g16561 ( new_n18910 , new_n18907_1 , new_n18908 );
xnor g16562 ( new_n18911 , new_n18868 , new_n18871 );
xor  g16563 ( new_n18912 , new_n18884 , new_n18887_1 );
nor  g16564 ( new_n18913 , new_n18911 , new_n18912 );
xnor g16565 ( new_n18914 , new_n18911 , new_n18912 );
and  g16566 ( new_n18915 , new_n9287_1 , new_n9351 );
nor  g16567 ( new_n18916 , new_n9352 , new_n9391 );
nor  g16568 ( new_n18917 , new_n18915 , new_n18916 );
nor  g16569 ( new_n18918 , new_n18914 , new_n18917 );
nor  g16570 ( new_n18919_1 , new_n18913 , new_n18918 );
nor  g16571 ( new_n18920 , new_n18910 , new_n18919_1 );
nor  g16572 ( new_n18921 , new_n18909 , new_n18920 );
nor  g16573 ( new_n18922 , new_n18906 , new_n18921 );
nor  g16574 ( new_n18923 , new_n18905 , new_n18922 );
nor  g16575 ( new_n18924 , new_n18902 , new_n18923 );
nor  g16576 ( new_n18925 , new_n18901_1 , new_n18924 );
xnor g16577 ( n6022 , new_n18897 , new_n18925 );
xnor g16578 ( n6031 , new_n18567 , new_n18584_1 );
not  g16579 ( new_n18928 , new_n8139_1 );
and  g16580 ( new_n18929 , new_n10873 , new_n16241 );
xnor g16581 ( new_n18930 , n17458 , new_n18929 );
xnor g16582 ( new_n18931 , new_n8719 , new_n18930 );
nor  g16583 ( new_n18932 , n15077 , new_n16242 );
and  g16584 ( new_n18933 , new_n16243_1 , new_n16279_1 );
nor  g16585 ( new_n18934 , new_n18932 , new_n18933 );
xnor g16586 ( new_n18935 , new_n18931 , new_n18934 );
xnor g16587 ( new_n18936 , n12702 , new_n18935 );
and  g16588 ( new_n18937 , new_n5611 , new_n16280 );
and  g16589 ( new_n18938 , new_n16281 , new_n16323 );
nor  g16590 ( new_n18939 , new_n18937 , new_n18938 );
xor  g16591 ( new_n18940_1 , new_n18936 , new_n18939 );
xnor g16592 ( new_n18941 , new_n18928 , new_n18940_1 );
nor  g16593 ( new_n18942 , new_n8144 , new_n16324 );
nor  g16594 ( new_n18943 , new_n16325 , new_n16363 );
nor  g16595 ( new_n18944 , new_n18942 , new_n18943 );
xnor g16596 ( n6044 , new_n18941 , new_n18944 );
and  g16597 ( new_n18946 , new_n9077 , new_n9119 );
and  g16598 ( new_n18947 , new_n9120 , new_n9177 );
nor  g16599 ( new_n18948 , new_n18946 , new_n18947 );
and  g16600 ( new_n18949 , new_n10679 , new_n9076 );
xnor g16601 ( new_n18950 , new_n18949 , new_n17629 );
xnor g16602 ( new_n18951 , new_n18948 , new_n18950 );
nor  g16603 ( new_n18952 , new_n4536 , new_n18951 );
xnor g16604 ( new_n18953 , new_n4536 , new_n18951 );
nor  g16605 ( new_n18954 , new_n9061 , new_n9178 );
nor  g16606 ( new_n18955 , new_n9179 , new_n9221 );
nor  g16607 ( new_n18956 , new_n18954 , new_n18955 );
nor  g16608 ( new_n18957 , new_n18953 , new_n18956 );
nor  g16609 ( new_n18958 , new_n18952 , new_n18957 );
not  g16610 ( new_n18959 , new_n18958 );
nor  g16611 ( new_n18960 , new_n18949 , new_n17629 );
and  g16612 ( new_n18961 , new_n18948 , new_n18960 );
and  g16613 ( new_n18962_1 , new_n4417 , new_n18961 );
and  g16614 ( new_n18963 , new_n18959 , new_n18962_1 );
or   g16615 ( new_n18964 , new_n4417 , new_n18961 );
nor  g16616 ( new_n18965 , new_n18959 , new_n18964 );
or   g16617 ( n6046 , new_n18963 , new_n18965 );
xnor g16618 ( new_n18967 , n7437 , n17077 );
nor  g16619 ( new_n18968 , new_n2893 , n26510 );
xnor g16620 ( new_n18969 , n20700 , n26510 );
nor  g16621 ( new_n18970_1 , new_n2896 , n23068 );
and  g16622 ( new_n18971 , new_n18646 , new_n18663 );
or   g16623 ( new_n18972 , new_n18970_1 , new_n18971 );
and  g16624 ( new_n18973 , new_n18969 , new_n18972 );
or   g16625 ( new_n18974 , new_n18968 , new_n18973 );
xor  g16626 ( new_n18975 , new_n18967 , new_n18974 );
xnor g16627 ( new_n18976 , new_n6970 , n21997 );
nor  g16628 ( new_n18977_1 , new_n6973 , new_n8501 );
or   g16629 ( new_n18978 , n21934 , n25119 );
nor  g16630 ( new_n18979 , n1163 , n18901 );
and  g16631 ( new_n18980 , new_n18618 , new_n18629 );
nor  g16632 ( new_n18981 , new_n18979 , new_n18980 );
and  g16633 ( new_n18982_1 , new_n18978 , new_n18981 );
nor  g16634 ( new_n18983 , new_n18977_1 , new_n18982_1 );
xor  g16635 ( new_n18984 , new_n18976 , new_n18983 );
xor  g16636 ( new_n18985 , new_n7479 , new_n18984 );
xnor g16637 ( new_n18986 , n21934 , n25119 );
xnor g16638 ( new_n18987 , new_n18981 , new_n18986 );
nor  g16639 ( new_n18988 , new_n2430 , new_n18987 );
nor  g16640 ( new_n18989 , new_n2423 , new_n18630 );
and  g16641 ( new_n18990 , new_n18631 , new_n18644 );
nor  g16642 ( new_n18991 , new_n18989 , new_n18990 );
xnor g16643 ( new_n18992 , new_n2431 , new_n18987 );
and  g16644 ( new_n18993 , new_n18991 , new_n18992 );
nor  g16645 ( new_n18994 , new_n18988 , new_n18993 );
xor  g16646 ( new_n18995 , new_n18985 , new_n18994 );
xnor g16647 ( new_n18996 , new_n18975 , new_n18995 );
not  g16648 ( new_n18997 , new_n18996 );
xor  g16649 ( new_n18998 , new_n18969 , new_n18972 );
xnor g16650 ( new_n18999_1 , new_n18991 , new_n18992 );
and  g16651 ( new_n19000 , new_n18998 , new_n18999_1 );
nor  g16652 ( new_n19001 , new_n18645 , new_n18664 );
and  g16653 ( new_n19002 , new_n18666 , new_n18695 );
nor  g16654 ( new_n19003 , new_n19001 , new_n19002 );
not  g16655 ( new_n19004 , new_n18999_1 );
xnor g16656 ( new_n19005_1 , new_n18998 , new_n19004 );
and  g16657 ( new_n19006 , new_n19003 , new_n19005_1 );
nor  g16658 ( new_n19007 , new_n19000 , new_n19006 );
xnor g16659 ( n6084 , new_n18997 , new_n19007 );
xnor g16660 ( n6160 , new_n10141 , new_n18775 );
xnor g16661 ( n6171 , new_n18779 , new_n18780_1 );
nor  g16662 ( new_n19011 , new_n7923 , n22359 );
and  g16663 ( new_n19012 , new_n9849 , new_n14865 );
or   g16664 ( new_n19013 , new_n19011 , new_n19012 );
xor  g16665 ( new_n19014 , new_n9852 , new_n19013 );
xnor g16666 ( new_n19015 , n21905 , n26264 );
not  g16667 ( new_n19016 , n7841 );
nor  g16668 ( new_n19017 , new_n19016 , n22918 );
xnor g16669 ( new_n19018 , n7841 , n22918 );
not  g16670 ( new_n19019 , n16812 );
nor  g16671 ( new_n19020 , new_n19019 , n25923 );
xnor g16672 ( new_n19021 , n16812 , n25923 );
not  g16673 ( new_n19022 , n25068 );
nor  g16674 ( new_n19023 , n6790 , new_n19022 );
and  g16675 ( new_n19024 , new_n17658 , new_n17678 );
or   g16676 ( new_n19025 , new_n19023 , new_n19024 );
and  g16677 ( new_n19026 , new_n19021 , new_n19025 );
or   g16678 ( new_n19027 , new_n19020 , new_n19026 );
and  g16679 ( new_n19028 , new_n19018 , new_n19027 );
or   g16680 ( new_n19029 , new_n19017 , new_n19028 );
xor  g16681 ( new_n19030 , new_n19015 , new_n19029 );
xnor g16682 ( new_n19031 , new_n15187 , new_n19030 );
xor  g16683 ( new_n19032 , new_n19018 , new_n19027 );
nor  g16684 ( new_n19033_1 , new_n15192 , new_n19032 );
xnor g16685 ( new_n19034 , new_n14932 , new_n19032 );
xor  g16686 ( new_n19035 , new_n19021 , new_n19025 );
and  g16687 ( new_n19036 , new_n14936 , new_n19035 );
xnor g16688 ( new_n19037 , new_n14935 , new_n19035 );
and  g16689 ( new_n19038 , new_n14941 , new_n17679 );
and  g16690 ( new_n19039 , new_n17680 , new_n17703 );
or   g16691 ( new_n19040 , new_n19038 , new_n19039 );
and  g16692 ( new_n19041 , new_n19037 , new_n19040 );
nor  g16693 ( new_n19042_1 , new_n19036 , new_n19041 );
and  g16694 ( new_n19043 , new_n19034 , new_n19042_1 );
nor  g16695 ( new_n19044_1 , new_n19033_1 , new_n19043 );
xor  g16696 ( new_n19045 , new_n19031 , new_n19044_1 );
xnor g16697 ( new_n19046 , new_n19014 , new_n19045 );
xnor g16698 ( new_n19047 , new_n19034 , new_n19042_1 );
nor  g16699 ( new_n19048 , new_n14866 , new_n19047 );
xnor g16700 ( new_n19049 , new_n14866 , new_n19047 );
xor  g16701 ( new_n19050 , new_n19037 , new_n19040 );
nor  g16702 ( new_n19051 , new_n14868 , new_n19050 );
xnor g16703 ( new_n19052 , new_n14868 , new_n19050 );
nor  g16704 ( new_n19053 , new_n14871 , new_n17704 );
nor  g16705 ( new_n19054 , new_n17705 , new_n17729 );
nor  g16706 ( new_n19055 , new_n19053 , new_n19054 );
nor  g16707 ( new_n19056 , new_n19052 , new_n19055 );
nor  g16708 ( new_n19057 , new_n19051 , new_n19056 );
nor  g16709 ( new_n19058 , new_n19049 , new_n19057 );
nor  g16710 ( new_n19059 , new_n19048 , new_n19058 );
xnor g16711 ( n6183 , new_n19046 , new_n19059 );
xnor g16712 ( new_n19061 , n14345 , n14702 );
nor  g16713 ( new_n19062 , n2999 , new_n9088 );
xnor g16714 ( new_n19063 , n2999 , n11356 );
nor  g16715 ( new_n19064 , n2547 , new_n9091 );
xnor g16716 ( new_n19065 , n2547 , n3164 );
nor  g16717 ( new_n19066 , new_n10623 , n10611 );
and  g16718 ( new_n19067 , new_n13783_1 , new_n13792 );
nor  g16719 ( new_n19068 , new_n19066 , new_n19067 );
and  g16720 ( new_n19069 , new_n19065 , new_n19068 );
or   g16721 ( new_n19070 , new_n19064 , new_n19069 );
and  g16722 ( new_n19071 , new_n19063 , new_n19070 );
or   g16723 ( new_n19072 , new_n19062 , new_n19071 );
xor  g16724 ( new_n19073 , new_n19061 , new_n19072 );
xor  g16725 ( new_n19074 , new_n9011 , new_n19073 );
xor  g16726 ( new_n19075 , new_n19063 , new_n19070 );
nor  g16727 ( new_n19076 , new_n9015 , new_n19075 );
xnor g16728 ( new_n19077 , new_n9015 , new_n19075 );
not  g16729 ( new_n19078 , new_n9019 );
xnor g16730 ( new_n19079 , new_n19065 , new_n19068 );
and  g16731 ( new_n19080 , new_n19078 , new_n19079 );
xnor g16732 ( new_n19081_1 , new_n19078 , new_n19079 );
and  g16733 ( new_n19082 , new_n9023 , new_n13793 );
nor  g16734 ( new_n19083 , new_n13794 , new_n13808 );
nor  g16735 ( new_n19084 , new_n19082 , new_n19083 );
nor  g16736 ( new_n19085 , new_n19081_1 , new_n19084 );
nor  g16737 ( new_n19086 , new_n19080 , new_n19085 );
nor  g16738 ( new_n19087 , new_n19077 , new_n19086 );
nor  g16739 ( new_n19088 , new_n19076 , new_n19087 );
xor  g16740 ( n6189 , new_n19074 , new_n19088 );
xnor g16741 ( new_n19090 , n15167 , n20036 );
nor  g16742 ( new_n19091 , n11192 , new_n12134 );
or   g16743 ( new_n19092 , new_n4120 , n21095 );
nor  g16744 ( new_n19093 , new_n6492 , n9380 );
and  g16745 ( new_n19094 , new_n19092 , new_n19093 );
or   g16746 ( new_n19095 , new_n19091 , new_n19094 );
xor  g16747 ( new_n19096 , new_n19090 , new_n19095 );
xnor g16748 ( new_n19097 , new_n17713 , new_n19096 );
xnor g16749 ( new_n19098 , n8656 , n9380 );
nor  g16750 ( new_n19099 , new_n17717 , new_n19098 );
xnor g16751 ( new_n19100 , n11192 , n21095 );
xnor g16752 ( new_n19101 , new_n19093 , new_n19100 );
nor  g16753 ( new_n19102 , new_n19099 , new_n19101 );
xnor g16754 ( new_n19103 , new_n19099 , new_n19101 );
nor  g16755 ( new_n19104 , new_n17721_1 , new_n19103 );
nor  g16756 ( new_n19105 , new_n19102 , new_n19104 );
xnor g16757 ( n6223 , new_n19097 , new_n19105 );
xnor g16758 ( n6233 , new_n13798_1 , new_n13806 );
xnor g16759 ( n6245 , new_n18308 , new_n18311_1 );
xnor g16760 ( n6248 , new_n10133 , new_n10145 );
xnor g16761 ( new_n19110 , n16544 , n21839 );
nor  g16762 ( new_n19111 , new_n2887_1 , n27089 );
and  g16763 ( new_n19112 , new_n18719 , new_n18749 );
or   g16764 ( new_n19113 , new_n19111 , new_n19112 );
xor  g16765 ( new_n19114 , new_n19110 , new_n19113 );
xnor g16766 ( new_n19115 , new_n10102 , new_n19114 );
nor  g16767 ( new_n19116_1 , new_n10106 , new_n18750 );
nor  g16768 ( new_n19117 , new_n18751_1 , new_n18791 );
nor  g16769 ( new_n19118 , new_n19116_1 , new_n19117 );
xnor g16770 ( n6256 , new_n19115 , new_n19118 );
xnor g16771 ( n6271 , new_n14605 , new_n14620 );
nor  g16772 ( new_n19121 , n13549 , new_n7918 );
not  g16773 ( new_n19122 , n23493 );
nor  g16774 ( new_n19123 , n8405 , new_n19122 );
and  g16775 ( new_n19124 , new_n9852 , new_n19013 );
or   g16776 ( new_n19125_1 , new_n19123 , new_n19124 );
and  g16777 ( new_n19126 , new_n9855 , new_n19125_1 );
nor  g16778 ( new_n19127 , new_n19121 , new_n19126 );
nor  g16779 ( new_n19128 , new_n2674 , n13951 );
xnor g16780 ( new_n19129 , n2944 , n13951 );
nor  g16781 ( new_n19130 , new_n2677 , n22793 );
or   g16782 ( new_n19131 , new_n14631 , new_n14650 );
and  g16783 ( new_n19132 , new_n14629 , new_n19131 );
or   g16784 ( new_n19133 , new_n19130 , new_n19132 );
and  g16785 ( new_n19134 , new_n19129 , new_n19133 );
nor  g16786 ( new_n19135 , new_n19128 , new_n19134 );
and  g16787 ( new_n19136 , new_n19127 , new_n19135 );
nor  g16788 ( new_n19137 , new_n19130 , new_n19132 );
xnor g16789 ( new_n19138 , new_n19129 , new_n19137 );
xor  g16790 ( new_n19139 , new_n9855 , new_n19125_1 );
nor  g16791 ( new_n19140 , new_n19138 , new_n19139 );
not  g16792 ( new_n19141_1 , new_n19138 );
xnor g16793 ( new_n19142 , new_n19141_1 , new_n19139 );
and  g16794 ( new_n19143 , new_n14652 , new_n19014 );
xnor g16795 ( new_n19144_1 , new_n14653 , new_n19014 );
nor  g16796 ( new_n19145 , new_n14655 , new_n14866 );
nor  g16797 ( new_n19146 , new_n14867 , new_n14885 );
nor  g16798 ( new_n19147 , new_n19145 , new_n19146 );
and  g16799 ( new_n19148 , new_n19144_1 , new_n19147 );
nor  g16800 ( new_n19149 , new_n19143 , new_n19148 );
and  g16801 ( new_n19150 , new_n19142 , new_n19149 );
nor  g16802 ( new_n19151 , new_n19140 , new_n19150 );
xnor g16803 ( new_n19152 , new_n19127 , new_n19135 );
nor  g16804 ( new_n19153 , new_n19151 , new_n19152 );
nor  g16805 ( new_n19154 , new_n19136 , new_n19153 );
not  g16806 ( new_n19155 , new_n19154 );
nor  g16807 ( new_n19156 , n1881 , new_n14547_1 );
xnor g16808 ( new_n19157 , n1881 , n8827 );
nor  g16809 ( new_n19158 , n5834 , new_n12683 );
and  g16810 ( new_n19159 , new_n18556 , new_n18559 );
or   g16811 ( new_n19160 , new_n19158 , new_n19159 );
and  g16812 ( new_n19161 , new_n19157 , new_n19160 );
nor  g16813 ( new_n19162 , new_n19156 , new_n19161 );
not  g16814 ( new_n19163_1 , new_n19162 );
xnor g16815 ( new_n19164_1 , new_n19155 , new_n19163_1 );
xnor g16816 ( new_n19165 , new_n19151 , new_n19152 );
nor  g16817 ( new_n19166 , new_n19162 , new_n19165 );
not  g16818 ( new_n19167 , new_n19165 );
xnor g16819 ( new_n19168 , new_n19162 , new_n19167 );
xor  g16820 ( new_n19169 , new_n19157 , new_n19160 );
xnor g16821 ( new_n19170 , new_n19142 , new_n19149 );
and  g16822 ( new_n19171 , new_n19169 , new_n19170 );
xnor g16823 ( new_n19172 , new_n19144_1 , new_n19147 );
not  g16824 ( new_n19173 , new_n19172 );
nor  g16825 ( new_n19174_1 , new_n18560 , new_n19173 );
xnor g16826 ( new_n19175 , new_n18560 , new_n19172 );
and  g16827 ( new_n19176_1 , new_n14886 , new_n15139_1 );
and  g16828 ( new_n19177 , new_n15140 , new_n15159 );
nor  g16829 ( new_n19178 , new_n19176_1 , new_n19177 );
and  g16830 ( new_n19179 , new_n19175 , new_n19178 );
nor  g16831 ( new_n19180 , new_n19174_1 , new_n19179 );
not  g16832 ( new_n19181 , new_n19170 );
xnor g16833 ( new_n19182 , new_n19169 , new_n19181 );
and  g16834 ( new_n19183 , new_n19180 , new_n19182 );
nor  g16835 ( new_n19184 , new_n19171 , new_n19183 );
and  g16836 ( new_n19185 , new_n19168 , new_n19184 );
nor  g16837 ( new_n19186 , new_n19166 , new_n19185 );
xor  g16838 ( n6276 , new_n19164_1 , new_n19186 );
xnor g16839 ( n6308 , new_n18267 , new_n18268 );
xnor g16840 ( n6311 , new_n16436 , new_n16450 );
xnor g16841 ( n6323 , new_n16203 , new_n16217_1 );
nor  g16842 ( new_n19191 , new_n13508 , new_n5915 );
and  g16843 ( new_n19192 , new_n5916 , new_n5979 );
nor  g16844 ( new_n19193 , new_n19191 , new_n19192 );
not  g16845 ( new_n19194 , new_n19193 );
and  g16846 ( new_n19195 , new_n13550 , new_n13194 );
and  g16847 ( new_n19196_1 , new_n19194 , new_n19195 );
or   g16848 ( new_n19197 , new_n13550 , new_n13194 );
nor  g16849 ( new_n19198 , new_n19194 , new_n19197 );
nor  g16850 ( new_n19199 , new_n19196_1 , new_n19198 );
nor  g16851 ( new_n19200 , new_n17497 , new_n19199 );
xnor g16852 ( new_n19201 , new_n17497 , new_n19199 );
xnor g16853 ( new_n19202_1 , new_n13550 , new_n13193 );
xnor g16854 ( new_n19203 , new_n19194 , new_n19202_1 );
nor  g16855 ( new_n19204 , new_n17500_1 , new_n19203 );
xnor g16856 ( new_n19205 , new_n17500_1 , new_n19203 );
nor  g16857 ( new_n19206 , new_n5980_1 , new_n6088 );
nor  g16858 ( new_n19207 , new_n6089 , new_n6149 );
nor  g16859 ( new_n19208 , new_n19206 , new_n19207 );
nor  g16860 ( new_n19209 , new_n19205 , new_n19208 );
nor  g16861 ( new_n19210 , new_n19204 , new_n19209 );
nor  g16862 ( new_n19211 , new_n19201 , new_n19210 );
nor  g16863 ( new_n19212 , new_n19200 , new_n19211 );
nor  g16864 ( n6330 , new_n19196_1 , new_n19212 );
xnor g16865 ( n6339 , new_n8534 , new_n8568 );
xnor g16866 ( n6354 , new_n13749 , new_n13775_1 );
or   g16867 ( new_n19216 , n7335 , new_n3213 );
nor  g16868 ( new_n19217 , n5696 , new_n3220 );
xnor g16869 ( new_n19218 , n5696 , new_n3221 );
nor  g16870 ( new_n19219 , n13367 , new_n3226 );
xnor g16871 ( new_n19220_1 , n13367 , new_n3227 );
nor  g16872 ( new_n19221_1 , n932 , new_n3231 );
xnor g16873 ( new_n19222 , n932 , new_n3232 );
nor  g16874 ( new_n19223_1 , n6691 , new_n3236 );
xnor g16875 ( new_n19224_1 , n6691 , new_n3237 );
nor  g16876 ( new_n19225 , n3260 , new_n3241 );
xnor g16877 ( new_n19226 , n3260 , new_n3242 );
nor  g16878 ( new_n19227 , n20489 , new_n3246 );
nor  g16879 ( new_n19228_1 , n2355 , new_n3251 );
xnor g16880 ( new_n19229 , n2355 , new_n3252 );
nor  g16881 ( new_n19230 , n11121 , new_n3262 );
or   g16882 ( new_n19231 , new_n2448 , new_n3117 );
xor  g16883 ( new_n19232 , n11121 , new_n3262 );
and  g16884 ( new_n19233_1 , new_n19231 , new_n19232 );
or   g16885 ( new_n19234_1 , new_n19230 , new_n19233_1 );
and  g16886 ( new_n19235 , new_n19229 , new_n19234_1 );
or   g16887 ( new_n19236 , new_n19228_1 , new_n19235 );
xnor g16888 ( new_n19237 , n20489 , new_n3247 );
and  g16889 ( new_n19238 , new_n19236 , new_n19237 );
or   g16890 ( new_n19239 , new_n19227 , new_n19238 );
and  g16891 ( new_n19240 , new_n19226 , new_n19239 );
or   g16892 ( new_n19241 , new_n19225 , new_n19240 );
and  g16893 ( new_n19242 , new_n19224_1 , new_n19241 );
or   g16894 ( new_n19243 , new_n19223_1 , new_n19242 );
and  g16895 ( new_n19244_1 , new_n19222 , new_n19243 );
or   g16896 ( new_n19245 , new_n19221_1 , new_n19244_1 );
and  g16897 ( new_n19246 , new_n19220_1 , new_n19245 );
or   g16898 ( new_n19247 , new_n19219 , new_n19246 );
and  g16899 ( new_n19248 , new_n19218 , new_n19247 );
nor  g16900 ( new_n19249 , new_n19217 , new_n19248 );
and  g16901 ( new_n19250 , new_n19216 , new_n19249 );
and  g16902 ( new_n19251 , n7335 , new_n3213 );
or   g16903 ( new_n19252 , new_n3218 , new_n19251 );
nor  g16904 ( new_n19253 , new_n19250 , new_n19252 );
and  g16905 ( new_n19254 , new_n16628 , new_n19253 );
nor  g16906 ( new_n19255 , new_n16668 , new_n19253 );
xnor g16907 ( new_n19256 , new_n16668 , new_n19253 );
xnor g16908 ( new_n19257 , n7335 , new_n3214 );
xnor g16909 ( new_n19258 , new_n19249 , new_n19257 );
and  g16910 ( new_n19259 , new_n16671 , new_n19258 );
xnor g16911 ( new_n19260 , new_n16671 , new_n19258 );
xor  g16912 ( new_n19261 , new_n19218 , new_n19247 );
and  g16913 ( new_n19262 , new_n16677 , new_n19261 );
xnor g16914 ( new_n19263 , new_n16677 , new_n19261 );
not  g16915 ( new_n19264 , new_n16681 );
xor  g16916 ( new_n19265 , new_n19220_1 , new_n19245 );
and  g16917 ( new_n19266 , new_n19264 , new_n19265 );
xnor g16918 ( new_n19267 , new_n19264 , new_n19265 );
xor  g16919 ( new_n19268 , new_n19222 , new_n19243 );
and  g16920 ( new_n19269 , new_n16685 , new_n19268 );
xnor g16921 ( new_n19270_1 , new_n16685 , new_n19268 );
xor  g16922 ( new_n19271 , new_n19224_1 , new_n19241 );
and  g16923 ( new_n19272 , new_n16690 , new_n19271 );
xnor g16924 ( new_n19273 , new_n16690 , new_n19271 );
xor  g16925 ( new_n19274 , new_n19226 , new_n19239 );
and  g16926 ( new_n19275 , new_n16695 , new_n19274 );
xnor g16927 ( new_n19276 , new_n16695 , new_n19274 );
xor  g16928 ( new_n19277 , new_n19236 , new_n19237 );
and  g16929 ( new_n19278 , new_n16698 , new_n19277 );
xnor g16930 ( new_n19279 , new_n16701 , new_n19277 );
xor  g16931 ( new_n19280 , new_n19229 , new_n19234_1 );
nor  g16932 ( new_n19281 , new_n16704 , new_n19280 );
xor  g16933 ( new_n19282_1 , new_n16704 , new_n19280 );
nor  g16934 ( new_n19283 , new_n16709 , new_n19232 );
xor  g16935 ( new_n19284 , new_n19231 , new_n19232 );
nor  g16936 ( new_n19285 , new_n16708 , new_n19284 );
xnor g16937 ( new_n19286 , n12315 , n16217 );
nor  g16938 ( new_n19287 , new_n16715 , new_n19286 );
nor  g16939 ( new_n19288 , new_n19285 , new_n19287 );
nor  g16940 ( new_n19289 , new_n19283 , new_n19288 );
and  g16941 ( new_n19290 , new_n19282_1 , new_n19289 );
nor  g16942 ( new_n19291 , new_n19281 , new_n19290 );
and  g16943 ( new_n19292 , new_n19279 , new_n19291 );
nor  g16944 ( new_n19293 , new_n19278 , new_n19292 );
nor  g16945 ( new_n19294 , new_n19276 , new_n19293 );
nor  g16946 ( new_n19295 , new_n19275 , new_n19294 );
nor  g16947 ( new_n19296 , new_n19273 , new_n19295 );
nor  g16948 ( new_n19297 , new_n19272 , new_n19296 );
nor  g16949 ( new_n19298 , new_n19270_1 , new_n19297 );
nor  g16950 ( new_n19299 , new_n19269 , new_n19298 );
nor  g16951 ( new_n19300 , new_n19267 , new_n19299 );
nor  g16952 ( new_n19301 , new_n19266 , new_n19300 );
nor  g16953 ( new_n19302 , new_n19263 , new_n19301 );
nor  g16954 ( new_n19303 , new_n19262 , new_n19302 );
nor  g16955 ( new_n19304 , new_n19260 , new_n19303 );
nor  g16956 ( new_n19305 , new_n19259 , new_n19304 );
nor  g16957 ( new_n19306 , new_n19256 , new_n19305 );
nor  g16958 ( new_n19307 , new_n19255 , new_n19306 );
nor  g16959 ( new_n19308 , new_n19254 , new_n19307 );
nor  g16960 ( new_n19309 , new_n16628 , new_n19253 );
nor  g16961 ( new_n19310 , new_n19306 , new_n19309 );
nor  g16962 ( n6375 , new_n19308 , new_n19310 );
xnor g16963 ( n6383 , new_n18420 , new_n18434 );
xnor g16964 ( n6407 , new_n14118 , new_n14158 );
xnor g16965 ( n6431 , new_n8559 , new_n8560 );
xnor g16966 ( n6437 , new_n16059 , new_n16062_1 );
xnor g16967 ( n6457 , new_n4159 , new_n4161 );
xnor g16968 ( n6465 , new_n12070 , new_n12099 );
not  g16969 ( new_n19318 , new_n8339_1 );
and  g16970 ( new_n19319 , n3740 , new_n16930 );
and  g16971 ( new_n19320 , new_n5982 , new_n16929 );
nor  g16972 ( new_n19321 , n3740 , new_n16930 );
nor  g16973 ( new_n19322 , new_n19321 , new_n16935 );
or   g16974 ( new_n19323_1 , new_n19320 , new_n19322 );
nor  g16975 ( new_n19324 , new_n19319 , new_n19323_1 );
not  g16976 ( new_n19325 , new_n19324 );
xnor g16977 ( new_n19326 , new_n19318 , new_n19325 );
not  g16978 ( new_n19327_1 , new_n3472 );
nor  g16979 ( new_n19328 , new_n19327_1 , new_n17928 );
xnor g16980 ( new_n19329 , new_n19327_1 , new_n16936 );
nor  g16981 ( new_n19330 , new_n3476 , new_n17930 );
and  g16982 ( new_n19331 , new_n14033 , new_n14073 );
nor  g16983 ( new_n19332 , new_n19330 , new_n19331 );
and  g16984 ( new_n19333_1 , new_n19329 , new_n19332 );
nor  g16985 ( new_n19334 , new_n19328 , new_n19333_1 );
xnor g16986 ( new_n19335 , new_n19326 , new_n19334 );
not  g16987 ( new_n19336 , new_n19335 );
nor  g16988 ( new_n19337 , n2743 , new_n3598 );
nor  g16989 ( new_n19338 , new_n3537 , new_n3603 );
nor  g16990 ( new_n19339 , n7026 , new_n3602 );
nor  g16991 ( new_n19340 , new_n19339 , new_n14105 );
nor  g16992 ( new_n19341 , new_n19338 , new_n19340 );
nor  g16993 ( new_n19342 , new_n19337 , new_n19341 );
and  g16994 ( new_n19343 , new_n4797 , new_n3597 );
not  g16995 ( new_n19344 , new_n3598 );
nor  g16996 ( new_n19345 , new_n13254 , new_n19344 );
or   g16997 ( new_n19346 , new_n19343 , new_n19345 );
nor  g16998 ( new_n19347 , new_n19342 , new_n19346 );
xnor g16999 ( new_n19348_1 , new_n19336 , new_n19347 );
xnor g17000 ( new_n19349 , new_n19329 , new_n19332 );
not  g17001 ( new_n19350 , new_n19349 );
xnor g17002 ( new_n19351 , n2743 , new_n19344 );
xnor g17003 ( new_n19352 , new_n19341 , new_n19351 );
nor  g17004 ( new_n19353 , new_n19350 , new_n19352 );
xnor g17005 ( new_n19354_1 , new_n19350 , new_n19352 );
nor  g17006 ( new_n19355 , new_n14074 , new_n14106 );
and  g17007 ( new_n19356 , new_n14107_1 , new_n14162 );
nor  g17008 ( new_n19357_1 , new_n19355 , new_n19356 );
nor  g17009 ( new_n19358 , new_n19354_1 , new_n19357_1 );
nor  g17010 ( new_n19359 , new_n19353 , new_n19358 );
xnor g17011 ( n6470 , new_n19348_1 , new_n19359 );
xnor g17012 ( n6476 , new_n11387 , new_n11409 );
xnor g17013 ( n6506 , new_n17960 , new_n17968_1 );
nor  g17014 ( new_n19363 , new_n9332 , new_n9334 );
not  g17015 ( new_n19364 , new_n19363 );
nor  g17016 ( new_n19365 , new_n9340 , new_n19364 );
not  g17017 ( new_n19366 , new_n19365 );
nor  g17018 ( new_n19367_1 , new_n9327 , new_n19366 );
not  g17019 ( new_n19368 , new_n19367_1 );
nor  g17020 ( new_n19369 , new_n9322 , new_n19368 );
not  g17021 ( new_n19370 , new_n19369 );
nor  g17022 ( new_n19371 , new_n9317 , new_n19370 );
not  g17023 ( new_n19372 , new_n19371 );
nor  g17024 ( new_n19373 , new_n9312 , new_n19372 );
not  g17025 ( new_n19374 , new_n19373 );
nor  g17026 ( new_n19375 , new_n13829 , new_n19374 );
xnor g17027 ( new_n19376 , new_n13859 , new_n19375 );
xnor g17028 ( new_n19377 , new_n10057_1 , new_n19376 );
xnor g17029 ( new_n19378 , new_n13829 , new_n19373 );
nor  g17030 ( new_n19379 , new_n10063 , new_n19378 );
xnor g17031 ( new_n19380 , new_n10063 , new_n19378 );
xnor g17032 ( new_n19381 , new_n9312 , new_n19371 );
nor  g17033 ( new_n19382 , new_n9249 , new_n19381 );
xnor g17034 ( new_n19383 , new_n9249 , new_n19381 );
xnor g17035 ( new_n19384 , new_n9317 , new_n19369 );
nor  g17036 ( new_n19385_1 , new_n9251_1 , new_n19384 );
xnor g17037 ( new_n19386 , new_n9251_1 , new_n19384 );
xnor g17038 ( new_n19387 , new_n9322 , new_n19367_1 );
nor  g17039 ( new_n19388 , new_n9256 , new_n19387 );
xnor g17040 ( new_n19389_1 , new_n9255 , new_n19387 );
xnor g17041 ( new_n19390 , new_n9327 , new_n19365 );
nor  g17042 ( new_n19391 , new_n9261_1 , new_n19390 );
xnor g17043 ( new_n19392 , new_n9340 , new_n19363 );
nor  g17044 ( new_n19393 , new_n9266 , new_n19392 );
xnor g17045 ( new_n19394 , new_n9265 , new_n19392 );
nor  g17046 ( new_n19395 , new_n9272 , new_n9335 );
nor  g17047 ( new_n19396 , new_n9274 , new_n19395 );
nor  g17048 ( new_n19397 , new_n9300 , new_n9335 );
or   g17049 ( new_n19398 , new_n19363 , new_n19397 );
and  g17050 ( new_n19399 , new_n9237 , new_n19395 );
nor  g17051 ( new_n19400 , new_n19396 , new_n19399 );
and  g17052 ( new_n19401_1 , new_n19398 , new_n19400 );
or   g17053 ( new_n19402 , new_n19396 , new_n19401_1 );
and  g17054 ( new_n19403 , new_n19394 , new_n19402 );
or   g17055 ( new_n19404 , new_n19393 , new_n19403 );
xnor g17056 ( new_n19405 , new_n9260 , new_n19390 );
and  g17057 ( new_n19406 , new_n19404 , new_n19405 );
or   g17058 ( new_n19407 , new_n19391 , new_n19406 );
and  g17059 ( new_n19408 , new_n19389_1 , new_n19407 );
nor  g17060 ( new_n19409 , new_n19388 , new_n19408 );
nor  g17061 ( new_n19410 , new_n19386 , new_n19409 );
nor  g17062 ( new_n19411 , new_n19385_1 , new_n19410 );
nor  g17063 ( new_n19412 , new_n19383 , new_n19411 );
nor  g17064 ( new_n19413 , new_n19382 , new_n19412 );
nor  g17065 ( new_n19414_1 , new_n19380 , new_n19413 );
or   g17066 ( new_n19415 , new_n19379 , new_n19414_1 );
xor  g17067 ( new_n19416 , new_n19377 , new_n19415 );
xor  g17068 ( new_n19417 , new_n16280 , new_n19416 );
xnor g17069 ( new_n19418 , new_n19380 , new_n19413 );
nor  g17070 ( new_n19419 , new_n16282 , new_n19418 );
xnor g17071 ( new_n19420 , new_n16282 , new_n19418 );
xnor g17072 ( new_n19421 , new_n19383 , new_n19411 );
nor  g17073 ( new_n19422 , new_n16289 , new_n19421 );
xnor g17074 ( new_n19423 , new_n16289 , new_n19421 );
xnor g17075 ( new_n19424_1 , new_n19386 , new_n19409 );
nor  g17076 ( new_n19425 , new_n16294 , new_n19424_1 );
xnor g17077 ( new_n19426 , new_n16292 , new_n19424_1 );
xor  g17078 ( new_n19427 , new_n19389_1 , new_n19407 );
nor  g17079 ( new_n19428 , new_n16296 , new_n19427 );
xor  g17080 ( new_n19429 , new_n19404 , new_n19405 );
nor  g17081 ( new_n19430 , new_n16299 , new_n19429 );
xnor g17082 ( new_n19431 , new_n16299 , new_n19429 );
xor  g17083 ( new_n19432 , new_n19394 , new_n19402 );
nor  g17084 ( new_n19433 , new_n16302 , new_n19432 );
xnor g17085 ( new_n19434 , new_n16302 , new_n19432 );
xor  g17086 ( new_n19435 , new_n19398 , new_n19400 );
nor  g17087 ( new_n19436 , new_n16305 , new_n19435 );
xnor g17088 ( new_n19437 , new_n6628_1 , n13714 );
xnor g17089 ( new_n19438 , new_n9272 , new_n9334 );
and  g17090 ( new_n19439 , new_n19437 , new_n19438 );
xor  g17091 ( new_n19440 , new_n16305 , new_n19435 );
and  g17092 ( new_n19441 , new_n19439 , new_n19440 );
nor  g17093 ( new_n19442 , new_n19436 , new_n19441 );
nor  g17094 ( new_n19443 , new_n19434 , new_n19442 );
nor  g17095 ( new_n19444 , new_n19433 , new_n19443 );
nor  g17096 ( new_n19445 , new_n19431 , new_n19444 );
nor  g17097 ( new_n19446 , new_n19430 , new_n19445 );
xnor g17098 ( new_n19447 , new_n16296 , new_n19427 );
nor  g17099 ( new_n19448 , new_n19446 , new_n19447 );
nor  g17100 ( new_n19449 , new_n19428 , new_n19448 );
and  g17101 ( new_n19450_1 , new_n19426 , new_n19449 );
nor  g17102 ( new_n19451 , new_n19425 , new_n19450_1 );
nor  g17103 ( new_n19452 , new_n19423 , new_n19451 );
nor  g17104 ( new_n19453 , new_n19422 , new_n19452 );
nor  g17105 ( new_n19454_1 , new_n19420 , new_n19453 );
nor  g17106 ( new_n19455 , new_n19419 , new_n19454_1 );
xor  g17107 ( n6514 , new_n19417 , new_n19455 );
and  g17108 ( new_n19457 , new_n11288 , new_n11376 );
nor  g17109 ( new_n19458_1 , new_n11377 , new_n11413 );
nor  g17110 ( new_n19459 , new_n19457 , new_n19458_1 );
not  g17111 ( new_n19460 , new_n19459 );
xnor g17112 ( new_n19461 , new_n11794 , new_n11336 );
and  g17113 ( new_n19462 , new_n11375_1 , new_n19461 );
nor  g17114 ( new_n19463 , new_n11850 , new_n11336 );
or   g17115 ( new_n19464 , new_n19463 , new_n11375_1 );
nor  g17116 ( new_n19465 , new_n19461 , new_n19464 );
nor  g17117 ( new_n19466 , new_n19462 , new_n19465 );
xnor g17118 ( n6542 , new_n19460 , new_n19466 );
xnor g17119 ( n6558 , new_n15027 , new_n15040 );
xnor g17120 ( n6560 , new_n17479 , new_n17481 );
xnor g17121 ( new_n19470 , new_n4021 , new_n6277 );
nor  g17122 ( new_n19471 , new_n4106 , new_n6280 );
xnor g17123 ( new_n19472_1 , new_n4106 , new_n6282 );
nor  g17124 ( new_n19473 , n17090 , new_n12226 );
or   g17125 ( new_n19474 , new_n4030 , new_n6288 );
xnor g17126 ( new_n19475 , new_n4111 , new_n12226 );
and  g17127 ( new_n19476 , new_n19474 , new_n19475 );
nor  g17128 ( new_n19477_1 , new_n19473 , new_n19476 );
and  g17129 ( new_n19478 , new_n19472_1 , new_n19477_1 );
or   g17130 ( new_n19479 , new_n19471 , new_n19478 );
xor  g17131 ( new_n19480 , new_n19470 , new_n19479 );
xnor g17132 ( new_n19481 , new_n9673 , new_n19480 );
xor  g17133 ( new_n19482 , new_n19472_1 , new_n19477_1 );
nor  g17134 ( new_n19483 , new_n9678 , new_n19482 );
xnor g17135 ( new_n19484 , new_n9678 , new_n19482 );
xor  g17136 ( new_n19485 , new_n19474 , new_n19475 );
and  g17137 ( new_n19486 , new_n9683 , new_n19485 );
nor  g17138 ( new_n19487 , new_n9686 , new_n17509 );
xnor g17139 ( new_n19488 , new_n10808 , new_n19485 );
and  g17140 ( new_n19489 , new_n19487 , new_n19488 );
nor  g17141 ( new_n19490 , new_n19486 , new_n19489 );
nor  g17142 ( new_n19491 , new_n19484 , new_n19490 );
nor  g17143 ( new_n19492 , new_n19483 , new_n19491 );
xnor g17144 ( n6567 , new_n19481 , new_n19492 );
not  g17145 ( new_n19494_1 , new_n13408 );
nor  g17146 ( new_n19495 , n8324 , new_n19494_1 );
not  g17147 ( new_n19496_1 , new_n19495 );
nor  g17148 ( new_n19497 , n1279 , new_n19496_1 );
not  g17149 ( new_n19498 , new_n19497 );
nor  g17150 ( new_n19499 , n9445 , new_n19498 );
not  g17151 ( new_n19500 , new_n19499 );
nor  g17152 ( new_n19501 , n19454 , new_n19500 );
xnor g17153 ( new_n19502 , n1536 , new_n19501 );
xnor g17154 ( new_n19503 , new_n4473 , new_n19502 );
xnor g17155 ( new_n19504 , n19454 , new_n19499 );
nor  g17156 ( new_n19505 , new_n4482 , new_n19504 );
xnor g17157 ( new_n19506 , new_n4481 , new_n19504 );
xnor g17158 ( new_n19507 , n9445 , new_n19497 );
nor  g17159 ( new_n19508 , new_n4488 , new_n19507 );
xnor g17160 ( new_n19509 , new_n4487 , new_n19507 );
xnor g17161 ( new_n19510 , n1279 , new_n19495 );
nor  g17162 ( new_n19511 , new_n4493 , new_n19510 );
xnor g17163 ( new_n19512 , new_n4493 , new_n19510 );
nor  g17164 ( new_n19513 , new_n3963 , new_n13409_1 );
nor  g17165 ( new_n19514_1 , new_n13410 , new_n13431 );
nor  g17166 ( new_n19515_1 , new_n19513 , new_n19514_1 );
nor  g17167 ( new_n19516 , new_n19512 , new_n19515_1 );
or   g17168 ( new_n19517 , new_n19511 , new_n19516 );
and  g17169 ( new_n19518 , new_n19509 , new_n19517 );
or   g17170 ( new_n19519 , new_n19508 , new_n19518 );
and  g17171 ( new_n19520 , new_n19506 , new_n19519 );
nor  g17172 ( new_n19521 , new_n19505 , new_n19520 );
xnor g17173 ( new_n19522 , new_n19503 , new_n19521 );
not  g17174 ( new_n19523_1 , new_n19522 );
xnor g17175 ( new_n19524 , n23272 , new_n8079 );
nor  g17176 ( new_n19525 , n11481 , new_n8081 );
xnor g17177 ( new_n19526 , new_n4361 , new_n8081 );
nor  g17178 ( new_n19527 , n16439 , new_n8084 );
xnor g17179 ( new_n19528 , new_n4365 , new_n8084 );
nor  g17180 ( new_n19529 , n15241 , new_n8087 );
nor  g17181 ( new_n19530 , new_n4373 , new_n8093 );
and  g17182 ( new_n19531_1 , new_n13433 , new_n13450 );
nor  g17183 ( new_n19532 , new_n19530 , new_n19531_1 );
xnor g17184 ( new_n19533 , new_n4369 , new_n8087 );
and  g17185 ( new_n19534 , new_n19532 , new_n19533 );
or   g17186 ( new_n19535 , new_n19529 , new_n19534 );
and  g17187 ( new_n19536 , new_n19528 , new_n19535 );
or   g17188 ( new_n19537 , new_n19527 , new_n19536 );
and  g17189 ( new_n19538 , new_n19526 , new_n19537 );
nor  g17190 ( new_n19539_1 , new_n19525 , new_n19538 );
xor  g17191 ( new_n19540 , new_n19524 , new_n19539_1 );
xnor g17192 ( new_n19541 , new_n19523_1 , new_n19540 );
xor  g17193 ( new_n19542 , new_n19506 , new_n19519 );
xor  g17194 ( new_n19543 , new_n19526 , new_n19537 );
and  g17195 ( new_n19544 , new_n19542 , new_n19543 );
xnor g17196 ( new_n19545 , new_n19542 , new_n19543 );
xor  g17197 ( new_n19546 , new_n19509 , new_n19517 );
xor  g17198 ( new_n19547 , new_n19528 , new_n19535 );
and  g17199 ( new_n19548 , new_n19546 , new_n19547 );
xnor g17200 ( new_n19549 , new_n19546 , new_n19547 );
xnor g17201 ( new_n19550 , new_n19512 , new_n19515_1 );
xnor g17202 ( new_n19551 , new_n19532 , new_n19533 );
nor  g17203 ( new_n19552 , new_n19550 , new_n19551 );
xnor g17204 ( new_n19553 , new_n19550 , new_n19551 );
nor  g17205 ( new_n19554 , new_n13432 , new_n13451 );
nor  g17206 ( new_n19555 , new_n13452 , new_n13482 );
nor  g17207 ( new_n19556 , new_n19554 , new_n19555 );
nor  g17208 ( new_n19557 , new_n19553 , new_n19556 );
nor  g17209 ( new_n19558 , new_n19552 , new_n19557 );
nor  g17210 ( new_n19559 , new_n19549 , new_n19558 );
nor  g17211 ( new_n19560 , new_n19548 , new_n19559 );
nor  g17212 ( new_n19561 , new_n19545 , new_n19560 );
nor  g17213 ( new_n19562 , new_n19544 , new_n19561 );
xnor g17214 ( n6576 , new_n19541 , new_n19562 );
xnor g17215 ( new_n19564 , new_n16708 , new_n19284 );
xnor g17216 ( n6587 , new_n19287 , new_n19564 );
xnor g17217 ( n6612 , new_n18234 , new_n18280 );
nor  g17218 ( new_n19567 , new_n10685 , new_n16992 );
xnor g17219 ( new_n19568 , new_n10685 , new_n16992 );
nor  g17220 ( new_n19569 , new_n10676 , new_n16994_1 );
xnor g17221 ( new_n19570_1 , new_n10676 , new_n16994_1 );
nor  g17222 ( new_n19571 , new_n10667 , new_n16997 );
xnor g17223 ( new_n19572 , new_n10667 , new_n16997 );
nor  g17224 ( new_n19573 , new_n10658 , new_n17000 );
xnor g17225 ( new_n19574 , new_n10658 , new_n17000 );
nor  g17226 ( new_n19575_1 , new_n10649 , new_n17003 );
xnor g17227 ( new_n19576 , new_n10649 , new_n17003 );
nor  g17228 ( new_n19577 , new_n10639 , new_n17005 );
xnor g17229 ( new_n19578 , new_n10639 , new_n17005 );
nor  g17230 ( new_n19579 , new_n10629 , new_n14750 );
xnor g17231 ( new_n19580 , new_n10629 , new_n14750 );
nor  g17232 ( new_n19581 , new_n10620 , new_n14753 );
nor  g17233 ( new_n19582 , n18 , new_n10607 );
and  g17234 ( new_n19583 , new_n9099 , new_n19582 );
nor  g17235 ( new_n19584_1 , new_n14756 , new_n19582 );
nor  g17236 ( new_n19585 , new_n19583 , new_n19584_1 );
and  g17237 ( new_n19586 , new_n10611_1 , new_n19585 );
nor  g17238 ( new_n19587 , new_n19583 , new_n19586 );
xnor g17239 ( new_n19588 , new_n10620 , new_n14752 );
and  g17240 ( new_n19589 , new_n19587 , new_n19588 );
or   g17241 ( new_n19590 , new_n19581 , new_n19589 );
nor  g17242 ( new_n19591 , new_n19580 , new_n19590 );
nor  g17243 ( new_n19592 , new_n19579 , new_n19591 );
nor  g17244 ( new_n19593 , new_n19578 , new_n19592 );
nor  g17245 ( new_n19594 , new_n19577 , new_n19593 );
nor  g17246 ( new_n19595 , new_n19576 , new_n19594 );
nor  g17247 ( new_n19596 , new_n19575_1 , new_n19595 );
nor  g17248 ( new_n19597 , new_n19574 , new_n19596 );
nor  g17249 ( new_n19598 , new_n19573 , new_n19597 );
nor  g17250 ( new_n19599 , new_n19572 , new_n19598 );
nor  g17251 ( new_n19600 , new_n19571 , new_n19599 );
nor  g17252 ( new_n19601 , new_n19570_1 , new_n19600 );
nor  g17253 ( new_n19602_1 , new_n19569 , new_n19601 );
nor  g17254 ( new_n19603 , new_n19568 , new_n19602_1 );
nor  g17255 ( new_n19604 , new_n19567 , new_n19603 );
and  g17256 ( new_n19605 , new_n17625 , new_n16991 );
and  g17257 ( new_n19606 , new_n19605 , new_n17634 );
and  g17258 ( new_n19607 , new_n19604 , new_n19606 );
or   g17259 ( new_n19608_1 , new_n19605 , new_n17634 );
nor  g17260 ( new_n19609 , new_n19604 , new_n19608_1 );
nor  g17261 ( new_n19610 , new_n19607 , new_n19609 );
xnor g17262 ( new_n19611 , new_n19605 , new_n17181 );
xnor g17263 ( new_n19612 , new_n19604 , new_n19611 );
nor  g17264 ( new_n19613 , new_n18899 , new_n19612 );
xnor g17265 ( new_n19614 , new_n18899 , new_n19612 );
xor  g17266 ( new_n19615 , new_n19568 , new_n19602_1 );
and  g17267 ( new_n19616 , new_n18904 , new_n19615 );
xnor g17268 ( new_n19617_1 , new_n18904 , new_n19615 );
xor  g17269 ( new_n19618_1 , new_n19570_1 , new_n19600 );
and  g17270 ( new_n19619 , new_n18908 , new_n19618_1 );
xnor g17271 ( new_n19620 , new_n18908 , new_n19618_1 );
xor  g17272 ( new_n19621 , new_n19572 , new_n19598 );
and  g17273 ( new_n19622 , new_n18912 , new_n19621 );
xnor g17274 ( new_n19623_1 , new_n18912 , new_n19621 );
xor  g17275 ( new_n19624 , new_n19574 , new_n19596 );
and  g17276 ( new_n19625 , new_n9350 , new_n19624 );
xnor g17277 ( new_n19626 , new_n9350 , new_n19624 );
xor  g17278 ( new_n19627 , new_n19576 , new_n19594 );
and  g17279 ( new_n19628 , new_n9354 , new_n19627 );
xnor g17280 ( new_n19629 , new_n9354 , new_n19627 );
xor  g17281 ( new_n19630 , new_n19578 , new_n19592 );
and  g17282 ( new_n19631 , new_n9359 , new_n19630 );
xnor g17283 ( new_n19632 , new_n9359 , new_n19630 );
xor  g17284 ( new_n19633 , new_n19580 , new_n19590 );
and  g17285 ( new_n19634 , new_n9364_1 , new_n19633 );
xnor g17286 ( new_n19635 , new_n9364_1 , new_n19633 );
xor  g17287 ( new_n19636 , new_n19587 , new_n19588 );
nor  g17288 ( new_n19637 , new_n9370 , new_n19636 );
xnor g17289 ( new_n19638 , new_n9370 , new_n19636 );
xnor g17290 ( new_n19639 , new_n13147 , new_n19585 );
and  g17291 ( new_n19640 , new_n9373 , new_n19639 );
xnor g17292 ( new_n19641_1 , new_n6596_1 , new_n10607 );
nor  g17293 ( new_n19642 , new_n9377 , new_n19641_1 );
xnor g17294 ( new_n19643 , new_n9373 , new_n19639 );
nor  g17295 ( new_n19644 , new_n19642 , new_n19643 );
nor  g17296 ( new_n19645 , new_n19640 , new_n19644 );
nor  g17297 ( new_n19646 , new_n19638 , new_n19645 );
nor  g17298 ( new_n19647 , new_n19637 , new_n19646 );
nor  g17299 ( new_n19648_1 , new_n19635 , new_n19647 );
nor  g17300 ( new_n19649 , new_n19634 , new_n19648_1 );
nor  g17301 ( new_n19650 , new_n19632 , new_n19649 );
nor  g17302 ( new_n19651 , new_n19631 , new_n19650 );
nor  g17303 ( new_n19652_1 , new_n19629 , new_n19651 );
nor  g17304 ( new_n19653 , new_n19628 , new_n19652_1 );
nor  g17305 ( new_n19654 , new_n19626 , new_n19653 );
nor  g17306 ( new_n19655 , new_n19625 , new_n19654 );
nor  g17307 ( new_n19656 , new_n19623_1 , new_n19655 );
nor  g17308 ( new_n19657 , new_n19622 , new_n19656 );
nor  g17309 ( new_n19658 , new_n19620 , new_n19657 );
nor  g17310 ( new_n19659 , new_n19619 , new_n19658 );
nor  g17311 ( new_n19660 , new_n19617_1 , new_n19659 );
nor  g17312 ( new_n19661 , new_n19616 , new_n19660 );
nor  g17313 ( new_n19662 , new_n19614 , new_n19661 );
or   g17314 ( new_n19663 , new_n19613 , new_n19662 );
not  g17315 ( new_n19664_1 , new_n19663 );
xnor g17316 ( new_n19665 , new_n18895 , new_n19664_1 );
xnor g17317 ( n6628 , new_n19610 , new_n19665 );
xnor g17318 ( n6630 , new_n2815 , new_n2835 );
not  g17319 ( new_n19668 , n17911 );
xnor g17320 ( new_n19669 , new_n19668 , n25331 );
nor  g17321 ( new_n19670 , n18483 , n21997 );
and  g17322 ( new_n19671 , new_n18976 , new_n18983 );
or   g17323 ( new_n19672 , new_n19670 , new_n19671 );
xor  g17324 ( new_n19673 , new_n19669 , new_n19672 );
xnor g17325 ( new_n19674 , new_n7487 , new_n19673 );
nor  g17326 ( new_n19675 , new_n7479 , new_n18984 );
and  g17327 ( new_n19676 , new_n18985 , new_n18994 );
or   g17328 ( new_n19677 , new_n19675 , new_n19676 );
xor  g17329 ( new_n19678 , new_n19674 , new_n19677 );
xnor g17330 ( new_n19679 , n468 , n14130 );
nor  g17331 ( new_n19680_1 , new_n8280 , n16482 );
xnor g17332 ( new_n19681 , n5400 , n16482 );
nor  g17333 ( new_n19682 , n9942 , new_n8284 );
nor  g17334 ( new_n19683 , new_n8353 , n25643 );
xnor g17335 ( new_n19684 , n329 , n25643 );
nor  g17336 ( new_n19685 , n9557 , new_n13046 );
xnor g17337 ( new_n19686 , n9557 , n24170 );
nor  g17338 ( new_n19687 , n2409 , new_n5106 );
xnor g17339 ( new_n19688 , n2409 , n3136 );
nor  g17340 ( new_n19689 , new_n2359 , n8869 );
and  g17341 ( new_n19690 , new_n18605 , new_n18608 );
or   g17342 ( new_n19691 , new_n19689 , new_n19690 );
and  g17343 ( new_n19692 , new_n19688 , new_n19691 );
nor  g17344 ( new_n19693 , new_n19687 , new_n19692 );
and  g17345 ( new_n19694 , new_n19686 , new_n19693 );
or   g17346 ( new_n19695 , new_n19685 , new_n19694 );
and  g17347 ( new_n19696 , new_n19684 , new_n19695 );
or   g17348 ( new_n19697 , new_n19683 , new_n19696 );
xnor g17349 ( new_n19698 , n9942 , n23923 );
and  g17350 ( new_n19699 , new_n19697 , new_n19698 );
or   g17351 ( new_n19700 , new_n19682 , new_n19699 );
and  g17352 ( new_n19701_1 , new_n19681 , new_n19700 );
or   g17353 ( new_n19702 , new_n19680_1 , new_n19701_1 );
xor  g17354 ( new_n19703 , new_n19679 , new_n19702 );
xor  g17355 ( new_n19704 , new_n19678 , new_n19703 );
xor  g17356 ( new_n19705 , new_n19681 , new_n19700 );
nor  g17357 ( new_n19706 , new_n18995 , new_n19705 );
xnor g17358 ( new_n19707 , new_n18995 , new_n19705 );
not  g17359 ( new_n19708 , new_n19707 );
xor  g17360 ( new_n19709 , new_n19697 , new_n19698 );
and  g17361 ( new_n19710 , new_n18999_1 , new_n19709 );
xor  g17362 ( new_n19711 , new_n19684 , new_n19695 );
nor  g17363 ( new_n19712 , new_n18645 , new_n19711 );
xnor g17364 ( new_n19713 , new_n18645 , new_n19711 );
xnor g17365 ( new_n19714 , new_n19686 , new_n19693 );
and  g17366 ( new_n19715 , new_n18670 , new_n19714 );
xnor g17367 ( new_n19716 , new_n18670 , new_n19714 );
xor  g17368 ( new_n19717 , new_n19688 , new_n19691 );
and  g17369 ( new_n19718 , new_n18672 , new_n19717 );
xnor g17370 ( new_n19719 , new_n18672 , new_n19717 );
and  g17371 ( new_n19720 , new_n18676 , new_n18609 );
and  g17372 ( new_n19721 , new_n18610_1 , new_n18613 );
nor  g17373 ( new_n19722 , new_n19720 , new_n19721 );
nor  g17374 ( new_n19723 , new_n19719 , new_n19722 );
nor  g17375 ( new_n19724 , new_n19718 , new_n19723 );
nor  g17376 ( new_n19725 , new_n19716 , new_n19724 );
nor  g17377 ( new_n19726 , new_n19715 , new_n19725 );
nor  g17378 ( new_n19727 , new_n19713 , new_n19726 );
nor  g17379 ( new_n19728 , new_n19712 , new_n19727 );
xnor g17380 ( new_n19729 , new_n19004 , new_n19709 );
and  g17381 ( new_n19730 , new_n19728 , new_n19729 );
nor  g17382 ( new_n19731 , new_n19710 , new_n19730 );
and  g17383 ( new_n19732 , new_n19708 , new_n19731 );
nor  g17384 ( new_n19733 , new_n19706 , new_n19732 );
xor  g17385 ( n6634 , new_n19704 , new_n19733 );
xnor g17386 ( n6652 , new_n6563 , new_n6577 );
xnor g17387 ( n6655 , new_n12331 , new_n12344 );
xnor g17388 ( n6669 , new_n11874 , new_n11892 );
xnor g17389 ( n6671 , new_n9367 , new_n9385 );
xnor g17390 ( n6673 , new_n13279 , new_n13296 );
and  g17391 ( new_n19740 , new_n19460 , new_n19466 );
or   g17392 ( new_n19741 , new_n11793 , new_n11336 );
nor  g17393 ( new_n19742 , new_n19741 , new_n19464 );
or   g17394 ( n6674 , new_n19740 , new_n19742 );
xnor g17395 ( n6684 , new_n16206_1 , new_n16215_1 );
xor  g17396 ( n6706 , new_n12061 , new_n12106 );
xnor g17397 ( new_n19746 , n8614 , n12702 );
nor  g17398 ( new_n19747 , n15182 , n26797 );
xnor g17399 ( new_n19748 , n15182 , n26797 );
nor  g17400 ( new_n19749_1 , n23913 , n27037 );
xnor g17401 ( new_n19750 , n23913 , n27037 );
nor  g17402 ( new_n19751 , n8964 , n22554 );
xnor g17403 ( new_n19752 , n8964 , n22554 );
nor  g17404 ( new_n19753 , n20151 , n20429 );
xnor g17405 ( new_n19754 , n20151 , n20429 );
nor  g17406 ( new_n19755 , n3909 , n7693 );
xnor g17407 ( new_n19756_1 , n3909 , n7693 );
nor  g17408 ( new_n19757 , n10405 , n23974 );
xnor g17409 ( new_n19758 , new_n4021 , n23974 );
nor  g17410 ( new_n19759 , new_n8050 , new_n4106 );
or   g17411 ( new_n19760 , n2146 , n11302 );
nor  g17412 ( new_n19761 , n17090 , n22173 );
nor  g17413 ( new_n19762 , new_n15352 , new_n15353_1 );
nor  g17414 ( new_n19763 , new_n19761 , new_n19762 );
and  g17415 ( new_n19764 , new_n19760 , new_n19763 );
nor  g17416 ( new_n19765 , new_n19759 , new_n19764 );
and  g17417 ( new_n19766 , new_n19758 , new_n19765 );
nor  g17418 ( new_n19767_1 , new_n19757 , new_n19766 );
nor  g17419 ( new_n19768 , new_n19756_1 , new_n19767_1 );
nor  g17420 ( new_n19769 , new_n19755 , new_n19768 );
nor  g17421 ( new_n19770_1 , new_n19754 , new_n19769 );
nor  g17422 ( new_n19771 , new_n19753 , new_n19770_1 );
nor  g17423 ( new_n19772 , new_n19752 , new_n19771 );
nor  g17424 ( new_n19773 , new_n19751 , new_n19772 );
nor  g17425 ( new_n19774 , new_n19750 , new_n19773 );
nor  g17426 ( new_n19775 , new_n19749_1 , new_n19774 );
nor  g17427 ( new_n19776 , new_n19748 , new_n19775 );
nor  g17428 ( new_n19777 , new_n19747 , new_n19776 );
xnor g17429 ( new_n19778 , new_n19746 , new_n19777 );
nor  g17430 ( new_n19779 , new_n6152 , new_n19778 );
xnor g17431 ( new_n19780_1 , new_n6152 , new_n19778 );
xnor g17432 ( new_n19781 , new_n19748 , new_n19775 );
nor  g17433 ( new_n19782 , new_n13645 , new_n19781 );
xnor g17434 ( new_n19783 , new_n13645 , new_n19781 );
xnor g17435 ( new_n19784 , new_n19750 , new_n19773 );
nor  g17436 ( new_n19785 , new_n13648 , new_n19784 );
xnor g17437 ( new_n19786 , new_n13648 , new_n19784 );
xnor g17438 ( new_n19787 , new_n19752 , new_n19771 );
nor  g17439 ( new_n19788 , new_n13651 , new_n19787 );
xnor g17440 ( new_n19789_1 , new_n13651 , new_n19787 );
xnor g17441 ( new_n19790 , new_n19754 , new_n19769 );
nor  g17442 ( new_n19791 , new_n6164 , new_n19790 );
xnor g17443 ( new_n19792_1 , new_n6164 , new_n19790 );
xnor g17444 ( new_n19793 , new_n19756_1 , new_n19767_1 );
nor  g17445 ( new_n19794 , new_n6167 , new_n19793 );
xnor g17446 ( new_n19795 , new_n6167 , new_n19793 );
xnor g17447 ( new_n19796 , new_n19758 , new_n19765 );
not  g17448 ( new_n19797 , new_n19796 );
and  g17449 ( new_n19798_1 , n20169 , new_n19797 );
xnor g17450 ( new_n19799 , n20169 , new_n19797 );
xnor g17451 ( new_n19800 , n2146 , n11302 );
xnor g17452 ( new_n19801 , new_n19763 , new_n19800 );
nor  g17453 ( new_n19802 , new_n6173 , new_n19801 );
xnor g17454 ( new_n19803_1 , n8285 , new_n19801 );
and  g17455 ( new_n19804 , new_n15351 , new_n15354 );
or   g17456 ( new_n19805 , new_n15350 , new_n19804 );
and  g17457 ( new_n19806 , new_n19803_1 , new_n19805 );
nor  g17458 ( new_n19807 , new_n19802 , new_n19806 );
nor  g17459 ( new_n19808 , new_n19799 , new_n19807 );
nor  g17460 ( new_n19809 , new_n19798_1 , new_n19808 );
nor  g17461 ( new_n19810 , new_n19795 , new_n19809 );
nor  g17462 ( new_n19811 , new_n19794 , new_n19810 );
nor  g17463 ( new_n19812 , new_n19792_1 , new_n19811 );
nor  g17464 ( new_n19813 , new_n19791 , new_n19812 );
nor  g17465 ( new_n19814 , new_n19789_1 , new_n19813 );
nor  g17466 ( new_n19815 , new_n19788 , new_n19814 );
nor  g17467 ( new_n19816 , new_n19786 , new_n19815 );
nor  g17468 ( new_n19817 , new_n19785 , new_n19816 );
nor  g17469 ( new_n19818 , new_n19783 , new_n19817 );
nor  g17470 ( new_n19819 , new_n19782 , new_n19818 );
nor  g17471 ( new_n19820 , new_n19780_1 , new_n19819 );
nor  g17472 ( new_n19821 , new_n19779 , new_n19820 );
nor  g17473 ( new_n19822 , n8614 , n12702 );
nor  g17474 ( new_n19823 , new_n19746 , new_n19777 );
nor  g17475 ( new_n19824 , new_n19822 , new_n19823 );
xnor g17476 ( new_n19825 , new_n19821 , new_n19824 );
and  g17477 ( new_n19826 , new_n4477 , new_n19502 );
and  g17478 ( new_n19827 , new_n19503 , new_n19521 );
nor  g17479 ( new_n19828 , new_n19826 , new_n19827 );
not  g17480 ( new_n19829 , new_n19828 );
not  g17481 ( new_n19830 , new_n19501 );
nor  g17482 ( new_n19831 , n1536 , new_n19830 );
xnor g17483 ( new_n19832 , new_n4538 , new_n19831 );
xnor g17484 ( new_n19833 , new_n19829 , new_n19832 );
xnor g17485 ( new_n19834 , new_n19825 , new_n19833 );
xnor g17486 ( new_n19835 , new_n19780_1 , new_n19819 );
nor  g17487 ( new_n19836 , new_n19523_1 , new_n19835 );
xnor g17488 ( new_n19837 , new_n19523_1 , new_n19835 );
xnor g17489 ( new_n19838 , new_n19783 , new_n19817 );
not  g17490 ( new_n19839 , new_n19838 );
and  g17491 ( new_n19840 , new_n19542 , new_n19839 );
xnor g17492 ( new_n19841 , new_n19542 , new_n19839 );
xnor g17493 ( new_n19842 , new_n19786 , new_n19815 );
not  g17494 ( new_n19843 , new_n19842 );
and  g17495 ( new_n19844 , new_n19546 , new_n19843 );
xnor g17496 ( new_n19845 , new_n19546 , new_n19843 );
xnor g17497 ( new_n19846 , new_n19789_1 , new_n19813 );
nor  g17498 ( new_n19847 , new_n19550 , new_n19846 );
xnor g17499 ( new_n19848 , new_n19550 , new_n19846 );
xnor g17500 ( new_n19849 , new_n19792_1 , new_n19811 );
nor  g17501 ( new_n19850 , new_n13432 , new_n19849 );
xnor g17502 ( new_n19851 , new_n13432 , new_n19849 );
xnor g17503 ( new_n19852 , new_n19795 , new_n19809 );
nor  g17504 ( new_n19853 , new_n13454 , new_n19852 );
xnor g17505 ( new_n19854 , new_n13454 , new_n19852 );
xnor g17506 ( new_n19855 , new_n19799 , new_n19807 );
nor  g17507 ( new_n19856 , new_n13458 , new_n19855 );
xor  g17508 ( new_n19857 , new_n13458 , new_n19855 );
xor  g17509 ( new_n19858 , new_n19803_1 , new_n19805 );
nor  g17510 ( new_n19859 , new_n13462 , new_n19858 );
and  g17511 ( new_n19860 , new_n13466 , new_n15356 );
nor  g17512 ( new_n19861 , new_n15346 , new_n15357 );
nor  g17513 ( new_n19862 , new_n19860 , new_n19861 );
xor  g17514 ( new_n19863 , new_n13462 , new_n19858 );
and  g17515 ( new_n19864 , new_n19862 , new_n19863 );
nor  g17516 ( new_n19865 , new_n19859 , new_n19864 );
and  g17517 ( new_n19866 , new_n19857 , new_n19865 );
nor  g17518 ( new_n19867 , new_n19856 , new_n19866 );
nor  g17519 ( new_n19868 , new_n19854 , new_n19867 );
nor  g17520 ( new_n19869 , new_n19853 , new_n19868 );
nor  g17521 ( new_n19870 , new_n19851 , new_n19869 );
nor  g17522 ( new_n19871 , new_n19850 , new_n19870 );
nor  g17523 ( new_n19872 , new_n19848 , new_n19871 );
nor  g17524 ( new_n19873_1 , new_n19847 , new_n19872 );
nor  g17525 ( new_n19874 , new_n19845 , new_n19873_1 );
nor  g17526 ( new_n19875 , new_n19844 , new_n19874 );
nor  g17527 ( new_n19876 , new_n19841 , new_n19875 );
nor  g17528 ( new_n19877 , new_n19840 , new_n19876 );
nor  g17529 ( new_n19878 , new_n19837 , new_n19877 );
nor  g17530 ( new_n19879 , new_n19836 , new_n19878 );
xnor g17531 ( n6707 , new_n19834 , new_n19879 );
xnor g17532 ( n6736 , new_n12645 , new_n12872 );
xnor g17533 ( new_n19882 , n5101 , n23895 );
and  g17534 ( new_n19883 , n16507 , new_n5456 );
xnor g17535 ( new_n19884 , n16507 , n17351 );
and  g17536 ( new_n19885 , new_n5459 , n22470 );
xnor g17537 ( new_n19886 , n11736 , n22470 );
and  g17538 ( new_n19887 , n19116 , new_n5462 );
and  g17539 ( new_n19888 , n6861 , new_n5465 );
and  g17540 ( new_n19889 , new_n17514 , new_n17531 );
or   g17541 ( new_n19890 , new_n19888 , new_n19889 );
xnor g17542 ( new_n19891 , n19116 , n23200 );
and  g17543 ( new_n19892 , new_n19890 , new_n19891 );
or   g17544 ( new_n19893 , new_n19887 , new_n19892 );
and  g17545 ( new_n19894 , new_n19886 , new_n19893 );
or   g17546 ( new_n19895 , new_n19885 , new_n19894 );
and  g17547 ( new_n19896 , new_n19884 , new_n19895 );
or   g17548 ( new_n19897 , new_n19883 , new_n19896 );
xor  g17549 ( new_n19898 , new_n19882 , new_n19897 );
not  g17550 ( new_n19899 , new_n17539 );
nor  g17551 ( new_n19900 , n22660 , new_n19899 );
not  g17552 ( new_n19901 , new_n19900 );
nor  g17553 ( new_n19902 , n13490 , new_n19901 );
not  g17554 ( new_n19903 , new_n19902 );
nor  g17555 ( new_n19904 , n9655 , new_n19903 );
not  g17556 ( new_n19905_1 , new_n19904 );
nor  g17557 ( new_n19906 , n25345 , new_n19905_1 );
xnor g17558 ( new_n19907 , n13494 , new_n19906 );
xnor g17559 ( new_n19908 , n12650 , new_n19907 );
xnor g17560 ( new_n19909_1 , n25345 , new_n19904 );
nor  g17561 ( new_n19910 , new_n5560 , new_n19909_1 );
xnor g17562 ( new_n19911_1 , n10201 , new_n19909_1 );
xnor g17563 ( new_n19912 , n9655 , new_n19902 );
nor  g17564 ( new_n19913 , new_n5564_1 , new_n19912 );
xnor g17565 ( new_n19914 , new_n5564_1 , new_n19912 );
xnor g17566 ( new_n19915 , n13490 , new_n19900 );
nor  g17567 ( new_n19916_1 , new_n5568 , new_n19915 );
xnor g17568 ( new_n19917 , n18290 , new_n19915 );
nor  g17569 ( new_n19918 , new_n5572 , new_n17540 );
and  g17570 ( new_n19919 , new_n17541 , new_n17562 );
or   g17571 ( new_n19920 , new_n19918 , new_n19919 );
and  g17572 ( new_n19921 , new_n19917 , new_n19920 );
nor  g17573 ( new_n19922_1 , new_n19916_1 , new_n19921 );
nor  g17574 ( new_n19923_1 , new_n19914 , new_n19922_1 );
or   g17575 ( new_n19924 , new_n19913 , new_n19923_1 );
and  g17576 ( new_n19925 , new_n19911_1 , new_n19924 );
or   g17577 ( new_n19926 , new_n19910 , new_n19925 );
xor  g17578 ( new_n19927 , new_n19908 , new_n19926 );
xnor g17579 ( new_n19928 , new_n15563 , new_n19927 );
xor  g17580 ( new_n19929 , new_n19911_1 , new_n19924 );
nor  g17581 ( new_n19930_1 , new_n15567 , new_n19929 );
xnor g17582 ( new_n19931 , new_n19914 , new_n19922_1 );
nor  g17583 ( new_n19932 , new_n15574 , new_n19931 );
xnor g17584 ( new_n19933 , new_n15572 , new_n19931 );
xor  g17585 ( new_n19934 , new_n19917 , new_n19920 );
nor  g17586 ( new_n19935 , new_n15577 , new_n19934 );
xnor g17587 ( new_n19936 , new_n15577 , new_n19934 );
nor  g17588 ( new_n19937 , new_n15581 , new_n17563 );
nor  g17589 ( new_n19938 , new_n17564 , new_n17587 );
nor  g17590 ( new_n19939 , new_n19937 , new_n19938 );
nor  g17591 ( new_n19940 , new_n19936 , new_n19939 );
nor  g17592 ( new_n19941_1 , new_n19935 , new_n19940 );
and  g17593 ( new_n19942 , new_n19933 , new_n19941_1 );
nor  g17594 ( new_n19943 , new_n19932 , new_n19942 );
xnor g17595 ( new_n19944 , new_n15569 , new_n19929 );
and  g17596 ( new_n19945 , new_n19943 , new_n19944 );
nor  g17597 ( new_n19946 , new_n19930_1 , new_n19945 );
xnor g17598 ( new_n19947 , new_n19928 , new_n19946 );
xnor g17599 ( new_n19948 , new_n19898 , new_n19947 );
xor  g17600 ( new_n19949 , new_n19884 , new_n19895 );
xor  g17601 ( new_n19950 , new_n19943 , new_n19944 );
nor  g17602 ( new_n19951 , new_n19949 , new_n19950 );
xnor g17603 ( new_n19952 , new_n19949 , new_n19950 );
xor  g17604 ( new_n19953 , new_n19886 , new_n19893 );
xnor g17605 ( new_n19954 , new_n19933 , new_n19941_1 );
nor  g17606 ( new_n19955 , new_n19953 , new_n19954 );
not  g17607 ( new_n19956 , new_n19954 );
xnor g17608 ( new_n19957 , new_n19953 , new_n19956 );
xor  g17609 ( new_n19958 , new_n19890 , new_n19891 );
xnor g17610 ( new_n19959 , new_n19936 , new_n19939 );
not  g17611 ( new_n19960 , new_n19959 );
and  g17612 ( new_n19961 , new_n19958 , new_n19960 );
xnor g17613 ( new_n19962 , new_n19958 , new_n19959 );
not  g17614 ( new_n19963 , new_n17588 );
and  g17615 ( new_n19964 , new_n17532 , new_n19963 );
and  g17616 ( new_n19965 , new_n17589 , new_n17621 );
or   g17617 ( new_n19966 , new_n19964 , new_n19965 );
and  g17618 ( new_n19967 , new_n19962 , new_n19966 );
nor  g17619 ( new_n19968_1 , new_n19961 , new_n19967 );
and  g17620 ( new_n19969 , new_n19957 , new_n19968_1 );
nor  g17621 ( new_n19970 , new_n19955 , new_n19969 );
nor  g17622 ( new_n19971 , new_n19952 , new_n19970 );
nor  g17623 ( new_n19972 , new_n19951 , new_n19971 );
xor  g17624 ( n6791 , new_n19948 , new_n19972 );
xnor g17625 ( n6802 , new_n3700 , new_n3709 );
xnor g17626 ( n6826 , new_n15894 , new_n15917_1 );
xnor g17627 ( n6835 , new_n9945 , new_n9972 );
nor  g17628 ( new_n19977 , new_n10030 , new_n17829 );
xnor g17629 ( new_n19978 , new_n10030 , new_n17831 );
nor  g17630 ( new_n19979 , new_n17810 , new_n2925 );
xnor g17631 ( new_n19980 , n22379 , new_n2925 );
nor  g17632 ( new_n19981 , new_n2850 , new_n2972 );
xnor g17633 ( new_n19982 , new_n2850 , new_n2976 );
nor  g17634 ( new_n19983 , new_n2853_1 , new_n2979_1 );
xnor g17635 ( new_n19984 , new_n2853_1 , new_n2980 );
nor  g17636 ( new_n19985 , new_n2856 , new_n2985_1 );
nor  g17637 ( new_n19986 , n5213 , new_n2990 );
xnor g17638 ( new_n19987 , new_n2859 , new_n2990 );
nor  g17639 ( new_n19988_1 , n4665 , new_n2996 );
xnor g17640 ( new_n19989 , new_n2862 , new_n2996 );
nor  g17641 ( new_n19990 , new_n2866 , new_n3002 );
xnor g17642 ( new_n19991 , n19005 , new_n3002 );
nor  g17643 ( new_n19992 , new_n5287 , new_n3063 );
nor  g17644 ( new_n19993 , n4326 , new_n19992 );
xnor g17645 ( new_n19994 , new_n2869 , new_n19992 );
and  g17646 ( new_n19995 , new_n3008 , new_n19994 );
nor  g17647 ( new_n19996 , new_n19993 , new_n19995 );
and  g17648 ( new_n19997 , new_n19991 , new_n19996 );
nor  g17649 ( new_n19998 , new_n19990 , new_n19997 );
and  g17650 ( new_n19999 , new_n19989 , new_n19998 );
or   g17651 ( new_n20000 , new_n19988_1 , new_n19999 );
and  g17652 ( new_n20001 , new_n19987 , new_n20000 );
nor  g17653 ( new_n20002 , new_n19986 , new_n20001 );
xnor g17654 ( new_n20003 , new_n2856 , new_n2986 );
and  g17655 ( new_n20004_1 , new_n20002 , new_n20003 );
or   g17656 ( new_n20005 , new_n19985 , new_n20004_1 );
and  g17657 ( new_n20006 , new_n19984 , new_n20005 );
or   g17658 ( new_n20007 , new_n19983 , new_n20006 );
and  g17659 ( new_n20008 , new_n19982 , new_n20007 );
or   g17660 ( new_n20009 , new_n19981 , new_n20008 );
and  g17661 ( new_n20010 , new_n19980 , new_n20009 );
or   g17662 ( new_n20011 , new_n19979 , new_n20010 );
and  g17663 ( new_n20012 , new_n19978 , new_n20011 );
nor  g17664 ( new_n20013_1 , new_n19977 , new_n20012 );
nor  g17665 ( new_n20014 , new_n17823 , new_n20013_1 );
xnor g17666 ( new_n20015 , new_n17498 , new_n20014 );
xnor g17667 ( new_n20016 , new_n17823 , new_n20013_1 );
and  g17668 ( new_n20017_1 , new_n17500_1 , new_n20016 );
xnor g17669 ( new_n20018 , new_n17500_1 , new_n20016 );
xor  g17670 ( new_n20019 , new_n19978 , new_n20011 );
nor  g17671 ( new_n20020 , new_n12670_1 , new_n20019 );
xnor g17672 ( new_n20021 , new_n12670_1 , new_n20019 );
xor  g17673 ( new_n20022 , new_n19980 , new_n20009 );
nor  g17674 ( new_n20023 , new_n12698 , new_n20022 );
xnor g17675 ( new_n20024 , new_n12698 , new_n20022 );
not  g17676 ( new_n20025 , new_n6097 );
xor  g17677 ( new_n20026 , new_n19982 , new_n20007 );
nor  g17678 ( new_n20027 , new_n20025 , new_n20026 );
xnor g17679 ( new_n20028 , new_n20025 , new_n20026 );
xor  g17680 ( new_n20029 , new_n19984 , new_n20005 );
nor  g17681 ( new_n20030 , new_n12704 , new_n20029 );
xnor g17682 ( new_n20031 , new_n12704 , new_n20029 );
not  g17683 ( new_n20032 , new_n6107 );
xor  g17684 ( new_n20033_1 , new_n20002 , new_n20003 );
nor  g17685 ( new_n20034 , new_n20032 , new_n20033_1 );
xnor g17686 ( new_n20035 , new_n20032 , new_n20033_1 );
xor  g17687 ( new_n20036_1 , new_n19987 , new_n20000 );
and  g17688 ( new_n20037 , new_n6112 , new_n20036_1 );
xnor g17689 ( new_n20038 , new_n6112 , new_n20036_1 );
xnor g17690 ( new_n20039 , new_n19989 , new_n19998 );
not  g17691 ( new_n20040_1 , new_n20039 );
and  g17692 ( new_n20041 , new_n6116 , new_n20040_1 );
xnor g17693 ( new_n20042 , new_n6116 , new_n20040_1 );
xor  g17694 ( new_n20043 , new_n19991 , new_n19996 );
nor  g17695 ( new_n20044 , new_n6121 , new_n20043 );
xnor g17696 ( new_n20045 , new_n6121 , new_n20043 );
xnor g17697 ( new_n20046 , new_n3009 , new_n19994 );
and  g17698 ( new_n20047 , new_n6132 , new_n20046 );
nor  g17699 ( new_n20048 , new_n5794 , new_n5795 );
xnor g17700 ( new_n20049 , new_n6126 , new_n20046 );
and  g17701 ( new_n20050 , new_n20048 , new_n20049 );
nor  g17702 ( new_n20051 , new_n20047 , new_n20050 );
nor  g17703 ( new_n20052 , new_n20045 , new_n20051 );
nor  g17704 ( new_n20053 , new_n20044 , new_n20052 );
nor  g17705 ( new_n20054 , new_n20042 , new_n20053 );
nor  g17706 ( new_n20055 , new_n20041 , new_n20054 );
nor  g17707 ( new_n20056 , new_n20038 , new_n20055 );
nor  g17708 ( new_n20057 , new_n20037 , new_n20056 );
nor  g17709 ( new_n20058 , new_n20035 , new_n20057 );
nor  g17710 ( new_n20059 , new_n20034 , new_n20058 );
nor  g17711 ( new_n20060 , new_n20031 , new_n20059 );
nor  g17712 ( new_n20061_1 , new_n20030 , new_n20060 );
nor  g17713 ( new_n20062 , new_n20028 , new_n20061_1 );
nor  g17714 ( new_n20063 , new_n20027 , new_n20062 );
nor  g17715 ( new_n20064 , new_n20024 , new_n20063 );
nor  g17716 ( new_n20065 , new_n20023 , new_n20064 );
nor  g17717 ( new_n20066 , new_n20021 , new_n20065 );
nor  g17718 ( new_n20067 , new_n20020 , new_n20066 );
nor  g17719 ( new_n20068 , new_n20018 , new_n20067 );
nor  g17720 ( new_n20069_1 , new_n20017_1 , new_n20068 );
xnor g17721 ( n6853 , new_n20015 , new_n20069_1 );
xnor g17722 ( new_n20071 , new_n11042 , new_n14607 );
nor  g17723 ( new_n20072 , new_n11048 , new_n14612 );
xnor g17724 ( new_n20073 , new_n11048 , new_n14610 );
nor  g17725 ( new_n20074 , new_n4194 , new_n11050 );
nor  g17726 ( new_n20075 , new_n12737 , new_n12750 );
nor  g17727 ( new_n20076 , new_n20074 , new_n20075 );
and  g17728 ( new_n20077_1 , new_n20073 , new_n20076 );
or   g17729 ( new_n20078 , new_n20072 , new_n20077_1 );
xor  g17730 ( n6862 , new_n20071 , new_n20078 );
and  g17731 ( new_n20080 , new_n7110 , n22253 );
and  g17732 ( new_n20081 , new_n15505 , new_n15520 );
nor  g17733 ( new_n20082 , new_n20080 , new_n20081 );
not  g17734 ( new_n20083 , n25296 );
nor  g17735 ( new_n20084 , n23717 , new_n20083 );
and  g17736 ( new_n20085 , new_n11187 , new_n11202 );
nor  g17737 ( new_n20086_1 , new_n20084 , new_n20085 );
nor  g17738 ( new_n20087 , new_n17984 , new_n20086_1 );
and  g17739 ( new_n20088 , new_n11186 , new_n11203 );
nor  g17740 ( new_n20089 , new_n11204 , new_n11225 );
nor  g17741 ( new_n20090 , new_n20088 , new_n20089 );
xnor g17742 ( new_n20091 , new_n17984 , new_n20086_1 );
nor  g17743 ( new_n20092 , new_n20090 , new_n20091 );
nor  g17744 ( new_n20093 , new_n20087 , new_n20092 );
and  g17745 ( new_n20094 , new_n20082 , new_n20093 );
not  g17746 ( new_n20095 , new_n11226 );
and  g17747 ( new_n20096_1 , new_n20095 , new_n15521 );
and  g17748 ( new_n20097 , new_n15522 , new_n15541 );
nor  g17749 ( new_n20098 , new_n20096_1 , new_n20097 );
nor  g17750 ( new_n20099 , new_n20093 , new_n20098 );
nor  g17751 ( new_n20100 , new_n20094 , new_n20099 );
xnor g17752 ( new_n20101 , new_n20090 , new_n20091 );
not  g17753 ( new_n20102 , new_n20101 );
nor  g17754 ( new_n20103_1 , new_n20082 , new_n20102 );
not  g17755 ( new_n20104 , new_n20098 );
nor  g17756 ( new_n20105 , new_n20104 , new_n20101 );
nor  g17757 ( new_n20106 , new_n20103_1 , new_n20105 );
and  g17758 ( n6863 , new_n20100 , new_n20106 );
xnor g17759 ( n6867 , new_n6094 , new_n6147 );
xnor g17760 ( n6965 , new_n17440_1 , new_n17448 );
xnor g17761 ( n6967 , new_n7379 , new_n7419 );
xor  g17762 ( n6975 , new_n14113 , new_n14160 );
xor  g17763 ( n6983 , new_n19439 , new_n19440 );
xnor g17764 ( new_n20113 , new_n11028 , new_n14586 );
nor  g17765 ( new_n20114 , new_n11030 , new_n14592 );
xnor g17766 ( new_n20115 , new_n11033 , new_n14591 );
nor  g17767 ( new_n20116 , new_n11035 , new_n14596 );
xnor g17768 ( new_n20117 , new_n11037 , new_n14596 );
not  g17769 ( new_n20118 , new_n11039 );
nor  g17770 ( new_n20119 , new_n20118 , new_n14603_1 );
nor  g17771 ( new_n20120 , new_n11044_1 , new_n14607 );
and  g17772 ( new_n20121 , new_n20071 , new_n20078 );
or   g17773 ( new_n20122 , new_n20120 , new_n20121 );
xnor g17774 ( new_n20123 , new_n20118 , new_n14600 );
and  g17775 ( new_n20124 , new_n20122 , new_n20123 );
nor  g17776 ( new_n20125 , new_n20119 , new_n20124 );
and  g17777 ( new_n20126_1 , new_n20117 , new_n20125 );
nor  g17778 ( new_n20127 , new_n20116 , new_n20126_1 );
nor  g17779 ( new_n20128 , new_n20115 , new_n20127 );
nor  g17780 ( new_n20129 , new_n20114 , new_n20128 );
xnor g17781 ( n6985 , new_n20113 , new_n20129 );
xnor g17782 ( n6998 , new_n14369 , new_n14407 );
not  g17783 ( new_n20132 , new_n8886 );
xnor g17784 ( n7032 , new_n20132 , new_n10992 );
xnor g17785 ( n7038 , new_n19267 , new_n19299 );
xnor g17786 ( n7079 , new_n17276 , new_n17277 );
xnor g17787 ( n7190 , new_n7407 , new_n7408_1 );
xnor g17788 ( n7229 , new_n15473 , new_n15476 );
xnor g17789 ( n7230 , new_n8550_1 , new_n8562 );
xnor g17790 ( n7233 , new_n18581 , new_n18582_1 );
xnor g17791 ( n7236 , new_n12971 , new_n12979 );
xnor g17792 ( n7253 , new_n6946 , new_n15806 );
and  g17793 ( new_n20142 , new_n10870 , new_n18929 );
nor  g17794 ( new_n20143 , n12507 , new_n18930 );
and  g17795 ( new_n20144 , n12507 , new_n18930 );
nor  g17796 ( new_n20145 , new_n20144 , new_n18934 );
nor  g17797 ( new_n20146 , new_n20143 , new_n20145 );
nor  g17798 ( new_n20147 , new_n20142 , new_n20146 );
not  g17799 ( new_n20148 , new_n19375 );
nor  g17800 ( new_n20149_1 , new_n13859 , new_n20148 );
xnor g17801 ( new_n20150 , new_n13823 , new_n20149_1 );
nor  g17802 ( new_n20151_1 , new_n10095 , new_n20150 );
xnor g17803 ( new_n20152 , new_n10054 , new_n20150 );
nor  g17804 ( new_n20153 , new_n10058 , new_n19376 );
and  g17805 ( new_n20154 , new_n19377 , new_n19415 );
or   g17806 ( new_n20155 , new_n20153 , new_n20154 );
and  g17807 ( new_n20156 , new_n20152 , new_n20155 );
nor  g17808 ( new_n20157 , new_n20151_1 , new_n20156 );
xor  g17809 ( new_n20158 , new_n13810 , new_n13822 );
and  g17810 ( new_n20159 , new_n20158 , new_n20149_1 );
nor  g17811 ( new_n20160 , new_n13869 , new_n20159 );
and  g17812 ( new_n20161 , new_n13866 , new_n20159 );
nor  g17813 ( new_n20162 , new_n20160 , new_n20161 );
xnor g17814 ( new_n20163 , new_n10044 , new_n20162 );
xnor g17815 ( new_n20164 , new_n20157 , new_n20163 );
nor  g17816 ( new_n20165 , new_n20147 , new_n20164 );
not  g17817 ( new_n20166 , new_n20147 );
xnor g17818 ( new_n20167 , new_n20166 , new_n20164 );
xor  g17819 ( new_n20168 , new_n20152 , new_n20155 );
nor  g17820 ( new_n20169_1 , new_n18935 , new_n20168 );
nor  g17821 ( new_n20170 , new_n16280 , new_n19416 );
and  g17822 ( new_n20171 , new_n19417 , new_n19455 );
nor  g17823 ( new_n20172 , new_n20170 , new_n20171 );
xnor g17824 ( new_n20173 , new_n18935 , new_n20168 );
nor  g17825 ( new_n20174 , new_n20172 , new_n20173 );
nor  g17826 ( new_n20175 , new_n20169_1 , new_n20174 );
and  g17827 ( new_n20176 , new_n20167 , new_n20175 );
nor  g17828 ( new_n20177 , new_n20165 , new_n20176 );
not  g17829 ( new_n20178 , new_n20177 );
and  g17830 ( new_n20179_1 , new_n10044 , new_n20162 );
or   g17831 ( new_n20180 , new_n10044 , new_n20162 );
and  g17832 ( new_n20181 , new_n20157 , new_n20180 );
or   g17833 ( new_n20182 , new_n20161 , new_n20181 );
nor  g17834 ( new_n20183 , new_n20179_1 , new_n20182 );
xnor g17835 ( n7256 , new_n20178 , new_n20183 );
not  g17836 ( new_n20185 , new_n15180_1 );
nor  g17837 ( new_n20186 , n2416 , new_n12048 );
xnor g17838 ( new_n20187_1 , n2416 , n22764 );
not  g17839 ( new_n20188 , n26264 );
nor  g17840 ( new_n20189 , n21905 , new_n20188 );
and  g17841 ( new_n20190 , new_n19015 , new_n19029 );
or   g17842 ( new_n20191 , new_n20189 , new_n20190 );
and  g17843 ( new_n20192 , new_n20187_1 , new_n20191 );
nor  g17844 ( new_n20193 , new_n20186 , new_n20192 );
xor  g17845 ( new_n20194 , new_n20187_1 , new_n20191 );
and  g17846 ( new_n20195 , new_n15184 , new_n20194 );
xnor g17847 ( new_n20196 , new_n15182_1 , new_n20194 );
and  g17848 ( new_n20197 , new_n15189 , new_n19030 );
and  g17849 ( new_n20198 , new_n19031 , new_n19044_1 );
or   g17850 ( new_n20199 , new_n20197 , new_n20198 );
and  g17851 ( new_n20200 , new_n20196 , new_n20199 );
nor  g17852 ( new_n20201 , new_n20195 , new_n20200 );
xnor g17853 ( new_n20202 , new_n20193 , new_n20201 );
xnor g17854 ( new_n20203 , new_n20185 , new_n20202 );
xnor g17855 ( new_n20204 , new_n19127 , new_n20203 );
xor  g17856 ( new_n20205 , new_n20196 , new_n20199 );
nor  g17857 ( new_n20206 , new_n19139 , new_n20205 );
xnor g17858 ( new_n20207 , new_n19139 , new_n20205 );
nor  g17859 ( new_n20208 , new_n19014 , new_n19045 );
nor  g17860 ( new_n20209 , new_n19046 , new_n19059 );
nor  g17861 ( new_n20210 , new_n20208 , new_n20209 );
nor  g17862 ( new_n20211 , new_n20207 , new_n20210 );
nor  g17863 ( new_n20212 , new_n20206 , new_n20211 );
xnor g17864 ( n7268 , new_n20204 , new_n20212 );
not  g17865 ( new_n20214 , new_n10789 );
nor  g17866 ( new_n20215 , n752 , new_n20214 );
not  g17867 ( new_n20216 , new_n20215 );
nor  g17868 ( new_n20217 , n2175 , new_n20216 );
not  g17869 ( new_n20218 , new_n20217 );
nor  g17870 ( new_n20219 , n13026 , new_n20218 );
not  g17871 ( new_n20220 , new_n20219 );
nor  g17872 ( new_n20221 , n23912 , new_n20220 );
not  g17873 ( new_n20222 , n10514 );
xnor g17874 ( new_n20223 , n23912 , new_n20219 );
nor  g17875 ( new_n20224 , new_n20222 , new_n20223 );
not  g17876 ( new_n20225 , new_n20223 );
xnor g17877 ( new_n20226 , new_n20222 , new_n20225 );
xnor g17878 ( new_n20227 , n13026 , new_n20217 );
nor  g17879 ( new_n20228 , new_n11276 , new_n20227 );
not  g17880 ( new_n20229 , new_n20227 );
xnor g17881 ( new_n20230 , new_n11276 , new_n20229 );
xnor g17882 ( new_n20231 , n2175 , new_n20215 );
nor  g17883 ( new_n20232 , new_n11389 , new_n20231 );
not  g17884 ( new_n20233 , new_n20231 );
xnor g17885 ( new_n20234 , new_n11389 , new_n20233 );
nor  g17886 ( new_n20235_1 , new_n10824 , new_n10790 );
xnor g17887 ( new_n20236 , n20470 , new_n10790 );
nor  g17888 ( new_n20237 , new_n10837 , new_n10792_1 );
xnor g17889 ( new_n20238 , n21222 , new_n10792_1 );
not  g17890 ( new_n20239 , n9832 );
nor  g17891 ( new_n20240 , new_n20239 , new_n10795 );
xnor g17892 ( new_n20241 , n9832 , new_n10795 );
nor  g17893 ( new_n20242 , new_n9479 , new_n10798 );
xnor g17894 ( new_n20243 , n1558 , new_n10798 );
xnor g17895 ( new_n20244 , n5131 , new_n10782 );
and  g17896 ( new_n20245 , n21749 , new_n20244 );
xnor g17897 ( new_n20246 , n21749 , new_n10800 );
nor  g17898 ( new_n20247 , new_n9487 , new_n10806 );
nor  g17899 ( new_n20248 , n15506 , new_n9485 );
xnor g17900 ( new_n20249 , new_n9487 , new_n10805 );
and  g17901 ( new_n20250_1 , new_n20248 , new_n20249 );
or   g17902 ( new_n20251 , new_n20247 , new_n20250_1 );
and  g17903 ( new_n20252 , new_n20246 , new_n20251 );
or   g17904 ( new_n20253 , new_n20245 , new_n20252 );
and  g17905 ( new_n20254 , new_n20243 , new_n20253 );
or   g17906 ( new_n20255 , new_n20242 , new_n20254 );
and  g17907 ( new_n20256 , new_n20241 , new_n20255 );
or   g17908 ( new_n20257 , new_n20240 , new_n20256 );
and  g17909 ( new_n20258 , new_n20238 , new_n20257 );
or   g17910 ( new_n20259_1 , new_n20237 , new_n20258 );
and  g17911 ( new_n20260 , new_n20236 , new_n20259_1 );
or   g17912 ( new_n20261 , new_n20235_1 , new_n20260 );
and  g17913 ( new_n20262 , new_n20234 , new_n20261 );
or   g17914 ( new_n20263 , new_n20232 , new_n20262 );
and  g17915 ( new_n20264 , new_n20230 , new_n20263 );
or   g17916 ( new_n20265 , new_n20228 , new_n20264 );
and  g17917 ( new_n20266 , new_n20226 , new_n20265 );
nor  g17918 ( new_n20267 , new_n20224 , new_n20266 );
and  g17919 ( new_n20268 , new_n20221 , new_n20267 );
xor  g17920 ( new_n20269 , new_n20226 , new_n20265 );
nor  g17921 ( new_n20270 , n9872 , new_n20269 );
not  g17922 ( new_n20271 , n9872 );
xnor g17923 ( new_n20272 , new_n20271 , new_n20269 );
xor  g17924 ( new_n20273 , new_n20230 , new_n20263 );
nor  g17925 ( new_n20274 , n5842 , new_n20273 );
not  g17926 ( new_n20275 , n5842 );
xnor g17927 ( new_n20276 , new_n20275 , new_n20273 );
xor  g17928 ( new_n20277 , new_n20234 , new_n20261 );
nor  g17929 ( new_n20278 , n6379 , new_n20277 );
not  g17930 ( new_n20279_1 , n6379 );
xnor g17931 ( new_n20280 , new_n20279_1 , new_n20277 );
xor  g17932 ( new_n20281 , new_n20236 , new_n20259_1 );
nor  g17933 ( new_n20282 , n2102 , new_n20281 );
not  g17934 ( new_n20283 , n2102 );
xnor g17935 ( new_n20284 , new_n20283 , new_n20281 );
xor  g17936 ( new_n20285 , new_n20238 , new_n20257 );
nor  g17937 ( new_n20286 , n17954 , new_n20285 );
xor  g17938 ( new_n20287_1 , new_n20241 , new_n20255 );
nor  g17939 ( new_n20288 , n8256 , new_n20287_1 );
not  g17940 ( new_n20289 , n8256 );
xnor g17941 ( new_n20290 , new_n20289 , new_n20287_1 );
xor  g17942 ( new_n20291 , new_n20243 , new_n20253 );
nor  g17943 ( new_n20292 , n24150 , new_n20291 );
not  g17944 ( new_n20293 , n24150 );
xnor g17945 ( new_n20294 , new_n20293 , new_n20291 );
xor  g17946 ( new_n20295 , new_n20246 , new_n20251 );
nor  g17947 ( new_n20296 , n19584 , new_n20295 );
not  g17948 ( new_n20297 , n19584 );
xnor g17949 ( new_n20298 , new_n20297 , new_n20295 );
not  g17950 ( new_n20299 , n5060 );
xnor g17951 ( new_n20300 , new_n20248 , new_n20249 );
nor  g17952 ( new_n20301_1 , new_n20299 , new_n20300 );
not  g17953 ( new_n20302 , new_n20300 );
or   g17954 ( new_n20303 , n5060 , new_n20302 );
xnor g17955 ( new_n20304 , n15506 , n21138 );
and  g17956 ( new_n20305 , n15332 , new_n20304 );
and  g17957 ( new_n20306 , new_n20303 , new_n20305 );
nor  g17958 ( new_n20307 , new_n20301_1 , new_n20306 );
and  g17959 ( new_n20308 , new_n20298 , new_n20307 );
or   g17960 ( new_n20309 , new_n20296 , new_n20308 );
and  g17961 ( new_n20310 , new_n20294 , new_n20309 );
or   g17962 ( new_n20311 , new_n20292 , new_n20310 );
and  g17963 ( new_n20312 , new_n20290 , new_n20311 );
or   g17964 ( new_n20313 , new_n20288 , new_n20312 );
not  g17965 ( new_n20314 , n17954 );
xnor g17966 ( new_n20315 , new_n20314 , new_n20285 );
and  g17967 ( new_n20316 , new_n20313 , new_n20315 );
or   g17968 ( new_n20317 , new_n20286 , new_n20316 );
and  g17969 ( new_n20318 , new_n20284 , new_n20317 );
or   g17970 ( new_n20319 , new_n20282 , new_n20318 );
and  g17971 ( new_n20320 , new_n20280 , new_n20319 );
or   g17972 ( new_n20321 , new_n20278 , new_n20320 );
and  g17973 ( new_n20322 , new_n20276 , new_n20321 );
or   g17974 ( new_n20323 , new_n20274 , new_n20322 );
and  g17975 ( new_n20324 , new_n20272 , new_n20323 );
nor  g17976 ( new_n20325 , new_n20270 , new_n20324 );
not  g17977 ( new_n20326 , new_n20325 );
and  g17978 ( new_n20327 , new_n20268 , new_n20326 );
or   g17979 ( new_n20328 , new_n20221 , new_n20267 );
nor  g17980 ( new_n20329 , new_n20326 , new_n20328 );
nor  g17981 ( new_n20330_1 , new_n20327 , new_n20329 );
xnor g17982 ( new_n20331 , new_n14356 , new_n20330_1 );
not  g17983 ( new_n20332 , new_n20221 );
xnor g17984 ( new_n20333_1 , new_n20332 , new_n20267 );
xnor g17985 ( new_n20334 , new_n20326 , new_n20333_1 );
nor  g17986 ( new_n20335 , new_n14361 , new_n20334 );
xnor g17987 ( new_n20336 , new_n14361 , new_n20334 );
xor  g17988 ( new_n20337 , new_n20272 , new_n20323 );
nor  g17989 ( new_n20338 , new_n2655 , new_n20337 );
xnor g17990 ( new_n20339 , new_n2655 , new_n20337 );
xor  g17991 ( new_n20340 , new_n20276 , new_n20321 );
nor  g17992 ( new_n20341 , new_n2786 , new_n20340 );
xor  g17993 ( new_n20342 , new_n20280 , new_n20319 );
nor  g17994 ( new_n20343 , new_n2792 , new_n20342 );
xnor g17995 ( new_n20344 , new_n2792 , new_n20342 );
xor  g17996 ( new_n20345 , new_n20284 , new_n20317 );
nor  g17997 ( new_n20346 , new_n2797 , new_n20345 );
xnor g17998 ( new_n20347 , new_n2797 , new_n20345 );
xor  g17999 ( new_n20348 , new_n20313 , new_n20315 );
nor  g18000 ( new_n20349_1 , new_n2801 , new_n20348 );
xnor g18001 ( new_n20350 , new_n2801 , new_n20348 );
not  g18002 ( new_n20351 , new_n2806 );
xor  g18003 ( new_n20352 , new_n20290 , new_n20311 );
nor  g18004 ( new_n20353 , new_n20351 , new_n20352 );
xnor g18005 ( new_n20354 , new_n20351 , new_n20352 );
xor  g18006 ( new_n20355_1 , new_n20294 , new_n20309 );
nor  g18007 ( new_n20356 , new_n2812 , new_n20355_1 );
xnor g18008 ( new_n20357 , new_n2812 , new_n20355_1 );
xor  g18009 ( new_n20358 , new_n20298 , new_n20307 );
nor  g18010 ( new_n20359_1 , new_n2818 , new_n20358 );
xnor g18011 ( new_n20360 , new_n2818 , new_n20358 );
xnor g18012 ( new_n20361 , new_n20299 , new_n20302 );
xnor g18013 ( new_n20362 , new_n20305 , new_n20361 );
nor  g18014 ( new_n20363 , new_n2824 , new_n20362 );
xnor g18015 ( new_n20364 , new_n16103 , new_n20304 );
nor  g18016 ( new_n20365 , new_n2827 , new_n20364 );
xnor g18017 ( new_n20366_1 , new_n2824 , new_n20362 );
nor  g18018 ( new_n20367 , new_n20365 , new_n20366_1 );
nor  g18019 ( new_n20368 , new_n20363 , new_n20367 );
nor  g18020 ( new_n20369 , new_n20360 , new_n20368 );
nor  g18021 ( new_n20370 , new_n20359_1 , new_n20369 );
nor  g18022 ( new_n20371 , new_n20357 , new_n20370 );
nor  g18023 ( new_n20372 , new_n20356 , new_n20371 );
nor  g18024 ( new_n20373 , new_n20354 , new_n20372 );
nor  g18025 ( new_n20374 , new_n20353 , new_n20373 );
nor  g18026 ( new_n20375 , new_n20350 , new_n20374 );
nor  g18027 ( new_n20376 , new_n20349_1 , new_n20375 );
nor  g18028 ( new_n20377 , new_n20347 , new_n20376 );
nor  g18029 ( new_n20378 , new_n20346 , new_n20377 );
nor  g18030 ( new_n20379 , new_n20344 , new_n20378 );
nor  g18031 ( new_n20380 , new_n20343 , new_n20379 );
xnor g18032 ( new_n20381 , new_n2786 , new_n20340 );
nor  g18033 ( new_n20382 , new_n20380 , new_n20381 );
nor  g18034 ( new_n20383 , new_n20341 , new_n20382 );
nor  g18035 ( new_n20384 , new_n20339 , new_n20383 );
nor  g18036 ( new_n20385_1 , new_n20338 , new_n20384 );
nor  g18037 ( new_n20386 , new_n20336 , new_n20385_1 );
nor  g18038 ( new_n20387 , new_n20335 , new_n20386 );
xnor g18039 ( n7277 , new_n20331 , new_n20387 );
xor  g18040 ( n7280 , new_n13126 , new_n13133 );
xnor g18041 ( n7298 , new_n5728 , new_n5753 );
xnor g18042 ( n7308 , new_n18910 , new_n18919_1 );
xnor g18043 ( new_n20392 , new_n7242 , new_n19135 );
nor  g18044 ( new_n20393 , new_n7266 , new_n19141_1 );
xnor g18045 ( new_n20394 , new_n7266 , new_n19138 );
nor  g18046 ( new_n20395 , new_n14628 , new_n14653 );
nor  g18047 ( new_n20396 , new_n14654 , new_n14680_1 );
or   g18048 ( new_n20397 , new_n20395 , new_n20396 );
and  g18049 ( new_n20398 , new_n20394 , new_n20397 );
nor  g18050 ( new_n20399 , new_n20393 , new_n20398 );
xnor g18051 ( new_n20400 , new_n20392 , new_n20399 );
not  g18052 ( new_n20401 , new_n20400 );
xnor g18053 ( new_n20402_1 , new_n19163_1 , new_n20401 );
xor  g18054 ( new_n20403_1 , new_n20394 , new_n20397 );
nor  g18055 ( new_n20404 , new_n19169 , new_n20403_1 );
and  g18056 ( new_n20405 , new_n14682 , new_n18560 );
and  g18057 ( new_n20406 , new_n18561 , new_n18590 );
nor  g18058 ( new_n20407 , new_n20405 , new_n20406 );
xnor g18059 ( new_n20408 , new_n19169 , new_n20403_1 );
not  g18060 ( new_n20409_1 , new_n20408 );
and  g18061 ( new_n20410 , new_n20407 , new_n20409_1 );
nor  g18062 ( new_n20411_1 , new_n20404 , new_n20410 );
xnor g18063 ( n7313 , new_n20402_1 , new_n20411_1 );
xnor g18064 ( n7346 , new_n3689 , new_n3713 );
xnor g18065 ( new_n20414 , new_n13735 , new_n20086_1 );
nor  g18066 ( new_n20415 , new_n13739 , new_n20086_1 );
xnor g18067 ( new_n20416 , new_n13739 , new_n20086_1 );
nor  g18068 ( new_n20417 , new_n11203 , new_n13743 );
xnor g18069 ( new_n20418 , new_n11203 , new_n13743 );
nor  g18070 ( new_n20419 , new_n11206 , new_n13747 );
xnor g18071 ( new_n20420 , new_n11206 , new_n13747 );
nor  g18072 ( new_n20421 , new_n11210 , new_n13752 );
nor  g18073 ( new_n20422 , new_n6431_1 , new_n6551 );
and  g18074 ( new_n20423 , new_n6553 , new_n6583 );
nor  g18075 ( new_n20424_1 , new_n20422 , new_n20423 );
xnor g18076 ( new_n20425 , new_n11210 , new_n13751 );
and  g18077 ( new_n20426 , new_n20424_1 , new_n20425 );
nor  g18078 ( new_n20427 , new_n20421 , new_n20426 );
nor  g18079 ( new_n20428 , new_n20420 , new_n20427 );
nor  g18080 ( new_n20429_1 , new_n20419 , new_n20428 );
nor  g18081 ( new_n20430 , new_n20418 , new_n20429_1 );
nor  g18082 ( new_n20431 , new_n20417 , new_n20430 );
nor  g18083 ( new_n20432 , new_n20416 , new_n20431 );
nor  g18084 ( new_n20433 , new_n20415 , new_n20432 );
xor  g18085 ( n7349 , new_n20414 , new_n20433 );
xnor g18086 ( n7363 , new_n20339 , new_n20383 );
nor  g18087 ( new_n20436_1 , new_n8954 , n21839 );
and  g18088 ( new_n20437 , new_n19110 , new_n19113 );
nor  g18089 ( new_n20438 , new_n20436_1 , new_n20437 );
xnor g18090 ( new_n20439 , new_n10099 , new_n20438 );
nor  g18091 ( new_n20440 , new_n10102 , new_n19114 );
nor  g18092 ( new_n20441_1 , new_n19115 , new_n19118 );
nor  g18093 ( new_n20442 , new_n20440 , new_n20441_1 );
xnor g18094 ( n7390 , new_n20439 , new_n20442 );
xnor g18095 ( n7403 , new_n9044 , new_n9045 );
xnor g18096 ( n7408 , new_n9182_1 , new_n9219 );
xnor g18097 ( n7432 , new_n19426 , new_n19449 );
nor  g18098 ( new_n20447 , new_n15098 , new_n17497 );
nor  g18099 ( new_n20448 , new_n17499 , new_n17507 );
or   g18100 ( n7475 , new_n20447 , new_n20448 );
xnor g18101 ( n7477 , new_n5208 , new_n5209 );
xnor g18102 ( n7507 , new_n8874 , new_n8899 );
nor  g18103 ( new_n20452 , new_n5453 , new_n11803 );
xnor g18104 ( new_n20453 , new_n5453 , new_n11802 );
nor  g18105 ( new_n20454 , new_n5456 , new_n6863_1 );
and  g18106 ( new_n20455_1 , new_n6865 , new_n6908 );
or   g18107 ( new_n20456 , new_n20454 , new_n20455_1 );
and  g18108 ( new_n20457 , new_n20453 , new_n20456 );
nor  g18109 ( new_n20458 , new_n20452 , new_n20457 );
xnor g18110 ( new_n20459 , new_n11851 , new_n20458 );
xnor g18111 ( new_n20460 , new_n16853 , new_n20459 );
xor  g18112 ( new_n20461 , new_n20453 , new_n20456 );
nor  g18113 ( new_n20462 , new_n16857 , new_n20461 );
xnor g18114 ( new_n20463 , new_n16857 , new_n20461 );
nor  g18115 ( new_n20464 , new_n6833 , new_n6909 );
nor  g18116 ( new_n20465 , new_n6910 , new_n6964 );
nor  g18117 ( new_n20466 , new_n20464 , new_n20465 );
nor  g18118 ( new_n20467 , new_n20463 , new_n20466 );
nor  g18119 ( new_n20468 , new_n20462 , new_n20467 );
xnor g18120 ( n7514 , new_n20460 , new_n20468 );
xnor g18121 ( n7558 , new_n10744 , new_n10767 );
xnor g18122 ( n7572 , new_n11885 , new_n11886 );
xnor g18123 ( new_n20472 , new_n4015 , new_n6274 );
nor  g18124 ( new_n20473 , new_n4021 , new_n6276_1 );
and  g18125 ( new_n20474 , new_n19470 , new_n19479 );
or   g18126 ( new_n20475 , new_n20473 , new_n20474 );
xor  g18127 ( new_n20476 , new_n20472 , new_n20475 );
xnor g18128 ( new_n20477 , new_n9668 , new_n20476 );
nor  g18129 ( new_n20478_1 , new_n9673 , new_n19480 );
nor  g18130 ( new_n20479 , new_n19481 , new_n19492 );
nor  g18131 ( new_n20480 , new_n20478_1 , new_n20479 );
xnor g18132 ( n7575 , new_n20477 , new_n20480 );
xnor g18133 ( new_n20482 , new_n9600 , new_n20229 );
nor  g18134 ( new_n20483 , new_n9652 , new_n20233 );
xnor g18135 ( new_n20484 , new_n9652 , new_n20233 );
and  g18136 ( new_n20485 , new_n9657 , new_n10790 );
and  g18137 ( new_n20486 , new_n10791 , new_n10822 );
nor  g18138 ( new_n20487 , new_n20485 , new_n20486 );
nor  g18139 ( new_n20488 , new_n20484 , new_n20487 );
nor  g18140 ( new_n20489_1 , new_n20483 , new_n20488 );
xnor g18141 ( new_n20490_1 , new_n20482 , new_n20489_1 );
xnor g18142 ( new_n20491 , new_n11384 , new_n20490_1 );
xnor g18143 ( new_n20492 , new_n20484 , new_n20487 );
nor  g18144 ( new_n20493 , new_n11392 , new_n20492 );
xnor g18145 ( new_n20494 , new_n11392 , new_n20492 );
nor  g18146 ( new_n20495_1 , new_n10823 , new_n10834_1 );
nor  g18147 ( new_n20496 , new_n10835 , new_n10868 );
or   g18148 ( new_n20497 , new_n20495_1 , new_n20496 );
nor  g18149 ( new_n20498 , new_n20494 , new_n20497 );
nor  g18150 ( new_n20499 , new_n20493 , new_n20498 );
xor  g18151 ( n7585 , new_n20491 , new_n20499 );
not  g18152 ( new_n20501 , new_n19947 );
xnor g18153 ( new_n20502 , new_n7698_1 , new_n20501 );
nor  g18154 ( new_n20503 , new_n7705 , new_n19950 );
xnor g18155 ( new_n20504 , new_n7705 , new_n19950 );
nor  g18156 ( new_n20505 , new_n7710 , new_n19954 );
xnor g18157 ( new_n20506 , new_n7714 , new_n19956 );
nor  g18158 ( new_n20507 , new_n7717 , new_n19960 );
xnor g18159 ( new_n20508 , new_n7717 , new_n19960 );
nor  g18160 ( new_n20509 , new_n7721_1 , new_n19963 );
xnor g18161 ( new_n20510 , new_n7721_1 , new_n19963 );
nor  g18162 ( new_n20511 , new_n7725 , new_n17591 );
xnor g18163 ( new_n20512 , new_n7725 , new_n17591 );
nor  g18164 ( new_n20513 , new_n7730 , new_n17594 );
xnor g18165 ( new_n20514 , new_n7729 , new_n17595 );
not  g18166 ( new_n20515_1 , new_n17599 );
nor  g18167 ( new_n20516 , new_n7739 , new_n20515_1 );
xnor g18168 ( new_n20517 , new_n7739 , new_n20515_1 );
nor  g18169 ( new_n20518 , new_n7748 , new_n17605 );
nor  g18170 ( new_n20519 , new_n7743 , new_n20518 );
xnor g18171 ( new_n20520 , new_n7742 , new_n20518 );
and  g18172 ( new_n20521 , new_n17611 , new_n20520 );
nor  g18173 ( new_n20522 , new_n20519 , new_n20521 );
nor  g18174 ( new_n20523 , new_n20517 , new_n20522 );
nor  g18175 ( new_n20524 , new_n20516 , new_n20523 );
nor  g18176 ( new_n20525 , new_n20514 , new_n20524 );
nor  g18177 ( new_n20526 , new_n20513 , new_n20525 );
nor  g18178 ( new_n20527 , new_n20512 , new_n20526 );
nor  g18179 ( new_n20528 , new_n20511 , new_n20527 );
nor  g18180 ( new_n20529 , new_n20510 , new_n20528 );
nor  g18181 ( new_n20530 , new_n20509 , new_n20529 );
nor  g18182 ( new_n20531 , new_n20508 , new_n20530 );
nor  g18183 ( new_n20532 , new_n20507 , new_n20531 );
nor  g18184 ( new_n20533_1 , new_n20506 , new_n20532 );
nor  g18185 ( new_n20534 , new_n20505 , new_n20533_1 );
nor  g18186 ( new_n20535 , new_n20504 , new_n20534 );
nor  g18187 ( new_n20536 , new_n20503 , new_n20535 );
xnor g18188 ( n7588 , new_n20502 , new_n20536 );
not  g18189 ( new_n20538 , new_n6679 );
nor  g18190 ( new_n20539 , n21832 , new_n20538 );
not  g18191 ( new_n20540 , new_n20539 );
nor  g18192 ( new_n20541 , n21753 , new_n20540 );
not  g18193 ( new_n20542 , new_n20541 );
nor  g18194 ( new_n20543 , n10739 , new_n20542 );
not  g18195 ( new_n20544 , new_n20543 );
nor  g18196 ( new_n20545 , n13074 , new_n20544 );
xnor g18197 ( new_n20546 , n23463 , new_n20545 );
not  g18198 ( new_n20547 , new_n20546 );
xnor g18199 ( new_n20548 , n23250 , new_n20547 );
xnor g18200 ( new_n20549 , n13074 , new_n20543 );
nor  g18201 ( new_n20550 , n11455 , new_n20549 );
not  g18202 ( new_n20551 , new_n20549 );
xnor g18203 ( new_n20552 , n11455 , new_n20551 );
xnor g18204 ( new_n20553 , n10739 , new_n20541 );
nor  g18205 ( new_n20554 , n3945 , new_n20553 );
xnor g18206 ( new_n20555 , new_n15602_1 , new_n20553 );
xnor g18207 ( new_n20556 , n21753 , new_n20539 );
nor  g18208 ( new_n20557 , n5255 , new_n20556 );
not  g18209 ( new_n20558 , new_n20556 );
xnor g18210 ( new_n20559 , n5255 , new_n20558 );
nor  g18211 ( new_n20560 , n21649 , new_n6680 );
xnor g18212 ( new_n20561 , new_n5163 , new_n6680 );
nor  g18213 ( new_n20562 , n18274 , new_n6698 );
nor  g18214 ( new_n20563 , n3828 , new_n6711 );
xnor g18215 ( new_n20564 , n3828 , new_n6712 );
nor  g18216 ( new_n20565 , n23842 , new_n6706_1 );
or   g18217 ( new_n20566 , new_n3116 , new_n15011_1 );
xnor g18218 ( new_n20567 , new_n5172 , new_n6706_1 );
and  g18219 ( new_n20568 , new_n20566 , new_n20567 );
or   g18220 ( new_n20569 , new_n20565 , new_n20568 );
and  g18221 ( new_n20570 , new_n20564 , new_n20569 );
or   g18222 ( new_n20571 , new_n20563 , new_n20570 );
xnor g18223 ( new_n20572 , new_n5166 , new_n6698 );
and  g18224 ( new_n20573 , new_n20571 , new_n20572 );
or   g18225 ( new_n20574 , new_n20562 , new_n20573 );
and  g18226 ( new_n20575 , new_n20561 , new_n20574 );
or   g18227 ( new_n20576 , new_n20560 , new_n20575 );
and  g18228 ( new_n20577 , new_n20559 , new_n20576 );
or   g18229 ( new_n20578 , new_n20557 , new_n20577 );
and  g18230 ( new_n20579 , new_n20555 , new_n20578 );
or   g18231 ( new_n20580 , new_n20554 , new_n20579 );
and  g18232 ( new_n20581 , new_n20552 , new_n20580 );
or   g18233 ( new_n20582_1 , new_n20550 , new_n20581 );
xor  g18234 ( new_n20583 , new_n20548 , new_n20582_1 );
xnor g18235 ( new_n20584 , new_n14074 , new_n20583 );
xor  g18236 ( new_n20585 , new_n20552 , new_n20580 );
and  g18237 ( new_n20586 , new_n14108 , new_n20585 );
xnor g18238 ( new_n20587 , new_n14112 , new_n20585 );
xor  g18239 ( new_n20588 , new_n20555 , new_n20578 );
nor  g18240 ( new_n20589 , new_n14116 , new_n20588 );
xnor g18241 ( new_n20590_1 , new_n14115 , new_n20588 );
xor  g18242 ( new_n20591 , new_n20559 , new_n20576 );
nor  g18243 ( new_n20592 , new_n14122 , new_n20591 );
xor  g18244 ( new_n20593 , new_n20561 , new_n20574 );
nor  g18245 ( new_n20594 , new_n14125 , new_n20593 );
xor  g18246 ( new_n20595 , new_n20571 , new_n20572 );
nor  g18247 ( new_n20596 , new_n14130_1 , new_n20595 );
xnor g18248 ( new_n20597 , new_n14129 , new_n20595 );
xor  g18249 ( new_n20598 , new_n20564 , new_n20569 );
nor  g18250 ( new_n20599 , new_n14136_1 , new_n20598 );
xnor g18251 ( new_n20600 , new_n14135 , new_n20598 );
nor  g18252 ( new_n20601 , new_n14140 , new_n20567 );
xor  g18253 ( new_n20602_1 , new_n20566 , new_n20567 );
nor  g18254 ( new_n20603 , new_n14139 , new_n20602_1 );
xnor g18255 ( new_n20604_1 , n2387 , n21654 );
nor  g18256 ( new_n20605 , new_n14146 , new_n20604_1 );
nor  g18257 ( new_n20606 , new_n20603 , new_n20605 );
nor  g18258 ( new_n20607 , new_n20601 , new_n20606 );
and  g18259 ( new_n20608 , new_n20600 , new_n20607 );
or   g18260 ( new_n20609_1 , new_n20599 , new_n20608 );
and  g18261 ( new_n20610 , new_n20597 , new_n20609_1 );
nor  g18262 ( new_n20611 , new_n20596 , new_n20610 );
xnor g18263 ( new_n20612 , new_n14125 , new_n20593 );
nor  g18264 ( new_n20613 , new_n20611 , new_n20612 );
or   g18265 ( new_n20614 , new_n20594 , new_n20613 );
xnor g18266 ( new_n20615 , new_n14120 , new_n20591 );
and  g18267 ( new_n20616 , new_n20614 , new_n20615 );
or   g18268 ( new_n20617 , new_n20592 , new_n20616 );
and  g18269 ( new_n20618 , new_n20590_1 , new_n20617 );
nor  g18270 ( new_n20619 , new_n20589 , new_n20618 );
and  g18271 ( new_n20620 , new_n20587 , new_n20619 );
nor  g18272 ( new_n20621 , new_n20586 , new_n20620 );
xor  g18273 ( n7598 , new_n20584 , new_n20621 );
xnor g18274 ( n7607 , new_n17502 , new_n17505 );
xnor g18275 ( n7610 , new_n4991 , new_n5016 );
xnor g18276 ( n7616 , new_n3366_1 , new_n3377 );
xnor g18277 ( new_n20626 , n6105 , n10514 );
nor  g18278 ( new_n20627 , n3795 , n18649 );
xnor g18279 ( new_n20628 , n3795 , n18649 );
nor  g18280 ( new_n20629_1 , n6218 , n25464 );
xnor g18281 ( new_n20630 , n6218 , n25464 );
nor  g18282 ( new_n20631 , n4590 , n20470 );
xnor g18283 ( new_n20632 , n4590 , n20470 );
nor  g18284 ( new_n20633 , n21222 , n26752 );
xnor g18285 ( new_n20634 , n21222 , n26752 );
nor  g18286 ( new_n20635 , n6513 , n9832 );
xnor g18287 ( new_n20636 , new_n6334 , n9832 );
nor  g18288 ( new_n20637 , new_n9479 , new_n6336 );
or   g18289 ( new_n20638 , n1558 , n3918 );
nor  g18290 ( new_n20639 , n919 , n21749 );
nor  g18291 ( new_n20640 , new_n16095 , new_n16100 );
nor  g18292 ( new_n20641 , new_n20639 , new_n20640 );
and  g18293 ( new_n20642 , new_n20638 , new_n20641 );
nor  g18294 ( new_n20643 , new_n20637 , new_n20642 );
and  g18295 ( new_n20644 , new_n20636 , new_n20643 );
nor  g18296 ( new_n20645 , new_n20635 , new_n20644 );
nor  g18297 ( new_n20646 , new_n20634 , new_n20645 );
nor  g18298 ( new_n20647 , new_n20633 , new_n20646 );
nor  g18299 ( new_n20648 , new_n20632 , new_n20647 );
nor  g18300 ( new_n20649 , new_n20631 , new_n20648 );
nor  g18301 ( new_n20650 , new_n20630 , new_n20649 );
nor  g18302 ( new_n20651 , new_n20629_1 , new_n20650 );
nor  g18303 ( new_n20652 , new_n20628 , new_n20651 );
nor  g18304 ( new_n20653 , new_n20627 , new_n20652 );
xnor g18305 ( new_n20654 , new_n20626 , new_n20653 );
nor  g18306 ( new_n20655 , new_n20271 , new_n20654 );
xnor g18307 ( new_n20656 , new_n20271 , new_n20654 );
xnor g18308 ( new_n20657 , new_n20628 , new_n20651 );
nor  g18309 ( new_n20658_1 , new_n20275 , new_n20657 );
xnor g18310 ( new_n20659 , new_n20275 , new_n20657 );
xnor g18311 ( new_n20660 , new_n20630 , new_n20649 );
nor  g18312 ( new_n20661_1 , new_n20279_1 , new_n20660 );
xnor g18313 ( new_n20662 , new_n20279_1 , new_n20660 );
xnor g18314 ( new_n20663 , new_n20632 , new_n20647 );
nor  g18315 ( new_n20664 , new_n20283 , new_n20663 );
xnor g18316 ( new_n20665 , new_n20283 , new_n20663 );
xnor g18317 ( new_n20666 , new_n20634 , new_n20645 );
nor  g18318 ( new_n20667 , new_n20314 , new_n20666 );
xnor g18319 ( new_n20668 , new_n20314 , new_n20666 );
xnor g18320 ( new_n20669 , new_n20636 , new_n20643 );
nor  g18321 ( new_n20670 , new_n20289 , new_n20669 );
xnor g18322 ( new_n20671 , new_n20289 , new_n20669 );
xnor g18323 ( new_n20672 , n1558 , n3918 );
xnor g18324 ( new_n20673_1 , new_n20641 , new_n20672 );
nor  g18325 ( new_n20674 , new_n20293 , new_n20673_1 );
xnor g18326 ( new_n20675 , n24150 , new_n20673_1 );
nor  g18327 ( new_n20676 , new_n20297 , new_n16101 );
and  g18328 ( new_n20677 , new_n16102 , new_n16110_1 );
or   g18329 ( new_n20678_1 , new_n20676 , new_n20677 );
and  g18330 ( new_n20679 , new_n20675 , new_n20678_1 );
nor  g18331 ( new_n20680_1 , new_n20674 , new_n20679 );
nor  g18332 ( new_n20681 , new_n20671 , new_n20680_1 );
nor  g18333 ( new_n20682 , new_n20670 , new_n20681 );
nor  g18334 ( new_n20683 , new_n20668 , new_n20682 );
nor  g18335 ( new_n20684 , new_n20667 , new_n20683 );
nor  g18336 ( new_n20685_1 , new_n20665 , new_n20684 );
nor  g18337 ( new_n20686 , new_n20664 , new_n20685_1 );
nor  g18338 ( new_n20687 , new_n20662 , new_n20686 );
nor  g18339 ( new_n20688 , new_n20661_1 , new_n20687 );
nor  g18340 ( new_n20689 , new_n20659 , new_n20688 );
nor  g18341 ( new_n20690 , new_n20658_1 , new_n20689 );
nor  g18342 ( new_n20691_1 , new_n20656 , new_n20690 );
nor  g18343 ( new_n20692 , new_n20655 , new_n20691_1 );
nor  g18344 ( new_n20693 , n6105 , n10514 );
nor  g18345 ( new_n20694 , new_n20626 , new_n20653 );
nor  g18346 ( new_n20695 , new_n20693 , new_n20694 );
nor  g18347 ( new_n20696_1 , new_n20692 , new_n20695 );
xnor g18348 ( new_n20697 , new_n15335 , new_n20696_1 );
xnor g18349 ( new_n20698 , new_n20692 , new_n20695 );
nor  g18350 ( new_n20699 , new_n15227 , new_n20698 );
xnor g18351 ( new_n20700_1 , new_n15227 , new_n20698 );
xnor g18352 ( new_n20701 , new_n20656 , new_n20690 );
nor  g18353 ( new_n20702 , new_n15270 , new_n20701 );
xnor g18354 ( new_n20703 , new_n15270 , new_n20701 );
xnor g18355 ( new_n20704_1 , new_n20659 , new_n20688 );
nor  g18356 ( new_n20705_1 , new_n15274 , new_n20704_1 );
xnor g18357 ( new_n20706 , new_n15274 , new_n20704_1 );
xnor g18358 ( new_n20707 , new_n20662 , new_n20686 );
nor  g18359 ( new_n20708 , new_n15278 , new_n20707 );
xnor g18360 ( new_n20709_1 , new_n15278 , new_n20707 );
xnor g18361 ( new_n20710 , new_n20665 , new_n20684 );
nor  g18362 ( new_n20711 , new_n15282 , new_n20710 );
xnor g18363 ( new_n20712 , new_n15282 , new_n20710 );
xnor g18364 ( new_n20713_1 , new_n20668 , new_n20682 );
nor  g18365 ( new_n20714 , new_n15286 , new_n20713_1 );
xnor g18366 ( new_n20715 , new_n15286 , new_n20713_1 );
xnor g18367 ( new_n20716 , new_n20671 , new_n20680_1 );
nor  g18368 ( new_n20717 , new_n15291 , new_n20716 );
xnor g18369 ( new_n20718 , new_n15291 , new_n20716 );
xor  g18370 ( new_n20719 , new_n20675 , new_n20678_1 );
and  g18371 ( new_n20720 , new_n15296 , new_n20719 );
xnor g18372 ( new_n20721 , new_n15296 , new_n20719 );
nor  g18373 ( new_n20722_1 , new_n15301 , new_n16111 );
nor  g18374 ( new_n20723_1 , new_n16112 , new_n16119 );
nor  g18375 ( new_n20724 , new_n20722_1 , new_n20723_1 );
nor  g18376 ( new_n20725 , new_n20721 , new_n20724 );
nor  g18377 ( new_n20726 , new_n20720 , new_n20725 );
nor  g18378 ( new_n20727 , new_n20718 , new_n20726 );
nor  g18379 ( new_n20728 , new_n20717 , new_n20727 );
nor  g18380 ( new_n20729 , new_n20715 , new_n20728 );
nor  g18381 ( new_n20730 , new_n20714 , new_n20729 );
nor  g18382 ( new_n20731 , new_n20712 , new_n20730 );
nor  g18383 ( new_n20732 , new_n20711 , new_n20731 );
nor  g18384 ( new_n20733 , new_n20709_1 , new_n20732 );
nor  g18385 ( new_n20734 , new_n20708 , new_n20733 );
nor  g18386 ( new_n20735 , new_n20706 , new_n20734 );
nor  g18387 ( new_n20736 , new_n20705_1 , new_n20735 );
nor  g18388 ( new_n20737 , new_n20703 , new_n20736 );
nor  g18389 ( new_n20738 , new_n20702 , new_n20737 );
nor  g18390 ( new_n20739 , new_n20700_1 , new_n20738 );
nor  g18391 ( new_n20740 , new_n20699 , new_n20739 );
xnor g18392 ( n7630 , new_n20697 , new_n20740 );
nor  g18393 ( new_n20742 , new_n18300 , new_n18324 );
nor  g18394 ( new_n20743 , new_n18325 , new_n18333 );
nor  g18395 ( n7643 , new_n20742 , new_n20743 );
xnor g18396 ( n7647 , new_n11987 , new_n12010 );
xnor g18397 ( n7679 , new_n9941 , new_n9974 );
xnor g18398 ( n7686 , new_n19629 , new_n19651 );
xnor g18399 ( new_n20748_1 , new_n17816 , new_n17857 );
xnor g18400 ( n7698 , new_n17855_1 , new_n20748_1 );
xnor g18401 ( n7708 , new_n18906 , new_n18921 );
not  g18402 ( new_n20751 , n3324 );
xnor g18403 ( new_n20752 , new_n20751 , new_n17831 );
nor  g18404 ( new_n20753 , new_n19668 , new_n2925 );
xnor g18405 ( new_n20754 , n17911 , new_n2925 );
nor  g18406 ( new_n20755 , n21997 , new_n2976 );
xnor g18407 ( new_n20756 , new_n18472 , new_n2976 );
nor  g18408 ( new_n20757 , n25119 , new_n2980 );
and  g18409 ( new_n20758 , new_n8502 , new_n8526_1 );
or   g18410 ( new_n20759 , new_n20757 , new_n20758 );
and  g18411 ( new_n20760 , new_n20756 , new_n20759 );
nor  g18412 ( new_n20761_1 , new_n20755 , new_n20760 );
and  g18413 ( new_n20762 , new_n20754 , new_n20761_1 );
nor  g18414 ( new_n20763 , new_n20753 , new_n20762 );
xnor g18415 ( new_n20764 , new_n20752 , new_n20763 );
xnor g18416 ( new_n20765 , new_n4907 , new_n6023 );
nor  g18417 ( new_n20766 , n2858 , new_n6029 );
and  g18418 ( new_n20767 , new_n15874 , new_n15882 );
nor  g18419 ( new_n20768 , new_n20766 , new_n20767 );
xnor g18420 ( new_n20769 , new_n20765 , new_n20768 );
xnor g18421 ( new_n20770 , new_n20764 , new_n20769 );
not  g18422 ( new_n20771 , new_n15883 );
xor  g18423 ( new_n20772 , new_n20754 , new_n20761_1 );
nor  g18424 ( new_n20773 , new_n20771 , new_n20772 );
xnor g18425 ( new_n20774_1 , new_n20771 , new_n20772 );
xor  g18426 ( new_n20775 , new_n20756 , new_n20759 );
and  g18427 ( new_n20776 , new_n15885_1 , new_n20775 );
xnor g18428 ( new_n20777 , new_n15885_1 , new_n20775 );
nor  g18429 ( new_n20778 , new_n8500 , new_n8527 );
nor  g18430 ( new_n20779 , new_n8528 , new_n8570 );
nor  g18431 ( new_n20780 , new_n20778 , new_n20779 );
nor  g18432 ( new_n20781 , new_n20777 , new_n20780 );
nor  g18433 ( new_n20782 , new_n20776 , new_n20781 );
nor  g18434 ( new_n20783 , new_n20774_1 , new_n20782 );
nor  g18435 ( new_n20784 , new_n20773 , new_n20783 );
xnor g18436 ( n7780 , new_n20770 , new_n20784 );
nor  g18437 ( new_n20786 , new_n4471 , new_n2603 );
xnor g18438 ( new_n20787 , new_n4471 , new_n2603 );
nor  g18439 ( new_n20788_1 , new_n4431 , new_n2607 );
nor  g18440 ( new_n20789 , new_n9569 , new_n9598_1 );
nor  g18441 ( new_n20790 , new_n20788_1 , new_n20789 );
nor  g18442 ( new_n20791 , new_n20787 , new_n20790 );
nor  g18443 ( new_n20792 , new_n20786 , new_n20791 );
xnor g18444 ( new_n20793 , new_n14355 , new_n20792 );
not  g18445 ( new_n20794_1 , new_n20793 );
nor  g18446 ( new_n20795_1 , new_n10052 , new_n16940 );
xnor g18447 ( new_n20796 , new_n10052 , new_n16939 );
and  g18448 ( new_n20797 , new_n2723 , new_n9611 );
and  g18449 ( new_n20798 , new_n9612 , new_n9648_1 );
or   g18450 ( new_n20799 , new_n20797 , new_n20798 );
and  g18451 ( new_n20800 , new_n20796 , new_n20799 );
nor  g18452 ( new_n20801 , new_n20795_1 , new_n20800 );
not  g18453 ( new_n20802 , new_n20801 );
and  g18454 ( new_n20803_1 , new_n4312 , new_n16938 );
xnor g18455 ( new_n20804 , new_n10049 , new_n20803_1 );
xnor g18456 ( new_n20805 , new_n20802 , new_n20804 );
xnor g18457 ( new_n20806 , new_n20794_1 , new_n20805 );
xor  g18458 ( new_n20807 , new_n20787 , new_n20790 );
xor  g18459 ( new_n20808 , new_n20796 , new_n20799 );
nor  g18460 ( new_n20809 , new_n20807 , new_n20808 );
xnor g18461 ( new_n20810 , new_n20807 , new_n20808 );
nor  g18462 ( new_n20811 , new_n9599 , new_n9649 );
and  g18463 ( new_n20812 , new_n9650 , new_n9703 );
nor  g18464 ( new_n20813 , new_n20811 , new_n20812 );
nor  g18465 ( new_n20814 , new_n20810 , new_n20813 );
nor  g18466 ( new_n20815 , new_n20809 , new_n20814 );
xnor g18467 ( n7794 , new_n20806 , new_n20815 );
xnor g18468 ( n7811 , new_n17113 , new_n17118 );
xor  g18469 ( n7830 , new_n17061 , new_n17066 );
xnor g18470 ( n7834 , new_n20506 , new_n20532 );
xnor g18471 ( n7884 , new_n10850 , new_n10862 );
xnor g18472 ( n7937 , new_n3069 , new_n3070 );
xnor g18473 ( n7943 , new_n3037 , new_n3082 );
xor  g18474 ( n7950 , new_n9666 , new_n9697 );
xnor g18475 ( new_n20824 , new_n15180_1 , new_n19167 );
nor  g18476 ( new_n20825 , new_n15184 , new_n19170 );
nor  g18477 ( new_n20826_1 , new_n15189 , new_n19173 );
xnor g18478 ( new_n20827 , new_n15189 , new_n19173 );
nor  g18479 ( new_n20828 , new_n14886 , new_n15192 );
nor  g18480 ( new_n20829 , new_n14933 , new_n14979 );
nor  g18481 ( new_n20830 , new_n20828 , new_n20829 );
nor  g18482 ( new_n20831 , new_n20827 , new_n20830 );
nor  g18483 ( new_n20832 , new_n20826_1 , new_n20831 );
xnor g18484 ( new_n20833 , new_n15182_1 , new_n19181 );
nor  g18485 ( new_n20834 , new_n20832 , new_n20833 );
nor  g18486 ( new_n20835 , new_n20825 , new_n20834 );
xor  g18487 ( n7959 , new_n20824 , new_n20835 );
xnor g18488 ( n7968 , new_n17109 , new_n17122 );
xnor g18489 ( n7992 , new_n18070 , new_n18071_1 );
xnor g18490 ( new_n20839 , n9554 , new_n12681 );
nor  g18491 ( new_n20840 , new_n7773_1 , new_n12685 );
xnor g18492 ( new_n20841 , new_n7773_1 , new_n12687 );
nor  g18493 ( new_n20842 , n18227 , new_n10450 );
and  g18494 ( new_n20843 , new_n17082 , new_n17094 );
nor  g18495 ( new_n20844 , new_n20842 , new_n20843 );
and  g18496 ( new_n20845 , new_n20841 , new_n20844 );
nor  g18497 ( new_n20846 , new_n20840 , new_n20845 );
xnor g18498 ( new_n20847 , new_n20839 , new_n20846 );
xnor g18499 ( new_n20848 , new_n18231 , new_n20847 );
xnor g18500 ( new_n20849 , new_n20841 , new_n20844 );
nor  g18501 ( new_n20850 , new_n18235 , new_n20849 );
not  g18502 ( new_n20851 , new_n20849 );
xnor g18503 ( new_n20852 , new_n18236 , new_n20851 );
nor  g18504 ( new_n20853 , new_n17096 , new_n18240 );
xnor g18505 ( new_n20854 , new_n17095_1 , new_n18241_1 );
nor  g18506 ( new_n20855 , new_n17100 , new_n18245 );
xnor g18507 ( new_n20856 , new_n17099 , new_n18246 );
and  g18508 ( new_n20857 , new_n17104_1 , new_n18251 );
xnor g18509 ( new_n20858 , new_n17104_1 , new_n18251 );
nor  g18510 ( new_n20859 , new_n17107 , new_n12769 );
nor  g18511 ( new_n20860 , new_n12771 , new_n12774 );
nor  g18512 ( new_n20861 , new_n20859 , new_n20860 );
nor  g18513 ( new_n20862 , new_n20858 , new_n20861 );
nor  g18514 ( new_n20863 , new_n20857 , new_n20862 );
nor  g18515 ( new_n20864 , new_n20856 , new_n20863 );
nor  g18516 ( new_n20865 , new_n20855 , new_n20864 );
nor  g18517 ( new_n20866 , new_n20854 , new_n20865 );
nor  g18518 ( new_n20867 , new_n20853 , new_n20866 );
nor  g18519 ( new_n20868 , new_n20852 , new_n20867 );
nor  g18520 ( new_n20869_1 , new_n20850 , new_n20868 );
xnor g18521 ( n7999 , new_n20848 , new_n20869_1 );
xnor g18522 ( n8027 , new_n17712 , new_n17725 );
nor  g18523 ( new_n20872 , new_n14355 , new_n20792 );
not  g18524 ( new_n20873 , new_n20872 );
nor  g18525 ( new_n20874 , new_n6198 , new_n6244 );
xnor g18526 ( new_n20875 , n8614 , new_n6244 );
nor  g18527 ( new_n20876 , new_n6215 , new_n6250 );
nor  g18528 ( new_n20877 , n27037 , new_n6257 );
xnor g18529 ( new_n20878 , n27037 , new_n6256_1 );
nor  g18530 ( new_n20879_1 , n8964 , new_n6304 );
xnor g18531 ( new_n20880 , new_n6222 , new_n6304 );
nor  g18532 ( new_n20881 , new_n6227 , new_n6268 );
nor  g18533 ( new_n20882 , new_n4015 , new_n6273 );
and  g18534 ( new_n20883 , new_n20472 , new_n20475 );
or   g18535 ( new_n20884 , new_n20882 , new_n20883 );
xnor g18536 ( new_n20885 , new_n6227 , new_n6269 );
and  g18537 ( new_n20886 , new_n20884 , new_n20885 );
nor  g18538 ( new_n20887 , new_n20881 , new_n20886 );
and  g18539 ( new_n20888 , new_n20880 , new_n20887 );
or   g18540 ( new_n20889 , new_n20879_1 , new_n20888 );
and  g18541 ( new_n20890 , new_n20878 , new_n20889 );
nor  g18542 ( new_n20891 , new_n20877 , new_n20890 );
xnor g18543 ( new_n20892 , new_n6215 , new_n6251 );
and  g18544 ( new_n20893 , new_n20891 , new_n20892 );
or   g18545 ( new_n20894 , new_n20876 , new_n20893 );
and  g18546 ( new_n20895 , new_n20875 , new_n20894 );
nor  g18547 ( new_n20896 , new_n20874 , new_n20895 );
nor  g18548 ( new_n20897 , new_n6242 , new_n20896 );
nor  g18549 ( new_n20898 , new_n20873 , new_n20897 );
and  g18550 ( new_n20899 , new_n20873 , new_n20897 );
xnor g18551 ( new_n20900 , new_n6197 , new_n20896 );
nor  g18552 ( new_n20901 , new_n20793 , new_n20900 );
xnor g18553 ( new_n20902 , new_n20793 , new_n20900 );
not  g18554 ( new_n20903 , new_n20807 );
xor  g18555 ( new_n20904 , new_n20875 , new_n20894 );
nor  g18556 ( new_n20905 , new_n20903 , new_n20904 );
xnor g18557 ( new_n20906 , new_n20903 , new_n20904 );
xor  g18558 ( new_n20907 , new_n20891 , new_n20892 );
nor  g18559 ( new_n20908 , new_n9600 , new_n20907 );
xnor g18560 ( new_n20909 , new_n9600 , new_n20907 );
xor  g18561 ( new_n20910 , new_n20878 , new_n20889 );
and  g18562 ( new_n20911 , new_n9651 , new_n20910 );
xnor g18563 ( new_n20912 , new_n9651 , new_n20910 );
xnor g18564 ( new_n20913 , new_n20880 , new_n20887 );
nor  g18565 ( new_n20914 , new_n9660 , new_n20913 );
xnor g18566 ( new_n20915_1 , new_n9660 , new_n20913 );
xor  g18567 ( new_n20916 , new_n20884 , new_n20885 );
nor  g18568 ( new_n20917 , new_n9663 , new_n20916 );
xnor g18569 ( new_n20918 , new_n9663 , new_n20916 );
nor  g18570 ( new_n20919 , new_n9668 , new_n20476 );
nor  g18571 ( new_n20920 , new_n20477 , new_n20480 );
nor  g18572 ( new_n20921 , new_n20919 , new_n20920 );
nor  g18573 ( new_n20922 , new_n20918 , new_n20921 );
nor  g18574 ( new_n20923_1 , new_n20917 , new_n20922 );
nor  g18575 ( new_n20924 , new_n20915_1 , new_n20923_1 );
nor  g18576 ( new_n20925 , new_n20914 , new_n20924 );
nor  g18577 ( new_n20926 , new_n20912 , new_n20925 );
nor  g18578 ( new_n20927 , new_n20911 , new_n20926 );
nor  g18579 ( new_n20928 , new_n20909 , new_n20927 );
nor  g18580 ( new_n20929_1 , new_n20908 , new_n20928 );
nor  g18581 ( new_n20930 , new_n20906 , new_n20929_1 );
nor  g18582 ( new_n20931 , new_n20905 , new_n20930 );
nor  g18583 ( new_n20932 , new_n20902 , new_n20931 );
nor  g18584 ( new_n20933 , new_n20901 , new_n20932 );
nor  g18585 ( new_n20934 , new_n20899 , new_n20933 );
or   g18586 ( n8031 , new_n20898 , new_n20934 );
and  g18587 ( new_n20936_1 , n22626 , new_n16939 );
nor  g18588 ( new_n20937 , n22626 , new_n16939 );
nor  g18589 ( new_n20938 , new_n20937 , new_n16949 );
or   g18590 ( new_n20939 , new_n20803_1 , new_n20938 );
nor  g18591 ( new_n20940 , new_n20936_1 , new_n20939 );
not  g18592 ( new_n20941 , new_n20940 );
nor  g18593 ( new_n20942 , new_n19325 , new_n20941 );
xnor g18594 ( new_n20943 , new_n19325 , new_n20941 );
nor  g18595 ( new_n20944 , new_n16936 , new_n16950 );
not  g18596 ( new_n20945 , new_n16977 );
nor  g18597 ( new_n20946_1 , new_n16951_1 , new_n20945 );
nor  g18598 ( new_n20947 , new_n20944 , new_n20946_1 );
nor  g18599 ( new_n20948 , new_n20943 , new_n20947 );
nor  g18600 ( new_n20949 , new_n20942 , new_n20948 );
not  g18601 ( new_n20950 , new_n20949 );
or   g18602 ( new_n20951 , n9554 , new_n16992 );
and  g18603 ( new_n20952 , new_n20951 , new_n17022 );
and  g18604 ( new_n20953 , n9554 , new_n16992 );
or   g18605 ( new_n20954 , new_n19605 , new_n20953 );
nor  g18606 ( new_n20955 , new_n20952 , new_n20954 );
nor  g18607 ( new_n20956 , new_n20950 , new_n20955 );
not  g18608 ( new_n20957 , new_n20955 );
xnor g18609 ( new_n20958 , new_n20950 , new_n20957 );
xnor g18610 ( new_n20959 , new_n20943 , new_n20947 );
not  g18611 ( new_n20960 , new_n20959 );
nor  g18612 ( new_n20961 , new_n20957 , new_n20960 );
xnor g18613 ( new_n20962 , new_n20957 , new_n20960 );
nor  g18614 ( new_n20963 , new_n16978 , new_n17023 );
nor  g18615 ( new_n20964 , new_n17025 , new_n17080 );
nor  g18616 ( new_n20965 , new_n20963 , new_n20964 );
nor  g18617 ( new_n20966 , new_n20962 , new_n20965 );
or   g18618 ( new_n20967 , new_n20961 , new_n20966 );
and  g18619 ( new_n20968 , new_n20958 , new_n20967 );
nor  g18620 ( n8042 , new_n20956 , new_n20968 );
nor  g18621 ( new_n20970 , new_n9817 , new_n9910 );
nor  g18622 ( new_n20971 , new_n9911 , new_n9986 );
or   g18623 ( n8095 , new_n20970 , new_n20971 );
nor  g18624 ( new_n20973 , n4306 , new_n17625 );
xnor g18625 ( new_n20974 , n4306 , n23166 );
nor  g18626 ( new_n20975 , n3279 , new_n9079 );
xnor g18627 ( new_n20976 , n3279 , n10577 );
nor  g18628 ( new_n20977 , new_n9082 , n13914 );
xnor g18629 ( new_n20978 , n6381 , n13914 );
nor  g18630 ( new_n20979 , new_n9085 , n14702 );
and  g18631 ( new_n20980 , new_n19061 , new_n19072 );
or   g18632 ( new_n20981 , new_n20979 , new_n20980 );
and  g18633 ( new_n20982 , new_n20978 , new_n20981 );
or   g18634 ( new_n20983 , new_n20977 , new_n20982 );
and  g18635 ( new_n20984 , new_n20976 , new_n20983 );
or   g18636 ( new_n20985 , new_n20975 , new_n20984 );
and  g18637 ( new_n20986_1 , new_n20974 , new_n20985 );
nor  g18638 ( new_n20987 , new_n20973 , new_n20986_1 );
xnor g18639 ( new_n20988 , new_n8953 , new_n20987 );
xor  g18640 ( new_n20989 , new_n20974 , new_n20985 );
nor  g18641 ( new_n20990 , new_n8999 , new_n20989 );
xnor g18642 ( new_n20991 , new_n8999 , new_n20989 );
xor  g18643 ( new_n20992 , new_n20976 , new_n20983 );
nor  g18644 ( new_n20993 , new_n9003_1 , new_n20992 );
xnor g18645 ( new_n20994 , new_n9003_1 , new_n20992 );
xor  g18646 ( new_n20995 , new_n20978 , new_n20981 );
nor  g18647 ( new_n20996 , new_n9007 , new_n20995 );
xnor g18648 ( new_n20997 , new_n9007 , new_n20995 );
not  g18649 ( new_n20998 , new_n20997 );
and  g18650 ( new_n20999 , new_n9011 , new_n19073 );
and  g18651 ( new_n21000 , new_n19074 , new_n19088 );
nor  g18652 ( new_n21001 , new_n20999 , new_n21000 );
and  g18653 ( new_n21002 , new_n20998 , new_n21001 );
nor  g18654 ( new_n21003 , new_n20996 , new_n21002 );
nor  g18655 ( new_n21004 , new_n20994 , new_n21003 );
nor  g18656 ( new_n21005 , new_n20993 , new_n21004 );
nor  g18657 ( new_n21006 , new_n20991 , new_n21005 );
nor  g18658 ( new_n21007 , new_n20990 , new_n21006 );
xnor g18659 ( n8103 , new_n20988 , new_n21007 );
xnor g18660 ( n8109 , new_n18456 , new_n18467_1 );
nor  g18661 ( new_n21010 , new_n18878 , new_n18896 );
nor  g18662 ( new_n21011 , new_n18897 , new_n18925 );
or   g18663 ( n8127 , new_n21010 , new_n21011 );
xnor g18664 ( n8130 , new_n16480 , new_n16483 );
nor  g18665 ( new_n21014 , new_n3087 , n8856 );
xnor g18666 ( new_n21015 , n4319 , n8856 );
nor  g18667 ( new_n21016 , n14130 , new_n11610 );
xnor g18668 ( new_n21017_1 , n14130 , n23463 );
nor  g18669 ( new_n21018 , new_n3095 , n16482 );
xnor g18670 ( new_n21019 , n13074 , n16482 );
nor  g18671 ( new_n21020 , n9942 , new_n3099 );
and  g18672 ( new_n21021 , new_n2349 , new_n2379 );
or   g18673 ( new_n21022 , new_n21020 , new_n21021 );
and  g18674 ( new_n21023 , new_n21019 , new_n21022 );
or   g18675 ( new_n21024 , new_n21018 , new_n21023 );
and  g18676 ( new_n21025 , new_n21017_1 , new_n21024 );
or   g18677 ( new_n21026 , new_n21016 , new_n21025 );
and  g18678 ( new_n21027 , new_n21015 , new_n21026 );
nor  g18679 ( new_n21028 , new_n21014 , new_n21027 );
xnor g18680 ( new_n21029 , new_n7547 , new_n21028 );
nor  g18681 ( new_n21030 , new_n7550 , new_n21028 );
xnor g18682 ( new_n21031 , new_n7550 , new_n21028 );
xor  g18683 ( new_n21032 , new_n21015 , new_n21026 );
nor  g18684 ( new_n21033 , new_n7554 , new_n21032 );
xnor g18685 ( new_n21034_1 , new_n7554 , new_n21032 );
xor  g18686 ( new_n21035 , new_n21017_1 , new_n21024 );
nor  g18687 ( new_n21036 , new_n7558_1 , new_n21035 );
xnor g18688 ( new_n21037 , new_n7558_1 , new_n21035 );
not  g18689 ( new_n21038 , new_n21037 );
xor  g18690 ( new_n21039 , new_n21019 , new_n21022 );
and  g18691 ( new_n21040 , new_n7562 , new_n21039 );
xnor g18692 ( new_n21041 , new_n7562 , new_n21039 );
and  g18693 ( new_n21042 , new_n2380 , new_n2501 );
and  g18694 ( new_n21043 , new_n2502 , new_n2540 );
nor  g18695 ( new_n21044 , new_n21042 , new_n21043 );
nor  g18696 ( new_n21045 , new_n21041 , new_n21044 );
nor  g18697 ( new_n21046_1 , new_n21040 , new_n21045 );
and  g18698 ( new_n21047 , new_n21038 , new_n21046_1 );
nor  g18699 ( new_n21048 , new_n21036 , new_n21047 );
nor  g18700 ( new_n21049 , new_n21034_1 , new_n21048 );
nor  g18701 ( new_n21050 , new_n21033 , new_n21049 );
nor  g18702 ( new_n21051 , new_n21031 , new_n21050 );
nor  g18703 ( new_n21052 , new_n21030 , new_n21051 );
xnor g18704 ( n8135 , new_n21029 , new_n21052 );
xnor g18705 ( n8139 , new_n2529 , new_n7586 );
not  g18706 ( new_n21055 , new_n17865 );
nor  g18707 ( new_n21056 , n3018 , new_n21055 );
not  g18708 ( new_n21057 , new_n21056 );
nor  g18709 ( new_n21058 , n26660 , new_n21057 );
xnor g18710 ( new_n21059 , n13783 , new_n21058 );
xnor g18711 ( new_n21060 , new_n2981 , new_n21059 );
xnor g18712 ( new_n21061 , n26660 , new_n21056 );
and  g18713 ( new_n21062_1 , new_n2987 , new_n21061 );
xnor g18714 ( new_n21063 , new_n2987 , new_n21061 );
and  g18715 ( new_n21064 , new_n2992 , new_n17866 );
and  g18716 ( new_n21065 , new_n17867 , new_n17884 );
nor  g18717 ( new_n21066 , new_n21064 , new_n21065 );
nor  g18718 ( new_n21067 , new_n21063 , new_n21066 );
nor  g18719 ( new_n21068 , new_n21062_1 , new_n21067 );
xor  g18720 ( new_n21069 , new_n21060 , new_n21068 );
xnor g18721 ( new_n21070 , new_n6918 , new_n21069 );
xor  g18722 ( new_n21071 , new_n21063 , new_n21066 );
nor  g18723 ( new_n21072 , new_n6923 , new_n21071 );
xnor g18724 ( new_n21073 , new_n6923 , new_n21071 );
nor  g18725 ( new_n21074 , new_n6926 , new_n17885 );
nor  g18726 ( new_n21075 , new_n17886 , new_n17903 );
nor  g18727 ( new_n21076 , new_n21074 , new_n21075 );
nor  g18728 ( new_n21077 , new_n21073 , new_n21076 );
nor  g18729 ( new_n21078_1 , new_n21072 , new_n21077 );
xnor g18730 ( n8148 , new_n21070 , new_n21078_1 );
xor  g18731 ( n8149 , new_n17283 , new_n17284 );
xnor g18732 ( n8159 , new_n3903 , new_n3920 );
xnor g18733 ( n8179 , new_n2552 , new_n11560 );
xnor g18734 ( n8215 , new_n14613 , new_n14616 );
xnor g18735 ( n8267 , new_n18458 , new_n18465 );
xnor g18736 ( n8276 , new_n19487 , new_n19488 );
not  g18737 ( new_n21086 , new_n21058 );
nor  g18738 ( new_n21087 , n13783 , new_n21086 );
not  g18739 ( new_n21088 , new_n21087 );
nor  g18740 ( new_n21089 , n1654 , new_n21088 );
not  g18741 ( new_n21090 , new_n21089 );
nor  g18742 ( new_n21091 , n14440 , new_n21090 );
xnor g18743 ( new_n21092 , n22626 , new_n21091 );
nor  g18744 ( new_n21093_1 , new_n14785 , new_n21092 );
xnor g18745 ( new_n21094_1 , new_n14785 , new_n21092 );
xnor g18746 ( new_n21095_1 , n14440 , new_n21089 );
nor  g18747 ( new_n21096 , new_n2969 , new_n21095_1 );
xnor g18748 ( new_n21097 , new_n2969 , new_n21095_1 );
xnor g18749 ( new_n21098 , n1654 , new_n21087 );
and  g18750 ( new_n21099 , new_n2973 , new_n21098 );
and  g18751 ( new_n21100 , new_n2981 , new_n21059 );
nor  g18752 ( new_n21101 , new_n21060 , new_n21068 );
nor  g18753 ( new_n21102 , new_n21100 , new_n21101 );
xnor g18754 ( new_n21103 , new_n2973 , new_n21098 );
nor  g18755 ( new_n21104 , new_n21102 , new_n21103 );
or   g18756 ( new_n21105 , new_n21099 , new_n21104 );
nor  g18757 ( new_n21106 , new_n21097 , new_n21105 );
nor  g18758 ( new_n21107 , new_n21096 , new_n21106 );
nor  g18759 ( new_n21108 , new_n21094_1 , new_n21107 );
nor  g18760 ( new_n21109 , new_n21093_1 , new_n21108 );
not  g18761 ( new_n21110 , new_n21091 );
nor  g18762 ( new_n21111 , n22626 , new_n21110 );
xnor g18763 ( new_n21112 , new_n14810 , new_n21111 );
xnor g18764 ( new_n21113 , new_n21109 , new_n21112 );
nor  g18765 ( new_n21114 , new_n16852 , new_n21113 );
xnor g18766 ( new_n21115 , new_n16852 , new_n21113 );
xor  g18767 ( new_n21116 , new_n21094_1 , new_n21107 );
and  g18768 ( new_n21117 , new_n16857 , new_n21116 );
xnor g18769 ( new_n21118 , new_n16857 , new_n21116 );
xor  g18770 ( new_n21119 , new_n21097 , new_n21105 );
and  g18771 ( new_n21120 , new_n6833 , new_n21119 );
xor  g18772 ( new_n21121 , new_n21102 , new_n21103 );
nor  g18773 ( new_n21122 , new_n6913 , new_n21121 );
xnor g18774 ( new_n21123_1 , new_n6913 , new_n21121 );
nor  g18775 ( new_n21124 , new_n6918 , new_n21069 );
nor  g18776 ( new_n21125 , new_n21070 , new_n21078_1 );
nor  g18777 ( new_n21126 , new_n21124 , new_n21125 );
nor  g18778 ( new_n21127 , new_n21123_1 , new_n21126 );
nor  g18779 ( new_n21128 , new_n21122 , new_n21127 );
xnor g18780 ( new_n21129 , new_n6833 , new_n21119 );
nor  g18781 ( new_n21130 , new_n21128 , new_n21129 );
nor  g18782 ( new_n21131 , new_n21120 , new_n21130 );
nor  g18783 ( new_n21132 , new_n21118 , new_n21131 );
nor  g18784 ( new_n21133 , new_n21117 , new_n21132 );
nor  g18785 ( new_n21134_1 , new_n21115 , new_n21133 );
nor  g18786 ( new_n21135 , new_n21114 , new_n21134_1 );
and  g18787 ( new_n21136 , new_n16797 , new_n21135 );
or   g18788 ( new_n21137 , new_n14811 , new_n21111 );
nor  g18789 ( new_n21138_1 , new_n21109 , new_n21137 );
or   g18790 ( new_n21139 , new_n16797 , new_n21135 );
and  g18791 ( new_n21140 , new_n14811 , new_n21111 );
and  g18792 ( new_n21141 , new_n21109 , new_n21140 );
nor  g18793 ( new_n21142 , new_n21139 , new_n21141 );
nor  g18794 ( new_n21143 , new_n21138_1 , new_n21142 );
nor  g18795 ( n8288 , new_n21136 , new_n21143 );
xnor g18796 ( n8306 , new_n7400 , new_n11147 );
xor  g18797 ( n8320 , new_n7857 , new_n7910 );
xnor g18798 ( n8321 , new_n12279 , new_n12298 );
xnor g18799 ( n8339 , new_n16053 , new_n16066 );
xnor g18800 ( n8376 , new_n9009 , new_n9053 );
not  g18801 ( new_n21150 , new_n10134 );
xnor g18802 ( n8408 , new_n21150 , new_n18769 );
xnor g18803 ( n8417 , new_n14144 , new_n14145 );
xnor g18804 ( n8432 , new_n12709 , new_n12722 );
nor  g18805 ( new_n21154_1 , new_n10045 , new_n10049 );
and  g18806 ( new_n21155 , new_n10051 , new_n10098 );
nor  g18807 ( new_n21156 , new_n21154_1 , new_n21155 );
not  g18808 ( new_n21157_1 , new_n21156 );
and  g18809 ( new_n21158 , new_n10028 , new_n21157_1 );
nor  g18810 ( new_n21159 , new_n10028 , new_n10099 );
nor  g18811 ( new_n21160 , new_n10100 , new_n10163 );
nor  g18812 ( new_n21161 , new_n21159 , new_n21160 );
nor  g18813 ( new_n21162 , new_n21158 , new_n21161 );
nor  g18814 ( new_n21163 , new_n10028 , new_n21157_1 );
nor  g18815 ( new_n21164 , new_n21160 , new_n21163 );
nor  g18816 ( n8453 , new_n21162 , new_n21164 );
xnor g18817 ( n8480 , new_n13470 , new_n15345_1 );
xnor g18818 ( n8489 , new_n16200 , new_n16219_1 );
xnor g18819 ( n8505 , new_n21034_1 , new_n21048 );
xnor g18820 ( n8510 , new_n19168 , new_n19184 );
xnor g18821 ( n8519 , new_n8631 , new_n12002 );
xnor g18822 ( n8535 , new_n9688 , new_n9689_1 );
xnor g18823 ( n8550 , new_n18914 , new_n18917 );
xnor g18824 ( n8563 , new_n20045 , new_n20051 );
xnor g18825 ( n8594 , new_n13130 , new_n13131 );
xnor g18826 ( n8608 , new_n6934 , new_n6954 );
xnor g18827 ( n8620 , new_n4584 , new_n4585 );
xnor g18828 ( n8637 , new_n7371 , new_n7423 );
xnor g18829 ( n8662 , new_n16869 , new_n16870 );
xnor g18830 ( n8716 , new_n18503 , new_n18512 );
xnor g18831 ( new_n21180 , new_n7858 , new_n7861 );
xnor g18832 ( n8744 , new_n7908 , new_n21180 );
nor  g18833 ( new_n21182_1 , new_n7772 , new_n12681 );
or   g18834 ( new_n21183 , new_n20840 , new_n20845 );
and  g18835 ( new_n21184 , new_n20839 , new_n21183 );
nor  g18836 ( new_n21185 , new_n21182_1 , new_n21184 );
xnor g18837 ( new_n21186 , new_n15096 , new_n21185 );
nor  g18838 ( new_n21187 , new_n4907 , new_n6022_1 );
and  g18839 ( new_n21188 , new_n20765 , new_n20768 );
nor  g18840 ( new_n21189 , new_n21187 , new_n21188 );
xnor g18841 ( new_n21190 , new_n17495 , new_n21189 );
xnor g18842 ( new_n21191 , new_n21186 , new_n21190 );
not  g18843 ( new_n21192 , new_n20769 );
not  g18844 ( new_n21193_1 , new_n20847 );
nor  g18845 ( new_n21194 , new_n21192 , new_n21193_1 );
xnor g18846 ( new_n21195 , new_n21192 , new_n20847 );
nor  g18847 ( new_n21196 , new_n20771 , new_n20851 );
xnor g18848 ( new_n21197 , new_n15883 , new_n20851 );
nor  g18849 ( new_n21198 , new_n15885_1 , new_n17096 );
nor  g18850 ( new_n21199 , new_n17097 , new_n17128 );
nor  g18851 ( new_n21200 , new_n21198 , new_n21199 );
and  g18852 ( new_n21201 , new_n21197 , new_n21200 );
nor  g18853 ( new_n21202 , new_n21196 , new_n21201 );
and  g18854 ( new_n21203_1 , new_n21195 , new_n21202 );
nor  g18855 ( new_n21204 , new_n21194 , new_n21203_1 );
xnor g18856 ( n8803 , new_n21191 , new_n21204 );
and  g18857 ( new_n21206 , new_n5500 , new_n19906 );
nor  g18858 ( new_n21207 , new_n5610 , new_n19907 );
and  g18859 ( new_n21208 , new_n19908 , new_n19926 );
nor  g18860 ( new_n21209 , new_n21207 , new_n21208 );
xnor g18861 ( new_n21210 , new_n21206 , new_n21209 );
nor  g18862 ( new_n21211 , n4319 , n16544 );
or   g18863 ( new_n21212 , new_n15544 , new_n15561 );
and  g18864 ( new_n21213 , new_n15543 , new_n21212 );
nor  g18865 ( new_n21214 , new_n21211 , new_n21213 );
xnor g18866 ( new_n21215 , new_n21210 , new_n21214 );
nor  g18867 ( new_n21216 , new_n15563 , new_n19927 );
nor  g18868 ( new_n21217 , new_n19928 , new_n19946 );
nor  g18869 ( new_n21218 , new_n21216 , new_n21217 );
xnor g18870 ( new_n21219 , new_n21215 , new_n21218 );
not  g18871 ( new_n21220 , new_n21219 );
xnor g18872 ( new_n21221 , new_n7695 , new_n21220 );
nor  g18873 ( new_n21222_1 , new_n7698_1 , new_n20501 );
nor  g18874 ( new_n21223 , new_n20502 , new_n20536 );
nor  g18875 ( new_n21224 , new_n21222_1 , new_n21223 );
xnor g18876 ( n8809 , new_n21221 , new_n21224 );
nor  g18877 ( new_n21226_1 , new_n17496 , new_n21189 );
not  g18878 ( new_n21227 , new_n21226_1 );
nor  g18879 ( new_n21228 , n3324 , new_n17831 );
and  g18880 ( new_n21229 , new_n20752 , new_n20763 );
nor  g18881 ( new_n21230 , new_n21228 , new_n21229 );
and  g18882 ( new_n21231 , new_n17825 , new_n21230 );
xnor g18883 ( new_n21232 , new_n21227 , new_n21231 );
not  g18884 ( new_n21233 , new_n21190 );
xnor g18885 ( new_n21234 , new_n17823 , new_n21230 );
nor  g18886 ( new_n21235 , new_n21233 , new_n21234 );
xnor g18887 ( new_n21236 , new_n21233 , new_n21234 );
nor  g18888 ( new_n21237 , new_n20764 , new_n20769 );
nor  g18889 ( new_n21238_1 , new_n20770 , new_n20784 );
nor  g18890 ( new_n21239 , new_n21237 , new_n21238_1 );
nor  g18891 ( new_n21240 , new_n21236 , new_n21239 );
nor  g18892 ( new_n21241 , new_n21235 , new_n21240 );
xnor g18893 ( n8821 , new_n21232 , new_n21241 );
xnor g18894 ( n8824 , new_n15314 , new_n15315 );
xor  g18895 ( n8849 , new_n17445 , new_n17446 );
xnor g18896 ( n8861 , new_n13574 , new_n13582 );
xnor g18897 ( new_n21246 , n8856 , n22442 );
nor  g18898 ( new_n21247 , new_n8273 , n14130 );
and  g18899 ( new_n21248 , new_n19679 , new_n19702 );
or   g18900 ( new_n21249 , new_n21247 , new_n21248 );
xor  g18901 ( new_n21250 , new_n21246 , new_n21249 );
xnor g18902 ( new_n21251 , new_n7179 , n3324 );
nor  g18903 ( new_n21252 , n17911 , n25331 );
and  g18904 ( new_n21253 , new_n19669 , new_n19672 );
or   g18905 ( new_n21254_1 , new_n21252 , new_n21253 );
xor  g18906 ( new_n21255 , new_n21251 , new_n21254_1 );
xnor g18907 ( new_n21256 , new_n7522 , new_n21255 );
nor  g18908 ( new_n21257 , new_n7488 , new_n19673 );
and  g18909 ( new_n21258 , new_n19674 , new_n19677 );
nor  g18910 ( new_n21259 , new_n21257 , new_n21258 );
xnor g18911 ( new_n21260 , new_n21256 , new_n21259 );
xnor g18912 ( new_n21261 , new_n21250 , new_n21260 );
and  g18913 ( new_n21262 , new_n19678 , new_n19703 );
and  g18914 ( new_n21263 , new_n19704 , new_n19733 );
or   g18915 ( new_n21264 , new_n21262 , new_n21263 );
xor  g18916 ( n8862 , new_n21261 , new_n21264 );
xor  g18917 ( n8884 , new_n13475 , new_n13476 );
not  g18918 ( new_n21267 , new_n17910 );
xnor g18919 ( n8909 , new_n21267 , new_n18681 );
xnor g18920 ( n8911 , new_n11537 , new_n11578 );
xnor g18921 ( n8971 , new_n11087 , new_n11088 );
xnor g18922 ( n8982 , new_n20906 , new_n20929_1 );
xnor g18923 ( n8993 , new_n5425 , new_n5441 );
xor  g18924 ( n9012 , new_n14153 , new_n14154 );
nor  g18925 ( new_n21274 , new_n19821 , new_n19824 );
or   g18926 ( new_n21275 , new_n4453 , new_n19831 );
nor  g18927 ( new_n21276_1 , new_n19829 , new_n21275 );
xnor g18928 ( new_n21277 , new_n21274 , new_n21276_1 );
nor  g18929 ( new_n21278 , new_n19825 , new_n19833 );
nor  g18930 ( new_n21279 , new_n19834 , new_n19879 );
nor  g18931 ( new_n21280 , new_n21278 , new_n21279 );
xnor g18932 ( n9032 , new_n21277 , new_n21280 );
xor  g18933 ( n9042 , new_n15807 , new_n15808 );
xnor g18934 ( n9046 , new_n17043 , new_n17074 );
xnor g18935 ( n9047 , new_n8142 , new_n8200 );
xnor g18936 ( n9104 , new_n15034 , new_n15035 );
nor  g18937 ( new_n21286 , new_n20193 , new_n20201 );
nor  g18938 ( new_n21287_1 , new_n20185 , new_n21286 );
and  g18939 ( new_n21288 , new_n20193 , new_n20201 );
nor  g18940 ( new_n21289 , new_n15180_1 , new_n21288 );
nor  g18941 ( new_n21290 , new_n21287_1 , new_n21289 );
not  g18942 ( new_n21291 , new_n21290 );
xnor g18943 ( new_n21292 , new_n19127 , new_n21291 );
nor  g18944 ( new_n21293 , new_n19127 , new_n20203 );
nor  g18945 ( new_n21294 , new_n20204 , new_n20212 );
nor  g18946 ( new_n21295 , new_n21293 , new_n21294 );
xor  g18947 ( n9129 , new_n21292 , new_n21295 );
xnor g18948 ( n9146 , new_n18827 , new_n18858_1 );
xnor g18949 ( n9164 , new_n6702 , new_n8631 );
xor  g18950 ( n9166 , new_n12646 , new_n12647 );
xnor g18951 ( new_n21300 , new_n17815 , new_n17842 );
xnor g18952 ( n9182 , new_n17853 , new_n21300 );
xnor g18953 ( n9191 , new_n7136 , new_n7168 );
xnor g18954 ( n9217 , new_n11528 , new_n11583 );
xor  g18955 ( n9220 , new_n15968 , new_n15969 );
xnor g18956 ( n9261 , new_n18842 , new_n18848 );
xnor g18957 ( new_n21306 , n3324 , n22626 );
nor  g18958 ( new_n21307 , n14440 , new_n19668 );
and  g18959 ( new_n21308 , new_n18471 , new_n18491 );
or   g18960 ( new_n21309 , new_n21307 , new_n21308 );
xor  g18961 ( new_n21310 , new_n21306 , new_n21309 );
and  g18962 ( new_n21311 , new_n17846 , new_n21310 );
xnor g18963 ( new_n21312 , new_n17846 , new_n21310 );
and  g18964 ( new_n21313 , new_n3032 , new_n18492 );
and  g18965 ( new_n21314 , new_n18493 , new_n18518 );
nor  g18966 ( new_n21315 , new_n21313 , new_n21314 );
nor  g18967 ( new_n21316 , new_n21312 , new_n21315 );
nor  g18968 ( new_n21317_1 , new_n21311 , new_n21316 );
not  g18969 ( new_n21318 , new_n21317_1 );
nor  g18970 ( new_n21319 , new_n20751 , n22626 );
and  g18971 ( new_n21320 , new_n21306 , new_n21309 );
nor  g18972 ( new_n21321 , new_n21319 , new_n21320 );
xnor g18973 ( new_n21322 , new_n17842 , new_n21321 );
xnor g18974 ( n9287 , new_n21318 , new_n21322 );
xor  g18975 ( n9308 , new_n13965 , new_n13974 );
xnor g18976 ( n9344 , new_n4983 , new_n5020_1 );
xnor g18977 ( n9364 , new_n3694 , new_n3711 );
or   g18978 ( new_n21327 , new_n17841 , new_n21321 );
nor  g18979 ( new_n21328 , new_n21317_1 , new_n21327 );
and  g18980 ( new_n21329 , new_n17839 , new_n21328 );
and  g18981 ( new_n21330 , new_n17841 , new_n21321 );
and  g18982 ( new_n21331 , new_n21317_1 , new_n21330 );
and  g18983 ( new_n21332 , new_n17857 , new_n21331 );
or   g18984 ( n9371 , new_n21329 , new_n21332 );
xnor g18985 ( n9382 , new_n21150 , new_n10135 );
xor  g18986 ( n9403 , new_n20958 , new_n20967 );
xnor g18987 ( n9419 , new_n12628 , new_n12653 );
xnor g18988 ( n9423 , new_n20709_1 , new_n20732 );
xnor g18989 ( n9430 , new_n18499 , new_n18514 );
xnor g18990 ( new_n21339 , n23272 , n25120 );
and  g18991 ( new_n21340 , n8363 , new_n4361 );
xnor g18992 ( new_n21341 , n8363 , n11481 );
and  g18993 ( new_n21342 , n14680 , new_n4365 );
and  g18994 ( new_n21343 , new_n15482 , new_n15485 );
or   g18995 ( new_n21344 , new_n21342 , new_n21343 );
and  g18996 ( new_n21345 , new_n21341 , new_n21344 );
or   g18997 ( new_n21346 , new_n21340 , new_n21345 );
xor  g18998 ( new_n21347 , new_n21339 , new_n21346 );
xnor g18999 ( new_n21348 , new_n16950 , new_n21347 );
xor  g19000 ( new_n21349_1 , new_n21341 , new_n21344 );
and  g19001 ( new_n21350 , new_n16974 , new_n21349_1 );
xnor g19002 ( new_n21351 , new_n16974 , new_n21349_1 );
and  g19003 ( new_n21352 , new_n15486 , new_n15492 );
nor  g19004 ( new_n21353 , new_n15493 , new_n15496_1 );
nor  g19005 ( new_n21354 , new_n21352 , new_n21353 );
nor  g19006 ( new_n21355 , new_n21351 , new_n21354 );
nor  g19007 ( new_n21356 , new_n21350 , new_n21355 );
xor  g19008 ( new_n21357 , new_n21348 , new_n21356 );
xnor g19009 ( new_n21358 , new_n17024 , new_n21357 );
xor  g19010 ( new_n21359 , new_n21351 , new_n21354 );
nor  g19011 ( new_n21360 , new_n17026 , new_n21359 );
xnor g19012 ( new_n21361 , new_n17026 , new_n21359 );
nor  g19013 ( new_n21362 , new_n15498 , new_n17032 );
xnor g19014 ( new_n21363 , new_n15498 , new_n17032 );
nor  g19015 ( new_n21364 , new_n10576 , new_n17039 );
xnor g19016 ( new_n21365_1 , new_n10576 , new_n17039 );
nor  g19017 ( new_n21366 , new_n10578 , new_n17048 );
xnor g19018 ( new_n21367_1 , new_n10578 , new_n17048 );
nor  g19019 ( new_n21368 , new_n10582 , new_n17054 );
and  g19020 ( new_n21369 , new_n10584 , new_n14764 );
nor  g19021 ( new_n21370 , new_n14765 , new_n14777 );
nor  g19022 ( new_n21371 , new_n21369 , new_n21370 );
xnor g19023 ( new_n21372 , new_n10600 , new_n17051 );
nor  g19024 ( new_n21373 , new_n21371 , new_n21372 );
or   g19025 ( new_n21374 , new_n21368 , new_n21373 );
nor  g19026 ( new_n21375 , new_n21367_1 , new_n21374 );
nor  g19027 ( new_n21376 , new_n21366 , new_n21375 );
nor  g19028 ( new_n21377 , new_n21365_1 , new_n21376 );
nor  g19029 ( new_n21378 , new_n21364 , new_n21377 );
nor  g19030 ( new_n21379 , new_n21363 , new_n21378 );
nor  g19031 ( new_n21380 , new_n21362 , new_n21379 );
nor  g19032 ( new_n21381 , new_n21361 , new_n21380 );
or   g19033 ( new_n21382 , new_n21360 , new_n21381 );
xor  g19034 ( n9435 , new_n21358 , new_n21382 );
xnor g19035 ( n9451 , new_n15891 , new_n15919 );
xnor g19036 ( new_n21385 , n10763 , n12657 );
nor  g19037 ( new_n21386 , new_n2890 , n17077 );
and  g19038 ( new_n21387 , new_n18967 , new_n18974 );
or   g19039 ( new_n21388 , new_n21386 , new_n21387 );
xor  g19040 ( new_n21389 , new_n21385 , new_n21388 );
xnor g19041 ( new_n21390 , new_n19678 , new_n21389 );
nor  g19042 ( new_n21391 , new_n18975 , new_n18995 );
and  g19043 ( new_n21392 , new_n18997 , new_n19007 );
nor  g19044 ( new_n21393 , new_n21391 , new_n21392 );
xnor g19045 ( n9458 , new_n21390 , new_n21393 );
nor  g19046 ( new_n21395 , new_n10030 , n12507 );
xnor g19047 ( new_n21396_1 , n11220 , n12507 );
nor  g19048 ( new_n21397 , n15077 , new_n17810 );
and  g19049 ( new_n21398_1 , new_n14683 , new_n14702_1 );
or   g19050 ( new_n21399_1 , new_n21397 , new_n21398_1 );
and  g19051 ( new_n21400 , new_n21396_1 , new_n21399_1 );
nor  g19052 ( new_n21401 , new_n21395 , new_n21400 );
not  g19053 ( new_n21402 , new_n21401 );
xnor g19054 ( new_n21403 , new_n20401 , new_n21402 );
xor  g19055 ( new_n21404_1 , new_n21396_1 , new_n21399_1 );
nor  g19056 ( new_n21405 , new_n20403_1 , new_n21404_1 );
xnor g19057 ( new_n21406 , new_n20403_1 , new_n21404_1 );
nor  g19058 ( new_n21407 , new_n14682 , new_n14703 );
nor  g19059 ( new_n21408 , new_n14704_1 , new_n14734_1 );
nor  g19060 ( new_n21409 , new_n21407 , new_n21408 );
nor  g19061 ( new_n21410 , new_n21406 , new_n21409 );
nor  g19062 ( new_n21411 , new_n21405 , new_n21410 );
xnor g19063 ( n9459 , new_n21403 , new_n21411 );
xnor g19064 ( n9508 , new_n14976 , new_n14977_1 );
xnor g19065 ( n9552 , new_n12619 , new_n12657_1 );
xnor g19066 ( n9556 , new_n4587 , new_n4588_1 );
xnor g19067 ( n9558 , new_n8832 , new_n11060 );
xnor g19068 ( n9616 , new_n14145 , new_n20604_1 );
xnor g19069 ( n9622 , new_n8539 , new_n8566 );
xnor g19070 ( n9626 , new_n16397 , new_n16412 );
xnor g19071 ( n9633 , new_n4576 , new_n4594 );
not  g19072 ( new_n21421 , n23272 );
and  g19073 ( new_n21422 , new_n21421 , n25120 );
and  g19074 ( new_n21423 , new_n21339 , new_n21346 );
nor  g19075 ( new_n21424 , new_n21422 , new_n21423 );
not  g19076 ( new_n21425 , new_n21424 );
nor  g19077 ( new_n21426 , new_n20941 , new_n21425 );
xnor g19078 ( new_n21427 , new_n20941 , new_n21424 );
and  g19079 ( new_n21428 , new_n16950 , new_n21347 );
nor  g19080 ( new_n21429 , new_n21348 , new_n21356 );
nor  g19081 ( new_n21430 , new_n21428 , new_n21429 );
and  g19082 ( new_n21431 , new_n21427 , new_n21430 );
nor  g19083 ( new_n21432 , new_n21426 , new_n21431 );
not  g19084 ( new_n21433 , new_n21432 );
nor  g19085 ( new_n21434 , new_n5542 , new_n21433 );
xnor g19086 ( new_n21435 , new_n10165_1 , new_n21433 );
xnor g19087 ( new_n21436 , new_n21427 , new_n21430 );
not  g19088 ( new_n21437 , new_n21436 );
nor  g19089 ( new_n21438 , new_n10165_1 , new_n21437 );
xnor g19090 ( new_n21439 , new_n10165_1 , new_n21437 );
nor  g19091 ( new_n21440 , new_n5544 , new_n21357 );
and  g19092 ( new_n21441 , new_n5619 , new_n21359 );
xnor g19093 ( new_n21442 , new_n5619 , new_n21359 );
nor  g19094 ( new_n21443 , new_n5626 , new_n15497 );
nor  g19095 ( new_n21444 , new_n15499 , new_n15502 );
nor  g19096 ( new_n21445 , new_n21443 , new_n21444 );
nor  g19097 ( new_n21446_1 , new_n21442 , new_n21445 );
or   g19098 ( new_n21447 , new_n21441 , new_n21446_1 );
xnor g19099 ( new_n21448 , new_n5544 , new_n21357 );
nor  g19100 ( new_n21449 , new_n21447 , new_n21448 );
or   g19101 ( new_n21450 , new_n21440 , new_n21449 );
nor  g19102 ( new_n21451 , new_n21439 , new_n21450 );
or   g19103 ( new_n21452 , new_n21438 , new_n21451 );
and  g19104 ( new_n21453 , new_n21435 , new_n21452 );
nor  g19105 ( n9635 , new_n21434 , new_n21453 );
xnor g19106 ( n9648 , new_n19205 , new_n19208 );
xnor g19107 ( n9689 , new_n5003 , new_n16081 );
xnor g19108 ( n9695 , new_n10747 , new_n10765 );
xnor g19109 ( n9699 , new_n7560 , new_n7600 );
xnor g19110 ( new_n21459 , new_n14513 , new_n16500 );
nor  g19111 ( new_n21460 , new_n14513 , new_n16503 );
nor  g19112 ( new_n21461 , new_n15937 , new_n15975 );
nor  g19113 ( new_n21462 , new_n21460 , new_n21461 );
xor  g19114 ( n9726 , new_n21459 , new_n21462 );
xnor g19115 ( n9753 , new_n9963 , new_n13142 );
xnor g19116 ( n9761 , new_n3360 , new_n3379 );
xnor g19117 ( n9763 , new_n9931 , new_n9978 );
xnor g19118 ( n9767 , new_n13472 , new_n13473 );
xnor g19119 ( n9771 , new_n13376 , new_n13628 );
xor  g19120 ( n9778 , new_n21041 , new_n21044 );
xnor g19121 ( n9783 , new_n15696 , new_n15705 );
xnor g19122 ( n9803 , new_n6733 , new_n6735 );
and  g19123 ( new_n21472_1 , new_n11610 , new_n20545 );
and  g19124 ( new_n21473 , new_n3087 , new_n21472_1 );
xnor g19125 ( new_n21474 , n4319 , new_n21472_1 );
not  g19126 ( new_n21475 , new_n21474 );
nor  g19127 ( new_n21476 , new_n17789 , new_n21475 );
nor  g19128 ( new_n21477 , new_n17788 , new_n21474 );
nor  g19129 ( new_n21478 , new_n17793 , new_n20547 );
and  g19130 ( new_n21479 , new_n17793 , new_n20547 );
and  g19131 ( new_n21480 , new_n16564 , new_n20549 );
or   g19132 ( new_n21481 , new_n16564 , new_n20549 );
nor  g19133 ( new_n21482 , new_n16567 , new_n20553 );
nor  g19134 ( new_n21483 , new_n16570 , new_n20558 );
xnor g19135 ( new_n21484 , new_n16571 , new_n20556 );
and  g19136 ( new_n21485 , new_n6680 , new_n6696 );
nor  g19137 ( new_n21486 , new_n6697 , new_n6720 );
nor  g19138 ( new_n21487 , new_n21485 , new_n21486 );
nor  g19139 ( new_n21488 , new_n21484 , new_n21487 );
nor  g19140 ( new_n21489_1 , new_n21483 , new_n21488 );
xor  g19141 ( new_n21490 , new_n16567 , new_n20553 );
and  g19142 ( new_n21491 , new_n21489_1 , new_n21490 );
nor  g19143 ( new_n21492 , new_n21482 , new_n21491 );
and  g19144 ( new_n21493 , new_n21481 , new_n21492 );
nor  g19145 ( new_n21494 , new_n21480 , new_n21493 );
nor  g19146 ( new_n21495 , new_n21479 , new_n21494 );
nor  g19147 ( new_n21496 , new_n21478 , new_n21495 );
nor  g19148 ( new_n21497 , new_n21477 , new_n21496 );
nor  g19149 ( new_n21498 , new_n21476 , new_n21497 );
xnor g19150 ( new_n21499 , new_n17784_1 , new_n21498 );
xnor g19151 ( new_n21500 , new_n21473 , new_n21499 );
nor  g19152 ( new_n21501 , new_n3327 , new_n21500 );
xnor g19153 ( new_n21502 , new_n3327 , new_n21500 );
xnor g19154 ( new_n21503 , new_n17789 , new_n21474 );
xnor g19155 ( new_n21504 , new_n21496 , new_n21503 );
nor  g19156 ( new_n21505 , new_n3334 , new_n21504 );
xnor g19157 ( new_n21506 , new_n3334 , new_n21504 );
xnor g19158 ( new_n21507 , new_n17793 , new_n20546 );
xnor g19159 ( new_n21508 , new_n21494 , new_n21507 );
nor  g19160 ( new_n21509 , new_n3338 , new_n21508 );
xnor g19161 ( new_n21510 , new_n3338 , new_n21508 );
xnor g19162 ( new_n21511 , new_n16564 , new_n20549 );
xnor g19163 ( new_n21512 , new_n21492 , new_n21511 );
nor  g19164 ( new_n21513 , new_n3342 , new_n21512 );
xnor g19165 ( new_n21514 , new_n3342 , new_n21512 );
xnor g19166 ( new_n21515 , new_n21489_1 , new_n21490 );
nor  g19167 ( new_n21516 , new_n3346 , new_n21515 );
xnor g19168 ( new_n21517 , new_n3346 , new_n21515 );
xor  g19169 ( new_n21518 , new_n21484 , new_n21487 );
nor  g19170 ( new_n21519 , new_n3350 , new_n21518 );
xnor g19171 ( new_n21520 , new_n3350 , new_n21518 );
nor  g19172 ( new_n21521 , new_n3354 , new_n6721 );
nor  g19173 ( new_n21522 , new_n6722 , new_n6742 );
nor  g19174 ( new_n21523 , new_n21521 , new_n21522 );
nor  g19175 ( new_n21524 , new_n21520 , new_n21523 );
nor  g19176 ( new_n21525_1 , new_n21519 , new_n21524 );
nor  g19177 ( new_n21526 , new_n21517 , new_n21525_1 );
nor  g19178 ( new_n21527 , new_n21516 , new_n21526 );
nor  g19179 ( new_n21528 , new_n21514 , new_n21527 );
nor  g19180 ( new_n21529 , new_n21513 , new_n21528 );
nor  g19181 ( new_n21530 , new_n21510 , new_n21529 );
nor  g19182 ( new_n21531 , new_n21509 , new_n21530 );
nor  g19183 ( new_n21532 , new_n21506 , new_n21531 );
nor  g19184 ( new_n21533 , new_n21505 , new_n21532 );
nor  g19185 ( new_n21534 , new_n21502 , new_n21533 );
nor  g19186 ( new_n21535 , new_n21501 , new_n21534 );
not  g19187 ( new_n21536 , new_n21498 );
nor  g19188 ( new_n21537 , new_n17784_1 , new_n21536 );
xnor g19189 ( new_n21538_1 , new_n17744 , new_n21473 );
and  g19190 ( new_n21539 , new_n21537 , new_n21538_1 );
nor  g19191 ( new_n21540 , new_n21498 , new_n21538_1 );
nor  g19192 ( new_n21541 , new_n21539 , new_n21540 );
and  g19193 ( new_n21542 , new_n21535 , new_n21541 );
or   g19194 ( new_n21543 , new_n17745 , new_n21473 );
nor  g19195 ( new_n21544 , new_n21536 , new_n21543 );
xor  g19196 ( n9833 , new_n21542 , new_n21544 );
not  g19197 ( new_n21546 , new_n17217 );
nor  g19198 ( new_n21547 , n13775 , new_n21546 );
and  g19199 ( new_n21548 , new_n8646 , new_n21547 );
and  g19200 ( new_n21549_1 , new_n11842_1 , new_n21548 );
or   g19201 ( new_n21550 , new_n17781 , new_n21549_1 );
xnor g19202 ( new_n21551 , n25972 , new_n21548 );
and  g19203 ( new_n21552 , new_n17760 , new_n21551 );
xnor g19204 ( new_n21553 , new_n17760 , new_n21551 );
xnor g19205 ( new_n21554 , n21915 , new_n21547 );
and  g19206 ( new_n21555 , new_n17765 , new_n21554 );
xnor g19207 ( new_n21556 , new_n17764 , new_n21554 );
and  g19208 ( new_n21557 , new_n16534 , new_n17218 );
and  g19209 ( new_n21558 , new_n17219_1 , new_n17248 );
or   g19210 ( new_n21559 , new_n21557 , new_n21558 );
and  g19211 ( new_n21560 , new_n21556 , new_n21559 );
nor  g19212 ( new_n21561 , new_n21555 , new_n21560 );
nor  g19213 ( new_n21562 , new_n21553 , new_n21561 );
nor  g19214 ( new_n21563 , new_n21552 , new_n21562 );
not  g19215 ( new_n21564 , new_n21563 );
nor  g19216 ( new_n21565 , new_n21550 , new_n21564 );
not  g19217 ( new_n21566 , new_n17251_1 );
nor  g19218 ( new_n21567 , n3710 , new_n21566 );
and  g19219 ( new_n21568 , new_n8789 , new_n21567 );
and  g19220 ( new_n21569 , new_n8719 , new_n21568 );
xnor g19221 ( new_n21570 , new_n16496 , new_n21569 );
xnor g19222 ( new_n21571 , n12507 , new_n21568 );
nor  g19223 ( new_n21572 , new_n12818 , new_n21571 );
xnor g19224 ( new_n21573 , n15077 , new_n21567 );
nor  g19225 ( new_n21574 , new_n5304 , new_n21573 );
xnor g19226 ( new_n21575 , new_n5304 , new_n21573 );
and  g19227 ( new_n21576 , new_n5341 , new_n17252 );
and  g19228 ( new_n21577 , new_n17253 , new_n17256 );
nor  g19229 ( new_n21578 , new_n21576 , new_n21577 );
not  g19230 ( new_n21579 , new_n21578 );
nor  g19231 ( new_n21580 , new_n21575 , new_n21579 );
nor  g19232 ( new_n21581 , new_n21574 , new_n21580 );
xnor g19233 ( new_n21582 , new_n12818 , new_n21571 );
nor  g19234 ( new_n21583 , new_n21581 , new_n21582 );
nor  g19235 ( new_n21584 , new_n21572 , new_n21583 );
xnor g19236 ( new_n21585 , new_n21570 , new_n21584 );
xnor g19237 ( new_n21586 , new_n17782 , new_n21549_1 );
xnor g19238 ( new_n21587 , new_n21564 , new_n21586 );
nor  g19239 ( new_n21588 , new_n21585 , new_n21587 );
xnor g19240 ( new_n21589 , new_n21585 , new_n21587 );
xnor g19241 ( new_n21590 , new_n21553 , new_n21561 );
xnor g19242 ( new_n21591 , new_n21581 , new_n21582 );
not  g19243 ( new_n21592 , new_n21591 );
and  g19244 ( new_n21593 , new_n21590 , new_n21592 );
xnor g19245 ( new_n21594 , new_n21590 , new_n21592 );
xnor g19246 ( new_n21595 , new_n21575 , new_n21578 );
not  g19247 ( new_n21596 , new_n21595 );
xor  g19248 ( new_n21597 , new_n21556 , new_n21559 );
nor  g19249 ( new_n21598 , new_n21596 , new_n21597 );
xnor g19250 ( new_n21599_1 , new_n21596 , new_n21597 );
nor  g19251 ( new_n21600 , new_n17249 , new_n17257 );
nor  g19252 ( new_n21601 , new_n17258 , new_n17291 );
nor  g19253 ( new_n21602 , new_n21600 , new_n21601 );
nor  g19254 ( new_n21603 , new_n21599_1 , new_n21602 );
nor  g19255 ( new_n21604 , new_n21598 , new_n21603 );
nor  g19256 ( new_n21605 , new_n21594 , new_n21604 );
nor  g19257 ( new_n21606 , new_n21593 , new_n21605 );
nor  g19258 ( new_n21607 , new_n21589 , new_n21606 );
or   g19259 ( new_n21608 , new_n21588 , new_n21607 );
and  g19260 ( new_n21609 , new_n21565 , new_n21608 );
xor  g19261 ( new_n21610 , new_n21565 , new_n21608 );
or   g19262 ( new_n21611 , new_n15927 , new_n21569 );
nor  g19263 ( new_n21612 , new_n21611 , new_n21584 );
not  g19264 ( new_n21613 , new_n21612 );
nor  g19265 ( new_n21614 , new_n21610 , new_n21613 );
or   g19266 ( n9838 , new_n21609 , new_n21614 );
xnor g19267 ( n9867 , new_n19354_1 , new_n19357_1 );
nor  g19268 ( new_n21617 , new_n5686 , new_n18935 );
and  g19269 ( new_n21618 , new_n18936 , new_n18939 );
nor  g19270 ( new_n21619 , new_n21617 , new_n21618 );
nor  g19271 ( new_n21620 , new_n20166 , new_n21619 );
xnor g19272 ( new_n21621 , new_n20147 , new_n21619 );
nor  g19273 ( new_n21622 , new_n8134 , new_n21621 );
nor  g19274 ( new_n21623 , new_n18928 , new_n18940_1 );
nor  g19275 ( new_n21624 , new_n18941 , new_n18944 );
nor  g19276 ( new_n21625 , new_n21623 , new_n21624 );
xnor g19277 ( new_n21626 , new_n8134 , new_n21621 );
nor  g19278 ( new_n21627 , new_n21625 , new_n21626 );
nor  g19279 ( new_n21628_1 , new_n21622 , new_n21627 );
nor  g19280 ( new_n21629 , new_n21620 , new_n21628_1 );
nor  g19281 ( n9890 , new_n8028 , new_n21629 );
xor  g19282 ( n9917 , new_n17792 , new_n17801 );
xnor g19283 ( n9919 , new_n20420 , new_n20427 );
xnor g19284 ( n9938 , new_n17957 , new_n17970 );
xnor g19285 ( n9946 , new_n17612 , new_n17613 );
xnor g19286 ( new_n21635 , new_n4907 , n21784 );
nor  g19287 ( new_n21636 , n2858 , n5521 );
xnor g19288 ( new_n21637_1 , n2858 , n5521 );
nor  g19289 ( new_n21638 , n2659 , n11926 );
xnor g19290 ( new_n21639 , n2659 , n11926 );
nor  g19291 ( new_n21640 , n4325 , n24327 );
xnor g19292 ( new_n21641 , new_n5991 , n24327 );
nor  g19293 ( new_n21642 , new_n14435 , new_n4922 );
or   g19294 ( new_n21643 , n5337 , n22198 );
nor  g19295 ( new_n21644 , n626 , n20826 );
and  g19296 ( new_n21645_1 , new_n12790 , new_n12793 );
nor  g19297 ( new_n21646 , new_n21644 , new_n21645_1 );
and  g19298 ( new_n21647 , new_n21643 , new_n21646 );
nor  g19299 ( new_n21648 , new_n21642 , new_n21647 );
and  g19300 ( new_n21649_1 , new_n21641 , new_n21648 );
nor  g19301 ( new_n21650 , new_n21640 , new_n21649_1 );
nor  g19302 ( new_n21651 , new_n21639 , new_n21650 );
nor  g19303 ( new_n21652 , new_n21638 , new_n21651 );
nor  g19304 ( new_n21653 , new_n21637_1 , new_n21652 );
or   g19305 ( new_n21654_1 , new_n21636 , new_n21653 );
xor  g19306 ( new_n21655 , new_n21635 , new_n21654_1 );
xnor g19307 ( new_n21656 , new_n4837 , new_n21655 );
xnor g19308 ( new_n21657 , new_n21637_1 , new_n21652 );
nor  g19309 ( new_n21658 , new_n4841 , new_n21657 );
xnor g19310 ( new_n21659 , new_n4841 , new_n21657 );
xnor g19311 ( new_n21660 , new_n21639 , new_n21650 );
nor  g19312 ( new_n21661 , new_n4845 , new_n21660 );
xnor g19313 ( new_n21662 , new_n21641 , new_n21648 );
nor  g19314 ( new_n21663 , new_n4850_1 , new_n21662 );
not  g19315 ( new_n21664 , new_n21662 );
xnor g19316 ( new_n21665_1 , new_n4850_1 , new_n21664 );
xnor g19317 ( new_n21666 , n5337 , n22198 );
xnor g19318 ( new_n21667 , new_n21646 , new_n21666 );
nor  g19319 ( new_n21668 , new_n4854 , new_n21667 );
and  g19320 ( new_n21669 , new_n12789 , new_n12795 );
nor  g19321 ( new_n21670 , new_n4861 , new_n12796 );
nor  g19322 ( new_n21671 , new_n21669 , new_n21670 );
xor  g19323 ( new_n21672 , new_n4854 , new_n21667 );
and  g19324 ( new_n21673 , new_n21671 , new_n21672 );
or   g19325 ( new_n21674_1 , new_n21668 , new_n21673 );
and  g19326 ( new_n21675 , new_n21665_1 , new_n21674_1 );
nor  g19327 ( new_n21676 , new_n21663 , new_n21675 );
xnor g19328 ( new_n21677 , new_n4845 , new_n21660 );
nor  g19329 ( new_n21678 , new_n21676 , new_n21677 );
nor  g19330 ( new_n21679 , new_n21661 , new_n21678 );
nor  g19331 ( new_n21680_1 , new_n21659 , new_n21679 );
nor  g19332 ( new_n21681 , new_n21658 , new_n21680_1 );
xnor g19333 ( new_n21682 , new_n21656 , new_n21681 );
xnor g19334 ( new_n21683 , new_n17137 , new_n21682 );
xnor g19335 ( new_n21684 , new_n21659 , new_n21679 );
nor  g19336 ( new_n21685_1 , new_n16464 , new_n21684 );
xnor g19337 ( new_n21686 , new_n16464 , new_n21684 );
xnor g19338 ( new_n21687_1 , new_n21676 , new_n21677 );
nor  g19339 ( new_n21688 , new_n16469 , new_n21687_1 );
xnor g19340 ( new_n21689 , new_n16469 , new_n21687_1 );
xor  g19341 ( new_n21690 , new_n21665_1 , new_n21674_1 );
and  g19342 ( new_n21691 , new_n3771 , new_n21690 );
xnor g19343 ( new_n21692 , new_n3772 , new_n21690 );
xor  g19344 ( new_n21693 , new_n21671 , new_n21672 );
nor  g19345 ( new_n21694 , new_n3775 , new_n21693 );
and  g19346 ( new_n21695 , new_n3782 , new_n12797 );
and  g19347 ( new_n21696 , new_n12798 , new_n12806 );
nor  g19348 ( new_n21697 , new_n21695 , new_n21696 );
xnor g19349 ( new_n21698 , new_n3775 , new_n21693 );
nor  g19350 ( new_n21699 , new_n21697 , new_n21698 );
nor  g19351 ( new_n21700 , new_n21694 , new_n21699 );
and  g19352 ( new_n21701 , new_n21692 , new_n21700 );
nor  g19353 ( new_n21702 , new_n21691 , new_n21701 );
nor  g19354 ( new_n21703 , new_n21689 , new_n21702 );
nor  g19355 ( new_n21704 , new_n21688 , new_n21703 );
nor  g19356 ( new_n21705 , new_n21686 , new_n21704 );
nor  g19357 ( new_n21706 , new_n21685_1 , new_n21705 );
xor  g19358 ( n9968 , new_n21683 , new_n21706 );
nor  g19359 ( new_n21708 , new_n13678 , new_n20093 );
xor  g19360 ( new_n21709 , new_n13678 , new_n20093 );
nor  g19361 ( new_n21710 , new_n13678 , new_n20102 );
xnor g19362 ( new_n21711 , new_n13678 , new_n20101 );
and  g19363 ( new_n21712 , new_n11169 , new_n20095 );
and  g19364 ( new_n21713 , new_n11227 , new_n11267 );
nor  g19365 ( new_n21714 , new_n21712 , new_n21713 );
and  g19366 ( new_n21715 , new_n21711 , new_n21714 );
nor  g19367 ( new_n21716 , new_n21710 , new_n21715 );
and  g19368 ( new_n21717_1 , new_n21709 , new_n21716 );
nor  g19369 ( n10009 , new_n21708 , new_n21717_1 );
xnor g19370 ( n10010 , new_n20810 , new_n20813 );
and  g19371 ( new_n21720 , new_n10955 , new_n14513 );
and  g19372 ( new_n21721 , new_n14515 , new_n14544 );
nor  g19373 ( new_n21722 , new_n21720 , new_n21721 );
not  g19374 ( new_n21723 , new_n21722 );
nor  g19375 ( new_n21724 , new_n14586 , new_n21723 );
xnor g19376 ( new_n21725 , new_n14586 , new_n21722 );
and  g19377 ( new_n21726 , new_n14545 , new_n14586 );
and  g19378 ( new_n21727 , new_n14587 , new_n14626 );
or   g19379 ( new_n21728 , new_n21726 , new_n21727 );
and  g19380 ( new_n21729 , new_n21725 , new_n21728 );
nor  g19381 ( n10019 , new_n21724 , new_n21729 );
xnor g19382 ( n10021 , new_n14363 , new_n14411 );
xor  g19383 ( n10055 , new_n9553 , new_n9563 );
xnor g19384 ( n10101 , new_n10581 , new_n10603 );
xnor g19385 ( n10111 , new_n4556 , new_n4602 );
nor  g19386 ( new_n21735_1 , new_n20751 , n16544 );
xnor g19387 ( new_n21736 , n3324 , n16544 );
nor  g19388 ( new_n21737 , n6814 , new_n19668 );
xnor g19389 ( new_n21738 , n6814 , n17911 );
nor  g19390 ( new_n21739 , n19701 , new_n18472 );
xnor g19391 ( new_n21740 , n19701 , n21997 );
nor  g19392 ( new_n21741 , n23529 , new_n8501 );
xnor g19393 ( new_n21742 , n23529 , n25119 );
nor  g19394 ( new_n21743 , new_n8503 , n24620 );
xnor g19395 ( new_n21744 , n1163 , n24620 );
nor  g19396 ( new_n21745 , n5211 , new_n8506 );
or   g19397 ( new_n21746 , new_n8968 , n18537 );
nor  g19398 ( new_n21747 , n7057 , new_n8971_1 );
and  g19399 ( new_n21748 , new_n9442 , new_n9451_1 );
nor  g19400 ( new_n21749_1 , new_n21747 , new_n21748 );
and  g19401 ( new_n21750_1 , new_n21746 , new_n21749_1 );
or   g19402 ( new_n21751 , new_n21745 , new_n21750_1 );
and  g19403 ( new_n21752 , new_n21744 , new_n21751 );
or   g19404 ( new_n21753_1 , new_n21743 , new_n21752 );
and  g19405 ( new_n21754 , new_n21742 , new_n21753_1 );
or   g19406 ( new_n21755 , new_n21741 , new_n21754 );
and  g19407 ( new_n21756 , new_n21740 , new_n21755 );
or   g19408 ( new_n21757 , new_n21739 , new_n21756 );
and  g19409 ( new_n21758 , new_n21738 , new_n21757 );
or   g19410 ( new_n21759 , new_n21737 , new_n21758 );
and  g19411 ( new_n21760 , new_n21736 , new_n21759 );
nor  g19412 ( new_n21761 , new_n21735_1 , new_n21760 );
not  g19413 ( new_n21762 , new_n21761 );
xnor g19414 ( new_n21763 , new_n20950 , new_n21762 );
nor  g19415 ( new_n21764 , new_n20960 , new_n21762 );
nor  g19416 ( new_n21765_1 , new_n20959 , new_n21761 );
xor  g19417 ( new_n21766 , new_n21736 , new_n21759 );
nor  g19418 ( new_n21767 , new_n16979 , new_n21766 );
xnor g19419 ( new_n21768 , new_n16979 , new_n21766 );
xor  g19420 ( new_n21769 , new_n21738 , new_n21757 );
nor  g19421 ( new_n21770 , new_n17027 , new_n21769 );
xnor g19422 ( new_n21771 , new_n17027 , new_n21769 );
xor  g19423 ( new_n21772 , new_n21740 , new_n21755 );
nor  g19424 ( new_n21773 , new_n17034 , new_n21772 );
xnor g19425 ( new_n21774 , new_n17034 , new_n21772 );
xor  g19426 ( new_n21775 , new_n21742 , new_n21753_1 );
nor  g19427 ( new_n21776 , new_n17041 , new_n21775 );
xnor g19428 ( new_n21777 , new_n17041 , new_n21775 );
xor  g19429 ( new_n21778 , new_n21744 , new_n21751 );
nor  g19430 ( new_n21779_1 , new_n17046 , new_n21778 );
xnor g19431 ( new_n21780 , n5211 , n18537 );
xnor g19432 ( new_n21781 , new_n21749_1 , new_n21780 );
nor  g19433 ( new_n21782 , new_n17055 , new_n21781 );
xnor g19434 ( new_n21783 , new_n17052 , new_n21781 );
and  g19435 ( new_n21784_1 , new_n9441 , new_n9452 );
and  g19436 ( new_n21785 , new_n9453 , new_n9473 );
or   g19437 ( new_n21786 , new_n21784_1 , new_n21785 );
and  g19438 ( new_n21787 , new_n21783 , new_n21786 );
nor  g19439 ( new_n21788 , new_n21782 , new_n21787 );
xnor g19440 ( new_n21789 , new_n17045 , new_n21778 );
and  g19441 ( new_n21790 , new_n21788 , new_n21789 );
nor  g19442 ( new_n21791 , new_n21779_1 , new_n21790 );
nor  g19443 ( new_n21792 , new_n21777 , new_n21791 );
nor  g19444 ( new_n21793 , new_n21776 , new_n21792 );
nor  g19445 ( new_n21794 , new_n21774 , new_n21793 );
nor  g19446 ( new_n21795 , new_n21773 , new_n21794 );
nor  g19447 ( new_n21796 , new_n21771 , new_n21795 );
nor  g19448 ( new_n21797 , new_n21770 , new_n21796 );
nor  g19449 ( new_n21798 , new_n21768 , new_n21797 );
nor  g19450 ( new_n21799 , new_n21767 , new_n21798 );
not  g19451 ( new_n21800_1 , new_n21799 );
nor  g19452 ( new_n21801 , new_n21765_1 , new_n21800_1 );
nor  g19453 ( new_n21802 , new_n21764 , new_n21801 );
xnor g19454 ( n10165 , new_n21763 , new_n21802 );
xnor g19455 ( n10236 , new_n12873_1 , new_n12874 );
xnor g19456 ( n10239 , new_n14263 , new_n14285 );
xnor g19457 ( n10244 , new_n6375_1 , new_n6415 );
xnor g19458 ( n10261 , new_n17889_1 , new_n17901 );
xnor g19459 ( n10262 , new_n15525 , new_n15539_1 );
xnor g19460 ( n10287 , new_n16713 , new_n16714 );
nor  g19461 ( new_n21810 , new_n15096 , new_n21185 );
xnor g19462 ( new_n21811 , new_n21810 , new_n21227 );
nor  g19463 ( new_n21812 , new_n21186 , new_n21190 );
nor  g19464 ( new_n21813 , new_n21191 , new_n21204 );
nor  g19465 ( new_n21814 , new_n21812 , new_n21813 );
xnor g19466 ( n10295 , new_n21811 , new_n21814 );
xnor g19467 ( n10321 , new_n14722 , new_n14725 );
xnor g19468 ( n10326 , new_n14260 , new_n14287 );
xor  g19469 ( n10327 , new_n2820 , new_n2833 );
xnor g19470 ( new_n21819 , new_n20082 , new_n20102 );
xnor g19471 ( n10330 , new_n20104 , new_n21819 );
xnor g19472 ( n10340 , new_n20703 , new_n20736 );
xnor g19473 ( new_n21822 , new_n16708 , new_n16711 );
xnor g19474 ( n10345 , new_n16716 , new_n21822 );
nor  g19475 ( new_n21824 , new_n4897 , new_n13919 );
nor  g19476 ( new_n21825 , new_n21824 , new_n18896 );
not  g19477 ( new_n21826 , new_n4902 );
nor  g19478 ( new_n21827 , new_n21826 , new_n18899 );
xnor g19479 ( new_n21828 , new_n21826 , new_n18899 );
and  g19480 ( new_n21829 , new_n4904 , new_n18904 );
xnor g19481 ( new_n21830 , new_n4904 , new_n18904 );
and  g19482 ( new_n21831 , new_n4910 , new_n18908 );
xnor g19483 ( new_n21832_1 , new_n4910 , new_n18908 );
and  g19484 ( new_n21833 , new_n4914 , new_n18912 );
xnor g19485 ( new_n21834 , new_n4914 , new_n18912 );
nor  g19486 ( new_n21835 , new_n4920 , new_n9351 );
xnor g19487 ( new_n21836 , new_n4920 , new_n9351 );
nor  g19488 ( new_n21837 , new_n4925_1 , new_n9355 );
xnor g19489 ( new_n21838 , new_n4925_1 , new_n9355 );
nor  g19490 ( new_n21839_1 , new_n4930 , new_n9360 );
xnor g19491 ( new_n21840 , new_n4930 , new_n9360 );
nor  g19492 ( new_n21841 , new_n4950 , new_n9365 );
xnor g19493 ( new_n21842 , new_n4950 , new_n9365 );
nor  g19494 ( new_n21843 , new_n4936 , new_n9370 );
xnor g19495 ( new_n21844 , new_n4936 , new_n9370 );
nor  g19496 ( new_n21845 , new_n4943 , new_n9376 );
and  g19497 ( new_n21846 , new_n9373 , new_n21845 );
xnor g19498 ( new_n21847 , new_n9380_1 , new_n21845 );
and  g19499 ( new_n21848 , new_n4940 , new_n21847 );
nor  g19500 ( new_n21849 , new_n21846 , new_n21848 );
nor  g19501 ( new_n21850 , new_n21844 , new_n21849 );
nor  g19502 ( new_n21851 , new_n21843 , new_n21850 );
nor  g19503 ( new_n21852 , new_n21842 , new_n21851 );
nor  g19504 ( new_n21853 , new_n21841 , new_n21852 );
nor  g19505 ( new_n21854 , new_n21840 , new_n21853 );
nor  g19506 ( new_n21855 , new_n21839_1 , new_n21854 );
nor  g19507 ( new_n21856 , new_n21838 , new_n21855 );
nor  g19508 ( new_n21857 , new_n21837 , new_n21856 );
nor  g19509 ( new_n21858 , new_n21836 , new_n21857 );
nor  g19510 ( new_n21859 , new_n21835 , new_n21858 );
nor  g19511 ( new_n21860 , new_n21834 , new_n21859 );
nor  g19512 ( new_n21861 , new_n21833 , new_n21860 );
nor  g19513 ( new_n21862 , new_n21832_1 , new_n21861 );
nor  g19514 ( new_n21863 , new_n21831 , new_n21862 );
nor  g19515 ( new_n21864 , new_n21830 , new_n21863 );
nor  g19516 ( new_n21865 , new_n21829 , new_n21864 );
nor  g19517 ( new_n21866 , new_n21828 , new_n21865 );
nor  g19518 ( new_n21867 , new_n21827 , new_n21866 );
xnor g19519 ( new_n21868 , new_n21824 , new_n18895 );
and  g19520 ( new_n21869 , new_n21867 , new_n21868 );
nor  g19521 ( n10356 , new_n21825 , new_n21869 );
xor  g19522 ( n10385 , new_n19446 , new_n19447 );
nor  g19523 ( new_n21872 , new_n18895 , new_n19664_1 );
or   g19524 ( new_n21873 , new_n18896 , new_n19663 );
and  g19525 ( new_n21874_1 , new_n19609 , new_n21873 );
nor  g19526 ( new_n21875 , new_n21872 , new_n21874_1 );
nor  g19527 ( n10387 , new_n19607 , new_n21875 );
xnor g19528 ( n10388 , new_n19854 , new_n19867 );
xnor g19529 ( n10390 , new_n15280 , new_n15325 );
xnor g19530 ( n10404 , new_n9460_1 , new_n9461 );
xnor g19531 ( n10409 , new_n15700 , new_n15703 );
xnor g19532 ( n10420 , new_n8557 , new_n15907 );
xnor g19533 ( n10432 , new_n6946 , new_n17894 );
xnor g19534 ( new_n21883 , new_n20225 , new_n20903 );
nor  g19535 ( new_n21884 , new_n9600 , new_n20229 );
nor  g19536 ( new_n21885 , new_n20482 , new_n20489_1 );
nor  g19537 ( new_n21886 , new_n21884 , new_n21885 );
xnor g19538 ( new_n21887 , new_n21883 , new_n21886 );
xnor g19539 ( new_n21888 , new_n11380 , new_n21887 );
nor  g19540 ( new_n21889 , new_n11384 , new_n20490_1 );
nor  g19541 ( new_n21890 , new_n20491 , new_n20499 );
nor  g19542 ( new_n21891 , new_n21889 , new_n21890 );
xor  g19543 ( n10484 , new_n21888 , new_n21891 );
xnor g19544 ( n10489 , new_n11243 , new_n11256 );
xnor g19545 ( n10525 , new_n3641 , new_n13288 );
xor  g19546 ( new_n21895 , new_n11992 , new_n17271 );
xnor g19547 ( n10540 , new_n17279 , new_n21895 );
xnor g19548 ( n10561 , new_n15792 , new_n15816_1 );
xnor g19549 ( n10564 , new_n15272 , new_n15329 );
xnor g19550 ( n10588 , new_n9961 , new_n9963 );
xnor g19551 ( n10595 , new_n9964 , new_n9966 );
xor  g19552 ( n10617 , new_n20597 , new_n20609_1 );
xnor g19553 ( n10628 , new_n12254 , new_n12310 );
xnor g19554 ( new_n21903 , new_n5726 , new_n10549 );
nor  g19555 ( new_n21904 , new_n5729 , new_n10558 );
xnor g19556 ( new_n21905_1 , new_n5730 , new_n10557 );
and  g19557 ( new_n21906 , new_n5734 , new_n10561_1 );
xnor g19558 ( new_n21907 , new_n5734 , new_n10561_1 );
nor  g19559 ( new_n21908 , new_n5739 , new_n5769 );
nor  g19560 ( new_n21909 , new_n5779 , new_n21908 );
xnor g19561 ( new_n21910 , new_n5779 , new_n21908 );
nor  g19562 ( new_n21911 , new_n5746 , new_n21910 );
nor  g19563 ( new_n21912 , new_n21909 , new_n21911 );
nor  g19564 ( new_n21913 , new_n21907 , new_n21912 );
nor  g19565 ( new_n21914 , new_n21906 , new_n21913 );
nor  g19566 ( new_n21915_1 , new_n21905_1 , new_n21914 );
nor  g19567 ( new_n21916 , new_n21904 , new_n21915_1 );
xnor g19568 ( n10647 , new_n21903 , new_n21916 );
nor  g19569 ( new_n21918 , new_n8333 , new_n19318 );
not  g19570 ( new_n21919 , new_n21918 );
nor  g19571 ( new_n21920 , new_n3582_1 , new_n19344 );
and  g19572 ( new_n21921 , new_n3599 , new_n3661 );
or   g19573 ( new_n21922 , new_n19343 , new_n21921 );
or   g19574 ( new_n21923 , new_n21920 , new_n21922 );
nor  g19575 ( new_n21924 , new_n13257 , new_n21923 );
xnor g19576 ( new_n21925 , new_n21919 , new_n21924 );
not  g19577 ( new_n21926 , new_n8340 );
xor  g19578 ( new_n21927 , new_n13257 , new_n21923 );
nor  g19579 ( new_n21928 , new_n21926 , new_n21927 );
nor  g19580 ( new_n21929 , new_n3535 , new_n3662 );
nor  g19581 ( new_n21930 , new_n3663 , new_n3723 );
nor  g19582 ( new_n21931 , new_n21929 , new_n21930 );
xnor g19583 ( new_n21932 , new_n8340 , new_n21927 );
and  g19584 ( new_n21933 , new_n21931 , new_n21932 );
nor  g19585 ( new_n21934_1 , new_n21928 , new_n21933 );
xnor g19586 ( n10653 , new_n21925 , new_n21934_1 );
xnor g19587 ( n10692 , new_n9032_1 , new_n9033 );
xnor g19588 ( n10694 , new_n4302 , new_n14463 );
xnor g19589 ( n10701 , new_n19708 , new_n19731 );
xnor g19590 ( n10756 , new_n6118 , new_n6137 );
not  g19591 ( new_n21940 , n6659 );
nor  g19592 ( new_n21941 , n5101 , new_n21940 );
and  g19593 ( new_n21942 , new_n15666 , new_n15670 );
nor  g19594 ( new_n21943_1 , new_n21941 , new_n21942 );
not  g19595 ( new_n21944 , new_n21943_1 );
not  g19596 ( new_n21945 , n13419 );
and  g19597 ( new_n21946 , new_n21945 , new_n15671 );
nor  g19598 ( new_n21947 , new_n21945 , new_n15671 );
not  g19599 ( new_n21948 , n4967 );
and  g19600 ( new_n21949 , new_n21948 , new_n15626 );
nor  g19601 ( new_n21950 , new_n21948 , new_n15626 );
nor  g19602 ( new_n21951 , new_n21950 , new_n18822 );
nor  g19603 ( new_n21952 , new_n21949 , new_n21951 );
nor  g19604 ( new_n21953 , new_n21947 , new_n21952 );
nor  g19605 ( new_n21954 , new_n21946 , new_n21953 );
and  g19606 ( new_n21955 , new_n21944 , new_n21954 );
xnor g19607 ( new_n21956 , new_n3197 , new_n21955 );
xnor g19608 ( new_n21957_1 , new_n21943_1 , new_n21954 );
and  g19609 ( new_n21958 , new_n3329 , new_n21957_1 );
xnor g19610 ( new_n21959 , new_n3329 , new_n21957_1 );
xnor g19611 ( new_n21960_1 , new_n15672 , new_n21952 );
nor  g19612 ( new_n21961 , new_n3215 , new_n21960_1 );
xnor g19613 ( new_n21962 , new_n3215 , new_n21960_1 );
nor  g19614 ( new_n21963 , new_n3224 , new_n18823 );
nor  g19615 ( new_n21964 , new_n18824 , new_n18860 );
or   g19616 ( new_n21965 , new_n21963 , new_n21964 );
nor  g19617 ( new_n21966 , new_n21962 , new_n21965 );
nor  g19618 ( new_n21967 , new_n21961 , new_n21966 );
nor  g19619 ( new_n21968 , new_n21959 , new_n21967 );
nor  g19620 ( new_n21969 , new_n21958 , new_n21968 );
xnor g19621 ( n10775 , new_n21956 , new_n21969 );
xnor g19622 ( n10780 , new_n20517 , new_n20522 );
xnor g19623 ( new_n21972 , new_n16134 , n17095 );
nor  g19624 ( new_n21973 , n22274 , n22591 );
or   g19625 ( new_n21974 , new_n4122 , new_n9532 );
xnor g19626 ( new_n21975 , new_n4118 , n22591 );
and  g19627 ( new_n21976_1 , new_n21974 , new_n21975 );
or   g19628 ( new_n21977 , new_n21973 , new_n21976_1 );
xor  g19629 ( new_n21978 , new_n21972 , new_n21977 );
xnor g19630 ( new_n21979 , n21749 , new_n21978 );
nor  g19631 ( new_n21980 , new_n9485 , new_n8912 );
nor  g19632 ( new_n21981_1 , n7769 , new_n21980 );
xor  g19633 ( new_n21982 , new_n21974 , new_n21975 );
xnor g19634 ( new_n21983 , new_n9487 , new_n21980 );
not  g19635 ( new_n21984 , new_n21983 );
nor  g19636 ( new_n21985 , new_n21982 , new_n21984 );
nor  g19637 ( new_n21986_1 , new_n21981_1 , new_n21985 );
xnor g19638 ( new_n21987 , new_n21979 , new_n21986_1 );
xnor g19639 ( new_n21988 , new_n18061_1 , new_n21987 );
xnor g19640 ( new_n21989 , new_n21982 , new_n21983 );
and  g19641 ( new_n21990 , new_n18065 , new_n21989 );
nor  g19642 ( new_n21991 , new_n18068 , new_n8913 );
xnor g19643 ( new_n21992 , new_n18064 , new_n21989 );
and  g19644 ( new_n21993_1 , new_n21991 , new_n21992 );
or   g19645 ( new_n21994 , new_n21990 , new_n21993_1 );
xor  g19646 ( n10817 , new_n21988 , new_n21994 );
not  g19647 ( new_n21996 , new_n21210 );
and  g19648 ( new_n21997_1 , new_n21996 , new_n21214 );
and  g19649 ( new_n21998 , new_n21206 , new_n21209 );
nor  g19650 ( new_n21999 , new_n21996 , new_n21214 );
nor  g19651 ( new_n22000 , new_n21999 , new_n21218 );
or   g19652 ( new_n22001 , new_n21998 , new_n22000 );
nor  g19653 ( new_n22002 , new_n21997_1 , new_n22001 );
nor  g19654 ( new_n22003 , new_n7694 , new_n22002 );
nor  g19655 ( new_n22004 , new_n7694 , new_n21219 );
nor  g19656 ( new_n22005 , new_n21221 , new_n21224 );
nor  g19657 ( new_n22006 , new_n22004 , new_n22005 );
not  g19658 ( new_n22007 , new_n22002 );
xnor g19659 ( new_n22008 , new_n7694 , new_n22007 );
and  g19660 ( new_n22009 , new_n22006 , new_n22008 );
nor  g19661 ( n10834 , new_n22003 , new_n22009 );
xor  g19662 ( n10851 , new_n21435 , new_n21452 );
xnor g19663 ( n10874 , new_n20994 , new_n21003 );
xor  g19664 ( new_n22013 , new_n21620 , new_n21628_1 );
xnor g19665 ( n10924 , new_n8028 , new_n22013 );
nor  g19666 ( new_n22015 , new_n11021 , new_n11025_1 );
and  g19667 ( new_n22016_1 , new_n11027 , new_n11090 );
nor  g19668 ( n10943 , new_n22015 , new_n22016_1 );
xnor g19669 ( n10961 , new_n11752 , new_n11785 );
xnor g19670 ( n11005 , new_n10487 , new_n10499 );
xnor g19671 ( n11023 , new_n20774_1 , new_n20782 );
nor  g19672 ( new_n22021 , new_n7263 , new_n17749_1 );
xnor g19673 ( new_n22022 , new_n7263 , new_n17749_1 );
nor  g19674 ( new_n22023 , new_n7269 , new_n17751 );
xnor g19675 ( new_n22024 , new_n7269 , new_n17751 );
nor  g19676 ( new_n22025 , new_n14657 , new_n16518 );
xnor g19677 ( new_n22026 , new_n14657 , new_n16518 );
and  g19678 ( new_n22027_1 , new_n7278 , new_n11951 );
nor  g19679 ( new_n22028 , new_n11952 , new_n11976 );
nor  g19680 ( new_n22029 , new_n22027_1 , new_n22028 );
nor  g19681 ( new_n22030 , new_n22026 , new_n22029 );
or   g19682 ( new_n22031 , new_n22025 , new_n22030 );
nor  g19683 ( new_n22032 , new_n22024 , new_n22031 );
nor  g19684 ( new_n22033 , new_n22023 , new_n22032 );
nor  g19685 ( new_n22034 , new_n22022 , new_n22033 );
nor  g19686 ( new_n22035 , new_n22021 , new_n22034 );
or   g19687 ( new_n22036 , new_n7241 , new_n22035 );
nor  g19688 ( new_n22037 , new_n17776 , new_n22036 );
not  g19689 ( new_n22038 , new_n21585 );
xnor g19690 ( new_n22039 , new_n7241 , new_n22035 );
xnor g19691 ( new_n22040 , new_n17776 , new_n22039 );
and  g19692 ( new_n22041 , new_n22038 , new_n22040 );
xnor g19693 ( new_n22042 , new_n22038 , new_n22040 );
xnor g19694 ( new_n22043_1 , new_n22022 , new_n22033 );
nor  g19695 ( new_n22044 , new_n21591 , new_n22043_1 );
xnor g19696 ( new_n22045 , new_n21591 , new_n22043_1 );
xnor g19697 ( new_n22046 , new_n22024 , new_n22031 );
nor  g19698 ( new_n22047 , new_n21596 , new_n22046 );
xnor g19699 ( new_n22048 , new_n21596 , new_n22046 );
xor  g19700 ( new_n22049 , new_n22026 , new_n22029 );
nor  g19701 ( new_n22050_1 , new_n17257 , new_n22049 );
xnor g19702 ( new_n22051 , new_n17257 , new_n22049 );
nor  g19703 ( new_n22052 , new_n11946 , new_n11977 );
nor  g19704 ( new_n22053 , new_n11978 , new_n12014 );
nor  g19705 ( new_n22054 , new_n22052 , new_n22053 );
nor  g19706 ( new_n22055 , new_n22051 , new_n22054 );
nor  g19707 ( new_n22056 , new_n22050_1 , new_n22055 );
nor  g19708 ( new_n22057 , new_n22048 , new_n22056 );
nor  g19709 ( new_n22058 , new_n22047 , new_n22057 );
nor  g19710 ( new_n22059 , new_n22045 , new_n22058 );
nor  g19711 ( new_n22060 , new_n22044 , new_n22059 );
nor  g19712 ( new_n22061 , new_n22042 , new_n22060 );
or   g19713 ( new_n22062 , new_n22041 , new_n22061 );
and  g19714 ( new_n22063_1 , new_n22037 , new_n22062 );
xor  g19715 ( new_n22064 , new_n22037 , new_n22062 );
nor  g19716 ( new_n22065 , new_n21613 , new_n22064 );
or   g19717 ( n11025 , new_n22063_1 , new_n22065 );
xnor g19718 ( new_n22067 , n21915 , new_n16154 );
nor  g19719 ( new_n22068_1 , new_n6836 , new_n16157 );
xnor g19720 ( new_n22069 , n13775 , new_n16157 );
nor  g19721 ( new_n22070 , new_n6839 , new_n16160 );
xnor g19722 ( new_n22071 , n1293 , new_n16160 );
nor  g19723 ( new_n22072_1 , new_n6842 , new_n16163 );
and  g19724 ( new_n22073 , new_n18701 , new_n18704 );
or   g19725 ( new_n22074 , new_n22072_1 , new_n22073 );
and  g19726 ( new_n22075 , new_n22071 , new_n22074 );
or   g19727 ( new_n22076_1 , new_n22070 , new_n22075 );
and  g19728 ( new_n22077 , new_n22069 , new_n22076_1 );
or   g19729 ( new_n22078 , new_n22068_1 , new_n22077 );
xor  g19730 ( new_n22079 , new_n22067 , new_n22078 );
not  g19731 ( new_n22080 , new_n18707 );
nor  g19732 ( new_n22081 , n26752 , new_n22080 );
not  g19733 ( new_n22082 , new_n22081 );
nor  g19734 ( new_n22083 , n4590 , new_n22082 );
not  g19735 ( new_n22084 , new_n22083 );
nor  g19736 ( new_n22085 , n25464 , new_n22084 );
xnor g19737 ( new_n22086 , n3795 , new_n22085 );
xnor g19738 ( new_n22087 , new_n8788 , new_n22086 );
xnor g19739 ( new_n22088 , n25464 , new_n22083 );
nor  g19740 ( new_n22089 , new_n8795 , new_n22088 );
xnor g19741 ( new_n22090_1 , new_n8795 , new_n22088 );
xnor g19742 ( new_n22091 , n4590 , new_n22081 );
nor  g19743 ( new_n22092 , new_n8801 , new_n22091 );
xnor g19744 ( new_n22093 , new_n8801 , new_n22091 );
nor  g19745 ( new_n22094 , new_n8807 , new_n18708_1 );
nor  g19746 ( new_n22095 , new_n18709 , new_n18712 );
nor  g19747 ( new_n22096 , new_n22094 , new_n22095 );
nor  g19748 ( new_n22097 , new_n22093 , new_n22096 );
nor  g19749 ( new_n22098 , new_n22092 , new_n22097 );
nor  g19750 ( new_n22099 , new_n22090_1 , new_n22098 );
nor  g19751 ( new_n22100 , new_n22089 , new_n22099 );
xnor g19752 ( new_n22101 , new_n22087 , new_n22100 );
xnor g19753 ( new_n22102 , new_n22079 , new_n22101 );
xor  g19754 ( new_n22103 , new_n22069 , new_n22076_1 );
xnor g19755 ( new_n22104 , new_n22090_1 , new_n22098 );
nor  g19756 ( new_n22105 , new_n22103 , new_n22104 );
xnor g19757 ( new_n22106 , new_n22103 , new_n22104 );
xor  g19758 ( new_n22107_1 , new_n22071 , new_n22074 );
xnor g19759 ( new_n22108 , new_n22093 , new_n22096 );
nor  g19760 ( new_n22109 , new_n22107_1 , new_n22108 );
xnor g19761 ( new_n22110 , new_n22107_1 , new_n22108 );
nor  g19762 ( new_n22111 , new_n18705 , new_n18713 );
nor  g19763 ( new_n22112 , new_n18714 , new_n18717 );
nor  g19764 ( new_n22113_1 , new_n22111 , new_n22112 );
nor  g19765 ( new_n22114 , new_n22110 , new_n22113_1 );
nor  g19766 ( new_n22115 , new_n22109 , new_n22114 );
nor  g19767 ( new_n22116 , new_n22106 , new_n22115 );
nor  g19768 ( new_n22117 , new_n22105 , new_n22116 );
xnor g19769 ( n11063 , new_n22102 , new_n22117 );
xnor g19770 ( n11078 , new_n19857 , new_n19865 );
xnor g19771 ( n11080 , new_n20514 , new_n20524 );
xnor g19772 ( n11094 , new_n13571 , new_n13584 );
xnor g19773 ( n11101 , new_n21788 , new_n21789 );
xnor g19774 ( new_n22123 , new_n14139 , new_n20602_1 );
xnor g19775 ( n11103 , new_n20605 , new_n22123 );
xnor g19776 ( n11120 , new_n6556_1 , new_n6581 );
xor  g19777 ( n11127 , new_n5007 , new_n5010 );
xnor g19778 ( n11132 , new_n14727 , new_n14728 );
xnor g19779 ( n11134 , new_n11038 , new_n11083 );
xnor g19780 ( n11138 , new_n3706 , new_n3707 );
xnor g19781 ( n11182 , new_n10381 , new_n10391 );
xnor g19782 ( n11234 , new_n13556 , new_n13594 );
xnor g19783 ( new_n22132 , new_n18226 , new_n21186 );
nor  g19784 ( new_n22133 , new_n18230 , new_n21193_1 );
nor  g19785 ( new_n22134 , new_n20848 , new_n20869_1 );
nor  g19786 ( new_n22135 , new_n22133 , new_n22134 );
xnor g19787 ( n11245 , new_n22132 , new_n22135 );
xnor g19788 ( n11261 , new_n8627 , new_n8641 );
xnor g19789 ( n11275 , new_n22106 , new_n22115 );
nand g19790 ( n11290 , new_n13251 , new_n13310 );
xnor g19791 ( n11313 , new_n9379 , new_n9381 );
xnor g19792 ( new_n22141 , new_n15936_1 , new_n16494 );
xnor g19793 ( n11325 , new_n16508 , new_n22141 );
xnor g19794 ( n11326 , new_n13635 , new_n13636 );
xnor g19795 ( n11330 , new_n16692 , new_n16724 );
xnor g19796 ( n11347 , new_n11049 , new_n11077 );
xnor g19797 ( n11348 , new_n21844 , new_n21849 );
xnor g19798 ( n11352 , new_n14830 , new_n14838 );
nor  g19799 ( new_n22148 , n3324 , new_n8271 );
xnor g19800 ( new_n22149 , n3324 , n22442 );
nor  g19801 ( new_n22150_1 , new_n8273 , n17911 );
nor  g19802 ( new_n22151 , new_n8280 , n21997 );
and  g19803 ( new_n22152 , new_n16908 , new_n16915 );
or   g19804 ( new_n22153 , new_n22151 , new_n22152 );
xnor g19805 ( new_n22154 , n468 , n17911 );
and  g19806 ( new_n22155 , new_n22153 , new_n22154 );
or   g19807 ( new_n22156 , new_n22150_1 , new_n22155 );
and  g19808 ( new_n22157_1 , new_n22149 , new_n22156 );
nor  g19809 ( new_n22158 , new_n22148 , new_n22157_1 );
not  g19810 ( new_n22159 , new_n22158 );
and  g19811 ( new_n22160 , new_n17419 , new_n17425 );
nor  g19812 ( new_n22161 , new_n7649 , new_n22160 );
nor  g19813 ( new_n22162 , new_n17419 , new_n17425 );
nor  g19814 ( new_n22163 , new_n7650 , new_n22162 );
nor  g19815 ( new_n22164 , new_n22161 , new_n22163 );
xnor g19816 ( new_n22165 , new_n22159 , new_n22164 );
nor  g19817 ( new_n22166 , new_n17427 , new_n22159 );
nor  g19818 ( new_n22167 , new_n17428 , new_n22158 );
xor  g19819 ( new_n22168 , new_n22149 , new_n22156 );
nor  g19820 ( new_n22169 , new_n17430 , new_n22168 );
xnor g19821 ( new_n22170 , new_n17430 , new_n22168 );
not  g19822 ( new_n22171 , new_n22170 );
xor  g19823 ( new_n22172 , new_n22153 , new_n22154 );
and  g19824 ( new_n22173_1 , new_n17433 , new_n22172 );
xnor g19825 ( new_n22174 , new_n17432_1 , new_n22172 );
and  g19826 ( new_n22175 , new_n17436_1 , new_n16916 );
and  g19827 ( new_n22176 , new_n16917 , new_n16927 );
or   g19828 ( new_n22177 , new_n22175 , new_n22176 );
and  g19829 ( new_n22178 , new_n22174 , new_n22177 );
nor  g19830 ( new_n22179 , new_n22173_1 , new_n22178 );
and  g19831 ( new_n22180 , new_n22171 , new_n22179 );
nor  g19832 ( new_n22181 , new_n22169 , new_n22180 );
not  g19833 ( new_n22182 , new_n22181 );
nor  g19834 ( new_n22183 , new_n22167 , new_n22182 );
nor  g19835 ( new_n22184 , new_n22166 , new_n22183 );
xnor g19836 ( n11375 , new_n22165 , new_n22184 );
xnor g19837 ( n11379 , new_n7158 , new_n12337 );
nor  g19838 ( new_n22187 , n2570 , new_n11795 );
and  g19839 ( new_n22188 , new_n16122 , new_n16151 );
nor  g19840 ( new_n22189 , new_n22187 , new_n22188 );
xnor g19841 ( new_n22190 , new_n11846 , new_n22189 );
nor  g19842 ( new_n22191 , new_n11802 , new_n16152 );
nor  g19843 ( new_n22192 , new_n16153 , new_n16188 );
or   g19844 ( new_n22193 , new_n22191 , new_n22192 );
xor  g19845 ( new_n22194 , new_n22190 , new_n22193 );
xnor g19846 ( new_n22195 , new_n6356_1 , new_n22194 );
nor  g19847 ( new_n22196 , new_n6361 , new_n16189 );
nor  g19848 ( new_n22197 , new_n16190 , new_n16225 );
nor  g19849 ( new_n22198_1 , new_n22196 , new_n22197 );
xnor g19850 ( n11386 , new_n22195 , new_n22198_1 );
xnor g19851 ( n11391 , new_n18839 , new_n18850 );
xnor g19852 ( n11398 , new_n20832 , new_n20833 );
xnor g19853 ( n11403 , new_n12643 , new_n12644 );
xnor g19854 ( n11419 , new_n12082 , new_n12087 );
xnor g19855 ( n11439 , new_n18675 , new_n18690_1 );
xnor g19856 ( new_n22205 , n2570 , new_n11325_1 );
nor  g19857 ( new_n22206 , n17037 , n19033 );
xnor g19858 ( new_n22207 , n17037 , n19033 );
nor  g19859 ( new_n22208 , n655 , n5386 );
xnor g19860 ( new_n22209 , n655 , n5386 );
nor  g19861 ( new_n22210 , n18145 , n26191 );
xnor g19862 ( new_n22211 , n18145 , n26191 );
nor  g19863 ( new_n22212 , n10712 , n26512 );
xnor g19864 ( new_n22213_1 , n10712 , n26512 );
nor  g19865 ( new_n22214 , n19575 , n25126 );
xnor g19866 ( new_n22215 , new_n15732 , n25126 );
and  g19867 ( new_n22216 , n15378 , n19608 );
or   g19868 ( new_n22217 , n15378 , n19608 );
nor  g19869 ( new_n22218 , n1689 , n17095 );
and  g19870 ( new_n22219 , new_n21972 , new_n21977 );
nor  g19871 ( new_n22220 , new_n22218 , new_n22219 );
and  g19872 ( new_n22221 , new_n22217 , new_n22220 );
nor  g19873 ( new_n22222 , new_n22216 , new_n22221 );
and  g19874 ( new_n22223 , new_n22215 , new_n22222 );
nor  g19875 ( new_n22224 , new_n22214 , new_n22223 );
nor  g19876 ( new_n22225 , new_n22213_1 , new_n22224 );
nor  g19877 ( new_n22226 , new_n22212 , new_n22225 );
nor  g19878 ( new_n22227 , new_n22211 , new_n22226 );
nor  g19879 ( new_n22228 , new_n22210 , new_n22227 );
nor  g19880 ( new_n22229 , new_n22209 , new_n22228 );
nor  g19881 ( new_n22230 , new_n22208 , new_n22229 );
nor  g19882 ( new_n22231 , new_n22207 , new_n22230 );
or   g19883 ( new_n22232 , new_n22206 , new_n22231 );
xor  g19884 ( new_n22233 , new_n22205 , new_n22232 );
nor  g19885 ( new_n22234 , n10514 , new_n22233 );
xnor g19886 ( new_n22235 , new_n20222 , new_n22233 );
xnor g19887 ( new_n22236 , new_n22207 , new_n22230 );
nor  g19888 ( new_n22237 , new_n11276 , new_n22236 );
xnor g19889 ( new_n22238 , new_n11276 , new_n22236 );
xnor g19890 ( new_n22239 , new_n22209 , new_n22228 );
nor  g19891 ( new_n22240 , new_n11389 , new_n22239 );
xnor g19892 ( new_n22241 , new_n11389 , new_n22239 );
xnor g19893 ( new_n22242 , new_n22211 , new_n22226 );
nor  g19894 ( new_n22243 , new_n10824 , new_n22242 );
xnor g19895 ( new_n22244 , new_n10824 , new_n22242 );
xnor g19896 ( new_n22245 , new_n22213_1 , new_n22224 );
nor  g19897 ( new_n22246 , new_n10837 , new_n22245 );
xnor g19898 ( new_n22247 , new_n10837 , new_n22245 );
xnor g19899 ( new_n22248 , new_n22215 , new_n22222 );
nor  g19900 ( new_n22249 , new_n20239 , new_n22248 );
xnor g19901 ( new_n22250 , n9832 , new_n22248 );
xnor g19902 ( new_n22251 , new_n15736 , n19608 );
xnor g19903 ( new_n22252 , new_n22220 , new_n22251 );
nor  g19904 ( new_n22253_1 , n1558 , new_n22252 );
xnor g19905 ( new_n22254 , new_n9479 , new_n22252 );
nor  g19906 ( new_n22255 , n21749 , new_n21978 );
nor  g19907 ( new_n22256 , new_n21979 , new_n21986_1 );
or   g19908 ( new_n22257 , new_n22255 , new_n22256 );
and  g19909 ( new_n22258 , new_n22254 , new_n22257 );
nor  g19910 ( new_n22259 , new_n22253_1 , new_n22258 );
and  g19911 ( new_n22260 , new_n22250 , new_n22259 );
nor  g19912 ( new_n22261 , new_n22249 , new_n22260 );
nor  g19913 ( new_n22262 , new_n22247 , new_n22261 );
nor  g19914 ( new_n22263 , new_n22246 , new_n22262 );
nor  g19915 ( new_n22264 , new_n22244 , new_n22263 );
nor  g19916 ( new_n22265 , new_n22243 , new_n22264 );
nor  g19917 ( new_n22266 , new_n22241 , new_n22265 );
nor  g19918 ( new_n22267 , new_n22240 , new_n22266 );
nor  g19919 ( new_n22268 , new_n22238 , new_n22267 );
nor  g19920 ( new_n22269 , new_n22237 , new_n22268 );
and  g19921 ( new_n22270_1 , new_n22235 , new_n22269 );
nor  g19922 ( new_n22271 , new_n22234 , new_n22270_1 );
nor  g19923 ( new_n22272 , n2570 , n7569 );
and  g19924 ( new_n22273 , new_n22205 , new_n22232 );
or   g19925 ( new_n22274_1 , new_n22272 , new_n22273 );
xor  g19926 ( new_n22275 , new_n22271 , new_n22274_1 );
not  g19927 ( new_n22276 , new_n22085 );
nor  g19928 ( new_n22277 , n3795 , new_n22276 );
not  g19929 ( new_n22278 , new_n22277 );
nor  g19930 ( new_n22279 , n6105 , new_n22278 );
xnor g19931 ( new_n22280 , new_n11026 , new_n22279 );
xnor g19932 ( new_n22281 , n6105 , new_n22277 );
nor  g19933 ( new_n22282 , new_n8718 , new_n22281 );
xnor g19934 ( new_n22283_1 , new_n11032 , new_n22281 );
nor  g19935 ( new_n22284 , new_n8788 , new_n22086 );
nor  g19936 ( new_n22285 , new_n22087 , new_n22100 );
or   g19937 ( new_n22286 , new_n22284 , new_n22285 );
and  g19938 ( new_n22287 , new_n22283_1 , new_n22286 );
nor  g19939 ( new_n22288 , new_n22282 , new_n22287 );
xnor g19940 ( new_n22289 , new_n22280 , new_n22288 );
not  g19941 ( new_n22290_1 , new_n22289 );
xnor g19942 ( new_n22291 , new_n22275 , new_n22290_1 );
xnor g19943 ( new_n22292 , new_n22235 , new_n22269 );
nor  g19944 ( new_n22293 , new_n22284 , new_n22285 );
xnor g19945 ( new_n22294 , new_n22283_1 , new_n22293 );
and  g19946 ( new_n22295 , new_n22292 , new_n22294 );
xnor g19947 ( new_n22296 , new_n22292 , new_n22294 );
xnor g19948 ( new_n22297 , new_n22238 , new_n22267 );
nor  g19949 ( new_n22298 , new_n22101 , new_n22297 );
xnor g19950 ( new_n22299 , new_n22101 , new_n22297 );
xnor g19951 ( new_n22300 , new_n22241 , new_n22265 );
nor  g19952 ( new_n22301 , new_n22104 , new_n22300 );
xnor g19953 ( new_n22302 , new_n22104 , new_n22300 );
xnor g19954 ( new_n22303 , new_n22244 , new_n22263 );
nor  g19955 ( new_n22304 , new_n22108 , new_n22303 );
xnor g19956 ( new_n22305 , new_n22108 , new_n22303 );
xnor g19957 ( new_n22306 , new_n22247 , new_n22261 );
nor  g19958 ( new_n22307 , new_n18713 , new_n22306 );
xnor g19959 ( new_n22308 , new_n18713 , new_n22306 );
xnor g19960 ( new_n22309_1 , new_n22250 , new_n22259 );
nor  g19961 ( new_n22310 , new_n18039 , new_n22309_1 );
xnor g19962 ( new_n22311_1 , new_n18039 , new_n22309_1 );
xor  g19963 ( new_n22312 , new_n22254 , new_n22257 );
nor  g19964 ( new_n22313 , new_n18057 , new_n22312 );
not  g19965 ( new_n22314 , new_n18061_1 );
nor  g19966 ( new_n22315 , new_n22314 , new_n21987 );
and  g19967 ( new_n22316 , new_n21988 , new_n21994 );
nor  g19968 ( new_n22317_1 , new_n22315 , new_n22316 );
xnor g19969 ( new_n22318 , new_n18057 , new_n22312 );
not  g19970 ( new_n22319 , new_n22318 );
and  g19971 ( new_n22320 , new_n22317_1 , new_n22319 );
nor  g19972 ( new_n22321 , new_n22313 , new_n22320 );
nor  g19973 ( new_n22322 , new_n22311_1 , new_n22321 );
nor  g19974 ( new_n22323 , new_n22310 , new_n22322 );
nor  g19975 ( new_n22324 , new_n22308 , new_n22323 );
nor  g19976 ( new_n22325 , new_n22307 , new_n22324 );
nor  g19977 ( new_n22326 , new_n22305 , new_n22325 );
nor  g19978 ( new_n22327 , new_n22304 , new_n22326 );
nor  g19979 ( new_n22328 , new_n22302 , new_n22327 );
nor  g19980 ( new_n22329 , new_n22301 , new_n22328 );
nor  g19981 ( new_n22330 , new_n22299 , new_n22329 );
nor  g19982 ( new_n22331 , new_n22298 , new_n22330 );
nor  g19983 ( new_n22332_1 , new_n22296 , new_n22331 );
nor  g19984 ( new_n22333 , new_n22295 , new_n22332_1 );
xnor g19985 ( n11462 , new_n22291 , new_n22333 );
xnor g19986 ( n11470 , new_n19848 , new_n19871 );
xnor g19987 ( n11472 , new_n15143 , new_n15157 );
xnor g19988 ( new_n22337 , new_n7323 , new_n18533 );
xnor g19989 ( n11496 , new_n18547 , new_n22337 );
xnor g19990 ( n11506 , new_n19623_1 , new_n19655 );
xnor g19991 ( new_n22340 , new_n5710 , new_n21349_1 );
nor  g19992 ( new_n22341_1 , new_n5714 , new_n15486 );
xnor g19993 ( new_n22342 , new_n5714 , new_n15486 );
nor  g19994 ( new_n22343 , new_n5718 , new_n10526 );
xnor g19995 ( new_n22344 , new_n5718 , new_n10526 );
nor  g19996 ( new_n22345 , new_n5722 , new_n10544 );
xnor g19997 ( new_n22346 , new_n5722 , new_n10544 );
nor  g19998 ( new_n22347 , new_n5726 , new_n10549 );
nor  g19999 ( new_n22348 , new_n21903 , new_n21916 );
nor  g20000 ( new_n22349 , new_n22347 , new_n22348 );
nor  g20001 ( new_n22350 , new_n22346 , new_n22349 );
nor  g20002 ( new_n22351 , new_n22345 , new_n22350 );
nor  g20003 ( new_n22352 , new_n22344 , new_n22351 );
nor  g20004 ( new_n22353_1 , new_n22343 , new_n22352 );
nor  g20005 ( new_n22354 , new_n22342 , new_n22353_1 );
nor  g20006 ( new_n22355 , new_n22341_1 , new_n22354 );
xnor g20007 ( n11515 , new_n22340 , new_n22355 );
xnor g20008 ( n11538 , new_n20504 , new_n20534 );
xnor g20009 ( n11548 , new_n18330 , new_n18331 );
xnor g20010 ( n11564 , new_n18572_1 , new_n18577 );
nor  g20011 ( new_n22360 , n8856 , new_n8271 );
and  g20012 ( new_n22361 , new_n21246 , new_n21249 );
nor  g20013 ( new_n22362 , new_n22360 , new_n22361 );
nor  g20014 ( new_n22363 , n2272 , n3324 );
and  g20015 ( new_n22364 , new_n21251 , new_n21254_1 );
nor  g20016 ( new_n22365 , new_n22363 , new_n22364 );
nor  g20017 ( new_n22366 , new_n7500 , new_n22365 );
nor  g20018 ( new_n22367 , new_n7522 , new_n21255 );
nor  g20019 ( new_n22368 , new_n21256 , new_n21259 );
nor  g20020 ( new_n22369 , new_n22367 , new_n22368 );
xnor g20021 ( new_n22370 , new_n7499 , new_n22365 );
and  g20022 ( new_n22371 , new_n22369 , new_n22370 );
nor  g20023 ( new_n22372 , new_n22366 , new_n22371 );
not  g20024 ( new_n22373 , new_n22372 );
xnor g20025 ( new_n22374 , new_n22362 , new_n22373 );
xnor g20026 ( new_n22375 , new_n22369 , new_n22370 );
nor  g20027 ( new_n22376 , new_n22362 , new_n22375 );
not  g20028 ( new_n22377 , new_n22375 );
xnor g20029 ( new_n22378 , new_n22362 , new_n22377 );
not  g20030 ( new_n22379_1 , new_n21260 );
and  g20031 ( new_n22380 , new_n21250 , new_n22379_1 );
and  g20032 ( new_n22381 , new_n21261 , new_n21264 );
nor  g20033 ( new_n22382 , new_n22380 , new_n22381 );
and  g20034 ( new_n22383 , new_n22378 , new_n22382 );
nor  g20035 ( new_n22384 , new_n22376 , new_n22383 );
xnor g20036 ( n11591 , new_n22374 , new_n22384 );
or   g20037 ( new_n22386 , new_n8320_1 , new_n8327 );
nor  g20038 ( new_n22387 , new_n8329 , new_n21926 );
nor  g20039 ( new_n22388 , new_n8328 , new_n8340 );
nor  g20040 ( new_n22389 , new_n22388 , new_n8391 );
or   g20041 ( new_n22390 , new_n21918 , new_n22389 );
nor  g20042 ( new_n22391 , new_n22387 , new_n22390 );
and  g20043 ( n11607 , new_n22386 , new_n22391 );
xnor g20044 ( n11647 , new_n18249 , new_n18274_1 );
xor  g20045 ( n11674 , new_n22174 , new_n22177 );
xnor g20046 ( new_n22395 , new_n20185 , new_n19155 );
nor  g20047 ( new_n22396 , new_n20185 , new_n19167 );
and  g20048 ( new_n22397 , new_n20824 , new_n20835 );
or   g20049 ( new_n22398 , new_n22396 , new_n22397 );
xor  g20050 ( n11682 , new_n22395 , new_n22398 );
xor  g20051 ( n11710 , new_n21439 , new_n21450 );
xnor g20052 ( n11712 , new_n13565 , new_n13588 );
xnor g20053 ( n11724 , new_n21118 , new_n21131 );
xnor g20054 ( n11741 , new_n17720 , new_n17721_1 );
not  g20055 ( new_n22404 , new_n3064 );
xnor g20056 ( n11770 , new_n22404 , new_n17476 );
xnor g20057 ( n11771 , new_n8377 , new_n8378 );
xnor g20058 ( n11818 , new_n18411 , new_n18440 );
xnor g20059 ( n11837 , new_n21907 , new_n21912 );
not  g20060 ( new_n22409 , new_n15833 );
nor  g20061 ( new_n22410 , n7026 , new_n22409 );
xnor g20062 ( new_n22411 , n2743 , new_n22410 );
and  g20063 ( new_n22412 , new_n5914 , new_n22411 );
xnor g20064 ( new_n22413 , new_n5915 , new_n22411 );
and  g20065 ( new_n22414 , new_n5919 , new_n15834 );
and  g20066 ( new_n22415 , new_n15835 , new_n15872 );
or   g20067 ( new_n22416 , new_n22414 , new_n22415 );
and  g20068 ( new_n22417 , new_n22413 , new_n22416 );
nor  g20069 ( new_n22418 , new_n22412 , new_n22417 );
not  g20070 ( new_n22419 , new_n22418 );
and  g20071 ( new_n22420 , new_n13254 , new_n22410 );
xnor g20072 ( new_n22421 , new_n13193 , new_n22420 );
xnor g20073 ( new_n22422 , new_n22419 , new_n22421 );
xnor g20074 ( new_n22423 , new_n21190 , new_n22422 );
xor  g20075 ( new_n22424 , new_n22413 , new_n22416 );
nor  g20076 ( new_n22425 , new_n21192 , new_n22424 );
xnor g20077 ( new_n22426 , new_n21192 , new_n22424 );
nor  g20078 ( new_n22427 , new_n15873 , new_n15883 );
nor  g20079 ( new_n22428 , new_n15884_1 , new_n15923 );
nor  g20080 ( new_n22429 , new_n22427 , new_n22428 );
nor  g20081 ( new_n22430 , new_n22426 , new_n22429 );
nor  g20082 ( new_n22431 , new_n22425 , new_n22430 );
xnor g20083 ( n11842 , new_n22423 , new_n22431 );
xnor g20084 ( n11843 , new_n15434 , new_n15451 );
xnor g20085 ( n11905 , new_n18059_1 , new_n18075 );
xnor g20086 ( n11965 , new_n11246 , new_n11251 );
xnor g20087 ( n12000 , new_n17963_1 , new_n17966 );
xor  g20088 ( n12003 , new_n15993 , new_n15996 );
xnor g20089 ( n12011 , new_n16576 , new_n16577 );
xnor g20090 ( n12072 , new_n17056 , new_n17070_1 );
xor  g20091 ( n12131 , new_n10599 , new_n10601 );
xor  g20092 ( n12146 , new_n15941 , new_n15971 );
xnor g20093 ( n12157 , new_n16210 , new_n16213 );
xnor g20094 ( n12158 , new_n10108 , new_n10159 );
xnor g20095 ( n12179 , new_n21510 , new_n21529 );
xnor g20096 ( n12192 , new_n6370 , new_n6417 );
xnor g20097 ( n12223 , new_n21842 , new_n21851 );
xnor g20098 ( n12225 , new_n10112 , new_n10157 );
xnor g20099 ( n12228 , new_n21905_1 , new_n21914 );
xnor g20100 ( n12235 , new_n7199 , new_n13129 );
xnor g20101 ( n12302 , new_n9021 , new_n9047_1 );
xnor g20102 ( n12304 , new_n16331 , new_n16359 );
xnor g20103 ( new_n22452 , n1742 , n19196 );
nor  g20104 ( new_n22453 , n4858 , new_n11812 );
xnor g20105 ( new_n22454 , n4858 , n23586 );
nor  g20106 ( new_n22455 , n8244 , new_n15238 );
xnor g20107 ( new_n22456 , n8244 , n21226 );
nor  g20108 ( new_n22457 , new_n6170 , n9493 );
nor  g20109 ( new_n22458 , new_n12132 , n20036 );
and  g20110 ( new_n22459 , new_n19090 , new_n19095 );
nor  g20111 ( new_n22460 , new_n22458 , new_n22459 );
xnor g20112 ( new_n22461 , n4426 , n9493 );
and  g20113 ( new_n22462 , new_n22460 , new_n22461 );
or   g20114 ( new_n22463 , new_n22457 , new_n22462 );
and  g20115 ( new_n22464 , new_n22456 , new_n22463 );
or   g20116 ( new_n22465 , new_n22455 , new_n22464 );
and  g20117 ( new_n22466 , new_n22454 , new_n22465 );
or   g20118 ( new_n22467_1 , new_n22453 , new_n22466 );
xor  g20119 ( new_n22468 , new_n22452 , new_n22467_1 );
xnor g20120 ( new_n22469 , new_n19050 , new_n22468 );
xor  g20121 ( new_n22470_1 , new_n22454 , new_n22465 );
nor  g20122 ( new_n22471 , new_n17704 , new_n22470_1 );
xnor g20123 ( new_n22472 , new_n17704 , new_n22470_1 );
xor  g20124 ( new_n22473 , new_n22456 , new_n22463 );
nor  g20125 ( new_n22474 , new_n17706 , new_n22473 );
xnor g20126 ( new_n22475 , new_n17706 , new_n22473 );
xnor g20127 ( new_n22476 , new_n22460 , new_n22461 );
and  g20128 ( new_n22477 , new_n17711 , new_n22476 );
xnor g20129 ( new_n22478 , new_n17711 , new_n22476 );
and  g20130 ( new_n22479 , new_n17713 , new_n19096 );
nor  g20131 ( new_n22480 , new_n19097 , new_n19105 );
nor  g20132 ( new_n22481 , new_n22479 , new_n22480 );
nor  g20133 ( new_n22482 , new_n22478 , new_n22481 );
nor  g20134 ( new_n22483 , new_n22477 , new_n22482 );
nor  g20135 ( new_n22484_1 , new_n22475 , new_n22483 );
nor  g20136 ( new_n22485 , new_n22474 , new_n22484_1 );
nor  g20137 ( new_n22486 , new_n22472 , new_n22485 );
nor  g20138 ( new_n22487 , new_n22471 , new_n22486 );
xnor g20139 ( n12324 , new_n22469 , new_n22487 );
xnor g20140 ( n12325 , new_n20827 , new_n20830 );
xor  g20141 ( n12329 , new_n10377 , new_n10393 );
xnor g20142 ( n12330 , new_n8638_1 , new_n8639 );
xnor g20143 ( n12346 , new_n5716 , new_n5759 );
xnor g20144 ( n12349 , new_n7573 , new_n7592 );
xnor g20145 ( n12364 , new_n18845 , new_n18846 );
nor  g20146 ( new_n22495 , new_n5699 , new_n21424 );
xnor g20147 ( new_n22496 , new_n5699 , new_n21425 );
nor  g20148 ( new_n22497 , new_n5702 , new_n21424 );
xnor g20149 ( new_n22498 , new_n5702 , new_n21424 );
nor  g20150 ( new_n22499 , new_n5706 , new_n21347 );
xnor g20151 ( new_n22500 , new_n5706 , new_n21347 );
nor  g20152 ( new_n22501 , new_n5710 , new_n21349_1 );
nor  g20153 ( new_n22502 , new_n22340 , new_n22355 );
nor  g20154 ( new_n22503 , new_n22501 , new_n22502 );
nor  g20155 ( new_n22504 , new_n22500 , new_n22503 );
nor  g20156 ( new_n22505 , new_n22499 , new_n22504 );
nor  g20157 ( new_n22506 , new_n22498 , new_n22505 );
nor  g20158 ( new_n22507 , new_n22497 , new_n22506 );
and  g20159 ( new_n22508 , new_n22496 , new_n22507 );
nor  g20160 ( n12383 , new_n22495 , new_n22508 );
xnor g20161 ( n12397 , new_n8557 , new_n8558 );
xor  g20162 ( n12408 , new_n16706 , new_n16718 );
nor  g20163 ( new_n22512 , new_n15180_1 , new_n19155 );
and  g20164 ( new_n22513 , new_n22395 , new_n22398 );
nor  g20165 ( n12449 , new_n22512 , new_n22513 );
xnor g20166 ( n12461 , new_n20587 , new_n20619 );
not  g20167 ( new_n22516 , new_n16797 );
nor  g20168 ( new_n22517 , new_n11846 , new_n20458 );
nor  g20169 ( new_n22518 , new_n22516 , new_n22517 );
and  g20170 ( new_n22519 , new_n22516 , new_n22517 );
nor  g20171 ( new_n22520 , new_n16853 , new_n20459 );
nor  g20172 ( new_n22521 , new_n20460 , new_n20468 );
nor  g20173 ( new_n22522 , new_n22520 , new_n22521 );
nor  g20174 ( new_n22523 , new_n22519 , new_n22522 );
or   g20175 ( n12462 , new_n22518 , new_n22523 );
xor  g20176 ( n12467 , new_n21535 , new_n21541 );
nor  g20177 ( new_n22526 , n3324 , new_n15563 );
or   g20178 ( new_n22527 , new_n15568 , new_n15595 );
and  g20179 ( new_n22528 , new_n15565 , new_n22527 );
nor  g20180 ( new_n22529 , new_n22526 , new_n22528 );
not  g20181 ( new_n22530 , new_n22529 );
nor  g20182 ( new_n22531 , new_n21214 , new_n22530 );
nor  g20183 ( new_n22532 , new_n15665 , new_n15672 );
nor  g20184 ( new_n22533_1 , n13419 , new_n15671 );
nor  g20185 ( new_n22534 , new_n22532 , new_n22533_1 );
not  g20186 ( new_n22535 , new_n22534 );
nor  g20187 ( new_n22536 , new_n21944 , new_n22535 );
xnor g20188 ( new_n22537 , new_n21214 , new_n22529 );
xnor g20189 ( new_n22538 , new_n21943_1 , new_n22535 );
nor  g20190 ( new_n22539 , new_n22537 , new_n22538 );
xnor g20191 ( new_n22540 , new_n22537 , new_n22538 );
not  g20192 ( new_n22541 , new_n22540 );
nor  g20193 ( new_n22542 , new_n15597 , new_n15673 );
and  g20194 ( new_n22543 , new_n15674 , new_n15715 );
nor  g20195 ( new_n22544 , new_n22542 , new_n22543 );
and  g20196 ( new_n22545 , new_n22541 , new_n22544 );
nor  g20197 ( new_n22546 , new_n22539 , new_n22545 );
xor  g20198 ( new_n22547 , new_n22536 , new_n22546 );
xnor g20199 ( n12469 , new_n22531 , new_n22547 );
xnor g20200 ( n12515 , new_n10842 , new_n10866 );
nor  g20201 ( new_n22550 , n5140 , new_n11795 );
xnor g20202 ( new_n22551 , n5140 , n10250 );
nor  g20203 ( new_n22552 , n6204 , new_n6155 );
xnor g20204 ( new_n22553 , n6204 , n7674 );
nor  g20205 ( new_n22554_1 , n3349 , new_n6158 );
xnor g20206 ( new_n22555 , n3349 , n6397 );
nor  g20207 ( new_n22556 , n1742 , new_n6161 );
and  g20208 ( new_n22557 , new_n22452 , new_n22467_1 );
or   g20209 ( new_n22558 , new_n22556 , new_n22557 );
and  g20210 ( new_n22559 , new_n22555 , new_n22558 );
or   g20211 ( new_n22560 , new_n22554_1 , new_n22559 );
and  g20212 ( new_n22561 , new_n22553 , new_n22560 );
or   g20213 ( new_n22562 , new_n22552 , new_n22561 );
and  g20214 ( new_n22563 , new_n22551 , new_n22562 );
nor  g20215 ( new_n22564 , new_n22550 , new_n22563 );
xnor g20216 ( new_n22565 , new_n21291 , new_n22564 );
and  g20217 ( new_n22566 , new_n20203 , new_n22564 );
or   g20218 ( new_n22567 , new_n20203 , new_n22564 );
xor  g20219 ( new_n22568 , new_n22551 , new_n22562 );
nor  g20220 ( new_n22569 , new_n20205 , new_n22568 );
xnor g20221 ( new_n22570 , new_n20205 , new_n22568 );
xor  g20222 ( new_n22571 , new_n22553 , new_n22560 );
nor  g20223 ( new_n22572 , new_n19045 , new_n22571 );
xnor g20224 ( new_n22573 , new_n19045 , new_n22571 );
xor  g20225 ( new_n22574 , new_n22555 , new_n22558 );
nor  g20226 ( new_n22575 , new_n19047 , new_n22574 );
xnor g20227 ( new_n22576 , new_n19047 , new_n22574 );
nor  g20228 ( new_n22577 , new_n19050 , new_n22468 );
nor  g20229 ( new_n22578 , new_n22469 , new_n22487 );
nor  g20230 ( new_n22579 , new_n22577 , new_n22578 );
nor  g20231 ( new_n22580 , new_n22576 , new_n22579 );
nor  g20232 ( new_n22581 , new_n22575 , new_n22580 );
nor  g20233 ( new_n22582 , new_n22573 , new_n22581 );
nor  g20234 ( new_n22583 , new_n22572 , new_n22582 );
nor  g20235 ( new_n22584_1 , new_n22570 , new_n22583 );
nor  g20236 ( new_n22585 , new_n22569 , new_n22584_1 );
and  g20237 ( new_n22586 , new_n22567 , new_n22585 );
nor  g20238 ( new_n22587 , new_n22566 , new_n22586 );
xnor g20239 ( n12516 , new_n22565 , new_n22587 );
xnor g20240 ( n12540 , new_n7397 , new_n7410 );
xnor g20241 ( n12545 , new_n11564_1 , new_n11565 );
xnor g20242 ( n12552 , new_n19851 , new_n19869 );
xnor g20243 ( n12566 , new_n8167 , new_n8190 );
xnor g20244 ( n12569 , new_n13075 , new_n13091 );
xnor g20245 ( n12607 , new_n6359 , new_n6421 );
xnor g20246 ( n12620 , new_n9916 , new_n9984 );
xnor g20247 ( n12621 , new_n3679_1 , new_n3717 );
xnor g20248 ( n12654 , new_n17895 , new_n17896 );
xnor g20249 ( n12665 , new_n14745 , new_n19098 );
xnor g20250 ( n12670 , new_n16743_1 , new_n16753 );
xnor g20251 ( n12707 , new_n2522 , new_n7581 );
xnor g20252 ( n12725 , new_n7149_1 , new_n7161 );
xnor g20253 ( n12727 , new_n15680 , new_n15713 );
xor  g20254 ( n12740 , new_n9671 , new_n9695_1 );
xor  g20255 ( n12742 , new_n20172 , new_n20173 );
xnor g20256 ( n12746 , new_n2826_1 , new_n20364 );
xor  g20257 ( n12756 , new_n9204 , new_n9205 );
xnor g20258 ( n12783 , new_n7124 , new_n7174 );
xnor g20259 ( new_n22608 , new_n20203 , new_n22564 );
xnor g20260 ( n12801 , new_n22585 , new_n22608 );
xnor g20261 ( n12812 , new_n17377 , new_n17380 );
xnor g20262 ( n12816 , new_n15888 , new_n15921 );
nor  g20263 ( new_n22612 , n6659 , new_n16936 );
and  g20264 ( new_n22613 , new_n17929 , new_n17949 );
nor  g20265 ( new_n22614 , new_n22612 , new_n22613 );
not  g20266 ( new_n22615 , new_n22614 );
nor  g20267 ( new_n22616 , new_n19325 , new_n22615 );
xnor g20268 ( new_n22617 , new_n19324 , new_n22615 );
nor  g20269 ( new_n22618 , new_n22537 , new_n22617 );
xnor g20270 ( new_n22619_1 , new_n22537 , new_n22617 );
and  g20271 ( new_n22620_1 , new_n15597 , new_n17950 );
nor  g20272 ( new_n22621 , new_n17951 , new_n17974 );
nor  g20273 ( new_n22622 , new_n22620_1 , new_n22621 );
nor  g20274 ( new_n22623_1 , new_n22619_1 , new_n22622 );
nor  g20275 ( new_n22624 , new_n22618 , new_n22623_1 );
nor  g20276 ( new_n22625 , new_n22616 , new_n22624 );
nor  g20277 ( n12843 , new_n22531 , new_n22625 );
xnor g20278 ( n12864 , new_n20407 , new_n20409_1 );
nor  g20279 ( new_n22628 , new_n4839 , new_n21655 );
and  g20280 ( new_n22629 , new_n21656 , new_n21681 );
nor  g20281 ( new_n22630 , new_n22628 , new_n22629 );
nor  g20282 ( new_n22631_1 , n3740 , n21784 );
and  g20283 ( new_n22632 , new_n21635 , new_n21654_1 );
nor  g20284 ( new_n22633 , new_n22631_1 , new_n22632 );
xnor g20285 ( new_n22634 , new_n4901 , new_n22633 );
xnor g20286 ( new_n22635 , new_n22630 , new_n22634 );
not  g20287 ( new_n22636 , new_n22635 );
nor  g20288 ( new_n22637 , new_n18323_1 , new_n22636 );
nor  g20289 ( new_n22638 , new_n17136 , new_n21682 );
and  g20290 ( new_n22639 , new_n21683 , new_n21706 );
or   g20291 ( new_n22640 , new_n22638 , new_n22639 );
xnor g20292 ( new_n22641 , new_n18322 , new_n22636 );
and  g20293 ( new_n22642 , new_n22640 , new_n22641 );
nor  g20294 ( new_n22643 , new_n22637 , new_n22642 );
and  g20295 ( new_n22644 , new_n13919 , new_n22633 );
nor  g20296 ( new_n22645 , new_n13919 , new_n22633 );
nor  g20297 ( new_n22646 , new_n22630 , new_n22645 );
nor  g20298 ( new_n22647 , new_n22644 , new_n22646 );
and  g20299 ( n12865 , new_n22643 , new_n22647 );
xnor g20300 ( n12870 , new_n12707_1 , new_n12724 );
xnor g20301 ( n12873 , new_n20354 , new_n20372 );
not  g20302 ( new_n22651 , new_n21810 );
nor  g20303 ( new_n22652 , new_n18143_1 , new_n22651 );
xnor g20304 ( new_n22653 , new_n18144 , new_n21810 );
nor  g20305 ( new_n22654 , new_n18226 , new_n21186 );
nor  g20306 ( new_n22655 , new_n22132 , new_n22135 );
nor  g20307 ( new_n22656 , new_n22654 , new_n22655 );
nor  g20308 ( new_n22657 , new_n22653 , new_n22656 );
or   g20309 ( n12904 , new_n22652 , new_n22657 );
xor  g20310 ( n12941 , new_n10397 , new_n10398 );
xnor g20311 ( n12942 , new_n11129 , new_n11137 );
xnor g20312 ( new_n22661 , new_n5846 , new_n5844 );
xnor g20313 ( n12978 , new_n5849 , new_n22661 );
xnor g20314 ( n12980 , new_n7887 , new_n9709 );
not  g20315 ( new_n22664 , new_n6568 );
xnor g20316 ( n12985 , new_n4711 , new_n22664 );
xnor g20317 ( n12987 , new_n14257 , new_n14289 );
nor  g20318 ( new_n22667 , new_n12808 , n11220 );
and  g20319 ( new_n22668 , new_n16416 , new_n16431 );
nor  g20320 ( new_n22669 , new_n22667 , new_n22668 );
xnor g20321 ( new_n22670 , new_n14546_1 , new_n22669 );
and  g20322 ( new_n22671 , new_n14589 , new_n16432 );
and  g20323 ( new_n22672 , new_n16433_1 , new_n16452 );
nor  g20324 ( new_n22673 , new_n22671 , new_n22672 );
xnor g20325 ( n12992 , new_n22670 , new_n22673 );
nor  g20326 ( new_n22675 , n6659 , new_n21474 );
nor  g20327 ( new_n22676 , n23250 , new_n20546 );
and  g20328 ( new_n22677 , new_n20548 , new_n20582_1 );
nor  g20329 ( new_n22678 , new_n22676 , new_n22677 );
nor  g20330 ( new_n22679 , new_n21940 , new_n21475 );
nor  g20331 ( new_n22680 , new_n22678 , new_n22679 );
nor  g20332 ( new_n22681 , new_n22675 , new_n22680 );
nor  g20333 ( new_n22682 , new_n21473 , new_n22681 );
not  g20334 ( new_n22683 , new_n22682 );
xnor g20335 ( new_n22684 , new_n19336 , new_n22683 );
xnor g20336 ( new_n22685 , n6659 , new_n21475 );
xnor g20337 ( new_n22686 , new_n22678 , new_n22685 );
nor  g20338 ( new_n22687 , new_n19349 , new_n22686 );
nor  g20339 ( new_n22688 , new_n14075 , new_n20583 );
and  g20340 ( new_n22689 , new_n20584 , new_n20621 );
or   g20341 ( new_n22690 , new_n22688 , new_n22689 );
xnor g20342 ( new_n22691 , new_n19350 , new_n22686 );
and  g20343 ( new_n22692 , new_n22690 , new_n22691 );
nor  g20344 ( new_n22693 , new_n22687 , new_n22692 );
xnor g20345 ( n13005 , new_n22684 , new_n22693 );
xnor g20346 ( n13043 , new_n16307 , new_n19438 );
xnor g20347 ( n13048 , new_n17454 , new_n17455 );
xnor g20348 ( n13054 , new_n15112 , new_n15113 );
xnor g20349 ( n13082 , new_n17603 , new_n17615 );
xnor g20350 ( n13096 , new_n7140 , new_n7166 );
xnor g20351 ( n13116 , new_n17598 , new_n17617 );
xnor g20352 ( n13122 , new_n19420 , new_n19453 );
xnor g20353 ( n13141 , new_n6402 , new_n6403 );
xor  g20354 ( n13144 , new_n19282_1 , new_n19289 );
xnor g20355 ( n13168 , new_n19841 , new_n19875 );
xnor g20356 ( n13198 , new_n20510 , new_n20528 );
xnor g20357 ( n13199 , new_n14266 , new_n14283 );
xnor g20358 ( n13204 , new_n14385 , new_n14397 );
xnor g20359 ( n13209 , new_n10123 , new_n10150 );
xnor g20360 ( n13270 , new_n19077 , new_n19086 );
xnor g20361 ( n13273 , new_n12962 , new_n12983 );
xnor g20362 ( n13285 , new_n21506 , new_n21531 );
xnor g20363 ( n13338 , new_n20909 , new_n20927 );
xnor g20364 ( n13407 , new_n7873 , new_n7904 );
xnor g20365 ( new_n22714_1 , new_n4264 , new_n5432 );
xnor g20366 ( n13409 , new_n15955 , new_n22714_1 );
xnor g20367 ( n13456 , new_n5416 , new_n5445 );
nor  g20368 ( new_n22717 , new_n20221 , new_n20872 );
nor  g20369 ( new_n22718 , new_n20225 , new_n20903 );
nor  g20370 ( new_n22719 , new_n21883 , new_n21886 );
nor  g20371 ( new_n22720 , new_n22718 , new_n22719 );
or   g20372 ( new_n22721 , new_n20221 , new_n20793 );
and  g20373 ( new_n22722 , new_n22720 , new_n22721 );
and  g20374 ( new_n22723 , new_n22717 , new_n22722 );
xnor g20375 ( new_n22724 , new_n20332 , new_n20794_1 );
xnor g20376 ( new_n22725 , new_n22720 , new_n22724 );
and  g20377 ( new_n22726 , new_n11288 , new_n22725 );
xnor g20378 ( new_n22727 , new_n11288 , new_n22725 );
nor  g20379 ( new_n22728 , new_n11380 , new_n21887 );
nor  g20380 ( new_n22729 , new_n21888 , new_n21891 );
or   g20381 ( new_n22730 , new_n22728 , new_n22729 );
nor  g20382 ( new_n22731 , new_n22727 , new_n22730 );
nor  g20383 ( new_n22732 , new_n22726 , new_n22731 );
xnor g20384 ( new_n22733 , new_n20221 , new_n20873 );
and  g20385 ( new_n22734 , new_n22720 , new_n22733 );
nor  g20386 ( new_n22735 , new_n22722 , new_n22733 );
nor  g20387 ( new_n22736 , new_n22734 , new_n22735 );
nor  g20388 ( new_n22737 , new_n22732 , new_n22736 );
or   g20389 ( n13457 , new_n22723 , new_n22737 );
xnor g20390 ( n13477 , new_n12031 , new_n12039 );
xnor g20391 ( n13484 , new_n12348 , new_n12349_1 );
xnor g20392 ( n13486 , new_n20031 , new_n20059 );
xnor g20393 ( new_n22742 , new_n20957 , new_n21437 );
and  g20394 ( new_n22743 , new_n17024 , new_n21357 );
nor  g20395 ( new_n22744 , new_n21358 , new_n21382 );
nor  g20396 ( new_n22745 , new_n22743 , new_n22744 );
xor  g20397 ( n13487 , new_n22742 , new_n22745 );
xnor g20398 ( n13500 , new_n5194 , new_n5213_1 );
xor  g20399 ( n13501 , new_n4590_1 , new_n4592 );
xnor g20400 ( n13506 , new_n6388 , new_n6409 );
xnor g20401 ( n13548 , new_n6124 , new_n6135 );
xnor g20402 ( n13551 , new_n22305 , new_n22325 );
xnor g20403 ( n13602 , new_n4995 , new_n5014 );
xnor g20404 ( n13626 , new_n17111 , new_n17120 );
xnor g20405 ( n13683 , new_n8177 , new_n8186 );
xnor g20406 ( n13710 , new_n19620 , new_n19657 );
xnor g20407 ( n13722 , new_n19276 , new_n19293 );
xnor g20408 ( new_n22757 , new_n13870 , new_n13925 );
xnor g20409 ( n13754 , new_n13992 , new_n22757 );
xor  g20410 ( n13764 , new_n2805 , new_n2839 );
xnor g20411 ( new_n22760 , new_n14139 , new_n14142 );
xnor g20412 ( n13798 , new_n14147_1 , new_n22760 );
xnor g20413 ( n13835 , new_n17106_1 , new_n17124 );
xnor g20414 ( n13850 , new_n15535 , new_n15537 );
xnor g20415 ( n13922 , new_n7888 , new_n17605 );
xnor g20416 ( n13923 , new_n19049 , new_n19057 );
xnor g20417 ( n14004 , new_n11569 , new_n11570 );
xnor g20418 ( n14036 , new_n11748 , new_n11787 );
xnor g20419 ( n14059 , new_n20991 , new_n21005 );
xor  g20420 ( n14081 , new_n16922 , new_n16925 );
xnor g20421 ( n14095 , new_n18540 , new_n18543 );
xnor g20422 ( n14107 , new_n11603 , new_n6728 );
xnor g20423 ( n14121 , new_n8870 , new_n8901 );
xnor g20424 ( n14126 , new_n12000_1 , new_n12002 );
xnor g20425 ( n14136 , new_n19270_1 , new_n19297 );
not  g20426 ( new_n22775 , new_n22669 );
nor  g20427 ( new_n22776 , new_n14546_1 , new_n22775 );
nor  g20428 ( new_n22777 , new_n14545 , new_n22669 );
nor  g20429 ( new_n22778 , new_n22777 , new_n22673 );
nor  g20430 ( new_n22779_1 , new_n22776 , new_n22778 );
xnor g20431 ( new_n22780 , new_n21723 , new_n22775 );
xnor g20432 ( n14147 , new_n22779_1 , new_n22780 );
xnor g20433 ( n14174 , new_n20700_1 , new_n20738 );
xnor g20434 ( n14190 , new_n16197 , new_n16221 );
xnor g20435 ( n14211 , new_n5420 , new_n5443_1 );
xnor g20436 ( n14222 , new_n16404 , new_n16407_1 );
xnor g20437 ( n14267 , new_n13262 , new_n13306 );
xnor g20438 ( n14271 , new_n5738 , new_n5749 );
xnor g20439 ( n14277 , new_n9372_1 , new_n9383 );
xnor g20440 ( n14294 , new_n8372 , new_n8373 );
xnor g20441 ( n14310 , new_n22296 , new_n22331 );
xnor g20442 ( n14326 , new_n22346 , new_n22349 );
xnor g20443 ( n14342 , new_n12262 , new_n12306 );
xnor g20444 ( n14353 , new_n18063 , new_n18073 );
and  g20445 ( new_n22794 , new_n11593 , new_n20987 );
nor  g20446 ( new_n22795 , new_n8953 , new_n20987 );
nor  g20447 ( new_n22796 , new_n20988 , new_n21007 );
nor  g20448 ( new_n22797 , new_n22795 , new_n22796 );
nor  g20449 ( new_n22798 , new_n22794 , new_n22797 );
nor  g20450 ( new_n22799 , new_n11593 , new_n20987 );
nor  g20451 ( new_n22800 , new_n22796 , new_n22799 );
nor  g20452 ( n14364 , new_n22798 , new_n22800 );
xor  g20453 ( n14375 , new_n21442 , new_n21445 );
xnor g20454 ( n14412 , new_n21834 , new_n21859 );
or   g20455 ( new_n22804 , new_n6240 , new_n17339 );
nor  g20456 ( new_n22805 , new_n22804 , new_n17363 );
xnor g20457 ( new_n22806 , new_n11524 , new_n22805 );
and  g20458 ( new_n22807 , new_n17331 , new_n17364 );
nor  g20459 ( new_n22808 , new_n17365 , new_n17388 );
nor  g20460 ( new_n22809 , new_n22807 , new_n22808 );
not  g20461 ( new_n22810 , new_n22809 );
xnor g20462 ( n14414 , new_n22806 , new_n22810 );
xnor g20463 ( n14457 , new_n15308 , new_n15310 );
xnor g20464 ( n14464 , new_n4987 , new_n5018 );
xnor g20465 ( n14471 , new_n10846 , new_n10864 );
nor  g20466 ( new_n22815 , new_n8339_1 , new_n19324 );
nor  g20467 ( new_n22816 , new_n19326 , new_n19334 );
nor  g20468 ( new_n22817 , new_n22815 , new_n22816 );
not  g20469 ( new_n22818 , new_n22817 );
xnor g20470 ( new_n22819_1 , new_n22682 , new_n22818 );
nor  g20471 ( new_n22820 , new_n19335 , new_n22683 );
nor  g20472 ( new_n22821 , new_n19336 , new_n22682 );
nor  g20473 ( new_n22822 , new_n22821 , new_n22693 );
nor  g20474 ( new_n22823 , new_n22820 , new_n22822 );
xnor g20475 ( n14475 , new_n22819_1 , new_n22823 );
xnor g20476 ( n14541 , new_n12293 , new_n12294 );
nor  g20477 ( new_n22826 , new_n21227 , new_n21231 );
nor  g20478 ( new_n22827 , new_n21232 , new_n21241 );
or   g20479 ( n14546 , new_n22826 , new_n22827 );
xnor g20480 ( n14547 , new_n11064 , new_n11065 );
xnor g20481 ( n14593 , new_n12632 , new_n12651 );
xnor g20482 ( n14636 , new_n9362 , new_n9387 );
xnor g20483 ( n14701 , new_n22472 , new_n22485 );
xnor g20484 ( n14734 , new_n12080 , new_n12089 );
xnor g20485 ( n14746 , new_n7128 , new_n7172 );
xnor g20486 ( n14763 , new_n9685 , new_n9687 );
xnor g20487 ( n14772 , new_n22048 , new_n22056 );
xnor g20488 ( n14801 , new_n21447 , new_n21448 );
xnor g20489 ( n14819 , new_n21031 , new_n21050 );
xnor g20490 ( n14827 , new_n14373 , new_n14405 );
xnor g20491 ( n14839 , new_n20463 , new_n20466 );
xnor g20492 ( n14849 , new_n17115 , new_n17116 );
nor  g20493 ( new_n22842 , new_n14356 , new_n20330_1 );
nor  g20494 ( new_n22843_1 , new_n20331 , new_n20387 );
nor  g20495 ( new_n22844 , new_n22842 , new_n22843_1 );
nor  g20496 ( n14891 , new_n20327 , new_n22844 );
xnor g20497 ( n14931 , new_n15341 , new_n6532 );
and  g20498 ( new_n22847 , new_n11524 , new_n22805 );
and  g20499 ( new_n22848 , new_n22847 , new_n22810 );
or   g20500 ( new_n22849 , new_n11524 , new_n22805 );
nor  g20501 ( new_n22850 , new_n22849 , new_n22810 );
or   g20502 ( n14944 , new_n22848 , new_n22850 );
xnor g20503 ( n14977 , new_n8911_1 , new_n18069 );
xnor g20504 ( n14989 , new_n12614 , new_n12659 );
xnor g20505 ( n15002 , new_n10752 , new_n10760 );
xnor g20506 ( n15004 , new_n5746 , new_n21910 );
xnor g20507 ( n15011 , new_n9013 , new_n9051 );
xor  g20508 ( n15019 , new_n21962 , new_n21965 );
nor  g20509 ( new_n22858_1 , new_n15090 , new_n15098 );
nor  g20510 ( new_n22859 , new_n15099 , new_n15119 );
or   g20511 ( n15031 , new_n22858_1 , new_n22859 );
xnor g20512 ( n15033 , new_n17604 , new_n17606 );
xnor g20513 ( n15052 , new_n7200 , new_n11884 );
xnor g20514 ( n15082 , new_n19201 , new_n19210 );
xnor g20515 ( n15094 , new_n8171 , new_n8188 );
xor  g20516 ( n15118 , new_n11621 , new_n11624 );
xnor g20517 ( n15128 , new_n22653 , new_n22656 );
xnor g20518 ( n15139 , new_n18405_1 , new_n18444_1 );
xnor g20519 ( new_n22868 , new_n16495 , new_n16500 );
xnor g20520 ( n15145 , new_n16510 , new_n22868 );
xnor g20521 ( n15165 , new_n14594 , new_n14624 );
xnor g20522 ( n15176 , new_n5081 , new_n15032 );
xor  g20523 ( n15180 , new_n19862 , new_n19863 );
xnor g20524 ( n15205 , new_n15939 , new_n15973 );
not  g20525 ( new_n22874 , new_n5436 );
xnor g20526 ( n15230 , new_n4266_1 , new_n22874 );
xor  g20527 ( n15255 , new_n16748 , new_n16749 );
xnor g20528 ( n15275 , new_n9661 , new_n9699_1 );
xnor g20529 ( n15300 , new_n13763 , new_n13766 );
or   g20530 ( new_n22879_1 , new_n13194 , new_n22420 );
nor  g20531 ( new_n22880 , new_n22419 , new_n22879_1 );
and  g20532 ( new_n22881 , new_n13194 , new_n22420 );
and  g20533 ( new_n22882 , new_n22419 , new_n22881 );
nor  g20534 ( new_n22883 , new_n22880 , new_n22882 );
xnor g20535 ( new_n22884 , new_n21227 , new_n22883 );
nor  g20536 ( new_n22885 , new_n21190 , new_n22422 );
nor  g20537 ( new_n22886 , new_n22423 , new_n22431 );
nor  g20538 ( new_n22887 , new_n22885 , new_n22886 );
not  g20539 ( new_n22888 , new_n22887 );
xnor g20540 ( n15307 , new_n22884 , new_n22888 );
xnor g20541 ( n15327 , new_n19617_1 , new_n19659 );
xnor g20542 ( n15345 , new_n19638 , new_n19645 );
xnor g20543 ( n15353 , new_n12638 , new_n12649 );
xor  g20544 ( n15366 , new_n22496 , new_n22507 );
xnor g20545 ( n15382 , new_n22643 , new_n22647 );
xnor g20546 ( n15407 , new_n9194 , new_n9211 );
not  g20547 ( new_n22896 , new_n13377 );
xnor g20548 ( n15428 , new_n22896 , new_n14962 );
and  g20549 ( new_n22898 , new_n22271 , new_n22274_1 );
and  g20550 ( new_n22899 , new_n22275 , new_n22290_1 );
nor  g20551 ( new_n22900 , new_n22291 , new_n22333 );
nor  g20552 ( new_n22901 , new_n22899 , new_n22900 );
nor  g20553 ( new_n22902 , new_n22898 , new_n22901 );
or   g20554 ( new_n22903_1 , new_n11025_1 , new_n22279 );
nor  g20555 ( new_n22904 , new_n22903_1 , new_n22288 );
not  g20556 ( new_n22905 , new_n22904 );
nor  g20557 ( new_n22906 , new_n22898 , new_n22905 );
nor  g20558 ( new_n22907_1 , new_n22900 , new_n22906 );
nor  g20559 ( n15435 , new_n22902 , new_n22907_1 );
or   g20560 ( new_n22909 , new_n21919 , new_n21924 );
nor  g20561 ( new_n22910_1 , new_n22909 , new_n21934_1 );
and  g20562 ( new_n22911 , new_n21919 , new_n21924 );
and  g20563 ( new_n22912 , new_n22911 , new_n21934_1 );
or   g20564 ( n15438 , new_n22910_1 , new_n22912 );
xnor g20565 ( n15465 , new_n22302 , new_n22327 );
xnor g20566 ( n15467 , new_n6665 , new_n8556 );
xnor g20567 ( n15470 , new_n7843 , new_n7914 );
xnor g20568 ( n15477 , new_n14366 , new_n14409 );
xnor g20569 ( n15481 , new_n22573 , new_n22581 );
xnor g20570 ( n15496 , new_n14833 , new_n14836 );
xnor g20571 ( n15501 , new_n11983 , new_n12012 );
xnor g20572 ( n15555 , new_n18537_1 , new_n18545 );
xnor g20573 ( n15558 , new_n20852 , new_n20867 );
nor  g20574 ( new_n22923 , new_n22651 , new_n21226_1 );
nor  g20575 ( new_n22924 , new_n21811 , new_n21814 );
or   g20576 ( n15559 , new_n22923 , new_n22924 );
and  g20577 ( new_n22926 , n5101 , new_n5453 );
and  g20578 ( new_n22927 , new_n19882 , new_n19897 );
nor  g20579 ( new_n22928 , new_n22926 , new_n22927 );
not  g20580 ( new_n22929 , new_n22928 );
nor  g20581 ( new_n22930 , new_n22007 , new_n22929 );
and  g20582 ( new_n22931 , new_n19898 , new_n20501 );
and  g20583 ( new_n22932 , new_n19948 , new_n19972 );
nor  g20584 ( new_n22933 , new_n22931 , new_n22932 );
nor  g20585 ( new_n22934 , new_n21219 , new_n22928 );
nor  g20586 ( new_n22935 , new_n22933 , new_n22934 );
and  g20587 ( new_n22936 , new_n22007 , new_n22935 );
nor  g20588 ( new_n22937 , new_n21219 , new_n22929 );
nor  g20589 ( new_n22938 , new_n22935 , new_n22937 );
or   g20590 ( new_n22939_1 , new_n22936 , new_n22938 );
nor  g20591 ( n15570 , new_n22930 , new_n22939_1 );
xnor g20592 ( n15573 , new_n12250 , new_n12312 );
xnor g20593 ( n15588 , new_n11580_1 , new_n11581 );
xnor g20594 ( n15590 , new_n21038 , new_n21046_1 );
xnor g20595 ( n15598 , new_n21594 , new_n21604 );
xnor g20596 ( n15614 , new_n9357 , new_n9389 );
xnor g20597 ( n15662 , new_n22042 , new_n22060 );
xnor g20598 ( n15716 , new_n3352 , new_n3383 );
xnor g20599 ( n15749 , new_n14254 , new_n14291 );
xnor g20600 ( n15762 , new_n18460 , new_n18463 );
xnor g20601 ( n15793 , new_n7887 , new_n7889 );
xnor g20602 ( n15812 , new_n21840 , new_n21853 );
xnor g20603 ( n15815 , new_n12258 , new_n12308 );
xnor g20604 ( n15816 , new_n8369 , new_n8370 );
xnor g20605 ( n15831 , new_n11878 , new_n11890 );
xnor g20606 ( n15846 , new_n9559 , new_n9561 );
xnor g20607 ( n15859 , new_n8427 , new_n8428 );
nor  g20608 ( new_n22957 , new_n21421 , new_n8079 );
and  g20609 ( new_n22958 , new_n19524 , new_n19539_1 );
nor  g20610 ( new_n22959 , new_n22957 , new_n22958 );
nor  g20611 ( new_n22960 , new_n8075 , new_n22959 );
xnor g20612 ( new_n22961 , new_n21276_1 , new_n22960 );
xnor g20613 ( new_n22962 , new_n8074 , new_n22959 );
nor  g20614 ( new_n22963 , new_n19833 , new_n22962 );
nor  g20615 ( new_n22964 , new_n19523_1 , new_n19540 );
nor  g20616 ( new_n22965 , new_n19541 , new_n19562 );
nor  g20617 ( new_n22966 , new_n22964 , new_n22965 );
xnor g20618 ( new_n22967 , new_n19833 , new_n22962 );
nor  g20619 ( new_n22968 , new_n22966 , new_n22967 );
nor  g20620 ( new_n22969 , new_n22963 , new_n22968 );
xnor g20621 ( n15869 , new_n22961 , new_n22969 );
xnor g20622 ( n15885 , new_n18563 , new_n18588 );
not  g20623 ( new_n22972 , new_n20696_1 );
and  g20624 ( new_n22973 , new_n15335 , new_n22972 );
and  g20625 ( new_n22974 , new_n22973 , new_n20740 );
and  g20626 ( new_n22975 , new_n20696_1 , new_n20739 );
or   g20627 ( n15889 , new_n22974 , new_n22975 );
xnor g20628 ( n15917 , new_n13634 , new_n18575 );
xnor g20629 ( n15922 , new_n13627 , new_n13628 );
not  g20630 ( new_n22979 , new_n7150 );
xnor g20631 ( n15947 , new_n22979 , new_n7151 );
and  g20632 ( new_n22981 , new_n7241 , new_n19135 );
and  g20633 ( new_n22982 , new_n20392 , new_n20399 );
nor  g20634 ( new_n22983 , new_n22981 , new_n22982 );
not  g20635 ( new_n22984 , new_n22983 );
xnor g20636 ( new_n22985 , new_n19163_1 , new_n22984 );
nor  g20637 ( new_n22986 , new_n19162 , new_n20400 );
nor  g20638 ( new_n22987 , new_n20402_1 , new_n20411_1 );
nor  g20639 ( new_n22988 , new_n22986 , new_n22987 );
xor  g20640 ( n15956 , new_n22985 , new_n22988 );
xor  g20641 ( n15958 , new_n13395 , new_n13398 );
nor  g20642 ( new_n22991 , new_n12059 , new_n16781 );
and  g20643 ( new_n22992 , new_n12063 , new_n16781 );
nor  g20644 ( new_n22993 , new_n22991 , new_n22992 );
nor  g20645 ( new_n22994 , new_n12059 , new_n16776 );
or   g20646 ( new_n22995 , new_n22994 , new_n16778 );
nor  g20647 ( n15986 , new_n22993 , new_n22995 );
xnor g20648 ( n16013 , new_n22426 , new_n22429 );
nor  g20649 ( new_n22998_1 , new_n20400 , new_n21401 );
nor  g20650 ( new_n22999 , new_n20401 , new_n21402 );
nor  g20651 ( new_n23000 , new_n22999 , new_n21411 );
nor  g20652 ( new_n23001 , new_n22998_1 , new_n23000 );
xnor g20653 ( new_n23002 , new_n21401 , new_n22984 );
xnor g20654 ( n16060 , new_n23001 , new_n23002 );
nor  g20655 ( new_n23004 , new_n11842_1 , new_n16152 );
xnor g20656 ( new_n23005 , n25972 , new_n16152 );
nor  g20657 ( new_n23006_1 , new_n8646 , new_n16154 );
and  g20658 ( new_n23007_1 , new_n22067 , new_n22078 );
or   g20659 ( new_n23008 , new_n23006_1 , new_n23007_1 );
and  g20660 ( new_n23009_1 , new_n23005 , new_n23008 );
nor  g20661 ( new_n23010 , new_n23004 , new_n23009_1 );
nor  g20662 ( new_n23011 , new_n22189 , new_n23010 );
xnor g20663 ( new_n23012 , new_n22189 , new_n23010 );
and  g20664 ( new_n23013 , new_n22290_1 , new_n23012 );
xnor g20665 ( new_n23014_1 , new_n22290_1 , new_n23012 );
not  g20666 ( new_n23015 , new_n22294 );
xor  g20667 ( new_n23016 , new_n23005 , new_n23008 );
nor  g20668 ( new_n23017 , new_n23015 , new_n23016 );
xnor g20669 ( new_n23018 , new_n23015 , new_n23016 );
nor  g20670 ( new_n23019 , new_n22079 , new_n22101 );
nor  g20671 ( new_n23020 , new_n22102 , new_n22117 );
nor  g20672 ( new_n23021 , new_n23019 , new_n23020 );
nor  g20673 ( new_n23022 , new_n23018 , new_n23021 );
nor  g20674 ( new_n23023 , new_n23017 , new_n23022 );
nor  g20675 ( new_n23024 , new_n23014_1 , new_n23023 );
nor  g20676 ( new_n23025 , new_n23013 , new_n23024 );
xnor g20677 ( new_n23026 , new_n23011 , new_n23025 );
xnor g20678 ( n16062 , new_n22905 , new_n23026 );
xnor g20679 ( n16068 , new_n22498 , new_n22505 );
xnor g20680 ( n16080 , new_n22727 , new_n22730 );
and  g20681 ( new_n23030 , new_n6356_1 , new_n22194 );
nor  g20682 ( new_n23031 , new_n22195 , new_n22198_1 );
nor  g20683 ( new_n23032 , new_n23030 , new_n23031 );
nor  g20684 ( new_n23033 , new_n11851 , new_n22189 );
and  g20685 ( new_n23034 , new_n22190 , new_n22193 );
nor  g20686 ( new_n23035_1 , new_n23033 , new_n23034 );
xnor g20687 ( n16098 , new_n23032 , new_n23035_1 );
xnor g20688 ( n16110 , new_n17317 , new_n17325 );
xnor g20689 ( n16142 , new_n14945 , new_n14974 );
xnor g20690 ( n16185 , new_n16341 , new_n16353 );
xnor g20691 ( n16196 , new_n12329_1 , new_n12346_1 );
xnor g20692 ( n16206 , new_n20424_1 , new_n20425 );
xor  g20693 ( n16215 , new_n20494 , new_n20497 );
xnor g20694 ( n16218 , new_n18680 , new_n18688 );
xnor g20695 ( n16219 , new_n3912 , new_n3913 );
xnor g20696 ( n16230 , new_n6949 , new_n6950 );
xor  g20697 ( n16243 , new_n8417_1 , new_n8425 );
xnor g20698 ( n16275 , new_n17059 , new_n17068_1 );
xnor g20699 ( n16279 , new_n10152 , new_n10153 );
nor  g20700 ( new_n23049 , new_n17498 , new_n20014 );
nor  g20701 ( new_n23050 , new_n20015 , new_n20069_1 );
or   g20702 ( n16322 , new_n23049 , new_n23050 );
xnor g20703 ( n16327 , new_n17036 , new_n17076 );
xnor g20704 ( n16350 , new_n20856 , new_n20863 );
xnor g20705 ( n16367 , new_n6665 , new_n6666 );
xnor g20706 ( n16379 , new_n18784 , new_n18785 );
xnor g20707 ( n16398 , new_n19632 , new_n19649 );
xnor g20708 ( n16406 , new_n13383 , new_n13385 );
xnor g20709 ( n16407 , new_n21589 , new_n21606 );
xnor g20710 ( n16419 , new_n23014_1 , new_n23023 );
xnor g20711 ( n16424 , new_n8347 , new_n8387 );
xnor g20712 ( new_n23061 , new_n13673 , new_n13739 );
xnor g20713 ( n16428 , new_n13779 , new_n23061 );
xnor g20714 ( n16433 , new_n11849 , new_n11906 );
xnor g20715 ( n16440 , new_n11857 , new_n11902 );
xnor g20716 ( n16445 , new_n17313 , new_n17327 );
xnor g20717 ( n16460 , new_n13936 , new_n13988 );
xnor g20718 ( n16481 , new_n19549 , new_n19558 );
nor  g20719 ( new_n23068_1 , new_n11021 , new_n14586 );
nor  g20720 ( new_n23069 , new_n11028 , new_n14586 );
nor  g20721 ( new_n23070 , new_n20113 , new_n20129 );
nor  g20722 ( new_n23071 , new_n23069 , new_n23070 );
xor  g20723 ( new_n23072 , new_n11021 , new_n14586 );
and  g20724 ( new_n23073 , new_n23071 , new_n23072 );
nor  g20725 ( n16493 , new_n23068_1 , new_n23073 );
xnor g20726 ( n16506 , new_n4728 , new_n4754 );
xnor g20727 ( n16516 , new_n12715 , new_n12716 );
xor  g20728 ( n16517 , new_n21697 , new_n21698 );
xnor g20729 ( n16527 , new_n15443 , new_n15444 );
xnor g20730 ( n16554 , new_n9156 , new_n10753 );
xnor g20731 ( n16583 , new_n5793 , new_n6130 );
xnor g20732 ( new_n23081 , new_n10028 , new_n21156 );
xnor g20733 ( n16584 , new_n21161 , new_n23081 );
xnor g20734 ( n16589 , new_n18833 , new_n18854 );
xor  g20735 ( n16596 , new_n19180 , new_n19182 );
xnor g20736 ( n16617 , new_n21828 , new_n21865 );
xnor g20737 ( n16630 , new_n7567 , new_n7596 );
xnor g20738 ( n16640 , new_n4940 , new_n21847 );
xnor g20739 ( n16656 , new_n2521 , new_n2522 );
xnor g20740 ( n16674 , new_n6915 , new_n6962 );
xnor g20741 ( n16682 , new_n13940 , new_n13986 );
xnor g20742 ( n16684 , new_n21774 , new_n21793 );
xnor g20743 ( n16688 , new_n10493 , new_n10497 );
xnor g20744 ( n16733 , new_n6397_1 , new_n6405 );
xnor g20745 ( n16798 , new_n7898 , new_n7900 );
xnor g20746 ( n16834 , new_n16447 , new_n16448 );
xnor g20747 ( n16837 , new_n3041 , new_n3080 );
xnor g20748 ( n16841 , new_n21406 , new_n21409 );
xnor g20749 ( n16885 , new_n5085 , new_n5086 );
xnor g20750 ( n16905 , new_n8137 , new_n8202 );
nor  g20751 ( new_n23100 , new_n21328 , new_n21331 );
xnor g20752 ( n16951 , new_n17839 , new_n23100 );
xor  g20753 ( n16954 , new_n15950 , new_n15959 );
xnor g20754 ( n16989 , new_n3704 , new_n8368 );
xnor g20755 ( n17006 , new_n18757 , new_n18787 );
xnor g20756 ( n17068 , new_n13289 , new_n13290 );
xnor g20757 ( n17070 , new_n14963 , new_n14964 );
xnor g20758 ( n17075 , new_n20021 , new_n20065 );
xnor g20759 ( n17084 , new_n16702 , new_n16720 );
xnor g20760 ( n17104 , new_n4746 , new_n4747_1 );
xnor g20761 ( n17106 , new_n13070 , new_n13093 );
xor  g20762 ( n17119 , new_n9681 , new_n9691 );
xnor g20763 ( n17130 , new_n12954 , new_n12987_1 );
xnor g20764 ( n17138 , new_n22308 , new_n22323 );
xnor g20765 ( n17163 , new_n21692 , new_n21700 );
xor  g20766 ( n17168 , new_n19728 , new_n19729 );
xnor g20767 ( n17202 , new_n11397 , new_n11405 );
xor  g20768 ( n17219 , new_n19003 , new_n19005_1 );
xnor g20769 ( n17232 , new_n18244 , new_n18276 );
xnor g20770 ( n17236 , new_n15069 , new_n15072 );
xor  g20771 ( n17243 , new_n10402 , new_n10403 );
xnor g20772 ( n17263 , new_n11056_1 , new_n11072 );
nor  g20773 ( new_n23122 , new_n19155 , new_n19162 );
and  g20774 ( new_n23123 , new_n19164_1 , new_n19186 );
nor  g20775 ( n17285 , new_n23122 , new_n23123 );
xnor g20776 ( n17320 , new_n11546 , new_n11574 );
xnor g20777 ( n17337 , new_n2795 , new_n2843 );
xnor g20778 ( n17344 , new_n21517 , new_n21525_1 );
xnor g20779 ( n17359 , new_n21502 , new_n21533 );
xnor g20780 ( n17387 , new_n13143 , new_n13969 );
xnor g20781 ( n17391 , new_n5081 , new_n5083 );
xnor g20782 ( n17392 , new_n18762 , new_n18782_1 );
xnor g20783 ( n17421 , new_n21771 , new_n21795 );
xnor g20784 ( n17432 , new_n6571 , new_n12037 );
xnor g20785 ( n17436 , new_n20712 , new_n20730 );
xnor g20786 ( n17440 , new_n4710 , new_n22979 );
xnor g20787 ( n17450 , new_n5794 , new_n8458 );
nor  g20788 ( new_n23137 , new_n7362 , new_n18553 );
nor  g20789 ( new_n23138 , new_n7322 , new_n7361 );
nor  g20790 ( new_n23139 , new_n7323 , new_n7362 );
nor  g20791 ( new_n23140 , new_n23139 , new_n7427 );
nor  g20792 ( new_n23141 , new_n23138 , new_n23140 );
nor  g20793 ( new_n23142 , new_n23137 , new_n23141 );
nor  g20794 ( new_n23143 , new_n7361 , new_n18552 );
nor  g20795 ( new_n23144 , new_n23140 , new_n23143 );
nor  g20796 ( n17461 , new_n23142 , new_n23144 );
xor  g20797 ( n17466 , new_n22690 , new_n22691 );
xnor g20798 ( n17493 , new_n13265 , new_n13304 );
xor  g20799 ( n17500 , new_n21197 , new_n21200 );
xnor g20800 ( n17524 , new_n22051 , new_n22054 );
xnor g20801 ( n17529 , new_n5720 , new_n5757 );
xnor g20802 ( new_n23151 , new_n10592 , new_n14770 );
xnor g20803 ( n17557 , new_n14773 , new_n23151 );
xnor g20804 ( n17583 , new_n16328 , new_n16361 );
xnor g20805 ( n17592 , new_n13956 , new_n13978 );
xnor g20806 ( n17638 , new_n8362 , new_n8375 );
xnor g20807 ( n17687 , new_n19545 , new_n19560 );
xnor g20808 ( n17721 , new_n13559 , new_n13592 );
xnor g20809 ( n17735 , new_n21361 , new_n21380 );
and  g20810 ( new_n23159 , new_n10050 , new_n20803_1 );
and  g20811 ( new_n23160_1 , new_n20802 , new_n23159 );
or   g20812 ( new_n23161 , new_n10050 , new_n20803_1 );
nor  g20813 ( new_n23162 , new_n20802 , new_n23161 );
nor  g20814 ( new_n23163 , new_n23160_1 , new_n23162 );
and  g20815 ( new_n23164 , new_n20872 , new_n23163 );
or   g20816 ( new_n23165 , new_n20872 , new_n23163 );
nor  g20817 ( new_n23166_1 , new_n20794_1 , new_n20805 );
nor  g20818 ( new_n23167 , new_n20806 , new_n20815 );
nor  g20819 ( new_n23168 , new_n23166_1 , new_n23167 );
and  g20820 ( new_n23169 , new_n23165 , new_n23168 );
or   g20821 ( new_n23170 , new_n23160_1 , new_n23169 );
nor  g20822 ( n17738 , new_n23164 , new_n23170 );
xor  g20823 ( n17746 , new_n15150 , new_n15153 );
xnor g20824 ( n17749 , new_n22478 , new_n22481 );
xnor g20825 ( n17820 , new_n18417 , new_n18436 );
xnor g20826 ( n17855 , new_n13961 , new_n13976 );
and  g20827 ( new_n23176 , new_n4897 , new_n13919 );
and  g20828 ( new_n23177 , new_n23176 , new_n4965 );
not  g20829 ( new_n23178 , new_n21824 );
nor  g20830 ( new_n23179 , new_n23178 , new_n4965 );
nor  g20831 ( new_n23180 , new_n23177 , new_n23179 );
and  g20832 ( new_n23181 , new_n4796 , new_n4966_1 );
and  g20833 ( new_n23182 , new_n4967_1 , new_n5028 );
or   g20834 ( new_n23183 , new_n23181 , new_n23182 );
and  g20835 ( new_n23184 , new_n23180 , new_n23183 );
nor  g20836 ( n17877 , new_n23177 , new_n23184 );
xnor g20837 ( n17889 , new_n15331 , new_n15332_1 );
and  g20838 ( new_n23187 , new_n22362 , new_n22372 );
nor  g20839 ( new_n23188 , new_n23187 , new_n22384 );
nor  g20840 ( new_n23189 , new_n22362 , new_n22372 );
nor  g20841 ( new_n23190 , new_n23189 , new_n22383 );
nor  g20842 ( n17912 , new_n23188 , new_n23190 );
xor  g20843 ( n17927 , new_n21783 , new_n21786 );
xnor g20844 ( n17931 , new_n21836 , new_n21857 );
xnor g20845 ( n17948 , new_n7891 , new_n7892 );
xor  g20846 ( n17956 , new_n15530 , new_n15533 );
nor  g20847 ( new_n23196 , new_n12442 , new_n12667 );
not  g20848 ( new_n23197 , new_n12592 );
nor  g20849 ( new_n23198 , new_n12442 , new_n23197 );
nor  g20850 ( new_n23199 , new_n23198 , new_n12666 );
nor  g20851 ( n17963 , new_n23196 , new_n23199 );
not  g20852 ( new_n23201 , new_n12948 );
nor  g20853 ( new_n23202 , new_n21940 , n25494 );
and  g20854 ( new_n23203 , new_n17293 , new_n17308 );
nor  g20855 ( new_n23204 , new_n23202 , new_n23203 );
and  g20856 ( new_n23205 , new_n23201 , new_n23204 );
nor  g20857 ( new_n23206 , new_n12952 , new_n23204 );
xnor g20858 ( new_n23207 , new_n12951 , new_n23204 );
and  g20859 ( new_n23208 , new_n12956_1 , new_n17309 );
and  g20860 ( new_n23209 , new_n17310 , new_n17329 );
nor  g20861 ( new_n23210 , new_n23208 , new_n23209 );
and  g20862 ( new_n23211 , new_n23207 , new_n23210 );
nor  g20863 ( new_n23212 , new_n23206 , new_n23211 );
nor  g20864 ( new_n23213 , new_n23205 , new_n23212 );
nor  g20865 ( new_n23214 , new_n23201 , new_n23204 );
nor  g20866 ( new_n23215 , new_n23211 , new_n23214 );
nor  g20867 ( n17976 , new_n23213 , new_n23215 );
xnor g20868 ( n17998 , new_n7132 , new_n7170 );
xnor g20869 ( n18025 , new_n2827 , new_n14391 );
xnor g20870 ( n18043 , new_n20380 , new_n20381 );
xnor g20871 ( n18045 , new_n21711 , new_n21714 );
xnor g20872 ( n18059 , new_n3907 , new_n3918_1 );
xnor g20873 ( n18061 , new_n20024 , new_n20063 );
xnor g20874 ( n18071 , new_n3336 , new_n3391 );
xnor g20875 ( n18143 , new_n9921 , new_n9982 );
xnor g20876 ( n18152 , new_n21195 , new_n21202 );
xnor g20877 ( n18193 , new_n7580 , new_n7588_1 );
xnor g20878 ( new_n23227 , new_n13392 , new_n11615_1 );
xnor g20879 ( n18232 , new_n11628 , new_n23227 );
xnor g20880 ( n18238 , new_n16697 , new_n16722_1 );
xnor g20881 ( n18241 , new_n18262 , new_n18265 );
xnor g20882 ( n18254 , new_n20718 , new_n20726 );
xnor g20883 ( n18288 , new_n21363 , new_n21378 );
xnor g20884 ( n18301 , new_n12066 , new_n12104 );
xnor g20885 ( n18304 , new_n21689 , new_n21702 );
xnor g20886 ( n18310 , new_n13259 , new_n13308 );
xnor g20887 ( n18311 , new_n6667 , new_n6669_1 );
xnor g20888 ( n18323 , new_n17435 , new_n17452 );
xnor g20889 ( n18332 , new_n5411 , new_n5447 );
xor  g20890 ( n18343 , new_n21867 , new_n21868 );
xnor g20891 ( n18350 , new_n19081_1 , new_n19084 );
xnor g20892 ( n18362 , new_n17898 , new_n17899 );
xnor g20893 ( n18377 , new_n4975 , new_n5024_1 );
xnor g20894 ( n18405 , new_n4082 , new_n4102 );
xnor g20895 ( n18414 , new_n16569 , new_n16579 );
xnor g20896 ( n18418 , new_n14462 , new_n14471_1 );
xnor g20897 ( n18437 , new_n8152 , new_n8196 );
xnor g20898 ( n18439 , new_n19837 , new_n19877 );
xnor g20899 ( n18445 , new_n11134_1 , new_n11135 );
xnor g20900 ( n18467 , new_n6920 , new_n6960 );
xnor g20901 ( n18482 , new_n18229 , new_n18282 );
xnor g20902 ( n18509 , new_n18565 , new_n18586 );
xnor g20903 ( n18513 , new_n9039 , new_n13804 );
xnor g20904 ( n18515 , new_n14970 , new_n14972 );
xnor g20905 ( n18572 , new_n15795 , new_n15814 );
and  g20906 ( new_n23255 , new_n23011 , new_n23025 );
nor  g20907 ( new_n23256 , new_n22905 , new_n23255 );
nor  g20908 ( new_n23257 , new_n23011 , new_n23025 );
nor  g20909 ( new_n23258 , new_n22904 , new_n23257 );
nor  g20910 ( n18574 , new_n23256 , new_n23258 );
xnor g20911 ( n18576 , new_n20858 , new_n20861 );
xnor g20912 ( n18582 , new_n22171 , new_n22179 );
xnor g20913 ( n18583 , new_n19635 , new_n19647 );
xnor g20914 ( n18610 , new_n20048 , new_n20049 );
xor  g20915 ( n18635 , new_n21725 , new_n21728 );
xnor g20916 ( n18653 , new_n6739 , new_n6740 );
xnor g20917 ( n18679 , new_n3669 , new_n3721 );
xnor g20918 ( n18693 , new_n20167 , new_n20175 );
xnor g20919 ( n18708 , new_n3045 , new_n3078 );
xnor g20920 ( new_n23269 , new_n22516 , new_n22517 );
xnor g20921 ( n18721 , new_n22522 , new_n23269 );
xnor g20922 ( n18725 , new_n18408 , new_n18442 );
xnor g20923 ( n18751 , new_n20508 , new_n20530 );
xnor g20924 ( n18780 , new_n16338 , new_n16355 );
xnor g20925 ( n18782 , new_n19260 , new_n19303 );
not  g20926 ( new_n23275 , new_n7547 );
and  g20927 ( new_n23276 , new_n7469 , new_n23275 );
nor  g20928 ( new_n23277 , new_n23276 , new_n7606 );
nor  g20929 ( new_n23278 , new_n7469 , new_n23275 );
nor  g20930 ( new_n23279 , new_n23278 , new_n7605 );
nor  g20931 ( n18802 , new_n23277 , new_n23279 );
xor  g20932 ( n18830 , new_n10859 , new_n10860 );
xor  g20933 ( n18831 , new_n12741 , new_n12746_1 );
xnor g20934 ( n18843 , new_n11881 , new_n11888 );
xnor g20935 ( n18858 , new_n3056 , new_n3074 );
xnor g20936 ( n18859 , new_n9950 , new_n9970 );
xnor g20937 ( n18864 , new_n17029 , new_n17078 );
xnor g20938 ( n18865 , new_n4541 , new_n4608 );
xnor g20939 ( n18886 , new_n21128 , new_n21129 );
xnor g20940 ( n18887 , new_n16350_1 , new_n16351 );
xnor g20941 ( n18919 , new_n8866 , new_n8903 );
xnor g20942 ( n18940 , new_n12284 , new_n12296 );
xor  g20943 ( n18945 , new_n22640 , new_n22641 );
xnor g20944 ( n18970 , new_n22342 , new_n22353_1 );
xnor g20945 ( new_n23294 , new_n12064 , new_n16776 );
xnor g20946 ( n18977 , new_n16781 , new_n23294 );
xnor g20947 ( n18982 , new_n15065 , new_n15074 );
xor  g20948 ( n18999 , new_n20614 , new_n20615 );
xnor g20949 ( n19044 , new_n5708 , new_n5763 );
xor  g20950 ( n19125 , new_n14768 , new_n14775 );
xnor g20951 ( n19141 , new_n5712 , new_n5761 );
xnor g20952 ( new_n23301 , new_n13933 , new_n17185 );
nor  g20953 ( new_n23302 , new_n13938 , new_n17188 );
xnor g20954 ( new_n23303 , new_n13938 , new_n17188 );
nor  g20955 ( new_n23304_1 , new_n13941 , new_n17193 );
nor  g20956 ( new_n23305_1 , new_n18454 , new_n18469 );
nor  g20957 ( new_n23306 , new_n23304_1 , new_n23305_1 );
nor  g20958 ( new_n23307 , new_n23303 , new_n23306 );
nor  g20959 ( new_n23308 , new_n23302 , new_n23307 );
xnor g20960 ( n19164 , new_n23301 , new_n23308 );
xnor g20961 ( n19174 , new_n8382 , new_n8383 );
xnor g20962 ( n19176 , new_n20777 , new_n20780 );
xnor g20963 ( n19202 , new_n21686 , new_n21704 );
xnor g20964 ( n19220 , new_n19957 , new_n19968_1 );
xor  g20965 ( n19221 , new_n7850 , new_n7912 );
xnor g20966 ( n19223 , new_n11253 , new_n11254 );
xor  g20967 ( n19224 , new_n17063 , new_n17064 );
xnor g20968 ( n19233 , new_n15469 , new_n15478 );
xnor g20969 ( n19244 , new_n12700 , new_n12730 );
xnor g20970 ( n19314 , new_n8862_1 , new_n8905 );
xnor g20971 ( n19315 , new_n10762 , new_n10763_1 );
xnor g20972 ( n19323 , new_n13272 , new_n13300 );
xnor g20973 ( n19333 , new_n21520 , new_n21523 );
nor  g20974 ( new_n23323 , new_n17177 , new_n17634 );
nor  g20975 ( new_n23324 , new_n9910 , new_n23323 );
nor  g20976 ( new_n23325 , new_n9914 , new_n17183 );
nor  g20977 ( new_n23326 , new_n17184 , new_n17204 );
nor  g20978 ( new_n23327 , new_n23325 , new_n23326 );
not  g20979 ( new_n23328 , new_n23323 );
xnor g20980 ( new_n23329 , new_n9910 , new_n23328 );
and  g20981 ( new_n23330 , new_n23327 , new_n23329 );
nor  g20982 ( n19348 , new_n23324 , new_n23330 );
xnor g20983 ( n19354 , new_n16670 , new_n16734 );
xnor g20984 ( n19367 , new_n11045 , new_n11079 );
xnor g20985 ( n19385 , new_n18902 , new_n18923 );
xnor g20986 ( new_n23335 , new_n16797 , new_n16849 );
xnor g20987 ( n19389 , new_n16878 , new_n23335 );
xnor g20988 ( n19401 , new_n16193 , new_n16223_1 );
xor  g20989 ( n19414 , new_n21959 , new_n21967 );
xnor g20990 ( n19424 , new_n17721_1 , new_n19103 );
xnor g20991 ( n19450 , new_n21115 , new_n21133 );
nor  g20992 ( new_n23341_1 , new_n13870 , new_n23328 );
xnor g20993 ( new_n23342_1 , new_n13870 , new_n23328 );
nor  g20994 ( new_n23343 , new_n13928 , new_n17183 );
xnor g20995 ( new_n23344 , new_n13928 , new_n17183 );
nor  g20996 ( new_n23345 , new_n13933 , new_n17185 );
nor  g20997 ( new_n23346 , new_n23301 , new_n23308 );
nor  g20998 ( new_n23347 , new_n23345 , new_n23346 );
nor  g20999 ( new_n23348 , new_n23344 , new_n23347 );
nor  g21000 ( new_n23349 , new_n23343 , new_n23348 );
nor  g21001 ( new_n23350 , new_n23342_1 , new_n23349 );
or   g21002 ( n19458 , new_n23341_1 , new_n23350 );
xnor g21003 ( n19467 , new_n15146_1 , new_n15155 );
xnor g21004 ( n19496 , new_n8147 , new_n8198 );
xor  g21005 ( n19523 , new_n15107 , new_n15115 );
xnor g21006 ( n19570 , new_n4561 , new_n4600 );
xnor g21007 ( n19602 , new_n11996 , new_n12006 );
xnor g21008 ( n19617 , new_n12334 , new_n12339 );
xnor g21009 ( n19623 , new_n13562 , new_n13590 );
xor  g21010 ( n19641 , new_n22006 , new_n22008 );
xnor g21011 ( n19648 , new_n21768 , new_n21797 );
xnor g21012 ( n19664 , new_n15799 , new_n15812_1 );
xnor g21013 ( n19736 , new_n19713 , new_n19726 );
nor  g21014 ( new_n23363 , new_n21955 , new_n21969 );
nor  g21015 ( new_n23364 , new_n3197 , new_n21955 );
nor  g21016 ( new_n23365 , new_n23364 , new_n21968 );
nor  g21017 ( n19749 , new_n23363 , new_n23365 );
xnor g21018 ( n19756 , new_n14827_1 , new_n14840 );
xnor g21019 ( n19767 , new_n12003_1 , new_n12004 );
xor  g21020 ( new_n23369_1 , new_n3327 , new_n3330 );
xnor g21021 ( n19780 , new_n3393 , new_n23369_1 );
xnor g21022 ( n19792 , new_n22541 , new_n22544 );
xnor g21023 ( n19798 , new_n20357 , new_n20370 );
xor  g21024 ( n19873 , new_n16442 , new_n16445_1 );
nor  g21025 ( new_n23374 , new_n18294 , new_n18313 );
not  g21026 ( new_n23375 , new_n18300 );
nor  g21027 ( new_n23376 , new_n18294 , new_n23375 );
nor  g21028 ( new_n23377 , new_n23376 , new_n18312 );
nor  g21029 ( n19909 , new_n23374 , new_n23377 );
xnor g21030 ( n19916 , new_n19716 , new_n19724 );
xnor g21031 ( n19923 , new_n20350 , new_n20374 );
xnor g21032 ( n19930 , new_n18754 , new_n18789 );
xnor g21033 ( n19968 , new_n6317 , new_n6423 );
xnor g21034 ( n19988 , new_n19279 , new_n19291 );
and  g21035 ( new_n23384 , new_n20438 , new_n21157_1 );
nor  g21036 ( new_n23385 , new_n10099 , new_n20438 );
nor  g21037 ( new_n23386 , new_n20439 , new_n20442 );
nor  g21038 ( new_n23387 , new_n23385 , new_n23386 );
nor  g21039 ( new_n23388 , new_n23384 , new_n23387 );
nor  g21040 ( new_n23389 , new_n20438 , new_n21157_1 );
nor  g21041 ( new_n23390 , new_n23386 , new_n23389 );
nor  g21042 ( n20004 , new_n23388 , new_n23390 );
xnor g21043 ( n20017 , new_n20512 , new_n20526 );
xnor g21044 ( n20033 , new_n18239 , new_n18278 );
xnor g21045 ( n20061 , new_n13770 , new_n13771 );
xnor g21046 ( n20069 , new_n17848 , new_n17851 );
nor  g21047 ( new_n23396 , new_n14346 , new_n14357 );
nor  g21048 ( new_n23397 , new_n14358 , new_n14413 );
or   g21049 ( n20086 , new_n23396 , new_n23397 );
xnor g21050 ( n20096 , new_n19175 , new_n19178 );
xnor g21051 ( n20103 , new_n13285_1 , new_n13292 );
xnor g21052 ( n20126 , new_n11542 , new_n11576 );
xnor g21053 ( n20149 , new_n20902 , new_n20931 );
xnor g21054 ( n20187 , new_n11861 , new_n11900 );
xnor g21055 ( n20279 , new_n17261 , new_n17289 );
and  g21056 ( new_n23405 , new_n22158 , new_n22164 );
nor  g21057 ( new_n23406 , new_n23405 , new_n22167 );
nor  g21058 ( new_n23407 , new_n22164 , new_n22182 );
nor  g21059 ( new_n23408 , new_n17427 , new_n22181 );
nor  g21060 ( new_n23409 , new_n23407 , new_n23408 );
and  g21061 ( n20287 , new_n23406 , new_n23409 );
xnor g21062 ( n20301 , new_n20207 , new_n20210 );
nor  g21063 ( new_n23412 , new_n8133 , new_n8204 );
nor  g21064 ( n20330 , new_n8028 , new_n23412 );
xnor g21065 ( n20333 , new_n11868 , new_n11896 );
and  g21066 ( new_n23415 , new_n10210 , new_n10346 );
and  g21067 ( new_n23416 , new_n23415 , new_n10410 );
or   g21068 ( new_n23417 , new_n10210 , new_n10346 );
nor  g21069 ( new_n23418 , new_n23417 , new_n10410 );
or   g21070 ( n20355 , new_n23416 , new_n23418 );
xnor g21071 ( n20366 , new_n5201 , new_n8418 );
xnor g21072 ( n20388 , new_n18953 , new_n18956 );
xnor g21073 ( n20402 , new_n21838 , new_n21855 );
xnor g21074 ( n20403 , new_n15293 , new_n15319 );
xnor g21075 ( n20424 , new_n3062 , new_n22404 );
xnor g21076 ( n20436 , new_n20042 , new_n20053 );
xor  g21077 ( n20441 , new_n8182 , new_n8184 );
xnor g21078 ( n20445 , new_n7552 , new_n7604 );
xnor g21079 ( n20450 , new_n4971 , new_n5026_1 );
xnor g21080 ( n20490 , new_n16365 , new_n16367_1 );
xor  g21081 ( n20495 , new_n19962 , new_n19966 );
and  g21082 ( new_n23431 , new_n15335 , new_n15337 );
and  g21083 ( new_n23432 , new_n15334 , new_n23431 );
or   g21084 ( new_n23433_1 , new_n15335 , new_n15337 );
nor  g21085 ( new_n23434_1 , new_n15334 , new_n23433_1 );
or   g21086 ( n20515 , new_n23432 , new_n23434_1 );
nor  g21087 ( new_n23436 , new_n22536 , new_n22546 );
nor  g21088 ( n20533 , new_n22531 , new_n23436 );
xnor g21089 ( n20582 , new_n17716 , new_n17723 );
xnor g21090 ( n20590 , new_n19423 , new_n19451 );
xnor g21091 ( n20602 , new_n3373 , new_n3375 );
xnor g21092 ( n20609 , new_n16347 , new_n16348 );
xnor g21093 ( n20623 , new_n6567_1 , new_n6575 );
xnor g21094 ( n20629 , new_n20336 , new_n20385_1 );
xnor g21095 ( n20661 , new_n13759 , new_n13768 );
xnor g21096 ( n20673 , new_n8461 , new_n8463 );
xnor g21097 ( n20678 , new_n20344 , new_n20378 );
nor  g21098 ( new_n23447 , new_n11793 , new_n14816 );
nor  g21099 ( new_n23448 , new_n23447 , new_n14847 );
and  g21100 ( new_n23449 , new_n11793 , new_n14816 );
or   g21101 ( new_n23450_1 , new_n14813 , new_n23449 );
nor  g21102 ( n20680 , new_n23448 , new_n23450_1 );
xnor g21103 ( n20685 , new_n4157 , new_n6401 );
xnor g21104 ( new_n23453 , new_n12948 , new_n23204 );
xnor g21105 ( n20691 , new_n23212 , new_n23453 );
xnor g21106 ( n20696 , new_n15802 , new_n15810 );
xnor g21107 ( n20704 , new_n22311_1 , new_n22321 );
xor  g21108 ( n20705 , new_n21371 , new_n21372 );
xnor g21109 ( n20709 , new_n9926_1 , new_n9980 );
xnor g21110 ( n20713 , new_n14708 , new_n14732 );
xnor g21111 ( n20722 , new_n8633 , new_n8634 );
not  g21112 ( new_n23461 , new_n19347 );
nor  g21113 ( new_n23462 , new_n23461 , new_n22817 );
nor  g21114 ( new_n23463_1 , new_n19336 , new_n19347 );
nor  g21115 ( new_n23464 , new_n19335 , new_n23461 );
nor  g21116 ( new_n23465 , new_n23464 , new_n19359 );
nor  g21117 ( new_n23466 , new_n23463_1 , new_n23465 );
nor  g21118 ( new_n23467 , new_n23462 , new_n23466 );
nor  g21119 ( new_n23468 , new_n19347 , new_n22818 );
nor  g21120 ( new_n23469 , new_n23465 , new_n23468 );
nor  g21121 ( n20723 , new_n23467 , new_n23469 );
xnor g21122 ( new_n23471_1 , new_n17428 , new_n22159 );
xnor g21123 ( n20748 , new_n22182 , new_n23471_1 );
xor  g21124 ( n20761 , new_n5429 , new_n5439_1 );
xnor g21125 ( n20774 , new_n20028 , new_n20061_1 );
xnor g21126 ( n20788 , new_n23342_1 , new_n23349 );
nor  g21127 ( new_n23476 , new_n21722 , new_n22669 );
nor  g21128 ( new_n23477 , new_n22779_1 , new_n23476 );
nor  g21129 ( new_n23478 , new_n21723 , new_n22775 );
nor  g21130 ( new_n23479 , new_n22778 , new_n23478 );
nor  g21131 ( n20795 , new_n23477 , new_n23479 );
xnor g21132 ( new_n23481 , new_n20082 , new_n20093 );
and  g21133 ( new_n23482 , new_n20082 , new_n20102 );
nor  g21134 ( new_n23483 , new_n20104 , new_n23482 );
nor  g21135 ( new_n23484 , new_n20103_1 , new_n23483 );
xnor g21136 ( n20803 , new_n23481 , new_n23484 );
xor  g21137 ( n20869 , new_n23180 , new_n23183 );
xnor g21138 ( n20879 , new_n22475 , new_n22483 );
xnor g21139 ( n20915 , new_n6384 , new_n6411 );
xnor g21140 ( new_n23489 , n2160 , n19282 );
nor  g21141 ( new_n23490 , new_n11674_1 , n12657 );
and  g21142 ( new_n23491 , new_n21385 , new_n21388 );
or   g21143 ( new_n23492 , new_n23490 , new_n23491 );
xor  g21144 ( new_n23493_1 , new_n23489 , new_n23492 );
nor  g21145 ( new_n23494 , new_n22379_1 , new_n23493_1 );
nor  g21146 ( new_n23495 , new_n19678 , new_n21389 );
nor  g21147 ( new_n23496 , new_n21390 , new_n21393 );
nor  g21148 ( new_n23497 , new_n23495 , new_n23496 );
xnor g21149 ( new_n23498 , new_n22379_1 , new_n23493_1 );
nor  g21150 ( new_n23499 , new_n23497 , new_n23498 );
nor  g21151 ( new_n23500 , new_n23494 , new_n23499 );
not  g21152 ( new_n23501 , new_n23500 );
nor  g21153 ( new_n23502 , new_n12808 , n19282 );
and  g21154 ( new_n23503 , new_n23489 , new_n23492 );
nor  g21155 ( new_n23504 , new_n23502 , new_n23503 );
and  g21156 ( new_n23505 , new_n22377 , new_n23504 );
and  g21157 ( new_n23506 , new_n23501 , new_n23505 );
and  g21158 ( new_n23507 , new_n22372 , new_n23506 );
or   g21159 ( new_n23508 , new_n22377 , new_n23504 );
nor  g21160 ( new_n23509 , new_n23501 , new_n23508 );
and  g21161 ( new_n23510 , new_n22373 , new_n23509 );
or   g21162 ( n20935 , new_n23507 , new_n23510 );
xnor g21163 ( n20936 , new_n21777 , new_n21791 );
xnor g21164 ( n21008 , new_n16762 , new_n16763 );
xnor g21165 ( n21017 , new_n19263 , new_n19301 );
and  g21166 ( new_n23515 , new_n21226_1 , new_n22883 );
nor  g21167 ( new_n23516 , new_n21226_1 , new_n22883 );
nor  g21168 ( new_n23517 , new_n23516 , new_n22888 );
or   g21169 ( new_n23518 , new_n22882 , new_n23517 );
nor  g21170 ( n21034 , new_n23515 , new_n23518 );
xor  g21171 ( n21046 , new_n21931 , new_n21932 );
xnor g21172 ( n21062 , new_n8545 , new_n8564 );
xor  g21173 ( new_n23522 , new_n22616 , new_n22624 );
xnor g21174 ( n21093 , new_n22531 , new_n23522 );
xnor g21175 ( n21094 , new_n7884_1 , new_n9725 );
xnor g21176 ( n21123 , new_n14599 , new_n14622 );
xnor g21177 ( n21154 , new_n17923 , new_n18686 );
xnor g21178 ( n21157 , new_n15431 , new_n15453 );
xnor g21179 ( n21168 , new_n20915_1 , new_n20923_1 );
xnor g21180 ( n21173 , new_n7398 , new_n7400 );
xnor g21181 ( n21176 , new_n4571 , new_n4596 );
xnor g21182 ( n21182 , new_n14272 , new_n14279 );
nor  g21183 ( new_n23532 , new_n20949 , new_n21762 );
nor  g21184 ( new_n23533 , new_n20950 , new_n21800_1 );
nor  g21185 ( new_n23534 , new_n23532 , new_n23533 );
nor  g21186 ( new_n23535 , new_n20960 , new_n21799 );
nor  g21187 ( new_n23536 , new_n21765_1 , new_n23535 );
and  g21188 ( n21193 , new_n23534 , new_n23536 );
xnor g21189 ( n21203 , new_n9468 , new_n9469 );
xnor g21190 ( n21225 , new_n2544 , new_n16346 );
xnor g21191 ( n21238 , new_n19614 , new_n19661 );
xnor g21192 ( n21254 , new_n13754_1 , new_n13773 );
xnor g21193 ( n21298 , new_n19845 , new_n19873_1 );
xnor g21194 ( n21302 , new_n9376 , new_n19641_1 );
xnor g21195 ( n21349 , new_n19719 , new_n19722 );
xnor g21196 ( n21365 , new_n15961 , new_n15962 );
xnor g21197 ( n21367 , new_n15104 , new_n15117 );
xnor g21198 ( n21396 , new_n11755 , new_n11783 );
xnor g21199 ( n21399 , new_n7556 , new_n7602 );
xnor g21200 ( n21404 , new_n3396 , new_n3401 );
xnor g21201 ( n21446 , new_n8454 , new_n8465 );
xnor g21202 ( n21472 , new_n11618 , new_n11626 );
xnor g21203 ( n21525 , new_n7375 , new_n7421_1 );
xnor g21204 ( n21549 , new_n17102 , new_n17126 );
xnor g21205 ( n21615 , new_n19553 , new_n19556 );
nor  g21206 ( new_n23555 , new_n7835 , new_n22164 );
xnor g21207 ( new_n23556 , new_n13394 , new_n22164 );
nor  g21208 ( new_n23557 , new_n13394 , new_n17427 );
and  g21209 ( new_n23558 , new_n17429 , new_n17457 );
or   g21210 ( new_n23559 , new_n23557 , new_n23558 );
and  g21211 ( new_n23560 , new_n23556 , new_n23559 );
nor  g21212 ( n21628 , new_n23555 , new_n23560 );
nor  g21213 ( new_n23562 , new_n20955 , new_n21433 );
xnor g21214 ( new_n23563 , new_n20957 , new_n21433 );
nor  g21215 ( new_n23564 , new_n20957 , new_n21437 );
nor  g21216 ( new_n23565 , new_n22742 , new_n22745 );
or   g21217 ( new_n23566 , new_n23564 , new_n23565 );
and  g21218 ( new_n23567 , new_n23563 , new_n23566 );
nor  g21219 ( n21637 , new_n23562 , new_n23567 );
xnor g21220 ( n21645 , new_n21367_1 , new_n21374 );
xnor g21221 ( n21665 , new_n22664 , new_n12032 );
xnor g21222 ( n21680 , new_n14821 , new_n14844 );
xnor g21223 ( n21685 , new_n21830 , new_n21863 );
xnor g21224 ( n21717 , new_n18414_1 , new_n18438 );
xnor g21225 ( n21719 , new_n16746 , new_n16751 );
xnor g21226 ( n21750 , new_n18427 , new_n18430 );
xnor g21227 ( n21765 , new_n21625 , new_n21626 );
xnor g21228 ( n21800 , new_n23497 , new_n23498 );
xnor g21229 ( new_n23578 , new_n4296 , new_n4299 );
xnor g21230 ( n21820 , new_n4304 , new_n23578 );
xnor g21231 ( n21874 , new_n19273 , new_n19295 );
xnor g21232 ( n21943 , new_n13282 , new_n13294 );
xnor g21233 ( n21960 , new_n15945 , new_n15966 );
xnor g21234 ( n21976 , new_n7157 , new_n7159 );
xnor g21235 ( n21986 , new_n11235 , new_n11263 );
xnor g21236 ( n22016 , new_n11041 , new_n11081 );
xnor g21237 ( n22027 , new_n18423 , new_n18432 );
xnor g21238 ( n22050 , new_n13080 , new_n13089 );
xnor g21239 ( n22063 , new_n4157 , new_n4158 );
xnor g21240 ( n22076 , new_n20918 , new_n20921 );
nor  g21241 ( new_n23590 , new_n13736 , new_n20086_1 );
and  g21242 ( new_n23591 , new_n20414 , new_n20433 );
nor  g21243 ( n22090 , new_n23590 , new_n23591 );
xnor g21244 ( n22107 , new_n22344 , new_n22351 );
xnor g21245 ( n22113 , new_n17593 , new_n17619 );
nor  g21246 ( new_n23595 , new_n13673 , new_n13735 );
nor  g21247 ( new_n23596 , new_n23595 , new_n13781_1 );
nor  g21248 ( new_n23597 , new_n13674 , new_n13736 );
nor  g21249 ( new_n23598 , new_n23597 , new_n13780 );
nor  g21250 ( n22124 , new_n23596 , new_n23598 );
nor  g21251 ( new_n23600 , new_n19162 , new_n22984 );
and  g21252 ( new_n23601 , new_n22985 , new_n22988 );
nor  g21253 ( n22126 , new_n23600 , new_n23601 );
nor  g21254 ( new_n23603 , new_n23506 , new_n23509 );
xnor g21255 ( n22130 , new_n22373 , new_n23603 );
xor  g21256 ( n22144 , new_n17798 , new_n17799 );
xnor g21257 ( n22150 , new_n22732 , new_n22736 );
xnor g21258 ( n22157 , new_n19484 , new_n19490 );
xnor g21259 ( n22213 , new_n23303 , new_n23306 );
xnor g21260 ( n22283 , new_n10388_1 , new_n10389 );
xor  g21261 ( n22311 , new_n20122 , new_n20123 );
xnor g21262 ( n22317 , new_n8858 , new_n8907 );
xnor g21263 ( n22341 , new_n17371 , new_n17384 );
nor  g21264 ( new_n23613 , new_n7182 , new_n7194 );
and  g21265 ( new_n23614 , new_n7178 , new_n23613 );
nand g21266 ( new_n23615 , new_n7182 , new_n7194 );
nor  g21267 ( new_n23616 , new_n7178 , new_n23615 );
nor  g21268 ( new_n23617 , new_n23614 , new_n23616 );
xnor g21269 ( n22353 , new_n18081 , new_n23617 );
xnor g21270 ( n22444 , new_n17374 , new_n17382 );
xnor g21271 ( n22467 , new_n10141 , new_n10143 );
xnor g21272 ( n22484 , new_n8885 , new_n20132 );
xnor g21273 ( n22489 , new_n4546 , new_n4606 );
xnor g21274 ( n22494 , new_n8344 , new_n8389 );
xnor g21275 ( n22533 , new_n10373 , new_n10395 );
xnor g21276 ( n22584 , new_n22317_1 , new_n22319 );
nor  g21277 ( new_n23626 , new_n17783 , new_n17805 );
nor  g21278 ( n22589 , new_n17744 , new_n23626 );
xnor g21279 ( n22620 , new_n23344 , new_n23347 );
xnor g21280 ( n22623 , new_n8459 , new_n8460 );
xnor g21281 ( n22697 , new_n16860 , new_n16874 );
xnor g21282 ( n22714 , new_n8879 , new_n8897 );
xnor g21283 ( n22761 , new_n11854 , new_n11904 );
xnor g21284 ( n22779 , new_n18836 , new_n18852 );
xnor g21285 ( n22787 , new_n22299 , new_n22329 );
xnor g21286 ( n22819 , new_n2506 , new_n2538 );
xnor g21287 ( n22858 , new_n4586 , new_n9203 );
xnor g21288 ( new_n23637_1 , new_n11592 , new_n20987 );
xnor g21289 ( n22870 , new_n22797 , new_n23637_1 );
xor  g21290 ( n22891 , new_n9676 , new_n9693 );
xor  g21291 ( n22897 , new_n19431 , new_n19444 );
xnor g21292 ( n22903 , new_n10104 , new_n10161 );
xnor g21293 ( n22907 , new_n14251 , new_n14293 );
xnor g21294 ( n22910 , new_n7163 , new_n7164 );
xnor g21295 ( n22914 , new_n12315_1 , new_n12321 );
xnor g21296 ( n22939 , new_n5853 , new_n5769 );
xnor g21297 ( new_n23646 , new_n4417 , new_n18961 );
xnor g21298 ( n22998 , new_n18959 , new_n23646 );
xnor g21299 ( n23006 , new_n8892 , new_n8893 );
xnor g21300 ( n23007 , new_n12739 , new_n12748 );
xnor g21301 ( n23009 , new_n17987 , new_n17990 );
xnor g21302 ( n23014 , new_n16675 , new_n16732 );
xor  g21303 ( n23047 , new_n23563 , new_n23566 );
xnor g21304 ( n23058 , new_n17438 , new_n17450_1 );
and  g21305 ( n23066 , new_n18446 , new_n18451 );
and  g21306 ( new_n23655 , new_n10209 , new_n18339 );
nor  g21307 ( new_n23656 , new_n18341 , new_n23655 );
xor  g21308 ( n23067 , new_n18336 , new_n23656 );
xor  g21309 ( n23238 , new_n15952 , new_n15957 );
xnor g21310 ( n23247 , new_n17187 , new_n17202_1 );
xor  g21311 ( n23248 , new_n14958 , new_n14966 );
xnor g21312 ( n23270 , new_n17270 , new_n17281 );
xnor g21313 ( n23289 , new_n22378 , new_n22382 );
xnor g21314 ( n23305 , new_n5406 , new_n5449 );
xnor g21315 ( n23341 , new_n20721 , new_n20724 );
xnor g21316 ( n23342 , new_n4943 , new_n9376 );
and  g21317 ( new_n23666 , new_n23275 , new_n21028 );
nor  g21318 ( new_n23667 , new_n23666 , new_n21052 );
nor  g21319 ( new_n23668 , new_n23275 , new_n21028 );
nor  g21320 ( new_n23669_1 , new_n23668 , new_n21051 );
nor  g21321 ( n23355 , new_n23667 , new_n23669_1 );
xnor g21322 ( n23371 , new_n19052 , new_n19055 );
xnor g21323 ( n23401 , new_n15284 , new_n15323 );
xnor g21324 ( n23414 , new_n13086 , new_n13087 );
xnor g21325 ( n23429 , new_n17264 , new_n17287 );
nor  g21326 ( new_n23675 , new_n21274 , new_n21280 );
not  g21327 ( new_n23676 , new_n21276_1 );
nor  g21328 ( new_n23677 , new_n21274 , new_n23676 );
nor  g21329 ( new_n23678 , new_n21279 , new_n23677 );
nor  g21330 ( n23433 , new_n23675 , new_n23678 );
xnor g21331 ( n23434 , new_n18256 , new_n18270 );
nor  g21332 ( new_n23681 , new_n21402 , new_n22984 );
nor  g21333 ( new_n23682 , new_n23001 , new_n23681 );
nor  g21334 ( new_n23683 , new_n21401 , new_n22983 );
nor  g21335 ( new_n23684_1 , new_n23000 , new_n23683 );
nor  g21336 ( n23450 , new_n23682 , new_n23684_1 );
xnor g21337 ( n23471 , new_n16679 , new_n16730 );
xnor g21338 ( n23480 , new_n20706 , new_n20734 );
xor  g21339 ( n23546 , new_n17646 , new_n17651 );
xnor g21340 ( n23550 , new_n20360 , new_n20368 );
xnor g21341 ( n23585 , new_n7387 , new_n7415 );
xor  g21342 ( n23588 , new_n19434 , new_n19442 );
xor  g21343 ( n23619 , new_n20611 , new_n20612 );
xnor g21344 ( n23624 , new_n3061 , new_n3072 );
xnor g21345 ( n23628 , new_n11768 , new_n11775_1 );
xnor g21346 ( n23637 , new_n21514 , new_n21527 );
xnor g21347 ( n23663 , new_n22110 , new_n22113_1 );
xnor g21348 ( n23669 , new_n11764 , new_n11777 );
xnor g21349 ( n23684 , new_n12958 , new_n12985_1 );
xnor g21350 ( n23690 , new_n18768 , new_n18777 );
xnor g21351 ( n23714 , new_n21832_1 , new_n21861 );
nor  g21352 ( n23719 , new_n23032 , new_n23035_1 );
xnor g21353 ( n23748 , new_n20998 , new_n21001 );
xnor g21354 ( n23856 , new_n7198 , new_n10855 );
xnor g21355 ( n23883 , new_n7412 , new_n7413 );
xnor g21356 ( new_n23705 , new_n5809 , new_n14273 );
xnor g21357 ( n23888 , new_n14276 , new_n23705 );
xnor g21358 ( n23899 , new_n3356 , new_n3381 );
xnor g21359 ( n23903 , new_n9461 , new_n14772_1 );
xnor g21360 ( n23924 , new_n12702_1 , new_n12728 );
xnor g21361 ( n23935 , new_n16409 , new_n16410 );
xnor g21362 ( n23942 , new_n12966 , new_n12981 );
xnor g21363 ( n23954 , new_n17475 , new_n17483 );
xnor g21364 ( n23958 , new_n18496_1 , new_n18516 );
xor  g21365 ( n23986 , new_n21991 , new_n21992 );
xor  g21366 ( n24002 , new_n16760 , new_n16765 );
xnor g21367 ( n24039 , new_n12868 , new_n12876 );
xnor g21368 ( n24052 , new_n22966 , new_n22967 );
xnor g21369 ( n24092 , new_n20038 , new_n20055 );
xnor g21370 ( n24096 , new_n15448 , new_n15449 );
xnor g21371 ( n24097 , new_n12072_1 , new_n12097 );
xnor g21372 ( n24105 , new_n11758 , new_n11781 );
xnor g21373 ( n24119 , new_n17954_1 , new_n17972 );
xnor g21374 ( n24133 , new_n14824 , new_n14842 );
xnor g21375 ( n24141 , new_n19626 , new_n19653 );
xnor g21376 ( new_n23725 , new_n20873 , new_n20897 );
xnor g21377 ( n24145 , new_n20933 , new_n23725 );
xnor g21378 ( n24146 , new_n21599_1 , new_n21602 );
xnor g21379 ( n24155 , new_n12609 , new_n12661 );
xnor g21380 ( n24160 , new_n23207 , new_n23210 );
xnor g21381 ( n24167 , new_n9185 , new_n9217_1 );
and  g21382 ( n24172 , new_n20178 , new_n20183 );
xnor g21383 ( n24177 , new_n14269 , new_n14281 );
xor  g21384 ( n24228 , new_n23071 , new_n23072 );
xnor g21385 ( n24258 , new_n17368 , new_n17386 );
nor  g21386 ( new_n23735 , new_n7182 , new_n18081 );
and  g21387 ( new_n23736 , new_n18083 , new_n23616 );
nor  g21388 ( new_n23737 , new_n23614 , new_n23736 );
nor  g21389 ( n24260 , new_n23735 , new_n23737 );
xnor g21390 ( n24289 , new_n18830_1 , new_n18856 );
xnor g21391 ( n24297 , new_n4738 , new_n4749 );
xnor g21392 ( n24307 , new_n3909_1 , new_n11773 );
xnor g21393 ( n24342 , new_n2520 , new_n2532 );
xnor g21394 ( n24345 , new_n15947_1 , new_n15964 );
xnor g21395 ( n24347 , new_n9459_1 , new_n9471 );
xnor g21396 ( n24373 , new_n4979 , new_n5022 );
xnor g21397 ( n24406 , new_n21267 , new_n17911_1 );
xnor g21398 ( n24415 , new_n13626_1 , new_n13638 );
xnor g21399 ( n24421 , new_n10756_1 , new_n10758 );
xnor g21400 ( n24431 , new_n13457_1 , new_n13480 );
xnor g21401 ( n24472 , new_n11871 , new_n11894 );
and  g21402 ( new_n23751 , new_n21918 , new_n22389 );
nor  g21403 ( new_n23752 , new_n22391 , new_n23751 );
xor  g21404 ( n24476 , new_n22386 , new_n23752 );
xnor g21405 ( n24483 , new_n10116 , new_n10155 );
xnor g21406 ( n24501 , new_n13376 , new_n22896 );
xnor g21407 ( n24512 , new_n18008 , new_n18011 );
xnor g21408 ( n24558 , new_n4751 , new_n4752 );
xnor g21409 ( n24576 , new_n2826_1 , new_n2829 );
xnor g21410 ( n24579 , new_n2830 , new_n2831 );
xnor g21411 ( n24602 , new_n20115 , new_n20127 );
xnor g21412 ( n24604 , new_n14123 , new_n14156 );
xnor g21413 ( n24626 , new_n22500 , new_n22503 );
xnor g21414 ( n24629 , new_n21610 , new_n21612 );
xnor g21415 ( n24636 , new_n21365_1 , new_n21376 );
xnor g21416 ( n24715 , new_n21123_1 , new_n21126 );
xnor g21417 ( n24723 , new_n20018 , new_n20067 );
xnor g21418 ( new_n23767 , new_n16627 , new_n16666 );
xnor g21419 ( n24749 , new_n16736 , new_n23767 );
xnor g21420 ( n24758 , new_n20035 , new_n20057 );
xnor g21421 ( n24784 , new_n22576 , new_n22579 );
xnor g21422 ( n24807 , new_n16116 , new_n16117 );
xnor g21423 ( n24826 , new_n7889 , new_n9720 );
xnor g21424 ( n24840 , new_n7564 , new_n7598_1 );
xnor g21425 ( n24841 , new_n9955 , new_n9968_1 );
xnor g21426 ( n24853 , new_n5199 , new_n5211_1 );
xnor g21427 ( n24857 , new_n3051 , new_n3076_1 );
xnor g21428 ( n24887 , new_n6393 , new_n6407_1 );
xor  g21429 ( n24934 , new_n9200 , new_n9207 );
xnor g21430 ( n24998 , new_n7367 , new_n7425 );
xnor g21431 ( n25006 , new_n11555 , new_n11567 );
xnor g21432 ( n25032 , new_n20418 , new_n20429_1 );
xnor g21433 ( n25062 , new_n16050 , new_n16068_1 );
xnor g21434 ( new_n23783 , new_n16627 , new_n19253 );
xnor g21435 ( n25083 , new_n19307 , new_n23783 );
xor  g21436 ( n25097 , new_n12974 , new_n12977 );
xnor g21437 ( n25133 , new_n17641 , new_n17644 );
xnor g21438 ( n25155 , new_n18253 , new_n18272 );
xnor g21439 ( new_n23788 , new_n22377 , new_n23504 );
xnor g21440 ( n25181 , new_n23501 , new_n23788 );
xnor g21441 ( n25200 , new_n20416 , new_n20431 );
nor  g21442 ( new_n23791 , new_n21138_1 , new_n21141 );
xnor g21443 ( new_n23792 , new_n16797 , new_n21135 );
xnor g21444 ( n25209 , new_n23791 , new_n23792 );
xnor g21445 ( n25215 , new_n15037 , new_n15038 );
xor  g21446 ( n25244 , new_n18084 , new_n18087 );
xnor g21447 ( n25254 , new_n17708 , new_n17727 );
xor  g21448 ( n25256 , new_n20590_1 , new_n20617 );
nor  g21449 ( new_n23798 , new_n21220 , new_n22929 );
nor  g21450 ( new_n23799 , new_n22935 , new_n23798 );
xnor g21451 ( new_n23800 , new_n22007 , new_n22928 );
xnor g21452 ( n25293 , new_n23799 , new_n23800 );
xor  g21453 ( n25328 , new_n20600 , new_n20607 );
xnor g21454 ( n25332 , new_n4301 , new_n11060 );
nor  g21455 ( new_n23804 , new_n21291 , new_n22564 );
nor  g21456 ( new_n23805 , new_n23804 , new_n22587 );
and  g21457 ( new_n23806 , new_n21291 , new_n22564 );
nor  g21458 ( new_n23807 , new_n23806 , new_n22586 );
nor  g21459 ( n25337 , new_n23805 , new_n23807 );
xnor g21460 ( new_n23809 , new_n10840 , new_n11398_1 );
xnor g21461 ( n25356 , new_n11403_1 , new_n23809 );
xnor g21462 ( n25362 , new_n9031 , new_n9042_1 );
xnor g21463 ( n25412 , new_n14382 , new_n14399 );
xor  g21464 ( n25460 , new_n15311 , new_n15312 );
xnor g21465 ( n25468 , new_n7383 , new_n7417 );
xnor g21466 ( n25499 , new_n14379 , new_n14401 );
xnor g21467 ( n25513 , new_n19642 , new_n19643 );
xnor g21468 ( n25518 , new_n12074 , new_n12095 );
xnor g21469 ( n25532 , new_n13268 , new_n13302 );
xnor g21470 ( n25539 , new_n19952 , new_n19970 );
xnor g21471 ( n25550 , new_n16864 , new_n16872 );
xnor g21472 ( n25611 , new_n20715 , new_n20728 );
xnor g21473 ( new_n23822 , new_n5432 , new_n5433 );
xnor g21474 ( n25614 , new_n5437 , new_n23822 );
xnor g21475 ( n25619 , new_n12705 , new_n12726 );
nor  g21476 ( new_n23825 , new_n22682 , new_n22818 );
nor  g21477 ( new_n23826 , new_n23825 , new_n22823 );
nor  g21478 ( new_n23827 , new_n22683 , new_n22817 );
nor  g21479 ( new_n23828 , new_n23827 , new_n22822 );
nor  g21480 ( n25665 , new_n23826 , new_n23828 );
xnor g21481 ( n25706 , new_n9191_1 , new_n9213 );
xnor g21482 ( new_n23831_1 , new_n23461 , new_n22818 );
xnor g21483 ( n25719 , new_n23466 , new_n23831_1 );
xor  g21484 ( n25756 , new_n9655_1 , new_n9701 );
and  g21485 ( new_n23834 , new_n12904_1 , new_n23201 );
nor  g21486 ( new_n23835 , new_n23834 , new_n12989 );
nor  g21487 ( new_n23836 , new_n12904_1 , new_n23201 );
nor  g21488 ( new_n23837 , new_n23836 , new_n12988 );
nor  g21489 ( n25758 , new_n23835 , new_n23837 );
xnor g21490 ( n25773 , new_n5771 , new_n14772_1 );
xnor g21491 ( n25784 , new_n17611 , new_n20520 );
xnor g21492 ( n25792 , new_n8357 , new_n8380 );
xnor g21493 ( n25816 , new_n6925 , new_n6958 );
xnor g21494 ( n25826 , new_n6380 , new_n6413 );
xnor g21495 ( n25839 , new_n12285 , new_n12287 );
xnor g21496 ( n25840 , new_n13944 , new_n13984 );
xnor g21497 ( n25873 , new_n8162 , new_n8192 );
xor  g21498 ( n25934 , new_n23556 , new_n23559 );
xnor g21499 ( n25938 , new_n20912 , new_n20925 );
xnor g21500 ( n25985 , new_n21236 , new_n21239 );
xnor g21501 ( n25994 , new_n9033 , new_n13799 );
nor  g21502 ( new_n23851 , new_n18144 , new_n18224 );
nor  g21503 ( new_n23852 , new_n18225 , new_n18284 );
or   g21504 ( n26084 , new_n23851 , new_n23852 );
xnor g21505 ( n26096 , new_n22570 , new_n22583 );
or   g21506 ( new_n23855 , new_n11523 , new_n11585 );
nor  g21507 ( n26111 , new_n11502 , new_n23855 );
xnor g21508 ( n26113 , new_n11549 , new_n11572 );
xor  g21509 ( n26156 , new_n20073 , new_n20076 );
xnor g21510 ( n26159 , new_n17050 , new_n17072 );
xnor g21511 ( n26179 , new_n3674 , new_n3719 );
xor  g21512 ( n26220 , new_n13969 , new_n13970 );
xnor g21513 ( n26229 , new_n22619_1 , new_n22622 );
xnor g21514 ( n26237 , new_n12624 , new_n12655 );
xnor g21515 ( n26250 , new_n15693 , new_n15707 );
xor  g21516 ( n26274 , new_n20962 , new_n20965 );
xnor g21517 ( n26287 , new_n15685 , new_n15711 );
xnor g21518 ( new_n23867 , new_n20438 , new_n21156 );
xnor g21519 ( n26317 , new_n23387 , new_n23867 );
nor  g21520 ( new_n23869 , new_n18533 , new_n18553 );
nor  g21521 ( new_n23870 , new_n18549 , new_n23869 );
nor  g21522 ( new_n23871 , new_n18531 , new_n18552 );
nor  g21523 ( new_n23872 , new_n18548 , new_n23871 );
nor  g21524 ( n26353 , new_n23870 , new_n23872 );
xnor g21525 ( n26375 , new_n20117 , new_n20125 );
nor  g21526 ( new_n23875 , new_n21276_1 , new_n22960 );
nor  g21527 ( new_n23876 , new_n22961 , new_n22969 );
nor  g21528 ( n26396 , new_n23875 , new_n23876 );
xnor g21529 ( n26429 , new_n5435 , new_n22874 );
xnor g21530 ( n26431 , new_n14458 , new_n14473 );
xnor g21531 ( n26439 , new_n7120 , new_n7176 );
xnor g21532 ( n26492 , new_n20365 , new_n20366_1 );
xnor g21533 ( n26515 , new_n10147 , new_n10148 );
xnor g21534 ( n26538 , new_n2510 , new_n2536 );
xnor g21535 ( n26590 , new_n14955 , new_n14968 );
xnor g21536 ( n26598 , new_n16714 , new_n19286 );
xnor g21537 ( new_n23886 , new_n21220 , new_n22928 );
xnor g21538 ( n26605 , new_n22933 , new_n23886 );
xnor g21539 ( new_n23888_1 , new_n22898 , new_n22904 );
xnor g21540 ( n26656 , new_n22901 , new_n23888_1 );
xnor g21541 ( n26674 , new_n11561 , new_n11562 );
xnor g21542 ( n26675 , new_n9549 , new_n9565 );
xnor g21543 ( n26681 , new_n20347 , new_n20376 );
nor  g21544 ( new_n23893 , new_n5498 , new_n5698 );
nor  g21545 ( new_n23894 , new_n23893 , new_n5767 );
nor  g21546 ( new_n23895_1 , new_n5499 , new_n5699 );
nor  g21547 ( new_n23896 , new_n23895_1 , new_n5766 );
nor  g21548 ( n26696 , new_n23894 , new_n23896 );
xnor g21549 ( n26698 , new_n14712 , new_n14730 );
xnor g21550 ( n26707 , new_n5800 , new_n15442 );
xor  g21551 ( n26719 , new_n23327 , new_n23329 );
xnor g21552 ( n26727 , new_n9197 , new_n9209 );
nor  g21553 ( new_n23902 , new_n19127 , new_n21290 );
and  g21554 ( new_n23903_1 , new_n21292 , new_n21295 );
nor  g21555 ( n26729 , new_n23902 , new_n23903_1 );
xor  g21556 ( n26745 , new_n21312 , new_n21315 );
xnor g21557 ( n26775 , new_n7868 , new_n7906 );
xnor g21558 ( n26780 , new_n10483 , new_n10501 );
xor  g21559 ( n26794 , new_n21709 , new_n21716 );
xnor g21560 ( n26795 , new_n3340_1 , new_n3389 );
xnor g21561 ( n26801 , new_n10735 , new_n10773 );
xnor g21562 ( n26815 , new_n11123 , new_n11141 );
xnor g21563 ( n26847 , new_n23018 , new_n23021 );
xnor g21564 ( new_n23913_1 , new_n7361 , new_n18553 );
xnor g21565 ( n26900 , new_n23141 , new_n23913_1 );
xor  g21566 ( n26902 , new_n18692 , new_n18693_1 );
xor  g21567 ( n26905 , new_n17320_1 , new_n17323 );
xnor g21568 ( n26921 , new_n8157 , new_n8194_1 );
xnor g21569 ( n26923 , new_n22045 , new_n22058 );
xnor g21570 ( n26929 , new_n10856 , new_n10857 );
xnor g21571 ( n26930 , new_n12599 , new_n12665_1 );
xnor g21572 ( n26943 , new_n15689 , new_n15709 );
xnor g21573 ( n26970 , new_n14376 , new_n14403 );
xnor g21574 ( n27004 , new_n20854 , new_n20865 );
xnor g21575 ( n27011 , new_n10353 , new_n10407 );
xnor g21576 ( n27019 , new_n19256 , new_n19305 );
xnor g21577 ( n27031 , new_n5001 , new_n5012 );
xnor g21578 ( new_n23927 , new_n20960 , new_n21761 );
xnor g21579 ( n27051 , new_n21800_1 , new_n23927 );
xor  g21580 ( n27072 , new_n17194 , new_n17197 );
xnor g21581 ( n27079 , new_n15276 , new_n15327_1 );
xnor g21582 ( n27096 , new_n4301 , new_n4302 );
xor  g21583 ( n27110 , new_n14138 , new_n14149 );
xnor g21584 ( n27112 , new_n13577 , new_n13580 );
xnor g21585 ( n27130 , new_n21612 , new_n22064 );
xnor g21586 ( n27145 , new_n16056 , new_n16064 );
nor  g21587 ( new_n23936 , new_n14513 , new_n16501 );
and  g21588 ( new_n23937 , new_n21459 , new_n21462 );
nor  g21589 ( n27158 , new_n23936 , new_n23937 );
xnor g21590 ( n27163 , new_n21073 , new_n21076 );
xnor g21591 ( new_n23940 , new_n20872 , new_n23163 );
xnor g21592 ( n27194 , new_n23168 , new_n23940 );
endmodule


