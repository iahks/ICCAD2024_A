// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Sun Aug 18 19:44:02 2024

module top_810026173_826291639_946996917_1246901 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83,
    pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81,
    pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181;
  wire new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n873, new_n875, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1123, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1132, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1157,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1164, new_n1166,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1175,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1371,
    new_n1373, new_n1375, new_n1376, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1412,
    new_n1415, new_n1416, new_n1417, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1426, new_n1427, new_n1433, new_n1434, new_n1435,
    new_n1438, new_n1439, new_n1440, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1447, new_n1448, new_n1449,
    new_n1450, new_n1451, new_n1452, new_n1453, new_n1455, new_n1459,
    new_n1461, new_n1466, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1476, new_n1477, new_n1482, new_n1486, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1497, new_n1498, new_n1499,
    new_n1500, new_n1503, new_n1508, new_n1509, new_n1510, new_n1511,
    new_n1512, new_n1513, new_n1514, new_n1522, new_n1525, new_n1528,
    new_n1536, new_n1539, new_n1541, new_n1542, new_n1548, new_n1550,
    new_n1555, new_n1556, new_n1559, new_n1562, new_n1563, new_n1569,
    new_n1575, new_n1579, new_n1584, new_n1588;
  nand_5 g0000(.A(pi25), .B(pi25), .Y(new_n276));
  nand_5     g0001(.A(pi85), .B(pi03), .Y(new_n277));
  or_6       g0002(.A(pi85), .B(pi03), .Y(new_n278));
  nand_5     g0003(.A(pi47), .B(pi30), .Y(new_n279));
  xor_4      g0004(.A(pi47), .B(pi30), .Y(new_n280));
  nand_5     g0005(.A(pi45), .B(pi19), .Y(new_n281));
  or_6       g0006(.A(pi56), .B(pi17), .Y(new_n282));
  xor_4      g0007(.A(pi56), .B(pi17), .Y(new_n283));
  nand_5     g0008(.A(pi63), .B(pi55), .Y(new_n284));
  nand_5     g0009(.A(new_n284), .B(new_n283), .Y(new_n285));
  nand_5     g0010(.A(new_n285), .B(new_n282), .Y(new_n286));
  nand_5 g0011(.A(new_n286), .B(new_n286), .Y(new_n287));
  xor_4      g0012(.A(pi45), .B(pi19), .Y(new_n288));
  nand_5     g0013(.A(new_n288), .B(new_n287), .Y(new_n289));
  nand_5     g0014(.A(new_n289), .B(new_n281), .Y(new_n290));
  nand_5     g0015(.A(new_n290), .B(new_n280), .Y(new_n291));
  nand_5     g0016(.A(new_n291), .B(new_n279), .Y(new_n292));
  nand_5     g0017(.A(new_n292), .B(new_n278), .Y(new_n293));
  nand_5     g0018(.A(new_n293), .B(new_n277), .Y(new_n294));
  nand_5     g0019(.A(new_n294), .B(pi77), .Y(new_n295));
  xor_4      g0020(.A(new_n295), .B(new_n276), .Y(new_n296));
  nand_5 g0021(.A(new_n296), .B(new_n296), .Y(new_n297));
  nand_5     g0022(.A(pi86), .B(pi60), .Y(new_n298));
  nand_5 g0023(.A(pi60), .B(pi60), .Y(new_n299));
  nand_5     g0024(.A(new_n299), .B(pi39), .Y(new_n300));
  nand_5     g0025(.A(new_n300), .B(new_n298), .Y(new_n301));
  nand_5     g0026(.A(pi60), .B(pi51), .Y(new_n302));
  nand_5     g0027(.A(new_n299), .B(pi06), .Y(new_n303));
  nand_5     g0028(.A(new_n303), .B(new_n302), .Y(new_n304));
  nand_5     g0029(.A(new_n304), .B(pi41), .Y(new_n305));
  xor_4      g0030(.A(new_n304), .B(pi41), .Y(new_n306));
  nand_5     g0031(.A(pi76), .B(pi60), .Y(new_n307));
  nand_5     g0032(.A(new_n299), .B(pi18), .Y(new_n308));
  nand_5     g0033(.A(new_n308), .B(new_n307), .Y(new_n309));
  nand_5     g0034(.A(new_n309), .B(pi79), .Y(new_n310));
  nand_5 g0035(.A(new_n310), .B(new_n310), .Y(new_n311));
  nand_5     g0036(.A(pi60), .B(pi32), .Y(new_n312));
  nand_5     g0037(.A(new_n299), .B(pi59), .Y(new_n313));
  nand_5     g0038(.A(new_n313), .B(new_n312), .Y(new_n314));
  or_6       g0039(.A(new_n314), .B(pi91), .Y(new_n315));
  or_6       g0040(.A(new_n315), .B(new_n311), .Y(new_n316));
  nand_5     g0041(.A(new_n314), .B(pi91), .Y(new_n317));
  or_6       g0042(.A(new_n317), .B(new_n310), .Y(new_n318));
  nand_5     g0043(.A(new_n318), .B(new_n316), .Y(new_n319));
  nand_5     g0044(.A(new_n319), .B(new_n306), .Y(new_n320));
  nand_5     g0045(.A(new_n320), .B(new_n305), .Y(new_n321));
  nand_5 g0046(.A(new_n316), .B(new_n316), .Y(new_n322));
  nand_5     g0047(.A(pi60), .B(pi08), .Y(new_n323));
  nand_5     g0048(.A(pi75), .B(new_n299), .Y(new_n324));
  nand_5     g0049(.A(new_n324), .B(new_n323), .Y(new_n325));
  nand_5 g0050(.A(new_n325), .B(new_n325), .Y(new_n326));
  nand_5     g0051(.A(new_n326), .B(new_n322), .Y(new_n327));
  or_6       g0052(.A(new_n327), .B(new_n321), .Y(new_n328));
  and_6      g0053(.A(new_n328), .B(new_n301), .Y(new_n329));
  nand_5 g0054(.A(new_n301), .B(new_n301), .Y(new_n330));
  nor_5      g0055(.A(new_n326), .B(new_n322), .Y(new_n331));
  nand_5     g0056(.A(new_n331), .B(new_n321), .Y(new_n332));
  nand_5     g0057(.A(new_n332), .B(new_n330), .Y(new_n333));
  nand_5     g0058(.A(pi82), .B(new_n299), .Y(new_n334));
  nand_5 g0059(.A(pi34), .B(pi34), .Y(new_n335));
  nand_5     g0060(.A(pi60), .B(new_n335), .Y(new_n336));
  nand_5     g0061(.A(new_n336), .B(new_n334), .Y(new_n337));
  nand_5 g0062(.A(new_n337), .B(new_n337), .Y(new_n338));
  nand_5     g0063(.A(new_n338), .B(new_n333), .Y(new_n339));
  nor_5      g0064(.A(new_n339), .B(new_n329), .Y(new_n340));
  nand_5 g0065(.A(pi04), .B(pi04), .Y(new_n341));
  nand_5 g0066(.A(pi39), .B(pi39), .Y(new_n342));
  nand_5 g0067(.A(pi82), .B(pi82), .Y(new_n343));
  nand_5     g0068(.A(new_n343), .B(new_n342), .Y(new_n344));
  xor_4      g0069(.A(new_n344), .B(new_n341), .Y(new_n345));
  nand_5     g0070(.A(new_n345), .B(new_n299), .Y(new_n346));
  nand_5 g0071(.A(pi02), .B(pi02), .Y(new_n347));
  nand_5     g0072(.A(pi86), .B(pi34), .Y(new_n348));
  or_6       g0073(.A(new_n348), .B(new_n347), .Y(new_n349));
  nand_5 g0074(.A(new_n349), .B(new_n349), .Y(new_n350));
  nand_5     g0075(.A(new_n348), .B(new_n347), .Y(new_n351));
  nand_5     g0076(.A(new_n351), .B(pi60), .Y(new_n352));
  or_6       g0077(.A(new_n352), .B(new_n350), .Y(new_n353));
  nand_5     g0078(.A(new_n353), .B(new_n346), .Y(new_n354));
  xnor_4     g0079(.A(new_n354), .B(new_n340), .Y(new_n355));
  xor_4      g0080(.A(new_n355), .B(new_n297), .Y(new_n356));
  nand_5 g0081(.A(new_n356), .B(new_n356), .Y(new_n357));
  xor_4      g0082(.A(new_n294), .B(pi77), .Y(new_n358));
  nand_5 g0083(.A(new_n358), .B(new_n358), .Y(new_n359));
  nand_5     g0084(.A(new_n333), .B(new_n328), .Y(new_n360));
  xor_4      g0085(.A(new_n360), .B(new_n337), .Y(new_n361));
  nand_5 g0086(.A(new_n361), .B(new_n361), .Y(new_n362));
  nand_5     g0087(.A(new_n362), .B(new_n359), .Y(new_n363));
  xor_4      g0088(.A(new_n361), .B(new_n359), .Y(new_n364));
  nand_5     g0089(.A(new_n278), .B(new_n277), .Y(new_n365));
  xor_4      g0090(.A(new_n365), .B(new_n292), .Y(new_n366));
  nand_5 g0091(.A(new_n366), .B(new_n366), .Y(new_n367));
  nand_5     g0092(.A(new_n332), .B(new_n328), .Y(new_n368));
  xor_4      g0093(.A(new_n368), .B(new_n301), .Y(new_n369));
  nand_5 g0094(.A(new_n369), .B(new_n369), .Y(new_n370));
  nand_5     g0095(.A(new_n370), .B(new_n367), .Y(new_n371));
  xor_4      g0096(.A(new_n369), .B(new_n366), .Y(new_n372));
  xor_4      g0097(.A(new_n290), .B(new_n280), .Y(new_n373));
  nand_5 g0098(.A(new_n373), .B(new_n373), .Y(new_n374));
  xor_4      g0099(.A(new_n288), .B(new_n286), .Y(new_n375));
  nand_5     g0100(.A(new_n317), .B(new_n315), .Y(new_n376));
  nand_5     g0101(.A(new_n376), .B(new_n311), .Y(new_n377));
  xor_4      g0102(.A(new_n284), .B(new_n283), .Y(new_n378));
  nand_5 g0103(.A(new_n378), .B(new_n378), .Y(new_n379));
  nand_5     g0104(.A(new_n379), .B(new_n376), .Y(new_n380));
  xor_4      g0105(.A(new_n379), .B(new_n376), .Y(new_n381));
  xor_4      g0106(.A(pi63), .B(pi55), .Y(new_n382));
  xor_4      g0107(.A(new_n309), .B(pi79), .Y(new_n383));
  nand_5     g0108(.A(new_n383), .B(new_n382), .Y(new_n384));
  nand_5     g0109(.A(new_n384), .B(new_n310), .Y(new_n385));
  nand_5     g0110(.A(new_n385), .B(new_n381), .Y(new_n386));
  nand_5     g0111(.A(new_n386), .B(new_n380), .Y(new_n387));
  nand_5     g0112(.A(new_n387), .B(new_n377), .Y(new_n388));
  nand_5     g0113(.A(new_n388), .B(new_n375), .Y(new_n389));
  xor_4      g0114(.A(new_n319), .B(new_n306), .Y(new_n390));
  nand_5 g0115(.A(new_n375), .B(new_n375), .Y(new_n391));
  xor_4      g0116(.A(new_n388), .B(new_n391), .Y(new_n392));
  or_6       g0117(.A(new_n392), .B(new_n390), .Y(new_n393));
  nand_5     g0118(.A(new_n393), .B(new_n389), .Y(new_n394));
  nand_5     g0119(.A(new_n394), .B(new_n374), .Y(new_n395));
  xor_4      g0120(.A(new_n394), .B(new_n373), .Y(new_n396));
  xor_4      g0121(.A(new_n326), .B(new_n316), .Y(new_n397));
  xor_4      g0122(.A(new_n397), .B(new_n321), .Y(new_n398));
  or_6       g0123(.A(new_n398), .B(new_n396), .Y(new_n399));
  nand_5     g0124(.A(new_n399), .B(new_n395), .Y(new_n400));
  nand_5 g0125(.A(new_n400), .B(new_n400), .Y(new_n401));
  nand_5     g0126(.A(new_n401), .B(new_n372), .Y(new_n402));
  nand_5     g0127(.A(new_n402), .B(new_n371), .Y(new_n403));
  or_6       g0128(.A(new_n403), .B(new_n364), .Y(new_n404));
  nand_5     g0129(.A(new_n404), .B(new_n363), .Y(new_n405));
  xor_4      g0130(.A(new_n405), .B(new_n357), .Y(po000));
  nand_5 g0131(.A(pi73), .B(pi73), .Y(new_n407));
  nand_5     g0132(.A(new_n407), .B(pi22), .Y(new_n408));
  nand_5     g0133(.A(new_n408), .B(pi76), .Y(new_n409));
  nand_5 g0134(.A(new_n408), .B(new_n408), .Y(new_n410));
  nand_5     g0135(.A(new_n410), .B(pi18), .Y(new_n411));
  nand_5     g0136(.A(new_n411), .B(new_n409), .Y(new_n412));
  xor_4      g0137(.A(new_n412), .B(pi16), .Y(new_n413));
  nand_5     g0138(.A(new_n413), .B(new_n382), .Y(new_n414));
  nand_5     g0139(.A(new_n414), .B(new_n378), .Y(new_n415));
  nand_5     g0140(.A(new_n412), .B(pi16), .Y(new_n416));
  nand_5     g0141(.A(new_n408), .B(pi32), .Y(new_n417));
  nand_5     g0142(.A(new_n410), .B(pi59), .Y(new_n418));
  nand_5     g0143(.A(new_n418), .B(new_n417), .Y(new_n419));
  xor_4      g0144(.A(new_n419), .B(pi57), .Y(new_n420));
  xor_4      g0145(.A(new_n420), .B(new_n416), .Y(new_n421));
  nor_5      g0146(.A(pi63), .B(pi55), .Y(new_n422));
  nand_5 g0147(.A(new_n413), .B(new_n413), .Y(new_n423));
  or_6       g0148(.A(new_n423), .B(new_n422), .Y(new_n424));
  nand_5 g0149(.A(new_n424), .B(new_n424), .Y(new_n425));
  nand_5     g0150(.A(new_n425), .B(new_n283), .Y(new_n426));
  nand_5     g0151(.A(new_n426), .B(new_n421), .Y(new_n427));
  nand_5     g0152(.A(new_n427), .B(new_n415), .Y(new_n428));
  xor_4      g0153(.A(new_n428), .B(new_n375), .Y(new_n429));
  nand_5     g0154(.A(new_n408), .B(pi51), .Y(new_n430));
  nand_5     g0155(.A(new_n410), .B(pi06), .Y(new_n431));
  nand_5     g0156(.A(new_n431), .B(new_n430), .Y(new_n432));
  xor_4      g0157(.A(new_n432), .B(pi07), .Y(new_n433));
  nand_5     g0158(.A(new_n419), .B(pi57), .Y(new_n434));
  nand_5 g0159(.A(new_n416), .B(new_n416), .Y(new_n435));
  nand_5     g0160(.A(new_n420), .B(new_n435), .Y(new_n436));
  nand_5     g0161(.A(new_n436), .B(new_n434), .Y(new_n437));
  xor_4      g0162(.A(new_n437), .B(new_n433), .Y(new_n438));
  xor_4      g0163(.A(new_n438), .B(new_n429), .Y(po001));
  nand_5 g0164(.A(pi84), .B(pi84), .Y(new_n440));
  nand_5     g0165(.A(new_n335), .B(new_n347), .Y(new_n441));
  or_6       g0166(.A(new_n441), .B(new_n407), .Y(new_n442));
  or_6       g0167(.A(new_n442), .B(pi13), .Y(new_n443));
  nand_5 g0168(.A(new_n443), .B(new_n443), .Y(new_n444));
  nand_5     g0169(.A(new_n444), .B(new_n440), .Y(new_n445));
  nand_5 g0170(.A(new_n445), .B(new_n445), .Y(new_n446));
  nand_5 g0171(.A(pi20), .B(pi20), .Y(new_n447));
  nand_5 g0172(.A(pi78), .B(pi78), .Y(new_n448));
  nand_5     g0173(.A(new_n448), .B(new_n341), .Y(new_n449));
  xor_4      g0174(.A(new_n449), .B(new_n447), .Y(new_n450));
  nand_5     g0175(.A(new_n450), .B(new_n410), .Y(new_n451));
  nand_5     g0176(.A(new_n408), .B(pi84), .Y(new_n452));
  or_6       g0177(.A(new_n452), .B(new_n444), .Y(new_n453));
  nand_5     g0178(.A(new_n453), .B(new_n451), .Y(new_n454));
  or_6       g0179(.A(new_n454), .B(new_n446), .Y(new_n455));
  nand_5 g0180(.A(new_n455), .B(new_n455), .Y(new_n456));
  nand_5 g0181(.A(new_n449), .B(new_n449), .Y(new_n457));
  nand_5     g0182(.A(pi78), .B(pi04), .Y(new_n458));
  nand_5     g0183(.A(new_n458), .B(new_n410), .Y(new_n459));
  nor_5      g0184(.A(new_n459), .B(new_n457), .Y(new_n460));
  nand_5 g0185(.A(pi13), .B(pi13), .Y(new_n461));
  nand_5     g0186(.A(new_n408), .B(new_n461), .Y(new_n462));
  nand_5     g0187(.A(new_n462), .B(new_n442), .Y(new_n463));
  or_6       g0188(.A(new_n463), .B(new_n460), .Y(new_n464));
  nand_5     g0189(.A(new_n464), .B(new_n443), .Y(new_n465));
  nand_5 g0190(.A(new_n465), .B(new_n465), .Y(new_n466));
  xor_4      g0191(.A(pi34), .B(pi02), .Y(new_n467));
  nor_5      g0192(.A(new_n467), .B(new_n407), .Y(new_n468));
  nand_5     g0193(.A(new_n410), .B(new_n341), .Y(new_n469));
  or_6       g0194(.A(pi73), .B(pi22), .Y(new_n470));
  or_6       g0195(.A(new_n470), .B(new_n347), .Y(new_n471));
  nand_5     g0196(.A(new_n471), .B(new_n469), .Y(new_n472));
  or_6       g0197(.A(new_n472), .B(new_n468), .Y(new_n473));
  nand_5 g0198(.A(new_n473), .B(new_n473), .Y(new_n474));
  nor_5      g0199(.A(new_n408), .B(pi82), .Y(new_n475));
  or_6       g0200(.A(new_n470), .B(pi34), .Y(new_n476));
  nand_5     g0201(.A(pi73), .B(pi34), .Y(new_n477));
  nand_5     g0202(.A(new_n477), .B(new_n476), .Y(new_n478));
  or_6       g0203(.A(new_n478), .B(new_n475), .Y(new_n479));
  nand_5     g0204(.A(new_n408), .B(pi86), .Y(new_n480));
  nand_5     g0205(.A(new_n410), .B(pi39), .Y(new_n481));
  nand_5     g0206(.A(new_n481), .B(new_n480), .Y(new_n482));
  or_6       g0207(.A(new_n482), .B(pi85), .Y(new_n483));
  xor_4      g0208(.A(new_n482), .B(pi85), .Y(new_n484));
  nand_5     g0209(.A(new_n408), .B(pi08), .Y(new_n485));
  nand_5     g0210(.A(new_n410), .B(pi75), .Y(new_n486));
  nand_5     g0211(.A(new_n486), .B(new_n485), .Y(new_n487));
  nand_5     g0212(.A(new_n487), .B(pi30), .Y(new_n488));
  or_6       g0213(.A(new_n432), .B(pi19), .Y(new_n489));
  or_6       g0214(.A(new_n419), .B(pi56), .Y(new_n490));
  nand_5     g0215(.A(new_n412), .B(pi63), .Y(new_n491));
  nand_5     g0216(.A(new_n419), .B(pi56), .Y(new_n492));
  nand_5     g0217(.A(new_n492), .B(new_n490), .Y(new_n493));
  nand_5 g0218(.A(new_n493), .B(new_n493), .Y(new_n494));
  nand_5     g0219(.A(new_n494), .B(new_n491), .Y(new_n495));
  nand_5     g0220(.A(new_n495), .B(new_n490), .Y(new_n496));
  xor_4      g0221(.A(new_n432), .B(pi19), .Y(new_n497));
  nand_5     g0222(.A(new_n497), .B(new_n496), .Y(new_n498));
  nand_5     g0223(.A(new_n498), .B(new_n489), .Y(new_n499));
  nand_5 g0224(.A(pi30), .B(pi30), .Y(new_n500));
  xor_4      g0225(.A(new_n487), .B(new_n500), .Y(new_n501));
  or_6       g0226(.A(new_n501), .B(new_n499), .Y(new_n502));
  and_6      g0227(.A(new_n502), .B(new_n488), .Y(new_n503));
  nand_5     g0228(.A(new_n503), .B(new_n484), .Y(new_n504));
  nand_5     g0229(.A(new_n504), .B(new_n483), .Y(new_n505));
  nand_5     g0230(.A(new_n505), .B(new_n479), .Y(new_n506));
  or_6       g0231(.A(new_n505), .B(new_n479), .Y(new_n507));
  xor_4      g0232(.A(new_n503), .B(new_n484), .Y(new_n508));
  nand_5 g0233(.A(new_n508), .B(new_n508), .Y(po064));
  xor_4      g0234(.A(new_n497), .B(new_n496), .Y(new_n510));
  or_6       g0235(.A(new_n412), .B(pi63), .Y(new_n511));
  nand_5 g0236(.A(new_n511), .B(new_n511), .Y(new_n512));
  nand_5     g0237(.A(new_n512), .B(new_n490), .Y(new_n513));
  nand_5     g0238(.A(new_n511), .B(new_n492), .Y(new_n514));
  nand_5     g0239(.A(new_n514), .B(new_n513), .Y(new_n515));
  xnor_4     g0240(.A(new_n515), .B(new_n497), .Y(po053));
  nand_5     g0241(.A(po053), .B(new_n510), .Y(new_n517));
  xor_4      g0242(.A(new_n501), .B(new_n499), .Y(po176));
  or_6       g0243(.A(po176), .B(new_n517), .Y(new_n519));
  nand_5     g0244(.A(new_n519), .B(po064), .Y(new_n520));
  nand_5     g0245(.A(new_n520), .B(new_n507), .Y(new_n521));
  nand_5     g0246(.A(new_n521), .B(new_n506), .Y(new_n522));
  or_6       g0247(.A(new_n522), .B(new_n474), .Y(new_n523));
  or_6       g0248(.A(new_n523), .B(new_n466), .Y(new_n524));
  xor_4      g0249(.A(new_n524), .B(new_n456), .Y(po002));
  xor_4      g0250(.A(new_n383), .B(new_n382), .Y(po003));
  nand_5 g0251(.A(pi21), .B(pi21), .Y(new_n527));
  nand_5     g0252(.A(pi14), .B(pi08), .Y(new_n528));
  nand_5 g0253(.A(pi14), .B(pi14), .Y(new_n529));
  nand_5     g0254(.A(pi75), .B(new_n529), .Y(new_n530));
  nand_5     g0255(.A(new_n530), .B(new_n528), .Y(new_n531));
  or_6       g0256(.A(new_n531), .B(pi12), .Y(new_n532));
  xor_4      g0257(.A(new_n531), .B(pi12), .Y(new_n533));
  nand_5 g0258(.A(new_n533), .B(new_n533), .Y(new_n534));
  nand_5     g0259(.A(pi32), .B(pi14), .Y(new_n535));
  nand_5     g0260(.A(pi59), .B(new_n529), .Y(new_n536));
  nand_5     g0261(.A(new_n536), .B(new_n535), .Y(new_n537));
  nand_5     g0262(.A(new_n537), .B(pi28), .Y(new_n538));
  nand_5 g0263(.A(new_n538), .B(new_n538), .Y(new_n539));
  nand_5     g0264(.A(pi51), .B(pi14), .Y(new_n540));
  nand_5     g0265(.A(new_n529), .B(pi06), .Y(new_n541));
  nand_5     g0266(.A(new_n541), .B(new_n540), .Y(new_n542));
  or_6       g0267(.A(new_n542), .B(pi26), .Y(new_n543));
  or_6       g0268(.A(new_n543), .B(new_n539), .Y(new_n544));
  nand_5     g0269(.A(new_n542), .B(pi26), .Y(new_n545));
  or_6       g0270(.A(new_n545), .B(new_n538), .Y(new_n546));
  nand_5     g0271(.A(new_n546), .B(new_n544), .Y(new_n547));
  or_6       g0272(.A(new_n547), .B(new_n534), .Y(new_n548));
  nand_5     g0273(.A(new_n548), .B(new_n532), .Y(new_n549));
  nand_5     g0274(.A(pi86), .B(pi14), .Y(new_n550));
  nand_5     g0275(.A(pi39), .B(new_n529), .Y(new_n551));
  nand_5     g0276(.A(new_n551), .B(new_n550), .Y(new_n552));
  nand_5     g0277(.A(new_n552), .B(new_n549), .Y(new_n553));
  nand_5 g0278(.A(new_n544), .B(new_n544), .Y(new_n554));
  nand_5     g0279(.A(new_n554), .B(new_n532), .Y(new_n555));
  nand_5 g0280(.A(new_n552), .B(new_n552), .Y(new_n556));
  nand_5     g0281(.A(new_n556), .B(new_n544), .Y(new_n557));
  nand_5     g0282(.A(new_n557), .B(new_n555), .Y(new_n558));
  nand_5 g0283(.A(new_n558), .B(new_n558), .Y(new_n559));
  nand_5     g0284(.A(new_n559), .B(new_n553), .Y(new_n560));
  nand_5 g0285(.A(new_n560), .B(new_n560), .Y(new_n561));
  xor_4      g0286(.A(pi86), .B(pi34), .Y(new_n562));
  or_6       g0287(.A(new_n562), .B(new_n529), .Y(new_n563));
  nand_5     g0288(.A(pi82), .B(pi39), .Y(new_n564));
  nand_5     g0289(.A(new_n344), .B(new_n529), .Y(new_n565));
  nand_5 g0290(.A(new_n565), .B(new_n565), .Y(new_n566));
  nand_5     g0291(.A(new_n566), .B(new_n564), .Y(new_n567));
  nand_5     g0292(.A(new_n567), .B(new_n563), .Y(new_n568));
  nand_5     g0293(.A(new_n568), .B(new_n561), .Y(new_n569));
  nand_5     g0294(.A(pi14), .B(pi02), .Y(new_n570));
  nand_5 g0295(.A(new_n570), .B(new_n570), .Y(new_n571));
  nand_5     g0296(.A(new_n529), .B(pi04), .Y(new_n572));
  or_6       g0297(.A(new_n572), .B(new_n343), .Y(new_n573));
  nand_5     g0298(.A(new_n343), .B(new_n529), .Y(new_n574));
  nand_5 g0299(.A(new_n574), .B(new_n574), .Y(new_n575));
  nand_5     g0300(.A(new_n575), .B(new_n341), .Y(new_n576));
  nand_5     g0301(.A(new_n576), .B(new_n573), .Y(new_n577));
  or_6       g0302(.A(new_n577), .B(new_n571), .Y(new_n578));
  xor_4      g0303(.A(new_n578), .B(new_n569), .Y(new_n579));
  or_6       g0304(.A(new_n579), .B(new_n527), .Y(new_n580));
  nand_5     g0305(.A(pi34), .B(pi14), .Y(new_n581));
  nand_5     g0306(.A(new_n581), .B(new_n574), .Y(new_n582));
  xor_4      g0307(.A(new_n582), .B(new_n560), .Y(new_n583));
  nand_5 g0308(.A(new_n583), .B(new_n583), .Y(new_n584));
  nand_5     g0309(.A(new_n584), .B(pi69), .Y(new_n585));
  or_6       g0310(.A(pi87), .B(pi85), .Y(new_n586));
  nand_5     g0311(.A(pi62), .B(pi30), .Y(new_n587));
  xor_4      g0312(.A(pi62), .B(new_n500), .Y(new_n588));
  or_6       g0313(.A(pi71), .B(pi19), .Y(new_n589));
  nand_5     g0314(.A(pi71), .B(pi19), .Y(new_n590));
  or_6       g0315(.A(pi56), .B(pi43), .Y(new_n591));
  nand_5     g0316(.A(pi56), .B(pi43), .Y(new_n592));
  nand_5     g0317(.A(pi63), .B(pi40), .Y(new_n593));
  nand_5     g0318(.A(new_n593), .B(new_n592), .Y(new_n594));
  nand_5     g0319(.A(new_n594), .B(new_n591), .Y(new_n595));
  nand_5     g0320(.A(new_n595), .B(new_n590), .Y(new_n596));
  nand_5     g0321(.A(new_n596), .B(new_n589), .Y(new_n597));
  or_6       g0322(.A(new_n597), .B(new_n588), .Y(new_n598));
  nand_5     g0323(.A(new_n598), .B(new_n587), .Y(new_n599));
  nand_5     g0324(.A(new_n599), .B(new_n586), .Y(new_n600));
  nand_5     g0325(.A(pi87), .B(pi85), .Y(new_n601));
  nand_5     g0326(.A(new_n601), .B(new_n600), .Y(new_n602));
  xor_4      g0327(.A(new_n583), .B(pi69), .Y(new_n603));
  xor_4      g0328(.A(new_n603), .B(new_n602), .Y(new_n604));
  nand_5     g0329(.A(new_n601), .B(new_n586), .Y(new_n605));
  xor_4      g0330(.A(new_n605), .B(new_n599), .Y(new_n606));
  nand_5     g0331(.A(new_n549), .B(new_n544), .Y(new_n607));
  nand_5     g0332(.A(new_n607), .B(new_n555), .Y(new_n608));
  xor_4      g0333(.A(new_n608), .B(new_n552), .Y(new_n609));
  or_6       g0334(.A(new_n609), .B(new_n606), .Y(new_n610));
  xor_4      g0335(.A(new_n609), .B(new_n606), .Y(new_n611));
  nand_5 g0336(.A(new_n611), .B(new_n611), .Y(new_n612));
  xor_4      g0337(.A(new_n547), .B(new_n534), .Y(new_n613));
  nand_5 g0338(.A(new_n613), .B(new_n613), .Y(new_n614));
  xor_4      g0339(.A(new_n597), .B(new_n588), .Y(new_n615));
  or_6       g0340(.A(new_n615), .B(new_n614), .Y(new_n616));
  xor_4      g0341(.A(new_n615), .B(new_n613), .Y(new_n617));
  nand_5     g0342(.A(new_n545), .B(new_n543), .Y(new_n618));
  xor_4      g0343(.A(new_n618), .B(new_n539), .Y(new_n619));
  nand_5     g0344(.A(new_n589), .B(new_n590), .Y(new_n620));
  xor_4      g0345(.A(new_n620), .B(new_n595), .Y(new_n621));
  nand_5     g0346(.A(new_n621), .B(new_n619), .Y(new_n622));
  or_6       g0347(.A(new_n621), .B(new_n619), .Y(new_n623));
  nand_5 g0348(.A(new_n537), .B(new_n537), .Y(new_n624));
  xor_4      g0349(.A(new_n624), .B(pi28), .Y(new_n625));
  nand_5     g0350(.A(new_n592), .B(new_n591), .Y(new_n626));
  xor_4      g0351(.A(new_n626), .B(new_n593), .Y(new_n627));
  nand_5 g0352(.A(new_n627), .B(new_n627), .Y(new_n628));
  or_6       g0353(.A(new_n628), .B(new_n625), .Y(new_n629));
  nand_5     g0354(.A(pi76), .B(pi14), .Y(new_n630));
  nand_5     g0355(.A(pi18), .B(new_n529), .Y(new_n631));
  nand_5     g0356(.A(new_n631), .B(new_n630), .Y(new_n632));
  nand_5     g0357(.A(new_n632), .B(pi48), .Y(new_n633));
  nor_5      g0358(.A(new_n632), .B(pi48), .Y(new_n634));
  nand_5 g0359(.A(pi63), .B(pi63), .Y(new_n635));
  nand_5 g0360(.A(new_n632), .B(new_n632), .Y(new_n636));
  nand_5     g0361(.A(new_n636), .B(new_n635), .Y(new_n637));
  nand_5     g0362(.A(new_n632), .B(pi63), .Y(new_n638));
  nand_5     g0363(.A(new_n638), .B(new_n637), .Y(po125));
  nand_5 g0364(.A(po125), .B(po125), .Y(po058));
  xor_4      g0365(.A(pi48), .B(pi40), .Y(new_n641));
  xor_4      g0366(.A(new_n641), .B(po058), .Y(po037));
  or_6       g0367(.A(po037), .B(new_n634), .Y(new_n643));
  nand_5     g0368(.A(new_n643), .B(new_n633), .Y(new_n644));
  xor_4      g0369(.A(new_n628), .B(new_n625), .Y(new_n645));
  nand_5     g0370(.A(new_n645), .B(new_n644), .Y(new_n646));
  nand_5     g0371(.A(new_n646), .B(new_n629), .Y(new_n647));
  nand_5     g0372(.A(new_n647), .B(new_n623), .Y(new_n648));
  nand_5     g0373(.A(new_n648), .B(new_n622), .Y(new_n649));
  or_6       g0374(.A(new_n649), .B(new_n617), .Y(new_n650));
  nand_5     g0375(.A(new_n650), .B(new_n616), .Y(new_n651));
  or_6       g0376(.A(new_n651), .B(new_n612), .Y(new_n652));
  nand_5     g0377(.A(new_n652), .B(new_n610), .Y(new_n653));
  nand_5 g0378(.A(new_n653), .B(new_n653), .Y(new_n654));
  or_6       g0379(.A(new_n654), .B(new_n604), .Y(new_n655));
  or_6       g0380(.A(new_n655), .B(new_n585), .Y(new_n656));
  or_6       g0381(.A(new_n656), .B(new_n580), .Y(new_n657));
  or_6       g0382(.A(new_n584), .B(pi69), .Y(new_n658));
  or_6       g0383(.A(new_n603), .B(new_n602), .Y(new_n659));
  nand_5     g0384(.A(new_n659), .B(new_n658), .Y(new_n660));
  nand_5     g0385(.A(new_n660), .B(new_n655), .Y(new_n661));
  nand_5     g0386(.A(new_n661), .B(new_n656), .Y(new_n662));
  xor_4      g0387(.A(new_n579), .B(new_n527), .Y(new_n663));
  or_6       g0388(.A(new_n663), .B(new_n662), .Y(new_n664));
  nand_5     g0389(.A(new_n664), .B(new_n661), .Y(new_n665));
  nand_5     g0390(.A(new_n665), .B(new_n580), .Y(new_n666));
  nand_5     g0391(.A(new_n666), .B(new_n657), .Y(new_n667));
  nand_5 g0392(.A(pi81), .B(pi81), .Y(new_n668));
  nand_5     g0393(.A(new_n467), .B(pi14), .Y(new_n669));
  nand_5     g0394(.A(new_n669), .B(new_n572), .Y(new_n670));
  or_6       g0395(.A(new_n670), .B(new_n569), .Y(new_n671));
  nand_5     g0396(.A(new_n448), .B(new_n529), .Y(new_n672));
  nand_5     g0397(.A(new_n672), .B(new_n576), .Y(new_n673));
  nand_5     g0398(.A(new_n457), .B(new_n343), .Y(new_n674));
  nand_5     g0399(.A(new_n674), .B(new_n673), .Y(new_n675));
  nand_5     g0400(.A(pi14), .B(new_n461), .Y(new_n676));
  nand_5     g0401(.A(new_n676), .B(new_n675), .Y(new_n677));
  nand_5 g0402(.A(new_n677), .B(new_n677), .Y(new_n678));
  xor_4      g0403(.A(new_n678), .B(new_n671), .Y(new_n679));
  xor_4      g0404(.A(new_n679), .B(new_n668), .Y(new_n680));
  xnor_4     g0405(.A(new_n680), .B(new_n667), .Y(po004));
  nand_5 g0406(.A(new_n582), .B(new_n582), .Y(new_n682));
  xor_4      g0407(.A(new_n677), .B(new_n682), .Y(new_n683));
  or_6       g0408(.A(new_n683), .B(new_n671), .Y(new_n684));
  nand_5     g0409(.A(new_n457), .B(new_n447), .Y(new_n685));
  nand_5 g0410(.A(new_n685), .B(new_n685), .Y(new_n686));
  nand_5     g0411(.A(new_n575), .B(new_n686), .Y(new_n687));
  nand_5 g0412(.A(new_n687), .B(new_n687), .Y(new_n688));
  nor_5      g0413(.A(new_n447), .B(pi14), .Y(new_n689));
  nand_5     g0414(.A(new_n689), .B(new_n674), .Y(new_n690));
  nand_5     g0415(.A(pi84), .B(pi14), .Y(new_n691));
  nand_5     g0416(.A(new_n691), .B(new_n690), .Y(new_n692));
  or_6       g0417(.A(new_n692), .B(new_n688), .Y(new_n693));
  nand_5 g0418(.A(new_n693), .B(new_n693), .Y(new_n694));
  nand_5     g0419(.A(new_n694), .B(new_n682), .Y(new_n695));
  or_6       g0420(.A(new_n695), .B(new_n684), .Y(new_n696));
  nand_5     g0421(.A(new_n678), .B(new_n582), .Y(new_n697));
  or_6       g0422(.A(new_n694), .B(new_n697), .Y(new_n698));
  or_6       g0423(.A(new_n698), .B(new_n671), .Y(new_n699));
  nand_5     g0424(.A(new_n699), .B(new_n696), .Y(new_n700));
  nand_5 g0425(.A(pi66), .B(pi66), .Y(new_n701));
  nand_5     g0426(.A(new_n687), .B(new_n529), .Y(new_n702));
  nor_5      g0427(.A(new_n702), .B(new_n701), .Y(new_n703));
  nand_5     g0428(.A(new_n688), .B(new_n701), .Y(new_n704));
  nand_5     g0429(.A(pi14), .B(pi09), .Y(new_n705));
  nand_5     g0430(.A(new_n705), .B(new_n704), .Y(new_n706));
  or_6       g0431(.A(new_n706), .B(new_n703), .Y(new_n707));
  nand_5 g0432(.A(new_n707), .B(new_n707), .Y(new_n708));
  xor_4      g0433(.A(new_n708), .B(new_n700), .Y(new_n709));
  nand_5 g0434(.A(new_n709), .B(new_n709), .Y(new_n710));
  nand_5 g0435(.A(pi35), .B(pi35), .Y(new_n711));
  xor_4      g0436(.A(new_n693), .B(new_n684), .Y(new_n712));
  xor_4      g0437(.A(new_n712), .B(new_n711), .Y(new_n713));
  or_6       g0438(.A(new_n679), .B(new_n668), .Y(new_n714));
  or_6       g0439(.A(new_n714), .B(new_n657), .Y(new_n715));
  or_6       g0440(.A(new_n680), .B(new_n667), .Y(new_n716));
  nand_5     g0441(.A(new_n716), .B(new_n666), .Y(new_n717));
  nand_5     g0442(.A(new_n717), .B(new_n714), .Y(new_n718));
  nand_5     g0443(.A(new_n718), .B(new_n715), .Y(new_n719));
  nand_5 g0444(.A(new_n719), .B(new_n719), .Y(new_n720));
  nand_5     g0445(.A(new_n720), .B(new_n713), .Y(new_n721));
  or_6       g0446(.A(new_n712), .B(new_n711), .Y(new_n722));
  and_6      g0447(.A(new_n715), .B(new_n722), .Y(new_n723));
  nand_5     g0448(.A(new_n723), .B(new_n721), .Y(new_n724));
  nand_5     g0449(.A(new_n724), .B(new_n710), .Y(new_n725));
  or_6       g0450(.A(new_n715), .B(new_n722), .Y(new_n726));
  nand_5     g0451(.A(new_n726), .B(new_n709), .Y(new_n727));
  nand_5     g0452(.A(new_n727), .B(new_n725), .Y(new_n728));
  nand_5     g0453(.A(new_n708), .B(new_n699), .Y(new_n729));
  nand_5     g0454(.A(new_n729), .B(new_n696), .Y(new_n730));
  nand_5     g0455(.A(new_n686), .B(new_n701), .Y(new_n731));
  nand_5     g0456(.A(new_n731), .B(pi74), .Y(new_n732));
  nand_5     g0457(.A(new_n732), .B(new_n529), .Y(new_n733));
  nand_5 g0458(.A(pi31), .B(pi31), .Y(new_n734));
  nand_5     g0459(.A(new_n734), .B(pi14), .Y(new_n735));
  nand_5     g0460(.A(new_n735), .B(new_n733), .Y(new_n736));
  nand_5 g0461(.A(new_n736), .B(new_n736), .Y(new_n737));
  nand_5 g0462(.A(pi74), .B(pi74), .Y(new_n738));
  nand_5     g0463(.A(new_n701), .B(new_n447), .Y(new_n739));
  nand_5 g0464(.A(new_n739), .B(new_n739), .Y(new_n740));
  nand_5     g0465(.A(new_n740), .B(new_n738), .Y(new_n741));
  nand_5 g0466(.A(new_n741), .B(new_n741), .Y(new_n742));
  nand_5     g0467(.A(new_n742), .B(new_n688), .Y(new_n743));
  or_6       g0468(.A(new_n702), .B(new_n738), .Y(new_n744));
  nand_5     g0469(.A(new_n744), .B(new_n743), .Y(new_n745));
  or_6       g0470(.A(new_n745), .B(new_n737), .Y(new_n746));
  xor_4      g0471(.A(new_n746), .B(new_n730), .Y(new_n747));
  xor_4      g0472(.A(new_n747), .B(new_n728), .Y(po005));
  nand_5 g0473(.A(new_n398), .B(new_n398), .Y(new_n749));
  or_6       g0474(.A(pi37), .B(pi19), .Y(new_n750));
  xor_4      g0475(.A(pi37), .B(pi19), .Y(new_n751));
  nand_5     g0476(.A(pi56), .B(pi36), .Y(new_n752));
  nand_5     g0477(.A(new_n752), .B(new_n751), .Y(new_n753));
  nand_5     g0478(.A(new_n753), .B(new_n750), .Y(new_n754));
  xor_4      g0479(.A(pi54), .B(pi30), .Y(new_n755));
  xor_4      g0480(.A(new_n755), .B(new_n754), .Y(new_n756));
  nand_5     g0481(.A(new_n756), .B(new_n749), .Y(new_n757));
  xor_4      g0482(.A(new_n756), .B(new_n749), .Y(new_n758));
  or_6       g0483(.A(pi56), .B(pi36), .Y(new_n759));
  nand_5     g0484(.A(new_n759), .B(new_n752), .Y(new_n760));
  xor_4      g0485(.A(new_n376), .B(new_n311), .Y(new_n761));
  nand_5     g0486(.A(pi92), .B(pi63), .Y(new_n762));
  xor_4      g0487(.A(pi92), .B(pi63), .Y(new_n763));
  nand_5     g0488(.A(new_n763), .B(new_n383), .Y(new_n764));
  nand_5     g0489(.A(new_n764), .B(new_n762), .Y(new_n765));
  xor_4      g0490(.A(new_n765), .B(new_n761), .Y(new_n766));
  or_6       g0491(.A(new_n766), .B(new_n760), .Y(new_n767));
  nand_5     g0492(.A(new_n767), .B(new_n759), .Y(new_n768));
  xor_4      g0493(.A(new_n768), .B(new_n751), .Y(new_n769));
  nand_5 g0494(.A(new_n390), .B(new_n390), .Y(new_n770));
  nand_5     g0495(.A(new_n765), .B(new_n761), .Y(new_n771));
  nand_5     g0496(.A(new_n771), .B(new_n770), .Y(new_n772));
  or_6       g0497(.A(new_n772), .B(new_n769), .Y(new_n773));
  nor_5      g0498(.A(new_n768), .B(new_n751), .Y(new_n774));
  or_6       g0499(.A(new_n771), .B(new_n770), .Y(new_n775));
  nand_5     g0500(.A(new_n775), .B(new_n753), .Y(new_n776));
  or_6       g0501(.A(new_n776), .B(new_n774), .Y(new_n777));
  nand_5     g0502(.A(new_n777), .B(new_n773), .Y(new_n778));
  nand_5     g0503(.A(new_n778), .B(new_n758), .Y(new_n779));
  nand_5     g0504(.A(new_n779), .B(new_n757), .Y(new_n780));
  xor_4      g0505(.A(pi85), .B(pi27), .Y(new_n781));
  nand_5     g0506(.A(pi54), .B(pi30), .Y(new_n782));
  nand_5 g0507(.A(new_n754), .B(new_n754), .Y(new_n783));
  nand_5     g0508(.A(new_n755), .B(new_n783), .Y(new_n784));
  nand_5     g0509(.A(new_n784), .B(new_n782), .Y(new_n785));
  xor_4      g0510(.A(new_n785), .B(new_n781), .Y(new_n786));
  xor_4      g0511(.A(new_n786), .B(new_n370), .Y(new_n787));
  xnor_4     g0512(.A(new_n787), .B(new_n780), .Y(po006));
  nand_5 g0513(.A(pi09), .B(pi09), .Y(new_n789));
  nand_5     g0514(.A(new_n446), .B(new_n789), .Y(new_n790));
  or_6       g0515(.A(new_n790), .B(pi31), .Y(new_n791));
  or_6       g0516(.A(new_n469), .B(pi78), .Y(new_n792));
  or_6       g0517(.A(new_n792), .B(new_n741), .Y(new_n793));
  nand_5     g0518(.A(new_n793), .B(new_n791), .Y(new_n794));
  nand_5 g0519(.A(new_n794), .B(new_n794), .Y(new_n795));
  and_6      g0520(.A(new_n732), .B(new_n410), .Y(new_n796));
  nand_5     g0521(.A(new_n408), .B(new_n734), .Y(new_n797));
  nand_5     g0522(.A(new_n797), .B(new_n790), .Y(new_n798));
  or_6       g0523(.A(new_n798), .B(new_n796), .Y(new_n799));
  nand_5     g0524(.A(new_n799), .B(new_n795), .Y(new_n800));
  nand_5 g0525(.A(new_n800), .B(new_n800), .Y(new_n801));
  or_6       g0526(.A(new_n524), .B(new_n456), .Y(new_n802));
  nand_5     g0527(.A(new_n408), .B(new_n789), .Y(new_n803));
  nand_5     g0528(.A(new_n803), .B(new_n445), .Y(new_n804));
  nand_5     g0529(.A(new_n804), .B(new_n790), .Y(new_n805));
  nor_5      g0530(.A(new_n686), .B(new_n701), .Y(new_n806));
  nand_5     g0531(.A(new_n731), .B(new_n410), .Y(new_n807));
  or_6       g0532(.A(new_n807), .B(new_n806), .Y(new_n808));
  nand_5     g0533(.A(new_n808), .B(new_n805), .Y(new_n809));
  or_6       g0534(.A(new_n809), .B(new_n802), .Y(new_n810));
  xor_4      g0535(.A(new_n810), .B(new_n801), .Y(po007));
  xor_4      g0536(.A(new_n522), .B(new_n474), .Y(po008));
  xor_4      g0537(.A(new_n651), .B(new_n612), .Y(po009));
  nand_5 g0538(.A(new_n578), .B(new_n578), .Y(new_n814));
  nand_5     g0539(.A(new_n552), .B(pi85), .Y(new_n815));
  xor_4      g0540(.A(new_n552), .B(pi85), .Y(new_n816));
  nand_5 g0541(.A(new_n816), .B(new_n816), .Y(new_n817));
  nand_5 g0542(.A(new_n531), .B(new_n531), .Y(new_n818));
  nor_5      g0543(.A(new_n818), .B(new_n500), .Y(new_n819));
  or_6       g0544(.A(new_n542), .B(pi19), .Y(new_n820));
  xor_4      g0545(.A(new_n542), .B(pi19), .Y(new_n821));
  or_6       g0546(.A(new_n537), .B(pi56), .Y(new_n822));
  nand_5     g0547(.A(new_n537), .B(pi56), .Y(new_n823));
  nand_5     g0548(.A(new_n823), .B(new_n638), .Y(new_n824));
  nand_5     g0549(.A(new_n824), .B(new_n822), .Y(new_n825));
  nand_5     g0550(.A(new_n825), .B(new_n821), .Y(new_n826));
  nand_5     g0551(.A(new_n826), .B(new_n820), .Y(new_n827));
  xor_4      g0552(.A(new_n531), .B(new_n500), .Y(new_n828));
  nor_5      g0553(.A(new_n828), .B(new_n827), .Y(new_n829));
  nor_5      g0554(.A(new_n829), .B(new_n819), .Y(new_n830));
  or_6       g0555(.A(new_n830), .B(new_n817), .Y(new_n831));
  nand_5     g0556(.A(new_n831), .B(new_n815), .Y(new_n832));
  nand_5     g0557(.A(new_n832), .B(new_n582), .Y(new_n833));
  xor_4      g0558(.A(new_n833), .B(new_n814), .Y(po010));
  or_6       g0559(.A(new_n507), .B(new_n474), .Y(new_n835));
  or_6       g0560(.A(new_n835), .B(new_n466), .Y(new_n836));
  or_6       g0561(.A(new_n836), .B(new_n456), .Y(new_n837));
  or_6       g0562(.A(new_n837), .B(new_n809), .Y(new_n838));
  xor_4      g0563(.A(new_n838), .B(new_n801), .Y(po011));
  xor_4      g0564(.A(new_n382), .B(pi18), .Y(po012));
  xor_4      g0565(.A(new_n358), .B(new_n343), .Y(new_n841));
  nand_5     g0566(.A(new_n366), .B(new_n342), .Y(new_n842));
  nand_5     g0567(.A(new_n367), .B(pi39), .Y(new_n843));
  or_6       g0568(.A(new_n373), .B(pi75), .Y(new_n844));
  nand_5     g0569(.A(new_n373), .B(pi75), .Y(new_n845));
  nand_5     g0570(.A(new_n391), .B(pi06), .Y(new_n846));
  nand_5     g0571(.A(new_n382), .B(pi18), .Y(new_n847));
  nand_5 g0572(.A(new_n847), .B(new_n847), .Y(new_n848));
  nand_5     g0573(.A(new_n848), .B(pi59), .Y(new_n849));
  xor_4      g0574(.A(new_n847), .B(pi59), .Y(new_n850));
  or_6       g0575(.A(new_n850), .B(new_n378), .Y(new_n851));
  nand_5     g0576(.A(new_n851), .B(new_n849), .Y(new_n852));
  or_6       g0577(.A(new_n391), .B(pi06), .Y(new_n853));
  nand_5     g0578(.A(new_n853), .B(new_n852), .Y(new_n854));
  nand_5     g0579(.A(new_n854), .B(new_n846), .Y(new_n855));
  nand_5 g0580(.A(new_n855), .B(new_n855), .Y(new_n856));
  nand_5     g0581(.A(new_n856), .B(new_n845), .Y(new_n857));
  nand_5     g0582(.A(new_n857), .B(new_n844), .Y(new_n858));
  nand_5     g0583(.A(new_n858), .B(new_n843), .Y(new_n859));
  nand_5     g0584(.A(new_n859), .B(new_n842), .Y(new_n860));
  xor_4      g0585(.A(new_n860), .B(new_n841), .Y(new_n861));
  nand_5     g0586(.A(new_n853), .B(new_n846), .Y(new_n862));
  xor_4      g0587(.A(new_n862), .B(new_n852), .Y(po047));
  nor_5      g0588(.A(po047), .B(new_n861), .Y(new_n864));
  nand_5 g0589(.A(po047), .B(po047), .Y(po145));
  or_6       g0590(.A(new_n856), .B(new_n845), .Y(new_n866));
  or_6       g0591(.A(new_n855), .B(new_n844), .Y(new_n867));
  nand_5     g0592(.A(new_n867), .B(new_n858), .Y(new_n868));
  and_6      g0593(.A(new_n868), .B(new_n866), .Y(po162));
  nand_5     g0594(.A(new_n842), .B(new_n843), .Y(new_n870));
  nand_5     g0595(.A(new_n867), .B(new_n866), .Y(new_n871));
  xnor_4     g0596(.A(new_n871), .B(new_n870), .Y(po147));
  nand_5     g0597(.A(po147), .B(po162), .Y(new_n873));
  xnor_4     g0598(.A(new_n873), .B(new_n861), .Y(po099));
  nor_5      g0599(.A(po099), .B(po145), .Y(new_n875));
  nor_5      g0600(.A(new_n875), .B(new_n864), .Y(po013));
  xor_4      g0601(.A(new_n392), .B(new_n770), .Y(po014));
  nand_5     g0602(.A(pi72), .B(pi30), .Y(new_n878));
  nand_5     g0603(.A(pi29), .B(pi19), .Y(new_n879));
  nand_5     g0604(.A(pi56), .B(pi23), .Y(new_n880));
  xor_4      g0605(.A(pi56), .B(pi23), .Y(new_n881));
  and_6      g0606(.A(pi63), .B(pi10), .Y(new_n882));
  nand_5     g0607(.A(new_n882), .B(new_n881), .Y(new_n883));
  and_6      g0608(.A(new_n883), .B(new_n880), .Y(new_n884));
  xnor_4     g0609(.A(pi29), .B(pi19), .Y(new_n885));
  or_6       g0610(.A(new_n885), .B(new_n884), .Y(new_n886));
  nand_5     g0611(.A(new_n886), .B(new_n879), .Y(new_n887));
  xor_4      g0612(.A(pi72), .B(new_n500), .Y(new_n888));
  nand_5 g0613(.A(new_n888), .B(new_n888), .Y(new_n889));
  nand_5     g0614(.A(new_n889), .B(new_n887), .Y(new_n890));
  nand_5     g0615(.A(new_n890), .B(new_n878), .Y(new_n891));
  nand_5 g0616(.A(new_n891), .B(new_n891), .Y(new_n892));
  or_6       g0617(.A(new_n542), .B(pi11), .Y(new_n893));
  nand_5     g0618(.A(new_n537), .B(pi88), .Y(new_n894));
  nand_5 g0619(.A(new_n894), .B(new_n894), .Y(new_n895));
  xnor_4     g0620(.A(new_n542), .B(pi11), .Y(new_n896));
  or_6       g0621(.A(new_n896), .B(new_n895), .Y(new_n897));
  nand_5     g0622(.A(new_n897), .B(new_n893), .Y(new_n898));
  or_6       g0623(.A(new_n898), .B(new_n818), .Y(new_n899));
  xor_4      g0624(.A(new_n899), .B(new_n556), .Y(new_n900));
  nand_5     g0625(.A(pi85), .B(pi24), .Y(new_n901));
  or_6       g0626(.A(pi85), .B(pi24), .Y(new_n902));
  nand_5     g0627(.A(new_n902), .B(new_n901), .Y(new_n903));
  xor_4      g0628(.A(new_n903), .B(new_n900), .Y(new_n904));
  or_6       g0629(.A(new_n904), .B(new_n892), .Y(new_n905));
  xor_4      g0630(.A(new_n904), .B(new_n891), .Y(new_n906));
  xor_4      g0631(.A(new_n898), .B(new_n818), .Y(new_n907));
  xor_4      g0632(.A(new_n889), .B(new_n887), .Y(new_n908));
  or_6       g0633(.A(new_n908), .B(new_n907), .Y(new_n909));
  xor_4      g0634(.A(new_n908), .B(new_n907), .Y(new_n910));
  xor_4      g0635(.A(new_n896), .B(new_n894), .Y(new_n911));
  xor_4      g0636(.A(new_n885), .B(new_n884), .Y(new_n912));
  or_6       g0637(.A(new_n912), .B(new_n911), .Y(new_n913));
  xnor_4     g0638(.A(new_n912), .B(new_n911), .Y(new_n914));
  xor_4      g0639(.A(new_n537), .B(pi88), .Y(new_n915));
  nand_5 g0640(.A(new_n915), .B(new_n915), .Y(new_n916));
  nand_5     g0641(.A(pi33), .B(pi10), .Y(new_n917));
  or_6       g0642(.A(new_n917), .B(new_n638), .Y(new_n918));
  nand_5 g0643(.A(pi33), .B(pi33), .Y(new_n919));
  xor_4      g0644(.A(new_n919), .B(pi10), .Y(new_n920));
  nor_5      g0645(.A(new_n920), .B(po125), .Y(new_n921));
  nand_5     g0646(.A(new_n917), .B(new_n638), .Y(new_n922));
  or_6       g0647(.A(new_n922), .B(new_n921), .Y(new_n923));
  nand_5     g0648(.A(new_n923), .B(new_n918), .Y(new_n924));
  xor_4      g0649(.A(new_n924), .B(new_n881), .Y(new_n925));
  or_6       g0650(.A(new_n925), .B(new_n916), .Y(new_n926));
  nor_5      g0651(.A(new_n924), .B(new_n881), .Y(new_n927));
  nand_5     g0652(.A(new_n923), .B(new_n883), .Y(new_n928));
  or_6       g0653(.A(new_n928), .B(new_n927), .Y(new_n929));
  nand_5     g0654(.A(new_n929), .B(new_n926), .Y(new_n930));
  or_6       g0655(.A(new_n930), .B(new_n914), .Y(new_n931));
  nand_5     g0656(.A(new_n931), .B(new_n913), .Y(new_n932));
  nand_5     g0657(.A(new_n932), .B(new_n910), .Y(new_n933));
  nand_5     g0658(.A(new_n933), .B(new_n909), .Y(new_n934));
  or_6       g0659(.A(new_n934), .B(new_n906), .Y(new_n935));
  nand_5     g0660(.A(new_n935), .B(new_n905), .Y(new_n936));
  or_6       g0661(.A(new_n899), .B(new_n556), .Y(new_n937));
  nand_5     g0662(.A(new_n937), .B(new_n682), .Y(new_n938));
  or_6       g0663(.A(new_n937), .B(new_n682), .Y(new_n939));
  nand_5     g0664(.A(new_n939), .B(new_n938), .Y(new_n940));
  xor_4      g0665(.A(new_n940), .B(pi01), .Y(new_n941));
  nand_5     g0666(.A(new_n902), .B(new_n900), .Y(new_n942));
  nand_5     g0667(.A(new_n942), .B(new_n901), .Y(new_n943));
  xor_4      g0668(.A(new_n943), .B(new_n941), .Y(new_n944));
  xnor_4     g0669(.A(new_n944), .B(new_n936), .Y(po015));
  xnor_4     g0670(.A(new_n930), .B(new_n914), .Y(po016));
  nand_5     g0671(.A(new_n726), .B(new_n724), .Y(new_n947));
  xor_4      g0672(.A(new_n947), .B(new_n709), .Y(po017));
  xor_4      g0673(.A(new_n693), .B(pi89), .Y(new_n949));
  xor_4      g0674(.A(new_n678), .B(pi44), .Y(new_n950));
  nand_5 g0675(.A(new_n943), .B(new_n943), .Y(new_n951));
  nand_5     g0676(.A(new_n951), .B(new_n941), .Y(new_n952));
  or_6       g0677(.A(new_n944), .B(new_n936), .Y(new_n953));
  nand_5     g0678(.A(new_n953), .B(new_n952), .Y(new_n954));
  nand_5     g0679(.A(new_n938), .B(pi01), .Y(new_n955));
  and_6      g0680(.A(new_n955), .B(new_n939), .Y(new_n956));
  or_6       g0681(.A(new_n956), .B(new_n954), .Y(new_n957));
  nand_5     g0682(.A(new_n578), .B(pi58), .Y(new_n958));
  xor_4      g0683(.A(new_n958), .B(new_n957), .Y(new_n959));
  xor_4      g0684(.A(new_n956), .B(new_n954), .Y(new_n960));
  nand_5 g0685(.A(new_n960), .B(new_n960), .Y(new_n961));
  xor_4      g0686(.A(new_n814), .B(pi58), .Y(new_n962));
  nor_5      g0687(.A(new_n962), .B(new_n961), .Y(new_n963));
  or_6       g0688(.A(new_n963), .B(new_n959), .Y(new_n964));
  nand_5     g0689(.A(new_n964), .B(new_n950), .Y(new_n965));
  nand_5     g0690(.A(new_n678), .B(pi44), .Y(new_n966));
  or_6       g0691(.A(new_n958), .B(new_n957), .Y(new_n967));
  xnor_4     g0692(.A(new_n967), .B(new_n966), .Y(new_n968));
  nand_5     g0693(.A(new_n968), .B(new_n965), .Y(new_n969));
  xor_4      g0694(.A(new_n969), .B(new_n949), .Y(po018));
  nor_5      g0695(.A(new_n295), .B(new_n276), .Y(new_n971));
  xor_4      g0696(.A(new_n971), .B(pi80), .Y(new_n972));
  nand_5 g0697(.A(new_n972), .B(new_n972), .Y(new_n973));
  nand_5     g0698(.A(new_n973), .B(new_n448), .Y(new_n974));
  xor_4      g0699(.A(new_n972), .B(pi78), .Y(new_n975));
  nand_5     g0700(.A(new_n297), .B(new_n341), .Y(new_n976));
  nand_5     g0701(.A(new_n296), .B(pi04), .Y(new_n977));
  nand_5     g0702(.A(new_n359), .B(new_n343), .Y(new_n978));
  nand_5 g0703(.A(new_n860), .B(new_n860), .Y(new_n979));
  or_6       g0704(.A(new_n979), .B(new_n841), .Y(new_n980));
  nand_5     g0705(.A(new_n980), .B(new_n978), .Y(new_n981));
  nand_5     g0706(.A(new_n981), .B(new_n977), .Y(new_n982));
  nand_5     g0707(.A(new_n982), .B(new_n976), .Y(new_n983));
  nand_5     g0708(.A(new_n983), .B(new_n975), .Y(new_n984));
  nand_5     g0709(.A(new_n984), .B(new_n974), .Y(new_n985));
  nand_5 g0710(.A(pi38), .B(pi38), .Y(new_n986));
  nand_5     g0711(.A(new_n971), .B(pi80), .Y(new_n987));
  or_6       g0712(.A(new_n987), .B(new_n986), .Y(new_n988));
  nand_5     g0713(.A(new_n987), .B(new_n986), .Y(new_n989));
  nand_5     g0714(.A(new_n989), .B(new_n988), .Y(new_n990));
  xor_4      g0715(.A(new_n990), .B(pi20), .Y(new_n991));
  nor_5      g0716(.A(new_n991), .B(new_n985), .Y(new_n992));
  nand_5     g0717(.A(new_n992), .B(pi66), .Y(new_n993));
  or_6       g0718(.A(new_n992), .B(pi66), .Y(new_n994));
  nand_5     g0719(.A(new_n994), .B(new_n993), .Y(new_n995));
  nand_5     g0720(.A(new_n988), .B(new_n447), .Y(new_n996));
  nand_5     g0721(.A(new_n996), .B(new_n989), .Y(new_n997));
  xor_4      g0722(.A(new_n997), .B(new_n995), .Y(new_n998));
  or_6       g0723(.A(new_n873), .B(new_n861), .Y(new_n999));
  nand_5     g0724(.A(new_n977), .B(new_n976), .Y(new_n1000));
  xor_4      g0725(.A(new_n1000), .B(new_n981), .Y(new_n1001));
  or_6       g0726(.A(new_n1001), .B(new_n999), .Y(new_n1002));
  xnor_4     g0727(.A(new_n983), .B(new_n975), .Y(new_n1003));
  or_6       g0728(.A(new_n1003), .B(new_n1002), .Y(new_n1004));
  xor_4      g0729(.A(new_n991), .B(new_n985), .Y(new_n1005));
  or_6       g0730(.A(new_n1005), .B(new_n1004), .Y(new_n1006));
  or_6       g0731(.A(new_n1006), .B(new_n998), .Y(new_n1007));
  or_6       g0732(.A(new_n1007), .B(po145), .Y(new_n1008));
  nand_5 g0733(.A(new_n1006), .B(new_n1006), .Y(new_n1009));
  nand_5     g0734(.A(new_n1009), .B(po047), .Y(new_n1010));
  nand_5     g0735(.A(new_n1010), .B(new_n998), .Y(new_n1011));
  nand_5     g0736(.A(new_n1011), .B(new_n1008), .Y(po019));
  or_6       g0737(.A(new_n619), .B(new_n391), .Y(new_n1013));
  nand_5     g0738(.A(new_n625), .B(new_n378), .Y(new_n1014));
  xor_4      g0739(.A(new_n625), .B(new_n378), .Y(new_n1015));
  or_6       g0740(.A(new_n632), .B(new_n382), .Y(new_n1016));
  nand_5 g0741(.A(pi48), .B(pi48), .Y(new_n1017));
  nand_5     g0742(.A(new_n632), .B(new_n382), .Y(new_n1018));
  nand_5     g0743(.A(new_n1018), .B(new_n1016), .Y(new_n1019));
  nand_5 g0744(.A(new_n1019), .B(new_n1019), .Y(new_n1020));
  nand_5     g0745(.A(new_n1020), .B(new_n1017), .Y(new_n1021));
  nand_5     g0746(.A(new_n1021), .B(new_n1016), .Y(new_n1022));
  nand_5     g0747(.A(new_n1022), .B(new_n1015), .Y(new_n1023));
  nand_5     g0748(.A(new_n1023), .B(new_n1014), .Y(new_n1024));
  xor_4      g0749(.A(new_n619), .B(new_n391), .Y(new_n1025));
  nand_5     g0750(.A(new_n1025), .B(new_n1024), .Y(new_n1026));
  nand_5     g0751(.A(new_n1026), .B(new_n1013), .Y(new_n1027));
  or_6       g0752(.A(new_n1027), .B(new_n374), .Y(new_n1028));
  xor_4      g0753(.A(new_n1027), .B(new_n373), .Y(new_n1029));
  or_6       g0754(.A(new_n1029), .B(new_n613), .Y(new_n1030));
  nand_5     g0755(.A(new_n1030), .B(new_n1028), .Y(new_n1031));
  xor_4      g0756(.A(new_n609), .B(new_n367), .Y(new_n1032));
  xnor_4     g0757(.A(new_n1032), .B(new_n1031), .Y(po020));
  xor_4      g0758(.A(new_n763), .B(new_n383), .Y(po021));
  xor_4      g0759(.A(new_n850), .B(new_n378), .Y(po022));
  nand_5 g0760(.A(new_n743), .B(new_n743), .Y(new_n1036));
  or_6       g0761(.A(new_n967), .B(new_n966), .Y(new_n1037));
  nand_5     g0762(.A(new_n1037), .B(new_n708), .Y(new_n1038));
  xor_4      g0763(.A(new_n1037), .B(new_n708), .Y(new_n1039));
  or_6       g0764(.A(new_n693), .B(pi89), .Y(new_n1040));
  nand_5 g0765(.A(new_n949), .B(new_n949), .Y(new_n1041));
  or_6       g0766(.A(new_n969), .B(new_n1041), .Y(new_n1042));
  nand_5     g0767(.A(new_n1042), .B(new_n1040), .Y(new_n1043));
  nand_5     g0768(.A(new_n1043), .B(new_n1039), .Y(new_n1044));
  nand_5     g0769(.A(new_n1044), .B(new_n1038), .Y(new_n1045));
  nand_5     g0770(.A(new_n1045), .B(new_n1036), .Y(new_n1046));
  nand_5 g0771(.A(new_n1046), .B(new_n1046), .Y(po023));
  nand_5 g0772(.A(new_n482), .B(new_n482), .Y(new_n1048));
  or_6       g0773(.A(new_n487), .B(pi70), .Y(new_n1049));
  xnor_4     g0774(.A(new_n487), .B(pi70), .Y(new_n1050));
  or_6       g0775(.A(new_n432), .B(pi07), .Y(new_n1051));
  nand_5 g0776(.A(new_n437), .B(new_n437), .Y(new_n1052));
  nand_5     g0777(.A(new_n1052), .B(new_n433), .Y(new_n1053));
  nand_5     g0778(.A(new_n1053), .B(new_n1051), .Y(new_n1054));
  nand_5 g0779(.A(new_n1054), .B(new_n1054), .Y(new_n1055));
  or_6       g0780(.A(new_n1055), .B(new_n1050), .Y(new_n1056));
  nand_5     g0781(.A(new_n1056), .B(new_n1049), .Y(new_n1057));
  or_6       g0782(.A(new_n1057), .B(new_n1048), .Y(new_n1058));
  or_6       g0783(.A(new_n1058), .B(new_n479), .Y(new_n1059));
  xor_4      g0784(.A(new_n1059), .B(new_n474), .Y(new_n1060));
  xor_4      g0785(.A(new_n1060), .B(pi65), .Y(new_n1061));
  nand_5 g0786(.A(new_n1061), .B(new_n1061), .Y(new_n1062));
  nand_5 g0787(.A(pi50), .B(pi50), .Y(new_n1063));
  or_6       g0788(.A(pi85), .B(pi46), .Y(new_n1064));
  xor_4      g0789(.A(pi85), .B(pi46), .Y(new_n1065));
  or_6       g0790(.A(pi64), .B(pi30), .Y(new_n1066));
  xor_4      g0791(.A(pi64), .B(pi30), .Y(new_n1067));
  or_6       g0792(.A(pi42), .B(pi19), .Y(new_n1068));
  nand_5     g0793(.A(pi67), .B(pi56), .Y(new_n1069));
  xor_4      g0794(.A(pi42), .B(pi19), .Y(new_n1070));
  nand_5     g0795(.A(new_n1070), .B(new_n1069), .Y(new_n1071));
  nand_5     g0796(.A(new_n1071), .B(new_n1068), .Y(new_n1072));
  nand_5     g0797(.A(new_n1072), .B(new_n1067), .Y(new_n1073));
  nand_5     g0798(.A(new_n1073), .B(new_n1066), .Y(new_n1074));
  nand_5     g0799(.A(new_n1074), .B(new_n1065), .Y(new_n1075));
  nand_5     g0800(.A(new_n1075), .B(new_n1064), .Y(new_n1076));
  or_6       g0801(.A(new_n1076), .B(new_n1063), .Y(new_n1077));
  xor_4      g0802(.A(new_n1058), .B(new_n479), .Y(new_n1078));
  xor_4      g0803(.A(new_n1057), .B(new_n1048), .Y(new_n1079));
  nand_5 g0804(.A(new_n1079), .B(new_n1079), .Y(new_n1080));
  xor_4      g0805(.A(new_n1074), .B(new_n1065), .Y(new_n1081));
  or_6       g0806(.A(new_n1081), .B(new_n1080), .Y(new_n1082));
  xor_4      g0807(.A(new_n1081), .B(new_n1080), .Y(new_n1083));
  xor_4      g0808(.A(new_n1054), .B(new_n1050), .Y(new_n1084));
  xor_4      g0809(.A(new_n1072), .B(new_n1067), .Y(new_n1085));
  nand_5 g0810(.A(new_n1085), .B(new_n1085), .Y(new_n1086));
  or_6       g0811(.A(new_n1086), .B(new_n1084), .Y(new_n1087));
  xor_4      g0812(.A(new_n1085), .B(new_n1084), .Y(new_n1088));
  nand_5 g0813(.A(new_n421), .B(new_n421), .Y(new_n1089));
  xor_4      g0814(.A(pi67), .B(pi56), .Y(new_n1090));
  or_6       g0815(.A(new_n1090), .B(new_n1089), .Y(new_n1091));
  nand_5 g0816(.A(pi61), .B(pi61), .Y(new_n1092));
  nand_5     g0817(.A(new_n635), .B(new_n1092), .Y(new_n1093));
  xor_4      g0818(.A(pi63), .B(new_n1092), .Y(new_n1094));
  or_6       g0819(.A(new_n1094), .B(new_n413), .Y(new_n1095));
  nand_5     g0820(.A(new_n1095), .B(new_n1093), .Y(new_n1096));
  nand_5 g0821(.A(new_n1096), .B(new_n1096), .Y(new_n1097));
  xor_4      g0822(.A(new_n1090), .B(new_n421), .Y(new_n1098));
  or_6       g0823(.A(new_n1098), .B(new_n1097), .Y(new_n1099));
  nand_5     g0824(.A(new_n1099), .B(new_n1091), .Y(new_n1100));
  xor_4      g0825(.A(new_n1070), .B(new_n1069), .Y(new_n1101));
  or_6       g0826(.A(new_n1101), .B(new_n1100), .Y(new_n1102));
  xor_4      g0827(.A(new_n1101), .B(new_n1100), .Y(new_n1103));
  nand_5     g0828(.A(new_n1103), .B(new_n438), .Y(new_n1104));
  nand_5     g0829(.A(new_n1104), .B(new_n1102), .Y(new_n1105));
  or_6       g0830(.A(new_n1105), .B(new_n1088), .Y(new_n1106));
  nand_5     g0831(.A(new_n1106), .B(new_n1087), .Y(new_n1107));
  nand_5 g0832(.A(new_n1107), .B(new_n1107), .Y(new_n1108));
  nand_5     g0833(.A(new_n1108), .B(new_n1083), .Y(new_n1109));
  nand_5     g0834(.A(new_n1109), .B(new_n1082), .Y(new_n1110));
  nand_5     g0835(.A(new_n1110), .B(new_n1078), .Y(new_n1111));
  or_6       g0836(.A(new_n1111), .B(new_n1077), .Y(new_n1112));
  or_6       g0837(.A(new_n1110), .B(new_n1078), .Y(new_n1113));
  nand_5     g0838(.A(new_n1113), .B(new_n1111), .Y(new_n1114));
  xor_4      g0839(.A(new_n1076), .B(new_n1063), .Y(new_n1115));
  or_6       g0840(.A(new_n1115), .B(new_n1114), .Y(new_n1116));
  nand_5     g0841(.A(new_n1116), .B(new_n1113), .Y(new_n1117));
  nand_5     g0842(.A(new_n1117), .B(new_n1077), .Y(new_n1118));
  nand_5     g0843(.A(new_n1118), .B(new_n1112), .Y(new_n1119));
  xor_4      g0844(.A(new_n1119), .B(new_n1062), .Y(po024));
  xor_4      g0845(.A(new_n1094), .B(new_n423), .Y(po025));
  xnor_4     g0846(.A(new_n778), .B(new_n758), .Y(po026));
  or_6       g0847(.A(new_n832), .B(new_n743), .Y(new_n1123));
  nand_5 g0848(.A(new_n1123), .B(new_n1123), .Y(po076));
  xor_4      g0849(.A(new_n830), .B(new_n817), .Y(po050));
  xor_4      g0850(.A(new_n825), .B(new_n821), .Y(new_n1126));
  nand_5 g0851(.A(new_n823), .B(new_n823), .Y(new_n1127));
  nand_5     g0852(.A(new_n1127), .B(new_n637), .Y(new_n1128));
  or_6       g0853(.A(new_n822), .B(new_n637), .Y(new_n1129));
  nand_5     g0854(.A(new_n1129), .B(new_n1128), .Y(new_n1130));
  xor_4      g0855(.A(new_n1130), .B(new_n821), .Y(po066));
  nand_5     g0856(.A(po066), .B(new_n1126), .Y(new_n1132));
  xor_4      g0857(.A(new_n828), .B(new_n827), .Y(po172));
  nand_5     g0858(.A(po172), .B(new_n1132), .Y(new_n1134));
  nand_5 g0859(.A(new_n1134), .B(new_n1134), .Y(new_n1135));
  nand_5     g0860(.A(new_n1135), .B(po050), .Y(new_n1136));
  nand_5     g0861(.A(new_n1136), .B(po076), .Y(new_n1137));
  or_6       g0862(.A(new_n832), .B(new_n582), .Y(new_n1138));
  nand_5     g0863(.A(new_n1136), .B(new_n833), .Y(new_n1139));
  nand_5     g0864(.A(new_n1139), .B(new_n1138), .Y(new_n1140));
  or_6       g0865(.A(new_n1140), .B(new_n814), .Y(new_n1141));
  or_6       g0866(.A(new_n1141), .B(new_n677), .Y(new_n1142));
  or_6       g0867(.A(new_n1142), .B(new_n694), .Y(new_n1143));
  or_6       g0868(.A(new_n1143), .B(new_n708), .Y(new_n1144));
  or_6       g0869(.A(new_n1144), .B(new_n736), .Y(new_n1145));
  nand_5     g0870(.A(new_n1145), .B(new_n1137), .Y(po027));
  or_6       g0871(.A(new_n1059), .B(new_n474), .Y(new_n1147));
  xor_4      g0872(.A(new_n1147), .B(new_n466), .Y(new_n1148));
  xor_4      g0873(.A(new_n1148), .B(pi90), .Y(new_n1149));
  nor_5      g0874(.A(new_n1119), .B(new_n1062), .Y(new_n1150));
  and_6      g0875(.A(new_n1060), .B(pi65), .Y(new_n1151));
  nand_5 g0876(.A(new_n1112), .B(new_n1112), .Y(new_n1152));
  xor_4      g0877(.A(new_n1152), .B(new_n1151), .Y(new_n1153));
  nor_5      g0878(.A(new_n1153), .B(new_n1150), .Y(new_n1154));
  xnor_4     g0879(.A(new_n1154), .B(new_n1149), .Y(po028));
  nand_5 g0880(.A(new_n510), .B(new_n510), .Y(po029));
  nand_5     g0881(.A(new_n775), .B(new_n772), .Y(new_n1157));
  xor_4      g0882(.A(new_n1157), .B(new_n769), .Y(po030));
  or_6       g0883(.A(new_n428), .B(new_n375), .Y(new_n1159));
  nand_5     g0884(.A(new_n438), .B(new_n429), .Y(new_n1160));
  nand_5     g0885(.A(new_n1160), .B(new_n1159), .Y(new_n1161));
  xor_4      g0886(.A(new_n1161), .B(new_n373), .Y(new_n1162));
  xor_4      g0887(.A(new_n1162), .B(new_n1084), .Y(po031));
  nand_5 g0888(.A(new_n746), .B(new_n746), .Y(new_n1164));
  xor_4      g0889(.A(new_n1144), .B(new_n1164), .Y(po032));
  nand_5     g0890(.A(new_n1138), .B(new_n833), .Y(new_n1166));
  xor_4      g0891(.A(new_n1166), .B(new_n1136), .Y(po033));
  xor_4      g0892(.A(new_n1079), .B(new_n366), .Y(new_n1168));
  nand_5     g0893(.A(new_n1161), .B(new_n373), .Y(new_n1169));
  nand_5     g0894(.A(new_n1162), .B(new_n1084), .Y(new_n1170));
  nand_5     g0895(.A(new_n1170), .B(new_n1169), .Y(new_n1171));
  xnor_4     g0896(.A(new_n1171), .B(new_n1168), .Y(po034));
  nor_5      g0897(.A(new_n1001), .B(po047), .Y(new_n1173));
  xnor_4     g0898(.A(new_n1001), .B(new_n999), .Y(po113));
  nor_5      g0899(.A(po113), .B(po145), .Y(new_n1175));
  nor_5      g0900(.A(new_n1175), .B(new_n1173), .Y(po035));
  xnor_4     g0901(.A(new_n1043), .B(new_n1039), .Y(po036));
  xor_4      g0902(.A(new_n749), .B(new_n396), .Y(po038));
  or_6       g0903(.A(new_n833), .B(new_n814), .Y(new_n1179));
  or_6       g0904(.A(new_n1179), .B(new_n677), .Y(new_n1180));
  or_6       g0905(.A(new_n1180), .B(new_n694), .Y(new_n1181));
  or_6       g0906(.A(new_n1181), .B(new_n708), .Y(new_n1182));
  xor_4      g0907(.A(new_n1182), .B(new_n1164), .Y(po040));
  nand_5     g0908(.A(new_n990), .B(new_n456), .Y(new_n1184));
  xor_4      g0909(.A(new_n990), .B(new_n455), .Y(new_n1185));
  nand_5     g0910(.A(new_n1148), .B(new_n972), .Y(new_n1186));
  or_6       g0911(.A(new_n1147), .B(new_n466), .Y(new_n1187));
  xor_4      g0912(.A(new_n1148), .B(new_n972), .Y(new_n1188));
  nand_5 g0913(.A(new_n1188), .B(new_n1188), .Y(new_n1189));
  or_6       g0914(.A(new_n1060), .B(new_n296), .Y(new_n1190));
  or_6       g0915(.A(new_n1078), .B(new_n358), .Y(new_n1191));
  xor_4      g0916(.A(new_n1078), .B(new_n358), .Y(new_n1192));
  nand_5     g0917(.A(new_n1080), .B(new_n366), .Y(new_n1193));
  or_6       g0918(.A(new_n1171), .B(new_n1168), .Y(new_n1194));
  nand_5     g0919(.A(new_n1194), .B(new_n1193), .Y(new_n1195));
  nand_5     g0920(.A(new_n1195), .B(new_n1192), .Y(new_n1196));
  nand_5     g0921(.A(new_n1196), .B(new_n1191), .Y(new_n1197));
  xor_4      g0922(.A(new_n1060), .B(new_n296), .Y(new_n1198));
  nand_5     g0923(.A(new_n1198), .B(new_n1197), .Y(new_n1199));
  nand_5     g0924(.A(new_n1199), .B(new_n1190), .Y(new_n1200));
  or_6       g0925(.A(new_n1200), .B(new_n1189), .Y(new_n1201));
  xnor_4     g0926(.A(new_n1201), .B(new_n1187), .Y(new_n1202));
  nand_5     g0927(.A(new_n1202), .B(new_n1186), .Y(new_n1203));
  or_6       g0928(.A(new_n1203), .B(new_n1185), .Y(new_n1204));
  nand_5     g0929(.A(new_n1204), .B(new_n1184), .Y(new_n1205));
  nand_5 g0930(.A(new_n809), .B(new_n809), .Y(new_n1206));
  or_6       g0931(.A(new_n1201), .B(new_n1187), .Y(new_n1207));
  nand_5     g0932(.A(new_n1207), .B(new_n988), .Y(new_n1208));
  xor_4      g0933(.A(new_n1208), .B(new_n1206), .Y(new_n1209));
  xnor_4     g0934(.A(new_n1209), .B(new_n1205), .Y(po041));
  xor_4      g0935(.A(new_n578), .B(new_n296), .Y(new_n1211));
  nand_5     g0936(.A(new_n582), .B(new_n358), .Y(new_n1212));
  xor_4      g0937(.A(new_n900), .B(new_n367), .Y(new_n1213));
  nand_5 g0938(.A(new_n1213), .B(new_n1213), .Y(new_n1214));
  or_6       g0939(.A(new_n907), .B(new_n373), .Y(new_n1215));
  or_6       g0940(.A(new_n911), .B(new_n391), .Y(new_n1216));
  xor_4      g0941(.A(new_n911), .B(new_n391), .Y(new_n1217));
  nand_5     g0942(.A(new_n916), .B(new_n378), .Y(new_n1218));
  xor_4      g0943(.A(new_n915), .B(new_n378), .Y(new_n1219));
  nand_5     g0944(.A(new_n1020), .B(pi33), .Y(new_n1220));
  nand_5     g0945(.A(new_n1220), .B(new_n1018), .Y(new_n1221));
  or_6       g0946(.A(new_n1221), .B(new_n1219), .Y(new_n1222));
  nand_5     g0947(.A(new_n1222), .B(new_n1218), .Y(new_n1223));
  nand_5     g0948(.A(new_n1223), .B(new_n1217), .Y(new_n1224));
  nand_5     g0949(.A(new_n1224), .B(new_n1216), .Y(new_n1225));
  xor_4      g0950(.A(new_n907), .B(new_n373), .Y(new_n1226));
  nand_5     g0951(.A(new_n1226), .B(new_n1225), .Y(new_n1227));
  nand_5     g0952(.A(new_n1227), .B(new_n1215), .Y(new_n1228));
  or_6       g0953(.A(new_n1228), .B(new_n1214), .Y(new_n1229));
  or_6       g0954(.A(new_n1229), .B(new_n937), .Y(new_n1230));
  or_6       g0955(.A(new_n1230), .B(new_n1212), .Y(new_n1231));
  nand_5 g0956(.A(new_n1231), .B(new_n1231), .Y(new_n1232));
  nand_5     g0957(.A(new_n1229), .B(new_n937), .Y(new_n1233));
  nand_5     g0958(.A(new_n900), .B(new_n367), .Y(new_n1234));
  nand_5     g0959(.A(new_n1234), .B(new_n1212), .Y(new_n1235));
  or_6       g0960(.A(new_n1235), .B(new_n1233), .Y(new_n1236));
  nor_5      g0961(.A(new_n582), .B(new_n358), .Y(new_n1237));
  nand_5     g0962(.A(new_n1237), .B(new_n1230), .Y(new_n1238));
  nand_5     g0963(.A(new_n1238), .B(new_n1236), .Y(new_n1239));
  nor_5      g0964(.A(new_n1239), .B(new_n1232), .Y(new_n1240));
  nand_5     g0965(.A(new_n1240), .B(new_n1211), .Y(new_n1241));
  nand_5     g0966(.A(new_n578), .B(new_n296), .Y(new_n1242));
  xor_4      g0967(.A(new_n1232), .B(new_n1242), .Y(new_n1243));
  nand_5     g0968(.A(new_n1243), .B(new_n1241), .Y(new_n1244));
  xor_4      g0969(.A(new_n972), .B(new_n678), .Y(new_n1245));
  nand_5     g0970(.A(new_n1245), .B(new_n1244), .Y(new_n1246));
  or_6       g0971(.A(new_n1231), .B(new_n1242), .Y(new_n1247));
  nand_5     g0972(.A(new_n972), .B(new_n678), .Y(new_n1248));
  xnor_4     g0973(.A(new_n1248), .B(new_n1247), .Y(new_n1249));
  nand_5     g0974(.A(new_n1249), .B(new_n1246), .Y(new_n1250));
  xor_4      g0975(.A(new_n990), .B(new_n693), .Y(new_n1251));
  xnor_4     g0976(.A(new_n1251), .B(new_n1250), .Y(po042));
  xor_4      g0977(.A(new_n990), .B(new_n712), .Y(new_n1253));
  nand_5 g0978(.A(new_n1253), .B(new_n1253), .Y(new_n1254));
  nand_5     g0979(.A(new_n973), .B(new_n679), .Y(new_n1255));
  xor_4      g0980(.A(new_n973), .B(new_n679), .Y(new_n1256));
  nand_5     g0981(.A(new_n579), .B(new_n297), .Y(new_n1257));
  xor_4      g0982(.A(new_n579), .B(new_n296), .Y(new_n1258));
  nand_5     g0983(.A(new_n584), .B(new_n358), .Y(new_n1259));
  nand_5     g0984(.A(new_n609), .B(new_n366), .Y(new_n1260));
  or_6       g0985(.A(new_n1032), .B(new_n1031), .Y(new_n1261));
  nand_5     g0986(.A(new_n1261), .B(new_n1260), .Y(new_n1262));
  nand_5 g0987(.A(new_n1262), .B(new_n1262), .Y(new_n1263));
  xor_4      g0988(.A(new_n583), .B(new_n359), .Y(new_n1264));
  nand_5     g0989(.A(new_n1264), .B(new_n1263), .Y(new_n1265));
  nand_5     g0990(.A(new_n1265), .B(new_n1259), .Y(new_n1266));
  or_6       g0991(.A(new_n1266), .B(new_n1258), .Y(new_n1267));
  nand_5     g0992(.A(new_n1267), .B(new_n1257), .Y(new_n1268));
  nand_5     g0993(.A(new_n1268), .B(new_n1256), .Y(new_n1269));
  nand_5     g0994(.A(new_n1269), .B(new_n1255), .Y(new_n1270));
  xor_4      g0995(.A(new_n1270), .B(new_n1254), .Y(po043));
  xnor_4     g0996(.A(new_n1005), .B(new_n1004), .Y(po044));
  nand_5     g0997(.A(pi60), .B(new_n347), .Y(new_n1273));
  nand_5     g0998(.A(new_n299), .B(pi04), .Y(new_n1274));
  and_6      g0999(.A(new_n1274), .B(new_n1273), .Y(new_n1275));
  nand_5     g1000(.A(new_n1275), .B(new_n340), .Y(new_n1276));
  or_6       g1001(.A(new_n344), .B(pi04), .Y(new_n1277));
  nand_5     g1002(.A(new_n1277), .B(pi78), .Y(new_n1278));
  or_6       g1003(.A(new_n674), .B(pi39), .Y(new_n1279));
  nand_5     g1004(.A(new_n1279), .B(new_n1278), .Y(new_n1280));
  nand_5     g1005(.A(new_n1280), .B(new_n299), .Y(new_n1281));
  nor_5      g1006(.A(new_n350), .B(pi13), .Y(new_n1282));
  nand_5     g1007(.A(new_n350), .B(pi13), .Y(new_n1283));
  nand_5     g1008(.A(new_n1283), .B(pi60), .Y(new_n1284));
  or_6       g1009(.A(new_n1284), .B(new_n1282), .Y(new_n1285));
  nand_5     g1010(.A(new_n1285), .B(new_n1281), .Y(new_n1286));
  xor_4      g1011(.A(new_n1286), .B(new_n321), .Y(new_n1287));
  or_6       g1012(.A(new_n1287), .B(new_n1276), .Y(new_n1288));
  xor_4      g1013(.A(new_n1283), .B(new_n440), .Y(new_n1289));
  nand_5     g1014(.A(new_n1289), .B(pi60), .Y(new_n1290));
  xor_4      g1015(.A(new_n1279), .B(new_n447), .Y(new_n1291));
  nand_5     g1016(.A(new_n1291), .B(new_n299), .Y(new_n1292));
  nand_5     g1017(.A(new_n1292), .B(new_n1290), .Y(new_n1293));
  xor_4      g1018(.A(new_n1293), .B(new_n1288), .Y(new_n1294));
  nand_5     g1019(.A(new_n1294), .B(pi84), .Y(new_n1295));
  or_6       g1020(.A(new_n1295), .B(pi09), .Y(new_n1296));
  nand_5     g1021(.A(new_n1296), .B(pi60), .Y(new_n1297));
  and_6      g1022(.A(new_n1295), .B(pi09), .Y(new_n1298));
  or_6       g1023(.A(new_n1298), .B(new_n1297), .Y(new_n1299));
  or_6       g1024(.A(new_n1294), .B(pi20), .Y(new_n1300));
  nand_5     g1025(.A(new_n1300), .B(pi66), .Y(new_n1301));
  nand_5     g1026(.A(new_n1301), .B(new_n299), .Y(new_n1302));
  nor_5      g1027(.A(new_n1300), .B(pi66), .Y(new_n1303));
  or_6       g1028(.A(new_n1303), .B(new_n1302), .Y(new_n1304));
  nand_5     g1029(.A(new_n1304), .B(new_n1299), .Y(new_n1305));
  nand_5 g1030(.A(new_n1305), .B(new_n1305), .Y(new_n1306));
  nand_5 g1031(.A(pi15), .B(pi15), .Y(new_n1307));
  xor_4      g1032(.A(new_n1294), .B(new_n1307), .Y(new_n1308));
  xor_4      g1033(.A(new_n1286), .B(new_n1276), .Y(new_n1309));
  nand_5 g1034(.A(new_n1309), .B(new_n1309), .Y(new_n1310));
  nand_5     g1035(.A(new_n1310), .B(pi53), .Y(new_n1311));
  nand_5 g1036(.A(new_n1311), .B(new_n1311), .Y(new_n1312));
  nand_5 g1037(.A(pi83), .B(pi83), .Y(new_n1313));
  xor_4      g1038(.A(new_n355), .B(new_n1313), .Y(new_n1314));
  nand_5     g1039(.A(pi85), .B(pi27), .Y(new_n1315));
  nand_5     g1040(.A(new_n785), .B(new_n781), .Y(new_n1316));
  nand_5     g1041(.A(new_n1316), .B(new_n1315), .Y(new_n1317));
  nand_5     g1042(.A(new_n1317), .B(pi05), .Y(new_n1318));
  or_6       g1043(.A(new_n786), .B(new_n370), .Y(new_n1319));
  nand_5     g1044(.A(new_n787), .B(new_n780), .Y(new_n1320));
  nand_5     g1045(.A(new_n1320), .B(new_n1319), .Y(new_n1321));
  and_6      g1046(.A(new_n1321), .B(new_n362), .Y(new_n1322));
  and_6      g1047(.A(new_n1322), .B(new_n1318), .Y(new_n1323));
  or_6       g1048(.A(new_n1321), .B(new_n362), .Y(new_n1324));
  nor_5      g1049(.A(new_n1317), .B(pi05), .Y(new_n1325));
  nand_5     g1050(.A(new_n1325), .B(new_n1324), .Y(new_n1326));
  or_6       g1051(.A(new_n1324), .B(new_n1318), .Y(new_n1327));
  nand_5     g1052(.A(new_n1327), .B(new_n1326), .Y(new_n1328));
  nor_5      g1053(.A(new_n1328), .B(new_n1323), .Y(new_n1329));
  nand_5     g1054(.A(new_n1329), .B(new_n1314), .Y(new_n1330));
  nor_5      g1055(.A(new_n355), .B(new_n1313), .Y(new_n1331));
  nand_5 g1056(.A(new_n1327), .B(new_n1327), .Y(new_n1332));
  nor_5      g1057(.A(new_n1332), .B(new_n1331), .Y(new_n1333));
  nand_5     g1058(.A(new_n1333), .B(new_n1330), .Y(new_n1334));
  nor_5      g1059(.A(new_n1334), .B(new_n1312), .Y(new_n1335));
  nand_5     g1060(.A(new_n1332), .B(new_n1331), .Y(new_n1336));
  or_6       g1061(.A(new_n1336), .B(new_n1311), .Y(new_n1337));
  nor_5      g1062(.A(new_n1310), .B(pi53), .Y(new_n1338));
  nand_5     g1063(.A(new_n1338), .B(new_n1336), .Y(new_n1339));
  nand_5     g1064(.A(new_n1339), .B(new_n1337), .Y(new_n1340));
  nor_5      g1065(.A(new_n1340), .B(new_n1335), .Y(new_n1341));
  nand_5     g1066(.A(new_n1341), .B(new_n1308), .Y(new_n1342));
  or_6       g1067(.A(new_n1294), .B(new_n1307), .Y(new_n1343));
  and_6      g1068(.A(new_n1337), .B(new_n1343), .Y(new_n1344));
  nand_5     g1069(.A(new_n1344), .B(new_n1342), .Y(new_n1345));
  nand_5     g1070(.A(new_n1345), .B(new_n1306), .Y(new_n1346));
  or_6       g1071(.A(new_n1337), .B(new_n1343), .Y(new_n1347));
  nand_5     g1072(.A(new_n1347), .B(new_n1305), .Y(new_n1348));
  nand_5     g1073(.A(new_n1348), .B(new_n1346), .Y(new_n1349));
  nand_5     g1074(.A(new_n742), .B(new_n299), .Y(new_n1350));
  or_6       g1075(.A(new_n1350), .B(new_n1349), .Y(new_n1351));
  nand_5 g1076(.A(new_n1351), .B(new_n1351), .Y(po045));
  xnor_4     g1077(.A(po176), .B(new_n517), .Y(po046));
  or_6       g1078(.A(new_n1248), .B(new_n1247), .Y(new_n1354));
  nand_5     g1079(.A(new_n1354), .B(new_n988), .Y(new_n1355));
  or_6       g1080(.A(new_n1355), .B(new_n707), .Y(new_n1356));
  nand_5     g1081(.A(new_n990), .B(new_n694), .Y(new_n1357));
  or_6       g1082(.A(new_n1251), .B(new_n1250), .Y(new_n1358));
  nand_5     g1083(.A(new_n1358), .B(new_n1357), .Y(new_n1359));
  xor_4      g1084(.A(new_n1355), .B(new_n708), .Y(new_n1360));
  nand_5 g1085(.A(new_n1360), .B(new_n1360), .Y(new_n1361));
  nand_5     g1086(.A(new_n1361), .B(new_n1359), .Y(new_n1362));
  nand_5     g1087(.A(new_n1362), .B(new_n1356), .Y(new_n1363));
  nand_5     g1088(.A(new_n1363), .B(new_n1036), .Y(new_n1364));
  nand_5 g1089(.A(new_n1364), .B(new_n1364), .Y(po048));
  xnor_4     g1090(.A(new_n1266), .B(new_n1258), .Y(po049));
  xor_4      g1091(.A(new_n1228), .B(new_n1214), .Y(po051));
  xor_4      g1092(.A(new_n1360), .B(new_n1359), .Y(po052));
  nand_5 g1093(.A(new_n1137), .B(new_n1137), .Y(po054));
  xor_4      g1094(.A(new_n1045), .B(new_n1164), .Y(po055));
  nand_5     g1095(.A(new_n838), .B(new_n794), .Y(new_n1371));
  nand_5 g1096(.A(new_n1371), .B(new_n1371), .Y(po056));
  nand_5     g1097(.A(new_n823), .B(new_n822), .Y(new_n1373));
  xor_4      g1098(.A(new_n1373), .B(new_n638), .Y(po057));
  xor_4      g1099(.A(new_n1317), .B(pi05), .Y(new_n1375));
  xor_4      g1100(.A(new_n1321), .B(new_n362), .Y(new_n1376));
  xor_4      g1101(.A(new_n1376), .B(new_n1375), .Y(po059));
  xor_4      g1102(.A(new_n654), .B(new_n604), .Y(po060));
  xor_4      g1103(.A(new_n964), .B(new_n950), .Y(po061));
  or_6       g1104(.A(new_n1297), .B(pi09), .Y(new_n1380));
  nand_5     g1105(.A(new_n1380), .B(new_n1302), .Y(new_n1381));
  nand_5     g1106(.A(pi60), .B(pi31), .Y(new_n1382));
  nand_5     g1107(.A(pi74), .B(new_n299), .Y(new_n1383));
  nand_5     g1108(.A(new_n1383), .B(new_n1382), .Y(new_n1384));
  nand_5 g1109(.A(new_n1384), .B(new_n1384), .Y(new_n1385));
  nand_5     g1110(.A(new_n1385), .B(new_n1381), .Y(new_n1386));
  nand_5 g1111(.A(new_n988), .B(new_n988), .Y(new_n1387));
  xor_4      g1112(.A(new_n1294), .B(new_n990), .Y(new_n1388));
  nand_5     g1113(.A(new_n1310), .B(new_n972), .Y(new_n1389));
  xor_4      g1114(.A(new_n1309), .B(new_n973), .Y(new_n1390));
  or_6       g1115(.A(new_n355), .B(new_n297), .Y(new_n1391));
  or_6       g1116(.A(new_n405), .B(new_n357), .Y(new_n1392));
  nand_5     g1117(.A(new_n1392), .B(new_n1391), .Y(new_n1393));
  nand_5     g1118(.A(new_n1393), .B(new_n1390), .Y(new_n1394));
  nand_5     g1119(.A(new_n1394), .B(new_n1389), .Y(new_n1395));
  nand_5     g1120(.A(new_n1395), .B(new_n1388), .Y(new_n1396));
  nand_5     g1121(.A(new_n1396), .B(new_n1387), .Y(new_n1397));
  nor_5      g1122(.A(new_n1396), .B(new_n1387), .Y(new_n1398));
  or_6       g1123(.A(new_n1294), .B(new_n990), .Y(new_n1399));
  nand_5     g1124(.A(new_n1397), .B(new_n1399), .Y(new_n1400));
  or_6       g1125(.A(new_n1400), .B(new_n1398), .Y(new_n1401));
  or_6       g1126(.A(new_n1401), .B(new_n1305), .Y(new_n1402));
  nand_5     g1127(.A(new_n1402), .B(new_n1397), .Y(new_n1403));
  nand_5 g1128(.A(new_n1403), .B(new_n1403), .Y(new_n1404));
  or_6       g1129(.A(new_n1404), .B(new_n1386), .Y(new_n1405));
  nand_5 g1130(.A(new_n1405), .B(new_n1405), .Y(po062));
  xnor_4     g1131(.A(new_n766), .B(new_n760), .Y(po063));
  xor_4      g1132(.A(new_n1140), .B(new_n814), .Y(po065));
  xnor_4     g1133(.A(new_n1268), .B(new_n1256), .Y(po067));
  xor_4      g1134(.A(new_n1393), .B(new_n1390), .Y(po068));
  xor_4      g1135(.A(new_n1200), .B(new_n1189), .Y(po069));
  or_6       g1136(.A(new_n1007), .B(new_n741), .Y(new_n1412));
  nand_5 g1137(.A(new_n1412), .B(new_n1412), .Y(po070));
  nand_5 g1138(.A(new_n1166), .B(new_n1166), .Y(po071));
  nand_5     g1139(.A(new_n1233), .B(new_n1230), .Y(new_n1415));
  nand_5     g1140(.A(new_n1415), .B(new_n1234), .Y(new_n1416));
  xor_4      g1141(.A(new_n582), .B(new_n358), .Y(new_n1417));
  xor_4      g1142(.A(new_n1417), .B(new_n1416), .Y(po072));
  xor_4      g1143(.A(new_n988), .B(new_n709), .Y(new_n1419));
  or_6       g1144(.A(new_n990), .B(new_n712), .Y(new_n1420));
  or_6       g1145(.A(new_n1270), .B(new_n1254), .Y(new_n1421));
  nand_5     g1146(.A(new_n1421), .B(new_n1420), .Y(new_n1422));
  xor_4      g1147(.A(new_n1422), .B(new_n1419), .Y(po073));
  xor_4      g1148(.A(new_n934), .B(new_n906), .Y(po074));
  xor_4      g1149(.A(new_n1103), .B(new_n438), .Y(po075));
  or_6       g1150(.A(new_n424), .B(new_n285), .Y(new_n1426));
  nand_5     g1151(.A(new_n1426), .B(new_n415), .Y(new_n1427));
  xor_4      g1152(.A(new_n1427), .B(new_n421), .Y(po077));
  xor_4      g1153(.A(new_n1395), .B(new_n1388), .Y(po078));
  xnor_4     g1154(.A(new_n1115), .B(new_n1114), .Y(po079));
  xor_4      g1155(.A(new_n1180), .B(new_n694), .Y(po080));
  xor_4      g1156(.A(new_n1245), .B(new_n1244), .Y(po081));
  or_6       g1157(.A(new_n1208), .B(new_n1206), .Y(new_n1433));
  nand_5     g1158(.A(new_n1209), .B(new_n1205), .Y(new_n1434));
  nand_5     g1159(.A(new_n1434), .B(new_n1433), .Y(new_n1435));
  xor_4      g1160(.A(new_n1435), .B(new_n801), .Y(po082));
  xnor_4     g1161(.A(new_n663), .B(new_n662), .Y(po083));
  nand_5     g1162(.A(new_n455), .B(pi49), .Y(new_n1438));
  xor_4      g1163(.A(new_n455), .B(pi49), .Y(new_n1439));
  nand_5     g1164(.A(new_n1152), .B(new_n1151), .Y(new_n1440));
  nand_5     g1165(.A(new_n1440), .B(new_n1187), .Y(new_n1441));
  nand_5     g1166(.A(new_n1441), .B(new_n1439), .Y(new_n1442));
  nand_5     g1167(.A(new_n1442), .B(new_n1438), .Y(new_n1443));
  or_6       g1168(.A(new_n1443), .B(new_n1206), .Y(new_n1444));
  xor_4      g1169(.A(new_n1443), .B(new_n1206), .Y(new_n1445));
  xor_4      g1170(.A(new_n1441), .B(new_n1439), .Y(new_n1446));
  nand_5 g1171(.A(new_n1446), .B(new_n1446), .Y(new_n1447));
  or_6       g1172(.A(new_n1148), .B(pi90), .Y(new_n1448));
  nand_5     g1173(.A(new_n1154), .B(new_n1149), .Y(new_n1449));
  nand_5     g1174(.A(new_n1449), .B(new_n1448), .Y(new_n1450));
  or_6       g1175(.A(new_n1450), .B(new_n1447), .Y(new_n1451));
  nand_5     g1176(.A(new_n1451), .B(new_n1445), .Y(new_n1452));
  nand_5     g1177(.A(new_n1452), .B(new_n1444), .Y(new_n1453));
  xor_4      g1178(.A(new_n1453), .B(new_n801), .Y(po084));
  nand_5     g1179(.A(new_n1453), .B(new_n794), .Y(new_n1455));
  nand_5 g1180(.A(new_n1455), .B(new_n1455), .Y(po085));
  xor_4      g1181(.A(new_n920), .B(po125), .Y(po086));
  xor_4      g1182(.A(new_n1029), .B(new_n613), .Y(po087));
  nor_5      g1183(.A(new_n1003), .B(po047), .Y(new_n1459));
  xnor_4     g1184(.A(new_n1003), .B(new_n1002), .Y(po117));
  nor_5      g1185(.A(po117), .B(po145), .Y(new_n1461));
  nor_5      g1186(.A(new_n1461), .B(new_n1459), .Y(po088));
  xor_4      g1187(.A(new_n809), .B(new_n802), .Y(po089));
  xor_4      g1188(.A(new_n1141), .B(new_n677), .Y(po090));
  xor_4      g1189(.A(new_n962), .B(new_n961), .Y(po091));
  or_6       g1190(.A(new_n1008), .B(new_n741), .Y(new_n1466));
  nand_5 g1191(.A(new_n1466), .B(new_n1466), .Y(po092));
  xnor_4     g1192(.A(new_n403), .B(new_n364), .Y(po093));
  nand_5     g1193(.A(new_n1164), .B(pi35), .Y(new_n1469));
  nand_5 g1194(.A(new_n747), .B(new_n747), .Y(new_n1470));
  nand_5     g1195(.A(new_n1470), .B(new_n711), .Y(new_n1471));
  nand_5     g1196(.A(new_n1471), .B(new_n1469), .Y(new_n1472));
  or_6       g1197(.A(new_n1472), .B(new_n728), .Y(new_n1473));
  nor_5      g1198(.A(new_n1473), .B(new_n737), .Y(po094));
  xor_4      g1199(.A(new_n1240), .B(new_n1211), .Y(po095));
  or_6       g1200(.A(new_n1385), .B(new_n1381), .Y(new_n1476));
  and_6      g1201(.A(new_n1476), .B(new_n1386), .Y(new_n1477));
  xor_4      g1202(.A(new_n1477), .B(new_n1403), .Y(po096));
  xor_4      g1203(.A(new_n1450), .B(new_n1447), .Y(po097));
  xnor_4     g1204(.A(new_n1203), .B(new_n1185), .Y(po098));
  nand_5 g1205(.A(new_n1126), .B(new_n1126), .Y(po100));
  or_6       g1206(.A(new_n736), .B(new_n730), .Y(new_n1482));
  xor_4      g1207(.A(new_n1482), .B(new_n1473), .Y(po101));
  xnor_4     g1208(.A(new_n1451), .B(new_n1445), .Y(po102));
  xor_4      g1209(.A(new_n720), .B(new_n713), .Y(po103));
  or_6       g1210(.A(new_n1453), .B(new_n799), .Y(new_n1486));
  nand_5     g1211(.A(new_n1486), .B(new_n1455), .Y(po104));
  xor_4      g1212(.A(new_n519), .B(po064), .Y(po105));
  xor_4      g1213(.A(new_n413), .B(new_n382), .Y(po106));
  xor_4      g1214(.A(new_n1179), .B(new_n677), .Y(po107));
  nand_5     g1215(.A(new_n997), .B(new_n993), .Y(new_n1491));
  nand_5     g1216(.A(new_n1491), .B(new_n994), .Y(new_n1492));
  nor_5      g1217(.A(new_n1492), .B(new_n738), .Y(new_n1493));
  nand_5     g1218(.A(new_n1493), .B(new_n1007), .Y(new_n1494));
  nand_5     g1219(.A(new_n1494), .B(new_n1412), .Y(po108));
  xor_4      g1220(.A(new_n835), .B(new_n466), .Y(po109));
  xor_4      g1221(.A(new_n1477), .B(new_n1349), .Y(new_n1497));
  or_6       g1222(.A(new_n1383), .B(new_n740), .Y(new_n1498));
  nand_5     g1223(.A(new_n1498), .B(new_n1382), .Y(new_n1499));
  nand_5     g1224(.A(new_n1499), .B(new_n1497), .Y(new_n1500));
  nand_5     g1225(.A(new_n1500), .B(new_n1351), .Y(po110));
  xor_4      g1226(.A(new_n837), .B(new_n809), .Y(po111));
  or_6       g1227(.A(new_n1476), .B(new_n1403), .Y(new_n1503));
  nand_5     g1228(.A(new_n1503), .B(new_n1405), .Y(po112));
  xor_4      g1229(.A(new_n1142), .B(new_n694), .Y(po114));
  nand_5     g1230(.A(new_n511), .B(new_n491), .Y(po123));
  nand_5 g1231(.A(po123), .B(po123), .Y(po115));
  nand_5     g1232(.A(new_n988), .B(new_n709), .Y(new_n1508));
  nand_5     g1233(.A(new_n1422), .B(new_n1419), .Y(new_n1509));
  nand_5     g1234(.A(new_n1509), .B(new_n1508), .Y(new_n1510));
  or_6       g1235(.A(new_n1510), .B(new_n1470), .Y(new_n1511));
  or_6       g1236(.A(new_n1511), .B(new_n737), .Y(new_n1512));
  nand_5 g1237(.A(new_n1482), .B(new_n1482), .Y(new_n1513));
  nand_5     g1238(.A(new_n1510), .B(new_n1513), .Y(new_n1514));
  nand_5     g1239(.A(new_n1514), .B(new_n1512), .Y(po116));
  xor_4      g1240(.A(new_n401), .B(new_n372), .Y(po118));
  xnor_4     g1241(.A(new_n1223), .B(new_n1217), .Y(po119));
  xor_4      g1242(.A(new_n1373), .B(new_n637), .Y(po120));
  xor_4      g1243(.A(new_n1135), .B(po050), .Y(po121));
  xor_4      g1244(.A(new_n1009), .B(new_n998), .Y(po122));
  xor_4      g1245(.A(new_n1181), .B(new_n708), .Y(po124));
  or_6       g1246(.A(new_n1045), .B(new_n736), .Y(new_n1522));
  nand_5     g1247(.A(new_n1522), .B(new_n1046), .Y(po126));
  xor_4      g1248(.A(new_n1143), .B(new_n708), .Y(po127));
  nand_5     g1249(.A(new_n1435), .B(new_n794), .Y(new_n1525));
  nand_5 g1250(.A(new_n1525), .B(new_n1525), .Y(po128));
  xor_4      g1251(.A(new_n385), .B(new_n381), .Y(po129));
  nand_5     g1252(.A(new_n1493), .B(new_n1008), .Y(new_n1528));
  nand_5     g1253(.A(new_n1528), .B(new_n1466), .Y(po130));
  and_6      g1254(.A(new_n507), .B(new_n506), .Y(po177));
  xnor_4     g1255(.A(po177), .B(new_n520), .Y(po131));
  xor_4      g1256(.A(new_n1341), .B(new_n1308), .Y(po132));
  xor_4      g1257(.A(new_n1264), .B(new_n1263), .Y(po133));
  xor_4      g1258(.A(new_n645), .B(new_n644), .Y(po134));
  nand_5 g1259(.A(new_n1497), .B(new_n1497), .Y(po135));
  or_6       g1260(.A(new_n838), .B(new_n799), .Y(new_n1536));
  nand_5     g1261(.A(new_n1536), .B(new_n1371), .Y(po136));
  xor_4      g1262(.A(new_n1108), .B(new_n1083), .Y(po137));
  xor_4      g1263(.A(new_n1492), .B(new_n738), .Y(new_n1539));
  xnor_4     g1264(.A(new_n1539), .B(new_n1007), .Y(po138));
  nand_5     g1265(.A(po138), .B(po047), .Y(new_n1541));
  nand_5     g1266(.A(new_n1539), .B(po145), .Y(new_n1542));
  nand_5     g1267(.A(new_n1542), .B(new_n1541), .Y(po139));
  xor_4      g1268(.A(new_n507), .B(new_n474), .Y(po140));
  xor_4      g1269(.A(new_n1329), .B(new_n1314), .Y(po141));
  xnor_4     g1270(.A(new_n1221), .B(new_n1219), .Y(po142));
  xnor_4     g1271(.A(new_n1025), .B(new_n1024), .Y(po143));
  or_6       g1272(.A(new_n1182), .B(new_n736), .Y(new_n1548));
  nand_5     g1273(.A(new_n1548), .B(new_n1123), .Y(po144));
  nand_5     g1274(.A(new_n810), .B(new_n794), .Y(new_n1550));
  nand_5 g1275(.A(new_n1550), .B(new_n1550), .Y(po146));
  xor_4      g1276(.A(new_n493), .B(new_n491), .Y(po148));
  xnor_4     g1277(.A(new_n1022), .B(new_n1015), .Y(po149));
  xor_4      g1278(.A(new_n1510), .B(new_n747), .Y(po150));
  nor_5      g1279(.A(new_n1005), .B(po047), .Y(new_n1555));
  nor_5      g1280(.A(po044), .B(po145), .Y(new_n1556));
  nor_5      g1281(.A(new_n1556), .B(new_n1555), .Y(po151));
  xor_4      g1282(.A(new_n1019), .B(new_n919), .Y(po152));
  nand_5     g1283(.A(new_n623), .B(new_n622), .Y(new_n1559));
  xnor_4     g1284(.A(new_n1559), .B(new_n647), .Y(po153));
  xnor_4     g1285(.A(new_n932), .B(new_n910), .Y(po154));
  or_6       g1286(.A(new_n1338), .B(new_n1312), .Y(new_n1562));
  nand_5     g1287(.A(new_n1336), .B(new_n1334), .Y(new_n1563));
  xor_4      g1288(.A(new_n1563), .B(new_n1562), .Y(po155));
  xnor_4     g1289(.A(new_n1105), .B(new_n1088), .Y(po156));
  xor_4      g1290(.A(po172), .B(new_n1132), .Y(po157));
  xnor_4     g1291(.A(new_n649), .B(new_n617), .Y(po158));
  xor_4      g1292(.A(po162), .B(po145), .Y(po159));
  or_6       g1293(.A(new_n810), .B(new_n799), .Y(new_n1569));
  nand_5     g1294(.A(new_n1569), .B(new_n1550), .Y(po160));
  xnor_4     g1295(.A(new_n1226), .B(new_n1225), .Y(po161));
  xor_4      g1296(.A(new_n511), .B(new_n493), .Y(po163));
  xor_4      g1297(.A(new_n1098), .B(new_n1096), .Y(po164));
  nand_5 g1298(.A(new_n1512), .B(new_n1512), .Y(po165));
  nand_5     g1299(.A(po162), .B(po145), .Y(new_n1575));
  xnor_4     g1300(.A(new_n1575), .B(po147), .Y(po166));
  xnor_4     g1301(.A(new_n1198), .B(new_n1197), .Y(po167));
  xor_4      g1302(.A(new_n523), .B(new_n466), .Y(po168));
  or_6       g1303(.A(new_n1435), .B(new_n799), .Y(new_n1579));
  nand_5     g1304(.A(new_n1579), .B(new_n1525), .Y(po169));
  xor_4      g1305(.A(new_n925), .B(new_n916), .Y(po170));
  xor_4      g1306(.A(new_n1363), .B(new_n1164), .Y(po173));
  xor_4      g1307(.A(new_n1019), .B(new_n1017), .Y(po174));
  nand_5     g1308(.A(new_n1347), .B(new_n1345), .Y(new_n1584));
  xor_4      g1309(.A(new_n1584), .B(new_n1305), .Y(po175));
  xor_4      g1310(.A(new_n1401), .B(new_n1306), .Y(po178));
  xor_4      g1311(.A(new_n836), .B(new_n456), .Y(po179));
  or_6       g1312(.A(new_n1363), .B(new_n736), .Y(new_n1588));
  nand_5     g1313(.A(new_n1588), .B(new_n1364), .Y(po180));
  xnor_4     g1314(.A(new_n1195), .B(new_n1192), .Y(po181));
  buf_8      g1315(.A(po012), .Y(po039));
  buf_8      g1316(.A(po022), .Y(po171));
endmodule


