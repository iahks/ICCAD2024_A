// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Mon Aug 12 17:50:58 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119;
  wire new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n384,
    new_n385, new_n386, new_n387, new_n388, new_n389, new_n390, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1875, new_n1876, new_n1877, new_n1878, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1890, new_n1891, new_n1892,
    new_n1893, new_n1894, new_n1895, new_n1896, new_n1897, new_n1898,
    new_n1899, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019,
    new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025,
    new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031,
    new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055,
    new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061,
    new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067,
    new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896,
    new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914,
    new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944,
    new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956,
    new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962,
    new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046,
    new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052,
    new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058,
    new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064,
    new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070,
    new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076,
    new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088,
    new_n3089, new_n3090, new_n3091, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3101, new_n3102, new_n3103, new_n3104, new_n3105, new_n3106,
    new_n3107, new_n3108, new_n3109, new_n3110, new_n3111, new_n3112,
    new_n3113, new_n3114, new_n3115, new_n3116, new_n3117, new_n3118,
    new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125,
    new_n3126, new_n3127, new_n3128, new_n3129, new_n3130, new_n3131,
    new_n3132, new_n3133, new_n3134, new_n3135, new_n3136, new_n3137,
    new_n3138, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143,
    new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149,
    new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3155,
    new_n3156, new_n3157, new_n3158, new_n3159, new_n3160, new_n3161,
    new_n3162, new_n3163, new_n3164, new_n3165, new_n3166, new_n3167,
    new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173,
    new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179,
    new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185,
    new_n3186, new_n3187, new_n3188, new_n3189, new_n3190, new_n3191,
    new_n3192, new_n3193, new_n3194, new_n3195, new_n3196, new_n3197,
    new_n3198, new_n3199, new_n3200, new_n3201, new_n3202, new_n3203,
    new_n3204, new_n3205, new_n3206, new_n3207, new_n3208, new_n3209,
    new_n3210, new_n3211, new_n3212, new_n3213, new_n3214, new_n3215,
    new_n3216, new_n3217, new_n3218, new_n3219, new_n3220, new_n3221,
    new_n3222, new_n3223, new_n3224, new_n3225, new_n3226, new_n3227,
    new_n3228, new_n3229, new_n3230, new_n3231, new_n3232, new_n3233,
    new_n3234, new_n3235, new_n3236, new_n3237, new_n3238, new_n3239,
    new_n3240, new_n3241, new_n3242, new_n3243, new_n3244, new_n3245,
    new_n3246, new_n3247, new_n3248, new_n3249, new_n3250, new_n3251,
    new_n3252, new_n3253, new_n3254, new_n3255, new_n3256, new_n3257,
    new_n3258, new_n3259, new_n3260, new_n3261, new_n3262, new_n3263,
    new_n3264, new_n3265, new_n3266, new_n3267, new_n3268, new_n3269,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3513, new_n3514, new_n3515, new_n3516, new_n3517,
    new_n3518, new_n3522, new_n3523, new_n3524, new_n3525, new_n3526,
    new_n3527, new_n3528, new_n3529, new_n3530, new_n3531, new_n3532,
    new_n3533, new_n3534, new_n3535, new_n3536, new_n3537, new_n3538,
    new_n3539, new_n3540, new_n3541, new_n3542, new_n3543, new_n3544,
    new_n3545, new_n3546, new_n3547, new_n3548, new_n3549, new_n3550,
    new_n3551, new_n3552, new_n3553, new_n3554, new_n3555, new_n3556,
    new_n3557, new_n3558, new_n3559, new_n3560, new_n3561, new_n3562,
    new_n3563, new_n3564, new_n3565, new_n3566, new_n3567, new_n3568,
    new_n3569, new_n3570, new_n3571, new_n3572, new_n3573, new_n3574,
    new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4214, new_n4215, new_n4216, new_n4217,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226, new_n4227, new_n4228, new_n4229,
    new_n4230, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4812, new_n4813,
    new_n4814, new_n4815, new_n4816, new_n4817, new_n4818, new_n4819,
    new_n4820, new_n4821, new_n4822, new_n4823, new_n4824, new_n4825,
    new_n4826, new_n4827, new_n4828, new_n4829, new_n4830, new_n4831,
    new_n4832, new_n4833, new_n4834, new_n4835, new_n4836, new_n4837,
    new_n4838, new_n4839, new_n4840, new_n4841, new_n4842, new_n4843,
    new_n4844, new_n4845, new_n4846, new_n4847, new_n4848, new_n4849,
    new_n4850, new_n4851, new_n4852, new_n4853, new_n4854, new_n4855,
    new_n4856, new_n4857, new_n4858, new_n4859, new_n4860, new_n4861,
    new_n4862, new_n4863, new_n4864, new_n4865, new_n4866, new_n4867,
    new_n4868, new_n4869, new_n4870, new_n4871, new_n4872, new_n4873,
    new_n4874, new_n4875, new_n4876, new_n4877, new_n4878, new_n4879,
    new_n4880, new_n4881, new_n4882, new_n4883, new_n4884, new_n4885,
    new_n4886, new_n4887, new_n4888, new_n4889, new_n4890, new_n4891,
    new_n4892, new_n4893, new_n4894, new_n4895, new_n4896, new_n4897,
    new_n4898, new_n4899, new_n4900, new_n4901, new_n4902, new_n4903,
    new_n4904, new_n4905, new_n4906, new_n4907, new_n4908, new_n4909,
    new_n4910, new_n4911, new_n4912, new_n4913, new_n4914, new_n4915,
    new_n4916, new_n4917, new_n4918, new_n4919, new_n4920, new_n4921,
    new_n4922, new_n4923, new_n4924, new_n4925, new_n4926, new_n4927,
    new_n4928, new_n4929, new_n4930, new_n4931, new_n4932, new_n4933,
    new_n4934, new_n4935, new_n4936, new_n4937, new_n4938, new_n4939,
    new_n4940, new_n4941, new_n4942, new_n4943, new_n4944, new_n4945,
    new_n4946, new_n4947, new_n4948, new_n4949, new_n4950, new_n4951,
    new_n4952, new_n4953, new_n4954, new_n4955, new_n4956, new_n4957,
    new_n4958, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970,
    new_n4971, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020,
    new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026,
    new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6377, new_n6378, new_n6379,
    new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385,
    new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391,
    new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397,
    new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429, new_n6430, new_n6431, new_n6432, new_n6433,
    new_n6434, new_n6435, new_n6436, new_n6437, new_n6438, new_n6439,
    new_n6440, new_n6441, new_n6442, new_n6443, new_n6444, new_n6445,
    new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451,
    new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457,
    new_n6458, new_n6459, new_n6460, new_n6461, new_n6462, new_n6463,
    new_n6464, new_n6465, new_n6466, new_n6467, new_n6468, new_n6469,
    new_n6470, new_n6471, new_n6472, new_n6473, new_n6474, new_n6475,
    new_n6476, new_n6477, new_n6478, new_n6479, new_n6480, new_n6481,
    new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487,
    new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493,
    new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558,
    new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6567, new_n6568, new_n6569, new_n6570,
    new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576,
    new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582,
    new_n6583, new_n6584, new_n6585, new_n6586, new_n6587, new_n6588,
    new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611, new_n6612,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687,
    new_n6688, new_n6689, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254,
    new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278,
    new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7917, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922,
    new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959, new_n7960, new_n7961, new_n7962, new_n7963, new_n7964,
    new_n7965, new_n7966, new_n7967, new_n7968, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637, new_n8638, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663,
    new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9652, new_n9653, new_n9654, new_n9655,
    new_n9656, new_n9657, new_n9658, new_n9659, new_n9660, new_n9661,
    new_n9662, new_n9663, new_n9664, new_n9665, new_n9666, new_n9667,
    new_n9668, new_n9669, new_n9670, new_n9671, new_n9672, new_n9673,
    new_n9674, new_n9675, new_n9676, new_n9677, new_n9678, new_n9679,
    new_n9680, new_n9681, new_n9682, new_n9683, new_n9684, new_n9685,
    new_n9686, new_n9687, new_n9688, new_n9689, new_n9690, new_n9691,
    new_n9692, new_n9693, new_n9694, new_n9695, new_n9696, new_n9697,
    new_n9698, new_n9699, new_n9700, new_n9701, new_n9702, new_n9703,
    new_n9704, new_n9705, new_n9706, new_n9707, new_n9708, new_n9709,
    new_n9710, new_n9711, new_n9712, new_n9713, new_n9714, new_n9715,
    new_n9716, new_n9717, new_n9718, new_n9719, new_n9720, new_n9721,
    new_n9722, new_n9723, new_n9724, new_n9725, new_n9726, new_n9727,
    new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733,
    new_n9734, new_n9735, new_n9736, new_n9737, new_n9738, new_n9739,
    new_n9740, new_n9741, new_n9742, new_n9743, new_n9744, new_n9745,
    new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751,
    new_n9752, new_n9753, new_n9754, new_n9755, new_n9756, new_n9757,
    new_n9758, new_n9759, new_n9760, new_n9761, new_n9762, new_n9763,
    new_n9764, new_n9765, new_n9766, new_n9767, new_n9768, new_n9769,
    new_n9770, new_n9771, new_n9772, new_n9773, new_n9774, new_n9775,
    new_n9776, new_n9777, new_n9778, new_n9779, new_n9780, new_n9781,
    new_n9782, new_n9783, new_n9784, new_n9785, new_n9786, new_n9787,
    new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793,
    new_n9794, new_n9795, new_n9796, new_n9797, new_n9798, new_n9799,
    new_n9800, new_n9801, new_n9802, new_n9803, new_n9804, new_n9805,
    new_n9806, new_n9807, new_n9808, new_n9809, new_n9810, new_n9811,
    new_n9812, new_n9813, new_n9814, new_n9815, new_n9816, new_n9817,
    new_n9818, new_n9819, new_n9820, new_n9829, new_n9830, new_n9831,
    new_n9832, new_n9833, new_n9834, new_n9835, new_n9836, new_n9837,
    new_n9838, new_n9839, new_n9840, new_n9841, new_n9842, new_n9843,
    new_n9844, new_n9845, new_n9846, new_n9847, new_n9848, new_n9849,
    new_n9850, new_n9851, new_n9852, new_n9853, new_n9854, new_n9855,
    new_n9856, new_n9857, new_n9858, new_n9859, new_n9860, new_n9861,
    new_n9862, new_n9863, new_n9864, new_n9865, new_n9866, new_n9867,
    new_n9868, new_n9869, new_n9870, new_n9871, new_n9872, new_n9873,
    new_n9874, new_n9875, new_n9876, new_n9877, new_n9878, new_n9879,
    new_n9880, new_n9881, new_n9882, new_n9883, new_n9884, new_n9885,
    new_n9886, new_n9887, new_n9888, new_n9889, new_n9890, new_n9891,
    new_n9892, new_n9893, new_n9894, new_n9895, new_n9896, new_n9897,
    new_n9898, new_n9899, new_n9900, new_n9901, new_n9902, new_n9903,
    new_n9904, new_n9905, new_n9906, new_n9907, new_n9908, new_n9909,
    new_n9910, new_n9911, new_n9912, new_n9913, new_n9914, new_n9915,
    new_n9916, new_n9917, new_n9918, new_n9919, new_n9920, new_n9921,
    new_n9922, new_n9923, new_n9924, new_n9925, new_n9926, new_n9927,
    new_n9928, new_n9929, new_n9930, new_n9931, new_n9932, new_n9933,
    new_n9934, new_n9935, new_n9936, new_n9937, new_n9938, new_n9939,
    new_n9940, new_n9941, new_n9942, new_n9943, new_n9944, new_n9945,
    new_n9946, new_n9947, new_n9948, new_n9949, new_n9950, new_n9951,
    new_n9952, new_n9953, new_n9954, new_n9955, new_n9956, new_n9957,
    new_n9958, new_n9959, new_n9960, new_n9961, new_n9962, new_n9963,
    new_n9964, new_n9965, new_n9966, new_n9967, new_n9968, new_n9969,
    new_n9970, new_n9971, new_n9972, new_n9973, new_n9974, new_n9975,
    new_n9976, new_n9977, new_n9978, new_n9979, new_n9980, new_n9981,
    new_n9982, new_n9983, new_n9984, new_n9985, new_n9986, new_n9987,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009, new_n10010, new_n10011,
    new_n10012, new_n10013, new_n10014, new_n10015, new_n10016, new_n10017,
    new_n10018, new_n10019, new_n10020, new_n10021, new_n10022, new_n10023,
    new_n10024, new_n10025, new_n10026, new_n10027, new_n10028, new_n10029,
    new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035,
    new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041,
    new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047,
    new_n10048, new_n10049, new_n10050, new_n10051, new_n10052, new_n10053,
    new_n10054, new_n10055, new_n10056, new_n10057, new_n10058, new_n10059,
    new_n10060, new_n10061, new_n10062, new_n10063, new_n10064, new_n10065,
    new_n10066, new_n10067, new_n10068, new_n10069, new_n10070, new_n10071,
    new_n10072, new_n10073, new_n10074, new_n10075, new_n10076, new_n10077,
    new_n10078, new_n10079, new_n10080, new_n10081, new_n10082, new_n10083,
    new_n10084, new_n10085, new_n10086, new_n10087, new_n10088, new_n10089,
    new_n10090, new_n10091, new_n10092, new_n10093, new_n10094, new_n10095,
    new_n10096, new_n10097, new_n10098, new_n10099, new_n10100, new_n10101,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111, new_n10112, new_n10113,
    new_n10114, new_n10115, new_n10116, new_n10117, new_n10118, new_n10119,
    new_n10120, new_n10121, new_n10122, new_n10123, new_n10124, new_n10125,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158, new_n10159, new_n10160, new_n10161,
    new_n10162, new_n10163, new_n10164, new_n10165, new_n10166, new_n10167,
    new_n10168, new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174, new_n10175, new_n10176, new_n10177, new_n10178, new_n10179,
    new_n10180, new_n10181, new_n10182, new_n10183, new_n10184, new_n10185,
    new_n10186, new_n10187, new_n10188, new_n10189, new_n10190, new_n10191,
    new_n10192, new_n10193, new_n10194, new_n10195, new_n10196, new_n10197,
    new_n10198, new_n10199, new_n10200, new_n10201, new_n10202, new_n10203,
    new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209,
    new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215,
    new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236, new_n10237, new_n10238, new_n10239,
    new_n10240, new_n10241, new_n10242, new_n10243, new_n10244, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250, new_n10251,
    new_n10252, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10263,
    new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274, new_n10275,
    new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283, new_n10284, new_n10285, new_n10286, new_n10287,
    new_n10288, new_n10289, new_n10290, new_n10291, new_n10292, new_n10293,
    new_n10294, new_n10295, new_n10296, new_n10297, new_n10298, new_n10299,
    new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305,
    new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311,
    new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317,
    new_n10318, new_n10319, new_n10320, new_n10323, new_n10324, new_n10325,
    new_n10326, new_n10327, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361,
    new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367,
    new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385,
    new_n10386, new_n10387, new_n10388, new_n10389, new_n10390, new_n10391,
    new_n10392, new_n10393, new_n10394, new_n10395, new_n10396, new_n10397,
    new_n10398, new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404, new_n10405, new_n10406, new_n10407, new_n10408, new_n10409,
    new_n10410, new_n10411, new_n10412, new_n10413, new_n10414, new_n10415,
    new_n10416, new_n10417, new_n10418, new_n10419, new_n10420, new_n10421,
    new_n10422, new_n10423, new_n10424, new_n10425, new_n10426, new_n10427,
    new_n10428, new_n10429, new_n10430, new_n10431, new_n10432, new_n10433,
    new_n10434, new_n10435, new_n10436, new_n10437, new_n10438, new_n10439,
    new_n10440, new_n10441, new_n10442, new_n10443, new_n10444, new_n10445,
    new_n10446, new_n10447, new_n10448, new_n10449, new_n10450, new_n10451,
    new_n10452, new_n10453, new_n10454, new_n10455, new_n10456, new_n10457,
    new_n10458, new_n10459, new_n10460, new_n10461, new_n10462, new_n10463,
    new_n10464, new_n10465, new_n10466, new_n10467, new_n10468, new_n10469,
    new_n10470, new_n10471, new_n10472, new_n10473, new_n10474, new_n10475,
    new_n10476, new_n10477, new_n10478, new_n10479, new_n10480, new_n10481,
    new_n10482, new_n10483, new_n10484, new_n10485, new_n10486, new_n10487,
    new_n10488, new_n10489, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10505, new_n10506, new_n10507, new_n10508, new_n10509, new_n10510,
    new_n10511, new_n10512, new_n10513, new_n10514, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525, new_n10526, new_n10527, new_n10528,
    new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534,
    new_n10535, new_n10536, new_n10537, new_n10538, new_n10539, new_n10540,
    new_n10541, new_n10542, new_n10543, new_n10544, new_n10545, new_n10546,
    new_n10547, new_n10548, new_n10549, new_n10550, new_n10551, new_n10552,
    new_n10553, new_n10554, new_n10555, new_n10556, new_n10557, new_n10558,
    new_n10559, new_n10560, new_n10561, new_n10562, new_n10563, new_n10564,
    new_n10565, new_n10566, new_n10567, new_n10568, new_n10569, new_n10570,
    new_n10571, new_n10572, new_n10573, new_n10574, new_n10575, new_n10576,
    new_n10577, new_n10578, new_n10579, new_n10580, new_n10581, new_n10582,
    new_n10583, new_n10584, new_n10585, new_n10586, new_n10587, new_n10588,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593, new_n10594,
    new_n10595, new_n10596, new_n10597, new_n10598, new_n10599, new_n10600,
    new_n10601, new_n10602, new_n10603, new_n10604, new_n10605, new_n10606,
    new_n10607, new_n10608, new_n10609, new_n10610, new_n10611, new_n10612,
    new_n10613, new_n10614, new_n10615, new_n10616, new_n10617, new_n10618,
    new_n10619, new_n10620, new_n10621, new_n10622, new_n10623, new_n10624,
    new_n10625, new_n10626, new_n10627, new_n10628, new_n10629, new_n10630,
    new_n10631, new_n10632, new_n10633, new_n10634, new_n10635, new_n10636,
    new_n10637, new_n10638, new_n10639, new_n10640, new_n10641, new_n10642,
    new_n10643, new_n10644, new_n10645, new_n10646, new_n10647, new_n10648,
    new_n10649, new_n10650, new_n10651, new_n10652, new_n10653, new_n10654,
    new_n10655, new_n10656, new_n10657, new_n10658, new_n10659, new_n10660,
    new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666,
    new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10675, new_n10676, new_n10677, new_n10678,
    new_n10679, new_n10680, new_n10681, new_n10682, new_n10683, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874;
  nand g00000 ( new_n377 , pi027 , pi236 );
  nand g00001 ( new_n378 , pi164 , pi213 );
  xor  g00002 ( new_n379 , new_n377 , new_n378 );
  nand g00003 ( new_n380 , pi147 , pi168 );
  xor  g00004 ( new_n381 , new_n379 , new_n380 );
  nand g00005 ( new_n382 , pi119 , pi131 );
  xor  g00006 ( po000 , new_n381 , new_n382 );
  nand g00007 ( new_n384 , pi008 , pi245 );
  nand g00008 ( new_n385 , pi027 , pi156 );
  nand g00009 ( new_n386 , pi026 , pi201 );
  nand g00010 ( new_n387 , new_n385 , new_n386 );
  nand g00011 ( new_n388 , pi027 , pi201 );
  nand g00012 ( new_n389 , pi026 , pi156 );
  or   g00013 ( new_n390 , new_n388 , new_n389 );
  nand g00014 ( new_n391 , new_n387 , new_n390 );
  xor  g00015 ( new_n392 , new_n384 , new_n391 );
  nand g00016 ( new_n393 , pi026 , pi245 );
  nand g00017 ( new_n394 , pi008 , pi049 );
  nand g00018 ( new_n395 , new_n393 , new_n394 );
  xor  g00019 ( new_n396 , new_n393 , new_n394 );
  nand g00020 ( new_n397 , new_n388 , new_n396 );
  nand g00021 ( new_n398 , new_n395 , new_n397 );
  xor  g00022 ( new_n399 , new_n392 , new_n398 );
  nand g00023 ( new_n400 , pi056 , pi171 );
  nand g00024 ( new_n401 , pi026 , pi049 );
  nand g00025 ( new_n402 , pi008 , pi171 );
  nand g00026 ( new_n403 , new_n401 , new_n402 );
  nand g00027 ( new_n404 , pi027 , pi245 );
  xor  g00028 ( new_n405 , new_n401 , new_n402 );
  nand g00029 ( new_n406 , new_n404 , new_n405 );
  nand g00030 ( new_n407 , new_n403 , new_n406 );
  nand g00031 ( new_n408 , new_n400 , new_n407 );
  xor  g00032 ( new_n409 , new_n388 , new_n396 );
  xor  g00033 ( new_n410 , new_n400 , new_n407 );
  nand g00034 ( new_n411 , new_n409 , new_n410 );
  nand g00035 ( new_n412 , new_n408 , new_n411 );
  nand g00036 ( new_n413 , pi049 , pi056 );
  nand g00037 ( new_n414 , pi136 , pi171 );
  nand g00038 ( new_n415 , new_n413 , new_n414 );
  nand g00039 ( new_n416 , pi049 , pi136 );
  or   g00040 ( new_n417 , new_n400 , new_n416 );
  nand g00041 ( new_n418 , new_n415 , new_n417 );
  xor  g00042 ( new_n419 , new_n412 , new_n418 );
  xor  g00043 ( new_n420 , new_n399 , new_n419 );
  not  g00044 ( new_n421 , new_n420 );
  nand g00045 ( new_n422 , pi107 , pi136 );
  not  g00046 ( new_n423 , new_n422 );
  nand g00047 ( new_n424 , pi027 , pi049 );
  nand g00048 ( new_n425 , pi008 , pi107 );
  nand g00049 ( new_n426 , new_n424 , new_n425 );
  nand g00050 ( new_n427 , pi026 , pi171 );
  or   g00051 ( new_n428 , new_n424 , new_n425 );
  nand g00052 ( new_n429 , new_n427 , new_n428 );
  nand g00053 ( new_n430 , new_n426 , new_n429 );
  nand g00054 ( new_n431 , pi056 , pi107 );
  or   g00055 ( new_n432 , new_n430 , new_n431 );
  xnor g00056 ( new_n433 , new_n404 , new_n405 );
  xor  g00057 ( new_n434 , new_n430 , new_n431 );
  nand g00058 ( new_n435 , new_n433 , new_n434 );
  nand g00059 ( new_n436 , new_n432 , new_n435 );
  nand g00060 ( new_n437 , new_n423 , new_n436 );
  xor  g00061 ( new_n438 , new_n409 , new_n410 );
  xor  g00062 ( new_n439 , new_n422 , new_n436 );
  or   g00063 ( new_n440 , new_n438 , new_n439 );
  nand g00064 ( new_n441 , new_n437 , new_n440 );
  nand g00065 ( new_n442 , new_n421 , new_n441 );
  nand g00066 ( new_n443 , pi008 , pi201 );
  nand g00067 ( new_n444 , pi027 , pi063 );
  xor  g00068 ( new_n445 , new_n443 , new_n444 );
  xor  g00069 ( new_n446 , new_n389 , new_n445 );
  not  g00070 ( new_n447 , new_n446 );
  nand g00071 ( new_n448 , pi056 , pi245 );
  xor  g00072 ( new_n449 , new_n390 , new_n448 );
  xor  g00073 ( new_n450 , new_n447 , new_n449 );
  nand g00074 ( new_n451 , pi096 , pi171 );
  nand g00075 ( new_n452 , pi107 , pi235 );
  xor  g00076 ( new_n453 , new_n451 , new_n452 );
  xor  g00077 ( new_n454 , new_n416 , new_n453 );
  nand g00078 ( new_n455 , new_n384 , new_n391 );
  nand g00079 ( new_n456 , new_n392 , new_n398 );
  nand g00080 ( new_n457 , new_n455 , new_n456 );
  xor  g00081 ( new_n458 , new_n454 , new_n457 );
  xor  g00082 ( new_n459 , new_n450 , new_n458 );
  nand g00083 ( new_n460 , new_n412 , new_n418 );
  nand g00084 ( new_n461 , new_n399 , new_n419 );
  nand g00085 ( new_n462 , new_n460 , new_n461 );
  xor  g00086 ( new_n463 , new_n417 , new_n462 );
  xnor g00087 ( new_n464 , new_n459 , new_n463 );
  xnor g00088 ( new_n465 , new_n442 , new_n464 );
  nand g00089 ( new_n466 , pi096 , pi107 );
  xnor g00090 ( new_n467 , new_n433 , new_n434 );
  not  g00091 ( new_n468 , new_n427 );
  not  g00092 ( new_n469 , new_n426 );
  nand g00093 ( new_n470 , pi027 , pi107 );
  nand g00094 ( new_n471 , new_n468 , new_n470 );
  nand g00095 ( new_n472 , new_n469 , new_n471 );
  nand g00096 ( new_n473 , new_n428 , new_n472 );
  nand g00097 ( new_n474 , new_n468 , new_n473 );
  nor  g00098 ( new_n475 , new_n467 , new_n474 );
  xor  g00099 ( new_n476 , new_n438 , new_n439 );
  nand g00100 ( new_n477 , new_n475 , new_n476 );
  nand g00101 ( new_n478 , new_n466 , new_n477 );
  xor  g00102 ( new_n479 , new_n420 , new_n441 );
  xor  g00103 ( new_n480 , new_n466 , new_n477 );
  nand g00104 ( new_n481 , new_n479 , new_n480 );
  nand g00105 ( new_n482 , new_n478 , new_n481 );
  xor  g00106 ( new_n483 , new_n465 , new_n482 );
  nand g00107 ( new_n484 , pi032 , pi039 );
  nand g00108 ( new_n485 , pi116 , pi206 );
  nand g00109 ( new_n486 , pi070 , pi164 );
  nand g00110 ( new_n487 , new_n485 , new_n486 );
  nand g00111 ( new_n488 , pi116 , pi164 );
  nand g00112 ( new_n489 , pi070 , pi206 );
  or   g00113 ( new_n490 , new_n488 , new_n489 );
  nand g00114 ( new_n491 , new_n487 , new_n490 );
  xor  g00115 ( new_n492 , new_n484 , new_n491 );
  nand g00116 ( new_n493 , pi032 , pi228 );
  nand g00117 ( new_n494 , pi039 , pi206 );
  nand g00118 ( new_n495 , new_n493 , new_n494 );
  xor  g00119 ( new_n496 , new_n493 , new_n494 );
  nand g00120 ( new_n497 , new_n488 , new_n496 );
  nand g00121 ( new_n498 , new_n495 , new_n497 );
  xor  g00122 ( new_n499 , new_n492 , new_n498 );
  nand g00123 ( new_n500 , pi145 , pi228 );
  nand g00124 ( new_n501 , pi148 , pi246 );
  and  g00125 ( new_n502 , new_n500 , new_n501 );
  nand g00126 ( new_n503 , pi145 , pi148 );
  nand g00127 ( new_n504 , pi228 , pi246 );
  nor  g00128 ( new_n505 , new_n503 , new_n504 );
  or   g00129 ( new_n506 , new_n502 , new_n505 );
  xnor g00130 ( new_n507 , new_n499 , new_n506 );
  nand g00131 ( new_n508 , pi032 , pi148 );
  nand g00132 ( new_n509 , pi039 , pi164 );
  nand g00133 ( new_n510 , new_n508 , new_n509 );
  nand g00134 ( new_n511 , pi206 , pi228 );
  xor  g00135 ( new_n512 , new_n508 , new_n509 );
  nand g00136 ( new_n513 , new_n511 , new_n512 );
  nand g00137 ( new_n514 , new_n510 , new_n513 );
  nand g00138 ( new_n515 , new_n503 , new_n514 );
  xor  g00139 ( new_n516 , new_n488 , new_n496 );
  xor  g00140 ( new_n517 , new_n503 , new_n514 );
  nand g00141 ( new_n518 , new_n516 , new_n517 );
  nand g00142 ( new_n519 , new_n515 , new_n518 );
  xor  g00143 ( new_n520 , new_n507 , new_n519 );
  nand g00144 ( new_n521 , pi163 , pi246 );
  nand g00145 ( new_n522 , pi145 , pi163 );
  nand g00146 ( new_n523 , pi148 , pi206 );
  nand g00147 ( new_n524 , pi032 , pi163 );
  nand g00148 ( new_n525 , new_n523 , new_n524 );
  nand g00149 ( new_n526 , pi164 , pi228 );
  xor  g00150 ( new_n527 , new_n523 , new_n524 );
  nand g00151 ( new_n528 , new_n526 , new_n527 );
  nand g00152 ( new_n529 , new_n525 , new_n528 );
  nand g00153 ( new_n530 , new_n522 , new_n529 );
  xor  g00154 ( new_n531 , new_n511 , new_n512 );
  xor  g00155 ( new_n532 , new_n522 , new_n529 );
  nand g00156 ( new_n533 , new_n531 , new_n532 );
  nand g00157 ( new_n534 , new_n530 , new_n533 );
  or   g00158 ( new_n535 , new_n521 , new_n534 );
  xnor g00159 ( new_n536 , new_n516 , new_n517 );
  xor  g00160 ( new_n537 , new_n521 , new_n534 );
  nand g00161 ( new_n538 , new_n536 , new_n537 );
  nand g00162 ( new_n539 , new_n535 , new_n538 );
  nand g00163 ( new_n540 , new_n520 , new_n539 );
  nand g00164 ( new_n541 , pi115 , pi164 );
  nand g00165 ( new_n542 , pi032 , pi116 );
  xor  g00166 ( new_n543 , new_n541 , new_n542 );
  xor  g00167 ( new_n544 , new_n489 , new_n543 );
  nand g00168 ( new_n545 , pi039 , pi145 );
  xor  g00169 ( new_n546 , new_n490 , new_n545 );
  xor  g00170 ( new_n547 , new_n544 , new_n546 );
  nand g00171 ( new_n548 , pi114 , pi148 );
  nand g00172 ( new_n549 , pi091 , pi163 );
  xor  g00173 ( new_n550 , new_n548 , new_n549 );
  xor  g00174 ( new_n551 , new_n504 , new_n550 );
  nand g00175 ( new_n552 , new_n484 , new_n491 );
  nand g00176 ( new_n553 , new_n492 , new_n498 );
  nand g00177 ( new_n554 , new_n552 , new_n553 );
  xor  g00178 ( new_n555 , new_n551 , new_n554 );
  xnor g00179 ( new_n556 , new_n547 , new_n555 );
  nor  g00180 ( new_n557 , new_n499 , new_n506 );
  nor  g00181 ( new_n558 , new_n507 , new_n519 );
  xor  g00182 ( new_n559 , new_n505 , new_n558 );
  nor  g00183 ( new_n560 , new_n557 , new_n559 );
  not  g00184 ( new_n561 , new_n560 );
  xor  g00185 ( new_n562 , new_n556 , new_n561 );
  xor  g00186 ( new_n563 , new_n540 , new_n562 );
  nand g00187 ( new_n564 , pi114 , pi163 );
  xor  g00188 ( new_n565 , new_n526 , new_n527 );
  nand g00189 ( new_n566 , pi163 , pi164 );
  nor  g00190 ( new_n567 , new_n523 , new_n566 );
  not  g00191 ( new_n568 , new_n567 );
  nor  g00192 ( new_n569 , new_n565 , new_n568 );
  not  g00193 ( new_n570 , new_n569 );
  xor  g00194 ( new_n571 , new_n531 , new_n532 );
  nor  g00195 ( new_n572 , new_n570 , new_n571 );
  xor  g00196 ( new_n573 , new_n536 , new_n537 );
  nand g00197 ( new_n574 , new_n572 , new_n573 );
  nand g00198 ( new_n575 , new_n564 , new_n574 );
  xnor g00199 ( new_n576 , new_n520 , new_n539 );
  xor  g00200 ( new_n577 , new_n564 , new_n574 );
  nand g00201 ( new_n578 , new_n576 , new_n577 );
  nand g00202 ( new_n579 , new_n575 , new_n578 );
  xor  g00203 ( new_n580 , new_n563 , new_n579 );
  xor  g00204 ( new_n581 , new_n483 , new_n580 );
  xor  g00205 ( new_n582 , new_n479 , new_n480 );
  xor  g00206 ( new_n583 , new_n576 , new_n577 );
  nor  g00207 ( new_n584 , new_n582 , new_n583 );
  xnor g00208 ( new_n585 , new_n582 , new_n583 );
  xnor g00209 ( new_n586 , new_n475 , new_n476 );
  xnor g00210 ( new_n587 , new_n467 , new_n474 );
  nand g00211 ( new_n588 , pi026 , pi107 );
  nand g00212 ( new_n589 , pi027 , pi171 );
  xor  g00213 ( new_n590 , new_n588 , new_n589 );
  not  g00214 ( new_n591 , new_n590 );
  nand g00215 ( new_n592 , pi148 , pi164 );
  nand g00216 ( new_n593 , pi163 , pi206 );
  nand g00217 ( new_n594 , new_n592 , new_n593 );
  nand g00218 ( new_n595 , new_n568 , new_n594 );
  nand g00219 ( new_n596 , new_n591 , new_n595 );
  nor  g00220 ( new_n597 , new_n470 , new_n566 );
  xor  g00221 ( new_n598 , new_n590 , new_n595 );
  or   g00222 ( new_n599 , new_n597 , new_n598 );
  nand g00223 ( new_n600 , new_n596 , new_n599 );
  nor  g00224 ( new_n601 , new_n469 , new_n471 );
  nor  g00225 ( new_n602 , new_n473 , new_n601 );
  not  g00226 ( new_n603 , new_n602 );
  nand g00227 ( new_n604 , new_n600 , new_n603 );
  xor  g00228 ( new_n605 , new_n565 , new_n567 );
  xor  g00229 ( new_n606 , new_n600 , new_n603 );
  nand g00230 ( new_n607 , new_n605 , new_n606 );
  nand g00231 ( new_n608 , new_n604 , new_n607 );
  nand g00232 ( new_n609 , new_n587 , new_n608 );
  xor  g00233 ( new_n610 , new_n569 , new_n571 );
  xor  g00234 ( new_n611 , new_n587 , new_n608 );
  nand g00235 ( new_n612 , new_n610 , new_n611 );
  nand g00236 ( new_n613 , new_n609 , new_n612 );
  nand g00237 ( new_n614 , new_n586 , new_n613 );
  xor  g00238 ( new_n615 , new_n572 , new_n573 );
  not  g00239 ( new_n616 , new_n615 );
  xor  g00240 ( new_n617 , new_n586 , new_n613 );
  nand g00241 ( new_n618 , new_n616 , new_n617 );
  nand g00242 ( new_n619 , new_n614 , new_n618 );
  nor  g00243 ( new_n620 , new_n585 , new_n619 );
  nor  g00244 ( new_n621 , new_n584 , new_n620 );
  xor  g00245 ( new_n622 , new_n581 , new_n621 );
  nand g00246 ( new_n623 , pi019 , pi149 );
  nand g00247 ( new_n624 , pi151 , pi167 );
  nand g00248 ( new_n625 , pi147 , pi181 );
  nand g00249 ( new_n626 , new_n624 , new_n625 );
  nand g00250 ( new_n627 , pi147 , pi167 );
  nand g00251 ( new_n628 , pi151 , pi181 );
  or   g00252 ( new_n629 , new_n627 , new_n628 );
  nand g00253 ( new_n630 , new_n626 , new_n629 );
  xor  g00254 ( new_n631 , new_n623 , new_n630 );
  nand g00255 ( new_n632 , pi149 , pi151 );
  nand g00256 ( new_n633 , new_n627 , new_n632 );
  nand g00257 ( new_n634 , pi019 , pi240 );
  xor  g00258 ( new_n635 , new_n627 , new_n632 );
  nand g00259 ( new_n636 , new_n634 , new_n635 );
  nand g00260 ( new_n637 , new_n633 , new_n636 );
  xor  g00261 ( new_n638 , new_n631 , new_n637 );
  nand g00262 ( new_n639 , pi097 , pi240 );
  nand g00263 ( new_n640 , pi075 , pi134 );
  and  g00264 ( new_n641 , new_n639 , new_n640 );
  nand g00265 ( new_n642 , pi097 , pi134 );
  nand g00266 ( new_n643 , pi075 , pi240 );
  nor  g00267 ( new_n644 , new_n642 , new_n643 );
  or   g00268 ( new_n645 , new_n641 , new_n644 );
  xnor g00269 ( new_n646 , new_n638 , new_n645 );
  nand g00270 ( new_n647 , pi019 , pi134 );
  nand g00271 ( new_n648 , pi151 , pi240 );
  nand g00272 ( new_n649 , new_n647 , new_n648 );
  nand g00273 ( new_n650 , pi147 , pi149 );
  xor  g00274 ( new_n651 , new_n647 , new_n648 );
  nand g00275 ( new_n652 , new_n650 , new_n651 );
  nand g00276 ( new_n653 , new_n649 , new_n652 );
  nand g00277 ( new_n654 , new_n642 , new_n653 );
  xor  g00278 ( new_n655 , new_n634 , new_n635 );
  xor  g00279 ( new_n656 , new_n642 , new_n653 );
  nand g00280 ( new_n657 , new_n655 , new_n656 );
  nand g00281 ( new_n658 , new_n654 , new_n657 );
  xor  g00282 ( new_n659 , new_n646 , new_n658 );
  nand g00283 ( new_n660 , pi075 , pi175 );
  not  g00284 ( new_n661 , new_n660 );
  nand g00285 ( new_n662 , pi147 , pi240 );
  nand g00286 ( new_n663 , pi019 , pi175 );
  nand g00287 ( new_n664 , new_n662 , new_n663 );
  nand g00288 ( new_n665 , pi134 , pi151 );
  or   g00289 ( new_n666 , new_n662 , new_n663 );
  nand g00290 ( new_n667 , new_n665 , new_n666 );
  nand g00291 ( new_n668 , new_n664 , new_n667 );
  nand g00292 ( new_n669 , pi097 , pi175 );
  or   g00293 ( new_n670 , new_n668 , new_n669 );
  xor  g00294 ( new_n671 , new_n650 , new_n651 );
  not  g00295 ( new_n672 , new_n671 );
  xor  g00296 ( new_n673 , new_n668 , new_n669 );
  nand g00297 ( new_n674 , new_n672 , new_n673 );
  nand g00298 ( new_n675 , new_n670 , new_n674 );
  nand g00299 ( new_n676 , new_n661 , new_n675 );
  xor  g00300 ( new_n677 , new_n655 , new_n656 );
  xor  g00301 ( new_n678 , new_n660 , new_n675 );
  or   g00302 ( new_n679 , new_n677 , new_n678 );
  nand g00303 ( new_n680 , new_n676 , new_n679 );
  nand g00304 ( new_n681 , new_n659 , new_n680 );
  nand g00305 ( new_n682 , pi019 , pi167 );
  nand g00306 ( new_n683 , pi147 , pi200 );
  xor  g00307 ( new_n684 , new_n682 , new_n683 );
  xor  g00308 ( new_n685 , new_n628 , new_n684 );
  nand g00309 ( new_n686 , pi097 , pi149 );
  xor  g00310 ( new_n687 , new_n629 , new_n686 );
  xor  g00311 ( new_n688 , new_n685 , new_n687 );
  nand g00312 ( new_n689 , pi093 , pi134 );
  nand g00313 ( new_n690 , pi166 , pi175 );
  xor  g00314 ( new_n691 , new_n689 , new_n690 );
  xor  g00315 ( new_n692 , new_n643 , new_n691 );
  nand g00316 ( new_n693 , new_n623 , new_n630 );
  nand g00317 ( new_n694 , new_n631 , new_n637 );
  nand g00318 ( new_n695 , new_n693 , new_n694 );
  xor  g00319 ( new_n696 , new_n692 , new_n695 );
  xnor g00320 ( new_n697 , new_n688 , new_n696 );
  nor  g00321 ( new_n698 , new_n638 , new_n645 );
  nor  g00322 ( new_n699 , new_n646 , new_n658 );
  xor  g00323 ( new_n700 , new_n644 , new_n699 );
  nor  g00324 ( new_n701 , new_n698 , new_n700 );
  xor  g00325 ( new_n702 , new_n697 , new_n701 );
  xor  g00326 ( new_n703 , new_n681 , new_n702 );
  nand g00327 ( new_n704 , pi093 , pi175 );
  xnor g00328 ( new_n705 , new_n659 , new_n680 );
  nor  g00329 ( new_n706 , new_n704 , new_n705 );
  xor  g00330 ( new_n707 , new_n671 , new_n673 );
  not  g00331 ( new_n708 , new_n665 );
  not  g00332 ( new_n709 , new_n664 );
  nand g00333 ( new_n710 , pi147 , pi175 );
  nand g00334 ( new_n711 , new_n708 , new_n710 );
  nand g00335 ( new_n712 , new_n709 , new_n711 );
  nand g00336 ( new_n713 , new_n666 , new_n712 );
  nand g00337 ( new_n714 , new_n708 , new_n713 );
  nor  g00338 ( new_n715 , new_n707 , new_n714 );
  xor  g00339 ( new_n716 , new_n677 , new_n678 );
  nand g00340 ( new_n717 , new_n715 , new_n716 );
  xor  g00341 ( new_n718 , new_n704 , new_n705 );
  not  g00342 ( new_n719 , new_n718 );
  nor  g00343 ( new_n720 , new_n717 , new_n719 );
  or   g00344 ( new_n721 , new_n706 , new_n720 );
  xor  g00345 ( new_n722 , new_n703 , new_n721 );
  xor  g00346 ( new_n723 , new_n622 , new_n722 );
  xor  g00347 ( new_n724 , new_n585 , new_n619 );
  xor  g00348 ( new_n725 , new_n717 , new_n719 );
  nand g00349 ( new_n726 , new_n724 , new_n725 );
  xor  g00350 ( new_n727 , new_n715 , new_n716 );
  xor  g00351 ( new_n728 , new_n707 , new_n714 );
  xnor g00352 ( new_n729 , new_n605 , new_n606 );
  nor  g00353 ( new_n730 , new_n709 , new_n711 );
  nor  g00354 ( new_n731 , new_n713 , new_n730 );
  nand g00355 ( new_n732 , new_n729 , new_n731 );
  xor  g00356 ( new_n733 , new_n729 , new_n731 );
  xor  g00357 ( new_n734 , new_n470 , new_n566 );
  not  g00358 ( new_n735 , new_n734 );
  nor  g00359 ( new_n736 , new_n710 , new_n735 );
  nand g00360 ( new_n737 , pi151 , pi175 );
  nand g00361 ( new_n738 , pi134 , pi147 );
  xor  g00362 ( new_n739 , new_n737 , new_n738 );
  nand g00363 ( new_n740 , new_n736 , new_n739 );
  xor  g00364 ( new_n741 , new_n597 , new_n598 );
  not  g00365 ( new_n742 , new_n741 );
  xor  g00366 ( new_n743 , new_n736 , new_n739 );
  nand g00367 ( new_n744 , new_n742 , new_n743 );
  nand g00368 ( new_n745 , new_n740 , new_n744 );
  nand g00369 ( new_n746 , new_n733 , new_n745 );
  nand g00370 ( new_n747 , new_n732 , new_n746 );
  nand g00371 ( new_n748 , new_n728 , new_n747 );
  xnor g00372 ( new_n749 , new_n610 , new_n611 );
  xor  g00373 ( new_n750 , new_n728 , new_n747 );
  nand g00374 ( new_n751 , new_n749 , new_n750 );
  nand g00375 ( new_n752 , new_n748 , new_n751 );
  nand g00376 ( new_n753 , new_n727 , new_n752 );
  xor  g00377 ( new_n754 , new_n615 , new_n617 );
  xor  g00378 ( new_n755 , new_n727 , new_n752 );
  nand g00379 ( new_n756 , new_n754 , new_n755 );
  nand g00380 ( new_n757 , new_n753 , new_n756 );
  xor  g00381 ( new_n758 , new_n724 , new_n725 );
  nand g00382 ( new_n759 , new_n757 , new_n758 );
  nand g00383 ( new_n760 , new_n726 , new_n759 );
  xor  g00384 ( new_n761 , new_n723 , new_n760 );
  nand g00385 ( new_n762 , pi080 , pi250 );
  nand g00386 ( new_n763 , pi045 , pi080 );
  nand g00387 ( new_n764 , pi119 , pi247 );
  nand g00388 ( new_n765 , new_n763 , new_n764 );
  nand g00389 ( new_n766 , pi016 , pi250 );
  xor  g00390 ( new_n767 , new_n763 , new_n764 );
  nand g00391 ( new_n768 , new_n766 , new_n767 );
  nand g00392 ( new_n769 , new_n765 , new_n768 );
  xor  g00393 ( new_n770 , new_n762 , new_n769 );
  nand g00394 ( new_n771 , pi045 , pi247 );
  nand g00395 ( new_n772 , pi119 , pi234 );
  nand g00396 ( new_n773 , new_n771 , new_n772 );
  nand g00397 ( new_n774 , pi045 , pi234 );
  nor  g00398 ( new_n775 , new_n764 , new_n774 );
  not  g00399 ( new_n776 , new_n775 );
  nand g00400 ( new_n777 , new_n773 , new_n776 );
  xor  g00401 ( new_n778 , new_n770 , new_n777 );
  nand g00402 ( new_n779 , pi054 , pi117 );
  nand g00403 ( new_n780 , pi016 , pi044 );
  and  g00404 ( new_n781 , new_n779 , new_n780 );
  nand g00405 ( new_n782 , pi044 , pi117 );
  nand g00406 ( new_n783 , pi016 , pi054 );
  nor  g00407 ( new_n784 , new_n782 , new_n783 );
  or   g00408 ( new_n785 , new_n781 , new_n784 );
  xnor g00409 ( new_n786 , new_n778 , new_n785 );
  nand g00410 ( new_n787 , pi080 , pi119 );
  nand g00411 ( new_n788 , pi016 , pi045 );
  nand g00412 ( new_n789 , new_n787 , new_n788 );
  nand g00413 ( new_n790 , pi117 , pi250 );
  xor  g00414 ( new_n791 , new_n787 , new_n788 );
  nand g00415 ( new_n792 , new_n790 , new_n791 );
  nand g00416 ( new_n793 , new_n789 , new_n792 );
  nand g00417 ( new_n794 , new_n782 , new_n793 );
  xor  g00418 ( new_n795 , new_n766 , new_n767 );
  xor  g00419 ( new_n796 , new_n782 , new_n793 );
  nand g00420 ( new_n797 , new_n795 , new_n796 );
  nand g00421 ( new_n798 , new_n794 , new_n797 );
  xor  g00422 ( new_n799 , new_n786 , new_n798 );
  xor  g00423 ( new_n800 , new_n795 , new_n796 );
  nand g00424 ( new_n801 , pi054 , pi103 );
  or   g00425 ( new_n802 , new_n800 , new_n801 );
  xor  g00426 ( new_n803 , new_n800 , new_n801 );
  nand g00427 ( new_n804 , pi044 , pi103 );
  nand g00428 ( new_n805 , pi045 , pi117 );
  nand g00429 ( new_n806 , pi103 , pi250 );
  nand g00430 ( new_n807 , new_n805 , new_n806 );
  nand g00431 ( new_n808 , pi016 , pi119 );
  xor  g00432 ( new_n809 , new_n805 , new_n806 );
  nand g00433 ( new_n810 , new_n808 , new_n809 );
  nand g00434 ( new_n811 , new_n807 , new_n810 );
  or   g00435 ( new_n812 , new_n804 , new_n811 );
  xor  g00436 ( new_n813 , new_n804 , new_n811 );
  xnor g00437 ( new_n814 , new_n790 , new_n791 );
  nand g00438 ( new_n815 , new_n813 , new_n814 );
  nand g00439 ( new_n816 , new_n812 , new_n815 );
  nand g00440 ( new_n817 , new_n803 , new_n816 );
  nand g00441 ( new_n818 , new_n802 , new_n817 );
  nand g00442 ( new_n819 , new_n799 , new_n818 );
  nand g00443 ( new_n820 , pi247 , pi250 );
  nand g00444 ( new_n821 , pi119 , pi214 );
  xor  g00445 ( new_n822 , new_n820 , new_n821 );
  xor  g00446 ( new_n823 , new_n774 , new_n822 );
  nand g00447 ( new_n824 , pi044 , pi080 );
  xor  g00448 ( new_n825 , new_n776 , new_n824 );
  not  g00449 ( new_n826 , new_n825 );
  xor  g00450 ( new_n827 , new_n823 , new_n826 );
  nand g00451 ( new_n828 , pi103 , pi248 );
  nand g00452 ( new_n829 , pi072 , pi117 );
  xor  g00453 ( new_n830 , new_n783 , new_n829 );
  xor  g00454 ( new_n831 , new_n828 , new_n830 );
  nand g00455 ( new_n832 , new_n762 , new_n769 );
  nand g00456 ( new_n833 , new_n770 , new_n777 );
  nand g00457 ( new_n834 , new_n832 , new_n833 );
  xor  g00458 ( new_n835 , new_n831 , new_n834 );
  xor  g00459 ( new_n836 , new_n827 , new_n835 );
  nor  g00460 ( new_n837 , new_n786 , new_n798 );
  nand g00461 ( new_n838 , new_n784 , new_n837 );
  nor  g00462 ( new_n839 , new_n778 , new_n785 );
  or   g00463 ( new_n840 , new_n784 , new_n839 );
  or   g00464 ( new_n841 , new_n837 , new_n840 );
  nand g00465 ( new_n842 , new_n838 , new_n841 );
  xor  g00466 ( new_n843 , new_n836 , new_n842 );
  xnor g00467 ( new_n844 , new_n819 , new_n843 );
  xor  g00468 ( new_n845 , new_n808 , new_n809 );
  nand g00469 ( new_n846 , pi103 , pi119 );
  nor  g00470 ( new_n847 , new_n805 , new_n846 );
  not  g00471 ( new_n848 , new_n847 );
  nor  g00472 ( new_n849 , new_n845 , new_n848 );
  not  g00473 ( new_n850 , new_n849 );
  xnor g00474 ( new_n851 , new_n813 , new_n814 );
  nor  g00475 ( new_n852 , new_n850 , new_n851 );
  xor  g00476 ( new_n853 , new_n803 , new_n816 );
  nand g00477 ( new_n854 , new_n852 , new_n853 );
  nand g00478 ( new_n855 , pi072 , pi103 );
  nand g00479 ( new_n856 , new_n854 , new_n855 );
  xor  g00480 ( new_n857 , new_n799 , new_n818 );
  not  g00481 ( new_n858 , new_n857 );
  xor  g00482 ( new_n859 , new_n854 , new_n855 );
  nand g00483 ( new_n860 , new_n858 , new_n859 );
  nand g00484 ( new_n861 , new_n856 , new_n860 );
  xor  g00485 ( new_n862 , new_n844 , new_n861 );
  not  g00486 ( new_n863 , new_n862 );
  xor  g00487 ( new_n864 , new_n761 , new_n863 );
  xor  g00488 ( new_n865 , new_n857 , new_n859 );
  xnor g00489 ( new_n866 , new_n852 , new_n853 );
  xnor g00490 ( new_n867 , new_n749 , new_n750 );
  xor  g00491 ( new_n868 , new_n850 , new_n851 );
  not  g00492 ( new_n869 , new_n868 );
  nand g00493 ( new_n870 , new_n867 , new_n869 );
  xor  g00494 ( new_n871 , new_n845 , new_n847 );
  xor  g00495 ( new_n872 , new_n710 , new_n734 );
  nor  g00496 ( new_n873 , new_n846 , new_n872 );
  not  g00497 ( new_n874 , new_n873 );
  nand g00498 ( new_n875 , pi045 , pi103 );
  nand g00499 ( new_n876 , pi117 , pi119 );
  nand g00500 ( new_n877 , new_n875 , new_n876 );
  nand g00501 ( new_n878 , new_n848 , new_n877 );
  nand g00502 ( new_n879 , new_n874 , new_n878 );
  xor  g00503 ( new_n880 , new_n741 , new_n743 );
  xor  g00504 ( new_n881 , new_n874 , new_n878 );
  nand g00505 ( new_n882 , new_n880 , new_n881 );
  nand g00506 ( new_n883 , new_n879 , new_n882 );
  nand g00507 ( new_n884 , new_n871 , new_n883 );
  xor  g00508 ( new_n885 , new_n733 , new_n745 );
  not  g00509 ( new_n886 , new_n885 );
  xor  g00510 ( new_n887 , new_n871 , new_n883 );
  nand g00511 ( new_n888 , new_n886 , new_n887 );
  nand g00512 ( new_n889 , new_n884 , new_n888 );
  xor  g00513 ( new_n890 , new_n867 , new_n869 );
  nand g00514 ( new_n891 , new_n889 , new_n890 );
  nand g00515 ( new_n892 , new_n870 , new_n891 );
  or   g00516 ( new_n893 , new_n866 , new_n892 );
  xor  g00517 ( new_n894 , new_n754 , new_n755 );
  xor  g00518 ( new_n895 , new_n866 , new_n892 );
  nand g00519 ( new_n896 , new_n894 , new_n895 );
  nand g00520 ( new_n897 , new_n893 , new_n896 );
  or   g00521 ( new_n898 , new_n865 , new_n897 );
  xor  g00522 ( new_n899 , new_n757 , new_n758 );
  not  g00523 ( new_n900 , new_n899 );
  xor  g00524 ( new_n901 , new_n865 , new_n897 );
  nand g00525 ( new_n902 , new_n900 , new_n901 );
  nand g00526 ( new_n903 , new_n898 , new_n902 );
  xnor g00527 ( po001 , new_n864 , new_n903 );
  nand g00528 ( new_n905 , pi042 , pi171 );
  nand g00529 ( new_n906 , pi107 , pi108 );
  xor  g00530 ( new_n907 , new_n905 , new_n906 );
  nand g00531 ( new_n908 , pi049 , pi051 );
  xor  g00532 ( new_n909 , new_n907 , new_n908 );
  nand g00533 ( new_n910 , pi051 , pi107 );
  nor  g00534 ( new_n911 , new_n905 , new_n910 );
  not  g00535 ( new_n912 , new_n911 );
  or   g00536 ( new_n913 , new_n909 , new_n912 );
  nand g00537 ( new_n914 , pi007 , pi107 );
  nand g00538 ( new_n915 , new_n905 , new_n906 );
  nand g00539 ( new_n916 , new_n907 , new_n908 );
  nand g00540 ( new_n917 , new_n915 , new_n916 );
  xor  g00541 ( new_n918 , new_n914 , new_n917 );
  nand g00542 ( new_n919 , pi108 , pi171 );
  nand g00543 ( new_n920 , pi051 , pi245 );
  nand g00544 ( new_n921 , pi042 , pi049 );
  xor  g00545 ( new_n922 , new_n920 , new_n921 );
  xor  g00546 ( new_n923 , new_n919 , new_n922 );
  xor  g00547 ( new_n924 , new_n918 , new_n923 );
  xor  g00548 ( new_n925 , new_n913 , new_n924 );
  nand g00549 ( new_n926 , pi148 , pi178 );
  nand g00550 ( new_n927 , pi061 , pi163 );
  xor  g00551 ( new_n928 , new_n926 , new_n927 );
  nand g00552 ( new_n929 , pi188 , pi228 );
  xor  g00553 ( new_n930 , new_n928 , new_n929 );
  nand g00554 ( new_n931 , pi163 , pi188 );
  nor  g00555 ( new_n932 , new_n926 , new_n931 );
  not  g00556 ( new_n933 , new_n932 );
  or   g00557 ( new_n934 , new_n930 , new_n933 );
  nand g00558 ( new_n935 , pi061 , pi148 );
  nand g00559 ( new_n936 , pi039 , pi188 );
  nand g00560 ( new_n937 , pi178 , pi228 );
  xor  g00561 ( new_n938 , new_n936 , new_n937 );
  xor  g00562 ( new_n939 , new_n935 , new_n938 );
  nand g00563 ( new_n940 , pi012 , pi163 );
  nand g00564 ( new_n941 , new_n926 , new_n927 );
  nand g00565 ( new_n942 , new_n928 , new_n929 );
  nand g00566 ( new_n943 , new_n941 , new_n942 );
  xor  g00567 ( new_n944 , new_n940 , new_n943 );
  xor  g00568 ( new_n945 , new_n939 , new_n944 );
  xor  g00569 ( new_n946 , new_n934 , new_n945 );
  xor  g00570 ( new_n947 , new_n925 , new_n946 );
  xor  g00571 ( new_n948 , new_n930 , new_n932 );
  xor  g00572 ( new_n949 , new_n909 , new_n912 );
  not  g00573 ( new_n950 , new_n949 );
  nor  g00574 ( new_n951 , new_n948 , new_n950 );
  xor  g00575 ( new_n952 , new_n948 , new_n949 );
  nand g00576 ( new_n953 , pi042 , pi107 );
  nand g00577 ( new_n954 , pi051 , pi171 );
  nand g00578 ( new_n955 , new_n953 , new_n954 );
  nand g00579 ( new_n956 , new_n912 , new_n955 );
  nand g00580 ( new_n957 , pi163 , pi178 );
  nand g00581 ( new_n958 , pi148 , pi188 );
  nand g00582 ( new_n959 , new_n957 , new_n958 );
  nand g00583 ( new_n960 , new_n933 , new_n959 );
  nand g00584 ( new_n961 , new_n956 , new_n960 );
  nor  g00585 ( new_n962 , new_n910 , new_n931 );
  not  g00586 ( new_n963 , new_n962 );
  xor  g00587 ( new_n964 , new_n956 , new_n960 );
  nand g00588 ( new_n965 , new_n963 , new_n964 );
  nand g00589 ( new_n966 , new_n961 , new_n965 );
  nor  g00590 ( new_n967 , new_n952 , new_n966 );
  nor  g00591 ( new_n968 , new_n951 , new_n967 );
  not  g00592 ( new_n969 , new_n968 );
  xor  g00593 ( new_n970 , new_n947 , new_n969 );
  nand g00594 ( new_n971 , pi162 , pi240 );
  nand g00595 ( new_n972 , pi175 , pi179 );
  nand g00596 ( new_n973 , new_n971 , new_n972 );
  nand g00597 ( new_n974 , pi033 , pi134 );
  or   g00598 ( new_n975 , new_n971 , new_n972 );
  nand g00599 ( new_n976 , new_n974 , new_n975 );
  nand g00600 ( new_n977 , new_n973 , new_n976 );
  nand g00601 ( new_n978 , pi048 , pi175 );
  xor  g00602 ( new_n979 , new_n977 , new_n978 );
  nand g00603 ( new_n980 , pi134 , pi179 );
  nand g00604 ( new_n981 , pi149 , pi162 );
  nand g00605 ( new_n982 , pi033 , pi240 );
  xor  g00606 ( new_n983 , new_n981 , new_n982 );
  xnor g00607 ( new_n984 , new_n980 , new_n983 );
  xnor g00608 ( new_n985 , new_n979 , new_n984 );
  not  g00609 ( new_n986 , new_n974 );
  not  g00610 ( new_n987 , new_n973 );
  nand g00611 ( new_n988 , pi162 , pi175 );
  nand g00612 ( new_n989 , new_n986 , new_n988 );
  nand g00613 ( new_n990 , new_n987 , new_n989 );
  nand g00614 ( new_n991 , new_n975 , new_n990 );
  nand g00615 ( new_n992 , new_n986 , new_n991 );
  xor  g00616 ( new_n993 , new_n985 , new_n992 );
  xor  g00617 ( new_n994 , new_n952 , new_n966 );
  nor  g00618 ( new_n995 , new_n987 , new_n989 );
  nor  g00619 ( new_n996 , new_n991 , new_n995 );
  nor  g00620 ( new_n997 , new_n994 , new_n996 );
  xnor g00621 ( new_n998 , new_n994 , new_n996 );
  xor  g00622 ( new_n999 , new_n910 , new_n931 );
  not  g00623 ( new_n1000 , new_n999 );
  nor  g00624 ( new_n1001 , new_n988 , new_n1000 );
  nand g00625 ( new_n1002 , pi134 , pi162 );
  nand g00626 ( new_n1003 , pi033 , pi175 );
  xor  g00627 ( new_n1004 , new_n1002 , new_n1003 );
  nand g00628 ( new_n1005 , new_n1001 , new_n1004 );
  xor  g00629 ( new_n1006 , new_n962 , new_n964 );
  xor  g00630 ( new_n1007 , new_n1001 , new_n1004 );
  nand g00631 ( new_n1008 , new_n1006 , new_n1007 );
  nand g00632 ( new_n1009 , new_n1005 , new_n1008 );
  nor  g00633 ( new_n1010 , new_n998 , new_n1009 );
  nor  g00634 ( new_n1011 , new_n997 , new_n1010 );
  xor  g00635 ( new_n1012 , new_n993 , new_n1011 );
  xor  g00636 ( new_n1013 , new_n970 , new_n1012 );
  nand g00637 ( new_n1014 , pi057 , pi117 );
  nand g00638 ( new_n1015 , pi103 , pi194 );
  xor  g00639 ( new_n1016 , new_n1014 , new_n1015 );
  nand g00640 ( new_n1017 , pi016 , pi143 );
  xor  g00641 ( new_n1018 , new_n1016 , new_n1017 );
  nand g00642 ( new_n1019 , pi103 , pi143 );
  nor  g00643 ( new_n1020 , new_n1014 , new_n1019 );
  not  g00644 ( new_n1021 , new_n1020 );
  or   g00645 ( new_n1022 , new_n1018 , new_n1021 );
  nand g00646 ( new_n1023 , pi080 , pi143 );
  nand g00647 ( new_n1024 , pi117 , pi194 );
  nand g00648 ( new_n1025 , pi016 , pi057 );
  xor  g00649 ( new_n1026 , new_n1024 , new_n1025 );
  xor  g00650 ( new_n1027 , new_n1023 , new_n1026 );
  nand g00651 ( new_n1028 , pi085 , pi103 );
  nand g00652 ( new_n1029 , new_n1014 , new_n1015 );
  nand g00653 ( new_n1030 , new_n1016 , new_n1017 );
  nand g00654 ( new_n1031 , new_n1029 , new_n1030 );
  xor  g00655 ( new_n1032 , new_n1028 , new_n1031 );
  xor  g00656 ( new_n1033 , new_n1027 , new_n1032 );
  xor  g00657 ( new_n1034 , new_n1022 , new_n1033 );
  xor  g00658 ( new_n1035 , new_n1018 , new_n1020 );
  xor  g00659 ( new_n1036 , new_n988 , new_n999 );
  or   g00660 ( new_n1037 , new_n1019 , new_n1036 );
  nand g00661 ( new_n1038 , pi057 , pi103 );
  nand g00662 ( new_n1039 , pi117 , pi143 );
  nand g00663 ( new_n1040 , new_n1038 , new_n1039 );
  nand g00664 ( new_n1041 , new_n1021 , new_n1040 );
  nand g00665 ( new_n1042 , new_n1037 , new_n1041 );
  xor  g00666 ( new_n1043 , new_n1006 , new_n1007 );
  not  g00667 ( new_n1044 , new_n1043 );
  xor  g00668 ( new_n1045 , new_n1037 , new_n1041 );
  nand g00669 ( new_n1046 , new_n1044 , new_n1045 );
  nand g00670 ( new_n1047 , new_n1042 , new_n1046 );
  or   g00671 ( new_n1048 , new_n1035 , new_n1047 );
  xnor g00672 ( new_n1049 , new_n998 , new_n1009 );
  xor  g00673 ( new_n1050 , new_n1035 , new_n1047 );
  nand g00674 ( new_n1051 , new_n1049 , new_n1050 );
  nand g00675 ( new_n1052 , new_n1048 , new_n1051 );
  xor  g00676 ( new_n1053 , new_n1034 , new_n1052 );
  xor  g00677 ( po002 , new_n1013 , new_n1053 );
  nand g00678 ( new_n1055 , pi142 , pi164 );
  nand g00679 ( new_n1056 , pi027 , pi087 );
  xor  g00680 ( new_n1057 , new_n1055 , new_n1056 );
  nand g00681 ( new_n1058 , pi138 , pi147 );
  xor  g00682 ( new_n1059 , new_n1057 , new_n1058 );
  nand g00683 ( new_n1060 , pi119 , pi160 );
  xor  g00684 ( po003 , new_n1059 , new_n1060 );
  nand g00685 ( new_n1062 , pi208 , pi222 );
  nand g00686 ( new_n1063 , pi125 , pi168 );
  xor  g00687 ( new_n1064 , new_n1062 , new_n1063 );
  nand g00688 ( new_n1065 , pi139 , pi249 );
  xor  g00689 ( new_n1066 , new_n1064 , new_n1065 );
  nand g00690 ( new_n1067 , pi168 , pi249 );
  nor  g00691 ( new_n1068 , new_n1062 , new_n1067 );
  not  g00692 ( new_n1069 , new_n1068 );
  or   g00693 ( new_n1070 , new_n1066 , new_n1069 );
  nand g00694 ( new_n1071 , pi125 , pi208 );
  nand g00695 ( new_n1072 , pi035 , pi249 );
  nand g00696 ( new_n1073 , pi139 , pi222 );
  xor  g00697 ( new_n1074 , new_n1072 , new_n1073 );
  xor  g00698 ( new_n1075 , new_n1071 , new_n1074 );
  nand g00699 ( new_n1076 , pi168 , pi176 );
  nand g00700 ( new_n1077 , new_n1062 , new_n1063 );
  nand g00701 ( new_n1078 , new_n1064 , new_n1065 );
  nand g00702 ( new_n1079 , new_n1077 , new_n1078 );
  xor  g00703 ( new_n1080 , new_n1076 , new_n1079 );
  xor  g00704 ( new_n1081 , new_n1075 , new_n1080 );
  xor  g00705 ( new_n1082 , new_n1070 , new_n1081 );
  nand g00706 ( new_n1083 , pi161 , pi242 );
  nand g00707 ( new_n1084 , pi236 , pi252 );
  nand g00708 ( new_n1085 , new_n1083 , new_n1084 );
  nand g00709 ( new_n1086 , pi140 , pi241 );
  or   g00710 ( new_n1087 , new_n1083 , new_n1084 );
  nand g00711 ( new_n1088 , new_n1086 , new_n1087 );
  nand g00712 ( new_n1089 , new_n1085 , new_n1088 );
  nand g00713 ( new_n1090 , pi121 , pi236 );
  xor  g00714 ( new_n1091 , new_n1089 , new_n1090 );
  nand g00715 ( new_n1092 , pi140 , pi161 );
  nand g00716 ( new_n1093 , pi141 , pi242 );
  nand g00717 ( new_n1094 , pi241 , pi252 );
  xor  g00718 ( new_n1095 , new_n1093 , new_n1094 );
  xnor g00719 ( new_n1096 , new_n1092 , new_n1095 );
  xnor g00720 ( new_n1097 , new_n1091 , new_n1096 );
  not  g00721 ( new_n1098 , new_n1086 );
  not  g00722 ( new_n1099 , new_n1085 );
  nand g00723 ( new_n1100 , pi236 , pi242 );
  nand g00724 ( new_n1101 , new_n1098 , new_n1100 );
  nand g00725 ( new_n1102 , new_n1099 , new_n1101 );
  nand g00726 ( new_n1103 , new_n1087 , new_n1102 );
  nand g00727 ( new_n1104 , new_n1098 , new_n1103 );
  xnor g00728 ( new_n1105 , new_n1097 , new_n1104 );
  nand g00729 ( new_n1106 , pi104 , pi111 );
  nand g00730 ( new_n1107 , pi013 , pi210 );
  nand g00731 ( new_n1108 , pi024 , pi212 );
  xor  g00732 ( new_n1109 , new_n1107 , new_n1108 );
  xor  g00733 ( new_n1110 , new_n1106 , new_n1109 );
  nand g00734 ( new_n1111 , pi104 , pi210 );
  nand g00735 ( new_n1112 , pi024 , pi213 );
  nand g00736 ( new_n1113 , new_n1111 , new_n1112 );
  nand g00737 ( new_n1114 , pi111 , pi212 );
  or   g00738 ( new_n1115 , new_n1111 , new_n1112 );
  nand g00739 ( new_n1116 , new_n1114 , new_n1115 );
  nand g00740 ( new_n1117 , new_n1113 , new_n1116 );
  nand g00741 ( new_n1118 , pi213 , pi224 );
  xor  g00742 ( new_n1119 , new_n1117 , new_n1118 );
  xor  g00743 ( new_n1120 , new_n1110 , new_n1119 );
  not  g00744 ( new_n1121 , new_n1114 );
  not  g00745 ( new_n1122 , new_n1113 );
  nand g00746 ( new_n1123 , pi210 , pi213 );
  nand g00747 ( new_n1124 , new_n1121 , new_n1123 );
  nand g00748 ( new_n1125 , new_n1122 , new_n1124 );
  nand g00749 ( new_n1126 , new_n1115 , new_n1125 );
  nand g00750 ( new_n1127 , new_n1121 , new_n1126 );
  xor  g00751 ( new_n1128 , new_n1120 , new_n1127 );
  xor  g00752 ( new_n1129 , new_n1105 , new_n1128 );
  nor  g00753 ( new_n1130 , new_n1099 , new_n1101 );
  or   g00754 ( new_n1131 , new_n1103 , new_n1130 );
  nor  g00755 ( new_n1132 , new_n1122 , new_n1124 );
  nor  g00756 ( new_n1133 , new_n1126 , new_n1132 );
  not  g00757 ( new_n1134 , new_n1133 );
  nand g00758 ( new_n1135 , new_n1131 , new_n1134 );
  nand g00759 ( new_n1136 , pi210 , pi212 );
  nand g00760 ( new_n1137 , pi111 , pi213 );
  xor  g00761 ( new_n1138 , new_n1136 , new_n1137 );
  nand g00762 ( new_n1139 , pi241 , pi242 );
  nand g00763 ( new_n1140 , pi140 , pi236 );
  xor  g00764 ( new_n1141 , new_n1139 , new_n1140 );
  or   g00765 ( new_n1142 , new_n1138 , new_n1141 );
  nor  g00766 ( new_n1143 , new_n1100 , new_n1123 );
  not  g00767 ( new_n1144 , new_n1143 );
  xor  g00768 ( new_n1145 , new_n1138 , new_n1141 );
  nand g00769 ( new_n1146 , new_n1144 , new_n1145 );
  nand g00770 ( new_n1147 , new_n1142 , new_n1146 );
  xor  g00771 ( new_n1148 , new_n1131 , new_n1134 );
  nand g00772 ( new_n1149 , new_n1147 , new_n1148 );
  nand g00773 ( new_n1150 , new_n1135 , new_n1149 );
  xor  g00774 ( new_n1151 , new_n1129 , new_n1150 );
  xor  g00775 ( new_n1152 , new_n1082 , new_n1151 );
  xor  g00776 ( new_n1153 , new_n1147 , new_n1148 );
  xor  g00777 ( new_n1154 , new_n1066 , new_n1069 );
  not  g00778 ( new_n1155 , new_n1154 );
  or   g00779 ( new_n1156 , new_n1153 , new_n1155 );
  xor  g00780 ( new_n1157 , new_n1153 , new_n1155 );
  xor  g00781 ( new_n1158 , new_n1100 , new_n1123 );
  not  g00782 ( new_n1159 , new_n1158 );
  or   g00783 ( new_n1160 , new_n1067 , new_n1159 );
  nand g00784 ( new_n1161 , pi168 , pi222 );
  nand g00785 ( new_n1162 , pi208 , pi249 );
  nand g00786 ( new_n1163 , new_n1161 , new_n1162 );
  nand g00787 ( new_n1164 , new_n1069 , new_n1163 );
  or   g00788 ( new_n1165 , new_n1160 , new_n1164 );
  xor  g00789 ( new_n1166 , new_n1143 , new_n1145 );
  xor  g00790 ( new_n1167 , new_n1160 , new_n1164 );
  nand g00791 ( new_n1168 , new_n1166 , new_n1167 );
  nand g00792 ( new_n1169 , new_n1165 , new_n1168 );
  nand g00793 ( new_n1170 , new_n1157 , new_n1169 );
  nand g00794 ( new_n1171 , new_n1156 , new_n1170 );
  xor  g00795 ( new_n1172 , new_n1152 , new_n1171 );
  nand g00796 ( new_n1173 , pi077 , pi100 );
  nand g00797 ( new_n1174 , pi133 , pi217 );
  nand g00798 ( new_n1175 , pi052 , pi227 );
  xor  g00799 ( new_n1176 , new_n1174 , new_n1175 );
  xor  g00800 ( new_n1177 , new_n1173 , new_n1176 );
  nand g00801 ( new_n1178 , pi077 , pi217 );
  nand g00802 ( new_n1179 , pi131 , pi227 );
  nand g00803 ( new_n1180 , new_n1178 , new_n1179 );
  nand g00804 ( new_n1181 , pi052 , pi100 );
  or   g00805 ( new_n1182 , new_n1178 , new_n1179 );
  nand g00806 ( new_n1183 , new_n1181 , new_n1182 );
  nand g00807 ( new_n1184 , new_n1180 , new_n1183 );
  nand g00808 ( new_n1185 , pi081 , pi131 );
  xor  g00809 ( new_n1186 , new_n1184 , new_n1185 );
  xor  g00810 ( new_n1187 , new_n1177 , new_n1186 );
  not  g00811 ( new_n1188 , new_n1181 );
  not  g00812 ( new_n1189 , new_n1180 );
  nand g00813 ( new_n1190 , pi131 , pi217 );
  nand g00814 ( new_n1191 , new_n1188 , new_n1190 );
  nand g00815 ( new_n1192 , new_n1189 , new_n1191 );
  nand g00816 ( new_n1193 , new_n1182 , new_n1192 );
  nand g00817 ( new_n1194 , new_n1188 , new_n1193 );
  xnor g00818 ( new_n1195 , new_n1187 , new_n1194 );
  xor  g00819 ( new_n1196 , new_n1067 , new_n1158 );
  nor  g00820 ( new_n1197 , new_n1190 , new_n1196 );
  nand g00821 ( new_n1198 , pi052 , pi217 );
  nand g00822 ( new_n1199 , pi100 , pi131 );
  xor  g00823 ( new_n1200 , new_n1198 , new_n1199 );
  or   g00824 ( new_n1201 , new_n1197 , new_n1200 );
  xor  g00825 ( new_n1202 , new_n1166 , new_n1167 );
  not  g00826 ( new_n1203 , new_n1202 );
  xor  g00827 ( new_n1204 , new_n1197 , new_n1200 );
  nand g00828 ( new_n1205 , new_n1203 , new_n1204 );
  nand g00829 ( new_n1206 , new_n1201 , new_n1205 );
  nor  g00830 ( new_n1207 , new_n1189 , new_n1191 );
  or   g00831 ( new_n1208 , new_n1193 , new_n1207 );
  nand g00832 ( new_n1209 , new_n1206 , new_n1208 );
  xnor g00833 ( new_n1210 , new_n1157 , new_n1169 );
  xor  g00834 ( new_n1211 , new_n1206 , new_n1208 );
  nand g00835 ( new_n1212 , new_n1210 , new_n1211 );
  nand g00836 ( new_n1213 , new_n1209 , new_n1212 );
  xor  g00837 ( new_n1214 , new_n1195 , new_n1213 );
  xor  g00838 ( po004 , new_n1172 , new_n1214 );
  nand g00839 ( new_n1216 , pi147 , pi192 );
  nand g00840 ( new_n1217 , pi019 , pi216 );
  nand g00841 ( new_n1218 , pi019 , pi041 );
  nand g00842 ( new_n1219 , pi076 , pi147 );
  nand g00843 ( new_n1220 , new_n1218 , new_n1219 );
  nand g00844 ( new_n1221 , pi151 , pi216 );
  xor  g00845 ( new_n1222 , new_n1218 , new_n1219 );
  nand g00846 ( new_n1223 , new_n1221 , new_n1222 );
  nand g00847 ( new_n1224 , new_n1220 , new_n1223 );
  nand g00848 ( new_n1225 , pi079 , pi147 );
  nand g00849 ( new_n1226 , pi076 , pi151 );
  nand g00850 ( new_n1227 , new_n1225 , new_n1226 );
  nand g00851 ( new_n1228 , pi079 , pi151 );
  or   g00852 ( new_n1229 , new_n1219 , new_n1228 );
  nand g00853 ( new_n1230 , new_n1227 , new_n1229 );
  xor  g00854 ( new_n1231 , new_n1224 , new_n1230 );
  xor  g00855 ( new_n1232 , new_n1217 , new_n1231 );
  nand g00856 ( new_n1233 , pi041 , pi097 );
  nand g00857 ( new_n1234 , pi075 , pi182 );
  nand g00858 ( new_n1235 , new_n1233 , new_n1234 );
  nand g00859 ( new_n1236 , pi097 , pi182 );
  nand g00860 ( new_n1237 , pi041 , pi075 );
  nor  g00861 ( new_n1238 , new_n1236 , new_n1237 );
  not  g00862 ( new_n1239 , new_n1238 );
  nand g00863 ( new_n1240 , new_n1235 , new_n1239 );
  xnor g00864 ( new_n1241 , new_n1232 , new_n1240 );
  nand g00865 ( new_n1242 , pi147 , pi216 );
  nand g00866 ( new_n1243 , pi041 , pi151 );
  nand g00867 ( new_n1244 , new_n1242 , new_n1243 );
  nand g00868 ( new_n1245 , pi019 , pi182 );
  xor  g00869 ( new_n1246 , new_n1242 , new_n1243 );
  nand g00870 ( new_n1247 , new_n1245 , new_n1246 );
  nand g00871 ( new_n1248 , new_n1244 , new_n1247 );
  nand g00872 ( new_n1249 , new_n1236 , new_n1248 );
  xor  g00873 ( new_n1250 , new_n1221 , new_n1222 );
  xor  g00874 ( new_n1251 , new_n1236 , new_n1248 );
  nand g00875 ( new_n1252 , new_n1250 , new_n1251 );
  nand g00876 ( new_n1253 , new_n1249 , new_n1252 );
  xor  g00877 ( new_n1254 , new_n1241 , new_n1253 );
  nand g00878 ( new_n1255 , pi075 , pi138 );
  not  g00879 ( new_n1256 , new_n1255 );
  nand g00880 ( new_n1257 , pi097 , pi138 );
  nand g00881 ( new_n1258 , pi151 , pi182 );
  nand g00882 ( new_n1259 , pi019 , pi138 );
  nand g00883 ( new_n1260 , new_n1258 , new_n1259 );
  nand g00884 ( new_n1261 , pi041 , pi147 );
  xor  g00885 ( new_n1262 , new_n1258 , new_n1259 );
  nand g00886 ( new_n1263 , new_n1261 , new_n1262 );
  nand g00887 ( new_n1264 , new_n1260 , new_n1263 );
  or   g00888 ( new_n1265 , new_n1257 , new_n1264 );
  xnor g00889 ( new_n1266 , new_n1245 , new_n1246 );
  xor  g00890 ( new_n1267 , new_n1257 , new_n1264 );
  nand g00891 ( new_n1268 , new_n1266 , new_n1267 );
  nand g00892 ( new_n1269 , new_n1265 , new_n1268 );
  nand g00893 ( new_n1270 , new_n1256 , new_n1269 );
  xor  g00894 ( new_n1271 , new_n1250 , new_n1251 );
  xor  g00895 ( new_n1272 , new_n1255 , new_n1269 );
  or   g00896 ( new_n1273 , new_n1271 , new_n1272 );
  nand g00897 ( new_n1274 , new_n1270 , new_n1273 );
  nand g00898 ( new_n1275 , new_n1254 , new_n1274 );
  nand g00899 ( new_n1276 , pi019 , pi076 );
  nand g00900 ( new_n1277 , pi147 , pi251 );
  xor  g00901 ( new_n1278 , new_n1276 , new_n1277 );
  xor  g00902 ( new_n1279 , new_n1228 , new_n1278 );
  nand g00903 ( new_n1280 , pi097 , pi216 );
  xor  g00904 ( new_n1281 , new_n1229 , new_n1280 );
  xor  g00905 ( new_n1282 , new_n1279 , new_n1281 );
  nand g00906 ( new_n1283 , pi138 , pi166 );
  nand g00907 ( new_n1284 , pi093 , pi182 );
  xor  g00908 ( new_n1285 , new_n1283 , new_n1284 );
  xor  g00909 ( new_n1286 , new_n1237 , new_n1285 );
  nand g00910 ( new_n1287 , new_n1224 , new_n1230 );
  nand g00911 ( new_n1288 , new_n1217 , new_n1231 );
  nand g00912 ( new_n1289 , new_n1287 , new_n1288 );
  xor  g00913 ( new_n1290 , new_n1286 , new_n1289 );
  xnor g00914 ( new_n1291 , new_n1282 , new_n1290 );
  nor  g00915 ( new_n1292 , new_n1241 , new_n1253 );
  and  g00916 ( new_n1293 , new_n1238 , new_n1292 );
  or   g00917 ( new_n1294 , new_n1232 , new_n1240 );
  nand g00918 ( new_n1295 , new_n1239 , new_n1294 );
  nor  g00919 ( new_n1296 , new_n1292 , new_n1295 );
  or   g00920 ( new_n1297 , new_n1293 , new_n1296 );
  xor  g00921 ( new_n1298 , new_n1291 , new_n1297 );
  xnor g00922 ( new_n1299 , new_n1275 , new_n1298 );
  xor  g00923 ( new_n1300 , new_n1261 , new_n1262 );
  or   g00924 ( new_n1301 , new_n1058 , new_n1258 );
  or   g00925 ( new_n1302 , new_n1300 , new_n1301 );
  xnor g00926 ( new_n1303 , new_n1266 , new_n1267 );
  nor  g00927 ( new_n1304 , new_n1302 , new_n1303 );
  xor  g00928 ( new_n1305 , new_n1271 , new_n1272 );
  nand g00929 ( new_n1306 , new_n1304 , new_n1305 );
  nand g00930 ( new_n1307 , pi093 , pi138 );
  nand g00931 ( new_n1308 , new_n1306 , new_n1307 );
  xnor g00932 ( new_n1309 , new_n1254 , new_n1274 );
  xor  g00933 ( new_n1310 , new_n1306 , new_n1307 );
  nand g00934 ( new_n1311 , new_n1309 , new_n1310 );
  nand g00935 ( new_n1312 , new_n1308 , new_n1311 );
  xor  g00936 ( new_n1313 , new_n1299 , new_n1312 );
  nand g00937 ( new_n1314 , pi071 , pi145 );
  nand g00938 ( new_n1315 , pi123 , pi164 );
  nand g00939 ( new_n1316 , pi169 , pi206 );
  nand g00940 ( new_n1317 , new_n1315 , new_n1316 );
  nand g00941 ( new_n1318 , pi032 , pi071 );
  xor  g00942 ( new_n1319 , new_n1315 , new_n1316 );
  nand g00943 ( new_n1320 , new_n1318 , new_n1319 );
  nand g00944 ( new_n1321 , new_n1317 , new_n1320 );
  nand g00945 ( new_n1322 , new_n1314 , new_n1321 );
  nand g00946 ( new_n1323 , pi032 , pi169 );
  nand g00947 ( new_n1324 , pi123 , pi206 );
  nand g00948 ( new_n1325 , pi099 , pi164 );
  xor  g00949 ( new_n1326 , new_n1324 , new_n1325 );
  xor  g00950 ( new_n1327 , new_n1323 , new_n1326 );
  xor  g00951 ( new_n1328 , new_n1314 , new_n1321 );
  nand g00952 ( new_n1329 , new_n1327 , new_n1328 );
  nand g00953 ( new_n1330 , new_n1322 , new_n1329 );
  nand g00954 ( new_n1331 , pi032 , pi123 );
  nand g00955 ( new_n1332 , new_n1324 , new_n1325 );
  nand g00956 ( new_n1333 , new_n1323 , new_n1326 );
  nand g00957 ( new_n1334 , new_n1332 , new_n1333 );
  xor  g00958 ( new_n1335 , new_n1331 , new_n1334 );
  nand g00959 ( new_n1336 , pi099 , pi206 );
  nand g00960 ( new_n1337 , pi023 , pi164 );
  nand g00961 ( new_n1338 , new_n1336 , new_n1337 );
  nand g00962 ( new_n1339 , pi023 , pi206 );
  nor  g00963 ( new_n1340 , new_n1325 , new_n1339 );
  not  g00964 ( new_n1341 , new_n1340 );
  nand g00965 ( new_n1342 , new_n1338 , new_n1341 );
  xor  g00966 ( new_n1343 , new_n1335 , new_n1342 );
  nand g00967 ( new_n1344 , pi071 , pi246 );
  nand g00968 ( new_n1345 , pi145 , pi169 );
  nand g00969 ( new_n1346 , new_n1344 , new_n1345 );
  nand g00970 ( new_n1347 , pi169 , pi246 );
  or   g00971 ( new_n1348 , new_n1314 , new_n1347 );
  nand g00972 ( new_n1349 , new_n1346 , new_n1348 );
  xor  g00973 ( new_n1350 , new_n1343 , new_n1349 );
  xnor g00974 ( new_n1351 , new_n1330 , new_n1350 );
  nand g00975 ( new_n1352 , pi142 , pi246 );
  nand g00976 ( new_n1353 , pi164 , pi169 );
  nand g00977 ( new_n1354 , pi032 , pi142 );
  nand g00978 ( new_n1355 , new_n1353 , new_n1354 );
  nand g00979 ( new_n1356 , pi071 , pi206 );
  or   g00980 ( new_n1357 , new_n1353 , new_n1354 );
  nand g00981 ( new_n1358 , new_n1356 , new_n1357 );
  nand g00982 ( new_n1359 , new_n1355 , new_n1358 );
  nand g00983 ( new_n1360 , pi142 , pi145 );
  nand g00984 ( new_n1361 , new_n1359 , new_n1360 );
  xor  g00985 ( new_n1362 , new_n1318 , new_n1319 );
  xor  g00986 ( new_n1363 , new_n1359 , new_n1360 );
  nand g00987 ( new_n1364 , new_n1362 , new_n1363 );
  nand g00988 ( new_n1365 , new_n1361 , new_n1364 );
  or   g00989 ( new_n1366 , new_n1352 , new_n1365 );
  xnor g00990 ( new_n1367 , new_n1327 , new_n1328 );
  xor  g00991 ( new_n1368 , new_n1352 , new_n1365 );
  nand g00992 ( new_n1369 , new_n1367 , new_n1368 );
  nand g00993 ( new_n1370 , new_n1366 , new_n1369 );
  xnor g00994 ( new_n1371 , new_n1351 , new_n1370 );
  xor  g00995 ( new_n1372 , new_n1362 , new_n1363 );
  not  g00996 ( new_n1373 , new_n1356 );
  not  g00997 ( new_n1374 , new_n1355 );
  nand g00998 ( new_n1375 , new_n1055 , new_n1373 );
  nand g00999 ( new_n1376 , new_n1374 , new_n1375 );
  nand g01000 ( new_n1377 , new_n1357 , new_n1376 );
  nand g01001 ( new_n1378 , new_n1373 , new_n1377 );
  nor  g01002 ( new_n1379 , new_n1372 , new_n1378 );
  xor  g01003 ( new_n1380 , new_n1367 , new_n1368 );
  nand g01004 ( new_n1381 , new_n1379 , new_n1380 );
  nand g01005 ( new_n1382 , pi114 , pi142 );
  xor  g01006 ( new_n1383 , new_n1381 , new_n1382 );
  xor  g01007 ( new_n1384 , new_n1371 , new_n1383 );
  xnor g01008 ( new_n1385 , new_n1379 , new_n1380 );
  nand g01009 ( new_n1386 , pi026 , pi219 );
  nand g01010 ( new_n1387 , pi008 , pi087 );
  xor  g01011 ( new_n1388 , new_n1386 , new_n1387 );
  nand g01012 ( new_n1389 , pi027 , pi102 );
  xor  g01013 ( new_n1390 , new_n1388 , new_n1389 );
  nor  g01014 ( new_n1391 , new_n1056 , new_n1386 );
  not  g01015 ( new_n1392 , new_n1391 );
  nor  g01016 ( new_n1393 , new_n1390 , new_n1392 );
  nand g01017 ( new_n1394 , pi056 , pi087 );
  nand g01018 ( new_n1395 , new_n1386 , new_n1387 );
  nand g01019 ( new_n1396 , new_n1388 , new_n1389 );
  nand g01020 ( new_n1397 , new_n1395 , new_n1396 );
  xor  g01021 ( new_n1398 , new_n1394 , new_n1397 );
  nand g01022 ( new_n1399 , pi008 , pi219 );
  nand g01023 ( new_n1400 , pi026 , pi102 );
  nand g01024 ( new_n1401 , pi001 , pi027 );
  xor  g01025 ( new_n1402 , new_n1400 , new_n1401 );
  xnor g01026 ( new_n1403 , new_n1399 , new_n1402 );
  xnor g01027 ( new_n1404 , new_n1398 , new_n1403 );
  xor  g01028 ( new_n1405 , new_n1393 , new_n1404 );
  nand g01029 ( new_n1406 , pi071 , pi164 );
  nand g01030 ( new_n1407 , pi142 , pi206 );
  xor  g01031 ( new_n1408 , new_n1406 , new_n1407 );
  not  g01032 ( new_n1409 , new_n1408 );
  nand g01033 ( new_n1410 , pi026 , pi087 );
  nand g01034 ( new_n1411 , pi027 , pi219 );
  nand g01035 ( new_n1412 , new_n1410 , new_n1411 );
  nand g01036 ( new_n1413 , new_n1392 , new_n1412 );
  nand g01037 ( new_n1414 , new_n1409 , new_n1413 );
  nor  g01038 ( new_n1415 , new_n1055 , new_n1056 );
  xor  g01039 ( new_n1416 , new_n1408 , new_n1413 );
  or   g01040 ( new_n1417 , new_n1415 , new_n1416 );
  nand g01041 ( new_n1418 , new_n1414 , new_n1417 );
  nor  g01042 ( new_n1419 , new_n1374 , new_n1375 );
  nor  g01043 ( new_n1420 , new_n1377 , new_n1419 );
  not  g01044 ( new_n1421 , new_n1420 );
  nand g01045 ( new_n1422 , new_n1418 , new_n1421 );
  xor  g01046 ( new_n1423 , new_n1390 , new_n1391 );
  xor  g01047 ( new_n1424 , new_n1418 , new_n1421 );
  nand g01048 ( new_n1425 , new_n1423 , new_n1424 );
  nand g01049 ( new_n1426 , new_n1422 , new_n1425 );
  nand g01050 ( new_n1427 , new_n1405 , new_n1426 );
  xor  g01051 ( new_n1428 , new_n1372 , new_n1378 );
  not  g01052 ( new_n1429 , new_n1428 );
  xor  g01053 ( new_n1430 , new_n1405 , new_n1426 );
  nand g01054 ( new_n1431 , new_n1429 , new_n1430 );
  nand g01055 ( new_n1432 , new_n1427 , new_n1431 );
  nand g01056 ( new_n1433 , new_n1385 , new_n1432 );
  not  g01057 ( new_n1434 , new_n1393 );
  nor  g01058 ( new_n1435 , new_n1434 , new_n1404 );
  nand g01059 ( new_n1436 , pi008 , pi102 );
  nand g01060 ( new_n1437 , pi001 , pi026 );
  nand g01061 ( new_n1438 , pi027 , pi122 );
  xor  g01062 ( new_n1439 , new_n1437 , new_n1438 );
  xor  g01063 ( new_n1440 , new_n1436 , new_n1439 );
  nand g01064 ( new_n1441 , pi056 , pi219 );
  nand g01065 ( new_n1442 , new_n1400 , new_n1401 );
  nand g01066 ( new_n1443 , new_n1399 , new_n1402 );
  nand g01067 ( new_n1444 , new_n1442 , new_n1443 );
  xor  g01068 ( new_n1445 , new_n1441 , new_n1444 );
  xor  g01069 ( new_n1446 , new_n1440 , new_n1445 );
  nand g01070 ( new_n1447 , pi087 , pi136 );
  xor  g01071 ( new_n1448 , new_n1446 , new_n1447 );
  or   g01072 ( new_n1449 , new_n1394 , new_n1397 );
  nand g01073 ( new_n1450 , new_n1398 , new_n1403 );
  nand g01074 ( new_n1451 , new_n1449 , new_n1450 );
  xor  g01075 ( new_n1452 , new_n1448 , new_n1451 );
  xnor g01076 ( new_n1453 , new_n1435 , new_n1452 );
  xor  g01077 ( new_n1454 , new_n1385 , new_n1432 );
  nand g01078 ( new_n1455 , new_n1453 , new_n1454 );
  nand g01079 ( new_n1456 , new_n1433 , new_n1455 );
  nand g01080 ( new_n1457 , pi001 , pi008 );
  nand g01081 ( new_n1458 , pi026 , pi122 );
  nand g01082 ( new_n1459 , pi027 , pi135 );
  nand g01083 ( new_n1460 , new_n1458 , new_n1459 );
  nand g01084 ( new_n1461 , pi026 , pi135 );
  or   g01085 ( new_n1462 , new_n1438 , new_n1461 );
  nand g01086 ( new_n1463 , new_n1460 , new_n1462 );
  xor  g01087 ( new_n1464 , new_n1457 , new_n1463 );
  nand g01088 ( new_n1465 , new_n1437 , new_n1438 );
  nand g01089 ( new_n1466 , new_n1436 , new_n1439 );
  nand g01090 ( new_n1467 , new_n1465 , new_n1466 );
  xor  g01091 ( new_n1468 , new_n1464 , new_n1467 );
  nand g01092 ( new_n1469 , pi056 , pi102 );
  nand g01093 ( new_n1470 , pi136 , pi219 );
  and  g01094 ( new_n1471 , new_n1469 , new_n1470 );
  nand g01095 ( new_n1472 , pi102 , pi136 );
  nor  g01096 ( new_n1473 , new_n1441 , new_n1472 );
  or   g01097 ( new_n1474 , new_n1471 , new_n1473 );
  xnor g01098 ( new_n1475 , new_n1468 , new_n1474 );
  nand g01099 ( new_n1476 , new_n1441 , new_n1444 );
  nand g01100 ( new_n1477 , new_n1440 , new_n1445 );
  nand g01101 ( new_n1478 , new_n1476 , new_n1477 );
  xor  g01102 ( new_n1479 , new_n1475 , new_n1478 );
  or   g01103 ( new_n1480 , new_n1446 , new_n1447 );
  nand g01104 ( new_n1481 , new_n1448 , new_n1451 );
  nand g01105 ( new_n1482 , new_n1480 , new_n1481 );
  xnor g01106 ( new_n1483 , new_n1479 , new_n1482 );
  nand g01107 ( new_n1484 , new_n1435 , new_n1452 );
  nand g01108 ( new_n1485 , pi087 , pi096 );
  xor  g01109 ( new_n1486 , new_n1484 , new_n1485 );
  xor  g01110 ( new_n1487 , new_n1483 , new_n1486 );
  xor  g01111 ( new_n1488 , new_n1456 , new_n1487 );
  xor  g01112 ( new_n1489 , new_n1384 , new_n1488 );
  xor  g01113 ( new_n1490 , new_n1309 , new_n1310 );
  or   g01114 ( new_n1491 , new_n1489 , new_n1490 );
  xor  g01115 ( new_n1492 , new_n1453 , new_n1454 );
  not  g01116 ( new_n1493 , new_n1492 );
  xor  g01117 ( new_n1494 , new_n1304 , new_n1305 );
  nor  g01118 ( new_n1495 , new_n1493 , new_n1494 );
  xor  g01119 ( new_n1496 , new_n1492 , new_n1494 );
  xor  g01120 ( new_n1497 , new_n1302 , new_n1303 );
  xor  g01121 ( new_n1498 , new_n1300 , new_n1301 );
  not  g01122 ( new_n1499 , new_n1057 );
  or   g01123 ( new_n1500 , new_n1499 , new_n1058 );
  nand g01124 ( new_n1501 , pi138 , pi151 );
  nand g01125 ( new_n1502 , pi147 , pi182 );
  nand g01126 ( new_n1503 , new_n1501 , new_n1502 );
  nand g01127 ( new_n1504 , new_n1301 , new_n1503 );
  or   g01128 ( new_n1505 , new_n1500 , new_n1504 );
  xor  g01129 ( new_n1506 , new_n1415 , new_n1416 );
  not  g01130 ( new_n1507 , new_n1506 );
  xor  g01131 ( new_n1508 , new_n1500 , new_n1504 );
  nand g01132 ( new_n1509 , new_n1507 , new_n1508 );
  nand g01133 ( new_n1510 , new_n1505 , new_n1509 );
  nand g01134 ( new_n1511 , new_n1498 , new_n1510 );
  xnor g01135 ( new_n1512 , new_n1423 , new_n1424 );
  xor  g01136 ( new_n1513 , new_n1498 , new_n1510 );
  nand g01137 ( new_n1514 , new_n1512 , new_n1513 );
  nand g01138 ( new_n1515 , new_n1511 , new_n1514 );
  nand g01139 ( new_n1516 , new_n1497 , new_n1515 );
  xor  g01140 ( new_n1517 , new_n1428 , new_n1430 );
  xor  g01141 ( new_n1518 , new_n1497 , new_n1515 );
  nand g01142 ( new_n1519 , new_n1517 , new_n1518 );
  nand g01143 ( new_n1520 , new_n1516 , new_n1519 );
  nor  g01144 ( new_n1521 , new_n1496 , new_n1520 );
  nor  g01145 ( new_n1522 , new_n1495 , new_n1521 );
  xor  g01146 ( new_n1523 , new_n1489 , new_n1490 );
  nand g01147 ( new_n1524 , new_n1522 , new_n1523 );
  nand g01148 ( new_n1525 , new_n1491 , new_n1524 );
  or   g01149 ( new_n1526 , new_n1313 , new_n1525 );
  nand g01150 ( new_n1527 , new_n1381 , new_n1382 );
  nand g01151 ( new_n1528 , new_n1371 , new_n1383 );
  nand g01152 ( new_n1529 , new_n1527 , new_n1528 );
  nand g01153 ( new_n1530 , new_n1351 , new_n1370 );
  nand g01154 ( new_n1531 , pi032 , pi099 );
  nand g01155 ( new_n1532 , pi155 , pi164 );
  xor  g01156 ( new_n1533 , new_n1339 , new_n1532 );
  xor  g01157 ( new_n1534 , new_n1531 , new_n1533 );
  nand g01158 ( new_n1535 , pi123 , pi145 );
  xor  g01159 ( new_n1536 , new_n1341 , new_n1535 );
  not  g01160 ( new_n1537 , new_n1536 );
  xor  g01161 ( new_n1538 , new_n1534 , new_n1537 );
  nand g01162 ( new_n1539 , pi071 , pi114 );
  nand g01163 ( new_n1540 , pi091 , pi142 );
  xor  g01164 ( new_n1541 , new_n1539 , new_n1540 );
  xor  g01165 ( new_n1542 , new_n1347 , new_n1541 );
  nand g01166 ( new_n1543 , new_n1331 , new_n1334 );
  nand g01167 ( new_n1544 , new_n1335 , new_n1342 );
  nand g01168 ( new_n1545 , new_n1543 , new_n1544 );
  xor  g01169 ( new_n1546 , new_n1542 , new_n1545 );
  xor  g01170 ( new_n1547 , new_n1538 , new_n1546 );
  nand g01171 ( new_n1548 , new_n1343 , new_n1349 );
  nand g01172 ( new_n1549 , new_n1330 , new_n1350 );
  nand g01173 ( new_n1550 , new_n1548 , new_n1549 );
  xor  g01174 ( new_n1551 , new_n1348 , new_n1550 );
  xnor g01175 ( new_n1552 , new_n1547 , new_n1551 );
  xnor g01176 ( new_n1553 , new_n1530 , new_n1552 );
  xor  g01177 ( new_n1554 , new_n1529 , new_n1553 );
  nand g01178 ( new_n1555 , new_n1484 , new_n1485 );
  nand g01179 ( new_n1556 , new_n1483 , new_n1486 );
  nand g01180 ( new_n1557 , new_n1555 , new_n1556 );
  nand g01181 ( new_n1558 , new_n1479 , new_n1482 );
  nand g01182 ( new_n1559 , pi008 , pi122 );
  nand g01183 ( new_n1560 , pi027 , pi059 );
  xor  g01184 ( new_n1561 , new_n1559 , new_n1560 );
  xor  g01185 ( new_n1562 , new_n1461 , new_n1561 );
  not  g01186 ( new_n1563 , new_n1562 );
  nand g01187 ( new_n1564 , pi001 , pi056 );
  xor  g01188 ( new_n1565 , new_n1462 , new_n1564 );
  xor  g01189 ( new_n1566 , new_n1563 , new_n1565 );
  nand g01190 ( new_n1567 , pi087 , pi235 );
  nand g01191 ( new_n1568 , pi096 , pi219 );
  xor  g01192 ( new_n1569 , new_n1472 , new_n1568 );
  xor  g01193 ( new_n1570 , new_n1567 , new_n1569 );
  nand g01194 ( new_n1571 , new_n1457 , new_n1463 );
  nand g01195 ( new_n1572 , new_n1464 , new_n1467 );
  nand g01196 ( new_n1573 , new_n1571 , new_n1572 );
  xor  g01197 ( new_n1574 , new_n1570 , new_n1573 );
  xor  g01198 ( new_n1575 , new_n1566 , new_n1574 );
  nor  g01199 ( new_n1576 , new_n1468 , new_n1474 );
  nor  g01200 ( new_n1577 , new_n1475 , new_n1478 );
  xor  g01201 ( new_n1578 , new_n1473 , new_n1577 );
  nor  g01202 ( new_n1579 , new_n1576 , new_n1578 );
  xor  g01203 ( new_n1580 , new_n1575 , new_n1579 );
  xor  g01204 ( new_n1581 , new_n1558 , new_n1580 );
  xor  g01205 ( new_n1582 , new_n1557 , new_n1581 );
  nand g01206 ( new_n1583 , new_n1456 , new_n1487 );
  nand g01207 ( new_n1584 , new_n1384 , new_n1488 );
  nand g01208 ( new_n1585 , new_n1583 , new_n1584 );
  xor  g01209 ( new_n1586 , new_n1582 , new_n1585 );
  xor  g01210 ( new_n1587 , new_n1554 , new_n1586 );
  not  g01211 ( new_n1588 , new_n1587 );
  xor  g01212 ( new_n1589 , new_n1313 , new_n1525 );
  nand g01213 ( new_n1590 , new_n1588 , new_n1589 );
  nand g01214 ( new_n1591 , new_n1526 , new_n1590 );
  xor  g01215 ( new_n1592 , new_n1216 , new_n1591 );
  nor  g01216 ( new_n1593 , new_n1275 , new_n1298 );
  nor  g01217 ( new_n1594 , new_n1299 , new_n1312 );
  nor  g01218 ( new_n1595 , new_n1593 , new_n1594 );
  nand g01219 ( new_n1596 , pi119 , pi137 );
  nand g01220 ( new_n1597 , pi009 , pi160 );
  xor  g01221 ( new_n1598 , new_n1596 , new_n1597 );
  nand g01222 ( new_n1599 , pi020 , pi044 );
  nand g01223 ( new_n1600 , pi054 , pi060 );
  or   g01224 ( new_n1601 , new_n1599 , new_n1600 );
  nand g01225 ( new_n1602 , pi045 , pi060 );
  nand g01226 ( new_n1603 , pi119 , pi223 );
  nand g01227 ( new_n1604 , new_n1602 , new_n1603 );
  nand g01228 ( new_n1605 , pi020 , pi250 );
  xor  g01229 ( new_n1606 , new_n1602 , new_n1603 );
  nand g01230 ( new_n1607 , new_n1605 , new_n1606 );
  nand g01231 ( new_n1608 , new_n1604 , new_n1607 );
  nand g01232 ( new_n1609 , new_n1599 , new_n1608 );
  nand g01233 ( new_n1610 , pi045 , pi223 );
  nand g01234 ( new_n1611 , pi060 , pi250 );
  nand g01235 ( new_n1612 , pi101 , pi119 );
  xor  g01236 ( new_n1613 , new_n1611 , new_n1612 );
  xor  g01237 ( new_n1614 , new_n1610 , new_n1613 );
  xor  g01238 ( new_n1615 , new_n1599 , new_n1608 );
  nand g01239 ( new_n1616 , new_n1614 , new_n1615 );
  nand g01240 ( new_n1617 , new_n1609 , new_n1616 );
  nand g01241 ( new_n1618 , pi044 , pi060 );
  nand g01242 ( new_n1619 , pi020 , pi054 );
  nand g01243 ( new_n1620 , new_n1618 , new_n1619 );
  nand g01244 ( new_n1621 , new_n1601 , new_n1620 );
  nand g01245 ( new_n1622 , new_n1617 , new_n1621 );
  nand g01246 ( new_n1623 , pi223 , pi250 );
  nand g01247 ( new_n1624 , new_n1611 , new_n1612 );
  nand g01248 ( new_n1625 , new_n1610 , new_n1613 );
  nand g01249 ( new_n1626 , new_n1624 , new_n1625 );
  nand g01250 ( new_n1627 , pi119 , pi225 );
  nand g01251 ( new_n1628 , pi045 , pi101 );
  nand g01252 ( new_n1629 , new_n1627 , new_n1628 );
  nand g01253 ( new_n1630 , pi045 , pi225 );
  or   g01254 ( new_n1631 , new_n1612 , new_n1630 );
  nand g01255 ( new_n1632 , new_n1629 , new_n1631 );
  xor  g01256 ( new_n1633 , new_n1626 , new_n1632 );
  xor  g01257 ( new_n1634 , new_n1623 , new_n1633 );
  xor  g01258 ( new_n1635 , new_n1617 , new_n1621 );
  nand g01259 ( new_n1636 , new_n1634 , new_n1635 );
  nand g01260 ( new_n1637 , new_n1622 , new_n1636 );
  or   g01261 ( new_n1638 , new_n1601 , new_n1637 );
  xor  g01262 ( new_n1639 , new_n1601 , new_n1637 );
  nand g01263 ( new_n1640 , pi101 , pi250 );
  nand g01264 ( new_n1641 , pi119 , pi177 );
  xor  g01265 ( new_n1642 , new_n1630 , new_n1641 );
  xor  g01266 ( new_n1643 , new_n1640 , new_n1642 );
  nand g01267 ( new_n1644 , pi044 , pi223 );
  xor  g01268 ( new_n1645 , new_n1631 , new_n1644 );
  not  g01269 ( new_n1646 , new_n1645 );
  xor  g01270 ( new_n1647 , new_n1643 , new_n1646 );
  nand g01271 ( new_n1648 , pi160 , pi248 );
  nand g01272 ( new_n1649 , pi020 , pi072 );
  xor  g01273 ( new_n1650 , new_n1648 , new_n1649 );
  xor  g01274 ( new_n1651 , new_n1600 , new_n1650 );
  nand g01275 ( new_n1652 , new_n1626 , new_n1632 );
  nand g01276 ( new_n1653 , new_n1623 , new_n1633 );
  nand g01277 ( new_n1654 , new_n1652 , new_n1653 );
  xor  g01278 ( new_n1655 , new_n1651 , new_n1654 );
  xor  g01279 ( new_n1656 , new_n1647 , new_n1655 );
  nand g01280 ( new_n1657 , new_n1639 , new_n1656 );
  nand g01281 ( new_n1658 , new_n1638 , new_n1657 );
  xor  g01282 ( new_n1659 , new_n1634 , new_n1635 );
  not  g01283 ( new_n1660 , new_n1659 );
  xor  g01284 ( new_n1661 , new_n1614 , new_n1615 );
  nand g01285 ( new_n1662 , pi054 , pi160 );
  or   g01286 ( new_n1663 , new_n1661 , new_n1662 );
  xor  g01287 ( new_n1664 , new_n1661 , new_n1662 );
  nand g01288 ( new_n1665 , pi060 , pi119 );
  nand g01289 ( new_n1666 , pi160 , pi250 );
  nand g01290 ( new_n1667 , new_n1665 , new_n1666 );
  nand g01291 ( new_n1668 , pi020 , pi045 );
  or   g01292 ( new_n1669 , new_n1665 , new_n1666 );
  nand g01293 ( new_n1670 , new_n1668 , new_n1669 );
  nand g01294 ( new_n1671 , new_n1667 , new_n1670 );
  nand g01295 ( new_n1672 , pi044 , pi160 );
  or   g01296 ( new_n1673 , new_n1671 , new_n1672 );
  xor  g01297 ( new_n1674 , new_n1605 , new_n1606 );
  not  g01298 ( new_n1675 , new_n1674 );
  xor  g01299 ( new_n1676 , new_n1671 , new_n1672 );
  nand g01300 ( new_n1677 , new_n1675 , new_n1676 );
  nand g01301 ( new_n1678 , new_n1673 , new_n1677 );
  nand g01302 ( new_n1679 , new_n1664 , new_n1678 );
  nand g01303 ( new_n1680 , new_n1663 , new_n1679 );
  nand g01304 ( new_n1681 , new_n1660 , new_n1680 );
  xnor g01305 ( new_n1682 , new_n1639 , new_n1656 );
  nor  g01306 ( new_n1683 , new_n1681 , new_n1682 );
  xor  g01307 ( new_n1684 , new_n1674 , new_n1676 );
  not  g01308 ( new_n1685 , new_n1668 );
  not  g01309 ( new_n1686 , new_n1667 );
  nand g01310 ( new_n1687 , new_n1060 , new_n1685 );
  nand g01311 ( new_n1688 , new_n1686 , new_n1687 );
  nand g01312 ( new_n1689 , new_n1669 , new_n1688 );
  nand g01313 ( new_n1690 , new_n1685 , new_n1689 );
  nor  g01314 ( new_n1691 , new_n1684 , new_n1690 );
  xor  g01315 ( new_n1692 , new_n1664 , new_n1678 );
  nand g01316 ( new_n1693 , new_n1691 , new_n1692 );
  nand g01317 ( new_n1694 , pi072 , pi160 );
  nand g01318 ( new_n1695 , new_n1693 , new_n1694 );
  xor  g01319 ( new_n1696 , new_n1659 , new_n1680 );
  xor  g01320 ( new_n1697 , new_n1693 , new_n1694 );
  nand g01321 ( new_n1698 , new_n1696 , new_n1697 );
  nand g01322 ( new_n1699 , new_n1695 , new_n1698 );
  xor  g01323 ( new_n1700 , new_n1681 , new_n1682 );
  not  g01324 ( new_n1701 , new_n1700 );
  nor  g01325 ( new_n1702 , new_n1699 , new_n1701 );
  or   g01326 ( new_n1703 , new_n1683 , new_n1702 );
  xor  g01327 ( new_n1704 , new_n1658 , new_n1703 );
  xor  g01328 ( new_n1705 , new_n1598 , new_n1704 );
  nand g01329 ( new_n1706 , pi096 , pi102 );
  nand g01330 ( new_n1707 , pi219 , pi235 );
  or   g01331 ( new_n1708 , new_n1462 , new_n1564 );
  nand g01332 ( new_n1709 , new_n1563 , new_n1565 );
  nand g01333 ( new_n1710 , new_n1708 , new_n1709 );
  xor  g01334 ( new_n1711 , new_n1707 , new_n1710 );
  xor  g01335 ( new_n1712 , new_n1706 , new_n1711 );
  xor  g01336 ( new_n1713 , new_n1705 , new_n1712 );
  nand g01337 ( new_n1714 , pi087 , pi110 );
  nand g01338 ( new_n1715 , pi027 , pi094 );
  nand g01339 ( new_n1716 , pi026 , pi059 );
  nand g01340 ( new_n1717 , pi008 , pi135 );
  xor  g01341 ( new_n1718 , new_n1716 , new_n1717 );
  nand g01342 ( new_n1719 , new_n1473 , new_n1577 );
  not  g01343 ( new_n1720 , new_n1579 );
  nand g01344 ( new_n1721 , new_n1575 , new_n1720 );
  nand g01345 ( new_n1722 , new_n1719 , new_n1721 );
  nand g01346 ( new_n1723 , new_n1539 , new_n1540 );
  nand g01347 ( new_n1724 , new_n1347 , new_n1541 );
  nand g01348 ( new_n1725 , new_n1723 , new_n1724 );
  xor  g01349 ( new_n1726 , new_n1722 , new_n1725 );
  nand g01350 ( new_n1727 , pi071 , pi091 );
  nand g01351 ( new_n1728 , pi114 , pi169 );
  xnor g01352 ( new_n1729 , new_n1727 , new_n1728 );
  nand g01353 ( new_n1730 , pi099 , pi145 );
  xor  g01354 ( new_n1731 , new_n1729 , new_n1730 );
  nand g01355 ( new_n1732 , new_n1542 , new_n1545 );
  not  g01356 ( new_n1733 , new_n1538 );
  nand g01357 ( new_n1734 , new_n1733 , new_n1546 );
  nand g01358 ( new_n1735 , new_n1732 , new_n1734 );
  nand g01359 ( new_n1736 , pi123 , pi246 );
  xor  g01360 ( new_n1737 , new_n1735 , new_n1736 );
  xor  g01361 ( new_n1738 , new_n1731 , new_n1737 );
  nand g01362 ( new_n1739 , new_n1339 , new_n1532 );
  nand g01363 ( new_n1740 , new_n1531 , new_n1533 );
  nand g01364 ( new_n1741 , new_n1739 , new_n1740 );
  nor  g01365 ( new_n1742 , new_n1341 , new_n1535 );
  nor  g01366 ( new_n1743 , new_n1534 , new_n1537 );
  or   g01367 ( new_n1744 , new_n1742 , new_n1743 );
  xor  g01368 ( new_n1745 , new_n1741 , new_n1744 );
  xor  g01369 ( new_n1746 , new_n1738 , new_n1745 );
  xor  g01370 ( new_n1747 , new_n1726 , new_n1746 );
  xor  g01371 ( new_n1748 , new_n1718 , new_n1747 );
  xor  g01372 ( new_n1749 , new_n1715 , new_n1748 );
  xor  g01373 ( new_n1750 , new_n1714 , new_n1749 );
  nand g01374 ( new_n1751 , new_n1472 , new_n1568 );
  nand g01375 ( new_n1752 , new_n1567 , new_n1569 );
  nand g01376 ( new_n1753 , new_n1751 , new_n1752 );
  nand g01377 ( new_n1754 , new_n1558 , new_n1580 );
  nand g01378 ( new_n1755 , new_n1557 , new_n1581 );
  nand g01379 ( new_n1756 , new_n1754 , new_n1755 );
  nand g01380 ( new_n1757 , pi056 , pi122 );
  nand g01381 ( new_n1758 , pi001 , pi136 );
  xor  g01382 ( new_n1759 , new_n1757 , new_n1758 );
  xor  g01383 ( new_n1760 , new_n1756 , new_n1759 );
  xor  g01384 ( new_n1761 , new_n1753 , new_n1760 );
  xor  g01385 ( new_n1762 , new_n1750 , new_n1761 );
  nand g01386 ( new_n1763 , new_n1570 , new_n1573 );
  not  g01387 ( new_n1764 , new_n1566 );
  nand g01388 ( new_n1765 , new_n1764 , new_n1574 );
  nand g01389 ( new_n1766 , new_n1763 , new_n1765 );
  nand g01390 ( new_n1767 , new_n1559 , new_n1560 );
  nand g01391 ( new_n1768 , new_n1461 , new_n1561 );
  nand g01392 ( new_n1769 , new_n1767 , new_n1768 );
  xor  g01393 ( new_n1770 , new_n1766 , new_n1769 );
  xor  g01394 ( new_n1771 , new_n1762 , new_n1770 );
  xor  g01395 ( new_n1772 , new_n1713 , new_n1771 );
  nand g01396 ( new_n1773 , new_n1630 , new_n1641 );
  nand g01397 ( new_n1774 , new_n1640 , new_n1642 );
  nand g01398 ( new_n1775 , new_n1773 , new_n1774 );
  nor  g01399 ( new_n1776 , new_n1631 , new_n1644 );
  nor  g01400 ( new_n1777 , new_n1643 , new_n1646 );
  or   g01401 ( new_n1778 , new_n1776 , new_n1777 );
  xor  g01402 ( new_n1779 , new_n1775 , new_n1778 );
  xor  g01403 ( new_n1780 , new_n1772 , new_n1779 );
  xor  g01404 ( new_n1781 , new_n1595 , new_n1780 );
  xor  g01405 ( new_n1782 , new_n1592 , new_n1781 );
  nand g01406 ( new_n1783 , pi151 , pi251 );
  nand g01407 ( new_n1784 , new_n1648 , new_n1649 );
  nand g01408 ( new_n1785 , new_n1600 , new_n1650 );
  nand g01409 ( new_n1786 , new_n1784 , new_n1785 );
  or   g01410 ( new_n1787 , new_n1651 , new_n1654 );
  nand g01411 ( new_n1788 , new_n1647 , new_n1655 );
  nand g01412 ( new_n1789 , new_n1787 , new_n1788 );
  xor  g01413 ( new_n1790 , new_n1786 , new_n1789 );
  xor  g01414 ( new_n1791 , new_n1783 , new_n1790 );
  xor  g01415 ( new_n1792 , new_n1699 , new_n1700 );
  xnor g01416 ( new_n1793 , new_n1691 , new_n1692 );
  xor  g01417 ( new_n1794 , new_n1684 , new_n1690 );
  xnor g01418 ( new_n1795 , new_n1512 , new_n1513 );
  nor  g01419 ( new_n1796 , new_n1059 , new_n1060 );
  nand g01420 ( new_n1797 , pi045 , pi160 );
  nand g01421 ( new_n1798 , pi020 , pi119 );
  xor  g01422 ( new_n1799 , new_n1797 , new_n1798 );
  or   g01423 ( new_n1800 , new_n1796 , new_n1799 );
  xor  g01424 ( new_n1801 , new_n1507 , new_n1508 );
  not  g01425 ( new_n1802 , new_n1801 );
  xor  g01426 ( new_n1803 , new_n1796 , new_n1799 );
  nand g01427 ( new_n1804 , new_n1802 , new_n1803 );
  nand g01428 ( new_n1805 , new_n1800 , new_n1804 );
  or   g01429 ( new_n1806 , new_n1795 , new_n1805 );
  xor  g01430 ( new_n1807 , new_n1795 , new_n1805 );
  nor  g01431 ( new_n1808 , new_n1686 , new_n1687 );
  nor  g01432 ( new_n1809 , new_n1689 , new_n1808 );
  nand g01433 ( new_n1810 , new_n1807 , new_n1809 );
  nand g01434 ( new_n1811 , new_n1806 , new_n1810 );
  or   g01435 ( new_n1812 , new_n1794 , new_n1811 );
  xor  g01436 ( new_n1813 , new_n1517 , new_n1518 );
  not  g01437 ( new_n1814 , new_n1813 );
  xor  g01438 ( new_n1815 , new_n1794 , new_n1811 );
  nand g01439 ( new_n1816 , new_n1814 , new_n1815 );
  nand g01440 ( new_n1817 , new_n1812 , new_n1816 );
  or   g01441 ( new_n1818 , new_n1793 , new_n1817 );
  xnor g01442 ( new_n1819 , new_n1496 , new_n1520 );
  xor  g01443 ( new_n1820 , new_n1793 , new_n1817 );
  nand g01444 ( new_n1821 , new_n1819 , new_n1820 );
  nand g01445 ( new_n1822 , new_n1818 , new_n1821 );
  xnor g01446 ( new_n1823 , new_n1696 , new_n1697 );
  or   g01447 ( new_n1824 , new_n1822 , new_n1823 );
  xor  g01448 ( new_n1825 , new_n1522 , new_n1523 );
  not  g01449 ( new_n1826 , new_n1825 );
  xor  g01450 ( new_n1827 , new_n1822 , new_n1823 );
  nand g01451 ( new_n1828 , new_n1826 , new_n1827 );
  nand g01452 ( new_n1829 , new_n1824 , new_n1828 );
  or   g01453 ( new_n1830 , new_n1792 , new_n1829 );
  xor  g01454 ( new_n1831 , new_n1587 , new_n1589 );
  xor  g01455 ( new_n1832 , new_n1792 , new_n1829 );
  nand g01456 ( new_n1833 , new_n1831 , new_n1832 );
  nand g01457 ( new_n1834 , new_n1830 , new_n1833 );
  nand g01458 ( new_n1835 , pi011 , pi138 );
  xor  g01459 ( new_n1836 , new_n1834 , new_n1835 );
  xor  g01460 ( new_n1837 , new_n1791 , new_n1836 );
  nor  g01461 ( new_n1838 , new_n1291 , new_n1297 );
  nor  g01462 ( new_n1839 , new_n1296 , new_n1838 );
  nand g01463 ( new_n1840 , pi045 , pi177 );
  nand g01464 ( new_n1841 , pi044 , pi101 );
  xor  g01465 ( new_n1842 , new_n1840 , new_n1841 );
  nand g01466 ( new_n1843 , pi054 , pi223 );
  or   g01467 ( new_n1844 , new_n1582 , new_n1585 );
  nand g01468 ( new_n1845 , new_n1554 , new_n1586 );
  nand g01469 ( new_n1846 , new_n1844 , new_n1845 );
  nand g01470 ( new_n1847 , pi075 , pi216 );
  nand g01471 ( new_n1848 , pi041 , pi093 );
  xor  g01472 ( new_n1849 , new_n1847 , new_n1848 );
  nand g01473 ( new_n1850 , pi076 , pi097 );
  nand g01474 ( new_n1851 , new_n1286 , new_n1289 );
  nand g01475 ( new_n1852 , new_n1282 , new_n1290 );
  nand g01476 ( new_n1853 , new_n1851 , new_n1852 );
  xor  g01477 ( new_n1854 , new_n1850 , new_n1853 );
  xor  g01478 ( new_n1855 , new_n1849 , new_n1854 );
  xor  g01479 ( new_n1856 , new_n1846 , new_n1855 );
  or   g01480 ( new_n1857 , new_n1348 , new_n1550 );
  nand g01481 ( new_n1858 , new_n1547 , new_n1551 );
  nand g01482 ( new_n1859 , new_n1857 , new_n1858 );
  nand g01483 ( new_n1860 , pi086 , pi164 );
  nand g01484 ( new_n1861 , new_n1283 , new_n1284 );
  nand g01485 ( new_n1862 , new_n1237 , new_n1285 );
  nand g01486 ( new_n1863 , new_n1861 , new_n1862 );
  nand g01487 ( new_n1864 , pi155 , pi206 );
  nand g01488 ( new_n1865 , pi023 , pi032 );
  xor  g01489 ( new_n1866 , new_n1864 , new_n1865 );
  xor  g01490 ( new_n1867 , new_n1863 , new_n1866 );
  xor  g01491 ( new_n1868 , new_n1860 , new_n1867 );
  xor  g01492 ( new_n1869 , new_n1859 , new_n1868 );
  nand g01493 ( new_n1870 , new_n1276 , new_n1277 );
  nand g01494 ( new_n1871 , new_n1228 , new_n1278 );
  nand g01495 ( new_n1872 , new_n1870 , new_n1871 );
  or   g01496 ( new_n1873 , new_n1229 , new_n1280 );
  not  g01497 ( new_n1874 , new_n1279 );
  nand g01498 ( new_n1875 , new_n1874 , new_n1281 );
  nand g01499 ( new_n1876 , new_n1873 , new_n1875 );
  xor  g01500 ( new_n1877 , new_n1872 , new_n1876 );
  nor  g01501 ( new_n1878 , new_n1530 , new_n1552 );
  nor  g01502 ( new_n1879 , new_n1529 , new_n1553 );
  nor  g01503 ( new_n1880 , new_n1878 , new_n1879 );
  nand g01504 ( new_n1881 , pi031 , pi142 );
  xor  g01505 ( new_n1882 , new_n1880 , new_n1881 );
  xor  g01506 ( new_n1883 , new_n1877 , new_n1882 );
  xor  g01507 ( new_n1884 , new_n1869 , new_n1883 );
  nand g01508 ( new_n1885 , pi166 , pi182 );
  nand g01509 ( new_n1886 , pi019 , pi079 );
  xor  g01510 ( new_n1887 , new_n1885 , new_n1886 );
  xor  g01511 ( new_n1888 , new_n1884 , new_n1887 );
  xor  g01512 ( new_n1889 , new_n1856 , new_n1888 );
  xor  g01513 ( new_n1890 , new_n1843 , new_n1889 );
  xor  g01514 ( new_n1891 , new_n1842 , new_n1890 );
  nand g01515 ( new_n1892 , pi225 , pi250 );
  nand g01516 ( new_n1893 , pi020 , pi248 );
  nand g01517 ( new_n1894 , pi060 , pi072 );
  xor  g01518 ( new_n1895 , new_n1893 , new_n1894 );
  xor  g01519 ( new_n1896 , new_n1892 , new_n1895 );
  xor  g01520 ( new_n1897 , new_n1891 , new_n1896 );
  xor  g01521 ( new_n1898 , new_n1839 , new_n1897 );
  xor  g01522 ( new_n1899 , new_n1837 , new_n1898 );
  xor  g01523 ( po005 , new_n1782 , new_n1899 );
  nand g01524 ( new_n1901 , pi067 , pi117 );
  nand g01525 ( new_n1902 , pi016 , pi053 );
  nor  g01526 ( new_n1903 , new_n1901 , new_n1902 );
  nand g01527 ( new_n1904 , pi080 , pi229 );
  nand g01528 ( new_n1905 , pi080 , pi092 );
  nand g01529 ( new_n1906 , pi016 , pi229 );
  nand g01530 ( new_n1907 , new_n1905 , new_n1906 );
  nand g01531 ( new_n1908 , pi190 , pi247 );
  xor  g01532 ( new_n1909 , new_n1905 , new_n1906 );
  nand g01533 ( new_n1910 , new_n1908 , new_n1909 );
  nand g01534 ( new_n1911 , new_n1907 , new_n1910 );
  xor  g01535 ( new_n1912 , new_n1904 , new_n1911 );
  nand g01536 ( new_n1913 , pi190 , pi234 );
  nand g01537 ( new_n1914 , pi092 , pi247 );
  nand g01538 ( new_n1915 , new_n1913 , new_n1914 );
  nand g01539 ( new_n1916 , pi092 , pi234 );
  or   g01540 ( new_n1917 , new_n1908 , new_n1916 );
  nand g01541 ( new_n1918 , new_n1915 , new_n1917 );
  xor  g01542 ( new_n1919 , new_n1912 , new_n1918 );
  nand g01543 ( new_n1920 , pi016 , pi067 );
  nand g01544 ( new_n1921 , pi053 , pi117 );
  and  g01545 ( new_n1922 , new_n1920 , new_n1921 );
  or   g01546 ( new_n1923 , new_n1903 , new_n1922 );
  xnor g01547 ( new_n1924 , new_n1919 , new_n1923 );
  nand g01548 ( new_n1925 , pi016 , pi092 );
  nand g01549 ( new_n1926 , pi080 , pi190 );
  nand g01550 ( new_n1927 , new_n1925 , new_n1926 );
  nand g01551 ( new_n1928 , pi117 , pi229 );
  xor  g01552 ( new_n1929 , new_n1925 , new_n1926 );
  nand g01553 ( new_n1930 , new_n1928 , new_n1929 );
  nand g01554 ( new_n1931 , new_n1927 , new_n1930 );
  nand g01555 ( new_n1932 , new_n1901 , new_n1931 );
  xor  g01556 ( new_n1933 , new_n1908 , new_n1909 );
  xor  g01557 ( new_n1934 , new_n1901 , new_n1931 );
  nand g01558 ( new_n1935 , new_n1933 , new_n1934 );
  nand g01559 ( new_n1936 , new_n1932 , new_n1935 );
  nor  g01560 ( new_n1937 , new_n1924 , new_n1936 );
  nand g01561 ( new_n1938 , new_n1903 , new_n1937 );
  nand g01562 ( new_n1939 , pi190 , pi214 );
  nand g01563 ( new_n1940 , pi229 , pi247 );
  xor  g01564 ( new_n1941 , new_n1939 , new_n1940 );
  xor  g01565 ( new_n1942 , new_n1916 , new_n1941 );
  nand g01566 ( new_n1943 , pi067 , pi080 );
  xor  g01567 ( new_n1944 , new_n1917 , new_n1943 );
  xor  g01568 ( new_n1945 , new_n1942 , new_n1944 );
  nand g01569 ( new_n1946 , pi030 , pi103 );
  nand g01570 ( new_n1947 , pi117 , pi185 );
  xor  g01571 ( new_n1948 , new_n1946 , new_n1947 );
  xor  g01572 ( new_n1949 , new_n1902 , new_n1948 );
  nand g01573 ( new_n1950 , new_n1904 , new_n1911 );
  nand g01574 ( new_n1951 , new_n1912 , new_n1918 );
  nand g01575 ( new_n1952 , new_n1950 , new_n1951 );
  xor  g01576 ( new_n1953 , new_n1949 , new_n1952 );
  xnor g01577 ( new_n1954 , new_n1945 , new_n1953 );
  nor  g01578 ( new_n1955 , new_n1919 , new_n1923 );
  xor  g01579 ( new_n1956 , new_n1903 , new_n1937 );
  nor  g01580 ( new_n1957 , new_n1955 , new_n1956 );
  not  g01581 ( new_n1958 , new_n1957 );
  nand g01582 ( new_n1959 , new_n1954 , new_n1958 );
  nand g01583 ( new_n1960 , new_n1938 , new_n1959 );
  xor  g01584 ( new_n1961 , new_n1924 , new_n1936 );
  xor  g01585 ( new_n1962 , new_n1933 , new_n1934 );
  nand g01586 ( new_n1963 , pi053 , pi103 );
  or   g01587 ( new_n1964 , new_n1962 , new_n1963 );
  xor  g01588 ( new_n1965 , new_n1962 , new_n1963 );
  nand g01589 ( new_n1966 , pi067 , pi103 );
  nand g01590 ( new_n1967 , pi092 , pi117 );
  nand g01591 ( new_n1968 , pi103 , pi229 );
  nand g01592 ( new_n1969 , new_n1967 , new_n1968 );
  xor  g01593 ( new_n1970 , new_n1967 , new_n1968 );
  nand g01594 ( new_n1971 , pi016 , pi190 );
  nand g01595 ( new_n1972 , new_n1970 , new_n1971 );
  nand g01596 ( new_n1973 , new_n1969 , new_n1972 );
  or   g01597 ( new_n1974 , new_n1966 , new_n1973 );
  xor  g01598 ( new_n1975 , new_n1966 , new_n1973 );
  xor  g01599 ( new_n1976 , new_n1928 , new_n1929 );
  not  g01600 ( new_n1977 , new_n1976 );
  nand g01601 ( new_n1978 , new_n1975 , new_n1977 );
  nand g01602 ( new_n1979 , new_n1974 , new_n1978 );
  nand g01603 ( new_n1980 , new_n1965 , new_n1979 );
  nand g01604 ( new_n1981 , new_n1964 , new_n1980 );
  nand g01605 ( new_n1982 , new_n1961 , new_n1981 );
  xor  g01606 ( new_n1983 , new_n1954 , new_n1957 );
  nand g01607 ( new_n1984 , new_n1982 , new_n1983 );
  xor  g01608 ( new_n1985 , new_n1970 , new_n1971 );
  nand g01609 ( new_n1986 , pi103 , pi190 );
  nor  g01610 ( new_n1987 , new_n1967 , new_n1986 );
  not  g01611 ( new_n1988 , new_n1987 );
  or   g01612 ( new_n1989 , new_n1985 , new_n1988 );
  xor  g01613 ( new_n1990 , new_n1975 , new_n1976 );
  nor  g01614 ( new_n1991 , new_n1989 , new_n1990 );
  xor  g01615 ( new_n1992 , new_n1965 , new_n1979 );
  nand g01616 ( new_n1993 , new_n1991 , new_n1992 );
  nand g01617 ( new_n1994 , pi103 , pi185 );
  nand g01618 ( new_n1995 , new_n1993 , new_n1994 );
  xnor g01619 ( new_n1996 , new_n1961 , new_n1981 );
  xor  g01620 ( new_n1997 , new_n1993 , new_n1994 );
  nand g01621 ( new_n1998 , new_n1996 , new_n1997 );
  nand g01622 ( new_n1999 , new_n1995 , new_n1998 );
  xor  g01623 ( new_n2000 , new_n1982 , new_n1983 );
  nand g01624 ( new_n2001 , new_n1999 , new_n2000 );
  nand g01625 ( new_n2002 , new_n1984 , new_n2001 );
  xor  g01626 ( new_n2003 , new_n1960 , new_n2002 );
  nand g01627 ( new_n2004 , pi006 , pi107 );
  nand g01628 ( new_n2005 , pi049 , pi158 );
  nand g01629 ( new_n2006 , pi245 , pi254 );
  nand g01630 ( new_n2007 , pi089 , pi171 );
  xor  g01631 ( new_n2008 , new_n2006 , new_n2007 );
  xnor g01632 ( new_n2009 , new_n2005 , new_n2008 );
  nand g01633 ( new_n2010 , pi049 , pi254 );
  nand g01634 ( new_n2011 , pi089 , pi107 );
  nand g01635 ( new_n2012 , new_n2010 , new_n2011 );
  nand g01636 ( new_n2013 , pi158 , pi171 );
  or   g01637 ( new_n2014 , new_n2010 , new_n2011 );
  nand g01638 ( new_n2015 , new_n2013 , new_n2014 );
  nand g01639 ( new_n2016 , new_n2012 , new_n2015 );
  nand g01640 ( new_n2017 , pi107 , pi154 );
  xor  g01641 ( new_n2018 , new_n2016 , new_n2017 );
  xnor g01642 ( new_n2019 , new_n2009 , new_n2018 );
  not  g01643 ( new_n2020 , new_n2013 );
  nand g01644 ( new_n2021 , pi107 , pi254 );
  nand g01645 ( new_n2022 , new_n2020 , new_n2021 );
  not  g01646 ( new_n2023 , new_n2022 );
  or   g01647 ( new_n2024 , new_n2012 , new_n2023 );
  nand g01648 ( new_n2025 , new_n2014 , new_n2024 );
  nand g01649 ( new_n2026 , new_n2020 , new_n2025 );
  nor  g01650 ( new_n2027 , new_n2019 , new_n2026 );
  nand g01651 ( new_n2028 , pi049 , pi089 );
  nand g01652 ( new_n2029 , pi158 , pi245 );
  nand g01653 ( new_n2030 , pi201 , pi254 );
  xor  g01654 ( new_n2031 , new_n2029 , new_n2030 );
  xor  g01655 ( new_n2032 , new_n2028 , new_n2031 );
  nand g01656 ( new_n2033 , pi154 , pi171 );
  nand g01657 ( new_n2034 , new_n2006 , new_n2007 );
  nand g01658 ( new_n2035 , new_n2005 , new_n2008 );
  nand g01659 ( new_n2036 , new_n2034 , new_n2035 );
  xor  g01660 ( new_n2037 , new_n2033 , new_n2036 );
  xor  g01661 ( new_n2038 , new_n2032 , new_n2037 );
  nand g01662 ( new_n2039 , pi095 , pi107 );
  or   g01663 ( new_n2040 , new_n2016 , new_n2017 );
  nand g01664 ( new_n2041 , new_n2009 , new_n2018 );
  nand g01665 ( new_n2042 , new_n2040 , new_n2041 );
  xor  g01666 ( new_n2043 , new_n2039 , new_n2042 );
  xor  g01667 ( new_n2044 , new_n2038 , new_n2043 );
  nand g01668 ( new_n2045 , new_n2027 , new_n2044 );
  nand g01669 ( new_n2046 , new_n2004 , new_n2045 );
  nand g01670 ( new_n2047 , new_n2033 , new_n2036 );
  nand g01671 ( new_n2048 , new_n2032 , new_n2037 );
  nand g01672 ( new_n2049 , new_n2047 , new_n2048 );
  nand g01673 ( new_n2050 , pi089 , pi245 );
  nand g01674 ( new_n2051 , pi156 , pi254 );
  nand g01675 ( new_n2052 , pi158 , pi201 );
  nand g01676 ( new_n2053 , new_n2051 , new_n2052 );
  nand g01677 ( new_n2054 , pi156 , pi158 );
  or   g01678 ( new_n2055 , new_n2030 , new_n2054 );
  nand g01679 ( new_n2056 , new_n2053 , new_n2055 );
  xor  g01680 ( new_n2057 , new_n2050 , new_n2056 );
  nand g01681 ( new_n2058 , new_n2029 , new_n2030 );
  nand g01682 ( new_n2059 , new_n2028 , new_n2031 );
  nand g01683 ( new_n2060 , new_n2058 , new_n2059 );
  xor  g01684 ( new_n2061 , new_n2057 , new_n2060 );
  nand g01685 ( new_n2062 , pi049 , pi154 );
  nand g01686 ( new_n2063 , pi095 , pi171 );
  nand g01687 ( new_n2064 , new_n2062 , new_n2063 );
  nand g01688 ( new_n2065 , pi049 , pi095 );
  or   g01689 ( new_n2066 , new_n2033 , new_n2065 );
  nand g01690 ( new_n2067 , new_n2064 , new_n2066 );
  xor  g01691 ( new_n2068 , new_n2061 , new_n2067 );
  xor  g01692 ( new_n2069 , new_n2049 , new_n2068 );
  not  g01693 ( new_n2070 , new_n2039 );
  nand g01694 ( new_n2071 , new_n2070 , new_n2042 );
  or   g01695 ( new_n2072 , new_n2038 , new_n2043 );
  nand g01696 ( new_n2073 , new_n2071 , new_n2072 );
  xor  g01697 ( new_n2074 , new_n2069 , new_n2073 );
  xor  g01698 ( new_n2075 , new_n2004 , new_n2045 );
  nand g01699 ( new_n2076 , new_n2074 , new_n2075 );
  nand g01700 ( new_n2077 , new_n2046 , new_n2076 );
  not  g01701 ( new_n2078 , new_n2069 );
  nand g01702 ( new_n2079 , new_n2078 , new_n2073 );
  nand g01703 ( new_n2080 , pi089 , pi201 );
  nand g01704 ( new_n2081 , pi063 , pi254 );
  xor  g01705 ( new_n2082 , new_n2080 , new_n2081 );
  xor  g01706 ( new_n2083 , new_n2054 , new_n2082 );
  not  g01707 ( new_n2084 , new_n2083 );
  nand g01708 ( new_n2085 , pi154 , pi245 );
  xor  g01709 ( new_n2086 , new_n2055 , new_n2085 );
  xor  g01710 ( new_n2087 , new_n2084 , new_n2086 );
  nand g01711 ( new_n2088 , pi006 , pi171 );
  nand g01712 ( new_n2089 , pi107 , pi209 );
  xor  g01713 ( new_n2090 , new_n2088 , new_n2089 );
  xor  g01714 ( new_n2091 , new_n2065 , new_n2090 );
  nand g01715 ( new_n2092 , new_n2050 , new_n2056 );
  nand g01716 ( new_n2093 , new_n2057 , new_n2060 );
  nand g01717 ( new_n2094 , new_n2092 , new_n2093 );
  xor  g01718 ( new_n2095 , new_n2091 , new_n2094 );
  xor  g01719 ( new_n2096 , new_n2087 , new_n2095 );
  nand g01720 ( new_n2097 , new_n2061 , new_n2067 );
  nand g01721 ( new_n2098 , new_n2049 , new_n2068 );
  nand g01722 ( new_n2099 , new_n2097 , new_n2098 );
  xor  g01723 ( new_n2100 , new_n2066 , new_n2099 );
  xnor g01724 ( new_n2101 , new_n2096 , new_n2100 );
  xor  g01725 ( new_n2102 , new_n2079 , new_n2101 );
  xnor g01726 ( new_n2103 , new_n2077 , new_n2102 );
  nand g01727 ( new_n2104 , pi039 , pi073 );
  nand g01728 ( new_n2105 , pi073 , pi228 );
  nand g01729 ( new_n2106 , pi116 , pi170 );
  nand g01730 ( new_n2107 , new_n2105 , new_n2106 );
  nand g01731 ( new_n2108 , pi004 , pi039 );
  xor  g01732 ( new_n2109 , new_n2105 , new_n2106 );
  nand g01733 ( new_n2110 , new_n2108 , new_n2109 );
  nand g01734 ( new_n2111 , new_n2107 , new_n2110 );
  xor  g01735 ( new_n2112 , new_n2104 , new_n2111 );
  nand g01736 ( new_n2113 , pi070 , pi170 );
  nand g01737 ( new_n2114 , pi004 , pi116 );
  nand g01738 ( new_n2115 , new_n2113 , new_n2114 );
  nand g01739 ( new_n2116 , pi004 , pi070 );
  nor  g01740 ( new_n2117 , new_n2106 , new_n2116 );
  not  g01741 ( new_n2118 , new_n2117 );
  nand g01742 ( new_n2119 , new_n2115 , new_n2118 );
  xor  g01743 ( new_n2120 , new_n2112 , new_n2119 );
  nand g01744 ( new_n2121 , pi130 , pi148 );
  nand g01745 ( new_n2122 , pi003 , pi228 );
  and  g01746 ( new_n2123 , new_n2121 , new_n2122 );
  nand g01747 ( new_n2124 , pi130 , pi228 );
  nand g01748 ( new_n2125 , pi003 , pi148 );
  nor  g01749 ( new_n2126 , new_n2124 , new_n2125 );
  or   g01750 ( new_n2127 , new_n2123 , new_n2126 );
  xnor g01751 ( new_n2128 , new_n2120 , new_n2127 );
  nand g01752 ( new_n2129 , pi004 , pi228 );
  nand g01753 ( new_n2130 , pi073 , pi148 );
  nand g01754 ( new_n2131 , new_n2129 , new_n2130 );
  nand g01755 ( new_n2132 , pi039 , pi170 );
  xor  g01756 ( new_n2133 , new_n2129 , new_n2130 );
  nand g01757 ( new_n2134 , new_n2132 , new_n2133 );
  nand g01758 ( new_n2135 , new_n2131 , new_n2134 );
  nand g01759 ( new_n2136 , new_n2125 , new_n2135 );
  xor  g01760 ( new_n2137 , new_n2108 , new_n2109 );
  xor  g01761 ( new_n2138 , new_n2125 , new_n2135 );
  nand g01762 ( new_n2139 , new_n2137 , new_n2138 );
  nand g01763 ( new_n2140 , new_n2136 , new_n2139 );
  xor  g01764 ( new_n2141 , new_n2128 , new_n2140 );
  nand g01765 ( new_n2142 , pi130 , pi163 );
  nand g01766 ( new_n2143 , pi170 , pi228 );
  nand g01767 ( new_n2144 , pi073 , pi163 );
  nand g01768 ( new_n2145 , new_n2143 , new_n2144 );
  nand g01769 ( new_n2146 , pi004 , pi148 );
  or   g01770 ( new_n2147 , new_n2143 , new_n2144 );
  nand g01771 ( new_n2148 , new_n2146 , new_n2147 );
  nand g01772 ( new_n2149 , new_n2145 , new_n2148 );
  nand g01773 ( new_n2150 , pi003 , pi163 );
  nand g01774 ( new_n2151 , new_n2149 , new_n2150 );
  xor  g01775 ( new_n2152 , new_n2132 , new_n2133 );
  xor  g01776 ( new_n2153 , new_n2149 , new_n2150 );
  nand g01777 ( new_n2154 , new_n2152 , new_n2153 );
  nand g01778 ( new_n2155 , new_n2151 , new_n2154 );
  or   g01779 ( new_n2156 , new_n2142 , new_n2155 );
  xnor g01780 ( new_n2157 , new_n2137 , new_n2138 );
  xor  g01781 ( new_n2158 , new_n2142 , new_n2155 );
  nand g01782 ( new_n2159 , new_n2157 , new_n2158 );
  nand g01783 ( new_n2160 , new_n2156 , new_n2159 );
  nand g01784 ( new_n2161 , new_n2141 , new_n2160 );
  nand g01785 ( new_n2162 , pi073 , pi116 );
  nand g01786 ( new_n2163 , pi115 , pi170 );
  xor  g01787 ( new_n2164 , new_n2162 , new_n2163 );
  xor  g01788 ( new_n2165 , new_n2116 , new_n2164 );
  nand g01789 ( new_n2166 , pi003 , pi039 );
  xor  g01790 ( new_n2167 , new_n2118 , new_n2166 );
  not  g01791 ( new_n2168 , new_n2167 );
  xor  g01792 ( new_n2169 , new_n2165 , new_n2168 );
  nand g01793 ( new_n2170 , pi124 , pi148 );
  nand g01794 ( new_n2171 , pi163 , pi215 );
  xor  g01795 ( new_n2172 , new_n2124 , new_n2171 );
  xor  g01796 ( new_n2173 , new_n2170 , new_n2172 );
  nand g01797 ( new_n2174 , new_n2104 , new_n2111 );
  nand g01798 ( new_n2175 , new_n2112 , new_n2119 );
  nand g01799 ( new_n2176 , new_n2174 , new_n2175 );
  xor  g01800 ( new_n2177 , new_n2173 , new_n2176 );
  xor  g01801 ( new_n2178 , new_n2169 , new_n2177 );
  nor  g01802 ( new_n2179 , new_n2128 , new_n2140 );
  nand g01803 ( new_n2180 , new_n2126 , new_n2179 );
  nor  g01804 ( new_n2181 , new_n2120 , new_n2127 );
  or   g01805 ( new_n2182 , new_n2126 , new_n2181 );
  or   g01806 ( new_n2183 , new_n2179 , new_n2182 );
  nand g01807 ( new_n2184 , new_n2180 , new_n2183 );
  xor  g01808 ( new_n2185 , new_n2178 , new_n2184 );
  xor  g01809 ( new_n2186 , new_n2161 , new_n2185 );
  xnor g01810 ( new_n2187 , new_n2141 , new_n2160 );
  nand g01811 ( new_n2188 , pi124 , pi163 );
  or   g01812 ( new_n2189 , new_n2187 , new_n2188 );
  xor  g01813 ( new_n2190 , new_n2152 , new_n2153 );
  not  g01814 ( new_n2191 , new_n2146 );
  not  g01815 ( new_n2192 , new_n2145 );
  nand g01816 ( new_n2193 , pi163 , pi170 );
  nand g01817 ( new_n2194 , new_n2191 , new_n2193 );
  nand g01818 ( new_n2195 , new_n2192 , new_n2194 );
  nand g01819 ( new_n2196 , new_n2147 , new_n2195 );
  nand g01820 ( new_n2197 , new_n2191 , new_n2196 );
  nor  g01821 ( new_n2198 , new_n2190 , new_n2197 );
  not  g01822 ( new_n2199 , new_n2198 );
  xnor g01823 ( new_n2200 , new_n2157 , new_n2158 );
  nor  g01824 ( new_n2201 , new_n2199 , new_n2200 );
  xor  g01825 ( new_n2202 , new_n2187 , new_n2188 );
  nand g01826 ( new_n2203 , new_n2201 , new_n2202 );
  nand g01827 ( new_n2204 , new_n2189 , new_n2203 );
  xor  g01828 ( new_n2205 , new_n2186 , new_n2204 );
  xor  g01829 ( new_n2206 , new_n2103 , new_n2205 );
  xor  g01830 ( new_n2207 , new_n2074 , new_n2075 );
  not  g01831 ( new_n2208 , new_n2207 );
  xor  g01832 ( new_n2209 , new_n2201 , new_n2202 );
  nand g01833 ( new_n2210 , new_n2208 , new_n2209 );
  not  g01834 ( new_n2211 , new_n2210 );
  xnor g01835 ( new_n2212 , new_n2027 , new_n2044 );
  xnor g01836 ( new_n2213 , new_n2019 , new_n2026 );
  and  g01837 ( new_n2214 , new_n2012 , new_n2023 );
  or   g01838 ( new_n2215 , new_n2025 , new_n2214 );
  nor  g01839 ( new_n2216 , new_n2192 , new_n2194 );
  nor  g01840 ( new_n2217 , new_n2196 , new_n2216 );
  not  g01841 ( new_n2218 , new_n2217 );
  nand g01842 ( new_n2219 , new_n2215 , new_n2218 );
  xor  g01843 ( new_n2220 , new_n2215 , new_n2217 );
  nor  g01844 ( new_n2221 , new_n2021 , new_n2193 );
  nand g01845 ( new_n2222 , pi171 , pi254 );
  nand g01846 ( new_n2223 , pi107 , pi158 );
  xor  g01847 ( new_n2224 , new_n2222 , new_n2223 );
  nand g01848 ( new_n2225 , new_n2221 , new_n2224 );
  nand g01849 ( new_n2226 , pi004 , pi163 );
  nand g01850 ( new_n2227 , pi148 , pi170 );
  xor  g01851 ( new_n2228 , new_n2226 , new_n2227 );
  xor  g01852 ( new_n2229 , new_n2221 , new_n2224 );
  nand g01853 ( new_n2230 , new_n2228 , new_n2229 );
  nand g01854 ( new_n2231 , new_n2225 , new_n2230 );
  or   g01855 ( new_n2232 , new_n2220 , new_n2231 );
  nand g01856 ( new_n2233 , new_n2219 , new_n2232 );
  nand g01857 ( new_n2234 , new_n2213 , new_n2233 );
  xor  g01858 ( new_n2235 , new_n2190 , new_n2197 );
  not  g01859 ( new_n2236 , new_n2235 );
  xor  g01860 ( new_n2237 , new_n2213 , new_n2233 );
  nand g01861 ( new_n2238 , new_n2236 , new_n2237 );
  nand g01862 ( new_n2239 , new_n2234 , new_n2238 );
  nand g01863 ( new_n2240 , new_n2212 , new_n2239 );
  xor  g01864 ( new_n2241 , new_n2198 , new_n2200 );
  xor  g01865 ( new_n2242 , new_n2212 , new_n2239 );
  nand g01866 ( new_n2243 , new_n2241 , new_n2242 );
  nand g01867 ( new_n2244 , new_n2240 , new_n2243 );
  xor  g01868 ( new_n2245 , new_n2207 , new_n2209 );
  nor  g01869 ( new_n2246 , new_n2244 , new_n2245 );
  nor  g01870 ( new_n2247 , new_n2211 , new_n2246 );
  xor  g01871 ( new_n2248 , new_n2206 , new_n2247 );
  nand g01872 ( new_n2249 , pi134 , pi172 );
  nand g01873 ( new_n2250 , pi062 , pi240 );
  nand g01874 ( new_n2251 , pi065 , pi149 );
  nand g01875 ( new_n2252 , new_n2250 , new_n2251 );
  nand g01876 ( new_n2253 , pi120 , pi134 );
  xor  g01877 ( new_n2254 , new_n2250 , new_n2251 );
  nand g01878 ( new_n2255 , new_n2253 , new_n2254 );
  nand g01879 ( new_n2256 , new_n2252 , new_n2255 );
  nand g01880 ( new_n2257 , new_n2249 , new_n2256 );
  nand g01881 ( new_n2258 , pi065 , pi167 );
  nand g01882 ( new_n2259 , pi120 , pi240 );
  nand g01883 ( new_n2260 , pi062 , pi149 );
  xor  g01884 ( new_n2261 , new_n2259 , new_n2260 );
  xor  g01885 ( new_n2262 , new_n2258 , new_n2261 );
  xor  g01886 ( new_n2263 , new_n2249 , new_n2256 );
  nand g01887 ( new_n2264 , new_n2262 , new_n2263 );
  nand g01888 ( new_n2265 , new_n2257 , new_n2264 );
  nand g01889 ( new_n2266 , pi120 , pi149 );
  nand g01890 ( new_n2267 , pi062 , pi167 );
  nand g01891 ( new_n2268 , pi065 , pi181 );
  nand g01892 ( new_n2269 , new_n2267 , new_n2268 );
  nand g01893 ( new_n2270 , pi062 , pi181 );
  or   g01894 ( new_n2271 , new_n2258 , new_n2270 );
  nand g01895 ( new_n2272 , new_n2269 , new_n2271 );
  xor  g01896 ( new_n2273 , new_n2266 , new_n2272 );
  nand g01897 ( new_n2274 , new_n2259 , new_n2260 );
  nand g01898 ( new_n2275 , new_n2258 , new_n2261 );
  nand g01899 ( new_n2276 , new_n2274 , new_n2275 );
  xor  g01900 ( new_n2277 , new_n2273 , new_n2276 );
  nand g01901 ( new_n2278 , pi172 , pi240 );
  nand g01902 ( new_n2279 , pi134 , pi198 );
  nand g01903 ( new_n2280 , new_n2278 , new_n2279 );
  nand g01904 ( new_n2281 , pi198 , pi240 );
  or   g01905 ( new_n2282 , new_n2249 , new_n2281 );
  nand g01906 ( new_n2283 , new_n2280 , new_n2282 );
  xor  g01907 ( new_n2284 , new_n2277 , new_n2283 );
  xor  g01908 ( new_n2285 , new_n2265 , new_n2284 );
  xor  g01909 ( new_n2286 , new_n2262 , new_n2263 );
  nand g01910 ( new_n2287 , pi175 , pi198 );
  or   g01911 ( new_n2288 , new_n2286 , new_n2287 );
  xor  g01912 ( new_n2289 , new_n2286 , new_n2287 );
  nand g01913 ( new_n2290 , pi120 , pi175 );
  nand g01914 ( new_n2291 , pi065 , pi240 );
  nand g01915 ( new_n2292 , new_n2290 , new_n2291 );
  nand g01916 ( new_n2293 , pi062 , pi134 );
  or   g01917 ( new_n2294 , new_n2290 , new_n2291 );
  nand g01918 ( new_n2295 , new_n2293 , new_n2294 );
  nand g01919 ( new_n2296 , new_n2292 , new_n2295 );
  nand g01920 ( new_n2297 , pi172 , pi175 );
  or   g01921 ( new_n2298 , new_n2296 , new_n2297 );
  xor  g01922 ( new_n2299 , new_n2296 , new_n2297 );
  xnor g01923 ( new_n2300 , new_n2253 , new_n2254 );
  nand g01924 ( new_n2301 , new_n2299 , new_n2300 );
  nand g01925 ( new_n2302 , new_n2298 , new_n2301 );
  nand g01926 ( new_n2303 , new_n2289 , new_n2302 );
  nand g01927 ( new_n2304 , new_n2288 , new_n2303 );
  xor  g01928 ( new_n2305 , new_n2285 , new_n2304 );
  xnor g01929 ( new_n2306 , new_n2299 , new_n2300 );
  not  g01930 ( new_n2307 , new_n2293 );
  not  g01931 ( new_n2308 , new_n2292 );
  nand g01932 ( new_n2309 , pi065 , pi175 );
  nand g01933 ( new_n2310 , new_n2307 , new_n2309 );
  nand g01934 ( new_n2311 , new_n2308 , new_n2310 );
  nand g01935 ( new_n2312 , new_n2294 , new_n2311 );
  nand g01936 ( new_n2313 , new_n2307 , new_n2312 );
  nor  g01937 ( new_n2314 , new_n2306 , new_n2313 );
  xor  g01938 ( new_n2315 , new_n2289 , new_n2302 );
  nand g01939 ( new_n2316 , new_n2314 , new_n2315 );
  nand g01940 ( new_n2317 , pi165 , pi175 );
  xor  g01941 ( new_n2318 , new_n2316 , new_n2317 );
  xor  g01942 ( new_n2319 , new_n2305 , new_n2318 );
  xor  g01943 ( new_n2320 , new_n2241 , new_n2242 );
  xor  g01944 ( new_n2321 , new_n2314 , new_n2315 );
  not  g01945 ( new_n2322 , new_n2321 );
  nor  g01946 ( new_n2323 , new_n2320 , new_n2322 );
  xor  g01947 ( new_n2324 , new_n2320 , new_n2321 );
  xor  g01948 ( new_n2325 , new_n2236 , new_n2237 );
  xor  g01949 ( new_n2326 , new_n2306 , new_n2313 );
  not  g01950 ( new_n2327 , new_n2326 );
  nand g01951 ( new_n2328 , new_n2325 , new_n2327 );
  xor  g01952 ( new_n2329 , new_n2325 , new_n2327 );
  xor  g01953 ( new_n2330 , new_n2220 , new_n2231 );
  nor  g01954 ( new_n2331 , new_n2308 , new_n2310 );
  nor  g01955 ( new_n2332 , new_n2312 , new_n2331 );
  not  g01956 ( new_n2333 , new_n2332 );
  nor  g01957 ( new_n2334 , new_n2330 , new_n2333 );
  xor  g01958 ( new_n2335 , new_n2330 , new_n2332 );
  xor  g01959 ( new_n2336 , new_n2021 , new_n2193 );
  not  g01960 ( new_n2337 , new_n2336 );
  nor  g01961 ( new_n2338 , new_n2309 , new_n2337 );
  nand g01962 ( new_n2339 , pi062 , pi175 );
  nand g01963 ( new_n2340 , pi065 , pi134 );
  xor  g01964 ( new_n2341 , new_n2339 , new_n2340 );
  or   g01965 ( new_n2342 , new_n2338 , new_n2341 );
  xor  g01966 ( new_n2343 , new_n2228 , new_n2229 );
  not  g01967 ( new_n2344 , new_n2343 );
  xor  g01968 ( new_n2345 , new_n2338 , new_n2341 );
  nand g01969 ( new_n2346 , new_n2344 , new_n2345 );
  nand g01970 ( new_n2347 , new_n2342 , new_n2346 );
  nor  g01971 ( new_n2348 , new_n2335 , new_n2347 );
  nor  g01972 ( new_n2349 , new_n2334 , new_n2348 );
  nand g01973 ( new_n2350 , new_n2329 , new_n2349 );
  nand g01974 ( new_n2351 , new_n2328 , new_n2350 );
  nor  g01975 ( new_n2352 , new_n2324 , new_n2351 );
  nor  g01976 ( new_n2353 , new_n2323 , new_n2352 );
  nand g01977 ( new_n2354 , new_n2319 , new_n2353 );
  xnor g01978 ( new_n2355 , new_n2244 , new_n2245 );
  xor  g01979 ( new_n2356 , new_n2319 , new_n2353 );
  nand g01980 ( new_n2357 , new_n2355 , new_n2356 );
  nand g01981 ( new_n2358 , new_n2354 , new_n2357 );
  nand g01982 ( new_n2359 , new_n2248 , new_n2358 );
  nand g01983 ( new_n2360 , new_n2316 , new_n2317 );
  nand g01984 ( new_n2361 , new_n2305 , new_n2318 );
  nand g01985 ( new_n2362 , new_n2360 , new_n2361 );
  not  g01986 ( new_n2363 , new_n2285 );
  nand g01987 ( new_n2364 , new_n2363 , new_n2304 );
  nand g01988 ( new_n2365 , pi065 , pi200 );
  nand g01989 ( new_n2366 , pi120 , pi167 );
  xor  g01990 ( new_n2367 , new_n2365 , new_n2366 );
  xor  g01991 ( new_n2368 , new_n2270 , new_n2367 );
  not  g01992 ( new_n2369 , new_n2368 );
  nand g01993 ( new_n2370 , pi149 , pi172 );
  xor  g01994 ( new_n2371 , new_n2271 , new_n2370 );
  xor  g01995 ( new_n2372 , new_n2369 , new_n2371 );
  nand g01996 ( new_n2373 , pi134 , pi165 );
  nand g01997 ( new_n2374 , pi175 , pi197 );
  xor  g01998 ( new_n2375 , new_n2373 , new_n2374 );
  xor  g01999 ( new_n2376 , new_n2281 , new_n2375 );
  nand g02000 ( new_n2377 , new_n2266 , new_n2272 );
  nand g02001 ( new_n2378 , new_n2273 , new_n2276 );
  nand g02002 ( new_n2379 , new_n2377 , new_n2378 );
  xor  g02003 ( new_n2380 , new_n2376 , new_n2379 );
  xor  g02004 ( new_n2381 , new_n2372 , new_n2380 );
  nand g02005 ( new_n2382 , new_n2277 , new_n2283 );
  nand g02006 ( new_n2383 , new_n2265 , new_n2284 );
  nand g02007 ( new_n2384 , new_n2382 , new_n2383 );
  xor  g02008 ( new_n2385 , new_n2282 , new_n2384 );
  xnor g02009 ( new_n2386 , new_n2381 , new_n2385 );
  xor  g02010 ( new_n2387 , new_n2364 , new_n2386 );
  xor  g02011 ( new_n2388 , new_n2362 , new_n2387 );
  xor  g02012 ( new_n2389 , new_n2248 , new_n2358 );
  nand g02013 ( new_n2390 , new_n2388 , new_n2389 );
  nand g02014 ( new_n2391 , new_n2359 , new_n2390 );
  nand g02015 ( new_n2392 , pi229 , pi234 );
  nand g02016 ( new_n2393 , new_n1939 , new_n1940 );
  nand g02017 ( new_n2394 , new_n1916 , new_n1941 );
  nand g02018 ( new_n2395 , new_n2393 , new_n2394 );
  xor  g02019 ( new_n2396 , new_n2392 , new_n2395 );
  xor  g02020 ( new_n2397 , new_n2391 , new_n2396 );
  nand g02021 ( new_n2398 , new_n1946 , new_n1947 );
  nand g02022 ( new_n2399 , new_n1902 , new_n1948 );
  nand g02023 ( new_n2400 , new_n2398 , new_n2399 );
  nand g02024 ( new_n2401 , pi067 , pi247 );
  nand g02025 ( new_n2402 , pi053 , pi080 );
  xor  g02026 ( new_n2403 , new_n2401 , new_n2402 );
  xor  g02027 ( new_n2404 , new_n2400 , new_n2403 );
  nand g02028 ( new_n2405 , new_n2364 , new_n2386 );
  nand g02029 ( new_n2406 , new_n2362 , new_n2387 );
  nand g02030 ( new_n2407 , new_n2405 , new_n2406 );
  nand g02031 ( new_n2408 , pi092 , pi214 );
  xor  g02032 ( new_n2409 , new_n2407 , new_n2408 );
  xor  g02033 ( new_n2410 , new_n2404 , new_n2409 );
  nand g02034 ( new_n2411 , pi062 , pi200 );
  nand g02035 ( new_n2412 , pi065 , pi203 );
  or   g02036 ( new_n2413 , new_n2282 , new_n2384 );
  nand g02037 ( new_n2414 , new_n2381 , new_n2385 );
  nand g02038 ( new_n2415 , new_n2413 , new_n2414 );
  xnor g02039 ( new_n2416 , new_n2412 , new_n2415 );
  xor  g02040 ( new_n2417 , new_n2411 , new_n2416 );
  nand g02041 ( new_n2418 , pi078 , pi175 );
  nand g02042 ( new_n2419 , new_n1949 , new_n1952 );
  nand g02043 ( new_n2420 , new_n1945 , new_n1953 );
  nand g02044 ( new_n2421 , new_n2419 , new_n2420 );
  xor  g02045 ( new_n2422 , new_n2418 , new_n2421 );
  xor  g02046 ( new_n2423 , new_n2417 , new_n2422 );
  nand g02047 ( new_n2424 , pi030 , pi117 );
  nand g02048 ( new_n2425 , pi016 , pi185 );
  or   g02049 ( new_n2426 , new_n1917 , new_n1943 );
  not  g02050 ( new_n2427 , new_n1942 );
  nand g02051 ( new_n2428 , new_n2427 , new_n1944 );
  nand g02052 ( new_n2429 , new_n2426 , new_n2428 );
  xor  g02053 ( new_n2430 , new_n2425 , new_n2429 );
  xor  g02054 ( new_n2431 , new_n2424 , new_n2430 );
  xor  g02055 ( new_n2432 , new_n2423 , new_n2431 );
  xor  g02056 ( new_n2433 , new_n2410 , new_n2432 );
  xor  g02057 ( new_n2434 , new_n2397 , new_n2433 );
  nand g02058 ( new_n2435 , pi134 , pi197 );
  nand g02059 ( new_n2436 , new_n2365 , new_n2366 );
  nand g02060 ( new_n2437 , new_n2270 , new_n2367 );
  nand g02061 ( new_n2438 , new_n2436 , new_n2437 );
  xor  g02062 ( new_n2439 , new_n2435 , new_n2438 );
  nand g02063 ( new_n2440 , pi000 , pi170 );
  nand g02064 ( new_n2441 , pi004 , pi115 );
  nand g02065 ( new_n2442 , pi070 , pi073 );
  xor  g02066 ( new_n2443 , new_n2441 , new_n2442 );
  nand g02067 ( new_n2444 , pi022 , pi163 );
  nand g02068 ( new_n2445 , new_n2376 , new_n2379 );
  not  g02069 ( new_n2446 , new_n2372 );
  nand g02070 ( new_n2447 , new_n2446 , new_n2380 );
  nand g02071 ( new_n2448 , new_n2445 , new_n2447 );
  xor  g02072 ( new_n2449 , new_n2444 , new_n2448 );
  xor  g02073 ( new_n2450 , new_n2443 , new_n2449 );
  xor  g02074 ( new_n2451 , new_n2440 , new_n2450 );
  xor  g02075 ( new_n2452 , new_n2439 , new_n2451 );
  xor  g02076 ( new_n2453 , new_n2434 , new_n2452 );
  xor  g02077 ( new_n2454 , new_n2003 , new_n2453 );
  nand g02078 ( new_n2455 , pi190 , pi202 );
  nand g02079 ( new_n2456 , pi103 , pi220 );
  xor  g02080 ( new_n2457 , new_n2455 , new_n2456 );
  nand g02081 ( new_n2458 , pi171 , pi209 );
  nand g02082 ( new_n2459 , new_n2091 , new_n2094 );
  not  g02083 ( new_n2460 , new_n2087 );
  nand g02084 ( new_n2461 , new_n2460 , new_n2095 );
  nand g02085 ( new_n2462 , new_n2459 , new_n2461 );
  xor  g02086 ( new_n2463 , new_n2458 , new_n2462 );
  xor  g02087 ( new_n2464 , new_n2457 , new_n2463 );
  nand g02088 ( new_n2465 , new_n2173 , new_n2176 );
  not  g02089 ( new_n2466 , new_n2169 );
  nand g02090 ( new_n2467 , new_n2466 , new_n2177 );
  nand g02091 ( new_n2468 , new_n2465 , new_n2467 );
  nand g02092 ( new_n2469 , new_n2079 , new_n2101 );
  nand g02093 ( new_n2470 , new_n2077 , new_n2102 );
  nand g02094 ( new_n2471 , new_n2469 , new_n2470 );
  xor  g02095 ( new_n2472 , new_n2468 , new_n2471 );
  nand g02096 ( new_n2473 , new_n2124 , new_n2171 );
  nand g02097 ( new_n2474 , new_n2170 , new_n2172 );
  nand g02098 ( new_n2475 , new_n2473 , new_n2474 );
  xor  g02099 ( new_n2476 , new_n2472 , new_n2475 );
  nor  g02100 ( new_n2477 , new_n2118 , new_n2166 );
  nor  g02101 ( new_n2478 , new_n2165 , new_n2168 );
  or   g02102 ( new_n2479 , new_n2477 , new_n2478 );
  nand g02103 ( new_n2480 , new_n2162 , new_n2163 );
  nand g02104 ( new_n2481 , new_n2116 , new_n2164 );
  nand g02105 ( new_n2482 , new_n2480 , new_n2481 );
  nand g02106 ( new_n2483 , pi003 , pi116 );
  xor  g02107 ( new_n2484 , new_n2482 , new_n2483 );
  or   g02108 ( new_n2485 , new_n2066 , new_n2099 );
  nand g02109 ( new_n2486 , new_n2096 , new_n2100 );
  nand g02110 ( new_n2487 , new_n2485 , new_n2486 );
  nand g02111 ( new_n2488 , pi154 , pi201 );
  nand g02112 ( new_n2489 , pi095 , pi245 );
  xor  g02113 ( new_n2490 , new_n2488 , new_n2489 );
  xor  g02114 ( new_n2491 , new_n2487 , new_n2490 );
  nand g02115 ( new_n2492 , pi063 , pi158 );
  nand g02116 ( new_n2493 , pi107 , pi153 );
  nand g02117 ( new_n2494 , pi089 , pi156 );
  nand g02118 ( new_n2495 , pi083 , pi254 );
  xor  g02119 ( new_n2496 , new_n2494 , new_n2495 );
  xor  g02120 ( new_n2497 , new_n2493 , new_n2496 );
  xor  g02121 ( new_n2498 , new_n2492 , new_n2497 );
  xor  g02122 ( new_n2499 , new_n2491 , new_n2498 );
  nand g02123 ( new_n2500 , pi039 , pi130 );
  nand g02124 ( new_n2501 , pi124 , pi228 );
  nand g02125 ( new_n2502 , pi148 , pi215 );
  xor  g02126 ( new_n2503 , new_n2501 , new_n2502 );
  xor  g02127 ( new_n2504 , new_n2500 , new_n2503 );
  xor  g02128 ( new_n2505 , new_n2499 , new_n2504 );
  xor  g02129 ( new_n2506 , new_n2484 , new_n2505 );
  xor  g02130 ( new_n2507 , new_n2479 , new_n2506 );
  xor  g02131 ( new_n2508 , new_n2476 , new_n2507 );
  nand g02132 ( new_n2509 , new_n2080 , new_n2081 );
  nand g02133 ( new_n2510 , new_n2054 , new_n2082 );
  nand g02134 ( new_n2511 , new_n2509 , new_n2510 );
  or   g02135 ( new_n2512 , new_n2055 , new_n2085 );
  nand g02136 ( new_n2513 , new_n2084 , new_n2086 );
  nand g02137 ( new_n2514 , new_n2512 , new_n2513 );
  nand g02138 ( new_n2515 , new_n2088 , new_n2089 );
  nand g02139 ( new_n2516 , new_n2065 , new_n2090 );
  nand g02140 ( new_n2517 , new_n2515 , new_n2516 );
  nand g02141 ( new_n2518 , pi006 , pi049 );
  xor  g02142 ( new_n2519 , new_n2517 , new_n2518 );
  xor  g02143 ( new_n2520 , new_n2514 , new_n2519 );
  xor  g02144 ( new_n2521 , new_n2511 , new_n2520 );
  xor  g02145 ( new_n2522 , new_n2508 , new_n2521 );
  xor  g02146 ( new_n2523 , new_n2464 , new_n2522 );
  nand g02147 ( new_n2524 , pi120 , pi181 );
  nand g02148 ( new_n2525 , new_n2373 , new_n2374 );
  nand g02149 ( new_n2526 , new_n2281 , new_n2375 );
  nand g02150 ( new_n2527 , new_n2525 , new_n2526 );
  or   g02151 ( new_n2528 , new_n2178 , new_n2184 );
  nand g02152 ( new_n2529 , new_n2183 , new_n2528 );
  xor  g02153 ( new_n2530 , new_n2527 , new_n2529 );
  or   g02154 ( new_n2531 , new_n2161 , new_n2185 );
  nand g02155 ( new_n2532 , new_n2186 , new_n2204 );
  nand g02156 ( new_n2533 , new_n2531 , new_n2532 );
  xor  g02157 ( new_n2534 , new_n2530 , new_n2533 );
  xor  g02158 ( new_n2535 , new_n2524 , new_n2534 );
  xor  g02159 ( new_n2536 , new_n1999 , new_n2000 );
  xor  g02160 ( new_n2537 , new_n2388 , new_n2389 );
  or   g02161 ( new_n2538 , new_n2536 , new_n2537 );
  xor  g02162 ( new_n2539 , new_n2536 , new_n2537 );
  xor  g02163 ( new_n2540 , new_n2355 , new_n2356 );
  xor  g02164 ( new_n2541 , new_n1996 , new_n1997 );
  or   g02165 ( new_n2542 , new_n2540 , new_n2541 );
  xor  g02166 ( new_n2543 , new_n2540 , new_n2541 );
  xor  g02167 ( new_n2544 , new_n2324 , new_n2351 );
  xor  g02168 ( new_n2545 , new_n1991 , new_n1992 );
  nand g02169 ( new_n2546 , new_n2544 , new_n2545 );
  xor  g02170 ( new_n2547 , new_n2544 , new_n2545 );
  xnor g02171 ( new_n2548 , new_n2329 , new_n2349 );
  xor  g02172 ( new_n2549 , new_n1989 , new_n1990 );
  nor  g02173 ( new_n2550 , new_n2548 , new_n2549 );
  xor  g02174 ( new_n2551 , new_n2548 , new_n2549 );
  not  g02175 ( new_n2552 , new_n2551 );
  xor  g02176 ( new_n2553 , new_n1985 , new_n1988 );
  xor  g02177 ( new_n2554 , new_n2309 , new_n2336 );
  or   g02178 ( new_n2555 , new_n1986 , new_n2554 );
  nand g02179 ( new_n2556 , pi092 , pi103 );
  nand g02180 ( new_n2557 , pi117 , pi190 );
  nand g02181 ( new_n2558 , new_n2556 , new_n2557 );
  nand g02182 ( new_n2559 , new_n1988 , new_n2558 );
  or   g02183 ( new_n2560 , new_n2555 , new_n2559 );
  xor  g02184 ( new_n2561 , new_n2343 , new_n2345 );
  xor  g02185 ( new_n2562 , new_n2555 , new_n2559 );
  nand g02186 ( new_n2563 , new_n2561 , new_n2562 );
  nand g02187 ( new_n2564 , new_n2560 , new_n2563 );
  nand g02188 ( new_n2565 , new_n2553 , new_n2564 );
  xor  g02189 ( new_n2566 , new_n2335 , new_n2347 );
  xor  g02190 ( new_n2567 , new_n2553 , new_n2564 );
  nand g02191 ( new_n2568 , new_n2566 , new_n2567 );
  nand g02192 ( new_n2569 , new_n2565 , new_n2568 );
  nor  g02193 ( new_n2570 , new_n2552 , new_n2569 );
  nor  g02194 ( new_n2571 , new_n2550 , new_n2570 );
  nand g02195 ( new_n2572 , new_n2547 , new_n2571 );
  nand g02196 ( new_n2573 , new_n2546 , new_n2572 );
  nand g02197 ( new_n2574 , new_n2543 , new_n2573 );
  nand g02198 ( new_n2575 , new_n2542 , new_n2574 );
  nand g02199 ( new_n2576 , new_n2539 , new_n2575 );
  nand g02200 ( new_n2577 , new_n2538 , new_n2576 );
  or   g02201 ( new_n2578 , new_n2271 , new_n2370 );
  nand g02202 ( new_n2579 , new_n2369 , new_n2371 );
  nand g02203 ( new_n2580 , new_n2578 , new_n2579 );
  nand g02204 ( new_n2581 , pi149 , pi198 );
  nand g02205 ( new_n2582 , pi165 , pi240 );
  xor  g02206 ( new_n2583 , new_n2581 , new_n2582 );
  xor  g02207 ( new_n2584 , new_n2580 , new_n2583 );
  xor  g02208 ( new_n2585 , new_n2577 , new_n2584 );
  xor  g02209 ( new_n2586 , new_n2535 , new_n2585 );
  nand g02210 ( new_n2587 , new_n2103 , new_n2205 );
  not  g02211 ( new_n2588 , new_n2247 );
  nand g02212 ( new_n2589 , new_n2206 , new_n2588 );
  nand g02213 ( new_n2590 , new_n2587 , new_n2589 );
  nand g02214 ( new_n2591 , pi167 , pi172 );
  xor  g02215 ( new_n2592 , new_n2590 , new_n2591 );
  xor  g02216 ( new_n2593 , new_n2586 , new_n2592 );
  xor  g02217 ( new_n2594 , new_n2523 , new_n2593 );
  xor  g02218 ( po006 , new_n2454 , new_n2594 );
  nand g02219 ( new_n2596 , pi120 , pi216 );
  nand g02220 ( new_n2597 , pi062 , pi076 );
  nand g02221 ( new_n2598 , pi065 , pi079 );
  nand g02222 ( new_n2599 , new_n2597 , new_n2598 );
  nand g02223 ( new_n2600 , pi065 , pi076 );
  nand g02224 ( new_n2601 , pi062 , pi079 );
  or   g02225 ( new_n2602 , new_n2600 , new_n2601 );
  nand g02226 ( new_n2603 , new_n2599 , new_n2602 );
  xor  g02227 ( new_n2604 , new_n2596 , new_n2603 );
  nand g02228 ( new_n2605 , pi041 , pi120 );
  nand g02229 ( new_n2606 , new_n2600 , new_n2605 );
  nand g02230 ( new_n2607 , pi062 , pi216 );
  xor  g02231 ( new_n2608 , new_n2600 , new_n2605 );
  nand g02232 ( new_n2609 , new_n2607 , new_n2608 );
  nand g02233 ( new_n2610 , new_n2606 , new_n2609 );
  xor  g02234 ( new_n2611 , new_n2604 , new_n2610 );
  nand g02235 ( new_n2612 , pi041 , pi172 );
  nand g02236 ( new_n2613 , pi182 , pi198 );
  and  g02237 ( new_n2614 , new_n2612 , new_n2613 );
  nand g02238 ( new_n2615 , pi172 , pi182 );
  nand g02239 ( new_n2616 , pi041 , pi198 );
  nor  g02240 ( new_n2617 , new_n2615 , new_n2616 );
  or   g02241 ( new_n2618 , new_n2614 , new_n2617 );
  xnor g02242 ( new_n2619 , new_n2611 , new_n2618 );
  nand g02243 ( new_n2620 , pi041 , pi062 );
  nand g02244 ( new_n2621 , pi065 , pi216 );
  nand g02245 ( new_n2622 , new_n2620 , new_n2621 );
  nand g02246 ( new_n2623 , pi120 , pi182 );
  xor  g02247 ( new_n2624 , new_n2620 , new_n2621 );
  nand g02248 ( new_n2625 , new_n2623 , new_n2624 );
  nand g02249 ( new_n2626 , new_n2622 , new_n2625 );
  nand g02250 ( new_n2627 , new_n2615 , new_n2626 );
  xor  g02251 ( new_n2628 , new_n2607 , new_n2608 );
  xor  g02252 ( new_n2629 , new_n2615 , new_n2626 );
  nand g02253 ( new_n2630 , new_n2628 , new_n2629 );
  nand g02254 ( new_n2631 , new_n2627 , new_n2630 );
  xor  g02255 ( new_n2632 , new_n2619 , new_n2631 );
  xor  g02256 ( new_n2633 , new_n2628 , new_n2629 );
  nand g02257 ( new_n2634 , pi138 , pi198 );
  or   g02258 ( new_n2635 , new_n2633 , new_n2634 );
  xor  g02259 ( new_n2636 , new_n2633 , new_n2634 );
  nand g02260 ( new_n2637 , pi138 , pi172 );
  nand g02261 ( new_n2638 , pi062 , pi182 );
  nand g02262 ( new_n2639 , pi120 , pi138 );
  nand g02263 ( new_n2640 , new_n2638 , new_n2639 );
  nand g02264 ( new_n2641 , pi041 , pi065 );
  xor  g02265 ( new_n2642 , new_n2638 , new_n2639 );
  nand g02266 ( new_n2643 , new_n2641 , new_n2642 );
  nand g02267 ( new_n2644 , new_n2640 , new_n2643 );
  or   g02268 ( new_n2645 , new_n2637 , new_n2644 );
  xnor g02269 ( new_n2646 , new_n2623 , new_n2624 );
  xor  g02270 ( new_n2647 , new_n2637 , new_n2644 );
  nand g02271 ( new_n2648 , new_n2646 , new_n2647 );
  nand g02272 ( new_n2649 , new_n2645 , new_n2648 );
  nand g02273 ( new_n2650 , new_n2636 , new_n2649 );
  nand g02274 ( new_n2651 , new_n2635 , new_n2650 );
  nand g02275 ( new_n2652 , new_n2632 , new_n2651 );
  nand g02276 ( new_n2653 , pi076 , pi120 );
  nand g02277 ( new_n2654 , pi065 , pi251 );
  xor  g02278 ( new_n2655 , new_n2653 , new_n2654 );
  xor  g02279 ( new_n2656 , new_n2601 , new_n2655 );
  not  g02280 ( new_n2657 , new_n2656 );
  nand g02281 ( new_n2658 , pi172 , pi216 );
  xor  g02282 ( new_n2659 , new_n2602 , new_n2658 );
  xor  g02283 ( new_n2660 , new_n2657 , new_n2659 );
  nand g02284 ( new_n2661 , pi138 , pi197 );
  nand g02285 ( new_n2662 , pi165 , pi182 );
  xor  g02286 ( new_n2663 , new_n2661 , new_n2662 );
  xor  g02287 ( new_n2664 , new_n2616 , new_n2663 );
  nand g02288 ( new_n2665 , new_n2596 , new_n2603 );
  nand g02289 ( new_n2666 , new_n2604 , new_n2610 );
  nand g02290 ( new_n2667 , new_n2665 , new_n2666 );
  xor  g02291 ( new_n2668 , new_n2664 , new_n2667 );
  xor  g02292 ( new_n2669 , new_n2660 , new_n2668 );
  nor  g02293 ( new_n2670 , new_n2619 , new_n2631 );
  nand g02294 ( new_n2671 , new_n2617 , new_n2670 );
  nor  g02295 ( new_n2672 , new_n2611 , new_n2618 );
  or   g02296 ( new_n2673 , new_n2617 , new_n2672 );
  or   g02297 ( new_n2674 , new_n2670 , new_n2673 );
  nand g02298 ( new_n2675 , new_n2671 , new_n2674 );
  xor  g02299 ( new_n2676 , new_n2669 , new_n2675 );
  xnor g02300 ( new_n2677 , new_n2652 , new_n2676 );
  nand g02301 ( new_n2678 , pi138 , pi165 );
  xor  g02302 ( new_n2679 , new_n2641 , new_n2642 );
  nand g02303 ( new_n2680 , pi065 , pi138 );
  nor  g02304 ( new_n2681 , new_n2638 , new_n2680 );
  not  g02305 ( new_n2682 , new_n2681 );
  or   g02306 ( new_n2683 , new_n2679 , new_n2682 );
  xnor g02307 ( new_n2684 , new_n2646 , new_n2647 );
  nor  g02308 ( new_n2685 , new_n2683 , new_n2684 );
  xor  g02309 ( new_n2686 , new_n2636 , new_n2649 );
  nand g02310 ( new_n2687 , new_n2685 , new_n2686 );
  nand g02311 ( new_n2688 , new_n2678 , new_n2687 );
  xnor g02312 ( new_n2689 , new_n2632 , new_n2651 );
  xor  g02313 ( new_n2690 , new_n2678 , new_n2687 );
  nand g02314 ( new_n2691 , new_n2689 , new_n2690 );
  nand g02315 ( new_n2692 , new_n2688 , new_n2691 );
  xor  g02316 ( new_n2693 , new_n2677 , new_n2692 );
  nand g02317 ( new_n2694 , pi001 , pi089 );
  nand g02318 ( new_n2695 , pi001 , pi158 );
  nand g02319 ( new_n2696 , pi122 , pi254 );
  nand g02320 ( new_n2697 , new_n2695 , new_n2696 );
  nand g02321 ( new_n2698 , pi089 , pi102 );
  xor  g02322 ( new_n2699 , new_n2695 , new_n2696 );
  nand g02323 ( new_n2700 , new_n2698 , new_n2699 );
  nand g02324 ( new_n2701 , new_n2697 , new_n2700 );
  xor  g02325 ( new_n2702 , new_n2694 , new_n2701 );
  nand g02326 ( new_n2703 , pi122 , pi158 );
  nand g02327 ( new_n2704 , pi135 , pi254 );
  nand g02328 ( new_n2705 , new_n2703 , new_n2704 );
  nand g02329 ( new_n2706 , pi135 , pi158 );
  nor  g02330 ( new_n2707 , new_n2696 , new_n2706 );
  not  g02331 ( new_n2708 , new_n2707 );
  nand g02332 ( new_n2709 , new_n2705 , new_n2708 );
  xor  g02333 ( new_n2710 , new_n2702 , new_n2709 );
  nand g02334 ( new_n2711 , pi095 , pi219 );
  nand g02335 ( new_n2712 , pi102 , pi154 );
  and  g02336 ( new_n2713 , new_n2711 , new_n2712 );
  nand g02337 ( new_n2714 , pi154 , pi219 );
  nand g02338 ( new_n2715 , pi095 , pi102 );
  nor  g02339 ( new_n2716 , new_n2714 , new_n2715 );
  or   g02340 ( new_n2717 , new_n2713 , new_n2716 );
  xnor g02341 ( new_n2718 , new_n2710 , new_n2717 );
  nand g02342 ( new_n2719 , pi102 , pi158 );
  nand g02343 ( new_n2720 , pi089 , pi219 );
  nand g02344 ( new_n2721 , new_n2719 , new_n2720 );
  nand g02345 ( new_n2722 , pi001 , pi254 );
  xor  g02346 ( new_n2723 , new_n2719 , new_n2720 );
  nand g02347 ( new_n2724 , new_n2722 , new_n2723 );
  nand g02348 ( new_n2725 , new_n2721 , new_n2724 );
  nand g02349 ( new_n2726 , new_n2714 , new_n2725 );
  xor  g02350 ( new_n2727 , new_n2698 , new_n2699 );
  xor  g02351 ( new_n2728 , new_n2714 , new_n2725 );
  nand g02352 ( new_n2729 , new_n2727 , new_n2728 );
  nand g02353 ( new_n2730 , new_n2726 , new_n2729 );
  xor  g02354 ( new_n2731 , new_n2718 , new_n2730 );
  xor  g02355 ( new_n2732 , new_n2727 , new_n2728 );
  nand g02356 ( new_n2733 , pi087 , pi095 );
  or   g02357 ( new_n2734 , new_n2732 , new_n2733 );
  xor  g02358 ( new_n2735 , new_n2732 , new_n2733 );
  nand g02359 ( new_n2736 , pi102 , pi254 );
  nand g02360 ( new_n2737 , pi087 , pi089 );
  nand g02361 ( new_n2738 , new_n2736 , new_n2737 );
  nand g02362 ( new_n2739 , pi158 , pi219 );
  or   g02363 ( new_n2740 , new_n2736 , new_n2737 );
  nand g02364 ( new_n2741 , new_n2739 , new_n2740 );
  nand g02365 ( new_n2742 , new_n2738 , new_n2741 );
  nand g02366 ( new_n2743 , pi087 , pi154 );
  or   g02367 ( new_n2744 , new_n2742 , new_n2743 );
  xor  g02368 ( new_n2745 , new_n2742 , new_n2743 );
  xnor g02369 ( new_n2746 , new_n2722 , new_n2723 );
  nand g02370 ( new_n2747 , new_n2745 , new_n2746 );
  nand g02371 ( new_n2748 , new_n2744 , new_n2747 );
  nand g02372 ( new_n2749 , new_n2735 , new_n2748 );
  nand g02373 ( new_n2750 , new_n2734 , new_n2749 );
  nand g02374 ( new_n2751 , new_n2731 , new_n2750 );
  nand g02375 ( new_n2752 , pi089 , pi122 );
  nand g02376 ( new_n2753 , pi059 , pi254 );
  xor  g02377 ( new_n2754 , new_n2752 , new_n2753 );
  xor  g02378 ( new_n2755 , new_n2706 , new_n2754 );
  nand g02379 ( new_n2756 , pi001 , pi154 );
  xor  g02380 ( new_n2757 , new_n2708 , new_n2756 );
  not  g02381 ( new_n2758 , new_n2757 );
  xor  g02382 ( new_n2759 , new_n2755 , new_n2758 );
  nand g02383 ( new_n2760 , pi087 , pi209 );
  nand g02384 ( new_n2761 , pi006 , pi219 );
  xor  g02385 ( new_n2762 , new_n2715 , new_n2761 );
  xor  g02386 ( new_n2763 , new_n2760 , new_n2762 );
  nand g02387 ( new_n2764 , new_n2694 , new_n2701 );
  nand g02388 ( new_n2765 , new_n2702 , new_n2709 );
  nand g02389 ( new_n2766 , new_n2764 , new_n2765 );
  xor  g02390 ( new_n2767 , new_n2763 , new_n2766 );
  xor  g02391 ( new_n2768 , new_n2759 , new_n2767 );
  nor  g02392 ( new_n2769 , new_n2718 , new_n2730 );
  nand g02393 ( new_n2770 , new_n2716 , new_n2769 );
  nor  g02394 ( new_n2771 , new_n2710 , new_n2717 );
  or   g02395 ( new_n2772 , new_n2716 , new_n2771 );
  or   g02396 ( new_n2773 , new_n2769 , new_n2772 );
  nand g02397 ( new_n2774 , new_n2770 , new_n2773 );
  xor  g02398 ( new_n2775 , new_n2768 , new_n2774 );
  xnor g02399 ( new_n2776 , new_n2751 , new_n2775 );
  xnor g02400 ( new_n2777 , new_n2745 , new_n2746 );
  not  g02401 ( new_n2778 , new_n2739 );
  not  g02402 ( new_n2779 , new_n2738 );
  nand g02403 ( new_n2780 , pi087 , pi254 );
  nand g02404 ( new_n2781 , new_n2778 , new_n2780 );
  nand g02405 ( new_n2782 , new_n2779 , new_n2781 );
  nand g02406 ( new_n2783 , new_n2740 , new_n2782 );
  nand g02407 ( new_n2784 , new_n2778 , new_n2783 );
  nor  g02408 ( new_n2785 , new_n2777 , new_n2784 );
  xor  g02409 ( new_n2786 , new_n2735 , new_n2748 );
  nand g02410 ( new_n2787 , new_n2785 , new_n2786 );
  nand g02411 ( new_n2788 , pi006 , pi087 );
  nand g02412 ( new_n2789 , new_n2787 , new_n2788 );
  xnor g02413 ( new_n2790 , new_n2731 , new_n2750 );
  xor  g02414 ( new_n2791 , new_n2787 , new_n2788 );
  nand g02415 ( new_n2792 , new_n2790 , new_n2791 );
  nand g02416 ( new_n2793 , new_n2789 , new_n2792 );
  xor  g02417 ( new_n2794 , new_n2776 , new_n2793 );
  nand g02418 ( new_n2795 , pi003 , pi071 );
  nand g02419 ( new_n2796 , pi004 , pi169 );
  nand g02420 ( new_n2797 , pi071 , pi073 );
  nand g02421 ( new_n2798 , new_n2796 , new_n2797 );
  nand g02422 ( new_n2799 , pi123 , pi170 );
  xor  g02423 ( new_n2800 , new_n2796 , new_n2797 );
  nand g02424 ( new_n2801 , new_n2799 , new_n2800 );
  nand g02425 ( new_n2802 , new_n2798 , new_n2801 );
  nand g02426 ( new_n2803 , new_n2795 , new_n2802 );
  nand g02427 ( new_n2804 , pi099 , pi170 );
  nand g02428 ( new_n2805 , pi073 , pi169 );
  nand g02429 ( new_n2806 , pi004 , pi123 );
  xor  g02430 ( new_n2807 , new_n2805 , new_n2806 );
  xor  g02431 ( new_n2808 , new_n2804 , new_n2807 );
  xor  g02432 ( new_n2809 , new_n2795 , new_n2802 );
  nand g02433 ( new_n2810 , new_n2808 , new_n2809 );
  nand g02434 ( new_n2811 , new_n2803 , new_n2810 );
  nand g02435 ( new_n2812 , pi073 , pi123 );
  nand g02436 ( new_n2813 , new_n2805 , new_n2806 );
  nand g02437 ( new_n2814 , new_n2804 , new_n2807 );
  nand g02438 ( new_n2815 , new_n2813 , new_n2814 );
  xor  g02439 ( new_n2816 , new_n2812 , new_n2815 );
  nand g02440 ( new_n2817 , pi004 , pi099 );
  nand g02441 ( new_n2818 , pi023 , pi170 );
  nand g02442 ( new_n2819 , new_n2817 , new_n2818 );
  nand g02443 ( new_n2820 , pi004 , pi023 );
  nor  g02444 ( new_n2821 , new_n2804 , new_n2820 );
  not  g02445 ( new_n2822 , new_n2821 );
  nand g02446 ( new_n2823 , new_n2819 , new_n2822 );
  xor  g02447 ( new_n2824 , new_n2816 , new_n2823 );
  nand g02448 ( new_n2825 , pi071 , pi130 );
  nand g02449 ( new_n2826 , pi003 , pi169 );
  nand g02450 ( new_n2827 , new_n2825 , new_n2826 );
  nand g02451 ( new_n2828 , pi130 , pi169 );
  or   g02452 ( new_n2829 , new_n2795 , new_n2828 );
  nand g02453 ( new_n2830 , new_n2827 , new_n2829 );
  xor  g02454 ( new_n2831 , new_n2824 , new_n2830 );
  xnor g02455 ( new_n2832 , new_n2811 , new_n2831 );
  xor  g02456 ( new_n2833 , new_n2808 , new_n2809 );
  nand g02457 ( new_n2834 , pi130 , pi142 );
  or   g02458 ( new_n2835 , new_n2833 , new_n2834 );
  xor  g02459 ( new_n2836 , new_n2833 , new_n2834 );
  nand g02460 ( new_n2837 , pi169 , pi170 );
  nand g02461 ( new_n2838 , pi073 , pi142 );
  nand g02462 ( new_n2839 , new_n2837 , new_n2838 );
  nand g02463 ( new_n2840 , pi004 , pi071 );
  or   g02464 ( new_n2841 , new_n2837 , new_n2838 );
  nand g02465 ( new_n2842 , new_n2840 , new_n2841 );
  nand g02466 ( new_n2843 , new_n2839 , new_n2842 );
  nand g02467 ( new_n2844 , pi003 , pi142 );
  or   g02468 ( new_n2845 , new_n2843 , new_n2844 );
  xor  g02469 ( new_n2846 , new_n2843 , new_n2844 );
  xnor g02470 ( new_n2847 , new_n2799 , new_n2800 );
  nand g02471 ( new_n2848 , new_n2846 , new_n2847 );
  nand g02472 ( new_n2849 , new_n2845 , new_n2848 );
  nand g02473 ( new_n2850 , new_n2836 , new_n2849 );
  nand g02474 ( new_n2851 , new_n2835 , new_n2850 );
  nand g02475 ( new_n2852 , new_n2832 , new_n2851 );
  nand g02476 ( new_n2853 , pi073 , pi099 );
  nand g02477 ( new_n2854 , pi155 , pi170 );
  xor  g02478 ( new_n2855 , new_n2853 , new_n2854 );
  xor  g02479 ( new_n2856 , new_n2820 , new_n2855 );
  nand g02480 ( new_n2857 , pi003 , pi123 );
  xor  g02481 ( new_n2858 , new_n2822 , new_n2857 );
  not  g02482 ( new_n2859 , new_n2858 );
  xor  g02483 ( new_n2860 , new_n2856 , new_n2859 );
  nand g02484 ( new_n2861 , pi142 , pi215 );
  nand g02485 ( new_n2862 , pi071 , pi124 );
  xor  g02486 ( new_n2863 , new_n2861 , new_n2862 );
  xor  g02487 ( new_n2864 , new_n2828 , new_n2863 );
  nand g02488 ( new_n2865 , new_n2812 , new_n2815 );
  nand g02489 ( new_n2866 , new_n2816 , new_n2823 );
  nand g02490 ( new_n2867 , new_n2865 , new_n2866 );
  xor  g02491 ( new_n2868 , new_n2864 , new_n2867 );
  xor  g02492 ( new_n2869 , new_n2860 , new_n2868 );
  not  g02493 ( new_n2870 , new_n2869 );
  nand g02494 ( new_n2871 , new_n2824 , new_n2830 );
  nand g02495 ( new_n2872 , new_n2811 , new_n2831 );
  nand g02496 ( new_n2873 , new_n2871 , new_n2872 );
  xor  g02497 ( new_n2874 , new_n2829 , new_n2873 );
  xor  g02498 ( new_n2875 , new_n2870 , new_n2874 );
  xnor g02499 ( new_n2876 , new_n2852 , new_n2875 );
  nand g02500 ( new_n2877 , pi124 , pi142 );
  xnor g02501 ( new_n2878 , new_n2846 , new_n2847 );
  not  g02502 ( new_n2879 , new_n2840 );
  not  g02503 ( new_n2880 , new_n2839 );
  nand g02504 ( new_n2881 , pi142 , pi170 );
  nand g02505 ( new_n2882 , new_n2879 , new_n2881 );
  nand g02506 ( new_n2883 , new_n2880 , new_n2882 );
  nand g02507 ( new_n2884 , new_n2841 , new_n2883 );
  nand g02508 ( new_n2885 , new_n2879 , new_n2884 );
  nor  g02509 ( new_n2886 , new_n2878 , new_n2885 );
  xor  g02510 ( new_n2887 , new_n2836 , new_n2849 );
  nand g02511 ( new_n2888 , new_n2886 , new_n2887 );
  nand g02512 ( new_n2889 , new_n2877 , new_n2888 );
  xnor g02513 ( new_n2890 , new_n2832 , new_n2851 );
  xor  g02514 ( new_n2891 , new_n2877 , new_n2888 );
  nand g02515 ( new_n2892 , new_n2890 , new_n2891 );
  nand g02516 ( new_n2893 , new_n2889 , new_n2892 );
  xor  g02517 ( new_n2894 , new_n2876 , new_n2893 );
  xor  g02518 ( new_n2895 , new_n2794 , new_n2894 );
  xor  g02519 ( new_n2896 , new_n2790 , new_n2791 );
  xor  g02520 ( new_n2897 , new_n2890 , new_n2891 );
  or   g02521 ( new_n2898 , new_n2896 , new_n2897 );
  xor  g02522 ( new_n2899 , new_n2896 , new_n2897 );
  xor  g02523 ( new_n2900 , new_n2785 , new_n2786 );
  xor  g02524 ( new_n2901 , new_n2886 , new_n2887 );
  nand g02525 ( new_n2902 , new_n2900 , new_n2901 );
  not  g02526 ( new_n2903 , new_n2902 );
  xnor g02527 ( new_n2904 , new_n2900 , new_n2901 );
  xnor g02528 ( new_n2905 , new_n2777 , new_n2784 );
  nor  g02529 ( new_n2906 , new_n2880 , new_n2882 );
  or   g02530 ( new_n2907 , new_n2884 , new_n2906 );
  nor  g02531 ( new_n2908 , new_n2779 , new_n2781 );
  nor  g02532 ( new_n2909 , new_n2783 , new_n2908 );
  not  g02533 ( new_n2910 , new_n2909 );
  nand g02534 ( new_n2911 , new_n2907 , new_n2910 );
  xor  g02535 ( new_n2912 , new_n2907 , new_n2909 );
  nor  g02536 ( new_n2913 , new_n2780 , new_n2881 );
  nand g02537 ( new_n2914 , pi087 , pi158 );
  nand g02538 ( new_n2915 , pi219 , pi254 );
  xor  g02539 ( new_n2916 , new_n2914 , new_n2915 );
  nand g02540 ( new_n2917 , new_n2913 , new_n2916 );
  nand g02541 ( new_n2918 , pi004 , pi142 );
  nand g02542 ( new_n2919 , pi071 , pi170 );
  xor  g02543 ( new_n2920 , new_n2918 , new_n2919 );
  xor  g02544 ( new_n2921 , new_n2913 , new_n2916 );
  nand g02545 ( new_n2922 , new_n2920 , new_n2921 );
  nand g02546 ( new_n2923 , new_n2917 , new_n2922 );
  or   g02547 ( new_n2924 , new_n2912 , new_n2923 );
  nand g02548 ( new_n2925 , new_n2911 , new_n2924 );
  nand g02549 ( new_n2926 , new_n2905 , new_n2925 );
  xor  g02550 ( new_n2927 , new_n2878 , new_n2885 );
  not  g02551 ( new_n2928 , new_n2927 );
  xor  g02552 ( new_n2929 , new_n2905 , new_n2925 );
  nand g02553 ( new_n2930 , new_n2928 , new_n2929 );
  nand g02554 ( new_n2931 , new_n2926 , new_n2930 );
  nor  g02555 ( new_n2932 , new_n2904 , new_n2931 );
  nor  g02556 ( new_n2933 , new_n2903 , new_n2932 );
  not  g02557 ( new_n2934 , new_n2933 );
  nand g02558 ( new_n2935 , new_n2899 , new_n2934 );
  nand g02559 ( new_n2936 , new_n2898 , new_n2935 );
  xor  g02560 ( new_n2937 , new_n2895 , new_n2936 );
  xor  g02561 ( new_n2938 , new_n2693 , new_n2937 );
  xor  g02562 ( new_n2939 , new_n2899 , new_n2933 );
  xor  g02563 ( new_n2940 , new_n2689 , new_n2690 );
  nor  g02564 ( new_n2941 , new_n2939 , new_n2940 );
  xnor g02565 ( new_n2942 , new_n2939 , new_n2940 );
  xor  g02566 ( new_n2943 , new_n2685 , new_n2686 );
  xor  g02567 ( new_n2944 , new_n2928 , new_n2929 );
  not  g02568 ( new_n2945 , new_n2944 );
  xor  g02569 ( new_n2946 , new_n2683 , new_n2684 );
  nor  g02570 ( new_n2947 , new_n2945 , new_n2946 );
  xor  g02571 ( new_n2948 , new_n2944 , new_n2946 );
  xor  g02572 ( new_n2949 , new_n2679 , new_n2681 );
  xor  g02573 ( new_n2950 , new_n2780 , new_n2881 );
  not  g02574 ( new_n2951 , new_n2950 );
  or   g02575 ( new_n2952 , new_n2680 , new_n2951 );
  nand g02576 ( new_n2953 , pi062 , pi138 );
  nand g02577 ( new_n2954 , pi065 , pi182 );
  nand g02578 ( new_n2955 , new_n2953 , new_n2954 );
  nand g02579 ( new_n2956 , new_n2682 , new_n2955 );
  nand g02580 ( new_n2957 , new_n2952 , new_n2956 );
  xor  g02581 ( new_n2958 , new_n2920 , new_n2921 );
  not  g02582 ( new_n2959 , new_n2958 );
  xor  g02583 ( new_n2960 , new_n2952 , new_n2956 );
  nand g02584 ( new_n2961 , new_n2959 , new_n2960 );
  nand g02585 ( new_n2962 , new_n2957 , new_n2961 );
  or   g02586 ( new_n2963 , new_n2949 , new_n2962 );
  xnor g02587 ( new_n2964 , new_n2912 , new_n2923 );
  xor  g02588 ( new_n2965 , new_n2949 , new_n2962 );
  nand g02589 ( new_n2966 , new_n2964 , new_n2965 );
  nand g02590 ( new_n2967 , new_n2963 , new_n2966 );
  nor  g02591 ( new_n2968 , new_n2948 , new_n2967 );
  nor  g02592 ( new_n2969 , new_n2947 , new_n2968 );
  or   g02593 ( new_n2970 , new_n2943 , new_n2969 );
  xor  g02594 ( new_n2971 , new_n2904 , new_n2931 );
  not  g02595 ( new_n2972 , new_n2971 );
  xor  g02596 ( new_n2973 , new_n2943 , new_n2969 );
  nand g02597 ( new_n2974 , new_n2972 , new_n2973 );
  nand g02598 ( new_n2975 , new_n2970 , new_n2974 );
  nor  g02599 ( new_n2976 , new_n2942 , new_n2975 );
  nor  g02600 ( new_n2977 , new_n2941 , new_n2976 );
  xnor g02601 ( new_n2978 , new_n2938 , new_n2977 );
  nand g02602 ( new_n2979 , pi101 , pi190 );
  nand g02603 ( new_n2980 , pi060 , pi229 );
  nand g02604 ( new_n2981 , pi092 , pi223 );
  xor  g02605 ( new_n2982 , new_n2980 , new_n2981 );
  xor  g02606 ( new_n2983 , new_n2979 , new_n2982 );
  nand g02607 ( new_n2984 , pi020 , pi067 );
  nand g02608 ( new_n2985 , pi060 , pi092 );
  nand g02609 ( new_n2986 , pi020 , pi229 );
  nand g02610 ( new_n2987 , new_n2985 , new_n2986 );
  nand g02611 ( new_n2988 , pi190 , pi223 );
  xor  g02612 ( new_n2989 , new_n2985 , new_n2986 );
  nand g02613 ( new_n2990 , new_n2988 , new_n2989 );
  nand g02614 ( new_n2991 , new_n2987 , new_n2990 );
  xor  g02615 ( new_n2992 , new_n2984 , new_n2991 );
  xor  g02616 ( new_n2993 , new_n2983 , new_n2992 );
  nand g02617 ( new_n2994 , pi053 , pi160 );
  or   g02618 ( new_n2995 , new_n2993 , new_n2994 );
  xor  g02619 ( new_n2996 , new_n2993 , new_n2994 );
  nand g02620 ( new_n2997 , pi060 , pi190 );
  nand g02621 ( new_n2998 , pi160 , pi229 );
  nand g02622 ( new_n2999 , new_n2997 , new_n2998 );
  nand g02623 ( new_n3000 , pi020 , pi092 );
  or   g02624 ( new_n3001 , new_n2997 , new_n2998 );
  nand g02625 ( new_n3002 , new_n3000 , new_n3001 );
  nand g02626 ( new_n3003 , new_n2999 , new_n3002 );
  nand g02627 ( new_n3004 , pi067 , pi160 );
  or   g02628 ( new_n3005 , new_n3003 , new_n3004 );
  xnor g02629 ( new_n3006 , new_n2988 , new_n2989 );
  xor  g02630 ( new_n3007 , new_n3003 , new_n3004 );
  nand g02631 ( new_n3008 , new_n3006 , new_n3007 );
  nand g02632 ( new_n3009 , new_n3005 , new_n3008 );
  nand g02633 ( new_n3010 , new_n2996 , new_n3009 );
  nand g02634 ( new_n3011 , new_n2995 , new_n3010 );
  nand g02635 ( new_n3012 , pi223 , pi229 );
  nand g02636 ( new_n3013 , new_n2980 , new_n2981 );
  nand g02637 ( new_n3014 , new_n2979 , new_n2982 );
  nand g02638 ( new_n3015 , new_n3013 , new_n3014 );
  nand g02639 ( new_n3016 , pi190 , pi225 );
  nand g02640 ( new_n3017 , pi092 , pi101 );
  nand g02641 ( new_n3018 , new_n3016 , new_n3017 );
  nand g02642 ( new_n3019 , pi092 , pi225 );
  or   g02643 ( new_n3020 , new_n2979 , new_n3019 );
  nand g02644 ( new_n3021 , new_n3018 , new_n3020 );
  xnor g02645 ( new_n3022 , new_n3015 , new_n3021 );
  xnor g02646 ( new_n3023 , new_n3012 , new_n3022 );
  nand g02647 ( new_n3024 , new_n2984 , new_n2991 );
  nand g02648 ( new_n3025 , new_n2983 , new_n2992 );
  nand g02649 ( new_n3026 , new_n3024 , new_n3025 );
  xor  g02650 ( new_n3027 , new_n3023 , new_n3026 );
  nand g02651 ( new_n3028 , pi060 , pi067 );
  nand g02652 ( new_n3029 , pi020 , pi053 );
  nand g02653 ( new_n3030 , new_n3028 , new_n3029 );
  nand g02654 ( new_n3031 , pi053 , pi060 );
  nor  g02655 ( new_n3032 , new_n2984 , new_n3031 );
  not  g02656 ( new_n3033 , new_n3032 );
  nand g02657 ( new_n3034 , new_n3030 , new_n3033 );
  xnor g02658 ( new_n3035 , new_n3027 , new_n3034 );
  nand g02659 ( new_n3036 , new_n3011 , new_n3035 );
  nand g02660 ( new_n3037 , new_n3023 , new_n3026 );
  nand g02661 ( new_n3038 , new_n3027 , new_n3034 );
  nand g02662 ( new_n3039 , new_n3037 , new_n3038 );
  nand g02663 ( new_n3040 , new_n3033 , new_n3039 );
  nor  g02664 ( new_n3041 , new_n3023 , new_n3026 );
  nand g02665 ( new_n3042 , new_n3041 , new_n3032 );
  nand g02666 ( new_n3043 , new_n3040 , new_n3042 );
  nand g02667 ( new_n3044 , pi177 , pi190 );
  nand g02668 ( new_n3045 , pi101 , pi229 );
  xor  g02669 ( new_n3046 , new_n3044 , new_n3045 );
  xor  g02670 ( new_n3047 , new_n3019 , new_n3046 );
  nand g02671 ( new_n3048 , pi067 , pi223 );
  xor  g02672 ( new_n3049 , new_n3020 , new_n3048 );
  xor  g02673 ( new_n3050 , new_n3047 , new_n3049 );
  nand g02674 ( new_n3051 , pi030 , pi160 );
  nand g02675 ( new_n3052 , pi020 , pi185 );
  xor  g02676 ( new_n3053 , new_n3051 , new_n3052 );
  xor  g02677 ( new_n3054 , new_n3031 , new_n3053 );
  nor  g02678 ( new_n3055 , new_n3015 , new_n3021 );
  nor  g02679 ( new_n3056 , new_n3012 , new_n3022 );
  nor  g02680 ( new_n3057 , new_n3055 , new_n3056 );
  xor  g02681 ( new_n3058 , new_n3054 , new_n3057 );
  xnor g02682 ( new_n3059 , new_n3050 , new_n3058 );
  xor  g02683 ( new_n3060 , new_n3043 , new_n3059 );
  xnor g02684 ( new_n3061 , new_n3036 , new_n3060 );
  nand g02685 ( new_n3062 , pi160 , pi185 );
  xor  g02686 ( new_n3063 , new_n3006 , new_n3007 );
  not  g02687 ( new_n3064 , new_n3063 );
  not  g02688 ( new_n3065 , new_n3000 );
  not  g02689 ( new_n3066 , new_n2999 );
  nand g02690 ( new_n3067 , pi160 , pi190 );
  nand g02691 ( new_n3068 , new_n3065 , new_n3067 );
  nand g02692 ( new_n3069 , new_n3066 , new_n3068 );
  nand g02693 ( new_n3070 , new_n3001 , new_n3069 );
  nand g02694 ( new_n3071 , new_n3065 , new_n3070 );
  nor  g02695 ( new_n3072 , new_n3064 , new_n3071 );
  xor  g02696 ( new_n3073 , new_n2996 , new_n3009 );
  nand g02697 ( new_n3074 , new_n3072 , new_n3073 );
  nand g02698 ( new_n3075 , new_n3062 , new_n3074 );
  xnor g02699 ( new_n3076 , new_n3011 , new_n3035 );
  xor  g02700 ( new_n3077 , new_n3062 , new_n3074 );
  nand g02701 ( new_n3078 , new_n3076 , new_n3077 );
  nand g02702 ( new_n3079 , new_n3075 , new_n3078 );
  xor  g02703 ( new_n3080 , new_n3061 , new_n3079 );
  xor  g02704 ( new_n3081 , new_n2978 , new_n3080 );
  xor  g02705 ( new_n3082 , new_n2942 , new_n2975 );
  not  g02706 ( new_n3083 , new_n3082 );
  xor  g02707 ( new_n3084 , new_n3076 , new_n3077 );
  or   g02708 ( new_n3085 , new_n3083 , new_n3084 );
  xor  g02709 ( new_n3086 , new_n3072 , new_n3073 );
  xor  g02710 ( new_n3087 , new_n3063 , new_n3071 );
  xor  g02711 ( new_n3088 , new_n2680 , new_n2950 );
  nor  g02712 ( new_n3089 , new_n3067 , new_n3088 );
  nand g02713 ( new_n3090 , pi092 , pi160 );
  nand g02714 ( new_n3091 , pi020 , pi190 );
  xor  g02715 ( new_n3092 , new_n3090 , new_n3091 );
  nand g02716 ( new_n3093 , new_n3089 , new_n3092 );
  xor  g02717 ( new_n3094 , new_n2958 , new_n2960 );
  xor  g02718 ( new_n3095 , new_n3089 , new_n3092 );
  nand g02719 ( new_n3096 , new_n3094 , new_n3095 );
  nand g02720 ( new_n3097 , new_n3093 , new_n3096 );
  nor  g02721 ( new_n3098 , new_n3066 , new_n3068 );
  nor  g02722 ( new_n3099 , new_n3070 , new_n3098 );
  or   g02723 ( new_n3100 , new_n3097 , new_n3099 );
  xor  g02724 ( new_n3101 , new_n2964 , new_n2965 );
  not  g02725 ( new_n3102 , new_n3101 );
  xor  g02726 ( new_n3103 , new_n3097 , new_n3099 );
  nand g02727 ( new_n3104 , new_n3102 , new_n3103 );
  nand g02728 ( new_n3105 , new_n3100 , new_n3104 );
  or   g02729 ( new_n3106 , new_n3087 , new_n3105 );
  xnor g02730 ( new_n3107 , new_n2948 , new_n2967 );
  xor  g02731 ( new_n3108 , new_n3087 , new_n3105 );
  nand g02732 ( new_n3109 , new_n3107 , new_n3108 );
  nand g02733 ( new_n3110 , new_n3106 , new_n3109 );
  nand g02734 ( new_n3111 , new_n3086 , new_n3110 );
  xor  g02735 ( new_n3112 , new_n2971 , new_n2973 );
  xor  g02736 ( new_n3113 , new_n3086 , new_n3110 );
  nand g02737 ( new_n3114 , new_n3112 , new_n3113 );
  nand g02738 ( new_n3115 , new_n3111 , new_n3114 );
  xor  g02739 ( new_n3116 , new_n3083 , new_n3084 );
  nand g02740 ( new_n3117 , new_n3115 , new_n3116 );
  nand g02741 ( new_n3118 , new_n3085 , new_n3117 );
  xor  g02742 ( po007 , new_n3081 , new_n3118 );
  nand g02743 ( new_n3120 , pi230 , pi236 );
  nand g02744 ( new_n3121 , pi173 , pi236 );
  nand g02745 ( new_n3122 , pi109 , pi161 );
  nand g02746 ( new_n3123 , new_n3121 , new_n3122 );
  nand g02747 ( new_n3124 , pi014 , pi241 );
  xor  g02748 ( new_n3125 , new_n3121 , new_n3122 );
  nand g02749 ( new_n3126 , new_n3124 , new_n3125 );
  nand g02750 ( new_n3127 , new_n3123 , new_n3126 );
  xor  g02751 ( new_n3128 , new_n3120 , new_n3127 );
  nand g02752 ( new_n3129 , pi014 , pi161 );
  nand g02753 ( new_n3130 , pi109 , pi141 );
  nand g02754 ( new_n3131 , pi173 , pi241 );
  xor  g02755 ( new_n3132 , new_n3130 , new_n3131 );
  xnor g02756 ( new_n3133 , new_n3129 , new_n3132 );
  xnor g02757 ( new_n3134 , new_n3128 , new_n3133 );
  nand g02758 ( new_n3135 , pi109 , pi236 );
  nor  g02759 ( new_n3136 , new_n3124 , new_n3125 );
  not  g02760 ( new_n3137 , new_n3136 );
  nor  g02761 ( new_n3138 , new_n3135 , new_n3137 );
  xor  g02762 ( new_n3139 , new_n3134 , new_n3138 );
  nand g02763 ( new_n3140 , pi207 , pi212 );
  nand g02764 ( new_n3141 , pi066 , pi213 );
  xor  g02765 ( new_n3142 , new_n3140 , new_n3141 );
  nand g02766 ( new_n3143 , pi104 , pi226 );
  xor  g02767 ( new_n3144 , new_n3142 , new_n3143 );
  nand g02768 ( new_n3145 , pi213 , pi226 );
  nor  g02769 ( new_n3146 , new_n3140 , new_n3145 );
  not  g02770 ( new_n3147 , new_n3146 );
  nor  g02771 ( new_n3148 , new_n3144 , new_n3147 );
  nand g02772 ( new_n3149 , pi066 , pi212 );
  nand g02773 ( new_n3150 , pi104 , pi207 );
  nand g02774 ( new_n3151 , pi013 , pi226 );
  xor  g02775 ( new_n3152 , new_n3150 , new_n3151 );
  xor  g02776 ( new_n3153 , new_n3149 , new_n3152 );
  nand g02777 ( new_n3154 , pi055 , pi213 );
  nand g02778 ( new_n3155 , new_n3140 , new_n3141 );
  nand g02779 ( new_n3156 , new_n3142 , new_n3143 );
  nand g02780 ( new_n3157 , new_n3155 , new_n3156 );
  xor  g02781 ( new_n3158 , new_n3154 , new_n3157 );
  xor  g02782 ( new_n3159 , new_n3153 , new_n3158 );
  not  g02783 ( new_n3160 , new_n3159 );
  xor  g02784 ( new_n3161 , new_n3148 , new_n3160 );
  xor  g02785 ( new_n3162 , new_n3139 , new_n3161 );
  xor  g02786 ( new_n3163 , new_n3144 , new_n3146 );
  nand g02787 ( new_n3164 , pi207 , pi213 );
  nand g02788 ( new_n3165 , pi212 , pi226 );
  nand g02789 ( new_n3166 , new_n3164 , new_n3165 );
  nand g02790 ( new_n3167 , new_n3147 , new_n3166 );
  nand g02791 ( new_n3168 , pi109 , pi241 );
  nand g02792 ( new_n3169 , pi014 , pi236 );
  nand g02793 ( new_n3170 , new_n3168 , new_n3169 );
  or   g02794 ( new_n3171 , new_n3124 , new_n3135 );
  nand g02795 ( new_n3172 , new_n3170 , new_n3171 );
  nand g02796 ( new_n3173 , new_n3167 , new_n3172 );
  nor  g02797 ( new_n3174 , new_n3135 , new_n3145 );
  not  g02798 ( new_n3175 , new_n3174 );
  xor  g02799 ( new_n3176 , new_n3167 , new_n3172 );
  nand g02800 ( new_n3177 , new_n3175 , new_n3176 );
  nand g02801 ( new_n3178 , new_n3173 , new_n3177 );
  nand g02802 ( new_n3179 , new_n3163 , new_n3178 );
  xor  g02803 ( new_n3180 , new_n3163 , new_n3178 );
  not  g02804 ( new_n3181 , new_n3138 );
  nand g02805 ( new_n3182 , new_n3126 , new_n3171 );
  or   g02806 ( new_n3183 , new_n3136 , new_n3182 );
  nand g02807 ( new_n3184 , new_n3181 , new_n3183 );
  nand g02808 ( new_n3185 , new_n3180 , new_n3184 );
  nand g02809 ( new_n3186 , new_n3179 , new_n3185 );
  xor  g02810 ( new_n3187 , new_n3162 , new_n3186 );
  nand g02811 ( new_n3188 , pi186 , pi208 );
  nand g02812 ( new_n3189 , pi058 , pi168 );
  xor  g02813 ( new_n3190 , new_n3188 , new_n3189 );
  nand g02814 ( new_n3191 , pi132 , pi139 );
  xor  g02815 ( new_n3192 , new_n3190 , new_n3191 );
  nand g02816 ( new_n3193 , pi132 , pi168 );
  or   g02817 ( new_n3194 , new_n3188 , new_n3193 );
  or   g02818 ( new_n3195 , new_n3192 , new_n3194 );
  nand g02819 ( new_n3196 , pi168 , pi211 );
  nand g02820 ( new_n3197 , new_n3188 , new_n3189 );
  nand g02821 ( new_n3198 , new_n3190 , new_n3191 );
  nand g02822 ( new_n3199 , new_n3197 , new_n3198 );
  xor  g02823 ( new_n3200 , new_n3196 , new_n3199 );
  nand g02824 ( new_n3201 , pi035 , pi132 );
  nand g02825 ( new_n3202 , pi058 , pi208 );
  nand g02826 ( new_n3203 , pi139 , pi186 );
  xor  g02827 ( new_n3204 , new_n3202 , new_n3203 );
  xnor g02828 ( new_n3205 , new_n3201 , new_n3204 );
  xnor g02829 ( new_n3206 , new_n3200 , new_n3205 );
  xor  g02830 ( new_n3207 , new_n3195 , new_n3206 );
  xor  g02831 ( new_n3208 , new_n3192 , new_n3194 );
  xor  g02832 ( new_n3209 , new_n3135 , new_n3145 );
  not  g02833 ( new_n3210 , new_n3209 );
  nor  g02834 ( new_n3211 , new_n3193 , new_n3210 );
  not  g02835 ( new_n3212 , new_n3211 );
  nand g02836 ( new_n3213 , pi168 , pi186 );
  nand g02837 ( new_n3214 , pi132 , pi208 );
  nand g02838 ( new_n3215 , new_n3213 , new_n3214 );
  nand g02839 ( new_n3216 , new_n3194 , new_n3215 );
  or   g02840 ( new_n3217 , new_n3212 , new_n3216 );
  xor  g02841 ( new_n3218 , new_n3174 , new_n3176 );
  xor  g02842 ( new_n3219 , new_n3212 , new_n3216 );
  nand g02843 ( new_n3220 , new_n3218 , new_n3219 );
  nand g02844 ( new_n3221 , new_n3217 , new_n3220 );
  nand g02845 ( new_n3222 , new_n3208 , new_n3221 );
  xnor g02846 ( new_n3223 , new_n3180 , new_n3184 );
  xor  g02847 ( new_n3224 , new_n3208 , new_n3221 );
  nand g02848 ( new_n3225 , new_n3223 , new_n3224 );
  nand g02849 ( new_n3226 , new_n3222 , new_n3225 );
  xor  g02850 ( new_n3227 , new_n3207 , new_n3226 );
  xor  g02851 ( new_n3228 , new_n3187 , new_n3227 );
  nand g02852 ( new_n3229 , pi052 , pi069 );
  nand g02853 ( new_n3230 , pi131 , pi244 );
  xor  g02854 ( new_n3231 , new_n3229 , new_n3230 );
  nand g02855 ( new_n3232 , pi029 , pi077 );
  xor  g02856 ( new_n3233 , new_n3231 , new_n3232 );
  nand g02857 ( new_n3234 , pi029 , pi131 );
  nor  g02858 ( new_n3235 , new_n3229 , new_n3234 );
  not  g02859 ( new_n3236 , new_n3235 );
  nor  g02860 ( new_n3237 , new_n3233 , new_n3236 );
  nand g02861 ( new_n3238 , pi029 , pi133 );
  nand g02862 ( new_n3239 , pi052 , pi244 );
  nand g02863 ( new_n3240 , pi069 , pi077 );
  xor  g02864 ( new_n3241 , new_n3239 , new_n3240 );
  xor  g02865 ( new_n3242 , new_n3238 , new_n3241 );
  nand g02866 ( new_n3243 , pi131 , pi150 );
  nand g02867 ( new_n3244 , new_n3229 , new_n3230 );
  nand g02868 ( new_n3245 , new_n3231 , new_n3232 );
  nand g02869 ( new_n3246 , new_n3244 , new_n3245 );
  xor  g02870 ( new_n3247 , new_n3243 , new_n3246 );
  xor  g02871 ( new_n3248 , new_n3242 , new_n3247 );
  xor  g02872 ( new_n3249 , new_n3237 , new_n3248 );
  xor  g02873 ( new_n3250 , new_n3233 , new_n3235 );
  xor  g02874 ( new_n3251 , new_n3193 , new_n3209 );
  nor  g02875 ( new_n3252 , new_n3234 , new_n3251 );
  not  g02876 ( new_n3253 , new_n3252 );
  nand g02877 ( new_n3254 , pi069 , pi131 );
  nand g02878 ( new_n3255 , pi029 , pi052 );
  nand g02879 ( new_n3256 , new_n3254 , new_n3255 );
  nand g02880 ( new_n3257 , new_n3236 , new_n3256 );
  nand g02881 ( new_n3258 , new_n3253 , new_n3257 );
  xnor g02882 ( new_n3259 , new_n3218 , new_n3219 );
  xor  g02883 ( new_n3260 , new_n3253 , new_n3257 );
  nand g02884 ( new_n3261 , new_n3259 , new_n3260 );
  nand g02885 ( new_n3262 , new_n3258 , new_n3261 );
  nand g02886 ( new_n3263 , new_n3250 , new_n3262 );
  xor  g02887 ( new_n3264 , new_n3223 , new_n3224 );
  not  g02888 ( new_n3265 , new_n3264 );
  xor  g02889 ( new_n3266 , new_n3250 , new_n3262 );
  nand g02890 ( new_n3267 , new_n3265 , new_n3266 );
  nand g02891 ( new_n3268 , new_n3263 , new_n3267 );
  xor  g02892 ( new_n3269 , new_n3249 , new_n3268 );
  xor  g02893 ( po008 , new_n3228 , new_n3269 );
  nand g02894 ( new_n3271 , pi013 , pi170 );
  nand g02895 ( new_n3272 , pi073 , pi212 );
  nand g02896 ( new_n3273 , pi004 , pi104 );
  xor  g02897 ( new_n3274 , new_n3272 , new_n3273 );
  xor  g02898 ( new_n3275 , new_n3271 , new_n3274 );
  nand g02899 ( new_n3276 , pi003 , pi213 );
  nand g02900 ( new_n3277 , pi104 , pi170 );
  nand g02901 ( new_n3278 , pi073 , pi213 );
  nand g02902 ( new_n3279 , new_n3277 , new_n3278 );
  nand g02903 ( new_n3280 , pi004 , pi212 );
  or   g02904 ( new_n3281 , new_n3277 , new_n3278 );
  nand g02905 ( new_n3282 , new_n3280 , new_n3281 );
  nand g02906 ( new_n3283 , new_n3279 , new_n3282 );
  xor  g02907 ( new_n3284 , new_n3276 , new_n3283 );
  xor  g02908 ( new_n3285 , new_n3275 , new_n3284 );
  not  g02909 ( new_n3286 , new_n3280 );
  not  g02910 ( new_n3287 , new_n3279 );
  nand g02911 ( new_n3288 , pi170 , pi213 );
  nand g02912 ( new_n3289 , new_n3286 , new_n3288 );
  nand g02913 ( new_n3290 , new_n3287 , new_n3289 );
  nand g02914 ( new_n3291 , new_n3281 , new_n3290 );
  nand g02915 ( new_n3292 , new_n3286 , new_n3291 );
  nor  g02916 ( new_n3293 , new_n3285 , new_n3292 );
  nand g02917 ( new_n3294 , pi073 , pi104 );
  nand g02918 ( new_n3295 , pi112 , pi170 );
  nand g02919 ( new_n3296 , pi004 , pi013 );
  xor  g02920 ( new_n3297 , new_n3295 , new_n3296 );
  xor  g02921 ( new_n3298 , new_n3294 , new_n3297 );
  nand g02922 ( new_n3299 , pi003 , pi212 );
  nand g02923 ( new_n3300 , new_n3272 , new_n3273 );
  nand g02924 ( new_n3301 , new_n3271 , new_n3274 );
  nand g02925 ( new_n3302 , new_n3300 , new_n3301 );
  xor  g02926 ( new_n3303 , new_n3299 , new_n3302 );
  xnor g02927 ( new_n3304 , new_n3298 , new_n3303 );
  nand g02928 ( new_n3305 , pi130 , pi213 );
  or   g02929 ( new_n3306 , new_n3276 , new_n3283 );
  not  g02930 ( new_n3307 , new_n3275 );
  nand g02931 ( new_n3308 , new_n3307 , new_n3284 );
  nand g02932 ( new_n3309 , new_n3306 , new_n3308 );
  xor  g02933 ( new_n3310 , new_n3305 , new_n3309 );
  xor  g02934 ( new_n3311 , new_n3304 , new_n3310 );
  xor  g02935 ( new_n3312 , new_n3293 , new_n3311 );
  nand g02936 ( new_n3313 , pi158 , pi241 );
  nand g02937 ( new_n3314 , pi089 , pi236 );
  xor  g02938 ( new_n3315 , new_n3313 , new_n3314 );
  nand g02939 ( new_n3316 , pi161 , pi254 );
  xor  g02940 ( new_n3317 , new_n3315 , new_n3316 );
  nand g02941 ( new_n3318 , pi236 , pi254 );
  or   g02942 ( new_n3319 , new_n3313 , new_n3318 );
  or   g02943 ( new_n3320 , new_n3317 , new_n3319 );
  nand g02944 ( new_n3321 , pi154 , pi236 );
  nand g02945 ( new_n3322 , new_n3313 , new_n3314 );
  nand g02946 ( new_n3323 , new_n3315 , new_n3316 );
  nand g02947 ( new_n3324 , new_n3322 , new_n3323 );
  xor  g02948 ( new_n3325 , new_n3321 , new_n3324 );
  nand g02949 ( new_n3326 , pi158 , pi161 );
  nand g02950 ( new_n3327 , pi089 , pi241 );
  nand g02951 ( new_n3328 , pi141 , pi254 );
  xor  g02952 ( new_n3329 , new_n3327 , new_n3328 );
  xnor g02953 ( new_n3330 , new_n3326 , new_n3329 );
  xnor g02954 ( new_n3331 , new_n3325 , new_n3330 );
  nor  g02955 ( new_n3332 , new_n3320 , new_n3331 );
  nand g02956 ( new_n3333 , pi141 , pi158 );
  nand g02957 ( new_n3334 , pi089 , pi161 );
  nand g02958 ( new_n3335 , pi090 , pi254 );
  xor  g02959 ( new_n3336 , new_n3334 , new_n3335 );
  xor  g02960 ( new_n3337 , new_n3333 , new_n3336 );
  nand g02961 ( new_n3338 , pi154 , pi241 );
  nand g02962 ( new_n3339 , new_n3327 , new_n3328 );
  nand g02963 ( new_n3340 , new_n3326 , new_n3329 );
  nand g02964 ( new_n3341 , new_n3339 , new_n3340 );
  xor  g02965 ( new_n3342 , new_n3338 , new_n3341 );
  xor  g02966 ( new_n3343 , new_n3337 , new_n3342 );
  nand g02967 ( new_n3344 , pi095 , pi236 );
  or   g02968 ( new_n3345 , new_n3321 , new_n3324 );
  nand g02969 ( new_n3346 , new_n3325 , new_n3330 );
  nand g02970 ( new_n3347 , new_n3345 , new_n3346 );
  xor  g02971 ( new_n3348 , new_n3344 , new_n3347 );
  xor  g02972 ( new_n3349 , new_n3343 , new_n3348 );
  xor  g02973 ( new_n3350 , new_n3332 , new_n3349 );
  xor  g02974 ( new_n3351 , new_n3320 , new_n3331 );
  xor  g02975 ( new_n3352 , new_n3285 , new_n3292 );
  nand g02976 ( new_n3353 , new_n3351 , new_n3352 );
  xor  g02977 ( new_n3354 , new_n3351 , new_n3352 );
  xor  g02978 ( new_n3355 , new_n3317 , new_n3319 );
  nor  g02979 ( new_n3356 , new_n3287 , new_n3289 );
  nor  g02980 ( new_n3357 , new_n3291 , new_n3356 );
  nand g02981 ( new_n3358 , new_n3355 , new_n3357 );
  nand g02982 ( new_n3359 , pi004 , pi213 );
  nand g02983 ( new_n3360 , pi170 , pi212 );
  xor  g02984 ( new_n3361 , new_n3359 , new_n3360 );
  not  g02985 ( new_n3362 , new_n3361 );
  nand g02986 ( new_n3363 , pi158 , pi236 );
  nand g02987 ( new_n3364 , pi241 , pi254 );
  nand g02988 ( new_n3365 , new_n3363 , new_n3364 );
  nand g02989 ( new_n3366 , new_n3319 , new_n3365 );
  nand g02990 ( new_n3367 , new_n3362 , new_n3366 );
  not  g02991 ( new_n3368 , new_n3367 );
  nor  g02992 ( new_n3369 , new_n3288 , new_n3318 );
  xor  g02993 ( new_n3370 , new_n3361 , new_n3366 );
  nor  g02994 ( new_n3371 , new_n3369 , new_n3370 );
  nor  g02995 ( new_n3372 , new_n3368 , new_n3371 );
  xor  g02996 ( new_n3373 , new_n3355 , new_n3357 );
  nand g02997 ( new_n3374 , new_n3372 , new_n3373 );
  nand g02998 ( new_n3375 , new_n3358 , new_n3374 );
  nand g02999 ( new_n3376 , new_n3354 , new_n3375 );
  nand g03000 ( new_n3377 , new_n3353 , new_n3376 );
  xor  g03001 ( new_n3378 , new_n3350 , new_n3377 );
  xnor g03002 ( new_n3379 , new_n3312 , new_n3378 );
  nand g03003 ( new_n3380 , pi062 , pi208 );
  nand g03004 ( new_n3381 , pi120 , pi168 );
  xor  g03005 ( new_n3382 , new_n3380 , new_n3381 );
  nand g03006 ( new_n3383 , pi065 , pi139 );
  xor  g03007 ( new_n3384 , new_n3382 , new_n3383 );
  nand g03008 ( new_n3385 , pi065 , pi168 );
  nor  g03009 ( new_n3386 , new_n3380 , new_n3385 );
  not  g03010 ( new_n3387 , new_n3386 );
  nor  g03011 ( new_n3388 , new_n3384 , new_n3387 );
  not  g03012 ( new_n3389 , new_n3388 );
  nand g03013 ( new_n3390 , pi168 , pi172 );
  nand g03014 ( new_n3391 , new_n3380 , new_n3381 );
  nand g03015 ( new_n3392 , new_n3382 , new_n3383 );
  nand g03016 ( new_n3393 , new_n3391 , new_n3392 );
  xor  g03017 ( new_n3394 , new_n3390 , new_n3393 );
  nand g03018 ( new_n3395 , pi120 , pi208 );
  nand g03019 ( new_n3396 , pi035 , pi065 );
  nand g03020 ( new_n3397 , pi062 , pi139 );
  xor  g03021 ( new_n3398 , new_n3396 , new_n3397 );
  xnor g03022 ( new_n3399 , new_n3395 , new_n3398 );
  xnor g03023 ( new_n3400 , new_n3394 , new_n3399 );
  nor  g03024 ( new_n3401 , new_n3389 , new_n3400 );
  nand g03025 ( new_n3402 , pi120 , pi139 );
  nand g03026 ( new_n3403 , pi035 , pi062 );
  nand g03027 ( new_n3404 , pi015 , pi065 );
  xor  g03028 ( new_n3405 , new_n3403 , new_n3404 );
  xor  g03029 ( new_n3406 , new_n3402 , new_n3405 );
  nand g03030 ( new_n3407 , pi172 , pi208 );
  nand g03031 ( new_n3408 , new_n3396 , new_n3397 );
  nand g03032 ( new_n3409 , new_n3395 , new_n3398 );
  nand g03033 ( new_n3410 , new_n3408 , new_n3409 );
  xor  g03034 ( new_n3411 , new_n3407 , new_n3410 );
  xor  g03035 ( new_n3412 , new_n3406 , new_n3411 );
  nand g03036 ( new_n3413 , pi168 , pi198 );
  or   g03037 ( new_n3414 , new_n3390 , new_n3393 );
  nand g03038 ( new_n3415 , new_n3394 , new_n3399 );
  nand g03039 ( new_n3416 , new_n3414 , new_n3415 );
  xor  g03040 ( new_n3417 , new_n3413 , new_n3416 );
  xor  g03041 ( new_n3418 , new_n3412 , new_n3417 );
  xnor g03042 ( new_n3419 , new_n3401 , new_n3418 );
  xor  g03043 ( new_n3420 , new_n3389 , new_n3400 );
  xor  g03044 ( new_n3421 , new_n3354 , new_n3375 );
  or   g03045 ( new_n3422 , new_n3420 , new_n3421 );
  xor  g03046 ( new_n3423 , new_n3372 , new_n3373 );
  xor  g03047 ( new_n3424 , new_n3384 , new_n3387 );
  nor  g03048 ( new_n3425 , new_n3423 , new_n3424 );
  xnor g03049 ( new_n3426 , new_n3423 , new_n3424 );
  xor  g03050 ( new_n3427 , new_n3288 , new_n3318 );
  not  g03051 ( new_n3428 , new_n3427 );
  or   g03052 ( new_n3429 , new_n3385 , new_n3428 );
  nand g03053 ( new_n3430 , pi062 , pi168 );
  nand g03054 ( new_n3431 , pi065 , pi208 );
  nand g03055 ( new_n3432 , new_n3430 , new_n3431 );
  nand g03056 ( new_n3433 , new_n3387 , new_n3432 );
  or   g03057 ( new_n3434 , new_n3429 , new_n3433 );
  xor  g03058 ( new_n3435 , new_n3369 , new_n3370 );
  not  g03059 ( new_n3436 , new_n3435 );
  xor  g03060 ( new_n3437 , new_n3429 , new_n3433 );
  nand g03061 ( new_n3438 , new_n3436 , new_n3437 );
  nand g03062 ( new_n3439 , new_n3434 , new_n3438 );
  nor  g03063 ( new_n3440 , new_n3426 , new_n3439 );
  or   g03064 ( new_n3441 , new_n3425 , new_n3440 );
  xor  g03065 ( new_n3442 , new_n3420 , new_n3421 );
  nand g03066 ( new_n3443 , new_n3441 , new_n3442 );
  nand g03067 ( new_n3444 , new_n3422 , new_n3443 );
  xor  g03068 ( new_n3445 , new_n3419 , new_n3444 );
  xor  g03069 ( new_n3446 , new_n3379 , new_n3445 );
  nand g03070 ( new_n3447 , pi052 , pi092 );
  nand g03071 ( new_n3448 , pi131 , pi229 );
  xor  g03072 ( new_n3449 , new_n3447 , new_n3448 );
  nand g03073 ( new_n3450 , pi077 , pi190 );
  xor  g03074 ( new_n3451 , new_n3449 , new_n3450 );
  nand g03075 ( new_n3452 , pi131 , pi190 );
  nor  g03076 ( new_n3453 , new_n3447 , new_n3452 );
  not  g03077 ( new_n3454 , new_n3453 );
  or   g03078 ( new_n3455 , new_n3451 , new_n3454 );
  nand g03079 ( new_n3456 , pi067 , pi131 );
  nand g03080 ( new_n3457 , new_n3447 , new_n3448 );
  nand g03081 ( new_n3458 , new_n3449 , new_n3450 );
  nand g03082 ( new_n3459 , new_n3457 , new_n3458 );
  xor  g03083 ( new_n3460 , new_n3456 , new_n3459 );
  nand g03084 ( new_n3461 , pi052 , pi229 );
  nand g03085 ( new_n3462 , pi133 , pi190 );
  nand g03086 ( new_n3463 , pi077 , pi092 );
  xor  g03087 ( new_n3464 , new_n3462 , new_n3463 );
  xnor g03088 ( new_n3465 , new_n3461 , new_n3464 );
  xnor g03089 ( new_n3466 , new_n3460 , new_n3465 );
  nor  g03090 ( new_n3467 , new_n3455 , new_n3466 );
  nand g03091 ( new_n3468 , pi077 , pi229 );
  nand g03092 ( new_n3469 , pi092 , pi133 );
  nand g03093 ( new_n3470 , pi189 , pi190 );
  xor  g03094 ( new_n3471 , new_n3469 , new_n3470 );
  xor  g03095 ( new_n3472 , new_n3468 , new_n3471 );
  nand g03096 ( new_n3473 , pi052 , pi067 );
  nand g03097 ( new_n3474 , new_n3462 , new_n3463 );
  nand g03098 ( new_n3475 , new_n3461 , new_n3464 );
  nand g03099 ( new_n3476 , new_n3474 , new_n3475 );
  xor  g03100 ( new_n3477 , new_n3473 , new_n3476 );
  xor  g03101 ( new_n3478 , new_n3472 , new_n3477 );
  nand g03102 ( new_n3479 , pi053 , pi131 );
  or   g03103 ( new_n3480 , new_n3456 , new_n3459 );
  nand g03104 ( new_n3481 , new_n3460 , new_n3465 );
  nand g03105 ( new_n3482 , new_n3480 , new_n3481 );
  xor  g03106 ( new_n3483 , new_n3479 , new_n3482 );
  xor  g03107 ( new_n3484 , new_n3478 , new_n3483 );
  xor  g03108 ( new_n3485 , new_n3467 , new_n3484 );
  xor  g03109 ( new_n3486 , new_n3441 , new_n3442 );
  not  g03110 ( new_n3487 , new_n3486 );
  xor  g03111 ( new_n3488 , new_n3455 , new_n3466 );
  nor  g03112 ( new_n3489 , new_n3487 , new_n3488 );
  xor  g03113 ( new_n3490 , new_n3486 , new_n3488 );
  xor  g03114 ( new_n3491 , new_n3451 , new_n3453 );
  xor  g03115 ( new_n3492 , new_n3385 , new_n3427 );
  or   g03116 ( new_n3493 , new_n3452 , new_n3492 );
  nand g03117 ( new_n3494 , pi092 , pi131 );
  nand g03118 ( new_n3495 , pi052 , pi190 );
  nand g03119 ( new_n3496 , new_n3494 , new_n3495 );
  nand g03120 ( new_n3497 , new_n3454 , new_n3496 );
  nand g03121 ( new_n3498 , new_n3493 , new_n3497 );
  xor  g03122 ( new_n3499 , new_n3436 , new_n3437 );
  not  g03123 ( new_n3500 , new_n3499 );
  xor  g03124 ( new_n3501 , new_n3493 , new_n3497 );
  nand g03125 ( new_n3502 , new_n3500 , new_n3501 );
  nand g03126 ( new_n3503 , new_n3498 , new_n3502 );
  or   g03127 ( new_n3504 , new_n3491 , new_n3503 );
  xnor g03128 ( new_n3505 , new_n3426 , new_n3439 );
  xor  g03129 ( new_n3506 , new_n3491 , new_n3503 );
  nand g03130 ( new_n3507 , new_n3505 , new_n3506 );
  nand g03131 ( new_n3508 , new_n3504 , new_n3507 );
  nor  g03132 ( new_n3509 , new_n3490 , new_n3508 );
  nor  g03133 ( new_n3510 , new_n3489 , new_n3509 );
  xor  g03134 ( new_n3511 , new_n3485 , new_n3510 );
  xor  g03135 ( po009 , new_n3446 , new_n3511 );
  nand g03136 ( new_n3513 , pi051 , pi236 );
  nand g03137 ( new_n3514 , pi188 , pi213 );
  xor  g03138 ( new_n3515 , new_n3513 , new_n3514 );
  nand g03139 ( new_n3516 , pi162 , pi168 );
  xor  g03140 ( new_n3517 , new_n3515 , new_n3516 );
  nand g03141 ( new_n3518 , pi131 , pi143 );
  xor  g03142 ( po010 , new_n3517 , new_n3518 );
  xor  g03143 ( po011 , new_n1825 , new_n1827 );
  xnor g03144 ( po012 , new_n3490 , new_n3508 );
  nand g03145 ( new_n3522 , pi223 , pi244 );
  nand g03146 ( new_n3523 , pi069 , pi101 );
  nand g03147 ( new_n3524 , pi029 , pi225 );
  nand g03148 ( new_n3525 , new_n3523 , new_n3524 );
  nand g03149 ( new_n3526 , pi029 , pi101 );
  nand g03150 ( new_n3527 , pi069 , pi225 );
  or   g03151 ( new_n3528 , new_n3526 , new_n3527 );
  nand g03152 ( new_n3529 , new_n3525 , new_n3528 );
  xor  g03153 ( new_n3530 , new_n3522 , new_n3529 );
  nand g03154 ( new_n3531 , pi069 , pi223 );
  nand g03155 ( new_n3532 , new_n3526 , new_n3531 );
  nand g03156 ( new_n3533 , pi060 , pi244 );
  xor  g03157 ( new_n3534 , new_n3526 , new_n3531 );
  nand g03158 ( new_n3535 , new_n3533 , new_n3534 );
  nand g03159 ( new_n3536 , new_n3532 , new_n3535 );
  xor  g03160 ( new_n3537 , new_n3530 , new_n3536 );
  nand g03161 ( new_n3538 , pi060 , pi150 );
  nand g03162 ( new_n3539 , pi020 , pi221 );
  nand g03163 ( new_n3540 , new_n3538 , new_n3539 );
  nand g03164 ( new_n3541 , pi020 , pi150 );
  nand g03165 ( new_n3542 , pi060 , pi221 );
  nor  g03166 ( new_n3543 , new_n3541 , new_n3542 );
  not  g03167 ( new_n3544 , new_n3543 );
  nand g03168 ( new_n3545 , new_n3540 , new_n3544 );
  xnor g03169 ( new_n3546 , new_n3537 , new_n3545 );
  nand g03170 ( new_n3547 , pi029 , pi223 );
  nand g03171 ( new_n3548 , pi020 , pi244 );
  nand g03172 ( new_n3549 , new_n3547 , new_n3548 );
  nand g03173 ( new_n3550 , pi060 , pi069 );
  xor  g03174 ( new_n3551 , new_n3547 , new_n3548 );
  nand g03175 ( new_n3552 , new_n3550 , new_n3551 );
  nand g03176 ( new_n3553 , new_n3549 , new_n3552 );
  nand g03177 ( new_n3554 , new_n3541 , new_n3553 );
  xor  g03178 ( new_n3555 , new_n3533 , new_n3534 );
  xor  g03179 ( new_n3556 , new_n3541 , new_n3553 );
  nand g03180 ( new_n3557 , new_n3555 , new_n3556 );
  nand g03181 ( new_n3558 , new_n3554 , new_n3557 );
  xor  g03182 ( new_n3559 , new_n3546 , new_n3558 );
  xor  g03183 ( new_n3560 , new_n3555 , new_n3556 );
  nand g03184 ( new_n3561 , pi160 , pi221 );
  nor  g03185 ( new_n3562 , new_n3560 , new_n3561 );
  xnor g03186 ( new_n3563 , new_n3560 , new_n3561 );
  nand g03187 ( new_n3564 , pi150 , pi160 );
  nand g03188 ( new_n3565 , pi020 , pi069 );
  nand g03189 ( new_n3566 , pi160 , pi244 );
  nand g03190 ( new_n3567 , new_n3565 , new_n3566 );
  nand g03191 ( new_n3568 , pi029 , pi060 );
  xor  g03192 ( new_n3569 , new_n3565 , new_n3566 );
  nand g03193 ( new_n3570 , new_n3568 , new_n3569 );
  nand g03194 ( new_n3571 , new_n3567 , new_n3570 );
  nand g03195 ( new_n3572 , new_n3564 , new_n3571 );
  xor  g03196 ( new_n3573 , new_n3550 , new_n3551 );
  xor  g03197 ( new_n3574 , new_n3564 , new_n3571 );
  nand g03198 ( new_n3575 , new_n3573 , new_n3574 );
  nand g03199 ( new_n3576 , new_n3572 , new_n3575 );
  nor  g03200 ( new_n3577 , new_n3563 , new_n3576 );
  nor  g03201 ( new_n3578 , new_n3562 , new_n3577 );
  not  g03202 ( new_n3579 , new_n3578 );
  nand g03203 ( new_n3580 , new_n3559 , new_n3579 );
  nand g03204 ( new_n3581 , pi029 , pi177 );
  nand g03205 ( new_n3582 , pi101 , pi244 );
  xor  g03206 ( new_n3583 , new_n3581 , new_n3582 );
  xor  g03207 ( new_n3584 , new_n3527 , new_n3583 );
  nand g03208 ( new_n3585 , pi150 , pi223 );
  xor  g03209 ( new_n3586 , new_n3528 , new_n3585 );
  xor  g03210 ( new_n3587 , new_n3584 , new_n3586 );
  nand g03211 ( new_n3588 , pi020 , pi196 );
  nand g03212 ( new_n3589 , pi160 , pi184 );
  xor  g03213 ( new_n3590 , new_n3588 , new_n3589 );
  xor  g03214 ( new_n3591 , new_n3542 , new_n3590 );
  nand g03215 ( new_n3592 , new_n3522 , new_n3529 );
  nand g03216 ( new_n3593 , new_n3530 , new_n3536 );
  nand g03217 ( new_n3594 , new_n3592 , new_n3593 );
  xor  g03218 ( new_n3595 , new_n3591 , new_n3594 );
  xnor g03219 ( new_n3596 , new_n3587 , new_n3595 );
  nor  g03220 ( new_n3597 , new_n3546 , new_n3558 );
  and  g03221 ( new_n3598 , new_n3543 , new_n3597 );
  or   g03222 ( new_n3599 , new_n3537 , new_n3545 );
  nand g03223 ( new_n3600 , new_n3544 , new_n3599 );
  nor  g03224 ( new_n3601 , new_n3597 , new_n3600 );
  or   g03225 ( new_n3602 , new_n3598 , new_n3601 );
  xor  g03226 ( new_n3603 , new_n3596 , new_n3602 );
  xnor g03227 ( new_n3604 , new_n3580 , new_n3603 );
  nand g03228 ( new_n3605 , pi160 , pi196 );
  xor  g03229 ( new_n3606 , new_n3568 , new_n3569 );
  nand g03230 ( new_n3607 , pi029 , pi160 );
  nor  g03231 ( new_n3608 , new_n3565 , new_n3607 );
  not  g03232 ( new_n3609 , new_n3608 );
  nor  g03233 ( new_n3610 , new_n3606 , new_n3609 );
  not  g03234 ( new_n3611 , new_n3610 );
  xor  g03235 ( new_n3612 , new_n3573 , new_n3574 );
  nor  g03236 ( new_n3613 , new_n3611 , new_n3612 );
  xor  g03237 ( new_n3614 , new_n3563 , new_n3576 );
  nand g03238 ( new_n3615 , new_n3613 , new_n3614 );
  nand g03239 ( new_n3616 , new_n3605 , new_n3615 );
  xor  g03240 ( new_n3617 , new_n3559 , new_n3578 );
  xor  g03241 ( new_n3618 , new_n3605 , new_n3615 );
  nand g03242 ( new_n3619 , new_n3617 , new_n3618 );
  nand g03243 ( new_n3620 , new_n3616 , new_n3619 );
  xor  g03244 ( new_n3621 , new_n3604 , new_n3620 );
  xor  g03245 ( new_n3622 , new_n3613 , new_n3614 );
  xor  g03246 ( new_n3623 , new_n3610 , new_n3612 );
  xor  g03247 ( new_n3624 , new_n3606 , new_n3608 );
  nand g03248 ( new_n3625 , pi169 , pi226 );
  nand g03249 ( new_n3626 , pi071 , pi207 );
  nand g03250 ( new_n3627 , pi066 , pi142 );
  xor  g03251 ( new_n3628 , new_n3626 , new_n3627 );
  xor  g03252 ( new_n3629 , new_n3625 , new_n3628 );
  nand g03253 ( new_n3630 , pi142 , pi207 );
  nand g03254 ( new_n3631 , pi071 , pi226 );
  nor  g03255 ( new_n3632 , new_n3630 , new_n3631 );
  xor  g03256 ( new_n3633 , new_n3629 , new_n3632 );
  xor  g03257 ( new_n3634 , new_n3630 , new_n3631 );
  nand g03258 ( new_n3635 , pi142 , pi226 );
  nand g03259 ( new_n3636 , pi087 , pi109 );
  nor  g03260 ( new_n3637 , new_n3635 , new_n3636 );
  nor  g03261 ( new_n3638 , new_n3634 , new_n3637 );
  nand g03262 ( new_n3639 , pi109 , pi219 );
  nand g03263 ( new_n3640 , pi014 , pi087 );
  xor  g03264 ( new_n3641 , new_n3639 , new_n3640 );
  xnor g03265 ( new_n3642 , new_n3634 , new_n3637 );
  nor  g03266 ( new_n3643 , new_n3641 , new_n3642 );
  nor  g03267 ( new_n3644 , new_n3638 , new_n3643 );
  nand g03268 ( new_n3645 , pi087 , pi173 );
  nand g03269 ( new_n3646 , pi102 , pi109 );
  nand g03270 ( new_n3647 , new_n3645 , new_n3646 );
  not  g03271 ( new_n3648 , new_n3647 );
  nand g03272 ( new_n3649 , pi014 , pi219 );
  not  g03273 ( new_n3650 , new_n3649 );
  nand g03274 ( new_n3651 , new_n3636 , new_n3650 );
  nor  g03275 ( new_n3652 , new_n3648 , new_n3651 );
  nand g03276 ( new_n3653 , new_n3648 , new_n3651 );
  or   g03277 ( new_n3654 , new_n3645 , new_n3646 );
  nand g03278 ( new_n3655 , new_n3653 , new_n3654 );
  nor  g03279 ( new_n3656 , new_n3652 , new_n3655 );
  xor  g03280 ( new_n3657 , new_n3644 , new_n3656 );
  xnor g03281 ( new_n3658 , new_n3633 , new_n3657 );
  nand g03282 ( new_n3659 , pi041 , pi132 );
  nand g03283 ( new_n3660 , pi182 , pi186 );
  nand g03284 ( new_n3661 , pi058 , pi138 );
  xor  g03285 ( new_n3662 , new_n3660 , new_n3661 );
  xor  g03286 ( new_n3663 , new_n3659 , new_n3662 );
  nand g03287 ( new_n3664 , pi132 , pi138 );
  or   g03288 ( new_n3665 , new_n3660 , new_n3664 );
  xor  g03289 ( new_n3666 , new_n3663 , new_n3665 );
  xor  g03290 ( new_n3667 , new_n3635 , new_n3636 );
  not  g03291 ( new_n3668 , new_n3667 );
  nor  g03292 ( new_n3669 , new_n3664 , new_n3668 );
  not  g03293 ( new_n3670 , new_n3669 );
  nand g03294 ( new_n3671 , pi138 , pi186 );
  nand g03295 ( new_n3672 , pi132 , pi182 );
  nand g03296 ( new_n3673 , new_n3671 , new_n3672 );
  nand g03297 ( new_n3674 , new_n3665 , new_n3673 );
  or   g03298 ( new_n3675 , new_n3670 , new_n3674 );
  xnor g03299 ( new_n3676 , new_n3641 , new_n3642 );
  xor  g03300 ( new_n3677 , new_n3670 , new_n3674 );
  nand g03301 ( new_n3678 , new_n3676 , new_n3677 );
  nand g03302 ( new_n3679 , new_n3675 , new_n3678 );
  xor  g03303 ( new_n3680 , new_n3666 , new_n3679 );
  xnor g03304 ( new_n3681 , new_n3658 , new_n3680 );
  nand g03305 ( new_n3682 , new_n3624 , new_n3681 );
  xor  g03306 ( new_n3683 , new_n3664 , new_n3667 );
  nor  g03307 ( new_n3684 , new_n3607 , new_n3683 );
  not  g03308 ( new_n3685 , new_n3684 );
  nand g03309 ( new_n3686 , pi020 , pi029 );
  nand g03310 ( new_n3687 , pi069 , pi160 );
  nand g03311 ( new_n3688 , new_n3686 , new_n3687 );
  nand g03312 ( new_n3689 , new_n3609 , new_n3688 );
  nand g03313 ( new_n3690 , new_n3685 , new_n3689 );
  xnor g03314 ( new_n3691 , new_n3676 , new_n3677 );
  xor  g03315 ( new_n3692 , new_n3685 , new_n3689 );
  nand g03316 ( new_n3693 , new_n3691 , new_n3692 );
  nand g03317 ( new_n3694 , new_n3690 , new_n3693 );
  xor  g03318 ( new_n3695 , new_n3624 , new_n3681 );
  nand g03319 ( new_n3696 , new_n3694 , new_n3695 );
  nand g03320 ( new_n3697 , new_n3682 , new_n3696 );
  or   g03321 ( new_n3698 , new_n3623 , new_n3697 );
  or   g03322 ( new_n3699 , new_n3663 , new_n3665 );
  nand g03323 ( new_n3700 , pi058 , pi182 );
  nand g03324 ( new_n3701 , pi132 , pi216 );
  nand g03325 ( new_n3702 , pi041 , pi186 );
  xor  g03326 ( new_n3703 , new_n3701 , new_n3702 );
  xnor g03327 ( new_n3704 , new_n3700 , new_n3703 );
  nand g03328 ( new_n3705 , pi138 , pi211 );
  nand g03329 ( new_n3706 , new_n3660 , new_n3661 );
  nand g03330 ( new_n3707 , new_n3659 , new_n3662 );
  nand g03331 ( new_n3708 , new_n3706 , new_n3707 );
  xor  g03332 ( new_n3709 , new_n3705 , new_n3708 );
  xnor g03333 ( new_n3710 , new_n3704 , new_n3709 );
  xor  g03334 ( new_n3711 , new_n3699 , new_n3710 );
  nand g03335 ( new_n3712 , new_n3649 , new_n3654 );
  nand g03336 ( new_n3713 , new_n3647 , new_n3712 );
  nand g03337 ( new_n3714 , pi087 , pi230 );
  xor  g03338 ( new_n3715 , new_n3713 , new_n3714 );
  nand g03339 ( new_n3716 , pi001 , pi109 );
  nand g03340 ( new_n3717 , pi173 , pi219 );
  nand g03341 ( new_n3718 , pi014 , pi102 );
  xor  g03342 ( new_n3719 , new_n3717 , new_n3718 );
  xnor g03343 ( new_n3720 , new_n3716 , new_n3719 );
  xnor g03344 ( new_n3721 , new_n3715 , new_n3720 );
  nand g03345 ( new_n3722 , new_n3650 , new_n3655 );
  xor  g03346 ( new_n3723 , new_n3721 , new_n3722 );
  not  g03347 ( new_n3724 , new_n3723 );
  not  g03348 ( new_n3725 , new_n3632 );
  nor  g03349 ( new_n3726 , new_n3629 , new_n3725 );
  nand g03350 ( new_n3727 , pi169 , pi207 );
  nand g03351 ( new_n3728 , pi066 , pi071 );
  nand g03352 ( new_n3729 , pi123 , pi226 );
  xor  g03353 ( new_n3730 , new_n3728 , new_n3729 );
  xnor g03354 ( new_n3731 , new_n3727 , new_n3730 );
  nand g03355 ( new_n3732 , pi055 , pi142 );
  nand g03356 ( new_n3733 , new_n3626 , new_n3627 );
  nand g03357 ( new_n3734 , new_n3625 , new_n3628 );
  nand g03358 ( new_n3735 , new_n3733 , new_n3734 );
  xor  g03359 ( new_n3736 , new_n3732 , new_n3735 );
  xnor g03360 ( new_n3737 , new_n3731 , new_n3736 );
  xor  g03361 ( new_n3738 , new_n3726 , new_n3737 );
  or   g03362 ( new_n3739 , new_n3644 , new_n3656 );
  nand g03363 ( new_n3740 , new_n3633 , new_n3657 );
  nand g03364 ( new_n3741 , new_n3739 , new_n3740 );
  xor  g03365 ( new_n3742 , new_n3738 , new_n3741 );
  xor  g03366 ( new_n3743 , new_n3724 , new_n3742 );
  not  g03367 ( new_n3744 , new_n3743 );
  xor  g03368 ( new_n3745 , new_n3711 , new_n3744 );
  nand g03369 ( new_n3746 , new_n3666 , new_n3679 );
  nand g03370 ( new_n3747 , new_n3658 , new_n3680 );
  nand g03371 ( new_n3748 , new_n3746 , new_n3747 );
  xor  g03372 ( new_n3749 , new_n3745 , new_n3748 );
  xor  g03373 ( new_n3750 , new_n3623 , new_n3697 );
  nand g03374 ( new_n3751 , new_n3749 , new_n3750 );
  nand g03375 ( new_n3752 , new_n3698 , new_n3751 );
  or   g03376 ( new_n3753 , new_n3622 , new_n3752 );
  not  g03377 ( new_n3754 , new_n3726 );
  nor  g03378 ( new_n3755 , new_n3754 , new_n3737 );
  nand g03379 ( new_n3756 , pi123 , pi207 );
  nand g03380 ( new_n3757 , pi099 , pi226 );
  nand g03381 ( new_n3758 , pi066 , pi169 );
  xor  g03382 ( new_n3759 , new_n3757 , new_n3758 );
  xor  g03383 ( new_n3760 , new_n3756 , new_n3759 );
  nand g03384 ( new_n3761 , pi055 , pi071 );
  nand g03385 ( new_n3762 , new_n3728 , new_n3729 );
  nand g03386 ( new_n3763 , new_n3727 , new_n3730 );
  nand g03387 ( new_n3764 , new_n3762 , new_n3763 );
  xor  g03388 ( new_n3765 , new_n3761 , new_n3764 );
  xor  g03389 ( new_n3766 , new_n3760 , new_n3765 );
  nand g03390 ( new_n3767 , pi002 , pi142 );
  or   g03391 ( new_n3768 , new_n3732 , new_n3735 );
  nand g03392 ( new_n3769 , new_n3731 , new_n3736 );
  nand g03393 ( new_n3770 , new_n3768 , new_n3769 );
  xor  g03394 ( new_n3771 , new_n3767 , new_n3770 );
  xor  g03395 ( new_n3772 , new_n3766 , new_n3771 );
  xnor g03396 ( new_n3773 , new_n3755 , new_n3772 );
  nor  g03397 ( new_n3774 , new_n3721 , new_n3722 );
  nand g03398 ( new_n3775 , pi050 , pi087 );
  or   g03399 ( new_n3776 , new_n3713 , new_n3714 );
  nand g03400 ( new_n3777 , new_n3715 , new_n3720 );
  nand g03401 ( new_n3778 , new_n3776 , new_n3777 );
  xor  g03402 ( new_n3779 , new_n3775 , new_n3778 );
  nand g03403 ( new_n3780 , pi102 , pi173 );
  nand g03404 ( new_n3781 , pi001 , pi014 );
  nand g03405 ( new_n3782 , pi109 , pi122 );
  xor  g03406 ( new_n3783 , new_n3781 , new_n3782 );
  xor  g03407 ( new_n3784 , new_n3780 , new_n3783 );
  nand g03408 ( new_n3785 , pi219 , pi230 );
  nand g03409 ( new_n3786 , new_n3717 , new_n3718 );
  nand g03410 ( new_n3787 , new_n3716 , new_n3719 );
  nand g03411 ( new_n3788 , new_n3786 , new_n3787 );
  xor  g03412 ( new_n3789 , new_n3785 , new_n3788 );
  xor  g03413 ( new_n3790 , new_n3784 , new_n3789 );
  xor  g03414 ( new_n3791 , new_n3779 , new_n3790 );
  xnor g03415 ( new_n3792 , new_n3774 , new_n3791 );
  nand g03416 ( new_n3793 , new_n3738 , new_n3741 );
  nand g03417 ( new_n3794 , new_n3724 , new_n3742 );
  nand g03418 ( new_n3795 , new_n3793 , new_n3794 );
  xor  g03419 ( new_n3796 , new_n3792 , new_n3795 );
  xnor g03420 ( new_n3797 , new_n3773 , new_n3796 );
  nor  g03421 ( new_n3798 , new_n3699 , new_n3710 );
  nand g03422 ( new_n3799 , pi076 , pi132 );
  nand g03423 ( new_n3800 , pi186 , pi216 );
  nand g03424 ( new_n3801 , pi041 , pi058 );
  xor  g03425 ( new_n3802 , new_n3800 , new_n3801 );
  xor  g03426 ( new_n3803 , new_n3799 , new_n3802 );
  nand g03427 ( new_n3804 , pi182 , pi211 );
  nand g03428 ( new_n3805 , new_n3701 , new_n3702 );
  nand g03429 ( new_n3806 , new_n3700 , new_n3703 );
  nand g03430 ( new_n3807 , new_n3805 , new_n3806 );
  xor  g03431 ( new_n3808 , new_n3804 , new_n3807 );
  xor  g03432 ( new_n3809 , new_n3803 , new_n3808 );
  nand g03433 ( new_n3810 , pi138 , pi199 );
  or   g03434 ( new_n3811 , new_n3705 , new_n3708 );
  nand g03435 ( new_n3812 , new_n3704 , new_n3709 );
  nand g03436 ( new_n3813 , new_n3811 , new_n3812 );
  xor  g03437 ( new_n3814 , new_n3810 , new_n3813 );
  xor  g03438 ( new_n3815 , new_n3809 , new_n3814 );
  xor  g03439 ( new_n3816 , new_n3798 , new_n3815 );
  nor  g03440 ( new_n3817 , new_n3711 , new_n3744 );
  not  g03441 ( new_n3818 , new_n3745 );
  nor  g03442 ( new_n3819 , new_n3818 , new_n3748 );
  nor  g03443 ( new_n3820 , new_n3817 , new_n3819 );
  xor  g03444 ( new_n3821 , new_n3816 , new_n3820 );
  xor  g03445 ( new_n3822 , new_n3797 , new_n3821 );
  not  g03446 ( new_n3823 , new_n3822 );
  xor  g03447 ( new_n3824 , new_n3622 , new_n3752 );
  nand g03448 ( new_n3825 , new_n3823 , new_n3824 );
  nand g03449 ( new_n3826 , new_n3753 , new_n3825 );
  xor  g03450 ( new_n3827 , new_n3617 , new_n3618 );
  or   g03451 ( new_n3828 , new_n3826 , new_n3827 );
  nand g03452 ( new_n3829 , new_n3792 , new_n3795 );
  nand g03453 ( new_n3830 , new_n3773 , new_n3796 );
  nand g03454 ( new_n3831 , new_n3829 , new_n3830 );
  and  g03455 ( new_n3832 , new_n3755 , new_n3772 );
  nand g03456 ( new_n3833 , pi025 , pi142 );
  nand g03457 ( new_n3834 , pi066 , pi123 );
  nand g03458 ( new_n3835 , pi023 , pi226 );
  nand g03459 ( new_n3836 , pi099 , pi207 );
  nand g03460 ( new_n3837 , new_n3835 , new_n3836 );
  nand g03461 ( new_n3838 , pi023 , pi207 );
  or   g03462 ( new_n3839 , new_n3757 , new_n3838 );
  nand g03463 ( new_n3840 , new_n3837 , new_n3839 );
  xor  g03464 ( new_n3841 , new_n3834 , new_n3840 );
  nand g03465 ( new_n3842 , new_n3757 , new_n3758 );
  nand g03466 ( new_n3843 , new_n3756 , new_n3759 );
  nand g03467 ( new_n3844 , new_n3842 , new_n3843 );
  xor  g03468 ( new_n3845 , new_n3841 , new_n3844 );
  nand g03469 ( new_n3846 , new_n3761 , new_n3764 );
  nand g03470 ( new_n3847 , new_n3760 , new_n3765 );
  nand g03471 ( new_n3848 , new_n3846 , new_n3847 );
  nand g03472 ( new_n3849 , pi002 , pi071 );
  nand g03473 ( new_n3850 , pi055 , pi169 );
  nand g03474 ( new_n3851 , new_n3849 , new_n3850 );
  nand g03475 ( new_n3852 , pi002 , pi169 );
  or   g03476 ( new_n3853 , new_n3761 , new_n3852 );
  nand g03477 ( new_n3854 , new_n3851 , new_n3853 );
  xor  g03478 ( new_n3855 , new_n3848 , new_n3854 );
  xor  g03479 ( new_n3856 , new_n3845 , new_n3855 );
  not  g03480 ( new_n3857 , new_n3767 );
  nand g03481 ( new_n3858 , new_n3857 , new_n3770 );
  or   g03482 ( new_n3859 , new_n3766 , new_n3771 );
  nand g03483 ( new_n3860 , new_n3858 , new_n3859 );
  xor  g03484 ( new_n3861 , new_n3856 , new_n3860 );
  xor  g03485 ( new_n3862 , new_n3833 , new_n3861 );
  xor  g03486 ( new_n3863 , new_n3832 , new_n3862 );
  nand g03487 ( new_n3864 , pi001 , pi173 );
  nand g03488 ( new_n3865 , new_n3781 , new_n3782 );
  nand g03489 ( new_n3866 , new_n3780 , new_n3783 );
  nand g03490 ( new_n3867 , new_n3865 , new_n3866 );
  xor  g03491 ( new_n3868 , new_n3864 , new_n3867 );
  nand g03492 ( new_n3869 , pi014 , pi122 );
  nand g03493 ( new_n3870 , pi109 , pi135 );
  nand g03494 ( new_n3871 , new_n3869 , new_n3870 );
  nand g03495 ( new_n3872 , pi014 , pi135 );
  nor  g03496 ( new_n3873 , new_n3782 , new_n3872 );
  not  g03497 ( new_n3874 , new_n3873 );
  nand g03498 ( new_n3875 , new_n3871 , new_n3874 );
  xor  g03499 ( new_n3876 , new_n3868 , new_n3875 );
  nand g03500 ( new_n3877 , pi102 , pi230 );
  nand g03501 ( new_n3878 , pi050 , pi219 );
  and  g03502 ( new_n3879 , new_n3877 , new_n3878 );
  nand g03503 ( new_n3880 , pi050 , pi102 );
  nor  g03504 ( new_n3881 , new_n3785 , new_n3880 );
  or   g03505 ( new_n3882 , new_n3879 , new_n3881 );
  xnor g03506 ( new_n3883 , new_n3876 , new_n3882 );
  nand g03507 ( new_n3884 , new_n3785 , new_n3788 );
  nand g03508 ( new_n3885 , new_n3784 , new_n3789 );
  nand g03509 ( new_n3886 , new_n3884 , new_n3885 );
  xor  g03510 ( new_n3887 , new_n3883 , new_n3886 );
  not  g03511 ( new_n3888 , new_n3775 );
  nand g03512 ( new_n3889 , new_n3888 , new_n3778 );
  or   g03513 ( new_n3890 , new_n3779 , new_n3790 );
  nand g03514 ( new_n3891 , new_n3889 , new_n3890 );
  xnor g03515 ( new_n3892 , new_n3887 , new_n3891 );
  nand g03516 ( new_n3893 , new_n3774 , new_n3791 );
  nand g03517 ( new_n3894 , pi087 , pi253 );
  xor  g03518 ( new_n3895 , new_n3893 , new_n3894 );
  xor  g03519 ( new_n3896 , new_n3892 , new_n3895 );
  xor  g03520 ( new_n3897 , new_n3863 , new_n3896 );
  xor  g03521 ( new_n3898 , new_n3831 , new_n3897 );
  nand g03522 ( new_n3899 , new_n3798 , new_n3815 );
  nand g03523 ( new_n3900 , pi138 , pi195 );
  nand g03524 ( new_n3901 , pi058 , pi216 );
  nand g03525 ( new_n3902 , pi076 , pi186 );
  nand g03526 ( new_n3903 , pi079 , pi132 );
  nand g03527 ( new_n3904 , new_n3902 , new_n3903 );
  nand g03528 ( new_n3905 , pi079 , pi186 );
  or   g03529 ( new_n3906 , new_n3799 , new_n3905 );
  nand g03530 ( new_n3907 , new_n3904 , new_n3906 );
  xor  g03531 ( new_n3908 , new_n3901 , new_n3907 );
  nand g03532 ( new_n3909 , new_n3800 , new_n3801 );
  nand g03533 ( new_n3910 , new_n3799 , new_n3802 );
  nand g03534 ( new_n3911 , new_n3909 , new_n3910 );
  xor  g03535 ( new_n3912 , new_n3908 , new_n3911 );
  nand g03536 ( new_n3913 , pi041 , pi211 );
  nand g03537 ( new_n3914 , pi182 , pi199 );
  nand g03538 ( new_n3915 , new_n3913 , new_n3914 );
  nand g03539 ( new_n3916 , pi041 , pi199 );
  nor  g03540 ( new_n3917 , new_n3804 , new_n3916 );
  not  g03541 ( new_n3918 , new_n3917 );
  nand g03542 ( new_n3919 , new_n3915 , new_n3918 );
  xnor g03543 ( new_n3920 , new_n3912 , new_n3919 );
  nand g03544 ( new_n3921 , new_n3804 , new_n3807 );
  nand g03545 ( new_n3922 , new_n3803 , new_n3808 );
  nand g03546 ( new_n3923 , new_n3921 , new_n3922 );
  xor  g03547 ( new_n3924 , new_n3920 , new_n3923 );
  not  g03548 ( new_n3925 , new_n3810 );
  nand g03549 ( new_n3926 , new_n3925 , new_n3813 );
  or   g03550 ( new_n3927 , new_n3809 , new_n3814 );
  nand g03551 ( new_n3928 , new_n3926 , new_n3927 );
  xnor g03552 ( new_n3929 , new_n3924 , new_n3928 );
  xor  g03553 ( new_n3930 , new_n3900 , new_n3929 );
  not  g03554 ( new_n3931 , new_n3930 );
  xor  g03555 ( new_n3932 , new_n3899 , new_n3931 );
  nand g03556 ( new_n3933 , new_n3816 , new_n3820 );
  nand g03557 ( new_n3934 , new_n3797 , new_n3821 );
  nand g03558 ( new_n3935 , new_n3933 , new_n3934 );
  xor  g03559 ( new_n3936 , new_n3932 , new_n3935 );
  xor  g03560 ( new_n3937 , new_n3898 , new_n3936 );
  xor  g03561 ( new_n3938 , new_n3826 , new_n3827 );
  nand g03562 ( new_n3939 , new_n3937 , new_n3938 );
  nand g03563 ( new_n3940 , new_n3828 , new_n3939 );
  nand g03564 ( new_n3941 , new_n3621 , new_n3940 );
  not  g03565 ( new_n3942 , new_n3856 );
  nand g03566 ( new_n3943 , new_n3942 , new_n3860 );
  nand g03567 ( new_n3944 , pi066 , pi099 );
  nand g03568 ( new_n3945 , pi155 , pi226 );
  xor  g03569 ( new_n3946 , new_n3838 , new_n3945 );
  xor  g03570 ( new_n3947 , new_n3944 , new_n3946 );
  nand g03571 ( new_n3948 , pi055 , pi123 );
  xor  g03572 ( new_n3949 , new_n3839 , new_n3948 );
  xor  g03573 ( new_n3950 , new_n3947 , new_n3949 );
  nand g03574 ( new_n3951 , pi025 , pi071 );
  nand g03575 ( new_n3952 , pi142 , pi239 );
  xor  g03576 ( new_n3953 , new_n3951 , new_n3952 );
  xor  g03577 ( new_n3954 , new_n3852 , new_n3953 );
  nand g03578 ( new_n3955 , new_n3834 , new_n3840 );
  nand g03579 ( new_n3956 , new_n3841 , new_n3844 );
  nand g03580 ( new_n3957 , new_n3955 , new_n3956 );
  xor  g03581 ( new_n3958 , new_n3954 , new_n3957 );
  xor  g03582 ( new_n3959 , new_n3950 , new_n3958 );
  nand g03583 ( new_n3960 , new_n3848 , new_n3854 );
  nand g03584 ( new_n3961 , new_n3845 , new_n3855 );
  nand g03585 ( new_n3962 , new_n3960 , new_n3961 );
  xor  g03586 ( new_n3963 , new_n3853 , new_n3962 );
  xor  g03587 ( new_n3964 , new_n3959 , new_n3963 );
  xor  g03588 ( new_n3965 , new_n3943 , new_n3964 );
  or   g03589 ( new_n3966 , new_n3833 , new_n3861 );
  nand g03590 ( new_n3967 , new_n3832 , new_n3862 );
  nand g03591 ( new_n3968 , new_n3966 , new_n3967 );
  xor  g03592 ( new_n3969 , new_n3965 , new_n3968 );
  nand g03593 ( new_n3970 , new_n3887 , new_n3891 );
  nand g03594 ( new_n3971 , pi122 , pi173 );
  nand g03595 ( new_n3972 , pi059 , pi109 );
  xor  g03596 ( new_n3973 , new_n3971 , new_n3972 );
  xor  g03597 ( new_n3974 , new_n3872 , new_n3973 );
  nand g03598 ( new_n3975 , pi001 , pi230 );
  xor  g03599 ( new_n3976 , new_n3874 , new_n3975 );
  not  g03600 ( new_n3977 , new_n3976 );
  xor  g03601 ( new_n3978 , new_n3974 , new_n3977 );
  nand g03602 ( new_n3979 , pi074 , pi087 );
  nand g03603 ( new_n3980 , pi219 , pi253 );
  xor  g03604 ( new_n3981 , new_n3979 , new_n3980 );
  xor  g03605 ( new_n3982 , new_n3880 , new_n3981 );
  nand g03606 ( new_n3983 , new_n3864 , new_n3867 );
  nand g03607 ( new_n3984 , new_n3868 , new_n3875 );
  nand g03608 ( new_n3985 , new_n3983 , new_n3984 );
  xor  g03609 ( new_n3986 , new_n3982 , new_n3985 );
  xor  g03610 ( new_n3987 , new_n3978 , new_n3986 );
  nor  g03611 ( new_n3988 , new_n3876 , new_n3882 );
  nor  g03612 ( new_n3989 , new_n3883 , new_n3886 );
  xor  g03613 ( new_n3990 , new_n3881 , new_n3989 );
  nor  g03614 ( new_n3991 , new_n3988 , new_n3990 );
  not  g03615 ( new_n3992 , new_n3991 );
  xor  g03616 ( new_n3993 , new_n3987 , new_n3992 );
  xor  g03617 ( new_n3994 , new_n3970 , new_n3993 );
  nand g03618 ( new_n3995 , new_n3893 , new_n3894 );
  nand g03619 ( new_n3996 , new_n3892 , new_n3895 );
  nand g03620 ( new_n3997 , new_n3995 , new_n3996 );
  xor  g03621 ( new_n3998 , new_n3994 , new_n3997 );
  xor  g03622 ( new_n3999 , new_n3969 , new_n3998 );
  not  g03623 ( new_n4000 , new_n3863 );
  nor  g03624 ( new_n4001 , new_n4000 , new_n3896 );
  nor  g03625 ( new_n4002 , new_n3831 , new_n3897 );
  nor  g03626 ( new_n4003 , new_n4001 , new_n4002 );
  not  g03627 ( new_n4004 , new_n4003 );
  xor  g03628 ( new_n4005 , new_n3999 , new_n4004 );
  nand g03629 ( new_n4006 , new_n3924 , new_n3928 );
  nand g03630 ( new_n4007 , pi132 , pi251 );
  nand g03631 ( new_n4008 , pi058 , pi076 );
  xor  g03632 ( new_n4009 , new_n3905 , new_n4008 );
  xor  g03633 ( new_n4010 , new_n4007 , new_n4009 );
  nand g03634 ( new_n4011 , pi211 , pi216 );
  xor  g03635 ( new_n4012 , new_n3906 , new_n4011 );
  not  g03636 ( new_n4013 , new_n4012 );
  xor  g03637 ( new_n4014 , new_n4010 , new_n4013 );
  nand g03638 ( new_n4015 , pi138 , pi218 );
  nand g03639 ( new_n4016 , pi182 , pi195 );
  xor  g03640 ( new_n4017 , new_n4015 , new_n4016 );
  xor  g03641 ( new_n4018 , new_n3916 , new_n4017 );
  nand g03642 ( new_n4019 , new_n3901 , new_n3907 );
  nand g03643 ( new_n4020 , new_n3908 , new_n3911 );
  nand g03644 ( new_n4021 , new_n4019 , new_n4020 );
  xor  g03645 ( new_n4022 , new_n4018 , new_n4021 );
  xor  g03646 ( new_n4023 , new_n4014 , new_n4022 );
  nor  g03647 ( new_n4024 , new_n3920 , new_n3923 );
  and  g03648 ( new_n4025 , new_n3917 , new_n4024 );
  or   g03649 ( new_n4026 , new_n3912 , new_n3919 );
  nand g03650 ( new_n4027 , new_n3918 , new_n4026 );
  nor  g03651 ( new_n4028 , new_n4024 , new_n4027 );
  or   g03652 ( new_n4029 , new_n4025 , new_n4028 );
  xor  g03653 ( new_n4030 , new_n4023 , new_n4029 );
  xor  g03654 ( new_n4031 , new_n4006 , new_n4030 );
  nor  g03655 ( new_n4032 , new_n3900 , new_n3929 );
  nor  g03656 ( new_n4033 , new_n3899 , new_n3931 );
  or   g03657 ( new_n4034 , new_n4032 , new_n4033 );
  xor  g03658 ( new_n4035 , new_n4031 , new_n4034 );
  nand g03659 ( new_n4036 , new_n3932 , new_n3935 );
  nand g03660 ( new_n4037 , new_n3898 , new_n3936 );
  nand g03661 ( new_n4038 , new_n4036 , new_n4037 );
  xor  g03662 ( new_n4039 , new_n4035 , new_n4038 );
  xor  g03663 ( new_n4040 , new_n4005 , new_n4039 );
  xor  g03664 ( new_n4041 , new_n3621 , new_n3940 );
  nand g03665 ( new_n4042 , new_n4040 , new_n4041 );
  nand g03666 ( new_n4043 , new_n3941 , new_n4042 );
  or   g03667 ( new_n4044 , new_n4035 , new_n4038 );
  not  g03668 ( new_n4045 , new_n4005 );
  nand g03669 ( new_n4046 , new_n4045 , new_n4039 );
  nand g03670 ( new_n4047 , new_n4044 , new_n4046 );
  nand g03671 ( new_n4048 , new_n3969 , new_n3998 );
  nand g03672 ( new_n4049 , new_n3999 , new_n4004 );
  nand g03673 ( new_n4050 , new_n4048 , new_n4049 );
  nor  g03674 ( new_n4051 , new_n4023 , new_n4029 );
  nor  g03675 ( new_n4052 , new_n4028 , new_n4051 );
  nand g03676 ( new_n4053 , pi037 , pi138 );
  xor  g03677 ( new_n4054 , new_n4052 , new_n4053 );
  xor  g03678 ( new_n4055 , new_n4050 , new_n4054 );
  nand g03679 ( new_n4056 , new_n3591 , new_n3594 );
  nand g03680 ( new_n4057 , new_n3587 , new_n3595 );
  nand g03681 ( new_n4058 , new_n4056 , new_n4057 );
  nand g03682 ( new_n4059 , new_n3588 , new_n3589 );
  nand g03683 ( new_n4060 , new_n3542 , new_n3590 );
  nand g03684 ( new_n4061 , new_n4059 , new_n4060 );
  xor  g03685 ( new_n4062 , new_n4058 , new_n4061 );
  nand g03686 ( new_n4063 , pi069 , pi177 );
  nand g03687 ( new_n4064 , pi101 , pi150 );
  nand g03688 ( new_n4065 , pi221 , pi223 );
  xor  g03689 ( new_n4066 , new_n4064 , new_n4065 );
  xor  g03690 ( new_n4067 , new_n4063 , new_n4066 );
  xor  g03691 ( new_n4068 , new_n4062 , new_n4067 );
  or   g03692 ( new_n4069 , new_n4006 , new_n4030 );
  nand g03693 ( new_n4070 , new_n4031 , new_n4034 );
  nand g03694 ( new_n4071 , new_n4069 , new_n4070 );
  nand g03695 ( new_n4072 , pi060 , pi196 );
  nand g03696 ( new_n4073 , pi225 , pi244 );
  xor  g03697 ( new_n4074 , new_n4072 , new_n4073 );
  xor  g03698 ( new_n4075 , new_n4071 , new_n4074 );
  xor  g03699 ( new_n4076 , new_n4068 , new_n4075 );
  nand g03700 ( new_n4077 , pi020 , pi184 );
  nand g03701 ( new_n4078 , new_n3581 , new_n3582 );
  nand g03702 ( new_n4079 , new_n3527 , new_n3583 );
  nand g03703 ( new_n4080 , new_n4078 , new_n4079 );
  xor  g03704 ( new_n4081 , new_n4077 , new_n4080 );
  nand g03705 ( new_n4082 , pi132 , pi192 );
  nand g03706 ( new_n4083 , pi186 , pi251 );
  xor  g03707 ( new_n4084 , new_n4082 , new_n4083 );
  xor  g03708 ( new_n4085 , new_n4081 , new_n4084 );
  xor  g03709 ( new_n4086 , new_n4076 , new_n4085 );
  xor  g03710 ( new_n4087 , new_n4055 , new_n4086 );
  nand g03711 ( new_n4088 , pi041 , pi195 );
  nand g03712 ( new_n4089 , pi076 , pi211 );
  or   g03713 ( new_n4090 , new_n4018 , new_n4021 );
  nand g03714 ( new_n4091 , new_n4014 , new_n4022 );
  nand g03715 ( new_n4092 , new_n4090 , new_n4091 );
  xor  g03716 ( new_n4093 , new_n4089 , new_n4092 );
  xor  g03717 ( new_n4094 , new_n4088 , new_n4093 );
  xor  g03718 ( new_n4095 , new_n4087 , new_n4094 );
  nand g03719 ( new_n4096 , new_n3853 , new_n3962 );
  nand g03720 ( new_n4097 , new_n3959 , new_n3963 );
  nand g03721 ( new_n4098 , new_n4096 , new_n4097 );
  nand g03722 ( new_n4099 , pi086 , pi226 );
  nand g03723 ( new_n4100 , new_n4015 , new_n4016 );
  nand g03724 ( new_n4101 , new_n3916 , new_n4017 );
  nand g03725 ( new_n4102 , new_n4100 , new_n4101 );
  nand g03726 ( new_n4103 , pi155 , pi207 );
  nand g03727 ( new_n4104 , pi023 , pi066 );
  xnor g03728 ( new_n4105 , new_n4103 , new_n4104 );
  xor  g03729 ( new_n4106 , new_n4102 , new_n4105 );
  xor  g03730 ( new_n4107 , new_n4099 , new_n4106 );
  xor  g03731 ( new_n4108 , new_n4098 , new_n4107 );
  nor  g03732 ( new_n4109 , new_n3906 , new_n4011 );
  nor  g03733 ( new_n4110 , new_n4010 , new_n4013 );
  or   g03734 ( new_n4111 , new_n4109 , new_n4110 );
  or   g03735 ( new_n4112 , new_n3943 , new_n3964 );
  nand g03736 ( new_n4113 , new_n3965 , new_n3968 );
  nand g03737 ( new_n4114 , new_n4112 , new_n4113 );
  nand g03738 ( new_n4115 , pi142 , pi243 );
  xor  g03739 ( new_n4116 , new_n4114 , new_n4115 );
  xor  g03740 ( new_n4117 , new_n4111 , new_n4116 );
  xor  g03741 ( new_n4118 , new_n4108 , new_n4117 );
  nand g03742 ( new_n4119 , pi182 , pi218 );
  nand g03743 ( new_n4120 , new_n3905 , new_n4008 );
  nand g03744 ( new_n4121 , new_n4007 , new_n4009 );
  nand g03745 ( new_n4122 , new_n4120 , new_n4121 );
  xor  g03746 ( new_n4123 , new_n4119 , new_n4122 );
  nand g03747 ( new_n4124 , pi058 , pi079 );
  nand g03748 ( new_n4125 , pi199 , pi216 );
  xor  g03749 ( new_n4126 , new_n4124 , new_n4125 );
  xor  g03750 ( new_n4127 , new_n4123 , new_n4126 );
  xor  g03751 ( new_n4128 , new_n4118 , new_n4127 );
  xor  g03752 ( new_n4129 , new_n4095 , new_n4128 );
  nand g03753 ( new_n4130 , new_n3881 , new_n3989 );
  nand g03754 ( new_n4131 , new_n3987 , new_n3992 );
  nand g03755 ( new_n4132 , new_n4130 , new_n4131 );
  nand g03756 ( new_n4133 , pi014 , pi059 );
  nand g03757 ( new_n4134 , pi135 , pi173 );
  xor  g03758 ( new_n4135 , new_n4133 , new_n4134 );
  xor  g03759 ( new_n4136 , new_n4132 , new_n4135 );
  xor  g03760 ( new_n4137 , new_n4129 , new_n4136 );
  xor  g03761 ( new_n4138 , new_n4047 , new_n4137 );
  xor  g03762 ( new_n4139 , new_n4043 , new_n4138 );
  nor  g03763 ( new_n4140 , new_n3580 , new_n3603 );
  nor  g03764 ( new_n4141 , new_n3604 , new_n3620 );
  nor  g03765 ( new_n4142 , new_n4140 , new_n4141 );
  or   g03766 ( new_n4143 , new_n3528 , new_n3585 );
  not  g03767 ( new_n4144 , new_n3584 );
  nand g03768 ( new_n4145 , new_n4144 , new_n3586 );
  nand g03769 ( new_n4146 , new_n4143 , new_n4145 );
  nand g03770 ( new_n4147 , pi122 , pi230 );
  nand g03771 ( new_n4148 , pi001 , pi050 );
  xor  g03772 ( new_n4149 , new_n4147 , new_n4148 );
  nand g03773 ( new_n4150 , new_n3838 , new_n3945 );
  nand g03774 ( new_n4151 , new_n3944 , new_n3946 );
  nand g03775 ( new_n4152 , new_n4150 , new_n4151 );
  nand g03776 ( new_n4153 , pi055 , pi099 );
  nand g03777 ( new_n4154 , pi002 , pi123 );
  xor  g03778 ( new_n4155 , new_n4153 , new_n4154 );
  xor  g03779 ( new_n4156 , new_n4152 , new_n4155 );
  nand g03780 ( new_n4157 , pi071 , pi239 );
  nand g03781 ( new_n4158 , pi025 , pi169 );
  xnor g03782 ( new_n4159 , new_n4157 , new_n4158 );
  or   g03783 ( new_n4160 , new_n3839 , new_n3948 );
  not  g03784 ( new_n4161 , new_n3947 );
  nand g03785 ( new_n4162 , new_n4161 , new_n3949 );
  nand g03786 ( new_n4163 , new_n4160 , new_n4162 );
  xor  g03787 ( new_n4164 , new_n4159 , new_n4163 );
  nand g03788 ( new_n4165 , new_n3951 , new_n3952 );
  nand g03789 ( new_n4166 , new_n3852 , new_n3953 );
  nand g03790 ( new_n4167 , new_n4165 , new_n4166 );
  nand g03791 ( new_n4168 , new_n3954 , new_n3957 );
  nand g03792 ( new_n4169 , new_n3950 , new_n3958 );
  nand g03793 ( new_n4170 , new_n4168 , new_n4169 );
  xor  g03794 ( new_n4171 , new_n4167 , new_n4170 );
  xor  g03795 ( new_n4172 , new_n4164 , new_n4171 );
  xor  g03796 ( new_n4173 , new_n4156 , new_n4172 );
  xor  g03797 ( new_n4174 , new_n4149 , new_n4173 );
  not  g03798 ( new_n4175 , new_n3993 );
  nor  g03799 ( new_n4176 , new_n3970 , new_n4175 );
  nor  g03800 ( new_n4177 , new_n3994 , new_n3997 );
  nor  g03801 ( new_n4178 , new_n4176 , new_n4177 );
  nand g03802 ( new_n4179 , pi087 , pi205 );
  xor  g03803 ( new_n4180 , new_n4178 , new_n4179 );
  xor  g03804 ( new_n4181 , new_n4174 , new_n4180 );
  nand g03805 ( new_n4182 , pi094 , pi109 );
  nand g03806 ( new_n4183 , pi029 , pi137 );
  nand g03807 ( new_n4184 , pi010 , pi160 );
  xor  g03808 ( new_n4185 , new_n4183 , new_n4184 );
  nand g03809 ( new_n4186 , new_n3979 , new_n3980 );
  nand g03810 ( new_n4187 , new_n3880 , new_n3981 );
  nand g03811 ( new_n4188 , new_n4186 , new_n4187 );
  nor  g03812 ( new_n4189 , new_n3874 , new_n3975 );
  nor  g03813 ( new_n4190 , new_n3974 , new_n3977 );
  or   g03814 ( new_n4191 , new_n4189 , new_n4190 );
  xor  g03815 ( new_n4192 , new_n4188 , new_n4191 );
  xor  g03816 ( new_n4193 , new_n4185 , new_n4192 );
  nor  g03817 ( new_n4194 , new_n3596 , new_n3602 );
  nor  g03818 ( new_n4195 , new_n3601 , new_n4194 );
  nand g03819 ( new_n4196 , new_n3971 , new_n3972 );
  nand g03820 ( new_n4197 , new_n3872 , new_n3973 );
  nand g03821 ( new_n4198 , new_n4196 , new_n4197 );
  nand g03822 ( new_n4199 , pi074 , pi219 );
  nand g03823 ( new_n4200 , pi102 , pi253 );
  xor  g03824 ( new_n4201 , new_n4199 , new_n4200 );
  or   g03825 ( new_n4202 , new_n3982 , new_n3985 );
  nand g03826 ( new_n4203 , new_n3978 , new_n3986 );
  nand g03827 ( new_n4204 , new_n4202 , new_n4203 );
  xor  g03828 ( new_n4205 , new_n4201 , new_n4204 );
  xor  g03829 ( new_n4206 , new_n4198 , new_n4205 );
  xor  g03830 ( new_n4207 , new_n4195 , new_n4206 );
  xor  g03831 ( new_n4208 , new_n4193 , new_n4207 );
  xor  g03832 ( new_n4209 , new_n4182 , new_n4208 );
  xor  g03833 ( new_n4210 , new_n4181 , new_n4209 );
  xor  g03834 ( new_n4211 , new_n4146 , new_n4210 );
  xor  g03835 ( new_n4212 , new_n4142 , new_n4211 );
  xor  g03836 ( po013 , new_n4139 , new_n4212 );
  nor  g03837 ( new_n4214 , new_n913 , new_n924 );
  nand g03838 ( new_n4215 , pi049 , pi108 );
  nand g03839 ( new_n4216 , pi042 , pi245 );
  nand g03840 ( new_n4217 , pi051 , pi201 );
  xor  g03841 ( new_n4218 , new_n4216 , new_n4217 );
  xor  g03842 ( new_n4219 , new_n4215 , new_n4218 );
  nand g03843 ( new_n4220 , pi007 , pi171 );
  nand g03844 ( new_n4221 , new_n920 , new_n921 );
  nand g03845 ( new_n4222 , new_n919 , new_n922 );
  nand g03846 ( new_n4223 , new_n4221 , new_n4222 );
  xor  g03847 ( new_n4224 , new_n4220 , new_n4223 );
  xor  g03848 ( new_n4225 , new_n4219 , new_n4224 );
  nand g03849 ( new_n4226 , pi107 , pi118 );
  or   g03850 ( new_n4227 , new_n914 , new_n917 );
  not  g03851 ( new_n4228 , new_n923 );
  nand g03852 ( new_n4229 , new_n918 , new_n4228 );
  nand g03853 ( new_n4230 , new_n4227 , new_n4229 );
  xor  g03854 ( new_n4231 , new_n4226 , new_n4230 );
  xor  g03855 ( new_n4232 , new_n4225 , new_n4231 );
  nand g03856 ( new_n4233 , new_n4214 , new_n4232 );
  nand g03857 ( new_n4234 , pi107 , pi113 );
  nand g03858 ( new_n4235 , new_n4233 , new_n4234 );
  nand g03859 ( new_n4236 , pi108 , pi245 );
  nand g03860 ( new_n4237 , pi042 , pi201 );
  nand g03861 ( new_n4238 , pi051 , pi156 );
  nand g03862 ( new_n4239 , new_n4237 , new_n4238 );
  nand g03863 ( new_n4240 , pi042 , pi156 );
  or   g03864 ( new_n4241 , new_n4217 , new_n4240 );
  nand g03865 ( new_n4242 , new_n4239 , new_n4241 );
  xor  g03866 ( new_n4243 , new_n4236 , new_n4242 );
  nand g03867 ( new_n4244 , new_n4216 , new_n4217 );
  nand g03868 ( new_n4245 , new_n4215 , new_n4218 );
  nand g03869 ( new_n4246 , new_n4244 , new_n4245 );
  xor  g03870 ( new_n4247 , new_n4243 , new_n4246 );
  nand g03871 ( new_n4248 , pi007 , pi049 );
  nand g03872 ( new_n4249 , pi118 , pi171 );
  and  g03873 ( new_n4250 , new_n4248 , new_n4249 );
  nand g03874 ( new_n4251 , pi049 , pi118 );
  nor  g03875 ( new_n4252 , new_n4220 , new_n4251 );
  or   g03876 ( new_n4253 , new_n4250 , new_n4252 );
  xnor g03877 ( new_n4254 , new_n4247 , new_n4253 );
  nand g03878 ( new_n4255 , new_n4220 , new_n4223 );
  nand g03879 ( new_n4256 , new_n4219 , new_n4224 );
  nand g03880 ( new_n4257 , new_n4255 , new_n4256 );
  xor  g03881 ( new_n4258 , new_n4254 , new_n4257 );
  not  g03882 ( new_n4259 , new_n4226 );
  nand g03883 ( new_n4260 , new_n4259 , new_n4230 );
  or   g03884 ( new_n4261 , new_n4225 , new_n4231 );
  nand g03885 ( new_n4262 , new_n4260 , new_n4261 );
  xnor g03886 ( new_n4263 , new_n4258 , new_n4262 );
  xor  g03887 ( new_n4264 , new_n4233 , new_n4234 );
  nand g03888 ( new_n4265 , new_n4263 , new_n4264 );
  nand g03889 ( new_n4266 , new_n4235 , new_n4265 );
  nand g03890 ( new_n4267 , new_n4258 , new_n4262 );
  nand g03891 ( new_n4268 , pi051 , pi063 );
  nand g03892 ( new_n4269 , pi108 , pi201 );
  xor  g03893 ( new_n4270 , new_n4268 , new_n4269 );
  xor  g03894 ( new_n4271 , new_n4240 , new_n4270 );
  not  g03895 ( new_n4272 , new_n4271 );
  nand g03896 ( new_n4273 , pi007 , pi245 );
  xor  g03897 ( new_n4274 , new_n4241 , new_n4273 );
  xor  g03898 ( new_n4275 , new_n4272 , new_n4274 );
  nand g03899 ( new_n4276 , pi038 , pi107 );
  nand g03900 ( new_n4277 , pi113 , pi171 );
  xor  g03901 ( new_n4278 , new_n4276 , new_n4277 );
  xor  g03902 ( new_n4279 , new_n4251 , new_n4278 );
  nand g03903 ( new_n4280 , new_n4236 , new_n4242 );
  nand g03904 ( new_n4281 , new_n4243 , new_n4246 );
  nand g03905 ( new_n4282 , new_n4280 , new_n4281 );
  xor  g03906 ( new_n4283 , new_n4279 , new_n4282 );
  xor  g03907 ( new_n4284 , new_n4275 , new_n4283 );
  nor  g03908 ( new_n4285 , new_n4247 , new_n4253 );
  nor  g03909 ( new_n4286 , new_n4254 , new_n4257 );
  xor  g03910 ( new_n4287 , new_n4252 , new_n4286 );
  nor  g03911 ( new_n4288 , new_n4285 , new_n4287 );
  xor  g03912 ( new_n4289 , new_n4284 , new_n4288 );
  xor  g03913 ( new_n4290 , new_n4267 , new_n4289 );
  xor  g03914 ( new_n4291 , new_n4266 , new_n4290 );
  nand g03915 ( new_n4292 , pi039 , pi061 );
  nand g03916 ( new_n4293 , pi116 , pi178 );
  nand g03917 ( new_n4294 , pi070 , pi188 );
  nand g03918 ( new_n4295 , new_n4293 , new_n4294 );
  nand g03919 ( new_n4296 , pi116 , pi188 );
  nand g03920 ( new_n4297 , pi070 , pi178 );
  or   g03921 ( new_n4298 , new_n4296 , new_n4297 );
  nand g03922 ( new_n4299 , new_n4295 , new_n4298 );
  xor  g03923 ( new_n4300 , new_n4292 , new_n4299 );
  nand g03924 ( new_n4301 , pi039 , pi178 );
  nand g03925 ( new_n4302 , new_n4296 , new_n4301 );
  nand g03926 ( new_n4303 , pi061 , pi228 );
  xor  g03927 ( new_n4304 , new_n4296 , new_n4301 );
  nand g03928 ( new_n4305 , new_n4303 , new_n4304 );
  nand g03929 ( new_n4306 , new_n4302 , new_n4305 );
  xor  g03930 ( new_n4307 , new_n4300 , new_n4306 );
  nand g03931 ( new_n4308 , pi012 , pi228 );
  nand g03932 ( new_n4309 , pi144 , pi148 );
  and  g03933 ( new_n4310 , new_n4308 , new_n4309 );
  nand g03934 ( new_n4311 , pi012 , pi148 );
  nand g03935 ( new_n4312 , pi144 , pi228 );
  nor  g03936 ( new_n4313 , new_n4311 , new_n4312 );
  or   g03937 ( new_n4314 , new_n4310 , new_n4313 );
  xnor g03938 ( new_n4315 , new_n4307 , new_n4314 );
  nand g03939 ( new_n4316 , new_n936 , new_n937 );
  nand g03940 ( new_n4317 , new_n935 , new_n938 );
  nand g03941 ( new_n4318 , new_n4316 , new_n4317 );
  nand g03942 ( new_n4319 , new_n4311 , new_n4318 );
  xor  g03943 ( new_n4320 , new_n4303 , new_n4304 );
  xor  g03944 ( new_n4321 , new_n4311 , new_n4318 );
  nand g03945 ( new_n4322 , new_n4320 , new_n4321 );
  nand g03946 ( new_n4323 , new_n4319 , new_n4322 );
  xor  g03947 ( new_n4324 , new_n4315 , new_n4323 );
  xor  g03948 ( new_n4325 , new_n4320 , new_n4321 );
  nand g03949 ( new_n4326 , pi144 , pi163 );
  nor  g03950 ( new_n4327 , new_n4325 , new_n4326 );
  xnor g03951 ( new_n4328 , new_n4325 , new_n4326 );
  nand g03952 ( new_n4329 , new_n940 , new_n943 );
  nand g03953 ( new_n4330 , new_n939 , new_n944 );
  nand g03954 ( new_n4331 , new_n4329 , new_n4330 );
  nor  g03955 ( new_n4332 , new_n4328 , new_n4331 );
  nor  g03956 ( new_n4333 , new_n4327 , new_n4332 );
  not  g03957 ( new_n4334 , new_n4333 );
  nand g03958 ( new_n4335 , new_n4324 , new_n4334 );
  nand g03959 ( new_n4336 , pi115 , pi188 );
  nand g03960 ( new_n4337 , pi061 , pi116 );
  xor  g03961 ( new_n4338 , new_n4336 , new_n4337 );
  xor  g03962 ( new_n4339 , new_n4297 , new_n4338 );
  nand g03963 ( new_n4340 , pi012 , pi039 );
  xor  g03964 ( new_n4341 , new_n4298 , new_n4340 );
  xor  g03965 ( new_n4342 , new_n4339 , new_n4341 );
  nand g03966 ( new_n4343 , pi098 , pi148 );
  nand g03967 ( new_n4344 , pi043 , pi163 );
  xor  g03968 ( new_n4345 , new_n4343 , new_n4344 );
  xor  g03969 ( new_n4346 , new_n4312 , new_n4345 );
  nand g03970 ( new_n4347 , new_n4292 , new_n4299 );
  nand g03971 ( new_n4348 , new_n4300 , new_n4306 );
  nand g03972 ( new_n4349 , new_n4347 , new_n4348 );
  xor  g03973 ( new_n4350 , new_n4346 , new_n4349 );
  xnor g03974 ( new_n4351 , new_n4342 , new_n4350 );
  nor  g03975 ( new_n4352 , new_n4307 , new_n4314 );
  nor  g03976 ( new_n4353 , new_n4315 , new_n4323 );
  xor  g03977 ( new_n4354 , new_n4313 , new_n4353 );
  nor  g03978 ( new_n4355 , new_n4352 , new_n4354 );
  not  g03979 ( new_n4356 , new_n4355 );
  xor  g03980 ( new_n4357 , new_n4351 , new_n4356 );
  xor  g03981 ( new_n4358 , new_n4335 , new_n4357 );
  nand g03982 ( new_n4359 , pi098 , pi163 );
  xor  g03983 ( new_n4360 , new_n4324 , new_n4333 );
  nand g03984 ( new_n4361 , new_n4359 , new_n4360 );
  nor  g03985 ( new_n4362 , new_n934 , new_n945 );
  xor  g03986 ( new_n4363 , new_n4328 , new_n4331 );
  nand g03987 ( new_n4364 , new_n4362 , new_n4363 );
  xor  g03988 ( new_n4365 , new_n4359 , new_n4360 );
  nand g03989 ( new_n4366 , new_n4364 , new_n4365 );
  nand g03990 ( new_n4367 , new_n4361 , new_n4366 );
  xor  g03991 ( new_n4368 , new_n4358 , new_n4367 );
  not  g03992 ( new_n4369 , new_n4368 );
  xor  g03993 ( new_n4370 , new_n4291 , new_n4369 );
  xor  g03994 ( new_n4371 , new_n4263 , new_n4264 );
  xor  g03995 ( new_n4372 , new_n4364 , new_n4365 );
  nor  g03996 ( new_n4373 , new_n4371 , new_n4372 );
  xnor g03997 ( new_n4374 , new_n4371 , new_n4372 );
  xor  g03998 ( new_n4375 , new_n4214 , new_n4232 );
  nand g03999 ( new_n4376 , new_n925 , new_n946 );
  nand g04000 ( new_n4377 , new_n947 , new_n969 );
  nand g04001 ( new_n4378 , new_n4376 , new_n4377 );
  or   g04002 ( new_n4379 , new_n4375 , new_n4378 );
  xnor g04003 ( new_n4380 , new_n4362 , new_n4363 );
  xor  g04004 ( new_n4381 , new_n4375 , new_n4378 );
  nand g04005 ( new_n4382 , new_n4380 , new_n4381 );
  nand g04006 ( new_n4383 , new_n4379 , new_n4382 );
  nor  g04007 ( new_n4384 , new_n4374 , new_n4383 );
  nor  g04008 ( new_n4385 , new_n4373 , new_n4384 );
  xnor g04009 ( new_n4386 , new_n4370 , new_n4385 );
  nand g04010 ( new_n4387 , pi149 , pi179 );
  nand g04011 ( new_n4388 , pi179 , pi240 );
  nand g04012 ( new_n4389 , pi033 , pi149 );
  nand g04013 ( new_n4390 , new_n4388 , new_n4389 );
  nand g04014 ( new_n4391 , pi162 , pi167 );
  xor  g04015 ( new_n4392 , new_n4388 , new_n4389 );
  nand g04016 ( new_n4393 , new_n4391 , new_n4392 );
  nand g04017 ( new_n4394 , new_n4390 , new_n4393 );
  xnor g04018 ( new_n4395 , new_n4387 , new_n4394 );
  nand g04019 ( new_n4396 , pi033 , pi167 );
  nand g04020 ( new_n4397 , pi162 , pi181 );
  nand g04021 ( new_n4398 , new_n4396 , new_n4397 );
  nand g04022 ( new_n4399 , pi033 , pi181 );
  or   g04023 ( new_n4400 , new_n4391 , new_n4399 );
  nand g04024 ( new_n4401 , new_n4398 , new_n4400 );
  xnor g04025 ( new_n4402 , new_n4395 , new_n4401 );
  nand g04026 ( new_n4403 , pi048 , pi240 );
  nand g04027 ( new_n4404 , pi134 , pi237 );
  and  g04028 ( new_n4405 , new_n4403 , new_n4404 );
  nand g04029 ( new_n4406 , pi048 , pi134 );
  nand g04030 ( new_n4407 , pi237 , pi240 );
  nor  g04031 ( new_n4408 , new_n4406 , new_n4407 );
  or   g04032 ( new_n4409 , new_n4405 , new_n4408 );
  xnor g04033 ( new_n4410 , new_n4402 , new_n4409 );
  nand g04034 ( new_n4411 , new_n981 , new_n982 );
  nand g04035 ( new_n4412 , new_n980 , new_n983 );
  nand g04036 ( new_n4413 , new_n4411 , new_n4412 );
  nand g04037 ( new_n4414 , new_n4406 , new_n4413 );
  xor  g04038 ( new_n4415 , new_n4391 , new_n4392 );
  xor  g04039 ( new_n4416 , new_n4406 , new_n4413 );
  nand g04040 ( new_n4417 , new_n4415 , new_n4416 );
  nand g04041 ( new_n4418 , new_n4414 , new_n4417 );
  xor  g04042 ( new_n4419 , new_n4410 , new_n4418 );
  nand g04043 ( new_n4420 , pi175 , pi237 );
  not  g04044 ( new_n4421 , new_n4420 );
  or   g04045 ( new_n4422 , new_n977 , new_n978 );
  nand g04046 ( new_n4423 , new_n979 , new_n984 );
  nand g04047 ( new_n4424 , new_n4422 , new_n4423 );
  nand g04048 ( new_n4425 , new_n4421 , new_n4424 );
  xor  g04049 ( new_n4426 , new_n4420 , new_n4424 );
  xor  g04050 ( new_n4427 , new_n4415 , new_n4416 );
  or   g04051 ( new_n4428 , new_n4426 , new_n4427 );
  nand g04052 ( new_n4429 , new_n4425 , new_n4428 );
  nand g04053 ( new_n4430 , new_n4419 , new_n4429 );
  nand g04054 ( new_n4431 , pi162 , pi200 );
  nand g04055 ( new_n4432 , pi167 , pi179 );
  xor  g04056 ( new_n4433 , new_n4431 , new_n4432 );
  xor  g04057 ( new_n4434 , new_n4399 , new_n4433 );
  nand g04058 ( new_n4435 , pi048 , pi149 );
  xor  g04059 ( new_n4436 , new_n4400 , new_n4435 );
  xor  g04060 ( new_n4437 , new_n4434 , new_n4436 );
  nand g04061 ( new_n4438 , pi134 , pi238 );
  nand g04062 ( new_n4439 , pi175 , pi193 );
  xor  g04063 ( new_n4440 , new_n4438 , new_n4439 );
  xor  g04064 ( new_n4441 , new_n4407 , new_n4440 );
  nor  g04065 ( new_n4442 , new_n4387 , new_n4394 );
  nor  g04066 ( new_n4443 , new_n4395 , new_n4401 );
  nor  g04067 ( new_n4444 , new_n4442 , new_n4443 );
  xor  g04068 ( new_n4445 , new_n4441 , new_n4444 );
  xnor g04069 ( new_n4446 , new_n4437 , new_n4445 );
  nor  g04070 ( new_n4447 , new_n4402 , new_n4409 );
  nor  g04071 ( new_n4448 , new_n4410 , new_n4418 );
  xor  g04072 ( new_n4449 , new_n4408 , new_n4448 );
  nor  g04073 ( new_n4450 , new_n4447 , new_n4449 );
  not  g04074 ( new_n4451 , new_n4450 );
  xor  g04075 ( new_n4452 , new_n4446 , new_n4451 );
  xor  g04076 ( new_n4453 , new_n4430 , new_n4452 );
  nand g04077 ( new_n4454 , pi175 , pi238 );
  nor  g04078 ( new_n4455 , new_n985 , new_n992 );
  xor  g04079 ( new_n4456 , new_n4426 , new_n4427 );
  nand g04080 ( new_n4457 , new_n4455 , new_n4456 );
  nand g04081 ( new_n4458 , new_n4454 , new_n4457 );
  xor  g04082 ( new_n4459 , new_n4419 , new_n4429 );
  not  g04083 ( new_n4460 , new_n4459 );
  xor  g04084 ( new_n4461 , new_n4454 , new_n4457 );
  nand g04085 ( new_n4462 , new_n4460 , new_n4461 );
  nand g04086 ( new_n4463 , new_n4458 , new_n4462 );
  xor  g04087 ( new_n4464 , new_n4453 , new_n4463 );
  xor  g04088 ( new_n4465 , new_n4386 , new_n4464 );
  xor  g04089 ( new_n4466 , new_n4459 , new_n4461 );
  xnor g04090 ( new_n4467 , new_n4455 , new_n4456 );
  or   g04091 ( new_n4468 , new_n993 , new_n1011 );
  not  g04092 ( new_n4469 , new_n970 );
  nand g04093 ( new_n4470 , new_n4469 , new_n1012 );
  nand g04094 ( new_n4471 , new_n4468 , new_n4470 );
  or   g04095 ( new_n4472 , new_n4467 , new_n4471 );
  xnor g04096 ( new_n4473 , new_n4380 , new_n4381 );
  xor  g04097 ( new_n4474 , new_n4467 , new_n4471 );
  nand g04098 ( new_n4475 , new_n4473 , new_n4474 );
  nand g04099 ( new_n4476 , new_n4472 , new_n4475 );
  nand g04100 ( new_n4477 , new_n4466 , new_n4476 );
  xor  g04101 ( new_n4478 , new_n4374 , new_n4383 );
  xor  g04102 ( new_n4479 , new_n4466 , new_n4476 );
  nand g04103 ( new_n4480 , new_n4478 , new_n4479 );
  nand g04104 ( new_n4481 , new_n4477 , new_n4480 );
  xor  g04105 ( new_n4482 , new_n4465 , new_n4481 );
  nand g04106 ( new_n4483 , pi080 , pi194 );
  nand g04107 ( new_n4484 , pi143 , pi247 );
  nand g04108 ( new_n4485 , pi057 , pi080 );
  nand g04109 ( new_n4486 , new_n4484 , new_n4485 );
  nand g04110 ( new_n4487 , pi016 , pi194 );
  xor  g04111 ( new_n4488 , new_n4484 , new_n4485 );
  nand g04112 ( new_n4489 , new_n4487 , new_n4488 );
  nand g04113 ( new_n4490 , new_n4486 , new_n4489 );
  xnor g04114 ( new_n4491 , new_n4483 , new_n4490 );
  nand g04115 ( new_n4492 , pi057 , pi247 );
  nand g04116 ( new_n4493 , pi143 , pi234 );
  nand g04117 ( new_n4494 , new_n4492 , new_n4493 );
  nand g04118 ( new_n4495 , pi057 , pi234 );
  or   g04119 ( new_n4496 , new_n4484 , new_n4495 );
  nand g04120 ( new_n4497 , new_n4494 , new_n4496 );
  xnor g04121 ( new_n4498 , new_n4491 , new_n4497 );
  nand g04122 ( new_n4499 , pi016 , pi085 );
  nand g04123 ( new_n4500 , pi117 , pi180 );
  and  g04124 ( new_n4501 , new_n4499 , new_n4500 );
  nand g04125 ( new_n4502 , pi085 , pi117 );
  nand g04126 ( new_n4503 , pi016 , pi180 );
  nor  g04127 ( new_n4504 , new_n4502 , new_n4503 );
  or   g04128 ( new_n4505 , new_n4501 , new_n4504 );
  xnor g04129 ( new_n4506 , new_n4498 , new_n4505 );
  nand g04130 ( new_n4507 , new_n1024 , new_n1025 );
  nand g04131 ( new_n4508 , new_n1023 , new_n1026 );
  nand g04132 ( new_n4509 , new_n4507 , new_n4508 );
  nand g04133 ( new_n4510 , new_n4502 , new_n4509 );
  xor  g04134 ( new_n4511 , new_n4487 , new_n4488 );
  xor  g04135 ( new_n4512 , new_n4502 , new_n4509 );
  nand g04136 ( new_n4513 , new_n4511 , new_n4512 );
  nand g04137 ( new_n4514 , new_n4510 , new_n4513 );
  xor  g04138 ( new_n4515 , new_n4506 , new_n4514 );
  nand g04139 ( new_n4516 , pi103 , pi180 );
  nand g04140 ( new_n4517 , new_n1028 , new_n1031 );
  nand g04141 ( new_n4518 , new_n1027 , new_n1032 );
  nand g04142 ( new_n4519 , new_n4517 , new_n4518 );
  or   g04143 ( new_n4520 , new_n4516 , new_n4519 );
  xnor g04144 ( new_n4521 , new_n4511 , new_n4512 );
  xor  g04145 ( new_n4522 , new_n4516 , new_n4519 );
  nand g04146 ( new_n4523 , new_n4521 , new_n4522 );
  nand g04147 ( new_n4524 , new_n4520 , new_n4523 );
  nand g04148 ( new_n4525 , new_n4515 , new_n4524 );
  nand g04149 ( new_n4526 , pi143 , pi214 );
  nand g04150 ( new_n4527 , pi194 , pi247 );
  xor  g04151 ( new_n4528 , new_n4526 , new_n4527 );
  xor  g04152 ( new_n4529 , new_n4495 , new_n4528 );
  nand g04153 ( new_n4530 , pi080 , pi085 );
  xor  g04154 ( new_n4531 , new_n4496 , new_n4530 );
  xor  g04155 ( new_n4532 , new_n4529 , new_n4531 );
  nand g04156 ( new_n4533 , pi036 , pi117 );
  nand g04157 ( new_n4534 , pi068 , pi103 );
  xor  g04158 ( new_n4535 , new_n4533 , new_n4534 );
  xor  g04159 ( new_n4536 , new_n4503 , new_n4535 );
  nor  g04160 ( new_n4537 , new_n4483 , new_n4490 );
  nor  g04161 ( new_n4538 , new_n4491 , new_n4497 );
  nor  g04162 ( new_n4539 , new_n4537 , new_n4538 );
  xor  g04163 ( new_n4540 , new_n4536 , new_n4539 );
  xnor g04164 ( new_n4541 , new_n4532 , new_n4540 );
  nor  g04165 ( new_n4542 , new_n4498 , new_n4505 );
  nor  g04166 ( new_n4543 , new_n4506 , new_n4514 );
  xor  g04167 ( new_n4544 , new_n4504 , new_n4543 );
  nor  g04168 ( new_n4545 , new_n4542 , new_n4544 );
  xor  g04169 ( new_n4546 , new_n4541 , new_n4545 );
  xor  g04170 ( new_n4547 , new_n4525 , new_n4546 );
  nand g04171 ( new_n4548 , pi036 , pi103 );
  nor  g04172 ( new_n4549 , new_n1022 , new_n1033 );
  xor  g04173 ( new_n4550 , new_n4521 , new_n4522 );
  nand g04174 ( new_n4551 , new_n4549 , new_n4550 );
  nand g04175 ( new_n4552 , new_n4548 , new_n4551 );
  xnor g04176 ( new_n4553 , new_n4515 , new_n4524 );
  xor  g04177 ( new_n4554 , new_n4548 , new_n4551 );
  nand g04178 ( new_n4555 , new_n4553 , new_n4554 );
  nand g04179 ( new_n4556 , new_n4552 , new_n4555 );
  xor  g04180 ( new_n4557 , new_n4547 , new_n4556 );
  xor  g04181 ( new_n4558 , new_n4553 , new_n4554 );
  xor  g04182 ( new_n4559 , new_n4549 , new_n4550 );
  nand g04183 ( new_n4560 , new_n1034 , new_n1052 );
  nand g04184 ( new_n4561 , new_n1013 , new_n1053 );
  nand g04185 ( new_n4562 , new_n4560 , new_n4561 );
  or   g04186 ( new_n4563 , new_n4559 , new_n4562 );
  xor  g04187 ( new_n4564 , new_n4473 , new_n4474 );
  not  g04188 ( new_n4565 , new_n4564 );
  xor  g04189 ( new_n4566 , new_n4559 , new_n4562 );
  nand g04190 ( new_n4567 , new_n4565 , new_n4566 );
  nand g04191 ( new_n4568 , new_n4563 , new_n4567 );
  nand g04192 ( new_n4569 , new_n4558 , new_n4568 );
  xor  g04193 ( new_n4570 , new_n4478 , new_n4479 );
  not  g04194 ( new_n4571 , new_n4570 );
  xor  g04195 ( new_n4572 , new_n4558 , new_n4568 );
  nand g04196 ( new_n4573 , new_n4571 , new_n4572 );
  nand g04197 ( new_n4574 , new_n4569 , new_n4573 );
  xor  g04198 ( new_n4575 , new_n4557 , new_n4574 );
  xor  g04199 ( po014 , new_n4482 , new_n4575 );
  nand g04200 ( new_n4577 , pi042 , pi241 );
  nand g04201 ( new_n4578 , pi108 , pi236 );
  xor  g04202 ( new_n4579 , new_n4577 , new_n4578 );
  nand g04203 ( new_n4580 , pi051 , pi161 );
  xor  g04204 ( new_n4581 , new_n4579 , new_n4580 );
  nor  g04205 ( new_n4582 , new_n3513 , new_n4577 );
  not  g04206 ( new_n4583 , new_n4582 );
  or   g04207 ( new_n4584 , new_n4581 , new_n4583 );
  nand g04208 ( new_n4585 , pi007 , pi236 );
  nand g04209 ( new_n4586 , new_n4577 , new_n4578 );
  nand g04210 ( new_n4587 , new_n4579 , new_n4580 );
  nand g04211 ( new_n4588 , new_n4586 , new_n4587 );
  xor  g04212 ( new_n4589 , new_n4585 , new_n4588 );
  nand g04213 ( new_n4590 , pi051 , pi141 );
  nand g04214 ( new_n4591 , pi108 , pi241 );
  nand g04215 ( new_n4592 , pi042 , pi161 );
  xor  g04216 ( new_n4593 , new_n4591 , new_n4592 );
  xor  g04217 ( new_n4594 , new_n4590 , new_n4593 );
  xor  g04218 ( new_n4595 , new_n4589 , new_n4594 );
  nor  g04219 ( new_n4596 , new_n4584 , new_n4595 );
  nand g04220 ( new_n4597 , pi108 , pi161 );
  nand g04221 ( new_n4598 , pi051 , pi090 );
  nand g04222 ( new_n4599 , pi042 , pi141 );
  xor  g04223 ( new_n4600 , new_n4598 , new_n4599 );
  xor  g04224 ( new_n4601 , new_n4597 , new_n4600 );
  nand g04225 ( new_n4602 , pi007 , pi241 );
  nand g04226 ( new_n4603 , new_n4591 , new_n4592 );
  nand g04227 ( new_n4604 , new_n4590 , new_n4593 );
  nand g04228 ( new_n4605 , new_n4603 , new_n4604 );
  xor  g04229 ( new_n4606 , new_n4602 , new_n4605 );
  xor  g04230 ( new_n4607 , new_n4601 , new_n4606 );
  nand g04231 ( new_n4608 , pi118 , pi236 );
  or   g04232 ( new_n4609 , new_n4585 , new_n4588 );
  not  g04233 ( new_n4610 , new_n4594 );
  nand g04234 ( new_n4611 , new_n4589 , new_n4610 );
  nand g04235 ( new_n4612 , new_n4609 , new_n4611 );
  xor  g04236 ( new_n4613 , new_n4608 , new_n4612 );
  xor  g04237 ( new_n4614 , new_n4607 , new_n4613 );
  xor  g04238 ( new_n4615 , new_n4596 , new_n4614 );
  nand g04239 ( new_n4616 , pi178 , pi212 );
  nand g04240 ( new_n4617 , pi061 , pi213 );
  xor  g04241 ( new_n4618 , new_n4616 , new_n4617 );
  nand g04242 ( new_n4619 , pi104 , pi188 );
  xor  g04243 ( new_n4620 , new_n4618 , new_n4619 );
  nor  g04244 ( new_n4621 , new_n3514 , new_n4616 );
  not  g04245 ( new_n4622 , new_n4621 );
  or   g04246 ( new_n4623 , new_n4620 , new_n4622 );
  nand g04247 ( new_n4624 , pi013 , pi188 );
  nand g04248 ( new_n4625 , pi061 , pi212 );
  nand g04249 ( new_n4626 , pi104 , pi178 );
  xor  g04250 ( new_n4627 , new_n4625 , new_n4626 );
  xor  g04251 ( new_n4628 , new_n4624 , new_n4627 );
  nand g04252 ( new_n4629 , pi012 , pi213 );
  nand g04253 ( new_n4630 , new_n4616 , new_n4617 );
  nand g04254 ( new_n4631 , new_n4618 , new_n4619 );
  nand g04255 ( new_n4632 , new_n4630 , new_n4631 );
  xor  g04256 ( new_n4633 , new_n4629 , new_n4632 );
  xor  g04257 ( new_n4634 , new_n4628 , new_n4633 );
  or   g04258 ( new_n4635 , new_n4623 , new_n4634 );
  nand g04259 ( new_n4636 , pi112 , pi188 );
  nand g04260 ( new_n4637 , pi061 , pi104 );
  nand g04261 ( new_n4638 , pi013 , pi178 );
  xor  g04262 ( new_n4639 , new_n4637 , new_n4638 );
  xor  g04263 ( new_n4640 , new_n4636 , new_n4639 );
  nand g04264 ( new_n4641 , pi012 , pi212 );
  nand g04265 ( new_n4642 , new_n4625 , new_n4626 );
  nand g04266 ( new_n4643 , new_n4624 , new_n4627 );
  nand g04267 ( new_n4644 , new_n4642 , new_n4643 );
  xor  g04268 ( new_n4645 , new_n4641 , new_n4644 );
  xnor g04269 ( new_n4646 , new_n4640 , new_n4645 );
  nand g04270 ( new_n4647 , pi144 , pi213 );
  nand g04271 ( new_n4648 , new_n4629 , new_n4632 );
  nand g04272 ( new_n4649 , new_n4628 , new_n4633 );
  nand g04273 ( new_n4650 , new_n4648 , new_n4649 );
  xor  g04274 ( new_n4651 , new_n4647 , new_n4650 );
  xnor g04275 ( new_n4652 , new_n4646 , new_n4651 );
  xor  g04276 ( new_n4653 , new_n4635 , new_n4652 );
  xor  g04277 ( new_n4654 , new_n4615 , new_n4653 );
  xor  g04278 ( new_n4655 , new_n4584 , new_n4595 );
  xor  g04279 ( new_n4656 , new_n4623 , new_n4634 );
  nand g04280 ( new_n4657 , new_n4655 , new_n4656 );
  not  g04281 ( new_n4658 , new_n4657 );
  xnor g04282 ( new_n4659 , new_n4655 , new_n4656 );
  xor  g04283 ( new_n4660 , new_n4620 , new_n4621 );
  nor  g04284 ( new_n4661 , new_n3513 , new_n3514 );
  not  g04285 ( new_n4662 , new_n4661 );
  nand g04286 ( new_n4663 , pi042 , pi236 );
  nand g04287 ( new_n4664 , pi051 , pi241 );
  nand g04288 ( new_n4665 , new_n4663 , new_n4664 );
  nand g04289 ( new_n4666 , new_n4583 , new_n4665 );
  nor  g04290 ( new_n4667 , new_n4662 , new_n4666 );
  xor  g04291 ( new_n4668 , new_n4661 , new_n4666 );
  nand g04292 ( new_n4669 , pi178 , pi213 );
  nand g04293 ( new_n4670 , pi188 , pi212 );
  nand g04294 ( new_n4671 , new_n4669 , new_n4670 );
  nand g04295 ( new_n4672 , new_n4622 , new_n4671 );
  nor  g04296 ( new_n4673 , new_n4668 , new_n4672 );
  nor  g04297 ( new_n4674 , new_n4667 , new_n4673 );
  nand g04298 ( new_n4675 , new_n4660 , new_n4674 );
  xor  g04299 ( new_n4676 , new_n4581 , new_n4582 );
  xor  g04300 ( new_n4677 , new_n4660 , new_n4674 );
  nand g04301 ( new_n4678 , new_n4676 , new_n4677 );
  nand g04302 ( new_n4679 , new_n4675 , new_n4678 );
  nor  g04303 ( new_n4680 , new_n4659 , new_n4679 );
  nor  g04304 ( new_n4681 , new_n4658 , new_n4680 );
  xor  g04305 ( new_n4682 , new_n4654 , new_n4681 );
  nand g04306 ( new_n4683 , pi033 , pi208 );
  nand g04307 ( new_n4684 , pi168 , pi179 );
  xor  g04308 ( new_n4685 , new_n4683 , new_n4684 );
  nand g04309 ( new_n4686 , pi139 , pi162 );
  xor  g04310 ( new_n4687 , new_n4685 , new_n4686 );
  nor  g04311 ( new_n4688 , new_n3516 , new_n4683 );
  not  g04312 ( new_n4689 , new_n4688 );
  or   g04313 ( new_n4690 , new_n4687 , new_n4689 );
  nand g04314 ( new_n4691 , pi048 , pi168 );
  nand g04315 ( new_n4692 , new_n4683 , new_n4684 );
  nand g04316 ( new_n4693 , new_n4685 , new_n4686 );
  nand g04317 ( new_n4694 , new_n4692 , new_n4693 );
  xor  g04318 ( new_n4695 , new_n4691 , new_n4694 );
  nand g04319 ( new_n4696 , pi179 , pi208 );
  nand g04320 ( new_n4697 , pi035 , pi162 );
  nand g04321 ( new_n4698 , pi033 , pi139 );
  xor  g04322 ( new_n4699 , new_n4697 , new_n4698 );
  xnor g04323 ( new_n4700 , new_n4696 , new_n4699 );
  xnor g04324 ( new_n4701 , new_n4695 , new_n4700 );
  nor  g04325 ( new_n4702 , new_n4690 , new_n4701 );
  nand g04326 ( new_n4703 , pi139 , pi179 );
  nand g04327 ( new_n4704 , pi033 , pi035 );
  nand g04328 ( new_n4705 , pi015 , pi162 );
  xor  g04329 ( new_n4706 , new_n4704 , new_n4705 );
  xor  g04330 ( new_n4707 , new_n4703 , new_n4706 );
  nand g04331 ( new_n4708 , pi048 , pi208 );
  nand g04332 ( new_n4709 , new_n4697 , new_n4698 );
  nand g04333 ( new_n4710 , new_n4696 , new_n4699 );
  nand g04334 ( new_n4711 , new_n4709 , new_n4710 );
  xor  g04335 ( new_n4712 , new_n4708 , new_n4711 );
  xor  g04336 ( new_n4713 , new_n4707 , new_n4712 );
  nand g04337 ( new_n4714 , pi168 , pi237 );
  or   g04338 ( new_n4715 , new_n4691 , new_n4694 );
  nand g04339 ( new_n4716 , new_n4695 , new_n4700 );
  nand g04340 ( new_n4717 , new_n4715 , new_n4716 );
  xor  g04341 ( new_n4718 , new_n4714 , new_n4717 );
  xor  g04342 ( new_n4719 , new_n4713 , new_n4718 );
  xor  g04343 ( new_n4720 , new_n4702 , new_n4719 );
  xor  g04344 ( new_n4721 , new_n4659 , new_n4679 );
  xor  g04345 ( new_n4722 , new_n4690 , new_n4701 );
  nor  g04346 ( new_n4723 , new_n4721 , new_n4722 );
  xnor g04347 ( new_n4724 , new_n4721 , new_n4722 );
  xor  g04348 ( new_n4725 , new_n4687 , new_n4688 );
  not  g04349 ( new_n4726 , new_n3515 );
  or   g04350 ( new_n4727 , new_n4726 , new_n3516 );
  nand g04351 ( new_n4728 , pi033 , pi168 );
  nand g04352 ( new_n4729 , pi162 , pi208 );
  nand g04353 ( new_n4730 , new_n4728 , new_n4729 );
  nand g04354 ( new_n4731 , new_n4689 , new_n4730 );
  nand g04355 ( new_n4732 , new_n4727 , new_n4731 );
  xor  g04356 ( new_n4733 , new_n4668 , new_n4672 );
  not  g04357 ( new_n4734 , new_n4733 );
  xor  g04358 ( new_n4735 , new_n4727 , new_n4731 );
  nand g04359 ( new_n4736 , new_n4734 , new_n4735 );
  nand g04360 ( new_n4737 , new_n4732 , new_n4736 );
  or   g04361 ( new_n4738 , new_n4725 , new_n4737 );
  xor  g04362 ( new_n4739 , new_n4676 , new_n4677 );
  not  g04363 ( new_n4740 , new_n4739 );
  xor  g04364 ( new_n4741 , new_n4725 , new_n4737 );
  nand g04365 ( new_n4742 , new_n4740 , new_n4741 );
  nand g04366 ( new_n4743 , new_n4738 , new_n4742 );
  nor  g04367 ( new_n4744 , new_n4724 , new_n4743 );
  nor  g04368 ( new_n4745 , new_n4723 , new_n4744 );
  xor  g04369 ( new_n4746 , new_n4720 , new_n4745 );
  xor  g04370 ( new_n4747 , new_n4682 , new_n4746 );
  nand g04371 ( new_n4748 , pi052 , pi057 );
  nand g04372 ( new_n4749 , pi131 , pi194 );
  xor  g04373 ( new_n4750 , new_n4748 , new_n4749 );
  nand g04374 ( new_n4751 , pi077 , pi143 );
  xor  g04375 ( new_n4752 , new_n4750 , new_n4751 );
  nand g04376 ( new_n4753 , pi057 , pi131 );
  nand g04377 ( new_n4754 , pi052 , pi143 );
  nor  g04378 ( new_n4755 , new_n4753 , new_n4754 );
  not  g04379 ( new_n4756 , new_n4755 );
  nor  g04380 ( new_n4757 , new_n4752 , new_n4756 );
  not  g04381 ( new_n4758 , new_n4757 );
  nand g04382 ( new_n4759 , pi085 , pi131 );
  nand g04383 ( new_n4760 , new_n4748 , new_n4749 );
  nand g04384 ( new_n4761 , new_n4750 , new_n4751 );
  nand g04385 ( new_n4762 , new_n4760 , new_n4761 );
  xor  g04386 ( new_n4763 , new_n4759 , new_n4762 );
  nand g04387 ( new_n4764 , pi057 , pi077 );
  nand g04388 ( new_n4765 , pi052 , pi194 );
  nand g04389 ( new_n4766 , pi133 , pi143 );
  xor  g04390 ( new_n4767 , new_n4765 , new_n4766 );
  xnor g04391 ( new_n4768 , new_n4764 , new_n4767 );
  xnor g04392 ( new_n4769 , new_n4763 , new_n4768 );
  nor  g04393 ( new_n4770 , new_n4758 , new_n4769 );
  nand g04394 ( new_n4771 , pi057 , pi133 );
  nand g04395 ( new_n4772 , pi143 , pi189 );
  nand g04396 ( new_n4773 , pi077 , pi194 );
  xor  g04397 ( new_n4774 , new_n4772 , new_n4773 );
  xor  g04398 ( new_n4775 , new_n4771 , new_n4774 );
  nand g04399 ( new_n4776 , pi052 , pi085 );
  nand g04400 ( new_n4777 , new_n4765 , new_n4766 );
  nand g04401 ( new_n4778 , new_n4764 , new_n4767 );
  nand g04402 ( new_n4779 , new_n4777 , new_n4778 );
  xor  g04403 ( new_n4780 , new_n4776 , new_n4779 );
  xor  g04404 ( new_n4781 , new_n4775 , new_n4780 );
  nand g04405 ( new_n4782 , pi131 , pi180 );
  xor  g04406 ( new_n4783 , new_n4781 , new_n4782 );
  or   g04407 ( new_n4784 , new_n4759 , new_n4762 );
  nand g04408 ( new_n4785 , new_n4763 , new_n4768 );
  nand g04409 ( new_n4786 , new_n4784 , new_n4785 );
  xor  g04410 ( new_n4787 , new_n4783 , new_n4786 );
  xor  g04411 ( new_n4788 , new_n4770 , new_n4787 );
  xor  g04412 ( new_n4789 , new_n4747 , new_n4788 );
  xor  g04413 ( new_n4790 , new_n4724 , new_n4743 );
  xor  g04414 ( new_n4791 , new_n4758 , new_n4769 );
  not  g04415 ( new_n4792 , new_n4791 );
  nand g04416 ( new_n4793 , new_n4790 , new_n4792 );
  xor  g04417 ( new_n4794 , new_n4790 , new_n4792 );
  xor  g04418 ( new_n4795 , new_n4739 , new_n4741 );
  xor  g04419 ( new_n4796 , new_n4752 , new_n4756 );
  not  g04420 ( new_n4797 , new_n4796 );
  nor  g04421 ( new_n4798 , new_n4795 , new_n4797 );
  xor  g04422 ( new_n4799 , new_n4795 , new_n4796 );
  nor  g04423 ( new_n4800 , new_n3517 , new_n3518 );
  xor  g04424 ( new_n4801 , new_n4753 , new_n4754 );
  or   g04425 ( new_n4802 , new_n4800 , new_n4801 );
  xor  g04426 ( new_n4803 , new_n4734 , new_n4735 );
  xor  g04427 ( new_n4804 , new_n4800 , new_n4801 );
  nand g04428 ( new_n4805 , new_n4803 , new_n4804 );
  nand g04429 ( new_n4806 , new_n4802 , new_n4805 );
  nor  g04430 ( new_n4807 , new_n4799 , new_n4806 );
  nor  g04431 ( new_n4808 , new_n4798 , new_n4807 );
  nand g04432 ( new_n4809 , new_n4794 , new_n4808 );
  nand g04433 ( new_n4810 , new_n4793 , new_n4809 );
  xor  g04434 ( po015 , new_n4789 , new_n4810 );
  nand g04435 ( new_n4812 , pi007 , pi087 );
  nand g04436 ( new_n4813 , pi087 , pi108 );
  nand g04437 ( new_n4814 , pi051 , pi102 );
  nand g04438 ( new_n4815 , new_n4813 , new_n4814 );
  nand g04439 ( new_n4816 , pi042 , pi219 );
  or   g04440 ( new_n4817 , new_n4813 , new_n4814 );
  nand g04441 ( new_n4818 , new_n4816 , new_n4817 );
  nand g04442 ( new_n4819 , new_n4815 , new_n4818 );
  xor  g04443 ( new_n4820 , new_n4812 , new_n4819 );
  nand g04444 ( new_n4821 , pi001 , pi051 );
  nand g04445 ( new_n4822 , pi108 , pi219 );
  nand g04446 ( new_n4823 , pi042 , pi102 );
  xor  g04447 ( new_n4824 , new_n4822 , new_n4823 );
  xnor g04448 ( new_n4825 , new_n4821 , new_n4824 );
  xnor g04449 ( new_n4826 , new_n4820 , new_n4825 );
  not  g04450 ( new_n4827 , new_n4816 );
  not  g04451 ( new_n4828 , new_n4815 );
  nand g04452 ( new_n4829 , pi051 , pi087 );
  nand g04453 ( new_n4830 , new_n4827 , new_n4829 );
  nand g04454 ( new_n4831 , new_n4828 , new_n4830 );
  nand g04455 ( new_n4832 , new_n4817 , new_n4831 );
  nand g04456 ( new_n4833 , new_n4827 , new_n4832 );
  xor  g04457 ( new_n4834 , new_n4826 , new_n4833 );
  nand g04458 ( new_n4835 , pi169 , pi188 );
  nand g04459 ( new_n4836 , pi061 , pi142 );
  nand g04460 ( new_n4837 , new_n4835 , new_n4836 );
  nand g04461 ( new_n4838 , pi071 , pi178 );
  or   g04462 ( new_n4839 , new_n4835 , new_n4836 );
  nand g04463 ( new_n4840 , new_n4838 , new_n4839 );
  nand g04464 ( new_n4841 , new_n4837 , new_n4840 );
  nand g04465 ( new_n4842 , pi012 , pi142 );
  xor  g04466 ( new_n4843 , new_n4841 , new_n4842 );
  nand g04467 ( new_n4844 , pi123 , pi188 );
  nand g04468 ( new_n4845 , pi061 , pi071 );
  nand g04469 ( new_n4846 , pi169 , pi178 );
  xor  g04470 ( new_n4847 , new_n4845 , new_n4846 );
  xor  g04471 ( new_n4848 , new_n4844 , new_n4847 );
  xor  g04472 ( new_n4849 , new_n4843 , new_n4848 );
  not  g04473 ( new_n4850 , new_n4838 );
  not  g04474 ( new_n4851 , new_n4837 );
  nand g04475 ( new_n4852 , pi142 , pi188 );
  nand g04476 ( new_n4853 , new_n4850 , new_n4852 );
  nand g04477 ( new_n4854 , new_n4851 , new_n4853 );
  nand g04478 ( new_n4855 , new_n4839 , new_n4854 );
  nand g04479 ( new_n4856 , new_n4850 , new_n4855 );
  xor  g04480 ( new_n4857 , new_n4849 , new_n4856 );
  xor  g04481 ( new_n4858 , new_n4834 , new_n4857 );
  nand g04482 ( new_n4859 , pi042 , pi087 );
  nand g04483 ( new_n4860 , pi051 , pi219 );
  xor  g04484 ( new_n4861 , new_n4859 , new_n4860 );
  nand g04485 ( new_n4862 , pi142 , pi178 );
  nand g04486 ( new_n4863 , pi071 , pi188 );
  xor  g04487 ( new_n4864 , new_n4862 , new_n4863 );
  or   g04488 ( new_n4865 , new_n4861 , new_n4864 );
  nor  g04489 ( new_n4866 , new_n4829 , new_n4852 );
  not  g04490 ( new_n4867 , new_n4866 );
  xor  g04491 ( new_n4868 , new_n4861 , new_n4864 );
  nand g04492 ( new_n4869 , new_n4867 , new_n4868 );
  nand g04493 ( new_n4870 , new_n4865 , new_n4869 );
  nor  g04494 ( new_n4871 , new_n4851 , new_n4853 );
  or   g04495 ( new_n4872 , new_n4855 , new_n4871 );
  or   g04496 ( new_n4873 , new_n4870 , new_n4872 );
  xor  g04497 ( new_n4874 , new_n4870 , new_n4872 );
  nor  g04498 ( new_n4875 , new_n4828 , new_n4830 );
  nor  g04499 ( new_n4876 , new_n4832 , new_n4875 );
  nand g04500 ( new_n4877 , new_n4874 , new_n4876 );
  nand g04501 ( new_n4878 , new_n4873 , new_n4877 );
  xor  g04502 ( new_n4879 , new_n4858 , new_n4878 );
  nand g04503 ( new_n4880 , pi033 , pi182 );
  nand g04504 ( new_n4881 , pi138 , pi179 );
  xor  g04505 ( new_n4882 , new_n4880 , new_n4881 );
  nand g04506 ( new_n4883 , pi041 , pi162 );
  xor  g04507 ( new_n4884 , new_n4882 , new_n4883 );
  nand g04508 ( new_n4885 , pi033 , pi138 );
  nand g04509 ( new_n4886 , pi162 , pi182 );
  nor  g04510 ( new_n4887 , new_n4885 , new_n4886 );
  not  g04511 ( new_n4888 , new_n4887 );
  nor  g04512 ( new_n4889 , new_n4884 , new_n4888 );
  nand g04513 ( new_n4890 , pi179 , pi182 );
  nand g04514 ( new_n4891 , pi033 , pi041 );
  nand g04515 ( new_n4892 , pi162 , pi216 );
  xor  g04516 ( new_n4893 , new_n4891 , new_n4892 );
  xor  g04517 ( new_n4894 , new_n4890 , new_n4893 );
  nand g04518 ( new_n4895 , pi048 , pi138 );
  nand g04519 ( new_n4896 , new_n4880 , new_n4881 );
  nand g04520 ( new_n4897 , new_n4882 , new_n4883 );
  nand g04521 ( new_n4898 , new_n4896 , new_n4897 );
  xor  g04522 ( new_n4899 , new_n4895 , new_n4898 );
  xor  g04523 ( new_n4900 , new_n4894 , new_n4899 );
  xor  g04524 ( new_n4901 , new_n4889 , new_n4900 );
  xnor g04525 ( new_n4902 , new_n4874 , new_n4876 );
  xor  g04526 ( new_n4903 , new_n4884 , new_n4887 );
  nor  g04527 ( new_n4904 , new_n4902 , new_n4903 );
  xnor g04528 ( new_n4905 , new_n4902 , new_n4903 );
  nand g04529 ( new_n4906 , pi138 , pi162 );
  xor  g04530 ( new_n4907 , new_n4829 , new_n4852 );
  not  g04531 ( new_n4908 , new_n4907 );
  nor  g04532 ( new_n4909 , new_n4906 , new_n4908 );
  xor  g04533 ( new_n4910 , new_n4885 , new_n4886 );
  or   g04534 ( new_n4911 , new_n4909 , new_n4910 );
  xor  g04535 ( new_n4912 , new_n4867 , new_n4868 );
  xor  g04536 ( new_n4913 , new_n4909 , new_n4910 );
  nand g04537 ( new_n4914 , new_n4912 , new_n4913 );
  nand g04538 ( new_n4915 , new_n4911 , new_n4914 );
  nor  g04539 ( new_n4916 , new_n4905 , new_n4915 );
  nor  g04540 ( new_n4917 , new_n4904 , new_n4916 );
  xor  g04541 ( new_n4918 , new_n4901 , new_n4917 );
  xor  g04542 ( new_n4919 , new_n4879 , new_n4918 );
  nand g04543 ( new_n4920 , pi020 , pi057 );
  nand g04544 ( new_n4921 , pi160 , pi194 );
  xor  g04545 ( new_n4922 , new_n4920 , new_n4921 );
  nand g04546 ( new_n4923 , pi060 , pi143 );
  xor  g04547 ( new_n4924 , new_n4922 , new_n4923 );
  nand g04548 ( new_n4925 , pi143 , pi160 );
  or   g04549 ( new_n4926 , new_n4920 , new_n4925 );
  nor  g04550 ( new_n4927 , new_n4924 , new_n4926 );
  nand g04551 ( new_n4928 , pi020 , pi194 );
  nand g04552 ( new_n4929 , pi143 , pi223 );
  nand g04553 ( new_n4930 , pi057 , pi060 );
  xor  g04554 ( new_n4931 , new_n4929 , new_n4930 );
  xor  g04555 ( new_n4932 , new_n4928 , new_n4931 );
  nand g04556 ( new_n4933 , pi085 , pi160 );
  nand g04557 ( new_n4934 , new_n4920 , new_n4921 );
  nand g04558 ( new_n4935 , new_n4922 , new_n4923 );
  nand g04559 ( new_n4936 , new_n4934 , new_n4935 );
  xor  g04560 ( new_n4937 , new_n4933 , new_n4936 );
  xor  g04561 ( new_n4938 , new_n4932 , new_n4937 );
  xor  g04562 ( new_n4939 , new_n4927 , new_n4938 );
  xor  g04563 ( new_n4940 , new_n4924 , new_n4926 );
  xor  g04564 ( new_n4941 , new_n4906 , new_n4907 );
  or   g04565 ( new_n4942 , new_n4925 , new_n4941 );
  nand g04566 ( new_n4943 , pi057 , pi160 );
  nand g04567 ( new_n4944 , pi020 , pi143 );
  nand g04568 ( new_n4945 , new_n4943 , new_n4944 );
  nand g04569 ( new_n4946 , new_n4926 , new_n4945 );
  or   g04570 ( new_n4947 , new_n4942 , new_n4946 );
  xnor g04571 ( new_n4948 , new_n4912 , new_n4913 );
  xor  g04572 ( new_n4949 , new_n4942 , new_n4946 );
  nand g04573 ( new_n4950 , new_n4948 , new_n4949 );
  nand g04574 ( new_n4951 , new_n4947 , new_n4950 );
  or   g04575 ( new_n4952 , new_n4940 , new_n4951 );
  xor  g04576 ( new_n4953 , new_n4905 , new_n4915 );
  not  g04577 ( new_n4954 , new_n4953 );
  xor  g04578 ( new_n4955 , new_n4940 , new_n4951 );
  nand g04579 ( new_n4956 , new_n4954 , new_n4955 );
  nand g04580 ( new_n4957 , new_n4952 , new_n4956 );
  xor  g04581 ( new_n4958 , new_n4939 , new_n4957 );
  xor  g04582 ( po016 , new_n4919 , new_n4958 );
  nand g04583 ( new_n4960 , pi163 , pi226 );
  nand g04584 ( new_n4961 , pi107 , pi109 );
  nor  g04585 ( new_n4962 , new_n4960 , new_n4961 );
  nand g04586 ( new_n4963 , pi148 , pi226 );
  nand g04587 ( new_n4964 , pi163 , pi207 );
  nand g04588 ( new_n4965 , new_n4963 , new_n4964 );
  nand g04589 ( new_n4966 , pi148 , pi207 );
  nor  g04590 ( new_n4967 , new_n4960 , new_n4966 );
  not  g04591 ( new_n4968 , new_n4967 );
  nand g04592 ( new_n4969 , new_n4965 , new_n4968 );
  xor  g04593 ( new_n4970 , new_n4962 , new_n4969 );
  nand g04594 ( new_n4971 , pi014 , pi107 );
  nand g04595 ( new_n4972 , pi109 , pi171 );
  nand g04596 ( new_n4973 , new_n4971 , new_n4972 );
  nand g04597 ( new_n4974 , pi014 , pi171 );
  nor  g04598 ( new_n4975 , new_n4961 , new_n4974 );
  not  g04599 ( new_n4976 , new_n4975 );
  nand g04600 ( new_n4977 , new_n4973 , new_n4976 );
  xor  g04601 ( new_n4978 , new_n4970 , new_n4977 );
  xor  g04602 ( new_n4979 , new_n4960 , new_n4961 );
  not  g04603 ( new_n4980 , new_n4979 );
  nand g04604 ( new_n4981 , pi132 , pi175 );
  or   g04605 ( new_n4982 , new_n4980 , new_n4981 );
  nand g04606 ( new_n4983 , pi175 , pi186 );
  nand g04607 ( new_n4984 , pi132 , pi134 );
  and  g04608 ( new_n4985 , new_n4983 , new_n4984 );
  nand g04609 ( new_n4986 , pi134 , pi186 );
  nor  g04610 ( new_n4987 , new_n4981 , new_n4986 );
  or   g04611 ( new_n4988 , new_n4985 , new_n4987 );
  xor  g04612 ( new_n4989 , new_n4982 , new_n4988 );
  xor  g04613 ( new_n4990 , new_n4978 , new_n4989 );
  xor  g04614 ( new_n4991 , new_n4979 , new_n4981 );
  nand g04615 ( new_n4992 , pi029 , pi103 );
  nor  g04616 ( new_n4993 , new_n4991 , new_n4992 );
  nand g04617 ( new_n4994 , pi029 , pi117 );
  nand g04618 ( new_n4995 , pi069 , pi103 );
  xor  g04619 ( new_n4996 , new_n4994 , new_n4995 );
  xor  g04620 ( new_n4997 , new_n4993 , new_n4996 );
  xor  g04621 ( po017 , new_n4990 , new_n4997 );
  xor  g04622 ( po018 , new_n3112 , new_n3113 );
  nand g04623 ( new_n5000 , pi141 , pi173 );
  nand g04624 ( new_n5001 , pi014 , pi090 );
  nand g04625 ( new_n5002 , pi047 , pi109 );
  nand g04626 ( new_n5003 , new_n5001 , new_n5002 );
  nand g04627 ( new_n5004 , pi090 , pi109 );
  nand g04628 ( new_n5005 , pi014 , pi047 );
  or   g04629 ( new_n5006 , new_n5004 , new_n5005 );
  nand g04630 ( new_n5007 , new_n5003 , new_n5006 );
  xor  g04631 ( new_n5008 , new_n5000 , new_n5007 );
  nand g04632 ( new_n5009 , pi014 , pi141 );
  nand g04633 ( new_n5010 , new_n5004 , new_n5009 );
  nand g04634 ( new_n5011 , pi161 , pi173 );
  xor  g04635 ( new_n5012 , new_n5004 , new_n5009 );
  nand g04636 ( new_n5013 , new_n5011 , new_n5012 );
  nand g04637 ( new_n5014 , new_n5010 , new_n5013 );
  xor  g04638 ( new_n5015 , new_n5008 , new_n5014 );
  nand g04639 ( new_n5016 , pi161 , pi230 );
  nand g04640 ( new_n5017 , pi050 , pi241 );
  and  g04641 ( new_n5018 , new_n5016 , new_n5017 );
  nand g04642 ( new_n5019 , pi230 , pi241 );
  nand g04643 ( new_n5020 , pi050 , pi161 );
  nor  g04644 ( new_n5021 , new_n5019 , new_n5020 );
  or   g04645 ( new_n5022 , new_n5018 , new_n5021 );
  xnor g04646 ( new_n5023 , new_n5015 , new_n5022 );
  nand g04647 ( new_n5024 , new_n3130 , new_n3131 );
  nand g04648 ( new_n5025 , new_n3129 , new_n3132 );
  nand g04649 ( new_n5026 , new_n5024 , new_n5025 );
  nand g04650 ( new_n5027 , new_n5019 , new_n5026 );
  xor  g04651 ( new_n5028 , new_n5011 , new_n5012 );
  xor  g04652 ( new_n5029 , new_n5019 , new_n5026 );
  nand g04653 ( new_n5030 , new_n5028 , new_n5029 );
  nand g04654 ( new_n5031 , new_n5027 , new_n5030 );
  xor  g04655 ( new_n5032 , new_n5023 , new_n5031 );
  xor  g04656 ( new_n5033 , new_n5028 , new_n5029 );
  nand g04657 ( new_n5034 , pi050 , pi236 );
  or   g04658 ( new_n5035 , new_n5033 , new_n5034 );
  xor  g04659 ( new_n5036 , new_n5033 , new_n5034 );
  or   g04660 ( new_n5037 , new_n3120 , new_n3127 );
  nand g04661 ( new_n5038 , new_n3128 , new_n3133 );
  nand g04662 ( new_n5039 , new_n5037 , new_n5038 );
  nand g04663 ( new_n5040 , new_n5036 , new_n5039 );
  nand g04664 ( new_n5041 , new_n5035 , new_n5040 );
  nand g04665 ( new_n5042 , new_n5032 , new_n5041 );
  nand g04666 ( new_n5043 , pi090 , pi173 );
  nand g04667 ( new_n5044 , pi018 , pi109 );
  xor  g04668 ( new_n5045 , new_n5043 , new_n5044 );
  xor  g04669 ( new_n5046 , new_n5005 , new_n5045 );
  nand g04670 ( new_n5047 , pi141 , pi230 );
  xor  g04671 ( new_n5048 , new_n5006 , new_n5047 );
  xor  g04672 ( new_n5049 , new_n5046 , new_n5048 );
  nand g04673 ( new_n5050 , pi241 , pi253 );
  nand g04674 ( new_n5051 , pi074 , pi236 );
  xor  g04675 ( new_n5052 , new_n5050 , new_n5051 );
  xor  g04676 ( new_n5053 , new_n5020 , new_n5052 );
  nand g04677 ( new_n5054 , new_n5000 , new_n5007 );
  nand g04678 ( new_n5055 , new_n5008 , new_n5014 );
  nand g04679 ( new_n5056 , new_n5054 , new_n5055 );
  xor  g04680 ( new_n5057 , new_n5053 , new_n5056 );
  xnor g04681 ( new_n5058 , new_n5049 , new_n5057 );
  nor  g04682 ( new_n5059 , new_n5015 , new_n5022 );
  nor  g04683 ( new_n5060 , new_n5023 , new_n5031 );
  xor  g04684 ( new_n5061 , new_n5021 , new_n5060 );
  nor  g04685 ( new_n5062 , new_n5059 , new_n5061 );
  xor  g04686 ( new_n5063 , new_n5058 , new_n5062 );
  xnor g04687 ( new_n5064 , new_n5042 , new_n5063 );
  nand g04688 ( new_n5065 , pi236 , pi253 );
  nor  g04689 ( new_n5066 , new_n3134 , new_n3181 );
  xor  g04690 ( new_n5067 , new_n5036 , new_n5039 );
  nand g04691 ( new_n5068 , new_n5066 , new_n5067 );
  nand g04692 ( new_n5069 , new_n5065 , new_n5068 );
  xnor g04693 ( new_n5070 , new_n5032 , new_n5041 );
  xor  g04694 ( new_n5071 , new_n5065 , new_n5068 );
  nand g04695 ( new_n5072 , new_n5070 , new_n5071 );
  nand g04696 ( new_n5073 , new_n5069 , new_n5072 );
  xnor g04697 ( new_n5074 , new_n5064 , new_n5073 );
  nand g04698 ( new_n5075 , pi013 , pi066 );
  nand g04699 ( new_n5076 , pi013 , pi207 );
  nand g04700 ( new_n5077 , pi066 , pi104 );
  nand g04701 ( new_n5078 , new_n5076 , new_n5077 );
  nand g04702 ( new_n5079 , pi112 , pi226 );
  xor  g04703 ( new_n5080 , new_n5076 , new_n5077 );
  nand g04704 ( new_n5081 , new_n5079 , new_n5080 );
  nand g04705 ( new_n5082 , new_n5078 , new_n5081 );
  nand g04706 ( new_n5083 , pi105 , pi226 );
  nand g04707 ( new_n5084 , pi112 , pi207 );
  nand g04708 ( new_n5085 , new_n5083 , new_n5084 );
  nand g04709 ( new_n5086 , pi105 , pi207 );
  or   g04710 ( new_n5087 , new_n5079 , new_n5086 );
  nand g04711 ( new_n5088 , new_n5085 , new_n5087 );
  xor  g04712 ( new_n5089 , new_n5082 , new_n5088 );
  xor  g04713 ( new_n5090 , new_n5075 , new_n5089 );
  nand g04714 ( new_n5091 , pi055 , pi104 );
  nand g04715 ( new_n5092 , pi002 , pi212 );
  nand g04716 ( new_n5093 , new_n5091 , new_n5092 );
  nand g04717 ( new_n5094 , pi055 , pi212 );
  nand g04718 ( new_n5095 , pi002 , pi104 );
  nor  g04719 ( new_n5096 , new_n5094 , new_n5095 );
  not  g04720 ( new_n5097 , new_n5096 );
  nand g04721 ( new_n5098 , new_n5093 , new_n5097 );
  xnor g04722 ( new_n5099 , new_n5090 , new_n5098 );
  nand g04723 ( new_n5100 , new_n3150 , new_n3151 );
  nand g04724 ( new_n5101 , new_n3149 , new_n3152 );
  nand g04725 ( new_n5102 , new_n5100 , new_n5101 );
  nand g04726 ( new_n5103 , new_n5094 , new_n5102 );
  xor  g04727 ( new_n5104 , new_n5079 , new_n5080 );
  xor  g04728 ( new_n5105 , new_n5094 , new_n5102 );
  nand g04729 ( new_n5106 , new_n5104 , new_n5105 );
  nand g04730 ( new_n5107 , new_n5103 , new_n5106 );
  xor  g04731 ( new_n5108 , new_n5099 , new_n5107 );
  nand g04732 ( new_n5109 , pi002 , pi213 );
  nand g04733 ( new_n5110 , new_n3154 , new_n3157 );
  nand g04734 ( new_n5111 , new_n3153 , new_n3158 );
  nand g04735 ( new_n5112 , new_n5110 , new_n5111 );
  or   g04736 ( new_n5113 , new_n5109 , new_n5112 );
  xor  g04737 ( new_n5114 , new_n5104 , new_n5105 );
  not  g04738 ( new_n5115 , new_n5114 );
  xor  g04739 ( new_n5116 , new_n5109 , new_n5112 );
  nand g04740 ( new_n5117 , new_n5115 , new_n5116 );
  nand g04741 ( new_n5118 , new_n5113 , new_n5117 );
  nand g04742 ( new_n5119 , new_n5108 , new_n5118 );
  nand g04743 ( new_n5120 , pi183 , pi226 );
  nand g04744 ( new_n5121 , pi066 , pi112 );
  xor  g04745 ( new_n5122 , new_n5120 , new_n5121 );
  xor  g04746 ( new_n5123 , new_n5086 , new_n5122 );
  nand g04747 ( new_n5124 , pi013 , pi055 );
  xor  g04748 ( new_n5125 , new_n5087 , new_n5124 );
  xor  g04749 ( new_n5126 , new_n5123 , new_n5125 );
  nand g04750 ( new_n5127 , pi025 , pi212 );
  nand g04751 ( new_n5128 , pi213 , pi239 );
  xor  g04752 ( new_n5129 , new_n5127 , new_n5128 );
  xor  g04753 ( new_n5130 , new_n5095 , new_n5129 );
  nand g04754 ( new_n5131 , new_n5082 , new_n5088 );
  nand g04755 ( new_n5132 , new_n5075 , new_n5089 );
  nand g04756 ( new_n5133 , new_n5131 , new_n5132 );
  xor  g04757 ( new_n5134 , new_n5130 , new_n5133 );
  xnor g04758 ( new_n5135 , new_n5126 , new_n5134 );
  nor  g04759 ( new_n5136 , new_n5099 , new_n5107 );
  and  g04760 ( new_n5137 , new_n5096 , new_n5136 );
  or   g04761 ( new_n5138 , new_n5090 , new_n5098 );
  nand g04762 ( new_n5139 , new_n5097 , new_n5138 );
  nor  g04763 ( new_n5140 , new_n5136 , new_n5139 );
  or   g04764 ( new_n5141 , new_n5137 , new_n5140 );
  xor  g04765 ( new_n5142 , new_n5135 , new_n5141 );
  xor  g04766 ( new_n5143 , new_n5119 , new_n5142 );
  nand g04767 ( new_n5144 , pi025 , pi213 );
  xnor g04768 ( new_n5145 , new_n5108 , new_n5118 );
  or   g04769 ( new_n5146 , new_n5144 , new_n5145 );
  nand g04770 ( new_n5147 , new_n3148 , new_n3160 );
  xor  g04771 ( new_n5148 , new_n5114 , new_n5116 );
  nor  g04772 ( new_n5149 , new_n5147 , new_n5148 );
  xor  g04773 ( new_n5150 , new_n5144 , new_n5145 );
  nand g04774 ( new_n5151 , new_n5149 , new_n5150 );
  nand g04775 ( new_n5152 , new_n5146 , new_n5151 );
  xor  g04776 ( new_n5153 , new_n5143 , new_n5152 );
  xor  g04777 ( new_n5154 , new_n5074 , new_n5153 );
  xnor g04778 ( new_n5155 , new_n5070 , new_n5071 );
  xor  g04779 ( new_n5156 , new_n5149 , new_n5150 );
  nand g04780 ( new_n5157 , new_n5155 , new_n5156 );
  xor  g04781 ( new_n5158 , new_n5155 , new_n5156 );
  xor  g04782 ( new_n5159 , new_n5066 , new_n5067 );
  xor  g04783 ( new_n5160 , new_n5147 , new_n5148 );
  nand g04784 ( new_n5161 , new_n5159 , new_n5160 );
  xor  g04785 ( new_n5162 , new_n5159 , new_n5160 );
  not  g04786 ( new_n5163 , new_n3161 );
  nor  g04787 ( new_n5164 , new_n3139 , new_n5163 );
  nor  g04788 ( new_n5165 , new_n3162 , new_n3186 );
  nor  g04789 ( new_n5166 , new_n5164 , new_n5165 );
  not  g04790 ( new_n5167 , new_n5166 );
  nand g04791 ( new_n5168 , new_n5162 , new_n5167 );
  nand g04792 ( new_n5169 , new_n5161 , new_n5168 );
  nand g04793 ( new_n5170 , new_n5158 , new_n5169 );
  nand g04794 ( new_n5171 , new_n5157 , new_n5170 );
  xnor g04795 ( new_n5172 , new_n5154 , new_n5171 );
  nand g04796 ( new_n5173 , pi035 , pi058 );
  nand g04797 ( new_n5174 , pi132 , pi204 );
  nand g04798 ( new_n5175 , pi015 , pi186 );
  nand g04799 ( new_n5176 , new_n5174 , new_n5175 );
  nand g04800 ( new_n5177 , pi015 , pi132 );
  nand g04801 ( new_n5178 , pi186 , pi204 );
  or   g04802 ( new_n5179 , new_n5177 , new_n5178 );
  nand g04803 ( new_n5180 , new_n5176 , new_n5179 );
  xor  g04804 ( new_n5181 , new_n5173 , new_n5180 );
  nand g04805 ( new_n5182 , pi035 , pi186 );
  nand g04806 ( new_n5183 , new_n5177 , new_n5182 );
  nand g04807 ( new_n5184 , pi058 , pi139 );
  xor  g04808 ( new_n5185 , new_n5177 , new_n5182 );
  nand g04809 ( new_n5186 , new_n5184 , new_n5185 );
  nand g04810 ( new_n5187 , new_n5183 , new_n5186 );
  xor  g04811 ( new_n5188 , new_n5181 , new_n5187 );
  nand g04812 ( new_n5189 , pi139 , pi211 );
  nand g04813 ( new_n5190 , pi199 , pi208 );
  and  g04814 ( new_n5191 , new_n5189 , new_n5190 );
  nand g04815 ( new_n5192 , pi208 , pi211 );
  nand g04816 ( new_n5193 , pi139 , pi199 );
  nor  g04817 ( new_n5194 , new_n5192 , new_n5193 );
  or   g04818 ( new_n5195 , new_n5191 , new_n5194 );
  xnor g04819 ( new_n5196 , new_n5188 , new_n5195 );
  nand g04820 ( new_n5197 , new_n3202 , new_n3203 );
  nand g04821 ( new_n5198 , new_n3201 , new_n3204 );
  nand g04822 ( new_n5199 , new_n5197 , new_n5198 );
  nand g04823 ( new_n5200 , new_n5192 , new_n5199 );
  xor  g04824 ( new_n5201 , new_n5184 , new_n5185 );
  xor  g04825 ( new_n5202 , new_n5192 , new_n5199 );
  nand g04826 ( new_n5203 , new_n5201 , new_n5202 );
  nand g04827 ( new_n5204 , new_n5200 , new_n5203 );
  xor  g04828 ( new_n5205 , new_n5196 , new_n5204 );
  xor  g04829 ( new_n5206 , new_n5201 , new_n5202 );
  nand g04830 ( new_n5207 , pi168 , pi199 );
  or   g04831 ( new_n5208 , new_n5206 , new_n5207 );
  xor  g04832 ( new_n5209 , new_n5206 , new_n5207 );
  or   g04833 ( new_n5210 , new_n3196 , new_n3199 );
  nand g04834 ( new_n5211 , new_n3200 , new_n3205 );
  nand g04835 ( new_n5212 , new_n5210 , new_n5211 );
  nand g04836 ( new_n5213 , new_n5209 , new_n5212 );
  nand g04837 ( new_n5214 , new_n5208 , new_n5213 );
  nand g04838 ( new_n5215 , new_n5205 , new_n5214 );
  nand g04839 ( new_n5216 , pi132 , pi146 );
  nand g04840 ( new_n5217 , pi015 , pi058 );
  xor  g04841 ( new_n5218 , new_n5216 , new_n5217 );
  xor  g04842 ( new_n5219 , new_n5178 , new_n5218 );
  nand g04843 ( new_n5220 , pi035 , pi211 );
  xor  g04844 ( new_n5221 , new_n5179 , new_n5220 );
  xor  g04845 ( new_n5222 , new_n5219 , new_n5221 );
  nand g04846 ( new_n5223 , pi195 , pi208 );
  nand g04847 ( new_n5224 , pi168 , pi218 );
  xor  g04848 ( new_n5225 , new_n5223 , new_n5224 );
  xor  g04849 ( new_n5226 , new_n5193 , new_n5225 );
  nand g04850 ( new_n5227 , new_n5173 , new_n5180 );
  nand g04851 ( new_n5228 , new_n5181 , new_n5187 );
  nand g04852 ( new_n5229 , new_n5227 , new_n5228 );
  xor  g04853 ( new_n5230 , new_n5226 , new_n5229 );
  xnor g04854 ( new_n5231 , new_n5222 , new_n5230 );
  nor  g04855 ( new_n5232 , new_n5188 , new_n5195 );
  nor  g04856 ( new_n5233 , new_n5196 , new_n5204 );
  xor  g04857 ( new_n5234 , new_n5194 , new_n5233 );
  nor  g04858 ( new_n5235 , new_n5232 , new_n5234 );
  xor  g04859 ( new_n5236 , new_n5231 , new_n5235 );
  nand g04860 ( new_n5237 , pi168 , pi195 );
  nor  g04861 ( new_n5238 , new_n3195 , new_n3206 );
  xor  g04862 ( new_n5239 , new_n5209 , new_n5212 );
  nand g04863 ( new_n5240 , new_n5238 , new_n5239 );
  nand g04864 ( new_n5241 , new_n5237 , new_n5240 );
  xnor g04865 ( new_n5242 , new_n5205 , new_n5214 );
  xor  g04866 ( new_n5243 , new_n5237 , new_n5240 );
  nand g04867 ( new_n5244 , new_n5242 , new_n5243 );
  nand g04868 ( new_n5245 , new_n5241 , new_n5244 );
  xor  g04869 ( new_n5246 , new_n5236 , new_n5245 );
  xor  g04870 ( new_n5247 , new_n5215 , new_n5246 );
  xor  g04871 ( new_n5248 , new_n5172 , new_n5247 );
  xor  g04872 ( new_n5249 , new_n5158 , new_n5169 );
  not  g04873 ( new_n5250 , new_n5249 );
  xor  g04874 ( new_n5251 , new_n5242 , new_n5243 );
  or   g04875 ( new_n5252 , new_n5250 , new_n5251 );
  xor  g04876 ( new_n5253 , new_n5250 , new_n5251 );
  xor  g04877 ( new_n5254 , new_n5162 , new_n5167 );
  xor  g04878 ( new_n5255 , new_n5238 , new_n5239 );
  nand g04879 ( new_n5256 , new_n5254 , new_n5255 );
  not  g04880 ( new_n5257 , new_n5256 );
  xnor g04881 ( new_n5258 , new_n5254 , new_n5255 );
  or   g04882 ( new_n5259 , new_n3207 , new_n3226 );
  not  g04883 ( new_n5260 , new_n3187 );
  nand g04884 ( new_n5261 , new_n5260 , new_n3227 );
  nand g04885 ( new_n5262 , new_n5259 , new_n5261 );
  nor  g04886 ( new_n5263 , new_n5258 , new_n5262 );
  nor  g04887 ( new_n5264 , new_n5257 , new_n5263 );
  not  g04888 ( new_n5265 , new_n5264 );
  nand g04889 ( new_n5266 , new_n5253 , new_n5265 );
  nand g04890 ( new_n5267 , new_n5252 , new_n5266 );
  xnor g04891 ( new_n5268 , new_n5248 , new_n5267 );
  nand g04892 ( new_n5269 , pi133 , pi244 );
  nand g04893 ( new_n5270 , pi069 , pi189 );
  nand g04894 ( new_n5271 , pi029 , pi064 );
  nand g04895 ( new_n5272 , new_n5270 , new_n5271 );
  nand g04896 ( new_n5273 , pi029 , pi189 );
  nand g04897 ( new_n5274 , pi064 , pi069 );
  or   g04898 ( new_n5275 , new_n5273 , new_n5274 );
  nand g04899 ( new_n5276 , new_n5272 , new_n5275 );
  xor  g04900 ( new_n5277 , new_n5269 , new_n5276 );
  nand g04901 ( new_n5278 , pi077 , pi244 );
  nand g04902 ( new_n5279 , pi069 , pi133 );
  nand g04903 ( new_n5280 , new_n5278 , new_n5279 );
  xor  g04904 ( new_n5281 , new_n5278 , new_n5279 );
  nand g04905 ( new_n5282 , new_n5273 , new_n5281 );
  nand g04906 ( new_n5283 , new_n5280 , new_n5282 );
  xor  g04907 ( new_n5284 , new_n5277 , new_n5283 );
  nand g04908 ( new_n5285 , pi077 , pi150 );
  nand g04909 ( new_n5286 , pi052 , pi221 );
  and  g04910 ( new_n5287 , new_n5285 , new_n5286 );
  nand g04911 ( new_n5288 , pi052 , pi150 );
  nand g04912 ( new_n5289 , pi077 , pi221 );
  nor  g04913 ( new_n5290 , new_n5288 , new_n5289 );
  or   g04914 ( new_n5291 , new_n5287 , new_n5290 );
  xnor g04915 ( new_n5292 , new_n5284 , new_n5291 );
  nand g04916 ( new_n5293 , new_n3239 , new_n3240 );
  nand g04917 ( new_n5294 , new_n3238 , new_n3241 );
  nand g04918 ( new_n5295 , new_n5293 , new_n5294 );
  nand g04919 ( new_n5296 , new_n5288 , new_n5295 );
  xor  g04920 ( new_n5297 , new_n5273 , new_n5281 );
  xor  g04921 ( new_n5298 , new_n5288 , new_n5295 );
  nand g04922 ( new_n5299 , new_n5297 , new_n5298 );
  nand g04923 ( new_n5300 , new_n5296 , new_n5299 );
  xor  g04924 ( new_n5301 , new_n5292 , new_n5300 );
  nand g04925 ( new_n5302 , pi131 , pi221 );
  nand g04926 ( new_n5303 , new_n3243 , new_n3246 );
  nand g04927 ( new_n5304 , new_n3242 , new_n3247 );
  nand g04928 ( new_n5305 , new_n5303 , new_n5304 );
  or   g04929 ( new_n5306 , new_n5302 , new_n5305 );
  xnor g04930 ( new_n5307 , new_n5297 , new_n5298 );
  xor  g04931 ( new_n5308 , new_n5302 , new_n5305 );
  nand g04932 ( new_n5309 , new_n5307 , new_n5308 );
  nand g04933 ( new_n5310 , new_n5306 , new_n5309 );
  nand g04934 ( new_n5311 , new_n5301 , new_n5310 );
  nand g04935 ( new_n5312 , pi029 , pi084 );
  nand g04936 ( new_n5313 , pi189 , pi244 );
  xor  g04937 ( new_n5314 , new_n5312 , new_n5313 );
  xor  g04938 ( new_n5315 , new_n5274 , new_n5314 );
  nand g04939 ( new_n5316 , pi133 , pi150 );
  xor  g04940 ( new_n5317 , new_n5275 , new_n5316 );
  xor  g04941 ( new_n5318 , new_n5315 , new_n5317 );
  nand g04942 ( new_n5319 , pi052 , pi196 );
  nand g04943 ( new_n5320 , pi131 , pi184 );
  xor  g04944 ( new_n5321 , new_n5319 , new_n5320 );
  xor  g04945 ( new_n5322 , new_n5289 , new_n5321 );
  nand g04946 ( new_n5323 , new_n5269 , new_n5276 );
  nand g04947 ( new_n5324 , new_n5277 , new_n5283 );
  nand g04948 ( new_n5325 , new_n5323 , new_n5324 );
  xor  g04949 ( new_n5326 , new_n5322 , new_n5325 );
  xnor g04950 ( new_n5327 , new_n5318 , new_n5326 );
  nor  g04951 ( new_n5328 , new_n5284 , new_n5291 );
  nor  g04952 ( new_n5329 , new_n5292 , new_n5300 );
  xor  g04953 ( new_n5330 , new_n5290 , new_n5329 );
  nor  g04954 ( new_n5331 , new_n5328 , new_n5330 );
  not  g04955 ( new_n5332 , new_n5331 );
  xor  g04956 ( new_n5333 , new_n5327 , new_n5332 );
  xor  g04957 ( new_n5334 , new_n5311 , new_n5333 );
  nand g04958 ( new_n5335 , pi131 , pi196 );
  not  g04959 ( new_n5336 , new_n3237 );
  nor  g04960 ( new_n5337 , new_n5336 , new_n3248 );
  xor  g04961 ( new_n5338 , new_n5307 , new_n5308 );
  nand g04962 ( new_n5339 , new_n5337 , new_n5338 );
  nand g04963 ( new_n5340 , new_n5335 , new_n5339 );
  xor  g04964 ( new_n5341 , new_n5301 , new_n5310 );
  not  g04965 ( new_n5342 , new_n5341 );
  xor  g04966 ( new_n5343 , new_n5335 , new_n5339 );
  nand g04967 ( new_n5344 , new_n5342 , new_n5343 );
  nand g04968 ( new_n5345 , new_n5340 , new_n5344 );
  xor  g04969 ( new_n5346 , new_n5334 , new_n5345 );
  xor  g04970 ( new_n5347 , new_n5268 , new_n5346 );
  xor  g04971 ( new_n5348 , new_n5253 , new_n5264 );
  xor  g04972 ( new_n5349 , new_n5337 , new_n5338 );
  or   g04973 ( new_n5350 , new_n3249 , new_n3268 );
  nand g04974 ( new_n5351 , new_n3228 , new_n3269 );
  nand g04975 ( new_n5352 , new_n5350 , new_n5351 );
  or   g04976 ( new_n5353 , new_n5349 , new_n5352 );
  xor  g04977 ( new_n5354 , new_n5258 , new_n5262 );
  not  g04978 ( new_n5355 , new_n5354 );
  xor  g04979 ( new_n5356 , new_n5349 , new_n5352 );
  nand g04980 ( new_n5357 , new_n5355 , new_n5356 );
  nand g04981 ( new_n5358 , new_n5353 , new_n5357 );
  or   g04982 ( new_n5359 , new_n5348 , new_n5358 );
  xor  g04983 ( new_n5360 , new_n5341 , new_n5343 );
  xor  g04984 ( new_n5361 , new_n5348 , new_n5358 );
  nand g04985 ( new_n5362 , new_n5360 , new_n5361 );
  nand g04986 ( new_n5363 , new_n5359 , new_n5362 );
  xor  g04987 ( po019 , new_n5347 , new_n5363 );
  xor  g04988 ( po020 , new_n3264 , new_n3266 );
  nand g04989 ( new_n5366 , pi028 , pi087 );
  nand g04990 ( new_n5367 , pi102 , pi113 );
  nand g04991 ( new_n5368 , pi001 , pi007 );
  nand g04992 ( new_n5369 , pi051 , pi122 );
  nand g04993 ( new_n5370 , pi042 , pi135 );
  or   g04994 ( new_n5371 , new_n5369 , new_n5370 );
  or   g04995 ( new_n5372 , new_n5368 , new_n5371 );
  nand g04996 ( new_n5373 , pi051 , pi059 );
  nand g04997 ( new_n5374 , pi108 , pi122 );
  xor  g04998 ( new_n5375 , new_n5373 , new_n5374 );
  xor  g04999 ( new_n5376 , new_n5370 , new_n5375 );
  not  g05000 ( new_n5377 , new_n5376 );
  xor  g05001 ( new_n5378 , new_n5368 , new_n5371 );
  nand g05002 ( new_n5379 , new_n5377 , new_n5378 );
  nand g05003 ( new_n5380 , new_n5372 , new_n5379 );
  xor  g05004 ( new_n5381 , new_n5367 , new_n5380 );
  nand g05005 ( new_n5382 , pi060 , pi180 );
  nand g05006 ( new_n5383 , pi020 , pi085 );
  nor  g05007 ( new_n5384 , new_n5382 , new_n5383 );
  nand g05008 ( new_n5385 , pi194 , pi223 );
  nand g05009 ( new_n5386 , pi143 , pi225 );
  nand g05010 ( new_n5387 , pi057 , pi101 );
  nand g05011 ( new_n5388 , new_n5386 , new_n5387 );
  nand g05012 ( new_n5389 , pi101 , pi143 );
  nand g05013 ( new_n5390 , pi057 , pi225 );
  or   g05014 ( new_n5391 , new_n5389 , new_n5390 );
  nand g05015 ( new_n5392 , new_n5388 , new_n5391 );
  xor  g05016 ( new_n5393 , new_n5385 , new_n5392 );
  nand g05017 ( new_n5394 , pi057 , pi223 );
  nand g05018 ( new_n5395 , new_n5389 , new_n5394 );
  nand g05019 ( new_n5396 , pi060 , pi194 );
  xor  g05020 ( new_n5397 , new_n5389 , new_n5394 );
  nand g05021 ( new_n5398 , new_n5396 , new_n5397 );
  nand g05022 ( new_n5399 , new_n5395 , new_n5398 );
  xor  g05023 ( new_n5400 , new_n5393 , new_n5399 );
  nand g05024 ( new_n5401 , pi020 , pi180 );
  nand g05025 ( new_n5402 , pi060 , pi085 );
  and  g05026 ( new_n5403 , new_n5401 , new_n5402 );
  or   g05027 ( new_n5404 , new_n5384 , new_n5403 );
  xnor g05028 ( new_n5405 , new_n5400 , new_n5404 );
  nand g05029 ( new_n5406 , new_n4929 , new_n4930 );
  nand g05030 ( new_n5407 , new_n4928 , new_n4931 );
  nand g05031 ( new_n5408 , new_n5406 , new_n5407 );
  nand g05032 ( new_n5409 , new_n5383 , new_n5408 );
  xor  g05033 ( new_n5410 , new_n5396 , new_n5397 );
  xor  g05034 ( new_n5411 , new_n5383 , new_n5408 );
  nand g05035 ( new_n5412 , new_n5410 , new_n5411 );
  nand g05036 ( new_n5413 , new_n5409 , new_n5412 );
  nor  g05037 ( new_n5414 , new_n5405 , new_n5413 );
  nand g05038 ( new_n5415 , new_n5384 , new_n5414 );
  nand g05039 ( new_n5416 , pi143 , pi177 );
  nand g05040 ( new_n5417 , pi101 , pi194 );
  xor  g05041 ( new_n5418 , new_n5416 , new_n5417 );
  xor  g05042 ( new_n5419 , new_n5390 , new_n5418 );
  nand g05043 ( new_n5420 , pi085 , pi223 );
  xor  g05044 ( new_n5421 , new_n5391 , new_n5420 );
  not  g05045 ( new_n5422 , new_n5421 );
  xor  g05046 ( new_n5423 , new_n5419 , new_n5422 );
  nand g05047 ( new_n5424 , pi068 , pi160 );
  nand g05048 ( new_n5425 , pi020 , pi036 );
  xor  g05049 ( new_n5426 , new_n5424 , new_n5425 );
  xor  g05050 ( new_n5427 , new_n5382 , new_n5426 );
  nand g05051 ( new_n5428 , new_n5385 , new_n5392 );
  nand g05052 ( new_n5429 , new_n5393 , new_n5399 );
  nand g05053 ( new_n5430 , new_n5428 , new_n5429 );
  xor  g05054 ( new_n5431 , new_n5427 , new_n5430 );
  xor  g05055 ( new_n5432 , new_n5423 , new_n5431 );
  nor  g05056 ( new_n5433 , new_n5400 , new_n5404 );
  xor  g05057 ( new_n5434 , new_n5384 , new_n5414 );
  nor  g05058 ( new_n5435 , new_n5433 , new_n5434 );
  not  g05059 ( new_n5436 , new_n5435 );
  nand g05060 ( new_n5437 , new_n5432 , new_n5436 );
  nand g05061 ( new_n5438 , new_n5415 , new_n5437 );
  nand g05062 ( new_n5439 , pi137 , pi143 );
  nand g05063 ( new_n5440 , pi046 , pi160 );
  xnor g05064 ( new_n5441 , new_n5439 , new_n5440 );
  xor  g05065 ( new_n5442 , new_n5438 , new_n5441 );
  nand g05066 ( new_n5443 , new_n5373 , new_n5374 );
  nand g05067 ( new_n5444 , new_n5370 , new_n5375 );
  nand g05068 ( new_n5445 , new_n5443 , new_n5444 );
  xor  g05069 ( new_n5446 , new_n5432 , new_n5435 );
  nand g05070 ( new_n5447 , pi036 , pi160 );
  not  g05071 ( new_n5448 , new_n4927 );
  nor  g05072 ( new_n5449 , new_n5448 , new_n4938 );
  xor  g05073 ( new_n5450 , new_n5410 , new_n5411 );
  nand g05074 ( new_n5451 , pi160 , pi180 );
  xnor g05075 ( new_n5452 , new_n5450 , new_n5451 );
  nand g05076 ( new_n5453 , new_n4933 , new_n4936 );
  nand g05077 ( new_n5454 , new_n4932 , new_n4937 );
  nand g05078 ( new_n5455 , new_n5453 , new_n5454 );
  xor  g05079 ( new_n5456 , new_n5452 , new_n5455 );
  nand g05080 ( new_n5457 , new_n5449 , new_n5456 );
  nand g05081 ( new_n5458 , new_n5447 , new_n5457 );
  xor  g05082 ( new_n5459 , new_n5405 , new_n5413 );
  nor  g05083 ( new_n5460 , new_n5450 , new_n5451 );
  nor  g05084 ( new_n5461 , new_n5452 , new_n5455 );
  nor  g05085 ( new_n5462 , new_n5460 , new_n5461 );
  xor  g05086 ( new_n5463 , new_n5459 , new_n5462 );
  xor  g05087 ( new_n5464 , new_n5447 , new_n5457 );
  nand g05088 ( new_n5465 , new_n5463 , new_n5464 );
  nand g05089 ( new_n5466 , new_n5458 , new_n5465 );
  nand g05090 ( new_n5467 , new_n5446 , new_n5466 );
  not  g05091 ( new_n5468 , new_n5462 );
  nand g05092 ( new_n5469 , new_n5459 , new_n5468 );
  xor  g05093 ( new_n5470 , new_n5446 , new_n5466 );
  nand g05094 ( new_n5471 , new_n5469 , new_n5470 );
  nand g05095 ( new_n5472 , new_n5467 , new_n5471 );
  xor  g05096 ( new_n5473 , new_n5445 , new_n5472 );
  xor  g05097 ( new_n5474 , new_n5442 , new_n5473 );
  nand g05098 ( new_n5475 , pi038 , pi219 );
  nand g05099 ( new_n5476 , pi038 , pi087 );
  nand g05100 ( new_n5477 , pi113 , pi219 );
  nand g05101 ( new_n5478 , new_n5476 , new_n5477 );
  nand g05102 ( new_n5479 , pi102 , pi118 );
  xor  g05103 ( new_n5480 , new_n5476 , new_n5477 );
  nand g05104 ( new_n5481 , new_n5479 , new_n5480 );
  nand g05105 ( new_n5482 , new_n5478 , new_n5481 );
  xor  g05106 ( new_n5483 , new_n5479 , new_n5480 );
  nand g05107 ( new_n5484 , pi001 , pi108 );
  nand g05108 ( new_n5485 , pi042 , pi122 );
  nand g05109 ( new_n5486 , pi051 , pi135 );
  nand g05110 ( new_n5487 , new_n5485 , new_n5486 );
  nand g05111 ( new_n5488 , new_n5371 , new_n5487 );
  nand g05112 ( new_n5489 , new_n5484 , new_n5488 );
  xor  g05113 ( new_n5490 , new_n5484 , new_n5488 );
  nand g05114 ( new_n5491 , pi102 , pi108 );
  nand g05115 ( new_n5492 , pi001 , pi042 );
  nand g05116 ( new_n5493 , new_n5491 , new_n5492 );
  xor  g05117 ( new_n5494 , new_n5491 , new_n5492 );
  nand g05118 ( new_n5495 , new_n5369 , new_n5494 );
  nand g05119 ( new_n5496 , new_n5493 , new_n5495 );
  nand g05120 ( new_n5497 , new_n5490 , new_n5496 );
  nand g05121 ( new_n5498 , new_n5489 , new_n5497 );
  or   g05122 ( new_n5499 , new_n5483 , new_n5498 );
  xor  g05123 ( new_n5500 , new_n5377 , new_n5378 );
  xor  g05124 ( new_n5501 , new_n5483 , new_n5498 );
  nand g05125 ( new_n5502 , new_n5500 , new_n5501 );
  nand g05126 ( new_n5503 , new_n5499 , new_n5502 );
  xor  g05127 ( new_n5504 , new_n5482 , new_n5503 );
  xor  g05128 ( new_n5505 , new_n5469 , new_n5470 );
  xor  g05129 ( new_n5506 , new_n5463 , new_n5464 );
  nand g05130 ( new_n5507 , pi048 , pi182 );
  nand g05131 ( new_n5508 , new_n4891 , new_n4892 );
  nand g05132 ( new_n5509 , new_n4890 , new_n4893 );
  nand g05133 ( new_n5510 , new_n5508 , new_n5509 );
  nand g05134 ( new_n5511 , new_n5507 , new_n5510 );
  nand g05135 ( new_n5512 , pi076 , pi162 );
  nand g05136 ( new_n5513 , pi033 , pi216 );
  nand g05137 ( new_n5514 , pi041 , pi179 );
  xor  g05138 ( new_n5515 , new_n5513 , new_n5514 );
  xor  g05139 ( new_n5516 , new_n5512 , new_n5515 );
  xor  g05140 ( new_n5517 , new_n5507 , new_n5510 );
  nand g05141 ( new_n5518 , new_n5516 , new_n5517 );
  nand g05142 ( new_n5519 , new_n5511 , new_n5518 );
  nand g05143 ( new_n5520 , pi179 , pi216 );
  nand g05144 ( new_n5521 , pi033 , pi076 );
  nand g05145 ( new_n5522 , pi079 , pi162 );
  nand g05146 ( new_n5523 , new_n5521 , new_n5522 );
  nand g05147 ( new_n5524 , pi033 , pi079 );
  or   g05148 ( new_n5525 , new_n5512 , new_n5524 );
  nand g05149 ( new_n5526 , new_n5523 , new_n5525 );
  xor  g05150 ( new_n5527 , new_n5520 , new_n5526 );
  nand g05151 ( new_n5528 , new_n5513 , new_n5514 );
  nand g05152 ( new_n5529 , new_n5512 , new_n5515 );
  nand g05153 ( new_n5530 , new_n5528 , new_n5529 );
  xor  g05154 ( new_n5531 , new_n5527 , new_n5530 );
  nand g05155 ( new_n5532 , pi041 , pi048 );
  nand g05156 ( new_n5533 , pi182 , pi237 );
  nand g05157 ( new_n5534 , new_n5532 , new_n5533 );
  nand g05158 ( new_n5535 , pi041 , pi237 );
  or   g05159 ( new_n5536 , new_n5507 , new_n5535 );
  nand g05160 ( new_n5537 , new_n5534 , new_n5536 );
  xor  g05161 ( new_n5538 , new_n5531 , new_n5537 );
  xnor g05162 ( new_n5539 , new_n5519 , new_n5538 );
  xor  g05163 ( new_n5540 , new_n5516 , new_n5517 );
  nand g05164 ( new_n5541 , pi138 , pi237 );
  nor  g05165 ( new_n5542 , new_n5540 , new_n5541 );
  xnor g05166 ( new_n5543 , new_n5540 , new_n5541 );
  nand g05167 ( new_n5544 , new_n4895 , new_n4898 );
  nand g05168 ( new_n5545 , new_n4894 , new_n4899 );
  nand g05169 ( new_n5546 , new_n5544 , new_n5545 );
  nor  g05170 ( new_n5547 , new_n5543 , new_n5546 );
  nor  g05171 ( new_n5548 , new_n5542 , new_n5547 );
  xor  g05172 ( new_n5549 , new_n5539 , new_n5548 );
  nand g05173 ( new_n5550 , pi138 , pi238 );
  not  g05174 ( new_n5551 , new_n4889 );
  nor  g05175 ( new_n5552 , new_n5551 , new_n4900 );
  xor  g05176 ( new_n5553 , new_n5543 , new_n5546 );
  nand g05177 ( new_n5554 , new_n5552 , new_n5553 );
  xor  g05178 ( new_n5555 , new_n5550 , new_n5554 );
  xor  g05179 ( new_n5556 , new_n5549 , new_n5555 );
  nand g05180 ( new_n5557 , pi061 , pi123 );
  nand g05181 ( new_n5558 , pi099 , pi178 );
  nand g05182 ( new_n5559 , pi023 , pi188 );
  nand g05183 ( new_n5560 , new_n5558 , new_n5559 );
  nand g05184 ( new_n5561 , pi099 , pi188 );
  nand g05185 ( new_n5562 , pi023 , pi178 );
  or   g05186 ( new_n5563 , new_n5561 , new_n5562 );
  nand g05187 ( new_n5564 , new_n5560 , new_n5563 );
  xor  g05188 ( new_n5565 , new_n5557 , new_n5564 );
  nand g05189 ( new_n5566 , pi061 , pi169 );
  nand g05190 ( new_n5567 , new_n5561 , new_n5566 );
  nand g05191 ( new_n5568 , pi123 , pi178 );
  xor  g05192 ( new_n5569 , new_n5561 , new_n5566 );
  nand g05193 ( new_n5570 , new_n5568 , new_n5569 );
  nand g05194 ( new_n5571 , new_n5567 , new_n5570 );
  xor  g05195 ( new_n5572 , new_n5565 , new_n5571 );
  nand g05196 ( new_n5573 , pi012 , pi169 );
  nand g05197 ( new_n5574 , pi071 , pi144 );
  and  g05198 ( new_n5575 , new_n5573 , new_n5574 );
  nand g05199 ( new_n5576 , pi012 , pi071 );
  nand g05200 ( new_n5577 , pi144 , pi169 );
  nor  g05201 ( new_n5578 , new_n5576 , new_n5577 );
  or   g05202 ( new_n5579 , new_n5575 , new_n5578 );
  xnor g05203 ( new_n5580 , new_n5572 , new_n5579 );
  nand g05204 ( new_n5581 , new_n4845 , new_n4846 );
  nand g05205 ( new_n5582 , new_n4844 , new_n4847 );
  nand g05206 ( new_n5583 , new_n5581 , new_n5582 );
  nand g05207 ( new_n5584 , new_n5576 , new_n5583 );
  xor  g05208 ( new_n5585 , new_n5568 , new_n5569 );
  xor  g05209 ( new_n5586 , new_n5576 , new_n5583 );
  nand g05210 ( new_n5587 , new_n5585 , new_n5586 );
  nand g05211 ( new_n5588 , new_n5584 , new_n5587 );
  xor  g05212 ( new_n5589 , new_n5580 , new_n5588 );
  nand g05213 ( new_n5590 , pi142 , pi144 );
  not  g05214 ( new_n5591 , new_n5590 );
  or   g05215 ( new_n5592 , new_n4841 , new_n4842 );
  not  g05216 ( new_n5593 , new_n4848 );
  nand g05217 ( new_n5594 , new_n4843 , new_n5593 );
  nand g05218 ( new_n5595 , new_n5592 , new_n5594 );
  nand g05219 ( new_n5596 , new_n5591 , new_n5595 );
  xor  g05220 ( new_n5597 , new_n5590 , new_n5595 );
  xor  g05221 ( new_n5598 , new_n5585 , new_n5586 );
  or   g05222 ( new_n5599 , new_n5597 , new_n5598 );
  nand g05223 ( new_n5600 , new_n5596 , new_n5599 );
  xor  g05224 ( new_n5601 , new_n5589 , new_n5600 );
  nor  g05225 ( new_n5602 , new_n4849 , new_n4856 );
  xor  g05226 ( new_n5603 , new_n5597 , new_n5598 );
  nand g05227 ( new_n5604 , new_n5602 , new_n5603 );
  nand g05228 ( new_n5605 , pi098 , pi142 );
  xor  g05229 ( new_n5606 , new_n5604 , new_n5605 );
  xor  g05230 ( new_n5607 , new_n5601 , new_n5606 );
  nor  g05231 ( new_n5608 , new_n4826 , new_n4833 );
  xor  g05232 ( new_n5609 , new_n5369 , new_n5494 );
  nand g05233 ( new_n5610 , pi007 , pi219 );
  nand g05234 ( new_n5611 , new_n4822 , new_n4823 );
  nand g05235 ( new_n5612 , new_n4821 , new_n4824 );
  nand g05236 ( new_n5613 , new_n5611 , new_n5612 );
  xor  g05237 ( new_n5614 , new_n5610 , new_n5613 );
  xnor g05238 ( new_n5615 , new_n5609 , new_n5614 );
  nand g05239 ( new_n5616 , pi087 , pi118 );
  or   g05240 ( new_n5617 , new_n4812 , new_n4819 );
  nand g05241 ( new_n5618 , new_n4820 , new_n4825 );
  nand g05242 ( new_n5619 , new_n5617 , new_n5618 );
  xor  g05243 ( new_n5620 , new_n5616 , new_n5619 );
  xnor g05244 ( new_n5621 , new_n5615 , new_n5620 );
  nand g05245 ( new_n5622 , new_n5608 , new_n5621 );
  nand g05246 ( new_n5623 , pi087 , pi113 );
  xor  g05247 ( new_n5624 , new_n5490 , new_n5496 );
  nand g05248 ( new_n5625 , pi118 , pi219 );
  nand g05249 ( new_n5626 , pi007 , pi102 );
  and  g05250 ( new_n5627 , new_n5625 , new_n5626 );
  nor  g05251 ( new_n5628 , new_n5479 , new_n5610 );
  or   g05252 ( new_n5629 , new_n5627 , new_n5628 );
  xnor g05253 ( new_n5630 , new_n5624 , new_n5629 );
  nand g05254 ( new_n5631 , new_n5610 , new_n5613 );
  nand g05255 ( new_n5632 , new_n5609 , new_n5614 );
  nand g05256 ( new_n5633 , new_n5631 , new_n5632 );
  xnor g05257 ( new_n5634 , new_n5630 , new_n5633 );
  not  g05258 ( new_n5635 , new_n5616 );
  nor  g05259 ( new_n5636 , new_n5635 , new_n5619 );
  nor  g05260 ( new_n5637 , new_n5615 , new_n5620 );
  nor  g05261 ( new_n5638 , new_n5636 , new_n5637 );
  xor  g05262 ( new_n5639 , new_n5634 , new_n5638 );
  xor  g05263 ( new_n5640 , new_n5623 , new_n5639 );
  not  g05264 ( new_n5641 , new_n5640 );
  xor  g05265 ( new_n5642 , new_n5622 , new_n5641 );
  xor  g05266 ( new_n5643 , new_n5607 , new_n5642 );
  xor  g05267 ( new_n5644 , new_n5608 , new_n5621 );
  xor  g05268 ( new_n5645 , new_n5602 , new_n5603 );
  nor  g05269 ( new_n5646 , new_n5644 , new_n5645 );
  xnor g05270 ( new_n5647 , new_n5644 , new_n5645 );
  nand g05271 ( new_n5648 , new_n4834 , new_n4857 );
  nand g05272 ( new_n5649 , new_n4858 , new_n4878 );
  nand g05273 ( new_n5650 , new_n5648 , new_n5649 );
  nor  g05274 ( new_n5651 , new_n5647 , new_n5650 );
  nor  g05275 ( new_n5652 , new_n5646 , new_n5651 );
  xor  g05276 ( new_n5653 , new_n5643 , new_n5652 );
  xnor g05277 ( new_n5654 , new_n5552 , new_n5553 );
  nand g05278 ( new_n5655 , new_n4901 , new_n4917 );
  not  g05279 ( new_n5656 , new_n4879 );
  nand g05280 ( new_n5657 , new_n5656 , new_n4918 );
  nand g05281 ( new_n5658 , new_n5655 , new_n5657 );
  or   g05282 ( new_n5659 , new_n5654 , new_n5658 );
  xnor g05283 ( new_n5660 , new_n5647 , new_n5650 );
  xor  g05284 ( new_n5661 , new_n5654 , new_n5658 );
  nand g05285 ( new_n5662 , new_n5660 , new_n5661 );
  nand g05286 ( new_n5663 , new_n5659 , new_n5662 );
  xor  g05287 ( new_n5664 , new_n5653 , new_n5663 );
  xor  g05288 ( new_n5665 , new_n5556 , new_n5664 );
  nand g05289 ( new_n5666 , new_n5506 , new_n5665 );
  xor  g05290 ( new_n5667 , new_n5506 , new_n5665 );
  xor  g05291 ( new_n5668 , new_n5449 , new_n5456 );
  or   g05292 ( new_n5669 , new_n4939 , new_n4957 );
  nand g05293 ( new_n5670 , new_n4919 , new_n4958 );
  nand g05294 ( new_n5671 , new_n5669 , new_n5670 );
  or   g05295 ( new_n5672 , new_n5668 , new_n5671 );
  xor  g05296 ( new_n5673 , new_n5660 , new_n5661 );
  not  g05297 ( new_n5674 , new_n5673 );
  xor  g05298 ( new_n5675 , new_n5668 , new_n5671 );
  nand g05299 ( new_n5676 , new_n5674 , new_n5675 );
  nand g05300 ( new_n5677 , new_n5672 , new_n5676 );
  nand g05301 ( new_n5678 , new_n5667 , new_n5677 );
  nand g05302 ( new_n5679 , new_n5666 , new_n5678 );
  nand g05303 ( new_n5680 , new_n5505 , new_n5679 );
  not  g05304 ( new_n5681 , new_n5638 );
  nor  g05305 ( new_n5682 , new_n5634 , new_n5681 );
  xor  g05306 ( new_n5683 , new_n5500 , new_n5501 );
  not  g05307 ( new_n5684 , new_n5683 );
  nor  g05308 ( new_n5685 , new_n5624 , new_n5629 );
  nor  g05309 ( new_n5686 , new_n5630 , new_n5633 );
  xor  g05310 ( new_n5687 , new_n5628 , new_n5686 );
  nor  g05311 ( new_n5688 , new_n5685 , new_n5687 );
  xor  g05312 ( new_n5689 , new_n5684 , new_n5688 );
  xor  g05313 ( new_n5690 , new_n5682 , new_n5689 );
  nor  g05314 ( new_n5691 , new_n5623 , new_n5639 );
  nor  g05315 ( new_n5692 , new_n5622 , new_n5641 );
  or   g05316 ( new_n5693 , new_n5691 , new_n5692 );
  xnor g05317 ( new_n5694 , new_n5690 , new_n5693 );
  nand g05318 ( new_n5695 , new_n5604 , new_n5605 );
  not  g05319 ( new_n5696 , new_n5601 );
  nand g05320 ( new_n5697 , new_n5696 , new_n5606 );
  nand g05321 ( new_n5698 , new_n5695 , new_n5697 );
  nand g05322 ( new_n5699 , new_n5589 , new_n5600 );
  nand g05323 ( new_n5700 , pi061 , pi099 );
  nand g05324 ( new_n5701 , pi155 , pi188 );
  xor  g05325 ( new_n5702 , new_n5700 , new_n5701 );
  xor  g05326 ( new_n5703 , new_n5562 , new_n5702 );
  not  g05327 ( new_n5704 , new_n5703 );
  nand g05328 ( new_n5705 , pi012 , pi123 );
  xor  g05329 ( new_n5706 , new_n5563 , new_n5705 );
  xor  g05330 ( new_n5707 , new_n5704 , new_n5706 );
  nand g05331 ( new_n5708 , pi071 , pi098 );
  nand g05332 ( new_n5709 , pi043 , pi142 );
  xor  g05333 ( new_n5710 , new_n5708 , new_n5709 );
  xor  g05334 ( new_n5711 , new_n5577 , new_n5710 );
  nand g05335 ( new_n5712 , new_n5557 , new_n5564 );
  nand g05336 ( new_n5713 , new_n5565 , new_n5571 );
  nand g05337 ( new_n5714 , new_n5712 , new_n5713 );
  xor  g05338 ( new_n5715 , new_n5711 , new_n5714 );
  xor  g05339 ( new_n5716 , new_n5707 , new_n5715 );
  nor  g05340 ( new_n5717 , new_n5572 , new_n5579 );
  nor  g05341 ( new_n5718 , new_n5580 , new_n5588 );
  xor  g05342 ( new_n5719 , new_n5578 , new_n5718 );
  nor  g05343 ( new_n5720 , new_n5717 , new_n5719 );
  xor  g05344 ( new_n5721 , new_n5716 , new_n5720 );
  xor  g05345 ( new_n5722 , new_n5699 , new_n5721 );
  xor  g05346 ( new_n5723 , new_n5698 , new_n5722 );
  xnor g05347 ( new_n5724 , new_n5694 , new_n5723 );
  nand g05348 ( new_n5725 , new_n5607 , new_n5642 );
  nand g05349 ( new_n5726 , new_n5643 , new_n5652 );
  nand g05350 ( new_n5727 , new_n5725 , new_n5726 );
  xor  g05351 ( new_n5728 , new_n5724 , new_n5727 );
  not  g05352 ( new_n5729 , new_n5548 );
  nand g05353 ( new_n5730 , new_n5539 , new_n5729 );
  nand g05354 ( new_n5731 , pi162 , pi251 );
  nand g05355 ( new_n5732 , pi076 , pi179 );
  xor  g05356 ( new_n5733 , new_n5731 , new_n5732 );
  xor  g05357 ( new_n5734 , new_n5524 , new_n5733 );
  not  g05358 ( new_n5735 , new_n5734 );
  nand g05359 ( new_n5736 , pi048 , pi216 );
  xor  g05360 ( new_n5737 , new_n5525 , new_n5736 );
  xor  g05361 ( new_n5738 , new_n5735 , new_n5737 );
  nand g05362 ( new_n5739 , pi182 , pi238 );
  nand g05363 ( new_n5740 , pi138 , pi193 );
  xor  g05364 ( new_n5741 , new_n5739 , new_n5740 );
  xor  g05365 ( new_n5742 , new_n5535 , new_n5741 );
  nand g05366 ( new_n5743 , new_n5520 , new_n5526 );
  nand g05367 ( new_n5744 , new_n5527 , new_n5530 );
  nand g05368 ( new_n5745 , new_n5743 , new_n5744 );
  xor  g05369 ( new_n5746 , new_n5742 , new_n5745 );
  xor  g05370 ( new_n5747 , new_n5738 , new_n5746 );
  nand g05371 ( new_n5748 , new_n5531 , new_n5537 );
  nand g05372 ( new_n5749 , new_n5519 , new_n5538 );
  nand g05373 ( new_n5750 , new_n5748 , new_n5749 );
  xor  g05374 ( new_n5751 , new_n5536 , new_n5750 );
  xnor g05375 ( new_n5752 , new_n5747 , new_n5751 );
  xnor g05376 ( new_n5753 , new_n5730 , new_n5752 );
  nand g05377 ( new_n5754 , new_n5550 , new_n5554 );
  nand g05378 ( new_n5755 , new_n5549 , new_n5555 );
  nand g05379 ( new_n5756 , new_n5754 , new_n5755 );
  xor  g05380 ( new_n5757 , new_n5753 , new_n5756 );
  xor  g05381 ( new_n5758 , new_n5728 , new_n5757 );
  or   g05382 ( new_n5759 , new_n5653 , new_n5663 );
  nand g05383 ( new_n5760 , new_n5556 , new_n5664 );
  nand g05384 ( new_n5761 , new_n5759 , new_n5760 );
  xor  g05385 ( new_n5762 , new_n5758 , new_n5761 );
  not  g05386 ( new_n5763 , new_n5762 );
  xor  g05387 ( new_n5764 , new_n5505 , new_n5679 );
  nand g05388 ( new_n5765 , new_n5763 , new_n5764 );
  nand g05389 ( new_n5766 , new_n5680 , new_n5765 );
  xor  g05390 ( new_n5767 , new_n5504 , new_n5766 );
  xor  g05391 ( new_n5768 , new_n5475 , new_n5767 );
  xor  g05392 ( new_n5769 , new_n5474 , new_n5768 );
  xor  g05393 ( new_n5770 , new_n5381 , new_n5769 );
  xor  g05394 ( new_n5771 , new_n5366 , new_n5770 );
  nand g05395 ( new_n5772 , new_n5628 , new_n5686 );
  or   g05396 ( new_n5773 , new_n5684 , new_n5688 );
  nand g05397 ( new_n5774 , new_n5772 , new_n5773 );
  nand g05398 ( new_n5775 , pi042 , pi059 );
  nand g05399 ( new_n5776 , pi108 , pi135 );
  xor  g05400 ( new_n5777 , new_n5775 , new_n5776 );
  xor  g05401 ( new_n5778 , new_n5774 , new_n5777 );
  nand g05402 ( new_n5779 , new_n5682 , new_n5689 );
  nand g05403 ( new_n5780 , new_n5690 , new_n5693 );
  nand g05404 ( new_n5781 , new_n5779 , new_n5780 );
  nand g05405 ( new_n5782 , pi051 , pi094 );
  xor  g05406 ( new_n5783 , new_n5781 , new_n5782 );
  xor  g05407 ( new_n5784 , new_n5778 , new_n5783 );
  nand g05408 ( new_n5785 , pi007 , pi122 );
  nand g05409 ( new_n5786 , pi001 , pi118 );
  xor  g05410 ( new_n5787 , new_n5785 , new_n5786 );
  nand g05411 ( new_n5788 , new_n5711 , new_n5714 );
  not  g05412 ( new_n5789 , new_n5707 );
  nand g05413 ( new_n5790 , new_n5789 , new_n5715 );
  nand g05414 ( new_n5791 , new_n5788 , new_n5790 );
  nand g05415 ( new_n5792 , pi123 , pi144 );
  nand g05416 ( new_n5793 , pi043 , pi071 );
  nand g05417 ( new_n5794 , pi098 , pi169 );
  xnor g05418 ( new_n5795 , new_n5793 , new_n5794 );
  xor  g05419 ( new_n5796 , new_n5792 , new_n5795 );
  xor  g05420 ( new_n5797 , new_n5791 , new_n5796 );
  nand g05421 ( new_n5798 , new_n5708 , new_n5709 );
  nand g05422 ( new_n5799 , new_n5577 , new_n5710 );
  nand g05423 ( new_n5800 , new_n5798 , new_n5799 );
  or   g05424 ( new_n5801 , new_n5563 , new_n5705 );
  nand g05425 ( new_n5802 , new_n5704 , new_n5706 );
  nand g05426 ( new_n5803 , new_n5801 , new_n5802 );
  xor  g05427 ( new_n5804 , new_n5800 , new_n5803 );
  nand g05428 ( new_n5805 , new_n5700 , new_n5701 );
  nand g05429 ( new_n5806 , new_n5562 , new_n5702 );
  nand g05430 ( new_n5807 , new_n5805 , new_n5806 );
  nand g05431 ( new_n5808 , pi012 , pi099 );
  xor  g05432 ( new_n5809 , new_n5807 , new_n5808 );
  xor  g05433 ( new_n5810 , new_n5804 , new_n5809 );
  xor  g05434 ( new_n5811 , new_n5797 , new_n5810 );
  xor  g05435 ( new_n5812 , new_n5787 , new_n5811 );
  xor  g05436 ( new_n5813 , new_n5784 , new_n5812 );
  xor  g05437 ( new_n5814 , new_n5771 , new_n5813 );
  nand g05438 ( new_n5815 , new_n5739 , new_n5740 );
  nand g05439 ( new_n5816 , new_n5535 , new_n5741 );
  nand g05440 ( new_n5817 , new_n5815 , new_n5816 );
  nand g05441 ( new_n5818 , pi216 , pi237 );
  nand g05442 ( new_n5819 , pi041 , pi238 );
  xor  g05443 ( new_n5820 , new_n5818 , new_n5819 );
  xor  g05444 ( new_n5821 , new_n5817 , new_n5820 );
  xor  g05445 ( new_n5822 , new_n5814 , new_n5821 );
  nand g05446 ( new_n5823 , new_n5699 , new_n5721 );
  nand g05447 ( new_n5824 , new_n5698 , new_n5722 );
  nand g05448 ( new_n5825 , new_n5823 , new_n5824 );
  nand g05449 ( new_n5826 , new_n5578 , new_n5718 );
  not  g05450 ( new_n5827 , new_n5720 );
  nand g05451 ( new_n5828 , new_n5716 , new_n5827 );
  nand g05452 ( new_n5829 , new_n5826 , new_n5828 );
  xor  g05453 ( new_n5830 , new_n5825 , new_n5829 );
  or   g05454 ( new_n5831 , new_n5525 , new_n5736 );
  nand g05455 ( new_n5832 , new_n5735 , new_n5737 );
  nand g05456 ( new_n5833 , new_n5831 , new_n5832 );
  nand g05457 ( new_n5834 , new_n5742 , new_n5745 );
  not  g05458 ( new_n5835 , new_n5738 );
  nand g05459 ( new_n5836 , new_n5835 , new_n5746 );
  nand g05460 ( new_n5837 , new_n5834 , new_n5836 );
  xor  g05461 ( new_n5838 , new_n5833 , new_n5837 );
  xor  g05462 ( new_n5839 , new_n5830 , new_n5838 );
  not  g05463 ( new_n5840 , new_n5757 );
  nor  g05464 ( new_n5841 , new_n5728 , new_n5840 );
  nor  g05465 ( new_n5842 , new_n5758 , new_n5761 );
  nor  g05466 ( new_n5843 , new_n5841 , new_n5842 );
  nor  g05467 ( new_n5844 , new_n5391 , new_n5420 );
  nor  g05468 ( new_n5845 , new_n5419 , new_n5422 );
  or   g05469 ( new_n5846 , new_n5844 , new_n5845 );
  nand g05470 ( new_n5847 , pi057 , pi177 );
  nand g05471 ( new_n5848 , pi194 , pi225 );
  xor  g05472 ( new_n5849 , new_n5847 , new_n5848 );
  xor  g05473 ( new_n5850 , new_n5846 , new_n5849 );
  xor  g05474 ( new_n5851 , new_n5843 , new_n5850 );
  nand g05475 ( new_n5852 , new_n5424 , new_n5425 );
  nand g05476 ( new_n5853 , new_n5382 , new_n5426 );
  nand g05477 ( new_n5854 , new_n5852 , new_n5853 );
  or   g05478 ( new_n5855 , new_n5427 , new_n5430 );
  nand g05479 ( new_n5856 , new_n5423 , new_n5431 );
  nand g05480 ( new_n5857 , new_n5855 , new_n5856 );
  xor  g05481 ( new_n5858 , new_n5854 , new_n5857 );
  nand g05482 ( new_n5859 , pi020 , pi068 );
  nand g05483 ( new_n5860 , pi085 , pi101 );
  xor  g05484 ( new_n5861 , new_n5859 , new_n5860 );
  xor  g05485 ( new_n5862 , new_n5858 , new_n5861 );
  nor  g05486 ( new_n5863 , new_n5730 , new_n5752 );
  nor  g05487 ( new_n5864 , new_n5753 , new_n5756 );
  nor  g05488 ( new_n5865 , new_n5863 , new_n5864 );
  nand g05489 ( new_n5866 , new_n5416 , new_n5417 );
  nand g05490 ( new_n5867 , new_n5390 , new_n5418 );
  nand g05491 ( new_n5868 , new_n5866 , new_n5867 );
  nand g05492 ( new_n5869 , pi180 , pi223 );
  xor  g05493 ( new_n5870 , new_n5868 , new_n5869 );
  xor  g05494 ( new_n5871 , new_n5865 , new_n5870 );
  xor  g05495 ( new_n5872 , new_n5862 , new_n5871 );
  nand g05496 ( new_n5873 , pi036 , pi060 );
  nand g05497 ( new_n5874 , pi138 , pi159 );
  nand g05498 ( new_n5875 , pi033 , pi251 );
  nand g05499 ( new_n5876 , pi162 , pi192 );
  or   g05500 ( new_n5877 , new_n5536 , new_n5750 );
  nand g05501 ( new_n5878 , new_n5747 , new_n5751 );
  nand g05502 ( new_n5879 , new_n5877 , new_n5878 );
  xor  g05503 ( new_n5880 , new_n5876 , new_n5879 );
  xor  g05504 ( new_n5881 , new_n5875 , new_n5880 );
  xor  g05505 ( new_n5882 , new_n5874 , new_n5881 );
  xor  g05506 ( new_n5883 , new_n5873 , new_n5882 );
  xor  g05507 ( new_n5884 , new_n5872 , new_n5883 );
  xor  g05508 ( new_n5885 , new_n5851 , new_n5884 );
  nand g05509 ( new_n5886 , pi048 , pi076 );
  nand g05510 ( new_n5887 , pi182 , pi193 );
  nand g05511 ( new_n5888 , new_n5731 , new_n5732 );
  nand g05512 ( new_n5889 , new_n5524 , new_n5733 );
  nand g05513 ( new_n5890 , new_n5888 , new_n5889 );
  xor  g05514 ( new_n5891 , new_n5887 , new_n5890 );
  xor  g05515 ( new_n5892 , new_n5886 , new_n5891 );
  xor  g05516 ( new_n5893 , new_n5885 , new_n5892 );
  xor  g05517 ( new_n5894 , new_n5839 , new_n5893 );
  nand g05518 ( new_n5895 , pi079 , pi179 );
  nand g05519 ( new_n5896 , pi086 , pi188 );
  nand g05520 ( new_n5897 , pi023 , pi061 );
  nand g05521 ( new_n5898 , pi155 , pi178 );
  xor  g05522 ( new_n5899 , new_n5897 , new_n5898 );
  nand g05523 ( new_n5900 , pi126 , pi142 );
  nand g05524 ( new_n5901 , new_n5694 , new_n5723 );
  or   g05525 ( new_n5902 , new_n5724 , new_n5727 );
  nand g05526 ( new_n5903 , new_n5901 , new_n5902 );
  xor  g05527 ( new_n5904 , new_n5900 , new_n5903 );
  xor  g05528 ( new_n5905 , new_n5899 , new_n5904 );
  xor  g05529 ( new_n5906 , new_n5896 , new_n5905 );
  xor  g05530 ( new_n5907 , new_n5895 , new_n5906 );
  xor  g05531 ( new_n5908 , new_n5894 , new_n5907 );
  xor  g05532 ( po021 , new_n5822 , new_n5908 );
  xor  g05533 ( po022 , new_n4799 , new_n4806 );
  xor  g05534 ( po023 , new_n2539 , new_n2575 );
  xor  g05535 ( po024 , new_n1813 , new_n1815 );
  xnor g05536 ( po025 , new_n3691 , new_n3692 );
  xor  g05537 ( po026 , new_n5360 , new_n5361 );
  nand g05538 ( new_n5915 , pi089 , pi141 );
  nand g05539 ( new_n5916 , new_n3334 , new_n3335 );
  nand g05540 ( new_n5917 , new_n3333 , new_n3336 );
  nand g05541 ( new_n5918 , new_n5916 , new_n5917 );
  xor  g05542 ( new_n5919 , new_n5915 , new_n5918 );
  nand g05543 ( new_n5920 , pi047 , pi254 );
  nand g05544 ( new_n5921 , pi090 , pi158 );
  nand g05545 ( new_n5922 , new_n5920 , new_n5921 );
  nand g05546 ( new_n5923 , pi047 , pi158 );
  nor  g05547 ( new_n5924 , new_n3335 , new_n5923 );
  not  g05548 ( new_n5925 , new_n5924 );
  nand g05549 ( new_n5926 , new_n5922 , new_n5925 );
  xor  g05550 ( new_n5927 , new_n5919 , new_n5926 );
  nand g05551 ( new_n5928 , new_n3338 , new_n3341 );
  nand g05552 ( new_n5929 , new_n3337 , new_n3342 );
  nand g05553 ( new_n5930 , new_n5928 , new_n5929 );
  nand g05554 ( new_n5931 , pi154 , pi161 );
  nand g05555 ( new_n5932 , pi095 , pi241 );
  nand g05556 ( new_n5933 , new_n5931 , new_n5932 );
  nand g05557 ( new_n5934 , pi095 , pi161 );
  or   g05558 ( new_n5935 , new_n3338 , new_n5934 );
  nand g05559 ( new_n5936 , new_n5933 , new_n5935 );
  xor  g05560 ( new_n5937 , new_n5930 , new_n5936 );
  xor  g05561 ( new_n5938 , new_n5927 , new_n5937 );
  not  g05562 ( new_n5939 , new_n5938 );
  not  g05563 ( new_n5940 , new_n3344 );
  nand g05564 ( new_n5941 , new_n5940 , new_n3347 );
  or   g05565 ( new_n5942 , new_n3343 , new_n3348 );
  nand g05566 ( new_n5943 , new_n5941 , new_n5942 );
  nand g05567 ( new_n5944 , new_n5939 , new_n5943 );
  nand g05568 ( new_n5945 , pi089 , pi090 );
  nand g05569 ( new_n5946 , pi018 , pi254 );
  xor  g05570 ( new_n5947 , new_n5945 , new_n5946 );
  xor  g05571 ( new_n5948 , new_n5923 , new_n5947 );
  nand g05572 ( new_n5949 , pi141 , pi154 );
  xor  g05573 ( new_n5950 , new_n5925 , new_n5949 );
  not  g05574 ( new_n5951 , new_n5950 );
  xor  g05575 ( new_n5952 , new_n5948 , new_n5951 );
  nand g05576 ( new_n5953 , pi006 , pi241 );
  nand g05577 ( new_n5954 , pi209 , pi236 );
  xor  g05578 ( new_n5955 , new_n5953 , new_n5954 );
  xor  g05579 ( new_n5956 , new_n5934 , new_n5955 );
  nand g05580 ( new_n5957 , new_n5915 , new_n5918 );
  nand g05581 ( new_n5958 , new_n5919 , new_n5926 );
  nand g05582 ( new_n5959 , new_n5957 , new_n5958 );
  xor  g05583 ( new_n5960 , new_n5956 , new_n5959 );
  xor  g05584 ( new_n5961 , new_n5952 , new_n5960 );
  nand g05585 ( new_n5962 , new_n5930 , new_n5936 );
  nand g05586 ( new_n5963 , new_n5927 , new_n5937 );
  nand g05587 ( new_n5964 , new_n5962 , new_n5963 );
  xor  g05588 ( new_n5965 , new_n5935 , new_n5964 );
  xnor g05589 ( new_n5966 , new_n5961 , new_n5965 );
  or   g05590 ( new_n5967 , new_n5944 , new_n5966 );
  xor  g05591 ( new_n5968 , new_n5944 , new_n5966 );
  nand g05592 ( new_n5969 , pi006 , pi236 );
  xor  g05593 ( new_n5970 , new_n5938 , new_n5943 );
  nor  g05594 ( new_n5971 , new_n5969 , new_n5970 );
  nand g05595 ( new_n5972 , new_n3332 , new_n3349 );
  xor  g05596 ( new_n5973 , new_n5969 , new_n5970 );
  not  g05597 ( new_n5974 , new_n5973 );
  nor  g05598 ( new_n5975 , new_n5972 , new_n5974 );
  or   g05599 ( new_n5976 , new_n5971 , new_n5975 );
  nand g05600 ( new_n5977 , new_n5968 , new_n5976 );
  nand g05601 ( new_n5978 , new_n5967 , new_n5977 );
  nand g05602 ( new_n5979 , pi133 , pi229 );
  nand g05603 ( new_n5980 , new_n3469 , new_n3470 );
  nand g05604 ( new_n5981 , new_n3468 , new_n3471 );
  nand g05605 ( new_n5982 , new_n5980 , new_n5981 );
  xor  g05606 ( new_n5983 , new_n5979 , new_n5982 );
  nand g05607 ( new_n5984 , pi092 , pi189 );
  nand g05608 ( new_n5985 , pi064 , pi190 );
  nand g05609 ( new_n5986 , new_n5984 , new_n5985 );
  nand g05610 ( new_n5987 , pi064 , pi092 );
  or   g05611 ( new_n5988 , new_n3470 , new_n5987 );
  nand g05612 ( new_n5989 , new_n5986 , new_n5988 );
  xor  g05613 ( new_n5990 , new_n5983 , new_n5989 );
  nand g05614 ( new_n5991 , pi067 , pi077 );
  nand g05615 ( new_n5992 , pi052 , pi053 );
  and  g05616 ( new_n5993 , new_n5991 , new_n5992 );
  nand g05617 ( new_n5994 , pi053 , pi077 );
  nor  g05618 ( new_n5995 , new_n3473 , new_n5994 );
  or   g05619 ( new_n5996 , new_n5993 , new_n5995 );
  xnor g05620 ( new_n5997 , new_n5990 , new_n5996 );
  nand g05621 ( new_n5998 , new_n3473 , new_n3476 );
  nand g05622 ( new_n5999 , new_n3472 , new_n3477 );
  nand g05623 ( new_n6000 , new_n5998 , new_n5999 );
  xor  g05624 ( new_n6001 , new_n5997 , new_n6000 );
  not  g05625 ( new_n6002 , new_n3479 );
  nand g05626 ( new_n6003 , new_n6002 , new_n3482 );
  or   g05627 ( new_n6004 , new_n3478 , new_n3483 );
  nand g05628 ( new_n6005 , new_n6003 , new_n6004 );
  nand g05629 ( new_n6006 , new_n6001 , new_n6005 );
  nand g05630 ( new_n6007 , pi189 , pi229 );
  nand g05631 ( new_n6008 , pi084 , pi190 );
  xor  g05632 ( new_n6009 , new_n6007 , new_n6008 );
  xor  g05633 ( new_n6010 , new_n5987 , new_n6009 );
  nand g05634 ( new_n6011 , pi067 , pi133 );
  xor  g05635 ( new_n6012 , new_n5988 , new_n6011 );
  xor  g05636 ( new_n6013 , new_n6010 , new_n6012 );
  nand g05637 ( new_n6014 , pi052 , pi185 );
  nand g05638 ( new_n6015 , pi030 , pi131 );
  xor  g05639 ( new_n6016 , new_n5994 , new_n6015 );
  xor  g05640 ( new_n6017 , new_n6014 , new_n6016 );
  nand g05641 ( new_n6018 , new_n5979 , new_n5982 );
  nand g05642 ( new_n6019 , new_n5983 , new_n5989 );
  nand g05643 ( new_n6020 , new_n6018 , new_n6019 );
  xor  g05644 ( new_n6021 , new_n6017 , new_n6020 );
  xnor g05645 ( new_n6022 , new_n6013 , new_n6021 );
  nor  g05646 ( new_n6023 , new_n5990 , new_n5996 );
  nor  g05647 ( new_n6024 , new_n5997 , new_n6000 );
  xor  g05648 ( new_n6025 , new_n5995 , new_n6024 );
  nor  g05649 ( new_n6026 , new_n6023 , new_n6025 );
  xor  g05650 ( new_n6027 , new_n6022 , new_n6026 );
  xnor g05651 ( new_n6028 , new_n6006 , new_n6027 );
  nand g05652 ( new_n6029 , new_n3467 , new_n3484 );
  nand g05653 ( new_n6030 , pi131 , pi185 );
  nand g05654 ( new_n6031 , new_n6029 , new_n6030 );
  xnor g05655 ( new_n6032 , new_n6001 , new_n6005 );
  xor  g05656 ( new_n6033 , new_n6029 , new_n6030 );
  nand g05657 ( new_n6034 , new_n6032 , new_n6033 );
  nand g05658 ( new_n6035 , new_n6031 , new_n6034 );
  xor  g05659 ( new_n6036 , new_n6028 , new_n6035 );
  nand g05660 ( new_n6037 , pi013 , pi073 );
  nand g05661 ( new_n6038 , pi004 , pi112 );
  nand g05662 ( new_n6039 , pi105 , pi170 );
  nand g05663 ( new_n6040 , new_n6038 , new_n6039 );
  nand g05664 ( new_n6041 , pi004 , pi105 );
  or   g05665 ( new_n6042 , new_n3295 , new_n6041 );
  nand g05666 ( new_n6043 , new_n6040 , new_n6042 );
  xor  g05667 ( new_n6044 , new_n6037 , new_n6043 );
  nand g05668 ( new_n6045 , new_n3295 , new_n3296 );
  nand g05669 ( new_n6046 , new_n3294 , new_n3297 );
  nand g05670 ( new_n6047 , new_n6045 , new_n6046 );
  xor  g05671 ( new_n6048 , new_n6044 , new_n6047 );
  nand g05672 ( new_n6049 , pi130 , pi212 );
  nand g05673 ( new_n6050 , pi003 , pi104 );
  nand g05674 ( new_n6051 , new_n6049 , new_n6050 );
  nand g05675 ( new_n6052 , pi104 , pi130 );
  nor  g05676 ( new_n6053 , new_n3299 , new_n6052 );
  not  g05677 ( new_n6054 , new_n6053 );
  nand g05678 ( new_n6055 , new_n6051 , new_n6054 );
  xnor g05679 ( new_n6056 , new_n6048 , new_n6055 );
  nand g05680 ( new_n6057 , new_n3299 , new_n3302 );
  nand g05681 ( new_n6058 , new_n3298 , new_n3303 );
  nand g05682 ( new_n6059 , new_n6057 , new_n6058 );
  xnor g05683 ( new_n6060 , new_n6056 , new_n6059 );
  not  g05684 ( new_n6061 , new_n3305 );
  nor  g05685 ( new_n6062 , new_n6061 , new_n3309 );
  nor  g05686 ( new_n6063 , new_n3304 , new_n3310 );
  nor  g05687 ( new_n6064 , new_n6062 , new_n6063 );
  not  g05688 ( new_n6065 , new_n6064 );
  nor  g05689 ( new_n6066 , new_n6060 , new_n6065 );
  not  g05690 ( new_n6067 , new_n6066 );
  nand g05691 ( new_n6068 , pi170 , pi183 );
  nand g05692 ( new_n6069 , pi073 , pi112 );
  xor  g05693 ( new_n6070 , new_n6068 , new_n6069 );
  xor  g05694 ( new_n6071 , new_n6041 , new_n6070 );
  nand g05695 ( new_n6072 , pi003 , pi013 );
  xor  g05696 ( new_n6073 , new_n6042 , new_n6072 );
  xor  g05697 ( new_n6074 , new_n6071 , new_n6073 );
  nand g05698 ( new_n6075 , pi213 , pi215 );
  nand g05699 ( new_n6076 , pi124 , pi212 );
  xor  g05700 ( new_n6077 , new_n6052 , new_n6076 );
  xor  g05701 ( new_n6078 , new_n6075 , new_n6077 );
  nand g05702 ( new_n6079 , new_n6037 , new_n6043 );
  nand g05703 ( new_n6080 , new_n6044 , new_n6047 );
  nand g05704 ( new_n6081 , new_n6079 , new_n6080 );
  xor  g05705 ( new_n6082 , new_n6078 , new_n6081 );
  xnor g05706 ( new_n6083 , new_n6074 , new_n6082 );
  nor  g05707 ( new_n6084 , new_n6056 , new_n6059 );
  and  g05708 ( new_n6085 , new_n6053 , new_n6084 );
  or   g05709 ( new_n6086 , new_n6048 , new_n6055 );
  nand g05710 ( new_n6087 , new_n6054 , new_n6086 );
  nor  g05711 ( new_n6088 , new_n6084 , new_n6087 );
  or   g05712 ( new_n6089 , new_n6085 , new_n6088 );
  xor  g05713 ( new_n6090 , new_n6083 , new_n6089 );
  xor  g05714 ( new_n6091 , new_n6067 , new_n6090 );
  nand g05715 ( new_n6092 , pi124 , pi213 );
  xor  g05716 ( new_n6093 , new_n6060 , new_n6064 );
  or   g05717 ( new_n6094 , new_n6092 , new_n6093 );
  not  g05718 ( new_n6095 , new_n3311 );
  nand g05719 ( new_n6096 , new_n3293 , new_n6095 );
  not  g05720 ( new_n6097 , new_n6096 );
  xor  g05721 ( new_n6098 , new_n6092 , new_n6093 );
  nand g05722 ( new_n6099 , new_n6097 , new_n6098 );
  nand g05723 ( new_n6100 , new_n6094 , new_n6099 );
  xor  g05724 ( new_n6101 , new_n6091 , new_n6100 );
  xor  g05725 ( new_n6102 , new_n5972 , new_n5974 );
  xor  g05726 ( new_n6103 , new_n6097 , new_n6098 );
  nand g05727 ( new_n6104 , new_n6102 , new_n6103 );
  not  g05728 ( new_n6105 , new_n6104 );
  xnor g05729 ( new_n6106 , new_n6102 , new_n6103 );
  or   g05730 ( new_n6107 , new_n3350 , new_n3377 );
  nand g05731 ( new_n6108 , new_n3312 , new_n3378 );
  nand g05732 ( new_n6109 , new_n6107 , new_n6108 );
  nor  g05733 ( new_n6110 , new_n6106 , new_n6109 );
  nor  g05734 ( new_n6111 , new_n6105 , new_n6110 );
  not  g05735 ( new_n6112 , new_n6111 );
  xor  g05736 ( new_n6113 , new_n6101 , new_n6112 );
  xor  g05737 ( new_n6114 , new_n5968 , new_n5976 );
  xnor g05738 ( new_n6115 , new_n6113 , new_n6114 );
  nand g05739 ( new_n6116 , new_n3407 , new_n3410 );
  nand g05740 ( new_n6117 , new_n3406 , new_n3411 );
  nand g05741 ( new_n6118 , new_n6116 , new_n6117 );
  nand g05742 ( new_n6119 , pi035 , pi120 );
  nand g05743 ( new_n6120 , new_n3403 , new_n3404 );
  nand g05744 ( new_n6121 , new_n3402 , new_n3405 );
  nand g05745 ( new_n6122 , new_n6120 , new_n6121 );
  xor  g05746 ( new_n6123 , new_n6119 , new_n6122 );
  nand g05747 ( new_n6124 , pi015 , pi062 );
  nand g05748 ( new_n6125 , pi065 , pi204 );
  nand g05749 ( new_n6126 , new_n6124 , new_n6125 );
  nand g05750 ( new_n6127 , pi062 , pi204 );
  nor  g05751 ( new_n6128 , new_n3404 , new_n6127 );
  not  g05752 ( new_n6129 , new_n6128 );
  nand g05753 ( new_n6130 , new_n6126 , new_n6129 );
  xor  g05754 ( new_n6131 , new_n6123 , new_n6130 );
  nand g05755 ( new_n6132 , pi139 , pi172 );
  nand g05756 ( new_n6133 , pi198 , pi208 );
  nand g05757 ( new_n6134 , new_n6132 , new_n6133 );
  nand g05758 ( new_n6135 , pi139 , pi198 );
  or   g05759 ( new_n6136 , new_n3407 , new_n6135 );
  nand g05760 ( new_n6137 , new_n6134 , new_n6136 );
  xor  g05761 ( new_n6138 , new_n6131 , new_n6137 );
  xor  g05762 ( new_n6139 , new_n6118 , new_n6138 );
  not  g05763 ( new_n6140 , new_n6139 );
  not  g05764 ( new_n6141 , new_n3413 );
  nand g05765 ( new_n6142 , new_n6141 , new_n3416 );
  or   g05766 ( new_n6143 , new_n3412 , new_n3417 );
  nand g05767 ( new_n6144 , new_n6142 , new_n6143 );
  nand g05768 ( new_n6145 , new_n6140 , new_n6144 );
  nand g05769 ( new_n6146 , pi015 , pi120 );
  nand g05770 ( new_n6147 , pi065 , pi146 );
  xor  g05771 ( new_n6148 , new_n6146 , new_n6147 );
  xor  g05772 ( new_n6149 , new_n6127 , new_n6148 );
  nand g05773 ( new_n6150 , pi035 , pi172 );
  xor  g05774 ( new_n6151 , new_n6129 , new_n6150 );
  not  g05775 ( new_n6152 , new_n6151 );
  xor  g05776 ( new_n6153 , new_n6149 , new_n6152 );
  nand g05777 ( new_n6154 , pi168 , pi197 );
  nand g05778 ( new_n6155 , pi165 , pi208 );
  xor  g05779 ( new_n6156 , new_n6154 , new_n6155 );
  xor  g05780 ( new_n6157 , new_n6135 , new_n6156 );
  nand g05781 ( new_n6158 , new_n6119 , new_n6122 );
  nand g05782 ( new_n6159 , new_n6123 , new_n6130 );
  nand g05783 ( new_n6160 , new_n6158 , new_n6159 );
  xor  g05784 ( new_n6161 , new_n6157 , new_n6160 );
  xor  g05785 ( new_n6162 , new_n6153 , new_n6161 );
  nand g05786 ( new_n6163 , new_n6131 , new_n6137 );
  nand g05787 ( new_n6164 , new_n6118 , new_n6138 );
  nand g05788 ( new_n6165 , new_n6163 , new_n6164 );
  xor  g05789 ( new_n6166 , new_n6136 , new_n6165 );
  xnor g05790 ( new_n6167 , new_n6162 , new_n6166 );
  xor  g05791 ( new_n6168 , new_n6145 , new_n6167 );
  nand g05792 ( new_n6169 , pi165 , pi168 );
  xor  g05793 ( new_n6170 , new_n6139 , new_n6144 );
  nor  g05794 ( new_n6171 , new_n6169 , new_n6170 );
  nand g05795 ( new_n6172 , new_n3401 , new_n3418 );
  xor  g05796 ( new_n6173 , new_n6169 , new_n6170 );
  not  g05797 ( new_n6174 , new_n6173 );
  nor  g05798 ( new_n6175 , new_n6172 , new_n6174 );
  or   g05799 ( new_n6176 , new_n6171 , new_n6175 );
  xor  g05800 ( new_n6177 , new_n6168 , new_n6176 );
  xor  g05801 ( new_n6178 , new_n6115 , new_n6177 );
  xor  g05802 ( new_n6179 , new_n6106 , new_n6109 );
  xor  g05803 ( new_n6180 , new_n6172 , new_n6174 );
  nand g05804 ( new_n6181 , new_n6179 , new_n6180 );
  or   g05805 ( new_n6182 , new_n3419 , new_n3444 );
  nand g05806 ( new_n6183 , new_n3379 , new_n3445 );
  nand g05807 ( new_n6184 , new_n6182 , new_n6183 );
  xor  g05808 ( new_n6185 , new_n6179 , new_n6180 );
  nand g05809 ( new_n6186 , new_n6184 , new_n6185 );
  nand g05810 ( new_n6187 , new_n6181 , new_n6186 );
  xor  g05811 ( new_n6188 , new_n6178 , new_n6187 );
  not  g05812 ( new_n6189 , new_n6188 );
  nand g05813 ( new_n6190 , new_n6036 , new_n6189 );
  xor  g05814 ( new_n6191 , new_n6036 , new_n6189 );
  not  g05815 ( new_n6192 , new_n6191 );
  xor  g05816 ( new_n6193 , new_n6184 , new_n6185 );
  xor  g05817 ( new_n6194 , new_n6032 , new_n6033 );
  not  g05818 ( new_n6195 , new_n6194 );
  nand g05819 ( new_n6196 , new_n6193 , new_n6195 );
  not  g05820 ( new_n6197 , new_n6196 );
  xor  g05821 ( new_n6198 , new_n6193 , new_n6194 );
  or   g05822 ( new_n6199 , new_n3485 , new_n3510 );
  not  g05823 ( new_n6200 , new_n3446 );
  nand g05824 ( new_n6201 , new_n6200 , new_n3511 );
  nand g05825 ( new_n6202 , new_n6199 , new_n6201 );
  nor  g05826 ( new_n6203 , new_n6198 , new_n6202 );
  nor  g05827 ( new_n6204 , new_n6197 , new_n6203 );
  or   g05828 ( new_n6205 , new_n6192 , new_n6204 );
  nand g05829 ( new_n6206 , new_n6190 , new_n6205 );
  nand g05830 ( new_n6207 , pi015 , pi172 );
  nand g05831 ( new_n6208 , new_n6157 , new_n6160 );
  not  g05832 ( new_n6209 , new_n6153 );
  nand g05833 ( new_n6210 , new_n6209 , new_n6161 );
  nand g05834 ( new_n6211 , new_n6208 , new_n6210 );
  xor  g05835 ( new_n6212 , new_n6207 , new_n6211 );
  xor  g05836 ( new_n6213 , new_n6206 , new_n6212 );
  xor  g05837 ( new_n6214 , new_n5978 , new_n6213 );
  nand g05838 ( new_n6215 , pi090 , pi154 );
  nand g05839 ( new_n6216 , pi095 , pi141 );
  xor  g05840 ( new_n6217 , new_n6215 , new_n6216 );
  or   g05841 ( new_n6218 , new_n6042 , new_n6072 );
  not  g05842 ( new_n6219 , new_n6071 );
  nand g05843 ( new_n6220 , new_n6219 , new_n6073 );
  nand g05844 ( new_n6221 , new_n6218 , new_n6220 );
  nand g05845 ( new_n6222 , new_n6068 , new_n6069 );
  nand g05846 ( new_n6223 , new_n6041 , new_n6070 );
  nand g05847 ( new_n6224 , new_n6222 , new_n6223 );
  xor  g05848 ( new_n6225 , new_n6221 , new_n6224 );
  nand g05849 ( new_n6226 , pi104 , pi124 );
  nand g05850 ( new_n6227 , pi212 , pi215 );
  xor  g05851 ( new_n6228 , new_n6226 , new_n6227 );
  xor  g05852 ( new_n6229 , new_n6225 , new_n6228 );
  nand g05853 ( new_n6230 , pi013 , pi130 );
  nand g05854 ( new_n6231 , new_n6052 , new_n6076 );
  nand g05855 ( new_n6232 , new_n6075 , new_n6077 );
  nand g05856 ( new_n6233 , new_n6231 , new_n6232 );
  xor  g05857 ( new_n6234 , new_n6230 , new_n6233 );
  nand g05858 ( new_n6235 , pi003 , pi112 );
  xor  g05859 ( new_n6236 , new_n6234 , new_n6235 );
  xor  g05860 ( new_n6237 , new_n6229 , new_n6236 );
  xor  g05861 ( new_n6238 , new_n6217 , new_n6237 );
  nand g05862 ( new_n6239 , new_n6078 , new_n6081 );
  nand g05863 ( new_n6240 , new_n6074 , new_n6082 );
  nand g05864 ( new_n6241 , new_n6239 , new_n6240 );
  nand g05865 ( new_n6242 , pi018 , pi158 );
  xor  g05866 ( new_n6243 , new_n6241 , new_n6242 );
  xor  g05867 ( new_n6244 , new_n6238 , new_n6243 );
  or   g05868 ( new_n6245 , new_n5935 , new_n5964 );
  nand g05869 ( new_n6246 , new_n5961 , new_n5965 );
  nand g05870 ( new_n6247 , new_n6245 , new_n6246 );
  nand g05871 ( new_n6248 , pi153 , pi236 );
  xor  g05872 ( new_n6249 , new_n6247 , new_n6248 );
  xor  g05873 ( new_n6250 , new_n6244 , new_n6249 );
  nor  g05874 ( new_n6251 , new_n6006 , new_n6027 );
  nor  g05875 ( new_n6252 , new_n6028 , new_n6035 );
  nor  g05876 ( new_n6253 , new_n6251 , new_n6252 );
  nand g05877 ( new_n6254 , pi006 , pi161 );
  nor  g05878 ( new_n6255 , new_n5925 , new_n5949 );
  nor  g05879 ( new_n6256 , new_n5948 , new_n5951 );
  or   g05880 ( new_n6257 , new_n6255 , new_n6256 );
  xor  g05881 ( new_n6258 , new_n6254 , new_n6257 );
  nand g05882 ( new_n6259 , new_n5956 , new_n5959 );
  not  g05883 ( new_n6260 , new_n5952 );
  nand g05884 ( new_n6261 , new_n6260 , new_n5960 );
  nand g05885 ( new_n6262 , new_n6259 , new_n6261 );
  nand g05886 ( new_n6263 , new_n5953 , new_n5954 );
  nand g05887 ( new_n6264 , new_n5934 , new_n5955 );
  nand g05888 ( new_n6265 , new_n6263 , new_n6264 );
  xor  g05889 ( new_n6266 , new_n6262 , new_n6265 );
  nand g05890 ( new_n6267 , new_n5945 , new_n5946 );
  nand g05891 ( new_n6268 , new_n5923 , new_n5947 );
  nand g05892 ( new_n6269 , new_n6267 , new_n6268 );
  xor  g05893 ( new_n6270 , new_n6266 , new_n6269 );
  nand g05894 ( new_n6271 , pi209 , pi241 );
  nand g05895 ( new_n6272 , pi034 , pi190 );
  nand g05896 ( new_n6273 , pi131 , pi220 );
  xor  g05897 ( new_n6274 , new_n6272 , new_n6273 );
  nand g05898 ( new_n6275 , new_n5995 , new_n6024 );
  not  g05899 ( new_n6276 , new_n6026 );
  nand g05900 ( new_n6277 , new_n6022 , new_n6276 );
  nand g05901 ( new_n6278 , new_n6275 , new_n6277 );
  xor  g05902 ( new_n6279 , new_n6274 , new_n6278 );
  xor  g05903 ( new_n6280 , new_n6271 , new_n6279 );
  xor  g05904 ( new_n6281 , new_n6270 , new_n6280 );
  xor  g05905 ( new_n6282 , new_n6258 , new_n6281 );
  nand g05906 ( new_n6283 , pi047 , pi089 );
  nand g05907 ( new_n6284 , pi128 , pi254 );
  xor  g05908 ( new_n6285 , new_n6283 , new_n6284 );
  xor  g05909 ( new_n6286 , new_n6282 , new_n6285 );
  xor  g05910 ( new_n6287 , new_n6253 , new_n6286 );
  xor  g05911 ( new_n6288 , new_n6250 , new_n6287 );
  nand g05912 ( new_n6289 , new_n6101 , new_n6112 );
  nand g05913 ( new_n6290 , new_n6113 , new_n6114 );
  nand g05914 ( new_n6291 , new_n6289 , new_n6290 );
  nand g05915 ( new_n6292 , pi035 , pi198 );
  nand g05916 ( new_n6293 , pi139 , pi165 );
  xor  g05917 ( new_n6294 , new_n6292 , new_n6293 );
  xor  g05918 ( new_n6295 , new_n6291 , new_n6294 );
  nand g05919 ( new_n6296 , pi120 , pi204 );
  not  g05920 ( new_n6297 , new_n6177 );
  nand g05921 ( new_n6298 , new_n6115 , new_n6297 );
  or   g05922 ( new_n6299 , new_n6178 , new_n6187 );
  nand g05923 ( new_n6300 , new_n6298 , new_n6299 );
  nand g05924 ( new_n6301 , pi064 , pi229 );
  nand g05925 ( new_n6302 , pi077 , pi185 );
  nand g05926 ( new_n6303 , pi030 , pi052 );
  xor  g05927 ( new_n6304 , new_n6302 , new_n6303 );
  xor  g05928 ( new_n6305 , new_n6301 , new_n6304 );
  xor  g05929 ( new_n6306 , new_n6300 , new_n6305 );
  nand g05930 ( new_n6307 , new_n6017 , new_n6020 );
  nand g05931 ( new_n6308 , new_n6013 , new_n6021 );
  nand g05932 ( new_n6309 , new_n6307 , new_n6308 );
  nand g05933 ( new_n6310 , new_n5994 , new_n6015 );
  nand g05934 ( new_n6311 , new_n6014 , new_n6016 );
  nand g05935 ( new_n6312 , new_n6310 , new_n6311 );
  xor  g05936 ( new_n6313 , new_n6309 , new_n6312 );
  nand g05937 ( new_n6314 , pi067 , pi189 );
  nand g05938 ( new_n6315 , pi053 , pi133 );
  xor  g05939 ( new_n6316 , new_n6314 , new_n6315 );
  xor  g05940 ( new_n6317 , new_n6313 , new_n6316 );
  or   g05941 ( new_n6318 , new_n6145 , new_n6167 );
  nand g05942 ( new_n6319 , new_n6168 , new_n6176 );
  nand g05943 ( new_n6320 , new_n6318 , new_n6319 );
  nand g05944 ( new_n6321 , pi084 , pi092 );
  xor  g05945 ( new_n6322 , new_n6320 , new_n6321 );
  xor  g05946 ( new_n6323 , new_n6317 , new_n6322 );
  nand g05947 ( new_n6324 , pi062 , pi146 );
  nand g05948 ( new_n6325 , pi078 , pi168 );
  xor  g05949 ( new_n6326 , new_n6324 , new_n6325 );
  nand g05950 ( new_n6327 , pi065 , pi152 );
  or   g05951 ( new_n6328 , new_n6136 , new_n6165 );
  nand g05952 ( new_n6329 , new_n6162 , new_n6166 );
  nand g05953 ( new_n6330 , new_n6328 , new_n6329 );
  xor  g05954 ( new_n6331 , new_n6327 , new_n6330 );
  xor  g05955 ( new_n6332 , new_n6326 , new_n6331 );
  nand g05956 ( new_n6333 , new_n6007 , new_n6008 );
  nand g05957 ( new_n6334 , new_n5987 , new_n6009 );
  nand g05958 ( new_n6335 , new_n6333 , new_n6334 );
  or   g05959 ( new_n6336 , new_n5988 , new_n6011 );
  not  g05960 ( new_n6337 , new_n6010 );
  nand g05961 ( new_n6338 , new_n6337 , new_n6012 );
  nand g05962 ( new_n6339 , new_n6336 , new_n6338 );
  xor  g05963 ( new_n6340 , new_n6335 , new_n6339 );
  xor  g05964 ( new_n6341 , new_n6332 , new_n6340 );
  xor  g05965 ( new_n6342 , new_n6323 , new_n6341 );
  xor  g05966 ( new_n6343 , new_n6306 , new_n6342 );
  xor  g05967 ( new_n6344 , new_n6296 , new_n6343 );
  xor  g05968 ( new_n6345 , new_n6295 , new_n6344 );
  nand g05969 ( new_n6346 , pi022 , pi213 );
  or   g05970 ( new_n6347 , new_n6067 , new_n6090 );
  nand g05971 ( new_n6348 , new_n6091 , new_n6100 );
  nand g05972 ( new_n6349 , new_n6347 , new_n6348 );
  xor  g05973 ( new_n6350 , new_n6346 , new_n6349 );
  nand g05974 ( new_n6351 , new_n6154 , new_n6155 );
  nand g05975 ( new_n6352 , new_n6135 , new_n6156 );
  nand g05976 ( new_n6353 , new_n6351 , new_n6352 );
  nor  g05977 ( new_n6354 , new_n6083 , new_n6089 );
  nor  g05978 ( new_n6355 , new_n6088 , new_n6354 );
  xor  g05979 ( new_n6356 , new_n6353 , new_n6355 );
  nand g05980 ( new_n6357 , pi004 , pi183 );
  nand g05981 ( new_n6358 , pi073 , pi105 );
  xor  g05982 ( new_n6359 , new_n6357 , new_n6358 );
  nand g05983 ( new_n6360 , pi088 , pi170 );
  xor  g05984 ( new_n6361 , new_n6359 , new_n6360 );
  xor  g05985 ( new_n6362 , new_n6356 , new_n6361 );
  xor  g05986 ( new_n6363 , new_n6350 , new_n6362 );
  nand g05987 ( new_n6364 , pi197 , pi208 );
  nand g05988 ( new_n6365 , new_n6146 , new_n6147 );
  nand g05989 ( new_n6366 , new_n6127 , new_n6148 );
  nand g05990 ( new_n6367 , new_n6365 , new_n6366 );
  nor  g05991 ( new_n6368 , new_n6129 , new_n6150 );
  nor  g05992 ( new_n6369 , new_n6149 , new_n6152 );
  or   g05993 ( new_n6370 , new_n6368 , new_n6369 );
  xor  g05994 ( new_n6371 , new_n6367 , new_n6370 );
  xor  g05995 ( new_n6372 , new_n6364 , new_n6371 );
  xor  g05996 ( new_n6373 , new_n6363 , new_n6372 );
  xor  g05997 ( new_n6374 , new_n6345 , new_n6373 );
  xor  g05998 ( new_n6375 , new_n6288 , new_n6374 );
  xor  g05999 ( po027 , new_n6214 , new_n6375 );
  nand g06000 ( new_n6377 , pi108 , pi141 );
  nand g06001 ( new_n6378 , new_n4598 , new_n4599 );
  nand g06002 ( new_n6379 , new_n4597 , new_n4600 );
  nand g06003 ( new_n6380 , new_n6378 , new_n6379 );
  xnor g06004 ( new_n6381 , new_n6377 , new_n6380 );
  nand g06005 ( new_n6382 , pi042 , pi090 );
  nand g06006 ( new_n6383 , pi047 , pi051 );
  nand g06007 ( new_n6384 , new_n6382 , new_n6383 );
  nand g06008 ( new_n6385 , pi042 , pi047 );
  or   g06009 ( new_n6386 , new_n4598 , new_n6385 );
  nand g06010 ( new_n6387 , new_n6384 , new_n6386 );
  xnor g06011 ( new_n6388 , new_n6381 , new_n6387 );
  nand g06012 ( new_n6389 , pi007 , pi161 );
  nand g06013 ( new_n6390 , pi118 , pi241 );
  and  g06014 ( new_n6391 , new_n6389 , new_n6390 );
  nand g06015 ( new_n6392 , pi118 , pi161 );
  nor  g06016 ( new_n6393 , new_n4602 , new_n6392 );
  or   g06017 ( new_n6394 , new_n6391 , new_n6393 );
  xnor g06018 ( new_n6395 , new_n6388 , new_n6394 );
  nand g06019 ( new_n6396 , new_n4602 , new_n4605 );
  nand g06020 ( new_n6397 , new_n4601 , new_n4606 );
  nand g06021 ( new_n6398 , new_n6396 , new_n6397 );
  xor  g06022 ( new_n6399 , new_n6395 , new_n6398 );
  not  g06023 ( new_n6400 , new_n4608 );
  nand g06024 ( new_n6401 , new_n6400 , new_n4612 );
  or   g06025 ( new_n6402 , new_n4607 , new_n4613 );
  nand g06026 ( new_n6403 , new_n6401 , new_n6402 );
  xnor g06027 ( new_n6404 , new_n6399 , new_n6403 );
  nand g06028 ( new_n6405 , new_n4596 , new_n4614 );
  nand g06029 ( new_n6406 , pi113 , pi236 );
  xor  g06030 ( new_n6407 , new_n6405 , new_n6406 );
  xnor g06031 ( new_n6408 , new_n6404 , new_n6407 );
  or   g06032 ( new_n6409 , new_n4635 , new_n4652 );
  nand g06033 ( new_n6410 , pi013 , pi061 );
  nand g06034 ( new_n6411 , pi105 , pi188 );
  nand g06035 ( new_n6412 , pi112 , pi178 );
  nand g06036 ( new_n6413 , new_n6411 , new_n6412 );
  nand g06037 ( new_n6414 , pi105 , pi178 );
  or   g06038 ( new_n6415 , new_n4636 , new_n6414 );
  nand g06039 ( new_n6416 , new_n6413 , new_n6415 );
  xor  g06040 ( new_n6417 , new_n6410 , new_n6416 );
  nand g06041 ( new_n6418 , new_n4637 , new_n4638 );
  nand g06042 ( new_n6419 , new_n4636 , new_n4639 );
  nand g06043 ( new_n6420 , new_n6418 , new_n6419 );
  xor  g06044 ( new_n6421 , new_n6417 , new_n6420 );
  nand g06045 ( new_n6422 , pi012 , pi104 );
  nand g06046 ( new_n6423 , pi144 , pi212 );
  and  g06047 ( new_n6424 , new_n6422 , new_n6423 );
  nand g06048 ( new_n6425 , pi104 , pi144 );
  nor  g06049 ( new_n6426 , new_n4641 , new_n6425 );
  or   g06050 ( new_n6427 , new_n6424 , new_n6426 );
  xnor g06051 ( new_n6428 , new_n6421 , new_n6427 );
  nand g06052 ( new_n6429 , new_n4641 , new_n4644 );
  nand g06053 ( new_n6430 , new_n4640 , new_n4645 );
  nand g06054 ( new_n6431 , new_n6429 , new_n6430 );
  xor  g06055 ( new_n6432 , new_n6428 , new_n6431 );
  or   g06056 ( new_n6433 , new_n4647 , new_n4650 );
  nand g06057 ( new_n6434 , new_n4646 , new_n4651 );
  nand g06058 ( new_n6435 , new_n6433 , new_n6434 );
  xnor g06059 ( new_n6436 , new_n6432 , new_n6435 );
  nand g06060 ( new_n6437 , pi098 , pi213 );
  xor  g06061 ( new_n6438 , new_n6436 , new_n6437 );
  xor  g06062 ( new_n6439 , new_n6409 , new_n6438 );
  xor  g06063 ( new_n6440 , new_n6408 , new_n6439 );
  nand g06064 ( new_n6441 , new_n4615 , new_n4653 );
  not  g06065 ( new_n6442 , new_n4681 );
  nand g06066 ( new_n6443 , new_n4654 , new_n6442 );
  nand g06067 ( new_n6444 , new_n6441 , new_n6443 );
  xnor g06068 ( new_n6445 , new_n6440 , new_n6444 );
  nand g06069 ( new_n6446 , pi035 , pi179 );
  nand g06070 ( new_n6447 , pi015 , pi033 );
  nand g06071 ( new_n6448 , pi162 , pi204 );
  nand g06072 ( new_n6449 , new_n6447 , new_n6448 );
  nand g06073 ( new_n6450 , pi033 , pi204 );
  or   g06074 ( new_n6451 , new_n4705 , new_n6450 );
  nand g06075 ( new_n6452 , new_n6449 , new_n6451 );
  xor  g06076 ( new_n6453 , new_n6446 , new_n6452 );
  nand g06077 ( new_n6454 , new_n4704 , new_n4705 );
  nand g06078 ( new_n6455 , new_n4703 , new_n4706 );
  nand g06079 ( new_n6456 , new_n6454 , new_n6455 );
  xor  g06080 ( new_n6457 , new_n6453 , new_n6456 );
  nand g06081 ( new_n6458 , pi048 , pi139 );
  nand g06082 ( new_n6459 , pi208 , pi237 );
  and  g06083 ( new_n6460 , new_n6458 , new_n6459 );
  nand g06084 ( new_n6461 , pi139 , pi237 );
  nor  g06085 ( new_n6462 , new_n4708 , new_n6461 );
  or   g06086 ( new_n6463 , new_n6460 , new_n6462 );
  xnor g06087 ( new_n6464 , new_n6457 , new_n6463 );
  nand g06088 ( new_n6465 , new_n4708 , new_n4711 );
  nand g06089 ( new_n6466 , new_n4707 , new_n4712 );
  nand g06090 ( new_n6467 , new_n6465 , new_n6466 );
  xor  g06091 ( new_n6468 , new_n6464 , new_n6467 );
  not  g06092 ( new_n6469 , new_n4714 );
  nand g06093 ( new_n6470 , new_n6469 , new_n4717 );
  or   g06094 ( new_n6471 , new_n4713 , new_n4718 );
  nand g06095 ( new_n6472 , new_n6470 , new_n6471 );
  xnor g06096 ( new_n6473 , new_n6468 , new_n6472 );
  nand g06097 ( new_n6474 , new_n4702 , new_n4719 );
  nand g06098 ( new_n6475 , pi168 , pi238 );
  xor  g06099 ( new_n6476 , new_n6474 , new_n6475 );
  xor  g06100 ( new_n6477 , new_n6473 , new_n6476 );
  or   g06101 ( new_n6478 , new_n4720 , new_n4745 );
  nand g06102 ( new_n6479 , new_n4682 , new_n4746 );
  nand g06103 ( new_n6480 , new_n6478 , new_n6479 );
  xor  g06104 ( new_n6481 , new_n6477 , new_n6480 );
  xor  g06105 ( new_n6482 , new_n6445 , new_n6481 );
  nand g06106 ( new_n6483 , pi133 , pi194 );
  nand g06107 ( new_n6484 , pi064 , pi143 );
  nand g06108 ( new_n6485 , pi057 , pi189 );
  nand g06109 ( new_n6486 , new_n6484 , new_n6485 );
  nand g06110 ( new_n6487 , pi057 , pi064 );
  or   g06111 ( new_n6488 , new_n4772 , new_n6487 );
  nand g06112 ( new_n6489 , new_n6486 , new_n6488 );
  xor  g06113 ( new_n6490 , new_n6483 , new_n6489 );
  nand g06114 ( new_n6491 , new_n4772 , new_n4773 );
  nand g06115 ( new_n6492 , new_n4771 , new_n4774 );
  nand g06116 ( new_n6493 , new_n6491 , new_n6492 );
  xor  g06117 ( new_n6494 , new_n6490 , new_n6493 );
  nand g06118 ( new_n6495 , pi077 , pi085 );
  nand g06119 ( new_n6496 , pi052 , pi180 );
  nand g06120 ( new_n6497 , new_n6495 , new_n6496 );
  nand g06121 ( new_n6498 , pi077 , pi180 );
  nor  g06122 ( new_n6499 , new_n4776 , new_n6498 );
  not  g06123 ( new_n6500 , new_n6499 );
  nand g06124 ( new_n6501 , new_n6497 , new_n6500 );
  xnor g06125 ( new_n6502 , new_n6494 , new_n6501 );
  nand g06126 ( new_n6503 , new_n4776 , new_n4779 );
  nand g06127 ( new_n6504 , new_n4775 , new_n4780 );
  nand g06128 ( new_n6505 , new_n6503 , new_n6504 );
  xor  g06129 ( new_n6506 , new_n6502 , new_n6505 );
  or   g06130 ( new_n6507 , new_n4781 , new_n4782 );
  nand g06131 ( new_n6508 , new_n4783 , new_n4786 );
  nand g06132 ( new_n6509 , new_n6507 , new_n6508 );
  xnor g06133 ( new_n6510 , new_n6506 , new_n6509 );
  nand g06134 ( new_n6511 , new_n4770 , new_n4787 );
  nand g06135 ( new_n6512 , pi036 , pi131 );
  xor  g06136 ( new_n6513 , new_n6511 , new_n6512 );
  xor  g06137 ( new_n6514 , new_n6510 , new_n6513 );
  not  g06138 ( new_n6515 , new_n4788 );
  nor  g06139 ( new_n6516 , new_n4747 , new_n6515 );
  nor  g06140 ( new_n6517 , new_n4789 , new_n4810 );
  nor  g06141 ( new_n6518 , new_n6516 , new_n6517 );
  xor  g06142 ( new_n6519 , new_n6514 , new_n6518 );
  xor  g06143 ( po028 , new_n6482 , new_n6519 );
  xnor g06144 ( po029 , new_n880 , new_n881 );
  xor  g06145 ( po030 , new_n1819 , new_n1820 );
  nand g06146 ( new_n6523 , pi163 , pi210 );
  nand g06147 ( new_n6524 , pi107 , pi242 );
  xor  g06148 ( new_n6525 , new_n6523 , new_n6524 );
  nand g06149 ( new_n6526 , pi175 , pi249 );
  xor  g06150 ( new_n6527 , new_n6525 , new_n6526 );
  nand g06151 ( new_n6528 , pi103 , pi217 );
  xor  g06152 ( po031 , new_n6527 , new_n6528 );
  xor  g06153 ( po032 , new_n2551 , new_n2569 );
  nand g06154 ( new_n6531 , pi140 , pi171 );
  nand g06155 ( new_n6532 , pi107 , pi252 );
  xor  g06156 ( new_n6533 , new_n6531 , new_n6532 );
  nand g06157 ( new_n6534 , pi049 , pi242 );
  xor  g06158 ( new_n6535 , new_n6533 , new_n6534 );
  nor  g06159 ( new_n6536 , new_n6524 , new_n6531 );
  xor  g06160 ( new_n6537 , new_n6535 , new_n6536 );
  not  g06161 ( new_n6538 , new_n6523 );
  nand g06162 ( new_n6539 , pi111 , pi148 );
  nor  g06163 ( new_n6540 , new_n6538 , new_n6539 );
  nand g06164 ( new_n6541 , pi210 , pi228 );
  nand g06165 ( new_n6542 , pi024 , pi163 );
  nand g06166 ( new_n6543 , new_n6541 , new_n6542 );
  or   g06167 ( new_n6544 , new_n6541 , new_n6542 );
  and  g06168 ( new_n6545 , new_n6543 , new_n6544 );
  or   g06169 ( new_n6546 , new_n6540 , new_n6545 );
  nand g06170 ( new_n6547 , new_n6540 , new_n6543 );
  nand g06171 ( new_n6548 , new_n6546 , new_n6547 );
  xor  g06172 ( new_n6549 , new_n6537 , new_n6548 );
  or   g06173 ( new_n6550 , new_n6523 , new_n6524 );
  nand g06174 ( new_n6551 , pi148 , pi210 );
  nand g06175 ( new_n6552 , pi111 , pi163 );
  nand g06176 ( new_n6553 , new_n6551 , new_n6552 );
  or   g06177 ( new_n6554 , new_n6523 , new_n6539 );
  nand g06178 ( new_n6555 , new_n6553 , new_n6554 );
  nor  g06179 ( new_n6556 , new_n6550 , new_n6555 );
  xnor g06180 ( new_n6557 , new_n6550 , new_n6555 );
  not  g06181 ( new_n6558 , new_n6536 );
  nand g06182 ( new_n6559 , pi107 , pi140 );
  nand g06183 ( new_n6560 , pi171 , pi242 );
  nand g06184 ( new_n6561 , new_n6559 , new_n6560 );
  nand g06185 ( new_n6562 , new_n6558 , new_n6561 );
  nor  g06186 ( new_n6563 , new_n6557 , new_n6562 );
  nor  g06187 ( new_n6564 , new_n6556 , new_n6563 );
  not  g06188 ( new_n6565 , new_n6564 );
  xor  g06189 ( new_n6566 , new_n6549 , new_n6565 );
  not  g06190 ( new_n6567 , new_n6525 );
  nor  g06191 ( new_n6568 , new_n6567 , new_n6526 );
  nand g06192 ( new_n6569 , pi134 , pi249 );
  nand g06193 ( new_n6570 , pi175 , pi222 );
  xor  g06194 ( new_n6571 , new_n6569 , new_n6570 );
  or   g06195 ( new_n6572 , new_n6568 , new_n6571 );
  xor  g06196 ( new_n6573 , new_n6557 , new_n6562 );
  not  g06197 ( new_n6574 , new_n6573 );
  xor  g06198 ( new_n6575 , new_n6568 , new_n6571 );
  nand g06199 ( new_n6576 , new_n6574 , new_n6575 );
  nand g06200 ( new_n6577 , new_n6572 , new_n6576 );
  nand g06201 ( new_n6578 , pi240 , pi249 );
  nand g06202 ( new_n6579 , pi125 , pi175 );
  nand g06203 ( new_n6580 , new_n6578 , new_n6579 );
  not  g06204 ( new_n6581 , new_n6580 );
  nand g06205 ( new_n6582 , pi134 , pi222 );
  not  g06206 ( new_n6583 , new_n6582 );
  nand g06207 ( new_n6584 , new_n6526 , new_n6583 );
  nor  g06208 ( new_n6585 , new_n6581 , new_n6584 );
  nand g06209 ( new_n6586 , new_n6581 , new_n6584 );
  or   g06210 ( new_n6587 , new_n6578 , new_n6579 );
  nand g06211 ( new_n6588 , new_n6586 , new_n6587 );
  or   g06212 ( new_n6589 , new_n6585 , new_n6588 );
  xor  g06213 ( new_n6590 , new_n6577 , new_n6589 );
  not  g06214 ( new_n6591 , new_n6590 );
  xor  g06215 ( new_n6592 , new_n6566 , new_n6591 );
  or   g06216 ( new_n6593 , new_n6527 , new_n6528 );
  nand g06217 ( new_n6594 , pi100 , pi103 );
  nand g06218 ( new_n6595 , pi117 , pi217 );
  nand g06219 ( new_n6596 , new_n6594 , new_n6595 );
  nand g06220 ( new_n6597 , pi100 , pi117 );
  or   g06221 ( new_n6598 , new_n6528 , new_n6597 );
  nand g06222 ( new_n6599 , new_n6596 , new_n6598 );
  or   g06223 ( new_n6600 , new_n6593 , new_n6599 );
  xor  g06224 ( new_n6601 , new_n6573 , new_n6575 );
  xor  g06225 ( new_n6602 , new_n6593 , new_n6599 );
  nand g06226 ( new_n6603 , new_n6601 , new_n6602 );
  nand g06227 ( new_n6604 , new_n6600 , new_n6603 );
  not  g06228 ( new_n6605 , new_n6528 );
  nor  g06229 ( new_n6606 , new_n6605 , new_n6597 );
  nand g06230 ( new_n6607 , pi103 , pi227 );
  nand g06231 ( new_n6608 , pi016 , pi217 );
  nand g06232 ( new_n6609 , new_n6607 , new_n6608 );
  or   g06233 ( new_n6610 , new_n6607 , new_n6608 );
  and  g06234 ( new_n6611 , new_n6609 , new_n6610 );
  nor  g06235 ( new_n6612 , new_n6606 , new_n6611 );
  not  g06236 ( new_n6613 , new_n6612 );
  nand g06237 ( new_n6614 , new_n6606 , new_n6609 );
  and  g06238 ( new_n6615 , new_n6613 , new_n6614 );
  xor  g06239 ( new_n6616 , new_n6604 , new_n6615 );
  xnor g06240 ( po033 , new_n6592 , new_n6616 );
  xor  g06241 ( po034 , new_n4564 , new_n4566 );
  xor  g06242 ( po035 , new_n4040 , new_n4041 );
  nand g06243 ( new_n6620 , pi080 , pi227 );
  nand g06244 ( new_n6621 , pi217 , pi234 );
  nand g06245 ( new_n6622 , pi100 , pi247 );
  nand g06246 ( new_n6623 , new_n6621 , new_n6622 );
  nand g06247 ( new_n6624 , pi217 , pi247 );
  nand g06248 ( new_n6625 , pi100 , pi234 );
  or   g06249 ( new_n6626 , new_n6624 , new_n6625 );
  nand g06250 ( new_n6627 , new_n6623 , new_n6626 );
  xor  g06251 ( new_n6628 , new_n6620 , new_n6627 );
  nand g06252 ( new_n6629 , pi016 , pi227 );
  nand g06253 ( new_n6630 , pi080 , pi100 );
  nand g06254 ( new_n6631 , new_n6629 , new_n6630 );
  xor  g06255 ( new_n6632 , new_n6629 , new_n6630 );
  nand g06256 ( new_n6633 , new_n6624 , new_n6632 );
  nand g06257 ( new_n6634 , new_n6631 , new_n6633 );
  xor  g06258 ( new_n6635 , new_n6628 , new_n6634 );
  nand g06259 ( new_n6636 , pi016 , pi081 );
  nand g06260 ( new_n6637 , pi106 , pi117 );
  nand g06261 ( new_n6638 , new_n6636 , new_n6637 );
  nand g06262 ( new_n6639 , pi016 , pi106 );
  nand g06263 ( new_n6640 , pi081 , pi117 );
  nor  g06264 ( new_n6641 , new_n6639 , new_n6640 );
  not  g06265 ( new_n6642 , new_n6641 );
  nand g06266 ( new_n6643 , new_n6638 , new_n6642 );
  xnor g06267 ( new_n6644 , new_n6635 , new_n6643 );
  nand g06268 ( new_n6645 , pi016 , pi100 );
  nand g06269 ( new_n6646 , pi080 , pi217 );
  nand g06270 ( new_n6647 , new_n6645 , new_n6646 );
  nand g06271 ( new_n6648 , pi117 , pi227 );
  xor  g06272 ( new_n6649 , new_n6645 , new_n6646 );
  nand g06273 ( new_n6650 , new_n6648 , new_n6649 );
  nand g06274 ( new_n6651 , new_n6647 , new_n6650 );
  nand g06275 ( new_n6652 , new_n6640 , new_n6651 );
  xor  g06276 ( new_n6653 , new_n6624 , new_n6632 );
  xor  g06277 ( new_n6654 , new_n6640 , new_n6651 );
  nand g06278 ( new_n6655 , new_n6653 , new_n6654 );
  nand g06279 ( new_n6656 , new_n6652 , new_n6655 );
  xor  g06280 ( new_n6657 , new_n6644 , new_n6656 );
  xor  g06281 ( new_n6658 , new_n6653 , new_n6654 );
  nand g06282 ( new_n6659 , pi103 , pi106 );
  or   g06283 ( new_n6660 , new_n6658 , new_n6659 );
  xor  g06284 ( new_n6661 , new_n6658 , new_n6659 );
  nand g06285 ( new_n6662 , pi081 , pi103 );
  nand g06286 ( new_n6663 , new_n6597 , new_n6610 );
  nand g06287 ( new_n6664 , new_n6609 , new_n6663 );
  or   g06288 ( new_n6665 , new_n6662 , new_n6664 );
  xnor g06289 ( new_n6666 , new_n6648 , new_n6649 );
  xor  g06290 ( new_n6667 , new_n6662 , new_n6664 );
  nand g06291 ( new_n6668 , new_n6666 , new_n6667 );
  nand g06292 ( new_n6669 , new_n6665 , new_n6668 );
  nand g06293 ( new_n6670 , new_n6661 , new_n6669 );
  nand g06294 ( new_n6671 , new_n6660 , new_n6670 );
  nand g06295 ( new_n6672 , new_n6657 , new_n6671 );
  nand g06296 ( new_n6673 , pi214 , pi217 );
  nand g06297 ( new_n6674 , pi227 , pi247 );
  xor  g06298 ( new_n6675 , new_n6673 , new_n6674 );
  xor  g06299 ( new_n6676 , new_n6625 , new_n6675 );
  nand g06300 ( new_n6677 , pi080 , pi081 );
  xor  g06301 ( new_n6678 , new_n6626 , new_n6677 );
  xor  g06302 ( new_n6679 , new_n6676 , new_n6678 );
  nand g06303 ( new_n6680 , pi117 , pi233 );
  nand g06304 ( new_n6681 , pi103 , pi187 );
  xor  g06305 ( new_n6682 , new_n6680 , new_n6681 );
  xor  g06306 ( new_n6683 , new_n6639 , new_n6682 );
  nand g06307 ( new_n6684 , new_n6620 , new_n6627 );
  nand g06308 ( new_n6685 , new_n6628 , new_n6634 );
  nand g06309 ( new_n6686 , new_n6684 , new_n6685 );
  xor  g06310 ( new_n6687 , new_n6683 , new_n6686 );
  xnor g06311 ( new_n6688 , new_n6679 , new_n6687 );
  nor  g06312 ( new_n6689 , new_n6644 , new_n6656 );
  and  g06313 ( new_n6690 , new_n6641 , new_n6689 );
  or   g06314 ( new_n6691 , new_n6635 , new_n6643 );
  nand g06315 ( new_n6692 , new_n6642 , new_n6691 );
  nor  g06316 ( new_n6693 , new_n6689 , new_n6692 );
  or   g06317 ( new_n6694 , new_n6690 , new_n6693 );
  xor  g06318 ( new_n6695 , new_n6688 , new_n6694 );
  xnor g06319 ( new_n6696 , new_n6672 , new_n6695 );
  nand g06320 ( new_n6697 , pi103 , pi233 );
  xor  g06321 ( new_n6698 , new_n6666 , new_n6667 );
  nor  g06322 ( new_n6699 , new_n6598 , new_n6613 );
  nand g06323 ( new_n6700 , new_n6698 , new_n6699 );
  not  g06324 ( new_n6701 , new_n6700 );
  xor  g06325 ( new_n6702 , new_n6661 , new_n6669 );
  nand g06326 ( new_n6703 , new_n6701 , new_n6702 );
  nand g06327 ( new_n6704 , new_n6697 , new_n6703 );
  xnor g06328 ( new_n6705 , new_n6657 , new_n6671 );
  xor  g06329 ( new_n6706 , new_n6697 , new_n6703 );
  nand g06330 ( new_n6707 , new_n6705 , new_n6706 );
  nand g06331 ( new_n6708 , new_n6704 , new_n6707 );
  xor  g06332 ( new_n6709 , new_n6696 , new_n6708 );
  or   g06333 ( new_n6710 , new_n6535 , new_n6558 );
  nand g06334 ( new_n6711 , pi107 , pi121 );
  nand g06335 ( new_n6712 , new_n6531 , new_n6532 );
  nand g06336 ( new_n6713 , new_n6533 , new_n6534 );
  nand g06337 ( new_n6714 , new_n6712 , new_n6713 );
  xor  g06338 ( new_n6715 , new_n6711 , new_n6714 );
  nand g06339 ( new_n6716 , pi171 , pi252 );
  nand g06340 ( new_n6717 , pi242 , pi245 );
  nand g06341 ( new_n6718 , pi049 , pi140 );
  xor  g06342 ( new_n6719 , new_n6717 , new_n6718 );
  xnor g06343 ( new_n6720 , new_n6716 , new_n6719 );
  xnor g06344 ( new_n6721 , new_n6715 , new_n6720 );
  nor  g06345 ( new_n6722 , new_n6710 , new_n6721 );
  nand g06346 ( new_n6723 , pi049 , pi252 );
  nand g06347 ( new_n6724 , pi201 , pi242 );
  nand g06348 ( new_n6725 , pi140 , pi245 );
  xor  g06349 ( new_n6726 , new_n6724 , new_n6725 );
  xor  g06350 ( new_n6727 , new_n6723 , new_n6726 );
  nand g06351 ( new_n6728 , pi121 , pi171 );
  nand g06352 ( new_n6729 , new_n6717 , new_n6718 );
  nand g06353 ( new_n6730 , new_n6716 , new_n6719 );
  nand g06354 ( new_n6731 , new_n6729 , new_n6730 );
  xor  g06355 ( new_n6732 , new_n6728 , new_n6731 );
  xor  g06356 ( new_n6733 , new_n6727 , new_n6732 );
  nand g06357 ( new_n6734 , pi107 , pi231 );
  or   g06358 ( new_n6735 , new_n6711 , new_n6714 );
  nand g06359 ( new_n6736 , new_n6715 , new_n6720 );
  nand g06360 ( new_n6737 , new_n6735 , new_n6736 );
  xor  g06361 ( new_n6738 , new_n6734 , new_n6737 );
  xor  g06362 ( new_n6739 , new_n6733 , new_n6738 );
  xnor g06363 ( new_n6740 , new_n6722 , new_n6739 );
  nand g06364 ( new_n6741 , pi039 , pi210 );
  nand g06365 ( new_n6742 , pi111 , pi228 );
  nand g06366 ( new_n6743 , pi024 , pi148 );
  xor  g06367 ( new_n6744 , new_n6742 , new_n6743 );
  xor  g06368 ( new_n6745 , new_n6741 , new_n6744 );
  nand g06369 ( new_n6746 , new_n6539 , new_n6544 );
  nand g06370 ( new_n6747 , new_n6543 , new_n6746 );
  nand g06371 ( new_n6748 , pi163 , pi224 );
  xor  g06372 ( new_n6749 , new_n6747 , new_n6748 );
  xor  g06373 ( new_n6750 , new_n6745 , new_n6749 );
  nor  g06374 ( new_n6751 , new_n6546 , new_n6554 );
  not  g06375 ( new_n6752 , new_n6751 );
  nor  g06376 ( new_n6753 , new_n6750 , new_n6752 );
  nand g06377 ( new_n6754 , pi116 , pi210 );
  nand g06378 ( new_n6755 , pi024 , pi228 );
  nand g06379 ( new_n6756 , pi039 , pi111 );
  xor  g06380 ( new_n6757 , new_n6755 , new_n6756 );
  xor  g06381 ( new_n6758 , new_n6754 , new_n6757 );
  nand g06382 ( new_n6759 , pi148 , pi224 );
  nand g06383 ( new_n6760 , new_n6742 , new_n6743 );
  nand g06384 ( new_n6761 , new_n6741 , new_n6744 );
  nand g06385 ( new_n6762 , new_n6760 , new_n6761 );
  xor  g06386 ( new_n6763 , new_n6759 , new_n6762 );
  xnor g06387 ( new_n6764 , new_n6758 , new_n6763 );
  nand g06388 ( new_n6765 , pi163 , pi255 );
  nand g06389 ( new_n6766 , new_n6747 , new_n6748 );
  nand g06390 ( new_n6767 , new_n6745 , new_n6749 );
  nand g06391 ( new_n6768 , new_n6766 , new_n6767 );
  xor  g06392 ( new_n6769 , new_n6765 , new_n6768 );
  xnor g06393 ( new_n6770 , new_n6764 , new_n6769 );
  xor  g06394 ( new_n6771 , new_n6753 , new_n6770 );
  xor  g06395 ( new_n6772 , new_n6710 , new_n6721 );
  or   g06396 ( new_n6773 , new_n6537 , new_n6548 );
  nand g06397 ( new_n6774 , new_n6549 , new_n6565 );
  nand g06398 ( new_n6775 , new_n6773 , new_n6774 );
  or   g06399 ( new_n6776 , new_n6772 , new_n6775 );
  xor  g06400 ( new_n6777 , new_n6750 , new_n6752 );
  not  g06401 ( new_n6778 , new_n6777 );
  xor  g06402 ( new_n6779 , new_n6772 , new_n6775 );
  nand g06403 ( new_n6780 , new_n6778 , new_n6779 );
  nand g06404 ( new_n6781 , new_n6776 , new_n6780 );
  xor  g06405 ( new_n6782 , new_n6771 , new_n6781 );
  xnor g06406 ( new_n6783 , new_n6740 , new_n6782 );
  nand g06407 ( new_n6784 , pi149 , pi249 );
  nand g06408 ( new_n6785 , pi222 , pi240 );
  nand g06409 ( new_n6786 , pi125 , pi134 );
  xor  g06410 ( new_n6787 , new_n6785 , new_n6786 );
  xnor g06411 ( new_n6788 , new_n6784 , new_n6787 );
  nand g06412 ( new_n6789 , new_n6582 , new_n6587 );
  nand g06413 ( new_n6790 , new_n6580 , new_n6789 );
  nand g06414 ( new_n6791 , pi175 , pi176 );
  xor  g06415 ( new_n6792 , new_n6790 , new_n6791 );
  xor  g06416 ( new_n6793 , new_n6788 , new_n6792 );
  not  g06417 ( new_n6794 , new_n6793 );
  nand g06418 ( new_n6795 , new_n6583 , new_n6588 );
  nor  g06419 ( new_n6796 , new_n6794 , new_n6795 );
  nand g06420 ( new_n6797 , pi167 , pi249 );
  nand g06421 ( new_n6798 , pi125 , pi240 );
  nand g06422 ( new_n6799 , pi149 , pi222 );
  xor  g06423 ( new_n6800 , new_n6798 , new_n6799 );
  xor  g06424 ( new_n6801 , new_n6797 , new_n6800 );
  nand g06425 ( new_n6802 , pi134 , pi176 );
  nand g06426 ( new_n6803 , new_n6785 , new_n6786 );
  nand g06427 ( new_n6804 , new_n6784 , new_n6787 );
  nand g06428 ( new_n6805 , new_n6803 , new_n6804 );
  xor  g06429 ( new_n6806 , new_n6802 , new_n6805 );
  xor  g06430 ( new_n6807 , new_n6801 , new_n6806 );
  nand g06431 ( new_n6808 , pi040 , pi175 );
  xor  g06432 ( new_n6809 , new_n6807 , new_n6808 );
  or   g06433 ( new_n6810 , new_n6790 , new_n6791 );
  nand g06434 ( new_n6811 , new_n6788 , new_n6792 );
  nand g06435 ( new_n6812 , new_n6810 , new_n6811 );
  xor  g06436 ( new_n6813 , new_n6809 , new_n6812 );
  xor  g06437 ( new_n6814 , new_n6796 , new_n6813 );
  nor  g06438 ( new_n6815 , new_n6783 , new_n6814 );
  xor  g06439 ( new_n6816 , new_n6783 , new_n6814 );
  not  g06440 ( new_n6817 , new_n6816 );
  xor  g06441 ( new_n6818 , new_n6793 , new_n6795 );
  nand g06442 ( new_n6819 , new_n6577 , new_n6589 );
  or   g06443 ( new_n6820 , new_n6566 , new_n6591 );
  nand g06444 ( new_n6821 , new_n6819 , new_n6820 );
  or   g06445 ( new_n6822 , new_n6818 , new_n6821 );
  xor  g06446 ( new_n6823 , new_n6777 , new_n6779 );
  xor  g06447 ( new_n6824 , new_n6818 , new_n6821 );
  nand g06448 ( new_n6825 , new_n6823 , new_n6824 );
  nand g06449 ( new_n6826 , new_n6822 , new_n6825 );
  nor  g06450 ( new_n6827 , new_n6817 , new_n6826 );
  nor  g06451 ( new_n6828 , new_n6815 , new_n6827 );
  nand g06452 ( new_n6829 , pi125 , pi149 );
  nand g06453 ( new_n6830 , pi167 , pi222 );
  nand g06454 ( new_n6831 , pi181 , pi249 );
  nand g06455 ( new_n6832 , new_n6830 , new_n6831 );
  nand g06456 ( new_n6833 , pi181 , pi222 );
  or   g06457 ( new_n6834 , new_n6797 , new_n6833 );
  nand g06458 ( new_n6835 , new_n6832 , new_n6834 );
  xor  g06459 ( new_n6836 , new_n6829 , new_n6835 );
  nand g06460 ( new_n6837 , new_n6798 , new_n6799 );
  nand g06461 ( new_n6838 , new_n6797 , new_n6800 );
  nand g06462 ( new_n6839 , new_n6837 , new_n6838 );
  xor  g06463 ( new_n6840 , new_n6836 , new_n6839 );
  nand g06464 ( new_n6841 , new_n6802 , new_n6805 );
  nand g06465 ( new_n6842 , new_n6801 , new_n6806 );
  nand g06466 ( new_n6843 , new_n6841 , new_n6842 );
  nand g06467 ( new_n6844 , pi176 , pi240 );
  nand g06468 ( new_n6845 , pi040 , pi134 );
  nand g06469 ( new_n6846 , new_n6844 , new_n6845 );
  nand g06470 ( new_n6847 , pi040 , pi240 );
  or   g06471 ( new_n6848 , new_n6802 , new_n6847 );
  nand g06472 ( new_n6849 , new_n6846 , new_n6848 );
  xor  g06473 ( new_n6850 , new_n6843 , new_n6849 );
  xnor g06474 ( new_n6851 , new_n6840 , new_n6850 );
  or   g06475 ( new_n6852 , new_n6807 , new_n6808 );
  nand g06476 ( new_n6853 , new_n6809 , new_n6812 );
  nand g06477 ( new_n6854 , new_n6852 , new_n6853 );
  xnor g06478 ( new_n6855 , new_n6851 , new_n6854 );
  nand g06479 ( new_n6856 , new_n6796 , new_n6813 );
  nand g06480 ( new_n6857 , pi174 , pi175 );
  xor  g06481 ( new_n6858 , new_n6856 , new_n6857 );
  xnor g06482 ( new_n6859 , new_n6855 , new_n6858 );
  not  g06483 ( new_n6860 , new_n6753 );
  nor  g06484 ( new_n6861 , new_n6860 , new_n6770 );
  nand g06485 ( new_n6862 , pi127 , pi163 );
  nand g06486 ( new_n6863 , pi024 , pi039 );
  nand g06487 ( new_n6864 , pi111 , pi116 );
  nand g06488 ( new_n6865 , pi070 , pi210 );
  nand g06489 ( new_n6866 , new_n6864 , new_n6865 );
  nand g06490 ( new_n6867 , pi070 , pi111 );
  or   g06491 ( new_n6868 , new_n6754 , new_n6867 );
  nand g06492 ( new_n6869 , new_n6866 , new_n6868 );
  xor  g06493 ( new_n6870 , new_n6863 , new_n6869 );
  nand g06494 ( new_n6871 , new_n6755 , new_n6756 );
  nand g06495 ( new_n6872 , new_n6754 , new_n6757 );
  nand g06496 ( new_n6873 , new_n6871 , new_n6872 );
  xor  g06497 ( new_n6874 , new_n6870 , new_n6873 );
  nand g06498 ( new_n6875 , pi224 , pi228 );
  nand g06499 ( new_n6876 , pi148 , pi255 );
  and  g06500 ( new_n6877 , new_n6875 , new_n6876 );
  nand g06501 ( new_n6878 , pi228 , pi255 );
  nor  g06502 ( new_n6879 , new_n6759 , new_n6878 );
  or   g06503 ( new_n6880 , new_n6877 , new_n6879 );
  xnor g06504 ( new_n6881 , new_n6874 , new_n6880 );
  nand g06505 ( new_n6882 , new_n6759 , new_n6762 );
  nand g06506 ( new_n6883 , new_n6758 , new_n6763 );
  nand g06507 ( new_n6884 , new_n6882 , new_n6883 );
  xor  g06508 ( new_n6885 , new_n6881 , new_n6884 );
  or   g06509 ( new_n6886 , new_n6765 , new_n6768 );
  nand g06510 ( new_n6887 , new_n6764 , new_n6769 );
  nand g06511 ( new_n6888 , new_n6886 , new_n6887 );
  xnor g06512 ( new_n6889 , new_n6885 , new_n6888 );
  xor  g06513 ( new_n6890 , new_n6862 , new_n6889 );
  xnor g06514 ( new_n6891 , new_n6861 , new_n6890 );
  nand g06515 ( new_n6892 , new_n6722 , new_n6739 );
  not  g06516 ( new_n6893 , new_n6892 );
  nand g06517 ( new_n6894 , pi005 , pi107 );
  nand g06518 ( new_n6895 , pi245 , pi252 );
  nand g06519 ( new_n6896 , new_n6724 , new_n6725 );
  nand g06520 ( new_n6897 , new_n6723 , new_n6726 );
  nand g06521 ( new_n6898 , new_n6896 , new_n6897 );
  xor  g06522 ( new_n6899 , new_n6895 , new_n6898 );
  nand g06523 ( new_n6900 , pi140 , pi201 );
  nand g06524 ( new_n6901 , pi156 , pi242 );
  nand g06525 ( new_n6902 , new_n6900 , new_n6901 );
  nand g06526 ( new_n6903 , pi140 , pi156 );
  nor  g06527 ( new_n6904 , new_n6724 , new_n6903 );
  not  g06528 ( new_n6905 , new_n6904 );
  nand g06529 ( new_n6906 , new_n6902 , new_n6905 );
  xor  g06530 ( new_n6907 , new_n6899 , new_n6906 );
  nand g06531 ( new_n6908 , pi171 , pi231 );
  nand g06532 ( new_n6909 , pi049 , pi121 );
  and  g06533 ( new_n6910 , new_n6908 , new_n6909 );
  nand g06534 ( new_n6911 , pi049 , pi231 );
  nor  g06535 ( new_n6912 , new_n6728 , new_n6911 );
  or   g06536 ( new_n6913 , new_n6910 , new_n6912 );
  xnor g06537 ( new_n6914 , new_n6907 , new_n6913 );
  nand g06538 ( new_n6915 , new_n6728 , new_n6731 );
  nand g06539 ( new_n6916 , new_n6727 , new_n6732 );
  nand g06540 ( new_n6917 , new_n6915 , new_n6916 );
  xor  g06541 ( new_n6918 , new_n6914 , new_n6917 );
  not  g06542 ( new_n6919 , new_n6734 );
  nand g06543 ( new_n6920 , new_n6919 , new_n6737 );
  or   g06544 ( new_n6921 , new_n6733 , new_n6738 );
  nand g06545 ( new_n6922 , new_n6920 , new_n6921 );
  xnor g06546 ( new_n6923 , new_n6918 , new_n6922 );
  xor  g06547 ( new_n6924 , new_n6894 , new_n6923 );
  xor  g06548 ( new_n6925 , new_n6893 , new_n6924 );
  xor  g06549 ( new_n6926 , new_n6891 , new_n6925 );
  nand g06550 ( new_n6927 , new_n6771 , new_n6781 );
  nand g06551 ( new_n6928 , new_n6740 , new_n6782 );
  nand g06552 ( new_n6929 , new_n6927 , new_n6928 );
  xor  g06553 ( new_n6930 , new_n6926 , new_n6929 );
  xor  g06554 ( new_n6931 , new_n6859 , new_n6930 );
  xor  g06555 ( new_n6932 , new_n6828 , new_n6931 );
  not  g06556 ( new_n6933 , new_n6932 );
  xor  g06557 ( new_n6934 , new_n6705 , new_n6706 );
  or   g06558 ( new_n6935 , new_n6933 , new_n6934 );
  xor  g06559 ( new_n6936 , new_n6933 , new_n6934 );
  xor  g06560 ( new_n6937 , new_n6700 , new_n6702 );
  xnor g06561 ( new_n6938 , new_n6698 , new_n6699 );
  or   g06562 ( new_n6939 , new_n6604 , new_n6615 );
  nand g06563 ( new_n6940 , new_n6592 , new_n6616 );
  nand g06564 ( new_n6941 , new_n6939 , new_n6940 );
  nand g06565 ( new_n6942 , new_n6938 , new_n6941 );
  xor  g06566 ( new_n6943 , new_n6823 , new_n6824 );
  not  g06567 ( new_n6944 , new_n6943 );
  xor  g06568 ( new_n6945 , new_n6938 , new_n6941 );
  nand g06569 ( new_n6946 , new_n6944 , new_n6945 );
  nand g06570 ( new_n6947 , new_n6942 , new_n6946 );
  or   g06571 ( new_n6948 , new_n6937 , new_n6947 );
  xor  g06572 ( new_n6949 , new_n6816 , new_n6826 );
  xor  g06573 ( new_n6950 , new_n6937 , new_n6947 );
  nand g06574 ( new_n6951 , new_n6949 , new_n6950 );
  nand g06575 ( new_n6952 , new_n6948 , new_n6951 );
  nand g06576 ( new_n6953 , new_n6936 , new_n6952 );
  nand g06577 ( new_n6954 , new_n6935 , new_n6953 );
  or   g06578 ( new_n6955 , new_n6709 , new_n6954 );
  not  g06579 ( new_n6956 , new_n6925 );
  nor  g06580 ( new_n6957 , new_n6891 , new_n6956 );
  nor  g06581 ( new_n6958 , new_n6926 , new_n6929 );
  nor  g06582 ( new_n6959 , new_n6957 , new_n6958 );
  nand g06583 ( new_n6960 , new_n6885 , new_n6888 );
  nand g06584 ( new_n6961 , pi115 , pi210 );
  nand g06585 ( new_n6962 , pi024 , pi116 );
  xor  g06586 ( new_n6963 , new_n6961 , new_n6962 );
  xor  g06587 ( new_n6964 , new_n6867 , new_n6963 );
  not  g06588 ( new_n6965 , new_n6964 );
  nand g06589 ( new_n6966 , pi039 , pi224 );
  xor  g06590 ( new_n6967 , new_n6868 , new_n6966 );
  xor  g06591 ( new_n6968 , new_n6965 , new_n6967 );
  nand g06592 ( new_n6969 , pi163 , pi232 );
  nand g06593 ( new_n6970 , pi127 , pi148 );
  xor  g06594 ( new_n6971 , new_n6969 , new_n6970 );
  xor  g06595 ( new_n6972 , new_n6878 , new_n6971 );
  nand g06596 ( new_n6973 , new_n6863 , new_n6869 );
  nand g06597 ( new_n6974 , new_n6870 , new_n6873 );
  nand g06598 ( new_n6975 , new_n6973 , new_n6974 );
  xor  g06599 ( new_n6976 , new_n6972 , new_n6975 );
  xor  g06600 ( new_n6977 , new_n6968 , new_n6976 );
  nor  g06601 ( new_n6978 , new_n6881 , new_n6884 );
  nand g06602 ( new_n6979 , new_n6879 , new_n6978 );
  nor  g06603 ( new_n6980 , new_n6874 , new_n6880 );
  or   g06604 ( new_n6981 , new_n6879 , new_n6980 );
  or   g06605 ( new_n6982 , new_n6978 , new_n6981 );
  nand g06606 ( new_n6983 , new_n6979 , new_n6982 );
  xor  g06607 ( new_n6984 , new_n6977 , new_n6983 );
  xor  g06608 ( new_n6985 , new_n6960 , new_n6984 );
  or   g06609 ( new_n6986 , new_n6862 , new_n6889 );
  nand g06610 ( new_n6987 , new_n6861 , new_n6890 );
  nand g06611 ( new_n6988 , new_n6986 , new_n6987 );
  xor  g06612 ( new_n6989 , new_n6985 , new_n6988 );
  nand g06613 ( new_n6990 , new_n6918 , new_n6922 );
  nand g06614 ( new_n6991 , pi063 , pi242 );
  nand g06615 ( new_n6992 , pi201 , pi252 );
  xor  g06616 ( new_n6993 , new_n6991 , new_n6992 );
  xor  g06617 ( new_n6994 , new_n6903 , new_n6993 );
  nand g06618 ( new_n6995 , pi121 , pi245 );
  xor  g06619 ( new_n6996 , new_n6905 , new_n6995 );
  not  g06620 ( new_n6997 , new_n6996 );
  xor  g06621 ( new_n6998 , new_n6994 , new_n6997 );
  nand g06622 ( new_n6999 , pi021 , pi107 );
  nand g06623 ( new_n7000 , pi005 , pi171 );
  xor  g06624 ( new_n7001 , new_n6999 , new_n7000 );
  xor  g06625 ( new_n7002 , new_n6911 , new_n7001 );
  nand g06626 ( new_n7003 , new_n6895 , new_n6898 );
  nand g06627 ( new_n7004 , new_n6899 , new_n6906 );
  nand g06628 ( new_n7005 , new_n7003 , new_n7004 );
  xor  g06629 ( new_n7006 , new_n7002 , new_n7005 );
  xor  g06630 ( new_n7007 , new_n6998 , new_n7006 );
  nor  g06631 ( new_n7008 , new_n6914 , new_n6917 );
  nand g06632 ( new_n7009 , new_n6912 , new_n7008 );
  nor  g06633 ( new_n7010 , new_n6907 , new_n6913 );
  or   g06634 ( new_n7011 , new_n6912 , new_n7010 );
  or   g06635 ( new_n7012 , new_n7008 , new_n7011 );
  nand g06636 ( new_n7013 , new_n7009 , new_n7012 );
  xor  g06637 ( new_n7014 , new_n7007 , new_n7013 );
  xor  g06638 ( new_n7015 , new_n6990 , new_n7014 );
  or   g06639 ( new_n7016 , new_n6894 , new_n6923 );
  nand g06640 ( new_n7017 , new_n6893 , new_n6924 );
  nand g06641 ( new_n7018 , new_n7016 , new_n7017 );
  xor  g06642 ( new_n7019 , new_n7015 , new_n7018 );
  xor  g06643 ( new_n7020 , new_n6989 , new_n7019 );
  xnor g06644 ( new_n7021 , new_n6959 , new_n7020 );
  nand g06645 ( new_n7022 , new_n6851 , new_n6854 );
  nand g06646 ( new_n7023 , pi200 , pi249 );
  nand g06647 ( new_n7024 , pi125 , pi167 );
  xor  g06648 ( new_n7025 , new_n7023 , new_n7024 );
  xor  g06649 ( new_n7026 , new_n6833 , new_n7025 );
  not  g06650 ( new_n7027 , new_n7026 );
  nand g06651 ( new_n7028 , pi149 , pi176 );
  xor  g06652 ( new_n7029 , new_n6834 , new_n7028 );
  xor  g06653 ( new_n7030 , new_n7027 , new_n7029 );
  nand g06654 ( new_n7031 , pi157 , pi175 );
  nand g06655 ( new_n7032 , pi134 , pi174 );
  xor  g06656 ( new_n7033 , new_n7031 , new_n7032 );
  xor  g06657 ( new_n7034 , new_n6847 , new_n7033 );
  nand g06658 ( new_n7035 , new_n6829 , new_n6835 );
  nand g06659 ( new_n7036 , new_n6836 , new_n6839 );
  nand g06660 ( new_n7037 , new_n7035 , new_n7036 );
  xor  g06661 ( new_n7038 , new_n7034 , new_n7037 );
  xor  g06662 ( new_n7039 , new_n7030 , new_n7038 );
  not  g06663 ( new_n7040 , new_n7039 );
  nand g06664 ( new_n7041 , new_n6843 , new_n6849 );
  nand g06665 ( new_n7042 , new_n6840 , new_n6850 );
  nand g06666 ( new_n7043 , new_n7041 , new_n7042 );
  xor  g06667 ( new_n7044 , new_n6848 , new_n7043 );
  xor  g06668 ( new_n7045 , new_n7040 , new_n7044 );
  xnor g06669 ( new_n7046 , new_n7022 , new_n7045 );
  nand g06670 ( new_n7047 , new_n6856 , new_n6857 );
  nand g06671 ( new_n7048 , new_n6855 , new_n6858 );
  nand g06672 ( new_n7049 , new_n7047 , new_n7048 );
  xor  g06673 ( new_n7050 , new_n7046 , new_n7049 );
  xor  g06674 ( new_n7051 , new_n7021 , new_n7050 );
  nand g06675 ( new_n7052 , new_n6859 , new_n6930 );
  nand g06676 ( new_n7053 , new_n6828 , new_n6931 );
  nand g06677 ( new_n7054 , new_n7052 , new_n7053 );
  xor  g06678 ( new_n7055 , new_n7051 , new_n7054 );
  not  g06679 ( new_n7056 , new_n7055 );
  xor  g06680 ( new_n7057 , new_n6709 , new_n6954 );
  nand g06681 ( new_n7058 , new_n7056 , new_n7057 );
  nand g06682 ( new_n7059 , new_n6955 , new_n7058 );
  nand g06683 ( new_n7060 , pi021 , pi171 );
  nand g06684 ( new_n7061 , new_n6991 , new_n6992 );
  nand g06685 ( new_n7062 , new_n6903 , new_n6993 );
  nand g06686 ( new_n7063 , new_n7061 , new_n7062 );
  xor  g06687 ( new_n7064 , new_n7060 , new_n7063 );
  nor  g06688 ( new_n7065 , new_n6688 , new_n6694 );
  nor  g06689 ( new_n7066 , new_n6693 , new_n7065 );
  nand g06690 ( new_n7067 , pi039 , pi255 );
  nand g06691 ( new_n7068 , new_n6969 , new_n6970 );
  nand g06692 ( new_n7069 , new_n6878 , new_n6971 );
  nand g06693 ( new_n7070 , new_n7068 , new_n7069 );
  xor  g06694 ( new_n7071 , new_n7067 , new_n7070 );
  or   g06695 ( new_n7072 , new_n7007 , new_n7013 );
  nand g06696 ( new_n7073 , new_n7012 , new_n7072 );
  nand g06697 ( new_n7074 , pi121 , pi201 );
  nand g06698 ( new_n7075 , pi231 , pi245 );
  xor  g06699 ( new_n7076 , new_n7074 , new_n7075 );
  xor  g06700 ( new_n7077 , new_n7073 , new_n7076 );
  xor  g06701 ( new_n7078 , new_n7071 , new_n7077 );
  xor  g06702 ( new_n7079 , new_n7066 , new_n7078 );
  xor  g06703 ( new_n7080 , new_n7064 , new_n7079 );
  xor  g06704 ( new_n7081 , new_n7059 , new_n7080 );
  or   g06705 ( new_n7082 , new_n6990 , new_n7014 );
  nand g06706 ( new_n7083 , new_n7015 , new_n7018 );
  nand g06707 ( new_n7084 , new_n7082 , new_n7083 );
  nor  g06708 ( new_n7085 , new_n6672 , new_n6695 );
  nor  g06709 ( new_n7086 , new_n6696 , new_n6708 );
  or   g06710 ( new_n7087 , new_n7085 , new_n7086 );
  xor  g06711 ( new_n7088 , new_n7084 , new_n7087 );
  nor  g06712 ( new_n7089 , new_n6905 , new_n6995 );
  nor  g06713 ( new_n7090 , new_n6994 , new_n6997 );
  or   g06714 ( new_n7091 , new_n7089 , new_n7090 );
  xor  g06715 ( new_n7092 , new_n7088 , new_n7091 );
  nand g06716 ( new_n7093 , pi125 , pi181 );
  nand g06717 ( new_n7094 , pi000 , pi210 );
  nand g06718 ( new_n7095 , pi024 , pi070 );
  nand g06719 ( new_n7096 , pi111 , pi115 );
  xor  g06720 ( new_n7097 , new_n7095 , new_n7096 );
  nand g06721 ( new_n7098 , pi163 , pi191 );
  or   g06722 ( new_n7099 , new_n6989 , new_n7019 );
  nand g06723 ( new_n7100 , new_n6959 , new_n7020 );
  nand g06724 ( new_n7101 , new_n7099 , new_n7100 );
  xor  g06725 ( new_n7102 , new_n7098 , new_n7101 );
  xor  g06726 ( new_n7103 , new_n7097 , new_n7102 );
  xor  g06727 ( new_n7104 , new_n7094 , new_n7103 );
  xor  g06728 ( new_n7105 , new_n7093 , new_n7104 );
  nand g06729 ( new_n7106 , pi167 , pi176 );
  or   g06730 ( new_n7107 , new_n6834 , new_n7028 );
  nand g06731 ( new_n7108 , new_n7027 , new_n7029 );
  nand g06732 ( new_n7109 , new_n7107 , new_n7108 );
  xor  g06733 ( new_n7110 , new_n7106 , new_n7109 );
  or   g06734 ( new_n7111 , new_n6960 , new_n6984 );
  nand g06735 ( new_n7112 , new_n6985 , new_n6988 );
  nand g06736 ( new_n7113 , new_n7111 , new_n7112 );
  nand g06737 ( new_n7114 , pi134 , pi157 );
  nand g06738 ( new_n7115 , new_n7023 , new_n7024 );
  nand g06739 ( new_n7116 , new_n6833 , new_n7025 );
  nand g06740 ( new_n7117 , new_n7115 , new_n7116 );
  or   g06741 ( new_n7118 , new_n7034 , new_n7037 );
  nand g06742 ( new_n7119 , new_n7030 , new_n7038 );
  nand g06743 ( new_n7120 , new_n7118 , new_n7119 );
  xor  g06744 ( new_n7121 , new_n7117 , new_n7120 );
  xor  g06745 ( new_n7122 , new_n7114 , new_n7121 );
  xor  g06746 ( new_n7123 , new_n7113 , new_n7122 );
  xor  g06747 ( new_n7124 , new_n7110 , new_n7123 );
  or   g06748 ( new_n7125 , new_n6977 , new_n6983 );
  nand g06749 ( new_n7126 , new_n6982 , new_n7125 );
  nand g06750 ( new_n7127 , new_n7031 , new_n7032 );
  nand g06751 ( new_n7128 , new_n6847 , new_n7033 );
  nand g06752 ( new_n7129 , new_n7127 , new_n7128 );
  xor  g06753 ( new_n7130 , new_n7126 , new_n7129 );
  nand g06754 ( new_n7131 , pi040 , pi149 );
  nand g06755 ( new_n7132 , pi174 , pi240 );
  xor  g06756 ( new_n7133 , new_n7131 , new_n7132 );
  xor  g06757 ( new_n7134 , new_n7130 , new_n7133 );
  xor  g06758 ( new_n7135 , new_n7124 , new_n7134 );
  xor  g06759 ( new_n7136 , new_n7105 , new_n7135 );
  nand g06760 ( new_n7137 , pi117 , pi187 );
  nand g06761 ( new_n7138 , pi100 , pi214 );
  xor  g06762 ( new_n7139 , new_n7137 , new_n7138 );
  xor  g06763 ( new_n7140 , new_n7136 , new_n7139 );
  nand g06764 ( new_n7141 , new_n6673 , new_n6674 );
  nand g06765 ( new_n7142 , new_n6625 , new_n6675 );
  nand g06766 ( new_n7143 , new_n7141 , new_n7142 );
  nand g06767 ( new_n7144 , pi081 , pi247 );
  nand g06768 ( new_n7145 , pi080 , pi106 );
  xor  g06769 ( new_n7146 , new_n7144 , new_n7145 );
  xor  g06770 ( new_n7147 , new_n7143 , new_n7146 );
  nand g06771 ( new_n7148 , pi016 , pi233 );
  nor  g06772 ( new_n7149 , new_n7022 , new_n7045 );
  nor  g06773 ( new_n7150 , new_n7046 , new_n7049 );
  or   g06774 ( new_n7151 , new_n7149 , new_n7150 );
  nand g06775 ( new_n7152 , pi203 , pi249 );
  xor  g06776 ( new_n7153 , new_n7151 , new_n7152 );
  nand g06777 ( new_n7154 , new_n6848 , new_n7043 );
  nand g06778 ( new_n7155 , new_n7040 , new_n7044 );
  nand g06779 ( new_n7156 , new_n7154 , new_n7155 );
  nand g06780 ( new_n7157 , new_n6683 , new_n6686 );
  nand g06781 ( new_n7158 , new_n6679 , new_n6687 );
  nand g06782 ( new_n7159 , new_n7157 , new_n7158 );
  nand g06783 ( new_n7160 , new_n6680 , new_n6681 );
  nand g06784 ( new_n7161 , new_n6639 , new_n6682 );
  nand g06785 ( new_n7162 , new_n7160 , new_n7161 );
  nand g06786 ( new_n7163 , pi200 , pi222 );
  nand g06787 ( new_n7164 , pi017 , pi175 );
  xor  g06788 ( new_n7165 , new_n7163 , new_n7164 );
  xor  g06789 ( new_n7166 , new_n7162 , new_n7165 );
  xor  g06790 ( new_n7167 , new_n7159 , new_n7166 );
  xor  g06791 ( new_n7168 , new_n7156 , new_n7167 );
  xor  g06792 ( new_n7169 , new_n7153 , new_n7168 );
  xor  g06793 ( new_n7170 , new_n7148 , new_n7169 );
  xor  g06794 ( new_n7171 , new_n7147 , new_n7170 );
  or   g06795 ( new_n7172 , new_n6626 , new_n6677 );
  not  g06796 ( new_n7173 , new_n6676 );
  nand g06797 ( new_n7174 , new_n7173 , new_n6678 );
  nand g06798 ( new_n7175 , new_n7172 , new_n7174 );
  nand g06799 ( new_n7176 , pi227 , pi234 );
  xor  g06800 ( new_n7177 , new_n7175 , new_n7176 );
  xor  g06801 ( new_n7178 , new_n7171 , new_n7177 );
  xor  g06802 ( new_n7179 , new_n7140 , new_n7178 );
  nand g06803 ( new_n7180 , new_n6999 , new_n7000 );
  nand g06804 ( new_n7181 , new_n6911 , new_n7001 );
  nand g06805 ( new_n7182 , new_n7180 , new_n7181 );
  or   g06806 ( new_n7183 , new_n7002 , new_n7005 );
  nand g06807 ( new_n7184 , new_n6998 , new_n7006 );
  nand g06808 ( new_n7185 , new_n7183 , new_n7184 );
  xor  g06809 ( new_n7186 , new_n7182 , new_n7185 );
  nand g06810 ( new_n7187 , pi005 , pi049 );
  xor  g06811 ( new_n7188 , new_n7186 , new_n7187 );
  xor  g06812 ( new_n7189 , new_n7179 , new_n7188 );
  xor  g06813 ( new_n7190 , new_n7092 , new_n7189 );
  nand g06814 ( new_n7191 , new_n7021 , new_n7050 );
  nand g06815 ( new_n7192 , new_n7051 , new_n7054 );
  nand g06816 ( new_n7193 , new_n7191 , new_n7192 );
  nand g06817 ( new_n7194 , pi202 , pi217 );
  nand g06818 ( new_n7195 , pi103 , pi129 );
  xor  g06819 ( new_n7196 , new_n7194 , new_n7195 );
  or   g06820 ( new_n7197 , new_n6972 , new_n6975 );
  nand g06821 ( new_n7198 , new_n6968 , new_n6976 );
  nand g06822 ( new_n7199 , new_n7197 , new_n7198 );
  xor  g06823 ( new_n7200 , new_n7196 , new_n7199 );
  nand g06824 ( new_n7201 , pi116 , pi224 );
  or   g06825 ( new_n7202 , new_n6868 , new_n6966 );
  nand g06826 ( new_n7203 , new_n6965 , new_n6967 );
  nand g06827 ( new_n7204 , new_n7202 , new_n7203 );
  nand g06828 ( new_n7205 , new_n6961 , new_n6962 );
  nand g06829 ( new_n7206 , new_n6867 , new_n6963 );
  nand g06830 ( new_n7207 , new_n7205 , new_n7206 );
  xor  g06831 ( new_n7208 , new_n7204 , new_n7207 );
  nand g06832 ( new_n7209 , pi148 , pi232 );
  nand g06833 ( new_n7210 , pi127 , pi228 );
  xor  g06834 ( new_n7211 , new_n7209 , new_n7210 );
  xor  g06835 ( new_n7212 , new_n7208 , new_n7211 );
  xor  g06836 ( new_n7213 , new_n7201 , new_n7212 );
  nand g06837 ( new_n7214 , pi063 , pi140 );
  nand g06838 ( new_n7215 , pi082 , pi107 );
  nand g06839 ( new_n7216 , pi156 , pi252 );
  nand g06840 ( new_n7217 , pi083 , pi242 );
  xor  g06841 ( new_n7218 , new_n7216 , new_n7217 );
  xor  g06842 ( new_n7219 , new_n7215 , new_n7218 );
  xor  g06843 ( new_n7220 , new_n7214 , new_n7219 );
  xor  g06844 ( new_n7221 , new_n7213 , new_n7220 );
  xor  g06845 ( new_n7222 , new_n7200 , new_n7221 );
  xor  g06846 ( new_n7223 , new_n7193 , new_n7222 );
  xor  g06847 ( new_n7224 , new_n7190 , new_n7223 );
  xor  g06848 ( po036 , new_n7081 , new_n7224 );
  xor  g06849 ( po037 , new_n6936 , new_n6952 );
  xnor g06850 ( po038 , new_n3259 , new_n3260 );
  nand g06851 ( new_n7228 , pi013 , pi145 );
  nand g06852 ( new_n7229 , pi112 , pi164 );
  nand g06853 ( new_n7230 , pi105 , pi206 );
  or   g06854 ( new_n7231 , new_n7229 , new_n7230 );
  or   g06855 ( new_n7232 , new_n7228 , new_n7231 );
  nand g06856 ( new_n7233 , pi164 , pi183 );
  nand g06857 ( new_n7234 , pi032 , pi112 );
  xor  g06858 ( new_n7235 , new_n7233 , new_n7234 );
  xor  g06859 ( new_n7236 , new_n7230 , new_n7235 );
  not  g06860 ( new_n7237 , new_n7236 );
  xor  g06861 ( new_n7238 , new_n7228 , new_n7231 );
  nand g06862 ( new_n7239 , new_n7237 , new_n7238 );
  nand g06863 ( new_n7240 , new_n7232 , new_n7239 );
  nand g06864 ( new_n7241 , pi054 , pi077 );
  nand g06865 ( new_n7242 , pi044 , pi052 );
  nor  g06866 ( new_n7243 , new_n7241 , new_n7242 );
  nand g06867 ( new_n7244 , pi133 , pi250 );
  nand g06868 ( new_n7245 , pi045 , pi189 );
  nand g06869 ( new_n7246 , pi064 , pi119 );
  nand g06870 ( new_n7247 , new_n7245 , new_n7246 );
  nand g06871 ( new_n7248 , pi119 , pi189 );
  nand g06872 ( new_n7249 , pi045 , pi064 );
  or   g06873 ( new_n7250 , new_n7248 , new_n7249 );
  nand g06874 ( new_n7251 , new_n7247 , new_n7250 );
  xor  g06875 ( new_n7252 , new_n7244 , new_n7251 );
  nand g06876 ( new_n7253 , pi077 , pi250 );
  nand g06877 ( new_n7254 , new_n7248 , new_n7253 );
  nand g06878 ( new_n7255 , pi045 , pi133 );
  xor  g06879 ( new_n7256 , new_n7248 , new_n7253 );
  nand g06880 ( new_n7257 , new_n7255 , new_n7256 );
  nand g06881 ( new_n7258 , new_n7254 , new_n7257 );
  xor  g06882 ( new_n7259 , new_n7252 , new_n7258 );
  nand g06883 ( new_n7260 , pi044 , pi077 );
  nand g06884 ( new_n7261 , pi052 , pi054 );
  and  g06885 ( new_n7262 , new_n7260 , new_n7261 );
  or   g06886 ( new_n7263 , new_n7243 , new_n7262 );
  xnor g06887 ( new_n7264 , new_n7259 , new_n7263 );
  nand g06888 ( new_n7265 , pi119 , pi133 );
  nand g06889 ( new_n7266 , pi045 , pi077 );
  nand g06890 ( new_n7267 , new_n7265 , new_n7266 );
  nand g06891 ( new_n7268 , pi052 , pi250 );
  xor  g06892 ( new_n7269 , new_n7265 , new_n7266 );
  nand g06893 ( new_n7270 , new_n7268 , new_n7269 );
  nand g06894 ( new_n7271 , new_n7267 , new_n7270 );
  nand g06895 ( new_n7272 , new_n7242 , new_n7271 );
  xor  g06896 ( new_n7273 , new_n7255 , new_n7256 );
  xor  g06897 ( new_n7274 , new_n7242 , new_n7271 );
  nand g06898 ( new_n7275 , new_n7273 , new_n7274 );
  nand g06899 ( new_n7276 , new_n7272 , new_n7275 );
  nor  g06900 ( new_n7277 , new_n7264 , new_n7276 );
  nand g06901 ( new_n7278 , new_n7243 , new_n7277 );
  nand g06902 ( new_n7279 , pi189 , pi250 );
  nand g06903 ( new_n7280 , pi084 , pi119 );
  xor  g06904 ( new_n7281 , new_n7279 , new_n7280 );
  xor  g06905 ( new_n7282 , new_n7249 , new_n7281 );
  nand g06906 ( new_n7283 , pi044 , pi133 );
  xor  g06907 ( new_n7284 , new_n7250 , new_n7283 );
  xor  g06908 ( new_n7285 , new_n7282 , new_n7284 );
  nand g06909 ( new_n7286 , pi052 , pi072 );
  nand g06910 ( new_n7287 , pi131 , pi248 );
  xor  g06911 ( new_n7288 , new_n7286 , new_n7287 );
  xor  g06912 ( new_n7289 , new_n7241 , new_n7288 );
  nand g06913 ( new_n7290 , new_n7244 , new_n7251 );
  nand g06914 ( new_n7291 , new_n7252 , new_n7258 );
  nand g06915 ( new_n7292 , new_n7290 , new_n7291 );
  xor  g06916 ( new_n7293 , new_n7289 , new_n7292 );
  xnor g06917 ( new_n7294 , new_n7285 , new_n7293 );
  nor  g06918 ( new_n7295 , new_n7259 , new_n7263 );
  xor  g06919 ( new_n7296 , new_n7243 , new_n7277 );
  nor  g06920 ( new_n7297 , new_n7295 , new_n7296 );
  not  g06921 ( new_n7298 , new_n7297 );
  nand g06922 ( new_n7299 , new_n7294 , new_n7298 );
  nand g06923 ( new_n7300 , new_n7278 , new_n7299 );
  nand g06924 ( new_n7301 , pi235 , pi241 );
  xor  g06925 ( new_n7302 , new_n7264 , new_n7276 );
  nand g06926 ( new_n7303 , pi054 , pi131 );
  nand g06927 ( new_n7304 , pi044 , pi131 );
  nand g06928 ( new_n7305 , pi131 , pi250 );
  nand g06929 ( new_n7306 , pi045 , pi052 );
  nand g06930 ( new_n7307 , new_n7305 , new_n7306 );
  nand g06931 ( new_n7308 , pi077 , pi119 );
  xor  g06932 ( new_n7309 , new_n7305 , new_n7306 );
  nand g06933 ( new_n7310 , new_n7308 , new_n7309 );
  nand g06934 ( new_n7311 , new_n7307 , new_n7310 );
  nand g06935 ( new_n7312 , new_n7304 , new_n7311 );
  xor  g06936 ( new_n7313 , new_n7268 , new_n7269 );
  xor  g06937 ( new_n7314 , new_n7304 , new_n7311 );
  nand g06938 ( new_n7315 , new_n7313 , new_n7314 );
  nand g06939 ( new_n7316 , new_n7312 , new_n7315 );
  or   g06940 ( new_n7317 , new_n7303 , new_n7316 );
  xor  g06941 ( new_n7318 , new_n7303 , new_n7316 );
  xnor g06942 ( new_n7319 , new_n7273 , new_n7274 );
  nand g06943 ( new_n7320 , new_n7318 , new_n7319 );
  nand g06944 ( new_n7321 , new_n7317 , new_n7320 );
  xor  g06945 ( new_n7322 , new_n7302 , new_n7321 );
  nand g06946 ( new_n7323 , pi072 , pi131 );
  xor  g06947 ( new_n7324 , new_n7308 , new_n7309 );
  nand g06948 ( new_n7325 , pi045 , pi131 );
  nand g06949 ( new_n7326 , pi052 , pi119 );
  nor  g06950 ( new_n7327 , new_n7325 , new_n7326 );
  not  g06951 ( new_n7328 , new_n7327 );
  or   g06952 ( new_n7329 , new_n7324 , new_n7328 );
  xor  g06953 ( new_n7330 , new_n7313 , new_n7314 );
  nor  g06954 ( new_n7331 , new_n7329 , new_n7330 );
  xor  g06955 ( new_n7332 , new_n7318 , new_n7319 );
  nand g06956 ( new_n7333 , new_n7331 , new_n7332 );
  xor  g06957 ( new_n7334 , new_n7323 , new_n7333 );
  xor  g06958 ( new_n7335 , new_n7322 , new_n7334 );
  xor  g06959 ( new_n7336 , new_n7331 , new_n7332 );
  not  g06960 ( new_n7337 , new_n7336 );
  nand g06961 ( new_n7338 , pi104 , pi164 );
  nand g06962 ( new_n7339 , pi206 , pi212 );
  nand g06963 ( new_n7340 , pi032 , pi213 );
  xor  g06964 ( new_n7341 , new_n7339 , new_n7340 );
  xor  g06965 ( new_n7342 , new_n7338 , new_n7341 );
  or   g06966 ( new_n7343 , new_n378 , new_n7339 );
  or   g06967 ( new_n7344 , new_n7342 , new_n7343 );
  nand g06968 ( new_n7345 , pi032 , pi212 );
  nand g06969 ( new_n7346 , pi104 , pi206 );
  nand g06970 ( new_n7347 , pi013 , pi164 );
  xor  g06971 ( new_n7348 , new_n7346 , new_n7347 );
  xor  g06972 ( new_n7349 , new_n7345 , new_n7348 );
  nand g06973 ( new_n7350 , pi145 , pi213 );
  nand g06974 ( new_n7351 , new_n7339 , new_n7340 );
  nand g06975 ( new_n7352 , new_n7338 , new_n7341 );
  nand g06976 ( new_n7353 , new_n7351 , new_n7352 );
  xor  g06977 ( new_n7354 , new_n7350 , new_n7353 );
  xor  g06978 ( new_n7355 , new_n7349 , new_n7354 );
  nor  g06979 ( new_n7356 , new_n7344 , new_n7355 );
  nand g06980 ( new_n7357 , pi032 , pi104 );
  nand g06981 ( new_n7358 , pi013 , pi206 );
  xor  g06982 ( new_n7359 , new_n7357 , new_n7358 );
  xor  g06983 ( new_n7360 , new_n7229 , new_n7359 );
  nand g06984 ( new_n7361 , pi145 , pi212 );
  nand g06985 ( new_n7362 , new_n7346 , new_n7347 );
  nand g06986 ( new_n7363 , new_n7345 , new_n7348 );
  nand g06987 ( new_n7364 , new_n7362 , new_n7363 );
  xor  g06988 ( new_n7365 , new_n7361 , new_n7364 );
  xor  g06989 ( new_n7366 , new_n7360 , new_n7365 );
  nand g06990 ( new_n7367 , pi213 , pi246 );
  xnor g06991 ( new_n7368 , new_n7366 , new_n7367 );
  nand g06992 ( new_n7369 , new_n7350 , new_n7353 );
  nand g06993 ( new_n7370 , new_n7349 , new_n7354 );
  nand g06994 ( new_n7371 , new_n7369 , new_n7370 );
  xor  g06995 ( new_n7372 , new_n7368 , new_n7371 );
  xnor g06996 ( new_n7373 , new_n7356 , new_n7372 );
  nand g06997 ( new_n7374 , pi027 , pi161 );
  nand g06998 ( new_n7375 , pi008 , pi236 );
  nand g06999 ( new_n7376 , new_n7374 , new_n7375 );
  nand g07000 ( new_n7377 , pi026 , pi241 );
  or   g07001 ( new_n7378 , new_n7374 , new_n7375 );
  nand g07002 ( new_n7379 , new_n7377 , new_n7378 );
  nand g07003 ( new_n7380 , new_n7376 , new_n7379 );
  nand g07004 ( new_n7381 , pi056 , pi236 );
  xor  g07005 ( new_n7382 , new_n7380 , new_n7381 );
  nand g07006 ( new_n7383 , pi026 , pi161 );
  nand g07007 ( new_n7384 , pi027 , pi141 );
  nand g07008 ( new_n7385 , pi008 , pi241 );
  xor  g07009 ( new_n7386 , new_n7384 , new_n7385 );
  xor  g07010 ( new_n7387 , new_n7383 , new_n7386 );
  xor  g07011 ( new_n7388 , new_n7382 , new_n7387 );
  not  g07012 ( new_n7389 , new_n7377 );
  not  g07013 ( new_n7390 , new_n7376 );
  nand g07014 ( new_n7391 , new_n377 , new_n7389 );
  nand g07015 ( new_n7392 , new_n7390 , new_n7391 );
  nand g07016 ( new_n7393 , new_n7378 , new_n7392 );
  nand g07017 ( new_n7394 , new_n7389 , new_n7393 );
  nor  g07018 ( new_n7395 , new_n7388 , new_n7394 );
  nand g07019 ( new_n7396 , pi008 , pi161 );
  nand g07020 ( new_n7397 , pi027 , pi090 );
  nand g07021 ( new_n7398 , pi026 , pi141 );
  xor  g07022 ( new_n7399 , new_n7397 , new_n7398 );
  xor  g07023 ( new_n7400 , new_n7396 , new_n7399 );
  nand g07024 ( new_n7401 , pi056 , pi241 );
  nand g07025 ( new_n7402 , new_n7384 , new_n7385 );
  nand g07026 ( new_n7403 , new_n7383 , new_n7386 );
  nand g07027 ( new_n7404 , new_n7402 , new_n7403 );
  xor  g07028 ( new_n7405 , new_n7401 , new_n7404 );
  xor  g07029 ( new_n7406 , new_n7400 , new_n7405 );
  nand g07030 ( new_n7407 , pi136 , pi236 );
  xor  g07031 ( new_n7408 , new_n7406 , new_n7407 );
  or   g07032 ( new_n7409 , new_n7380 , new_n7381 );
  not  g07033 ( new_n7410 , new_n7387 );
  nand g07034 ( new_n7411 , new_n7382 , new_n7410 );
  nand g07035 ( new_n7412 , new_n7409 , new_n7411 );
  xor  g07036 ( new_n7413 , new_n7408 , new_n7412 );
  xnor g07037 ( new_n7414 , new_n7395 , new_n7413 );
  xor  g07038 ( new_n7415 , new_n7388 , new_n7394 );
  xor  g07039 ( new_n7416 , new_n7342 , new_n7343 );
  nor  g07040 ( new_n7417 , new_n7390 , new_n7391 );
  nor  g07041 ( new_n7418 , new_n7393 , new_n7417 );
  nand g07042 ( new_n7419 , new_n7416 , new_n7418 );
  xor  g07043 ( new_n7420 , new_n7416 , new_n7418 );
  nor  g07044 ( new_n7421 , new_n377 , new_n378 );
  nand g07045 ( new_n7422 , pi027 , pi241 );
  nand g07046 ( new_n7423 , pi026 , pi236 );
  xor  g07047 ( new_n7424 , new_n7422 , new_n7423 );
  nand g07048 ( new_n7425 , new_n7421 , new_n7424 );
  xnor g07049 ( new_n7426 , new_n7421 , new_n7424 );
  nand g07050 ( new_n7427 , pi206 , pi213 );
  nand g07051 ( new_n7428 , pi164 , pi212 );
  nand g07052 ( new_n7429 , new_n7427 , new_n7428 );
  nand g07053 ( new_n7430 , new_n7343 , new_n7429 );
  or   g07054 ( new_n7431 , new_n7426 , new_n7430 );
  nand g07055 ( new_n7432 , new_n7425 , new_n7431 );
  nand g07056 ( new_n7433 , new_n7420 , new_n7432 );
  nand g07057 ( new_n7434 , new_n7419 , new_n7433 );
  or   g07058 ( new_n7435 , new_n7415 , new_n7434 );
  xnor g07059 ( new_n7436 , new_n7344 , new_n7355 );
  xor  g07060 ( new_n7437 , new_n7415 , new_n7434 );
  nand g07061 ( new_n7438 , new_n7436 , new_n7437 );
  nand g07062 ( new_n7439 , new_n7435 , new_n7438 );
  xor  g07063 ( new_n7440 , new_n7414 , new_n7439 );
  xor  g07064 ( new_n7441 , new_n7373 , new_n7440 );
  nand g07065 ( new_n7442 , pi035 , pi147 );
  nand g07066 ( new_n7443 , pi019 , pi208 );
  nand g07067 ( new_n7444 , pi139 , pi151 );
  xor  g07068 ( new_n7445 , new_n7443 , new_n7444 );
  xnor g07069 ( new_n7446 , new_n7442 , new_n7445 );
  nand g07070 ( new_n7447 , pi019 , pi168 );
  nand g07071 ( new_n7448 , pi139 , pi147 );
  nand g07072 ( new_n7449 , new_n7447 , new_n7448 );
  nand g07073 ( new_n7450 , pi151 , pi208 );
  or   g07074 ( new_n7451 , new_n7447 , new_n7448 );
  nand g07075 ( new_n7452 , new_n7450 , new_n7451 );
  nand g07076 ( new_n7453 , new_n7449 , new_n7452 );
  nand g07077 ( new_n7454 , pi097 , pi168 );
  xor  g07078 ( new_n7455 , new_n7453 , new_n7454 );
  xnor g07079 ( new_n7456 , new_n7446 , new_n7455 );
  not  g07080 ( new_n7457 , new_n7450 );
  not  g07081 ( new_n7458 , new_n7449 );
  nand g07082 ( new_n7459 , new_n380 , new_n7457 );
  nand g07083 ( new_n7460 , new_n7458 , new_n7459 );
  nand g07084 ( new_n7461 , new_n7451 , new_n7460 );
  nand g07085 ( new_n7462 , new_n7457 , new_n7461 );
  nor  g07086 ( new_n7463 , new_n7456 , new_n7462 );
  nand g07087 ( new_n7464 , pi019 , pi139 );
  nand g07088 ( new_n7465 , pi035 , pi151 );
  nand g07089 ( new_n7466 , pi015 , pi147 );
  xor  g07090 ( new_n7467 , new_n7465 , new_n7466 );
  xor  g07091 ( new_n7468 , new_n7464 , new_n7467 );
  nand g07092 ( new_n7469 , pi097 , pi208 );
  nand g07093 ( new_n7470 , new_n7443 , new_n7444 );
  nand g07094 ( new_n7471 , new_n7442 , new_n7445 );
  nand g07095 ( new_n7472 , new_n7470 , new_n7471 );
  xor  g07096 ( new_n7473 , new_n7469 , new_n7472 );
  xor  g07097 ( new_n7474 , new_n7468 , new_n7473 );
  nand g07098 ( new_n7475 , pi075 , pi168 );
  or   g07099 ( new_n7476 , new_n7453 , new_n7454 );
  nand g07100 ( new_n7477 , new_n7446 , new_n7455 );
  nand g07101 ( new_n7478 , new_n7476 , new_n7477 );
  xor  g07102 ( new_n7479 , new_n7475 , new_n7478 );
  xor  g07103 ( new_n7480 , new_n7474 , new_n7479 );
  xor  g07104 ( new_n7481 , new_n7463 , new_n7480 );
  not  g07105 ( new_n7482 , new_n7481 );
  xor  g07106 ( new_n7483 , new_n7441 , new_n7482 );
  xor  g07107 ( new_n7484 , new_n7436 , new_n7437 );
  xor  g07108 ( new_n7485 , new_n7456 , new_n7462 );
  not  g07109 ( new_n7486 , new_n7485 );
  nand g07110 ( new_n7487 , new_n7484 , new_n7486 );
  xor  g07111 ( new_n7488 , new_n7484 , new_n7486 );
  xor  g07112 ( new_n7489 , new_n7420 , new_n7432 );
  nor  g07113 ( new_n7490 , new_n7458 , new_n7459 );
  nor  g07114 ( new_n7491 , new_n7461 , new_n7490 );
  or   g07115 ( new_n7492 , new_n7489 , new_n7491 );
  xor  g07116 ( new_n7493 , new_n7489 , new_n7491 );
  not  g07117 ( new_n7494 , new_n379 );
  nor  g07118 ( new_n7495 , new_n7494 , new_n380 );
  nand g07119 ( new_n7496 , pi151 , pi168 );
  nand g07120 ( new_n7497 , pi147 , pi208 );
  xor  g07121 ( new_n7498 , new_n7496 , new_n7497 );
  or   g07122 ( new_n7499 , new_n7495 , new_n7498 );
  xnor g07123 ( new_n7500 , new_n7426 , new_n7430 );
  xor  g07124 ( new_n7501 , new_n7495 , new_n7498 );
  nand g07125 ( new_n7502 , new_n7500 , new_n7501 );
  nand g07126 ( new_n7503 , new_n7499 , new_n7502 );
  nand g07127 ( new_n7504 , new_n7493 , new_n7503 );
  nand g07128 ( new_n7505 , new_n7492 , new_n7504 );
  nand g07129 ( new_n7506 , new_n7488 , new_n7505 );
  nand g07130 ( new_n7507 , new_n7487 , new_n7506 );
  xor  g07131 ( new_n7508 , new_n7483 , new_n7507 );
  nor  g07132 ( new_n7509 , new_n7337 , new_n7508 );
  xor  g07133 ( new_n7510 , new_n7337 , new_n7508 );
  not  g07134 ( new_n7511 , new_n7510 );
  xor  g07135 ( new_n7512 , new_n7329 , new_n7330 );
  not  g07136 ( new_n7513 , new_n7512 );
  xor  g07137 ( new_n7514 , new_n7488 , new_n7505 );
  nor  g07138 ( new_n7515 , new_n7513 , new_n7514 );
  xor  g07139 ( new_n7516 , new_n7512 , new_n7514 );
  xor  g07140 ( new_n7517 , new_n7493 , new_n7503 );
  nor  g07141 ( new_n7518 , new_n381 , new_n382 );
  xor  g07142 ( new_n7519 , new_n7325 , new_n7326 );
  or   g07143 ( new_n7520 , new_n7518 , new_n7519 );
  xor  g07144 ( new_n7521 , new_n7500 , new_n7501 );
  xor  g07145 ( new_n7522 , new_n7518 , new_n7519 );
  nand g07146 ( new_n7523 , new_n7521 , new_n7522 );
  nand g07147 ( new_n7524 , new_n7520 , new_n7523 );
  nand g07148 ( new_n7525 , new_n7517 , new_n7524 );
  xor  g07149 ( new_n7526 , new_n7324 , new_n7328 );
  not  g07150 ( new_n7527 , new_n7526 );
  xor  g07151 ( new_n7528 , new_n7517 , new_n7524 );
  nand g07152 ( new_n7529 , new_n7527 , new_n7528 );
  nand g07153 ( new_n7530 , new_n7525 , new_n7529 );
  nor  g07154 ( new_n7531 , new_n7516 , new_n7530 );
  nor  g07155 ( new_n7532 , new_n7515 , new_n7531 );
  nor  g07156 ( new_n7533 , new_n7511 , new_n7532 );
  or   g07157 ( new_n7534 , new_n7509 , new_n7533 );
  nand g07158 ( new_n7535 , new_n7335 , new_n7534 );
  nand g07159 ( new_n7536 , pi013 , pi032 );
  nand g07160 ( new_n7537 , pi112 , pi206 );
  nand g07161 ( new_n7538 , pi105 , pi164 );
  nand g07162 ( new_n7539 , new_n7537 , new_n7538 );
  nand g07163 ( new_n7540 , new_n7231 , new_n7539 );
  xor  g07164 ( new_n7541 , new_n7536 , new_n7540 );
  nand g07165 ( new_n7542 , new_n7357 , new_n7358 );
  nand g07166 ( new_n7543 , new_n7229 , new_n7359 );
  nand g07167 ( new_n7544 , new_n7542 , new_n7543 );
  xor  g07168 ( new_n7545 , new_n7541 , new_n7544 );
  nand g07169 ( new_n7546 , pi104 , pi145 );
  nand g07170 ( new_n7547 , pi212 , pi246 );
  and  g07171 ( new_n7548 , new_n7546 , new_n7547 );
  nand g07172 ( new_n7549 , pi104 , pi246 );
  nor  g07173 ( new_n7550 , new_n7361 , new_n7549 );
  or   g07174 ( new_n7551 , new_n7548 , new_n7550 );
  xnor g07175 ( new_n7552 , new_n7545 , new_n7551 );
  nand g07176 ( new_n7553 , new_n7361 , new_n7364 );
  nand g07177 ( new_n7554 , new_n7360 , new_n7365 );
  nand g07178 ( new_n7555 , new_n7553 , new_n7554 );
  xor  g07179 ( new_n7556 , new_n7552 , new_n7555 );
  nor  g07180 ( new_n7557 , new_n7366 , new_n7367 );
  nor  g07181 ( new_n7558 , new_n7368 , new_n7371 );
  nor  g07182 ( new_n7559 , new_n7557 , new_n7558 );
  xor  g07183 ( new_n7560 , new_n7556 , new_n7559 );
  nand g07184 ( new_n7561 , new_n7356 , new_n7372 );
  nand g07185 ( new_n7562 , pi114 , pi213 );
  xor  g07186 ( new_n7563 , new_n7561 , new_n7562 );
  xor  g07187 ( new_n7564 , new_n7560 , new_n7563 );
  nand g07188 ( new_n7565 , pi008 , pi141 );
  nand g07189 ( new_n7566 , pi026 , pi090 );
  nand g07190 ( new_n7567 , pi027 , pi047 );
  nand g07191 ( new_n7568 , new_n7566 , new_n7567 );
  nand g07192 ( new_n7569 , pi026 , pi047 );
  or   g07193 ( new_n7570 , new_n7397 , new_n7569 );
  nand g07194 ( new_n7571 , new_n7568 , new_n7570 );
  xor  g07195 ( new_n7572 , new_n7565 , new_n7571 );
  nand g07196 ( new_n7573 , new_n7397 , new_n7398 );
  nand g07197 ( new_n7574 , new_n7396 , new_n7399 );
  nand g07198 ( new_n7575 , new_n7573 , new_n7574 );
  xor  g07199 ( new_n7576 , new_n7572 , new_n7575 );
  nand g07200 ( new_n7577 , pi136 , pi241 );
  nand g07201 ( new_n7578 , pi056 , pi161 );
  and  g07202 ( new_n7579 , new_n7577 , new_n7578 );
  nand g07203 ( new_n7580 , pi136 , pi161 );
  nor  g07204 ( new_n7581 , new_n7401 , new_n7580 );
  or   g07205 ( new_n7582 , new_n7579 , new_n7581 );
  xnor g07206 ( new_n7583 , new_n7576 , new_n7582 );
  nand g07207 ( new_n7584 , new_n7401 , new_n7404 );
  nand g07208 ( new_n7585 , new_n7400 , new_n7405 );
  nand g07209 ( new_n7586 , new_n7584 , new_n7585 );
  xor  g07210 ( new_n7587 , new_n7583 , new_n7586 );
  or   g07211 ( new_n7588 , new_n7406 , new_n7407 );
  nand g07212 ( new_n7589 , new_n7408 , new_n7412 );
  nand g07213 ( new_n7590 , new_n7588 , new_n7589 );
  xnor g07214 ( new_n7591 , new_n7587 , new_n7590 );
  nand g07215 ( new_n7592 , new_n7395 , new_n7413 );
  nand g07216 ( new_n7593 , pi096 , pi236 );
  xor  g07217 ( new_n7594 , new_n7592 , new_n7593 );
  xor  g07218 ( new_n7595 , new_n7591 , new_n7594 );
  xnor g07219 ( new_n7596 , new_n7564 , new_n7595 );
  nand g07220 ( new_n7597 , new_n7414 , new_n7439 );
  nand g07221 ( new_n7598 , new_n7373 , new_n7440 );
  nand g07222 ( new_n7599 , new_n7597 , new_n7598 );
  xnor g07223 ( new_n7600 , new_n7596 , new_n7599 );
  nand g07224 ( new_n7601 , new_n7469 , new_n7472 );
  nand g07225 ( new_n7602 , new_n7468 , new_n7473 );
  nand g07226 ( new_n7603 , new_n7601 , new_n7602 );
  nand g07227 ( new_n7604 , pi019 , pi035 );
  nand g07228 ( new_n7605 , new_n7465 , new_n7466 );
  nand g07229 ( new_n7606 , new_n7464 , new_n7467 );
  nand g07230 ( new_n7607 , new_n7605 , new_n7606 );
  xor  g07231 ( new_n7608 , new_n7604 , new_n7607 );
  nand g07232 ( new_n7609 , pi015 , pi151 );
  nand g07233 ( new_n7610 , pi147 , pi204 );
  nand g07234 ( new_n7611 , new_n7609 , new_n7610 );
  nand g07235 ( new_n7612 , pi151 , pi204 );
  nor  g07236 ( new_n7613 , new_n7466 , new_n7612 );
  not  g07237 ( new_n7614 , new_n7613 );
  nand g07238 ( new_n7615 , new_n7611 , new_n7614 );
  xor  g07239 ( new_n7616 , new_n7608 , new_n7615 );
  nand g07240 ( new_n7617 , pi097 , pi139 );
  nand g07241 ( new_n7618 , pi075 , pi208 );
  nand g07242 ( new_n7619 , new_n7617 , new_n7618 );
  nand g07243 ( new_n7620 , pi075 , pi139 );
  or   g07244 ( new_n7621 , new_n7469 , new_n7620 );
  nand g07245 ( new_n7622 , new_n7619 , new_n7621 );
  xor  g07246 ( new_n7623 , new_n7616 , new_n7622 );
  xor  g07247 ( new_n7624 , new_n7603 , new_n7623 );
  not  g07248 ( new_n7625 , new_n7475 );
  nand g07249 ( new_n7626 , new_n7625 , new_n7478 );
  or   g07250 ( new_n7627 , new_n7474 , new_n7479 );
  nand g07251 ( new_n7628 , new_n7626 , new_n7627 );
  xor  g07252 ( new_n7629 , new_n7624 , new_n7628 );
  nand g07253 ( new_n7630 , new_n7463 , new_n7480 );
  nand g07254 ( new_n7631 , pi093 , pi168 );
  xor  g07255 ( new_n7632 , new_n7630 , new_n7631 );
  xor  g07256 ( new_n7633 , new_n7629 , new_n7632 );
  xor  g07257 ( new_n7634 , new_n7600 , new_n7633 );
  nand g07258 ( new_n7635 , new_n7441 , new_n7482 );
  nand g07259 ( new_n7636 , new_n7483 , new_n7507 );
  nand g07260 ( new_n7637 , new_n7635 , new_n7636 );
  xnor g07261 ( new_n7638 , new_n7634 , new_n7637 );
  xor  g07262 ( new_n7639 , new_n7335 , new_n7534 );
  nand g07263 ( new_n7640 , new_n7638 , new_n7639 );
  nand g07264 ( new_n7641 , new_n7535 , new_n7640 );
  nand g07265 ( new_n7642 , new_n7323 , new_n7333 );
  not  g07266 ( new_n7643 , new_n7322 );
  nand g07267 ( new_n7644 , new_n7643 , new_n7334 );
  nand g07268 ( new_n7645 , new_n7642 , new_n7644 );
  nand g07269 ( new_n7646 , new_n7302 , new_n7321 );
  xor  g07270 ( new_n7647 , new_n7294 , new_n7297 );
  xor  g07271 ( new_n7648 , new_n7646 , new_n7647 );
  xnor g07272 ( new_n7649 , new_n7645 , new_n7648 );
  or   g07273 ( new_n7650 , new_n7641 , new_n7649 );
  not  g07274 ( new_n7651 , new_n7559 );
  nand g07275 ( new_n7652 , new_n7556 , new_n7651 );
  xor  g07276 ( new_n7653 , new_n7236 , new_n7238 );
  nand g07277 ( new_n7654 , pi114 , pi212 );
  nand g07278 ( new_n7655 , pi091 , pi213 );
  xor  g07279 ( new_n7656 , new_n7654 , new_n7655 );
  xor  g07280 ( new_n7657 , new_n7549 , new_n7656 );
  nand g07281 ( new_n7658 , new_n7536 , new_n7540 );
  nand g07282 ( new_n7659 , new_n7541 , new_n7544 );
  nand g07283 ( new_n7660 , new_n7658 , new_n7659 );
  xor  g07284 ( new_n7661 , new_n7657 , new_n7660 );
  xnor g07285 ( new_n7662 , new_n7653 , new_n7661 );
  nor  g07286 ( new_n7663 , new_n7545 , new_n7551 );
  nor  g07287 ( new_n7664 , new_n7552 , new_n7555 );
  xor  g07288 ( new_n7665 , new_n7550 , new_n7664 );
  nor  g07289 ( new_n7666 , new_n7663 , new_n7665 );
  xor  g07290 ( new_n7667 , new_n7662 , new_n7666 );
  xnor g07291 ( new_n7668 , new_n7652 , new_n7667 );
  nand g07292 ( new_n7669 , new_n7561 , new_n7562 );
  nand g07293 ( new_n7670 , new_n7560 , new_n7563 );
  nand g07294 ( new_n7671 , new_n7669 , new_n7670 );
  xnor g07295 ( new_n7672 , new_n7668 , new_n7671 );
  nand g07296 ( new_n7673 , new_n7587 , new_n7590 );
  nand g07297 ( new_n7674 , pi018 , pi027 );
  nand g07298 ( new_n7675 , pi008 , pi090 );
  xor  g07299 ( new_n7676 , new_n7674 , new_n7675 );
  xor  g07300 ( new_n7677 , new_n7569 , new_n7676 );
  nand g07301 ( new_n7678 , pi056 , pi141 );
  xor  g07302 ( new_n7679 , new_n7570 , new_n7678 );
  xor  g07303 ( new_n7680 , new_n7677 , new_n7679 );
  nand g07304 ( new_n7681 , pi096 , pi241 );
  nand g07305 ( new_n7682 , pi235 , pi236 );
  xor  g07306 ( new_n7683 , new_n7681 , new_n7682 );
  xor  g07307 ( new_n7684 , new_n7580 , new_n7683 );
  nand g07308 ( new_n7685 , new_n7565 , new_n7571 );
  nand g07309 ( new_n7686 , new_n7572 , new_n7575 );
  nand g07310 ( new_n7687 , new_n7685 , new_n7686 );
  xor  g07311 ( new_n7688 , new_n7684 , new_n7687 );
  xnor g07312 ( new_n7689 , new_n7680 , new_n7688 );
  nor  g07313 ( new_n7690 , new_n7576 , new_n7582 );
  nor  g07314 ( new_n7691 , new_n7583 , new_n7586 );
  xor  g07315 ( new_n7692 , new_n7581 , new_n7691 );
  nor  g07316 ( new_n7693 , new_n7690 , new_n7692 );
  xor  g07317 ( new_n7694 , new_n7689 , new_n7693 );
  xnor g07318 ( new_n7695 , new_n7673 , new_n7694 );
  nand g07319 ( new_n7696 , new_n7592 , new_n7593 );
  nand g07320 ( new_n7697 , new_n7591 , new_n7594 );
  nand g07321 ( new_n7698 , new_n7696 , new_n7697 );
  xor  g07322 ( new_n7699 , new_n7695 , new_n7698 );
  not  g07323 ( new_n7700 , new_n7699 );
  xor  g07324 ( new_n7701 , new_n7672 , new_n7700 );
  nor  g07325 ( new_n7702 , new_n7564 , new_n7595 );
  nor  g07326 ( new_n7703 , new_n7596 , new_n7599 );
  nor  g07327 ( new_n7704 , new_n7702 , new_n7703 );
  xor  g07328 ( new_n7705 , new_n7701 , new_n7704 );
  not  g07329 ( new_n7706 , new_n7624 );
  nand g07330 ( new_n7707 , new_n7706 , new_n7628 );
  nand g07331 ( new_n7708 , pi146 , pi147 );
  nand g07332 ( new_n7709 , pi015 , pi019 );
  xor  g07333 ( new_n7710 , new_n7708 , new_n7709 );
  xor  g07334 ( new_n7711 , new_n7612 , new_n7710 );
  nand g07335 ( new_n7712 , pi035 , pi097 );
  xor  g07336 ( new_n7713 , new_n7614 , new_n7712 );
  not  g07337 ( new_n7714 , new_n7713 );
  xor  g07338 ( new_n7715 , new_n7711 , new_n7714 );
  nand g07339 ( new_n7716 , pi093 , pi208 );
  nand g07340 ( new_n7717 , pi166 , pi168 );
  xor  g07341 ( new_n7718 , new_n7716 , new_n7717 );
  xor  g07342 ( new_n7719 , new_n7620 , new_n7718 );
  nand g07343 ( new_n7720 , new_n7604 , new_n7607 );
  nand g07344 ( new_n7721 , new_n7608 , new_n7615 );
  nand g07345 ( new_n7722 , new_n7720 , new_n7721 );
  xor  g07346 ( new_n7723 , new_n7719 , new_n7722 );
  xor  g07347 ( new_n7724 , new_n7715 , new_n7723 );
  nand g07348 ( new_n7725 , new_n7616 , new_n7622 );
  nand g07349 ( new_n7726 , new_n7603 , new_n7623 );
  nand g07350 ( new_n7727 , new_n7725 , new_n7726 );
  xor  g07351 ( new_n7728 , new_n7621 , new_n7727 );
  xnor g07352 ( new_n7729 , new_n7724 , new_n7728 );
  xnor g07353 ( new_n7730 , new_n7707 , new_n7729 );
  nand g07354 ( new_n7731 , new_n7630 , new_n7631 );
  nand g07355 ( new_n7732 , new_n7629 , new_n7632 );
  nand g07356 ( new_n7733 , new_n7731 , new_n7732 );
  xor  g07357 ( new_n7734 , new_n7730 , new_n7733 );
  not  g07358 ( new_n7735 , new_n7734 );
  xor  g07359 ( new_n7736 , new_n7705 , new_n7735 );
  nand g07360 ( new_n7737 , new_n7600 , new_n7633 );
  nand g07361 ( new_n7738 , new_n7634 , new_n7637 );
  nand g07362 ( new_n7739 , new_n7737 , new_n7738 );
  xor  g07363 ( new_n7740 , new_n7736 , new_n7739 );
  xor  g07364 ( new_n7741 , new_n7641 , new_n7649 );
  nand g07365 ( new_n7742 , new_n7740 , new_n7741 );
  nand g07366 ( new_n7743 , new_n7650 , new_n7742 );
  xor  g07367 ( new_n7744 , new_n7301 , new_n7743 );
  xor  g07368 ( new_n7745 , new_n7300 , new_n7744 );
  nand g07369 ( new_n7746 , pi009 , pi131 );
  nand g07370 ( new_n7747 , new_n7646 , new_n7647 );
  nand g07371 ( new_n7748 , new_n7645 , new_n7648 );
  nand g07372 ( new_n7749 , new_n7747 , new_n7748 );
  nand g07373 ( new_n7750 , pi034 , pi119 );
  xor  g07374 ( new_n7751 , new_n7749 , new_n7750 );
  xor  g07375 ( new_n7752 , new_n7746 , new_n7751 );
  nand g07376 ( new_n7753 , new_n7674 , new_n7675 );
  nand g07377 ( new_n7754 , new_n7569 , new_n7676 );
  nand g07378 ( new_n7755 , new_n7753 , new_n7754 );
  or   g07379 ( new_n7756 , new_n7570 , new_n7678 );
  not  g07380 ( new_n7757 , new_n7677 );
  nand g07381 ( new_n7758 , new_n7757 , new_n7679 );
  nand g07382 ( new_n7759 , new_n7756 , new_n7758 );
  nand g07383 ( new_n7760 , new_n7684 , new_n7687 );
  nand g07384 ( new_n7761 , new_n7680 , new_n7688 );
  nand g07385 ( new_n7762 , new_n7760 , new_n7761 );
  nand g07386 ( new_n7763 , new_n7681 , new_n7682 );
  nand g07387 ( new_n7764 , new_n7580 , new_n7683 );
  nand g07388 ( new_n7765 , new_n7763 , new_n7764 );
  xor  g07389 ( new_n7766 , new_n7762 , new_n7765 );
  nand g07390 ( new_n7767 , pi096 , pi161 );
  xor  g07391 ( new_n7768 , new_n7766 , new_n7767 );
  xor  g07392 ( new_n7769 , new_n7759 , new_n7768 );
  xor  g07393 ( new_n7770 , new_n7755 , new_n7769 );
  xor  g07394 ( new_n7771 , new_n7752 , new_n7770 );
  xor  g07395 ( new_n7772 , new_n7745 , new_n7771 );
  xor  g07396 ( new_n7773 , new_n7240 , new_n7772 );
  nand g07397 ( new_n7774 , new_n7654 , new_n7655 );
  nand g07398 ( new_n7775 , new_n7549 , new_n7656 );
  nand g07399 ( new_n7776 , new_n7774 , new_n7775 );
  nor  g07400 ( new_n7777 , new_n7673 , new_n7694 );
  nor  g07401 ( new_n7778 , new_n7695 , new_n7698 );
  nor  g07402 ( new_n7779 , new_n7777 , new_n7778 );
  xor  g07403 ( new_n7780 , new_n7776 , new_n7779 );
  nand g07404 ( new_n7781 , pi091 , pi212 );
  nand g07405 ( new_n7782 , pi104 , pi114 );
  xor  g07406 ( new_n7783 , new_n7781 , new_n7782 );
  nand g07407 ( new_n7784 , new_n7581 , new_n7691 );
  not  g07408 ( new_n7785 , new_n7693 );
  nand g07409 ( new_n7786 , new_n7689 , new_n7785 );
  nand g07410 ( new_n7787 , new_n7784 , new_n7786 );
  nand g07411 ( new_n7788 , pi056 , pi090 );
  nand g07412 ( new_n7789 , pi136 , pi141 );
  xor  g07413 ( new_n7790 , new_n7788 , new_n7789 );
  xor  g07414 ( new_n7791 , new_n7787 , new_n7790 );
  nand g07415 ( new_n7792 , pi008 , pi047 );
  nand g07416 ( new_n7793 , pi110 , pi236 );
  nand g07417 ( new_n7794 , pi018 , pi026 );
  nand g07418 ( new_n7795 , pi027 , pi128 );
  xor  g07419 ( new_n7796 , new_n7794 , new_n7795 );
  xor  g07420 ( new_n7797 , new_n7793 , new_n7796 );
  xor  g07421 ( new_n7798 , new_n7792 , new_n7797 );
  xor  g07422 ( new_n7799 , new_n7791 , new_n7798 );
  xor  g07423 ( new_n7800 , new_n7783 , new_n7799 );
  xor  g07424 ( new_n7801 , new_n7780 , new_n7800 );
  nand g07425 ( new_n7802 , pi088 , pi164 );
  nand g07426 ( new_n7803 , pi183 , pi206 );
  nand g07427 ( new_n7804 , pi032 , pi105 );
  xor  g07428 ( new_n7805 , new_n7803 , new_n7804 );
  nand g07429 ( new_n7806 , pi031 , pi213 );
  nand g07430 ( new_n7807 , new_n7672 , new_n7700 );
  nand g07431 ( new_n7808 , new_n7701 , new_n7704 );
  nand g07432 ( new_n7809 , new_n7807 , new_n7808 );
  xor  g07433 ( new_n7810 , new_n7806 , new_n7809 );
  xor  g07434 ( new_n7811 , new_n7805 , new_n7810 );
  xor  g07435 ( new_n7812 , new_n7802 , new_n7811 );
  nand g07436 ( new_n7813 , pi035 , pi075 );
  nand g07437 ( new_n7814 , pi093 , pi139 );
  xor  g07438 ( new_n7815 , new_n7813 , new_n7814 );
  nand g07439 ( new_n7816 , pi019 , pi204 );
  xor  g07440 ( new_n7817 , new_n7815 , new_n7816 );
  nand g07441 ( new_n7818 , pi166 , pi208 );
  nand g07442 ( new_n7819 , new_n7708 , new_n7709 );
  nand g07443 ( new_n7820 , new_n7612 , new_n7710 );
  nand g07444 ( new_n7821 , new_n7819 , new_n7820 );
  nor  g07445 ( new_n7822 , new_n7614 , new_n7712 );
  nor  g07446 ( new_n7823 , new_n7711 , new_n7714 );
  or   g07447 ( new_n7824 , new_n7822 , new_n7823 );
  xor  g07448 ( new_n7825 , new_n7821 , new_n7824 );
  xor  g07449 ( new_n7826 , new_n7818 , new_n7825 );
  xor  g07450 ( new_n7827 , new_n7817 , new_n7826 );
  xor  g07451 ( new_n7828 , new_n7812 , new_n7827 );
  nand g07452 ( new_n7829 , new_n7550 , new_n7664 );
  not  g07453 ( new_n7830 , new_n7666 );
  nand g07454 ( new_n7831 , new_n7662 , new_n7830 );
  nand g07455 ( new_n7832 , new_n7829 , new_n7831 );
  nor  g07456 ( new_n7833 , new_n7652 , new_n7667 );
  nor  g07457 ( new_n7834 , new_n7668 , new_n7671 );
  or   g07458 ( new_n7835 , new_n7833 , new_n7834 );
  xor  g07459 ( new_n7836 , new_n7832 , new_n7835 );
  nand g07460 ( new_n7837 , new_n7716 , new_n7717 );
  nand g07461 ( new_n7838 , new_n7620 , new_n7718 );
  nand g07462 ( new_n7839 , new_n7837 , new_n7838 );
  nand g07463 ( new_n7840 , pi015 , pi097 );
  nand g07464 ( new_n7841 , new_n7719 , new_n7722 );
  not  g07465 ( new_n7842 , new_n7715 );
  nand g07466 ( new_n7843 , new_n7842 , new_n7723 );
  nand g07467 ( new_n7844 , new_n7841 , new_n7843 );
  xor  g07468 ( new_n7845 , new_n7840 , new_n7844 );
  xor  g07469 ( new_n7846 , new_n7839 , new_n7845 );
  xor  g07470 ( new_n7847 , new_n7836 , new_n7846 );
  xor  g07471 ( new_n7848 , new_n7828 , new_n7847 );
  nand g07472 ( new_n7849 , pi045 , pi084 );
  nand g07473 ( new_n7850 , pi052 , pi248 );
  nand g07474 ( new_n7851 , pi072 , pi077 );
  xor  g07475 ( new_n7852 , new_n7850 , new_n7851 );
  xor  g07476 ( new_n7853 , new_n7849 , new_n7852 );
  xor  g07477 ( new_n7854 , new_n7848 , new_n7853 );
  nand g07478 ( new_n7855 , new_n7289 , new_n7292 );
  nand g07479 ( new_n7856 , new_n7285 , new_n7293 );
  nand g07480 ( new_n7857 , new_n7855 , new_n7856 );
  nand g07481 ( new_n7858 , new_n7286 , new_n7287 );
  nand g07482 ( new_n7859 , new_n7241 , new_n7288 );
  nand g07483 ( new_n7860 , new_n7858 , new_n7859 );
  xor  g07484 ( new_n7861 , new_n7857 , new_n7860 );
  nand g07485 ( new_n7862 , pi044 , pi189 );
  nand g07486 ( new_n7863 , pi054 , pi133 );
  xor  g07487 ( new_n7864 , new_n7862 , new_n7863 );
  xor  g07488 ( new_n7865 , new_n7861 , new_n7864 );
  nor  g07489 ( new_n7866 , new_n7707 , new_n7729 );
  nor  g07490 ( new_n7867 , new_n7730 , new_n7733 );
  nor  g07491 ( new_n7868 , new_n7866 , new_n7867 );
  nand g07492 ( new_n7869 , pi064 , pi250 );
  xor  g07493 ( new_n7870 , new_n7868 , new_n7869 );
  xor  g07494 ( new_n7871 , new_n7865 , new_n7870 );
  or   g07495 ( new_n7872 , new_n7621 , new_n7727 );
  nand g07496 ( new_n7873 , new_n7724 , new_n7728 );
  nand g07497 ( new_n7874 , new_n7872 , new_n7873 );
  nand g07498 ( new_n7875 , pi011 , pi168 );
  xor  g07499 ( new_n7876 , new_n7874 , new_n7875 );
  nand g07500 ( new_n7877 , pi147 , pi152 );
  nand g07501 ( new_n7878 , pi146 , pi151 );
  xor  g07502 ( new_n7879 , new_n7877 , new_n7878 );
  xor  g07503 ( new_n7880 , new_n7876 , new_n7879 );
  nand g07504 ( new_n7881 , new_n7279 , new_n7280 );
  nand g07505 ( new_n7882 , new_n7249 , new_n7281 );
  nand g07506 ( new_n7883 , new_n7881 , new_n7882 );
  or   g07507 ( new_n7884 , new_n7250 , new_n7283 );
  not  g07508 ( new_n7885 , new_n7282 );
  nand g07509 ( new_n7886 , new_n7885 , new_n7284 );
  nand g07510 ( new_n7887 , new_n7884 , new_n7886 );
  xor  g07511 ( new_n7888 , new_n7883 , new_n7887 );
  xor  g07512 ( new_n7889 , new_n7880 , new_n7888 );
  xor  g07513 ( new_n7890 , new_n7871 , new_n7889 );
  xor  g07514 ( new_n7891 , new_n7854 , new_n7890 );
  nand g07515 ( new_n7892 , pi013 , pi246 );
  nand g07516 ( new_n7893 , new_n7657 , new_n7660 );
  nand g07517 ( new_n7894 , new_n7653 , new_n7661 );
  nand g07518 ( new_n7895 , new_n7893 , new_n7894 );
  xor  g07519 ( new_n7896 , new_n7892 , new_n7895 );
  nand g07520 ( new_n7897 , pi112 , pi145 );
  xor  g07521 ( new_n7898 , new_n7896 , new_n7897 );
  xor  g07522 ( new_n7899 , new_n7891 , new_n7898 );
  xor  g07523 ( new_n7900 , new_n7801 , new_n7899 );
  nand g07524 ( new_n7901 , new_n7705 , new_n7735 );
  nand g07525 ( new_n7902 , new_n7736 , new_n7739 );
  nand g07526 ( new_n7903 , new_n7901 , new_n7902 );
  nand g07527 ( new_n7904 , new_n7233 , new_n7234 );
  nand g07528 ( new_n7905 , new_n7230 , new_n7235 );
  nand g07529 ( new_n7906 , new_n7904 , new_n7905 );
  xor  g07530 ( new_n7907 , new_n7903 , new_n7906 );
  xor  g07531 ( new_n7908 , new_n7900 , new_n7907 );
  xor  g07532 ( po039 , new_n7773 , new_n7908 );
  xor  g07533 ( po040 , new_n7638 , new_n7639 );
  nand g07534 ( new_n7911 , pi066 , pi163 );
  xor  g07535 ( new_n7912 , new_n4966 , new_n7911 );
  nand g07536 ( new_n7913 , pi226 , pi228 );
  xor  g07537 ( new_n7914 , new_n7912 , new_n7913 );
  or   g07538 ( new_n7915 , new_n4968 , new_n7914 );
  nand g07539 ( new_n7916 , pi207 , pi228 );
  nand g07540 ( new_n7917 , pi066 , pi148 );
  nand g07541 ( new_n7918 , pi039 , pi226 );
  xor  g07542 ( new_n7919 , new_n7917 , new_n7918 );
  xor  g07543 ( new_n7920 , new_n7916 , new_n7919 );
  nand g07544 ( new_n7921 , pi055 , pi163 );
  nand g07545 ( new_n7922 , new_n4966 , new_n7911 );
  nand g07546 ( new_n7923 , new_n7912 , new_n7913 );
  nand g07547 ( new_n7924 , new_n7922 , new_n7923 );
  xor  g07548 ( new_n7925 , new_n7921 , new_n7924 );
  xor  g07549 ( new_n7926 , new_n7920 , new_n7925 );
  or   g07550 ( new_n7927 , new_n7915 , new_n7926 );
  nand g07551 ( new_n7928 , pi002 , pi163 );
  nand g07552 ( new_n7929 , new_n7921 , new_n7924 );
  nand g07553 ( new_n7930 , new_n7920 , new_n7925 );
  nand g07554 ( new_n7931 , new_n7929 , new_n7930 );
  xor  g07555 ( new_n7932 , new_n7928 , new_n7931 );
  nand g07556 ( new_n7933 , pi116 , pi226 );
  nand g07557 ( new_n7934 , pi066 , pi228 );
  nand g07558 ( new_n7935 , pi039 , pi207 );
  xor  g07559 ( new_n7936 , new_n7934 , new_n7935 );
  xor  g07560 ( new_n7937 , new_n7933 , new_n7936 );
  nand g07561 ( new_n7938 , pi055 , pi148 );
  nand g07562 ( new_n7939 , new_n7917 , new_n7918 );
  nand g07563 ( new_n7940 , new_n7916 , new_n7919 );
  nand g07564 ( new_n7941 , new_n7939 , new_n7940 );
  xor  g07565 ( new_n7942 , new_n7938 , new_n7941 );
  xnor g07566 ( new_n7943 , new_n7937 , new_n7942 );
  xnor g07567 ( new_n7944 , new_n7932 , new_n7943 );
  xor  g07568 ( new_n7945 , new_n7927 , new_n7944 );
  nand g07569 ( new_n7946 , pi107 , pi173 );
  xor  g07570 ( new_n7947 , new_n4974 , new_n7946 );
  nand g07571 ( new_n7948 , pi049 , pi109 );
  xor  g07572 ( new_n7949 , new_n7947 , new_n7948 );
  or   g07573 ( new_n7950 , new_n4976 , new_n7949 );
  nand g07574 ( new_n7951 , pi171 , pi173 );
  nand g07575 ( new_n7952 , pi109 , pi245 );
  nand g07576 ( new_n7953 , pi014 , pi049 );
  xor  g07577 ( new_n7954 , new_n7952 , new_n7953 );
  xor  g07578 ( new_n7955 , new_n7951 , new_n7954 );
  nand g07579 ( new_n7956 , pi107 , pi230 );
  nand g07580 ( new_n7957 , new_n4974 , new_n7946 );
  nand g07581 ( new_n7958 , new_n7947 , new_n7948 );
  nand g07582 ( new_n7959 , new_n7957 , new_n7958 );
  xor  g07583 ( new_n7960 , new_n7956 , new_n7959 );
  xor  g07584 ( new_n7961 , new_n7955 , new_n7960 );
  nor  g07585 ( new_n7962 , new_n7950 , new_n7961 );
  nand g07586 ( new_n7963 , pi049 , pi173 );
  nand g07587 ( new_n7964 , pi014 , pi245 );
  nand g07588 ( new_n7965 , pi109 , pi201 );
  xor  g07589 ( new_n7966 , new_n7964 , new_n7965 );
  xor  g07590 ( new_n7967 , new_n7963 , new_n7966 );
  nand g07591 ( new_n7968 , pi171 , pi230 );
  nand g07592 ( new_n7969 , new_n7952 , new_n7953 );
  nand g07593 ( new_n7970 , new_n7951 , new_n7954 );
  nand g07594 ( new_n7971 , new_n7969 , new_n7970 );
  xor  g07595 ( new_n7972 , new_n7968 , new_n7971 );
  xnor g07596 ( new_n7973 , new_n7967 , new_n7972 );
  nand g07597 ( new_n7974 , pi050 , pi107 );
  nand g07598 ( new_n7975 , new_n7956 , new_n7959 );
  nand g07599 ( new_n7976 , new_n7955 , new_n7960 );
  nand g07600 ( new_n7977 , new_n7975 , new_n7976 );
  xor  g07601 ( new_n7978 , new_n7974 , new_n7977 );
  xor  g07602 ( new_n7979 , new_n7973 , new_n7978 );
  xor  g07603 ( new_n7980 , new_n7962 , new_n7979 );
  xor  g07604 ( new_n7981 , new_n7945 , new_n7980 );
  xor  g07605 ( new_n7982 , new_n7950 , new_n7961 );
  xor  g07606 ( new_n7983 , new_n7915 , new_n7926 );
  nand g07607 ( new_n7984 , new_n7982 , new_n7983 );
  not  g07608 ( new_n7985 , new_n7984 );
  xnor g07609 ( new_n7986 , new_n7982 , new_n7983 );
  xor  g07610 ( new_n7987 , new_n4975 , new_n7949 );
  not  g07611 ( new_n7988 , new_n4962 );
  nor  g07612 ( new_n7989 , new_n7988 , new_n4969 );
  nor  g07613 ( new_n7990 , new_n4970 , new_n4977 );
  nor  g07614 ( new_n7991 , new_n7989 , new_n7990 );
  nand g07615 ( new_n7992 , new_n7987 , new_n7991 );
  xor  g07616 ( new_n7993 , new_n4968 , new_n7914 );
  not  g07617 ( new_n7994 , new_n7993 );
  xor  g07618 ( new_n7995 , new_n7987 , new_n7991 );
  nand g07619 ( new_n7996 , new_n7994 , new_n7995 );
  nand g07620 ( new_n7997 , new_n7992 , new_n7996 );
  nor  g07621 ( new_n7998 , new_n7986 , new_n7997 );
  nor  g07622 ( new_n7999 , new_n7985 , new_n7998 );
  not  g07623 ( new_n8000 , new_n7999 );
  xor  g07624 ( new_n8001 , new_n7981 , new_n8000 );
  nand g07625 ( new_n8002 , pi058 , pi175 );
  xor  g07626 ( new_n8003 , new_n4986 , new_n8002 );
  nand g07627 ( new_n8004 , pi132 , pi240 );
  xor  g07628 ( new_n8005 , new_n8003 , new_n8004 );
  not  g07629 ( new_n8006 , new_n8005 );
  nand g07630 ( new_n8007 , new_n4987 , new_n8006 );
  nand g07631 ( new_n8008 , pi175 , pi211 );
  nand g07632 ( new_n8009 , new_n4986 , new_n8002 );
  nand g07633 ( new_n8010 , new_n8003 , new_n8004 );
  nand g07634 ( new_n8011 , new_n8009 , new_n8010 );
  xor  g07635 ( new_n8012 , new_n8008 , new_n8011 );
  nand g07636 ( new_n8013 , pi058 , pi134 );
  nand g07637 ( new_n8014 , pi132 , pi149 );
  nand g07638 ( new_n8015 , pi186 , pi240 );
  xor  g07639 ( new_n8016 , new_n8014 , new_n8015 );
  xor  g07640 ( new_n8017 , new_n8013 , new_n8016 );
  xor  g07641 ( new_n8018 , new_n8012 , new_n8017 );
  nor  g07642 ( new_n8019 , new_n8007 , new_n8018 );
  nand g07643 ( new_n8020 , pi058 , pi240 );
  nand g07644 ( new_n8021 , pi149 , pi186 );
  nand g07645 ( new_n8022 , pi132 , pi167 );
  xor  g07646 ( new_n8023 , new_n8021 , new_n8022 );
  xor  g07647 ( new_n8024 , new_n8020 , new_n8023 );
  nand g07648 ( new_n8025 , pi134 , pi211 );
  nand g07649 ( new_n8026 , new_n8014 , new_n8015 );
  nand g07650 ( new_n8027 , new_n8013 , new_n8016 );
  nand g07651 ( new_n8028 , new_n8026 , new_n8027 );
  xor  g07652 ( new_n8029 , new_n8025 , new_n8028 );
  xor  g07653 ( new_n8030 , new_n8024 , new_n8029 );
  nand g07654 ( new_n8031 , pi175 , pi199 );
  or   g07655 ( new_n8032 , new_n8008 , new_n8011 );
  not  g07656 ( new_n8033 , new_n8017 );
  nand g07657 ( new_n8034 , new_n8012 , new_n8033 );
  nand g07658 ( new_n8035 , new_n8032 , new_n8034 );
  xor  g07659 ( new_n8036 , new_n8031 , new_n8035 );
  xor  g07660 ( new_n8037 , new_n8030 , new_n8036 );
  xor  g07661 ( new_n8038 , new_n8019 , new_n8037 );
  xor  g07662 ( new_n8039 , new_n8001 , new_n8038 );
  xor  g07663 ( new_n8040 , new_n7986 , new_n7997 );
  xor  g07664 ( new_n8041 , new_n8007 , new_n8018 );
  nand g07665 ( new_n8042 , new_n8040 , new_n8041 );
  xor  g07666 ( new_n8043 , new_n8040 , new_n8041 );
  xor  g07667 ( new_n8044 , new_n4987 , new_n8005 );
  nand g07668 ( new_n8045 , new_n4982 , new_n4988 );
  not  g07669 ( new_n8046 , new_n4978 );
  nand g07670 ( new_n8047 , new_n8046 , new_n4989 );
  nand g07671 ( new_n8048 , new_n8045 , new_n8047 );
  or   g07672 ( new_n8049 , new_n8044 , new_n8048 );
  xor  g07673 ( new_n8050 , new_n7993 , new_n7995 );
  xor  g07674 ( new_n8051 , new_n8044 , new_n8048 );
  nand g07675 ( new_n8052 , new_n8050 , new_n8051 );
  nand g07676 ( new_n8053 , new_n8049 , new_n8052 );
  nand g07677 ( new_n8054 , new_n8043 , new_n8053 );
  nand g07678 ( new_n8055 , new_n8042 , new_n8054 );
  xor  g07679 ( new_n8056 , new_n8039 , new_n8055 );
  nand g07680 ( new_n8057 , pi103 , pi150 );
  nand g07681 ( new_n8058 , pi103 , pi244 );
  nand g07682 ( new_n8059 , pi016 , pi029 );
  nand g07683 ( new_n8060 , new_n8058 , new_n8059 );
  nand g07684 ( new_n8061 , pi069 , pi117 );
  or   g07685 ( new_n8062 , new_n8058 , new_n8059 );
  nand g07686 ( new_n8063 , new_n8061 , new_n8062 );
  nand g07687 ( new_n8064 , new_n8060 , new_n8063 );
  xor  g07688 ( new_n8065 , new_n8057 , new_n8064 );
  nand g07689 ( new_n8066 , pi016 , pi069 );
  nand g07690 ( new_n8067 , pi029 , pi080 );
  nand g07691 ( new_n8068 , pi117 , pi244 );
  xor  g07692 ( new_n8069 , new_n8067 , new_n8068 );
  xor  g07693 ( new_n8070 , new_n8066 , new_n8069 );
  xor  g07694 ( new_n8071 , new_n8065 , new_n8070 );
  not  g07695 ( new_n8072 , new_n8061 );
  not  g07696 ( new_n8073 , new_n8060 );
  nand g07697 ( new_n8074 , new_n4992 , new_n8072 );
  nand g07698 ( new_n8075 , new_n8073 , new_n8074 );
  nand g07699 ( new_n8076 , new_n8062 , new_n8075 );
  nand g07700 ( new_n8077 , new_n8072 , new_n8076 );
  nor  g07701 ( new_n8078 , new_n8071 , new_n8077 );
  nand g07702 ( new_n8079 , pi016 , pi244 );
  nand g07703 ( new_n8080 , pi069 , pi080 );
  nand g07704 ( new_n8081 , pi029 , pi247 );
  xor  g07705 ( new_n8082 , new_n8080 , new_n8081 );
  xor  g07706 ( new_n8083 , new_n8079 , new_n8082 );
  nand g07707 ( new_n8084 , pi117 , pi150 );
  nand g07708 ( new_n8085 , new_n8067 , new_n8068 );
  nand g07709 ( new_n8086 , new_n8066 , new_n8069 );
  nand g07710 ( new_n8087 , new_n8085 , new_n8086 );
  xor  g07711 ( new_n8088 , new_n8084 , new_n8087 );
  xnor g07712 ( new_n8089 , new_n8083 , new_n8088 );
  nand g07713 ( new_n8090 , pi103 , pi221 );
  or   g07714 ( new_n8091 , new_n8057 , new_n8064 );
  not  g07715 ( new_n8092 , new_n8070 );
  nand g07716 ( new_n8093 , new_n8065 , new_n8092 );
  nand g07717 ( new_n8094 , new_n8091 , new_n8093 );
  xor  g07718 ( new_n8095 , new_n8090 , new_n8094 );
  xor  g07719 ( new_n8096 , new_n8089 , new_n8095 );
  xor  g07720 ( new_n8097 , new_n8078 , new_n8096 );
  xor  g07721 ( new_n8098 , new_n8071 , new_n8077 );
  nor  g07722 ( new_n8099 , new_n8073 , new_n8074 );
  nor  g07723 ( new_n8100 , new_n8076 , new_n8099 );
  nand g07724 ( new_n8101 , new_n4993 , new_n4996 );
  nand g07725 ( new_n8102 , new_n4990 , new_n4997 );
  nand g07726 ( new_n8103 , new_n8101 , new_n8102 );
  nand g07727 ( new_n8104 , new_n8100 , new_n8103 );
  xor  g07728 ( new_n8105 , new_n8050 , new_n8051 );
  xor  g07729 ( new_n8106 , new_n8100 , new_n8103 );
  nand g07730 ( new_n8107 , new_n8105 , new_n8106 );
  nand g07731 ( new_n8108 , new_n8104 , new_n8107 );
  or   g07732 ( new_n8109 , new_n8098 , new_n8108 );
  xor  g07733 ( new_n8110 , new_n8043 , new_n8053 );
  not  g07734 ( new_n8111 , new_n8110 );
  xor  g07735 ( new_n8112 , new_n8098 , new_n8108 );
  nand g07736 ( new_n8113 , new_n8111 , new_n8112 );
  nand g07737 ( new_n8114 , new_n8109 , new_n8113 );
  xor  g07738 ( new_n8115 , new_n8097 , new_n8114 );
  xor  g07739 ( po041 , new_n8056 , new_n8115 );
  xor  g07740 ( po042 , new_n6943 , new_n6945 );
  xor  g07741 ( po043 , new_n4953 , new_n4955 );
  xor  g07742 ( po044 , new_n1019 , new_n1036 );
  xor  g07743 ( po045 , new_n2543 , new_n2573 );
  xor  g07744 ( po046 , new_n4925 , new_n4941 );
  nand g07745 ( new_n8122 , pi107 , pi205 );
  nand g07746 ( new_n8123 , pi171 , pi253 );
  nand g07747 ( new_n8124 , pi074 , pi107 );
  nand g07748 ( new_n8125 , new_n8123 , new_n8124 );
  nand g07749 ( new_n8126 , pi049 , pi050 );
  xor  g07750 ( new_n8127 , new_n8123 , new_n8124 );
  nand g07751 ( new_n8128 , new_n8126 , new_n8127 );
  nand g07752 ( new_n8129 , new_n8125 , new_n8128 );
  nand g07753 ( new_n8130 , pi074 , pi171 );
  nand g07754 ( new_n8131 , pi063 , pi109 );
  nand g07755 ( new_n8132 , pi173 , pi201 );
  nand g07756 ( new_n8133 , new_n8131 , new_n8132 );
  nand g07757 ( new_n8134 , pi014 , pi156 );
  xor  g07758 ( new_n8135 , new_n8131 , new_n8132 );
  nand g07759 ( new_n8136 , new_n8134 , new_n8135 );
  nand g07760 ( new_n8137 , new_n8133 , new_n8136 );
  xor  g07761 ( new_n8138 , new_n8130 , new_n8137 );
  xor  g07762 ( new_n8139 , new_n8129 , new_n8138 );
  nand g07763 ( new_n8140 , pi029 , pi202 );
  nand g07764 ( new_n8141 , pi080 , pi244 );
  nand g07765 ( new_n8142 , new_n8080 , new_n8081 );
  nand g07766 ( new_n8143 , new_n8079 , new_n8082 );
  nand g07767 ( new_n8144 , new_n8142 , new_n8143 );
  xor  g07768 ( new_n8145 , new_n8141 , new_n8144 );
  nand g07769 ( new_n8146 , pi069 , pi247 );
  nand g07770 ( new_n8147 , pi029 , pi234 );
  nand g07771 ( new_n8148 , new_n8146 , new_n8147 );
  nand g07772 ( new_n8149 , pi069 , pi234 );
  nor  g07773 ( new_n8150 , new_n8081 , new_n8149 );
  not  g07774 ( new_n8151 , new_n8150 );
  nand g07775 ( new_n8152 , new_n8148 , new_n8151 );
  xor  g07776 ( new_n8153 , new_n8145 , new_n8152 );
  nand g07777 ( new_n8154 , pi016 , pi150 );
  nand g07778 ( new_n8155 , pi117 , pi221 );
  nand g07779 ( new_n8156 , new_n8154 , new_n8155 );
  nand g07780 ( new_n8157 , pi016 , pi221 );
  or   g07781 ( new_n8158 , new_n8084 , new_n8157 );
  nand g07782 ( new_n8159 , new_n8156 , new_n8158 );
  xor  g07783 ( new_n8160 , new_n8153 , new_n8159 );
  nand g07784 ( new_n8161 , new_n8084 , new_n8087 );
  nand g07785 ( new_n8162 , new_n8083 , new_n8088 );
  nand g07786 ( new_n8163 , new_n8161 , new_n8162 );
  xor  g07787 ( new_n8164 , new_n8160 , new_n8163 );
  not  g07788 ( new_n8165 , new_n8090 );
  nor  g07789 ( new_n8166 , new_n8165 , new_n8094 );
  nor  g07790 ( new_n8167 , new_n8089 , new_n8095 );
  nor  g07791 ( new_n8168 , new_n8166 , new_n8167 );
  not  g07792 ( new_n8169 , new_n8168 );
  nor  g07793 ( new_n8170 , new_n8164 , new_n8169 );
  nand g07794 ( new_n8171 , pi244 , pi247 );
  nand g07795 ( new_n8172 , pi029 , pi214 );
  xor  g07796 ( new_n8173 , new_n8149 , new_n8172 );
  xor  g07797 ( new_n8174 , new_n8171 , new_n8173 );
  nand g07798 ( new_n8175 , pi080 , pi150 );
  xor  g07799 ( new_n8176 , new_n8151 , new_n8175 );
  not  g07800 ( new_n8177 , new_n8176 );
  xor  g07801 ( new_n8178 , new_n8174 , new_n8177 );
  nand g07802 ( new_n8179 , pi117 , pi196 );
  nand g07803 ( new_n8180 , pi103 , pi184 );
  xor  g07804 ( new_n8181 , new_n8179 , new_n8180 );
  xor  g07805 ( new_n8182 , new_n8157 , new_n8181 );
  nand g07806 ( new_n8183 , new_n8141 , new_n8144 );
  nand g07807 ( new_n8184 , new_n8145 , new_n8152 );
  nand g07808 ( new_n8185 , new_n8183 , new_n8184 );
  xor  g07809 ( new_n8186 , new_n8182 , new_n8185 );
  xor  g07810 ( new_n8187 , new_n8178 , new_n8186 );
  nand g07811 ( new_n8188 , new_n8153 , new_n8159 );
  nand g07812 ( new_n8189 , new_n8160 , new_n8163 );
  nand g07813 ( new_n8190 , new_n8188 , new_n8189 );
  xor  g07814 ( new_n8191 , new_n8158 , new_n8190 );
  xor  g07815 ( new_n8192 , new_n8187 , new_n8191 );
  nand g07816 ( new_n8193 , new_n8170 , new_n8192 );
  xor  g07817 ( new_n8194 , new_n8170 , new_n8192 );
  nand g07818 ( new_n8195 , pi103 , pi196 );
  xor  g07819 ( new_n8196 , new_n8164 , new_n8168 );
  or   g07820 ( new_n8197 , new_n8195 , new_n8196 );
  not  g07821 ( new_n8198 , new_n8078 );
  nor  g07822 ( new_n8199 , new_n8198 , new_n8096 );
  xor  g07823 ( new_n8200 , new_n8195 , new_n8196 );
  nand g07824 ( new_n8201 , new_n8199 , new_n8200 );
  nand g07825 ( new_n8202 , new_n8197 , new_n8201 );
  nand g07826 ( new_n8203 , new_n8194 , new_n8202 );
  nand g07827 ( new_n8204 , new_n8193 , new_n8203 );
  xor  g07828 ( new_n8205 , new_n8140 , new_n8204 );
  nand g07829 ( new_n8206 , pi010 , pi103 );
  xor  g07830 ( new_n8207 , new_n8205 , new_n8206 );
  or   g07831 ( new_n8208 , new_n8158 , new_n8190 );
  nand g07832 ( new_n8209 , new_n8187 , new_n8191 );
  nand g07833 ( new_n8210 , new_n8208 , new_n8209 );
  nand g07834 ( new_n8211 , pi049 , pi253 );
  nand g07835 ( new_n8212 , pi230 , pi245 );
  or   g07836 ( new_n8213 , new_n7965 , new_n8134 );
  or   g07837 ( new_n8214 , new_n8212 , new_n8213 );
  xor  g07838 ( new_n8215 , new_n8134 , new_n8135 );
  not  g07839 ( new_n8216 , new_n8215 );
  xor  g07840 ( new_n8217 , new_n8212 , new_n8213 );
  nand g07841 ( new_n8218 , new_n8216 , new_n8217 );
  nand g07842 ( new_n8219 , new_n8214 , new_n8218 );
  xor  g07843 ( new_n8220 , new_n8211 , new_n8219 );
  xor  g07844 ( new_n8221 , new_n8210 , new_n8220 );
  xor  g07845 ( new_n8222 , new_n8207 , new_n8221 );
  xor  g07846 ( new_n8223 , new_n8194 , new_n8202 );
  not  g07847 ( new_n8224 , new_n8223 );
  nand g07848 ( new_n8225 , new_n8019 , new_n8037 );
  nand g07849 ( new_n8226 , pi175 , pi195 );
  nand g07850 ( new_n8227 , new_n8225 , new_n8226 );
  nand g07851 ( new_n8228 , pi058 , pi149 );
  nand g07852 ( new_n8229 , new_n8021 , new_n8022 );
  nand g07853 ( new_n8230 , new_n8020 , new_n8023 );
  nand g07854 ( new_n8231 , new_n8229 , new_n8230 );
  xor  g07855 ( new_n8232 , new_n8228 , new_n8231 );
  nand g07856 ( new_n8233 , pi167 , pi186 );
  nand g07857 ( new_n8234 , pi132 , pi181 );
  nand g07858 ( new_n8235 , new_n8233 , new_n8234 );
  nand g07859 ( new_n8236 , pi181 , pi186 );
  nor  g07860 ( new_n8237 , new_n8022 , new_n8236 );
  not  g07861 ( new_n8238 , new_n8237 );
  nand g07862 ( new_n8239 , new_n8235 , new_n8238 );
  xor  g07863 ( new_n8240 , new_n8232 , new_n8239 );
  nand g07864 ( new_n8241 , pi211 , pi240 );
  nand g07865 ( new_n8242 , pi134 , pi199 );
  and  g07866 ( new_n8243 , new_n8241 , new_n8242 );
  nand g07867 ( new_n8244 , pi199 , pi240 );
  nor  g07868 ( new_n8245 , new_n8025 , new_n8244 );
  or   g07869 ( new_n8246 , new_n8243 , new_n8245 );
  xnor g07870 ( new_n8247 , new_n8240 , new_n8246 );
  nand g07871 ( new_n8248 , new_n8025 , new_n8028 );
  nand g07872 ( new_n8249 , new_n8024 , new_n8029 );
  nand g07873 ( new_n8250 , new_n8248 , new_n8249 );
  xor  g07874 ( new_n8251 , new_n8247 , new_n8250 );
  not  g07875 ( new_n8252 , new_n8031 );
  nand g07876 ( new_n8253 , new_n8252 , new_n8035 );
  or   g07877 ( new_n8254 , new_n8030 , new_n8036 );
  nand g07878 ( new_n8255 , new_n8253 , new_n8254 );
  xor  g07879 ( new_n8256 , new_n8251 , new_n8255 );
  not  g07880 ( new_n8257 , new_n8256 );
  xor  g07881 ( new_n8258 , new_n8225 , new_n8226 );
  nand g07882 ( new_n8259 , new_n8257 , new_n8258 );
  nand g07883 ( new_n8260 , new_n8227 , new_n8259 );
  nand g07884 ( new_n8261 , new_n8251 , new_n8255 );
  nand g07885 ( new_n8262 , pi132 , pi200 );
  nand g07886 ( new_n8263 , pi058 , pi167 );
  xor  g07887 ( new_n8264 , new_n8262 , new_n8263 );
  xor  g07888 ( new_n8265 , new_n8236 , new_n8264 );
  nand g07889 ( new_n8266 , pi149 , pi211 );
  xor  g07890 ( new_n8267 , new_n8238 , new_n8266 );
  not  g07891 ( new_n8268 , new_n8267 );
  xor  g07892 ( new_n8269 , new_n8265 , new_n8268 );
  nand g07893 ( new_n8270 , pi134 , pi195 );
  nand g07894 ( new_n8271 , pi175 , pi218 );
  xor  g07895 ( new_n8272 , new_n8270 , new_n8271 );
  xor  g07896 ( new_n8273 , new_n8244 , new_n8272 );
  nand g07897 ( new_n8274 , new_n8228 , new_n8231 );
  nand g07898 ( new_n8275 , new_n8232 , new_n8239 );
  nand g07899 ( new_n8276 , new_n8274 , new_n8275 );
  xor  g07900 ( new_n8277 , new_n8273 , new_n8276 );
  xor  g07901 ( new_n8278 , new_n8269 , new_n8277 );
  nor  g07902 ( new_n8279 , new_n8240 , new_n8246 );
  nor  g07903 ( new_n8280 , new_n8247 , new_n8250 );
  xor  g07904 ( new_n8281 , new_n8245 , new_n8280 );
  nor  g07905 ( new_n8282 , new_n8279 , new_n8281 );
  xor  g07906 ( new_n8283 , new_n8278 , new_n8282 );
  xor  g07907 ( new_n8284 , new_n8261 , new_n8283 );
  xor  g07908 ( new_n8285 , new_n8260 , new_n8284 );
  nand g07909 ( new_n8286 , pi173 , pi245 );
  nand g07910 ( new_n8287 , pi014 , pi201 );
  nand g07911 ( new_n8288 , pi109 , pi156 );
  nand g07912 ( new_n8289 , new_n8287 , new_n8288 );
  nand g07913 ( new_n8290 , new_n8213 , new_n8289 );
  xor  g07914 ( new_n8291 , new_n8286 , new_n8290 );
  nand g07915 ( new_n8292 , new_n7964 , new_n7965 );
  nand g07916 ( new_n8293 , new_n7963 , new_n7966 );
  nand g07917 ( new_n8294 , new_n8292 , new_n8293 );
  xor  g07918 ( new_n8295 , new_n8291 , new_n8294 );
  nand g07919 ( new_n8296 , pi049 , pi230 );
  nand g07920 ( new_n8297 , pi050 , pi171 );
  and  g07921 ( new_n8298 , new_n8296 , new_n8297 );
  nor  g07922 ( new_n8299 , new_n7968 , new_n8126 );
  or   g07923 ( new_n8300 , new_n8298 , new_n8299 );
  xnor g07924 ( new_n8301 , new_n8295 , new_n8300 );
  nand g07925 ( new_n8302 , new_n7968 , new_n7971 );
  nand g07926 ( new_n8303 , new_n7967 , new_n7972 );
  nand g07927 ( new_n8304 , new_n8302 , new_n8303 );
  xor  g07928 ( new_n8305 , new_n8301 , new_n8304 );
  or   g07929 ( new_n8306 , new_n7974 , new_n7977 );
  nand g07930 ( new_n8307 , new_n7973 , new_n7978 );
  nand g07931 ( new_n8308 , new_n8306 , new_n8307 );
  nand g07932 ( new_n8309 , new_n8305 , new_n8308 );
  xor  g07933 ( new_n8310 , new_n8215 , new_n8217 );
  xor  g07934 ( new_n8311 , new_n8126 , new_n8127 );
  nand g07935 ( new_n8312 , new_n8286 , new_n8290 );
  nand g07936 ( new_n8313 , new_n8291 , new_n8294 );
  nand g07937 ( new_n8314 , new_n8312 , new_n8313 );
  xor  g07938 ( new_n8315 , new_n8311 , new_n8314 );
  xnor g07939 ( new_n8316 , new_n8310 , new_n8315 );
  nor  g07940 ( new_n8317 , new_n8295 , new_n8300 );
  nor  g07941 ( new_n8318 , new_n8301 , new_n8304 );
  xor  g07942 ( new_n8319 , new_n8299 , new_n8318 );
  nor  g07943 ( new_n8320 , new_n8317 , new_n8319 );
  xor  g07944 ( new_n8321 , new_n8316 , new_n8320 );
  xnor g07945 ( new_n8322 , new_n8309 , new_n8321 );
  nand g07946 ( new_n8323 , new_n7962 , new_n7979 );
  nand g07947 ( new_n8324 , pi107 , pi253 );
  nand g07948 ( new_n8325 , new_n8323 , new_n8324 );
  xnor g07949 ( new_n8326 , new_n8305 , new_n8308 );
  xor  g07950 ( new_n8327 , new_n8323 , new_n8324 );
  nand g07951 ( new_n8328 , new_n8326 , new_n8327 );
  nand g07952 ( new_n8329 , new_n8325 , new_n8328 );
  xnor g07953 ( new_n8330 , new_n8322 , new_n8329 );
  nor  g07954 ( new_n8331 , new_n7927 , new_n7944 );
  not  g07955 ( new_n8332 , new_n8331 );
  nand g07956 ( new_n8333 , pi025 , pi163 );
  nand g07957 ( new_n8334 , new_n8332 , new_n8333 );
  nand g07958 ( new_n8335 , pi039 , pi066 );
  nand g07959 ( new_n8336 , pi116 , pi207 );
  nand g07960 ( new_n8337 , pi070 , pi226 );
  nand g07961 ( new_n8338 , new_n8336 , new_n8337 );
  nand g07962 ( new_n8339 , pi070 , pi207 );
  or   g07963 ( new_n8340 , new_n7933 , new_n8339 );
  nand g07964 ( new_n8341 , new_n8338 , new_n8340 );
  xor  g07965 ( new_n8342 , new_n8335 , new_n8341 );
  nand g07966 ( new_n8343 , new_n7934 , new_n7935 );
  nand g07967 ( new_n8344 , new_n7933 , new_n7936 );
  nand g07968 ( new_n8345 , new_n8343 , new_n8344 );
  xor  g07969 ( new_n8346 , new_n8342 , new_n8345 );
  nand g07970 ( new_n8347 , new_n7938 , new_n7941 );
  nand g07971 ( new_n8348 , new_n7937 , new_n7942 );
  nand g07972 ( new_n8349 , new_n8347 , new_n8348 );
  nand g07973 ( new_n8350 , pi055 , pi228 );
  nand g07974 ( new_n8351 , pi002 , pi148 );
  nand g07975 ( new_n8352 , new_n8350 , new_n8351 );
  nand g07976 ( new_n8353 , pi002 , pi228 );
  or   g07977 ( new_n8354 , new_n7938 , new_n8353 );
  nand g07978 ( new_n8355 , new_n8352 , new_n8354 );
  xor  g07979 ( new_n8356 , new_n8349 , new_n8355 );
  xor  g07980 ( new_n8357 , new_n8346 , new_n8356 );
  or   g07981 ( new_n8358 , new_n7928 , new_n7931 );
  nand g07982 ( new_n8359 , new_n7932 , new_n7943 );
  nand g07983 ( new_n8360 , new_n8358 , new_n8359 );
  xor  g07984 ( new_n8361 , new_n8357 , new_n8360 );
  xor  g07985 ( new_n8362 , new_n8332 , new_n8333 );
  nand g07986 ( new_n8363 , new_n8361 , new_n8362 );
  nand g07987 ( new_n8364 , new_n8334 , new_n8363 );
  not  g07988 ( new_n8365 , new_n8357 );
  nand g07989 ( new_n8366 , new_n8365 , new_n8360 );
  nand g07990 ( new_n8367 , pi115 , pi226 );
  nand g07991 ( new_n8368 , pi066 , pi116 );
  xor  g07992 ( new_n8369 , new_n8367 , new_n8368 );
  xor  g07993 ( new_n8370 , new_n8339 , new_n8369 );
  not  g07994 ( new_n8371 , new_n8370 );
  nand g07995 ( new_n8372 , pi039 , pi055 );
  xor  g07996 ( new_n8373 , new_n8340 , new_n8372 );
  xor  g07997 ( new_n8374 , new_n8371 , new_n8373 );
  nand g07998 ( new_n8375 , pi163 , pi239 );
  nand g07999 ( new_n8376 , pi025 , pi148 );
  xor  g08000 ( new_n8377 , new_n8375 , new_n8376 );
  xor  g08001 ( new_n8378 , new_n8353 , new_n8377 );
  nand g08002 ( new_n8379 , new_n8335 , new_n8341 );
  nand g08003 ( new_n8380 , new_n8342 , new_n8345 );
  nand g08004 ( new_n8381 , new_n8379 , new_n8380 );
  xor  g08005 ( new_n8382 , new_n8378 , new_n8381 );
  xor  g08006 ( new_n8383 , new_n8374 , new_n8382 );
  nand g08007 ( new_n8384 , new_n8349 , new_n8355 );
  nand g08008 ( new_n8385 , new_n8346 , new_n8356 );
  nand g08009 ( new_n8386 , new_n8384 , new_n8385 );
  xor  g08010 ( new_n8387 , new_n8354 , new_n8386 );
  xnor g08011 ( new_n8388 , new_n8383 , new_n8387 );
  xor  g08012 ( new_n8389 , new_n8366 , new_n8388 );
  xor  g08013 ( new_n8390 , new_n8364 , new_n8389 );
  xor  g08014 ( new_n8391 , new_n8330 , new_n8390 );
  xnor g08015 ( new_n8392 , new_n8361 , new_n8362 );
  nand g08016 ( new_n8393 , new_n7945 , new_n7980 );
  nand g08017 ( new_n8394 , new_n7981 , new_n8000 );
  nand g08018 ( new_n8395 , new_n8393 , new_n8394 );
  nand g08019 ( new_n8396 , new_n8392 , new_n8395 );
  xnor g08020 ( new_n8397 , new_n8326 , new_n8327 );
  xor  g08021 ( new_n8398 , new_n8392 , new_n8395 );
  nand g08022 ( new_n8399 , new_n8397 , new_n8398 );
  nand g08023 ( new_n8400 , new_n8396 , new_n8399 );
  xor  g08024 ( new_n8401 , new_n8391 , new_n8400 );
  xor  g08025 ( new_n8402 , new_n8256 , new_n8258 );
  nand g08026 ( new_n8403 , new_n8001 , new_n8038 );
  nand g08027 ( new_n8404 , new_n8039 , new_n8055 );
  nand g08028 ( new_n8405 , new_n8403 , new_n8404 );
  nand g08029 ( new_n8406 , new_n8402 , new_n8405 );
  xor  g08030 ( new_n8407 , new_n8397 , new_n8398 );
  xor  g08031 ( new_n8408 , new_n8402 , new_n8405 );
  nand g08032 ( new_n8409 , new_n8407 , new_n8408 );
  nand g08033 ( new_n8410 , new_n8406 , new_n8409 );
  xor  g08034 ( new_n8411 , new_n8401 , new_n8410 );
  xor  g08035 ( new_n8412 , new_n8285 , new_n8411 );
  nor  g08036 ( new_n8413 , new_n8224 , new_n8412 );
  xor  g08037 ( new_n8414 , new_n8223 , new_n8412 );
  xnor g08038 ( new_n8415 , new_n8199 , new_n8200 );
  nand g08039 ( new_n8416 , new_n8097 , new_n8114 );
  not  g08040 ( new_n8417 , new_n8056 );
  nand g08041 ( new_n8418 , new_n8417 , new_n8115 );
  nand g08042 ( new_n8419 , new_n8416 , new_n8418 );
  nand g08043 ( new_n8420 , new_n8415 , new_n8419 );
  xor  g08044 ( new_n8421 , new_n8407 , new_n8408 );
  not  g08045 ( new_n8422 , new_n8421 );
  xor  g08046 ( new_n8423 , new_n8415 , new_n8419 );
  nand g08047 ( new_n8424 , new_n8422 , new_n8423 );
  nand g08048 ( new_n8425 , new_n8420 , new_n8424 );
  nor  g08049 ( new_n8426 , new_n8414 , new_n8425 );
  nor  g08050 ( new_n8427 , new_n8413 , new_n8426 );
  nand g08051 ( new_n8428 , new_n8311 , new_n8314 );
  nand g08052 ( new_n8429 , new_n8310 , new_n8315 );
  nand g08053 ( new_n8430 , new_n8428 , new_n8429 );
  xor  g08054 ( new_n8431 , new_n8427 , new_n8430 );
  xor  g08055 ( new_n8432 , new_n8222 , new_n8431 );
  xor  g08056 ( new_n8433 , new_n8139 , new_n8432 );
  xor  g08057 ( new_n8434 , new_n8122 , new_n8433 );
  nand g08058 ( new_n8435 , pi014 , pi063 );
  nand g08059 ( new_n8436 , pi156 , pi173 );
  xor  g08060 ( new_n8437 , new_n8435 , new_n8436 );
  nand g08061 ( new_n8438 , new_n8378 , new_n8381 );
  not  g08062 ( new_n8439 , new_n8374 );
  nand g08063 ( new_n8440 , new_n8439 , new_n8382 );
  nand g08064 ( new_n8441 , new_n8438 , new_n8440 );
  nand g08065 ( new_n8442 , pi055 , pi116 );
  xor  g08066 ( new_n8443 , new_n8441 , new_n8442 );
  nand g08067 ( new_n8444 , new_n8367 , new_n8368 );
  nand g08068 ( new_n8445 , new_n8339 , new_n8369 );
  nand g08069 ( new_n8446 , new_n8444 , new_n8445 );
  nand g08070 ( new_n8447 , new_n8375 , new_n8376 );
  nand g08071 ( new_n8448 , new_n8353 , new_n8377 );
  nand g08072 ( new_n8449 , new_n8447 , new_n8448 );
  nand g08073 ( new_n8450 , pi002 , pi039 );
  xor  g08074 ( new_n8451 , new_n8449 , new_n8450 );
  xor  g08075 ( new_n8452 , new_n8446 , new_n8451 );
  or   g08076 ( new_n8453 , new_n8340 , new_n8372 );
  nand g08077 ( new_n8454 , new_n8371 , new_n8373 );
  nand g08078 ( new_n8455 , new_n8453 , new_n8454 );
  nand g08079 ( new_n8456 , pi148 , pi239 );
  nand g08080 ( new_n8457 , pi025 , pi228 );
  xnor g08081 ( new_n8458 , new_n8456 , new_n8457 );
  xor  g08082 ( new_n8459 , new_n8455 , new_n8458 );
  xor  g08083 ( new_n8460 , new_n8452 , new_n8459 );
  xor  g08084 ( new_n8461 , new_n8443 , new_n8460 );
  xor  g08085 ( new_n8462 , new_n8437 , new_n8461 );
  nor  g08086 ( new_n8463 , new_n8309 , new_n8321 );
  nor  g08087 ( new_n8464 , new_n8322 , new_n8329 );
  nor  g08088 ( new_n8465 , new_n8463 , new_n8464 );
  nand g08089 ( new_n8466 , pi083 , pi109 );
  xor  g08090 ( new_n8467 , new_n8465 , new_n8466 );
  xor  g08091 ( new_n8468 , new_n8462 , new_n8467 );
  nand g08092 ( new_n8469 , new_n8299 , new_n8318 );
  not  g08093 ( new_n8470 , new_n8320 );
  nand g08094 ( new_n8471 , new_n8316 , new_n8470 );
  nand g08095 ( new_n8472 , new_n8469 , new_n8471 );
  nand g08096 ( new_n8473 , pi201 , pi230 );
  nand g08097 ( new_n8474 , pi050 , pi245 );
  xor  g08098 ( new_n8475 , new_n8473 , new_n8474 );
  xor  g08099 ( new_n8476 , new_n8472 , new_n8475 );
  xor  g08100 ( new_n8477 , new_n8468 , new_n8476 );
  xor  g08101 ( new_n8478 , new_n8434 , new_n8477 );
  nand g08102 ( new_n8479 , pi186 , pi200 );
  nand g08103 ( new_n8480 , pi132 , pi203 );
  nand g08104 ( new_n8481 , new_n8245 , new_n8280 );
  not  g08105 ( new_n8482 , new_n8282 );
  nand g08106 ( new_n8483 , new_n8278 , new_n8482 );
  nand g08107 ( new_n8484 , new_n8481 , new_n8483 );
  xor  g08108 ( new_n8485 , new_n8480 , new_n8484 );
  nand g08109 ( new_n8486 , pi037 , pi175 );
  nand g08110 ( new_n8487 , new_n8261 , new_n8283 );
  nand g08111 ( new_n8488 , new_n8260 , new_n8284 );
  nand g08112 ( new_n8489 , new_n8487 , new_n8488 );
  xor  g08113 ( new_n8490 , new_n8486 , new_n8489 );
  xor  g08114 ( new_n8491 , new_n8485 , new_n8490 );
  xor  g08115 ( new_n8492 , new_n8479 , new_n8491 );
  nand g08116 ( new_n8493 , new_n8149 , new_n8172 );
  nand g08117 ( new_n8494 , new_n8171 , new_n8173 );
  nand g08118 ( new_n8495 , new_n8493 , new_n8494 );
  nor  g08119 ( new_n8496 , new_n8151 , new_n8175 );
  nor  g08120 ( new_n8497 , new_n8174 , new_n8177 );
  or   g08121 ( new_n8498 , new_n8496 , new_n8497 );
  xor  g08122 ( new_n8499 , new_n8495 , new_n8498 );
  xor  g08123 ( new_n8500 , new_n8492 , new_n8499 );
  xor  g08124 ( new_n8501 , new_n8478 , new_n8500 );
  or   g08125 ( new_n8502 , new_n8354 , new_n8386 );
  nand g08126 ( new_n8503 , new_n8383 , new_n8387 );
  nand g08127 ( new_n8504 , new_n8502 , new_n8503 );
  nand g08128 ( new_n8505 , new_n8366 , new_n8388 );
  nand g08129 ( new_n8506 , new_n8364 , new_n8389 );
  nand g08130 ( new_n8507 , new_n8505 , new_n8506 );
  xor  g08131 ( new_n8508 , new_n8504 , new_n8507 );
  nand g08132 ( new_n8509 , pi149 , pi199 );
  nand g08133 ( new_n8510 , pi195 , pi240 );
  xor  g08134 ( new_n8511 , new_n8509 , new_n8510 );
  nand g08135 ( new_n8512 , pi167 , pi211 );
  nand g08136 ( new_n8513 , new_n8273 , new_n8276 );
  not  g08137 ( new_n8514 , new_n8269 );
  nand g08138 ( new_n8515 , new_n8514 , new_n8277 );
  nand g08139 ( new_n8516 , new_n8513 , new_n8515 );
  xnor g08140 ( new_n8517 , new_n8512 , new_n8516 );
  xor  g08141 ( new_n8518 , new_n8511 , new_n8517 );
  xor  g08142 ( new_n8519 , new_n8508 , new_n8518 );
  nand g08143 ( new_n8520 , new_n8262 , new_n8263 );
  nand g08144 ( new_n8521 , new_n8236 , new_n8264 );
  nand g08145 ( new_n8522 , new_n8520 , new_n8521 );
  nand g08146 ( new_n8523 , pi134 , pi218 );
  nand g08147 ( new_n8524 , new_n8270 , new_n8271 );
  nand g08148 ( new_n8525 , new_n8244 , new_n8272 );
  nand g08149 ( new_n8526 , new_n8524 , new_n8525 );
  xor  g08150 ( new_n8527 , new_n8523 , new_n8526 );
  xor  g08151 ( new_n8528 , new_n8522 , new_n8527 );
  nor  g08152 ( new_n8529 , new_n8238 , new_n8266 );
  nor  g08153 ( new_n8530 , new_n8265 , new_n8268 );
  or   g08154 ( new_n8531 , new_n8529 , new_n8530 );
  nand g08155 ( new_n8532 , pi058 , pi181 );
  xor  g08156 ( new_n8533 , new_n8531 , new_n8532 );
  xor  g08157 ( new_n8534 , new_n8528 , new_n8533 );
  xor  g08158 ( new_n8535 , new_n8519 , new_n8534 );
  nand g08159 ( new_n8536 , pi069 , pi214 );
  nand g08160 ( new_n8537 , pi150 , pi247 );
  xor  g08161 ( new_n8538 , new_n8536 , new_n8537 );
  xor  g08162 ( new_n8539 , new_n8535 , new_n8538 );
  or   g08163 ( new_n8540 , new_n8401 , new_n8410 );
  nand g08164 ( new_n8541 , new_n8285 , new_n8411 );
  nand g08165 ( new_n8542 , new_n8540 , new_n8541 );
  nand g08166 ( new_n8543 , new_n8182 , new_n8185 );
  not  g08167 ( new_n8544 , new_n8178 );
  nand g08168 ( new_n8545 , new_n8544 , new_n8186 );
  nand g08169 ( new_n8546 , new_n8543 , new_n8545 );
  nand g08170 ( new_n8547 , new_n8179 , new_n8180 );
  nand g08171 ( new_n8548 , new_n8157 , new_n8181 );
  nand g08172 ( new_n8549 , new_n8547 , new_n8548 );
  xor  g08173 ( new_n8550 , new_n8546 , new_n8549 );
  nand g08174 ( new_n8551 , pi080 , pi221 );
  xor  g08175 ( new_n8552 , new_n8550 , new_n8551 );
  xor  g08176 ( new_n8553 , new_n8542 , new_n8552 );
  xor  g08177 ( new_n8554 , new_n8539 , new_n8553 );
  nand g08178 ( new_n8555 , pi000 , pi226 );
  nand g08179 ( new_n8556 , pi115 , pi207 );
  nand g08180 ( new_n8557 , pi066 , pi070 );
  xor  g08181 ( new_n8558 , new_n8556 , new_n8557 );
  nand g08182 ( new_n8559 , pi163 , pi243 );
  nand g08183 ( new_n8560 , new_n8330 , new_n8390 );
  not  g08184 ( new_n8561 , new_n8391 );
  or   g08185 ( new_n8562 , new_n8561 , new_n8400 );
  nand g08186 ( new_n8563 , new_n8560 , new_n8562 );
  xor  g08187 ( new_n8564 , new_n8559 , new_n8563 );
  xor  g08188 ( new_n8565 , new_n8558 , new_n8564 );
  xor  g08189 ( new_n8566 , new_n8555 , new_n8565 );
  nand g08190 ( new_n8567 , pi234 , pi244 );
  nand g08191 ( new_n8568 , pi117 , pi184 );
  nand g08192 ( new_n8569 , pi016 , pi196 );
  xor  g08193 ( new_n8570 , new_n8568 , new_n8569 );
  xor  g08194 ( new_n8571 , new_n8567 , new_n8570 );
  xor  g08195 ( new_n8572 , new_n8566 , new_n8571 );
  xor  g08196 ( new_n8573 , new_n8554 , new_n8572 );
  xor  g08197 ( po047 , new_n8501 , new_n8573 );
  xnor g08198 ( po048 , new_n4794 , new_n4808 );
  xor  g08199 ( po049 , new_n3094 , new_n3095 );
  nor  g08200 ( new_n8577 , new_n1097 , new_n1104 );
  nand g08201 ( new_n8578 , pi161 , pi252 );
  nand g08202 ( new_n8579 , pi090 , pi242 );
  nand g08203 ( new_n8580 , pi140 , pi141 );
  xor  g08204 ( new_n8581 , new_n8579 , new_n8580 );
  xor  g08205 ( new_n8582 , new_n8578 , new_n8581 );
  nand g08206 ( new_n8583 , pi121 , pi241 );
  nand g08207 ( new_n8584 , new_n1093 , new_n1094 );
  nand g08208 ( new_n8585 , new_n1092 , new_n1095 );
  nand g08209 ( new_n8586 , new_n8584 , new_n8585 );
  xor  g08210 ( new_n8587 , new_n8583 , new_n8586 );
  xor  g08211 ( new_n8588 , new_n8582 , new_n8587 );
  nand g08212 ( new_n8589 , pi231 , pi236 );
  or   g08213 ( new_n8590 , new_n1089 , new_n1090 );
  nand g08214 ( new_n8591 , new_n1091 , new_n1096 );
  nand g08215 ( new_n8592 , new_n8590 , new_n8591 );
  xor  g08216 ( new_n8593 , new_n8589 , new_n8592 );
  xor  g08217 ( new_n8594 , new_n8588 , new_n8593 );
  xor  g08218 ( new_n8595 , new_n8577 , new_n8594 );
  nor  g08219 ( new_n8596 , new_n1120 , new_n1127 );
  nand g08220 ( new_n8597 , pi024 , pi104 );
  nand g08221 ( new_n8598 , pi112 , pi210 );
  nand g08222 ( new_n8599 , pi013 , pi111 );
  xor  g08223 ( new_n8600 , new_n8598 , new_n8599 );
  xor  g08224 ( new_n8601 , new_n8597 , new_n8600 );
  nand g08225 ( new_n8602 , pi212 , pi224 );
  nand g08226 ( new_n8603 , new_n1107 , new_n1108 );
  nand g08227 ( new_n8604 , new_n1106 , new_n1109 );
  nand g08228 ( new_n8605 , new_n8603 , new_n8604 );
  xor  g08229 ( new_n8606 , new_n8602 , new_n8605 );
  xnor g08230 ( new_n8607 , new_n8601 , new_n8606 );
  nand g08231 ( new_n8608 , pi213 , pi255 );
  nand g08232 ( new_n8609 , new_n1117 , new_n1118 );
  nand g08233 ( new_n8610 , new_n1110 , new_n1119 );
  nand g08234 ( new_n8611 , new_n8609 , new_n8610 );
  xor  g08235 ( new_n8612 , new_n8608 , new_n8611 );
  xor  g08236 ( new_n8613 , new_n8607 , new_n8612 );
  xnor g08237 ( new_n8614 , new_n8596 , new_n8613 );
  not  g08238 ( new_n8615 , new_n1128 );
  nor  g08239 ( new_n8616 , new_n1105 , new_n8615 );
  nor  g08240 ( new_n8617 , new_n1129 , new_n1150 );
  nor  g08241 ( new_n8618 , new_n8616 , new_n8617 );
  xor  g08242 ( new_n8619 , new_n8614 , new_n8618 );
  xor  g08243 ( new_n8620 , new_n8595 , new_n8619 );
  or   g08244 ( new_n8621 , new_n1070 , new_n1081 );
  nand g08245 ( new_n8622 , pi015 , pi249 );
  nand g08246 ( new_n8623 , pi035 , pi222 );
  nand g08247 ( new_n8624 , pi125 , pi139 );
  xor  g08248 ( new_n8625 , new_n8623 , new_n8624 );
  xor  g08249 ( new_n8626 , new_n8622 , new_n8625 );
  nand g08250 ( new_n8627 , pi176 , pi208 );
  nand g08251 ( new_n8628 , new_n1072 , new_n1073 );
  nand g08252 ( new_n8629 , new_n1071 , new_n1074 );
  nand g08253 ( new_n8630 , new_n8628 , new_n8629 );
  xor  g08254 ( new_n8631 , new_n8627 , new_n8630 );
  xnor g08255 ( new_n8632 , new_n8626 , new_n8631 );
  nand g08256 ( new_n8633 , pi040 , pi168 );
  nand g08257 ( new_n8634 , new_n1076 , new_n1079 );
  nand g08258 ( new_n8635 , new_n1075 , new_n1080 );
  nand g08259 ( new_n8636 , new_n8634 , new_n8635 );
  xor  g08260 ( new_n8637 , new_n8633 , new_n8636 );
  xnor g08261 ( new_n8638 , new_n8632 , new_n8637 );
  xor  g08262 ( new_n8639 , new_n8621 , new_n8638 );
  nand g08263 ( new_n8640 , new_n1082 , new_n1151 );
  nand g08264 ( new_n8641 , new_n1152 , new_n1171 );
  nand g08265 ( new_n8642 , new_n8640 , new_n8641 );
  xor  g08266 ( new_n8643 , new_n8639 , new_n8642 );
  xnor g08267 ( new_n8644 , new_n8620 , new_n8643 );
  nor  g08268 ( new_n8645 , new_n1187 , new_n1194 );
  nand g08269 ( new_n8646 , pi106 , pi131 );
  nand g08270 ( new_n8647 , new_n1184 , new_n1185 );
  nand g08271 ( new_n8648 , new_n1177 , new_n1186 );
  nand g08272 ( new_n8649 , new_n8647 , new_n8648 );
  xor  g08273 ( new_n8650 , new_n8646 , new_n8649 );
  nand g08274 ( new_n8651 , pi100 , pi133 );
  nand g08275 ( new_n8652 , pi077 , pi227 );
  nand g08276 ( new_n8653 , pi189 , pi217 );
  xor  g08277 ( new_n8654 , new_n8652 , new_n8653 );
  xor  g08278 ( new_n8655 , new_n8651 , new_n8654 );
  nand g08279 ( new_n8656 , pi052 , pi081 );
  nand g08280 ( new_n8657 , new_n1174 , new_n1175 );
  nand g08281 ( new_n8658 , new_n1173 , new_n1176 );
  nand g08282 ( new_n8659 , new_n8657 , new_n8658 );
  xor  g08283 ( new_n8660 , new_n8656 , new_n8659 );
  xnor g08284 ( new_n8661 , new_n8655 , new_n8660 );
  xor  g08285 ( new_n8662 , new_n8650 , new_n8661 );
  xor  g08286 ( new_n8663 , new_n8645 , new_n8662 );
  not  g08287 ( new_n8664 , new_n8663 );
  xor  g08288 ( new_n8665 , new_n8644 , new_n8664 );
  nand g08289 ( new_n8666 , new_n1195 , new_n1213 );
  not  g08290 ( new_n8667 , new_n1172 );
  nand g08291 ( new_n8668 , new_n8667 , new_n1214 );
  nand g08292 ( new_n8669 , new_n8666 , new_n8668 );
  xnor g08293 ( po050 , new_n8665 , new_n8669 );
  nand g08294 ( new_n8671 , pi125 , pi216 );
  nand g08295 ( new_n8672 , pi076 , pi222 );
  nand g08296 ( new_n8673 , pi079 , pi249 );
  nand g08297 ( new_n8674 , new_n8672 , new_n8673 );
  nand g08298 ( new_n8675 , pi076 , pi249 );
  nand g08299 ( new_n8676 , pi079 , pi222 );
  or   g08300 ( new_n8677 , new_n8675 , new_n8676 );
  nand g08301 ( new_n8678 , new_n8674 , new_n8677 );
  xor  g08302 ( new_n8679 , new_n8671 , new_n8678 );
  nand g08303 ( new_n8680 , pi041 , pi125 );
  nand g08304 ( new_n8681 , new_n8675 , new_n8680 );
  nand g08305 ( new_n8682 , pi216 , pi222 );
  xor  g08306 ( new_n8683 , new_n8675 , new_n8680 );
  nand g08307 ( new_n8684 , new_n8682 , new_n8683 );
  nand g08308 ( new_n8685 , new_n8681 , new_n8684 );
  xor  g08309 ( new_n8686 , new_n8679 , new_n8685 );
  nand g08310 ( new_n8687 , pi176 , pi182 );
  nand g08311 ( new_n8688 , pi041 , pi222 );
  nand g08312 ( new_n8689 , pi216 , pi249 );
  nand g08313 ( new_n8690 , new_n8688 , new_n8689 );
  nand g08314 ( new_n8691 , pi125 , pi182 );
  xor  g08315 ( new_n8692 , new_n8688 , new_n8689 );
  nand g08316 ( new_n8693 , new_n8691 , new_n8692 );
  nand g08317 ( new_n8694 , new_n8690 , new_n8693 );
  nand g08318 ( new_n8695 , new_n8687 , new_n8694 );
  xor  g08319 ( new_n8696 , new_n8682 , new_n8683 );
  xor  g08320 ( new_n8697 , new_n8687 , new_n8694 );
  nand g08321 ( new_n8698 , new_n8696 , new_n8697 );
  nand g08322 ( new_n8699 , new_n8695 , new_n8698 );
  nand g08323 ( new_n8700 , pi041 , pi176 );
  nand g08324 ( new_n8701 , pi040 , pi182 );
  nand g08325 ( new_n8702 , new_n8700 , new_n8701 );
  nand g08326 ( new_n8703 , pi040 , pi041 );
  or   g08327 ( new_n8704 , new_n8687 , new_n8703 );
  nand g08328 ( new_n8705 , new_n8702 , new_n8704 );
  xor  g08329 ( new_n8706 , new_n8699 , new_n8705 );
  xor  g08330 ( new_n8707 , new_n8686 , new_n8706 );
  not  g08331 ( new_n8708 , new_n8707 );
  xor  g08332 ( new_n8709 , new_n8696 , new_n8697 );
  nand g08333 ( new_n8710 , pi040 , pi138 );
  or   g08334 ( new_n8711 , new_n8709 , new_n8710 );
  xor  g08335 ( new_n8712 , new_n8709 , new_n8710 );
  nand g08336 ( new_n8713 , pi041 , pi249 );
  nand g08337 ( new_n8714 , pi125 , pi138 );
  nand g08338 ( new_n8715 , new_n8713 , new_n8714 );
  nand g08339 ( new_n8716 , pi182 , pi222 );
  or   g08340 ( new_n8717 , new_n8713 , new_n8714 );
  nand g08341 ( new_n8718 , new_n8716 , new_n8717 );
  nand g08342 ( new_n8719 , new_n8715 , new_n8718 );
  nand g08343 ( new_n8720 , pi138 , pi176 );
  or   g08344 ( new_n8721 , new_n8719 , new_n8720 );
  xnor g08345 ( new_n8722 , new_n8691 , new_n8692 );
  xor  g08346 ( new_n8723 , new_n8719 , new_n8720 );
  nand g08347 ( new_n8724 , new_n8722 , new_n8723 );
  nand g08348 ( new_n8725 , new_n8721 , new_n8724 );
  nand g08349 ( new_n8726 , new_n8712 , new_n8725 );
  nand g08350 ( new_n8727 , new_n8711 , new_n8726 );
  nand g08351 ( new_n8728 , new_n8708 , new_n8727 );
  nand g08352 ( new_n8729 , pi076 , pi125 );
  nand g08353 ( new_n8730 , pi249 , pi251 );
  xor  g08354 ( new_n8731 , new_n8729 , new_n8730 );
  xor  g08355 ( new_n8732 , new_n8676 , new_n8731 );
  not  g08356 ( new_n8733 , new_n8732 );
  nand g08357 ( new_n8734 , pi176 , pi216 );
  xor  g08358 ( new_n8735 , new_n8677 , new_n8734 );
  xor  g08359 ( new_n8736 , new_n8733 , new_n8735 );
  nand g08360 ( new_n8737 , pi174 , pi182 );
  nand g08361 ( new_n8738 , pi138 , pi157 );
  xor  g08362 ( new_n8739 , new_n8737 , new_n8738 );
  xor  g08363 ( new_n8740 , new_n8703 , new_n8739 );
  nand g08364 ( new_n8741 , new_n8671 , new_n8678 );
  nand g08365 ( new_n8742 , new_n8679 , new_n8685 );
  nand g08366 ( new_n8743 , new_n8741 , new_n8742 );
  xor  g08367 ( new_n8744 , new_n8740 , new_n8743 );
  xor  g08368 ( new_n8745 , new_n8736 , new_n8744 );
  nand g08369 ( new_n8746 , new_n8699 , new_n8705 );
  nand g08370 ( new_n8747 , new_n8686 , new_n8706 );
  nand g08371 ( new_n8748 , new_n8746 , new_n8747 );
  xor  g08372 ( new_n8749 , new_n8704 , new_n8748 );
  xnor g08373 ( new_n8750 , new_n8745 , new_n8749 );
  xnor g08374 ( new_n8751 , new_n8728 , new_n8750 );
  nand g08375 ( new_n8752 , pi138 , pi174 );
  xor  g08376 ( new_n8753 , new_n8712 , new_n8725 );
  xnor g08377 ( new_n8754 , new_n8722 , new_n8723 );
  not  g08378 ( new_n8755 , new_n8716 );
  not  g08379 ( new_n8756 , new_n8715 );
  nand g08380 ( new_n8757 , pi138 , pi249 );
  nand g08381 ( new_n8758 , new_n8755 , new_n8757 );
  nand g08382 ( new_n8759 , new_n8756 , new_n8758 );
  nand g08383 ( new_n8760 , new_n8717 , new_n8759 );
  nand g08384 ( new_n8761 , new_n8755 , new_n8760 );
  nor  g08385 ( new_n8762 , new_n8754 , new_n8761 );
  nand g08386 ( new_n8763 , new_n8753 , new_n8762 );
  nand g08387 ( new_n8764 , new_n8752 , new_n8763 );
  xor  g08388 ( new_n8765 , new_n8707 , new_n8727 );
  xor  g08389 ( new_n8766 , new_n8752 , new_n8763 );
  nand g08390 ( new_n8767 , new_n8765 , new_n8766 );
  nand g08391 ( new_n8768 , new_n8764 , new_n8767 );
  xor  g08392 ( new_n8769 , new_n8751 , new_n8768 );
  nand g08393 ( new_n8770 , pi024 , pi123 );
  nand g08394 ( new_n8771 , pi023 , pi210 );
  nand g08395 ( new_n8772 , pi099 , pi111 );
  nand g08396 ( new_n8773 , new_n8771 , new_n8772 );
  nand g08397 ( new_n8774 , pi099 , pi210 );
  nand g08398 ( new_n8775 , pi023 , pi111 );
  or   g08399 ( new_n8776 , new_n8774 , new_n8775 );
  nand g08400 ( new_n8777 , new_n8773 , new_n8776 );
  xor  g08401 ( new_n8778 , new_n8770 , new_n8777 );
  nand g08402 ( new_n8779 , pi024 , pi169 );
  nand g08403 ( new_n8780 , pi111 , pi123 );
  nand g08404 ( new_n8781 , new_n8779 , new_n8780 );
  xor  g08405 ( new_n8782 , new_n8779 , new_n8780 );
  nand g08406 ( new_n8783 , new_n8774 , new_n8782 );
  nand g08407 ( new_n8784 , new_n8781 , new_n8783 );
  xor  g08408 ( new_n8785 , new_n8778 , new_n8784 );
  nand g08409 ( new_n8786 , pi169 , pi224 );
  nand g08410 ( new_n8787 , pi071 , pi255 );
  and  g08411 ( new_n8788 , new_n8786 , new_n8787 );
  nand g08412 ( new_n8789 , pi071 , pi224 );
  nand g08413 ( new_n8790 , pi169 , pi255 );
  nor  g08414 ( new_n8791 , new_n8789 , new_n8790 );
  or   g08415 ( new_n8792 , new_n8788 , new_n8791 );
  xnor g08416 ( new_n8793 , new_n8785 , new_n8792 );
  nand g08417 ( new_n8794 , pi111 , pi169 );
  nand g08418 ( new_n8795 , pi024 , pi071 );
  nand g08419 ( new_n8796 , new_n8794 , new_n8795 );
  nand g08420 ( new_n8797 , pi123 , pi210 );
  xor  g08421 ( new_n8798 , new_n8794 , new_n8795 );
  nand g08422 ( new_n8799 , new_n8797 , new_n8798 );
  nand g08423 ( new_n8800 , new_n8796 , new_n8799 );
  nand g08424 ( new_n8801 , new_n8789 , new_n8800 );
  xor  g08425 ( new_n8802 , new_n8774 , new_n8782 );
  xor  g08426 ( new_n8803 , new_n8789 , new_n8800 );
  nand g08427 ( new_n8804 , new_n8802 , new_n8803 );
  nand g08428 ( new_n8805 , new_n8801 , new_n8804 );
  xor  g08429 ( new_n8806 , new_n8793 , new_n8805 );
  nand g08430 ( new_n8807 , pi142 , pi255 );
  not  g08431 ( new_n8808 , new_n8807 );
  nand g08432 ( new_n8809 , pi169 , pi210 );
  nand g08433 ( new_n8810 , pi024 , pi142 );
  nand g08434 ( new_n8811 , new_n8809 , new_n8810 );
  nand g08435 ( new_n8812 , pi071 , pi111 );
  or   g08436 ( new_n8813 , new_n8809 , new_n8810 );
  nand g08437 ( new_n8814 , new_n8812 , new_n8813 );
  nand g08438 ( new_n8815 , new_n8811 , new_n8814 );
  nand g08439 ( new_n8816 , pi142 , pi224 );
  or   g08440 ( new_n8817 , new_n8815 , new_n8816 );
  xor  g08441 ( new_n8818 , new_n8815 , new_n8816 );
  xnor g08442 ( new_n8819 , new_n8797 , new_n8798 );
  nand g08443 ( new_n8820 , new_n8818 , new_n8819 );
  nand g08444 ( new_n8821 , new_n8817 , new_n8820 );
  nand g08445 ( new_n8822 , new_n8808 , new_n8821 );
  xor  g08446 ( new_n8823 , new_n8807 , new_n8821 );
  xor  g08447 ( new_n8824 , new_n8802 , new_n8803 );
  or   g08448 ( new_n8825 , new_n8823 , new_n8824 );
  nand g08449 ( new_n8826 , new_n8822 , new_n8825 );
  nand g08450 ( new_n8827 , new_n8806 , new_n8826 );
  nand g08451 ( new_n8828 , pi024 , pi099 );
  nand g08452 ( new_n8829 , pi155 , pi210 );
  xor  g08453 ( new_n8830 , new_n8775 , new_n8829 );
  xor  g08454 ( new_n8831 , new_n8828 , new_n8830 );
  nand g08455 ( new_n8832 , pi123 , pi224 );
  xor  g08456 ( new_n8833 , new_n8776 , new_n8832 );
  xor  g08457 ( new_n8834 , new_n8831 , new_n8833 );
  nand g08458 ( new_n8835 , pi071 , pi127 );
  nand g08459 ( new_n8836 , pi142 , pi232 );
  xor  g08460 ( new_n8837 , new_n8835 , new_n8836 );
  xor  g08461 ( new_n8838 , new_n8790 , new_n8837 );
  nand g08462 ( new_n8839 , new_n8770 , new_n8777 );
  nand g08463 ( new_n8840 , new_n8778 , new_n8784 );
  nand g08464 ( new_n8841 , new_n8839 , new_n8840 );
  xor  g08465 ( new_n8842 , new_n8838 , new_n8841 );
  xnor g08466 ( new_n8843 , new_n8834 , new_n8842 );
  nor  g08467 ( new_n8844 , new_n8793 , new_n8805 );
  nand g08468 ( new_n8845 , new_n8791 , new_n8844 );
  nor  g08469 ( new_n8846 , new_n8785 , new_n8792 );
  or   g08470 ( new_n8847 , new_n8791 , new_n8846 );
  or   g08471 ( new_n8848 , new_n8844 , new_n8847 );
  nand g08472 ( new_n8849 , new_n8845 , new_n8848 );
  xor  g08473 ( new_n8850 , new_n8843 , new_n8849 );
  xnor g08474 ( new_n8851 , new_n8827 , new_n8850 );
  nand g08475 ( new_n8852 , pi127 , pi142 );
  xnor g08476 ( new_n8853 , new_n8818 , new_n8819 );
  not  g08477 ( new_n8854 , new_n8812 );
  not  g08478 ( new_n8855 , new_n8811 );
  nand g08479 ( new_n8856 , pi142 , pi210 );
  nand g08480 ( new_n8857 , new_n8854 , new_n8856 );
  nand g08481 ( new_n8858 , new_n8855 , new_n8857 );
  nand g08482 ( new_n8859 , new_n8813 , new_n8858 );
  nand g08483 ( new_n8860 , new_n8854 , new_n8859 );
  nor  g08484 ( new_n8861 , new_n8853 , new_n8860 );
  xor  g08485 ( new_n8862 , new_n8823 , new_n8824 );
  nand g08486 ( new_n8863 , new_n8861 , new_n8862 );
  nand g08487 ( new_n8864 , new_n8852 , new_n8863 );
  xnor g08488 ( new_n8865 , new_n8806 , new_n8826 );
  xor  g08489 ( new_n8866 , new_n8852 , new_n8863 );
  nand g08490 ( new_n8867 , new_n8865 , new_n8866 );
  nand g08491 ( new_n8868 , new_n8864 , new_n8867 );
  xor  g08492 ( new_n8869 , new_n8851 , new_n8868 );
  nand g08493 ( new_n8870 , pi135 , pi140 );
  nand g08494 ( new_n8871 , pi122 , pi252 );
  nand g08495 ( new_n8872 , pi059 , pi242 );
  xor  g08496 ( new_n8873 , new_n8871 , new_n8872 );
  xor  g08497 ( new_n8874 , new_n8870 , new_n8873 );
  not  g08498 ( new_n8875 , new_n8874 );
  nand g08499 ( new_n8876 , pi001 , pi121 );
  nand g08500 ( new_n8877 , pi122 , pi242 );
  or   g08501 ( new_n8878 , new_n8870 , new_n8877 );
  xor  g08502 ( new_n8879 , new_n8876 , new_n8878 );
  xor  g08503 ( new_n8880 , new_n8875 , new_n8879 );
  nand g08504 ( new_n8881 , pi102 , pi231 );
  nand g08505 ( new_n8882 , pi021 , pi087 );
  nand g08506 ( new_n8883 , pi005 , pi219 );
  xor  g08507 ( new_n8884 , new_n8882 , new_n8883 );
  xor  g08508 ( new_n8885 , new_n8881 , new_n8884 );
  nand g08509 ( new_n8886 , pi001 , pi252 );
  nand g08510 ( new_n8887 , pi122 , pi140 );
  nand g08511 ( new_n8888 , pi135 , pi242 );
  nand g08512 ( new_n8889 , new_n8887 , new_n8888 );
  nand g08513 ( new_n8890 , new_n8878 , new_n8889 );
  nand g08514 ( new_n8891 , new_n8886 , new_n8890 );
  xor  g08515 ( new_n8892 , new_n8886 , new_n8890 );
  nand g08516 ( new_n8893 , pi001 , pi140 );
  nand g08517 ( new_n8894 , new_n8877 , new_n8893 );
  nand g08518 ( new_n8895 , pi102 , pi252 );
  xor  g08519 ( new_n8896 , new_n8877 , new_n8893 );
  nand g08520 ( new_n8897 , new_n8895 , new_n8896 );
  nand g08521 ( new_n8898 , new_n8894 , new_n8897 );
  nand g08522 ( new_n8899 , new_n8892 , new_n8898 );
  nand g08523 ( new_n8900 , new_n8891 , new_n8899 );
  xor  g08524 ( new_n8901 , new_n8885 , new_n8900 );
  xor  g08525 ( new_n8902 , new_n8880 , new_n8901 );
  not  g08526 ( new_n8903 , new_n8902 );
  nand g08527 ( new_n8904 , pi121 , pi219 );
  or   g08528 ( new_n8905 , new_n8881 , new_n8904 );
  nand g08529 ( new_n8906 , pi001 , pi242 );
  nand g08530 ( new_n8907 , pi219 , pi252 );
  nand g08531 ( new_n8908 , new_n8906 , new_n8907 );
  nand g08532 ( new_n8909 , pi102 , pi140 );
  xor  g08533 ( new_n8910 , new_n8906 , new_n8907 );
  nand g08534 ( new_n8911 , new_n8909 , new_n8910 );
  nand g08535 ( new_n8912 , new_n8908 , new_n8911 );
  nand g08536 ( new_n8913 , new_n8904 , new_n8912 );
  xor  g08537 ( new_n8914 , new_n8895 , new_n8896 );
  xor  g08538 ( new_n8915 , new_n8904 , new_n8912 );
  nand g08539 ( new_n8916 , new_n8914 , new_n8915 );
  nand g08540 ( new_n8917 , new_n8913 , new_n8916 );
  nand g08541 ( new_n8918 , pi102 , pi121 );
  nand g08542 ( new_n8919 , pi219 , pi231 );
  nand g08543 ( new_n8920 , new_n8918 , new_n8919 );
  nand g08544 ( new_n8921 , new_n8905 , new_n8920 );
  nand g08545 ( new_n8922 , new_n8917 , new_n8921 );
  xor  g08546 ( new_n8923 , new_n8892 , new_n8898 );
  xor  g08547 ( new_n8924 , new_n8917 , new_n8921 );
  nand g08548 ( new_n8925 , new_n8923 , new_n8924 );
  nand g08549 ( new_n8926 , new_n8922 , new_n8925 );
  xor  g08550 ( new_n8927 , new_n8905 , new_n8926 );
  xor  g08551 ( new_n8928 , new_n8903 , new_n8927 );
  xor  g08552 ( new_n8929 , new_n8923 , new_n8924 );
  not  g08553 ( new_n8930 , new_n8929 );
  nand g08554 ( new_n8931 , pi087 , pi231 );
  not  g08555 ( new_n8932 , new_n8931 );
  nand g08556 ( new_n8933 , pi102 , pi242 );
  nand g08557 ( new_n8934 , pi087 , pi252 );
  nand g08558 ( new_n8935 , new_n8933 , new_n8934 );
  nand g08559 ( new_n8936 , pi140 , pi219 );
  or   g08560 ( new_n8937 , new_n8933 , new_n8934 );
  nand g08561 ( new_n8938 , new_n8936 , new_n8937 );
  nand g08562 ( new_n8939 , new_n8935 , new_n8938 );
  nand g08563 ( new_n8940 , pi087 , pi121 );
  or   g08564 ( new_n8941 , new_n8939 , new_n8940 );
  xor  g08565 ( new_n8942 , new_n8939 , new_n8940 );
  xnor g08566 ( new_n8943 , new_n8909 , new_n8910 );
  nand g08567 ( new_n8944 , new_n8942 , new_n8943 );
  nand g08568 ( new_n8945 , new_n8941 , new_n8944 );
  nand g08569 ( new_n8946 , new_n8932 , new_n8945 );
  xor  g08570 ( new_n8947 , new_n8914 , new_n8915 );
  xor  g08571 ( new_n8948 , new_n8931 , new_n8945 );
  or   g08572 ( new_n8949 , new_n8947 , new_n8948 );
  nand g08573 ( new_n8950 , new_n8946 , new_n8949 );
  nand g08574 ( new_n8951 , new_n8930 , new_n8950 );
  xnor g08575 ( new_n8952 , new_n8942 , new_n8943 );
  not  g08576 ( new_n8953 , new_n8936 );
  not  g08577 ( new_n8954 , new_n8935 );
  nand g08578 ( new_n8955 , pi087 , pi242 );
  nand g08579 ( new_n8956 , new_n8953 , new_n8955 );
  nand g08580 ( new_n8957 , new_n8954 , new_n8956 );
  nand g08581 ( new_n8958 , new_n8937 , new_n8957 );
  nand g08582 ( new_n8959 , new_n8953 , new_n8958 );
  nor  g08583 ( new_n8960 , new_n8952 , new_n8959 );
  xor  g08584 ( new_n8961 , new_n8947 , new_n8948 );
  nand g08585 ( new_n8962 , new_n8960 , new_n8961 );
  nand g08586 ( new_n8963 , pi005 , pi087 );
  xor  g08587 ( new_n8964 , new_n8929 , new_n8950 );
  xnor g08588 ( new_n8965 , new_n8963 , new_n8964 );
  nor  g08589 ( new_n8966 , new_n8962 , new_n8965 );
  not  g08590 ( new_n8967 , new_n8966 );
  nor  g08591 ( new_n8968 , new_n8951 , new_n8967 );
  or   g08592 ( new_n8969 , new_n8963 , new_n8964 );
  nand g08593 ( new_n8970 , new_n8951 , new_n8969 );
  nor  g08594 ( new_n8971 , new_n8966 , new_n8970 );
  nor  g08595 ( new_n8972 , new_n8968 , new_n8971 );
  xor  g08596 ( new_n8973 , new_n8928 , new_n8972 );
  not  g08597 ( new_n8974 , new_n8973 );
  xor  g08598 ( new_n8975 , new_n8869 , new_n8974 );
  xnor g08599 ( new_n8976 , new_n8865 , new_n8866 );
  xor  g08600 ( new_n8977 , new_n8962 , new_n8965 );
  nand g08601 ( new_n8978 , new_n8976 , new_n8977 );
  xor  g08602 ( new_n8979 , new_n8976 , new_n8977 );
  xor  g08603 ( new_n8980 , new_n8960 , new_n8961 );
  xor  g08604 ( new_n8981 , new_n8861 , new_n8862 );
  nand g08605 ( new_n8982 , new_n8980 , new_n8981 );
  not  g08606 ( new_n8983 , new_n8982 );
  xnor g08607 ( new_n8984 , new_n8980 , new_n8981 );
  xnor g08608 ( new_n8985 , new_n8952 , new_n8959 );
  nor  g08609 ( new_n8986 , new_n8855 , new_n8857 );
  or   g08610 ( new_n8987 , new_n8859 , new_n8986 );
  nor  g08611 ( new_n8988 , new_n8954 , new_n8956 );
  nor  g08612 ( new_n8989 , new_n8958 , new_n8988 );
  not  g08613 ( new_n8990 , new_n8989 );
  nand g08614 ( new_n8991 , new_n8987 , new_n8990 );
  xor  g08615 ( new_n8992 , new_n8987 , new_n8989 );
  nand g08616 ( new_n8993 , pi111 , pi142 );
  nand g08617 ( new_n8994 , pi071 , pi210 );
  xor  g08618 ( new_n8995 , new_n8993 , new_n8994 );
  nor  g08619 ( new_n8996 , new_n8856 , new_n8955 );
  nand g08620 ( new_n8997 , new_n8995 , new_n8996 );
  nand g08621 ( new_n8998 , pi219 , pi242 );
  nand g08622 ( new_n8999 , pi087 , pi140 );
  xor  g08623 ( new_n9000 , new_n8998 , new_n8999 );
  xor  g08624 ( new_n9001 , new_n8995 , new_n8996 );
  nand g08625 ( new_n9002 , new_n9000 , new_n9001 );
  nand g08626 ( new_n9003 , new_n8997 , new_n9002 );
  or   g08627 ( new_n9004 , new_n8992 , new_n9003 );
  nand g08628 ( new_n9005 , new_n8991 , new_n9004 );
  nand g08629 ( new_n9006 , new_n8985 , new_n9005 );
  xor  g08630 ( new_n9007 , new_n8853 , new_n8860 );
  not  g08631 ( new_n9008 , new_n9007 );
  xor  g08632 ( new_n9009 , new_n8985 , new_n9005 );
  nand g08633 ( new_n9010 , new_n9008 , new_n9009 );
  nand g08634 ( new_n9011 , new_n9006 , new_n9010 );
  nor  g08635 ( new_n9012 , new_n8984 , new_n9011 );
  nor  g08636 ( new_n9013 , new_n8983 , new_n9012 );
  not  g08637 ( new_n9014 , new_n9013 );
  nand g08638 ( new_n9015 , new_n8979 , new_n9014 );
  nand g08639 ( new_n9016 , new_n8978 , new_n9015 );
  xor  g08640 ( new_n9017 , new_n8975 , new_n9016 );
  xor  g08641 ( new_n9018 , new_n8769 , new_n9017 );
  xor  g08642 ( new_n9019 , new_n8979 , new_n9013 );
  xor  g08643 ( new_n9020 , new_n8765 , new_n8766 );
  nor  g08644 ( new_n9021 , new_n9019 , new_n9020 );
  xnor g08645 ( new_n9022 , new_n9019 , new_n9020 );
  xor  g08646 ( new_n9023 , new_n8753 , new_n8762 );
  xor  g08647 ( new_n9024 , new_n8754 , new_n8761 );
  xor  g08648 ( new_n9025 , new_n9008 , new_n9009 );
  not  g08649 ( new_n9026 , new_n9025 );
  nor  g08650 ( new_n9027 , new_n9024 , new_n9026 );
  xor  g08651 ( new_n9028 , new_n9024 , new_n9025 );
  xor  g08652 ( new_n9029 , new_n8992 , new_n9003 );
  xor  g08653 ( new_n9030 , new_n8856 , new_n8955 );
  not  g08654 ( new_n9031 , new_n9030 );
  nor  g08655 ( new_n9032 , new_n8757 , new_n9031 );
  nand g08656 ( new_n9033 , pi138 , pi222 );
  nand g08657 ( new_n9034 , pi182 , pi249 );
  xor  g08658 ( new_n9035 , new_n9033 , new_n9034 );
  or   g08659 ( new_n9036 , new_n9032 , new_n9035 );
  xnor g08660 ( new_n9037 , new_n9000 , new_n9001 );
  xor  g08661 ( new_n9038 , new_n9032 , new_n9035 );
  nand g08662 ( new_n9039 , new_n9037 , new_n9038 );
  nand g08663 ( new_n9040 , new_n9036 , new_n9039 );
  or   g08664 ( new_n9041 , new_n9029 , new_n9040 );
  xor  g08665 ( new_n9042 , new_n9029 , new_n9040 );
  nor  g08666 ( new_n9043 , new_n8756 , new_n8758 );
  nor  g08667 ( new_n9044 , new_n8760 , new_n9043 );
  nand g08668 ( new_n9045 , new_n9042 , new_n9044 );
  nand g08669 ( new_n9046 , new_n9041 , new_n9045 );
  nor  g08670 ( new_n9047 , new_n9028 , new_n9046 );
  nor  g08671 ( new_n9048 , new_n9027 , new_n9047 );
  or   g08672 ( new_n9049 , new_n9023 , new_n9048 );
  xor  g08673 ( new_n9050 , new_n8984 , new_n9011 );
  not  g08674 ( new_n9051 , new_n9050 );
  xor  g08675 ( new_n9052 , new_n9023 , new_n9048 );
  nand g08676 ( new_n9053 , new_n9051 , new_n9052 );
  nand g08677 ( new_n9054 , new_n9049 , new_n9053 );
  nor  g08678 ( new_n9055 , new_n9022 , new_n9054 );
  nor  g08679 ( new_n9056 , new_n9021 , new_n9055 );
  xor  g08680 ( new_n9057 , new_n9018 , new_n9056 );
  nand g08681 ( new_n9058 , pi160 , pi233 );
  nand g08682 ( new_n9059 , pi060 , pi217 );
  nand g08683 ( new_n9060 , pi160 , pi227 );
  nand g08684 ( new_n9061 , pi020 , pi100 );
  xor  g08685 ( new_n9062 , new_n9060 , new_n9061 );
  xor  g08686 ( new_n9063 , new_n9059 , new_n9062 );
  nand g08687 ( new_n9064 , pi100 , pi160 );
  nand g08688 ( new_n9065 , pi020 , pi217 );
  nor  g08689 ( new_n9066 , new_n9064 , new_n9065 );
  not  g08690 ( new_n9067 , new_n9066 );
  nor  g08691 ( new_n9068 , new_n9063 , new_n9067 );
  not  g08692 ( new_n9069 , new_n9068 );
  nand g08693 ( new_n9070 , pi020 , pi227 );
  nand g08694 ( new_n9071 , pi217 , pi223 );
  nand g08695 ( new_n9072 , pi060 , pi100 );
  xor  g08696 ( new_n9073 , new_n9071 , new_n9072 );
  xnor g08697 ( new_n9074 , new_n9070 , new_n9073 );
  nand g08698 ( new_n9075 , pi081 , pi160 );
  nand g08699 ( new_n9076 , new_n9060 , new_n9061 );
  nand g08700 ( new_n9077 , new_n9059 , new_n9062 );
  nand g08701 ( new_n9078 , new_n9076 , new_n9077 );
  xor  g08702 ( new_n9079 , new_n9075 , new_n9078 );
  xnor g08703 ( new_n9080 , new_n9074 , new_n9079 );
  nor  g08704 ( new_n9081 , new_n9069 , new_n9080 );
  nand g08705 ( new_n9082 , pi060 , pi227 );
  nand g08706 ( new_n9083 , pi100 , pi223 );
  nand g08707 ( new_n9084 , pi101 , pi217 );
  xor  g08708 ( new_n9085 , new_n9083 , new_n9084 );
  xor  g08709 ( new_n9086 , new_n9082 , new_n9085 );
  nand g08710 ( new_n9087 , pi020 , pi081 );
  nand g08711 ( new_n9088 , new_n9071 , new_n9072 );
  nand g08712 ( new_n9089 , new_n9070 , new_n9073 );
  nand g08713 ( new_n9090 , new_n9088 , new_n9089 );
  xor  g08714 ( new_n9091 , new_n9087 , new_n9090 );
  xor  g08715 ( new_n9092 , new_n9086 , new_n9091 );
  nand g08716 ( new_n9093 , pi106 , pi160 );
  xor  g08717 ( new_n9094 , new_n9092 , new_n9093 );
  or   g08718 ( new_n9095 , new_n9075 , new_n9078 );
  nand g08719 ( new_n9096 , new_n9074 , new_n9079 );
  nand g08720 ( new_n9097 , new_n9095 , new_n9096 );
  xor  g08721 ( new_n9098 , new_n9094 , new_n9097 );
  nand g08722 ( new_n9099 , new_n9081 , new_n9098 );
  nand g08723 ( new_n9100 , new_n9058 , new_n9099 );
  nand g08724 ( new_n9101 , pi223 , pi227 );
  nand g08725 ( new_n9102 , pi217 , pi225 );
  nand g08726 ( new_n9103 , pi100 , pi101 );
  nand g08727 ( new_n9104 , new_n9102 , new_n9103 );
  nand g08728 ( new_n9105 , pi100 , pi225 );
  or   g08729 ( new_n9106 , new_n9084 , new_n9105 );
  nand g08730 ( new_n9107 , new_n9104 , new_n9106 );
  xor  g08731 ( new_n9108 , new_n9101 , new_n9107 );
  nand g08732 ( new_n9109 , new_n9083 , new_n9084 );
  nand g08733 ( new_n9110 , new_n9082 , new_n9085 );
  nand g08734 ( new_n9111 , new_n9109 , new_n9110 );
  xor  g08735 ( new_n9112 , new_n9108 , new_n9111 );
  nand g08736 ( new_n9113 , pi060 , pi081 );
  nand g08737 ( new_n9114 , pi020 , pi106 );
  and  g08738 ( new_n9115 , new_n9113 , new_n9114 );
  nand g08739 ( new_n9116 , pi060 , pi106 );
  nor  g08740 ( new_n9117 , new_n9087 , new_n9116 );
  or   g08741 ( new_n9118 , new_n9115 , new_n9117 );
  xnor g08742 ( new_n9119 , new_n9112 , new_n9118 );
  nand g08743 ( new_n9120 , new_n9087 , new_n9090 );
  nand g08744 ( new_n9121 , new_n9086 , new_n9091 );
  nand g08745 ( new_n9122 , new_n9120 , new_n9121 );
  xor  g08746 ( new_n9123 , new_n9119 , new_n9122 );
  or   g08747 ( new_n9124 , new_n9092 , new_n9093 );
  nand g08748 ( new_n9125 , new_n9094 , new_n9097 );
  nand g08749 ( new_n9126 , new_n9124 , new_n9125 );
  xnor g08750 ( new_n9127 , new_n9123 , new_n9126 );
  xor  g08751 ( new_n9128 , new_n9058 , new_n9099 );
  nand g08752 ( new_n9129 , new_n9127 , new_n9128 );
  nand g08753 ( new_n9130 , new_n9100 , new_n9129 );
  nand g08754 ( new_n9131 , new_n9123 , new_n9126 );
  nand g08755 ( new_n9132 , pi101 , pi227 );
  nand g08756 ( new_n9133 , pi177 , pi217 );
  xor  g08757 ( new_n9134 , new_n9132 , new_n9133 );
  xor  g08758 ( new_n9135 , new_n9105 , new_n9134 );
  nand g08759 ( new_n9136 , pi081 , pi223 );
  xor  g08760 ( new_n9137 , new_n9106 , new_n9136 );
  xor  g08761 ( new_n9138 , new_n9135 , new_n9137 );
  nand g08762 ( new_n9139 , pi020 , pi233 );
  nand g08763 ( new_n9140 , pi160 , pi187 );
  xor  g08764 ( new_n9141 , new_n9139 , new_n9140 );
  xor  g08765 ( new_n9142 , new_n9116 , new_n9141 );
  nand g08766 ( new_n9143 , new_n9101 , new_n9107 );
  nand g08767 ( new_n9144 , new_n9108 , new_n9111 );
  nand g08768 ( new_n9145 , new_n9143 , new_n9144 );
  xor  g08769 ( new_n9146 , new_n9142 , new_n9145 );
  xnor g08770 ( new_n9147 , new_n9138 , new_n9146 );
  nor  g08771 ( new_n9148 , new_n9112 , new_n9118 );
  nor  g08772 ( new_n9149 , new_n9119 , new_n9122 );
  xor  g08773 ( new_n9150 , new_n9117 , new_n9149 );
  nor  g08774 ( new_n9151 , new_n9148 , new_n9150 );
  xor  g08775 ( new_n9152 , new_n9147 , new_n9151 );
  xor  g08776 ( new_n9153 , new_n9131 , new_n9152 );
  xor  g08777 ( new_n9154 , new_n9130 , new_n9153 );
  or   g08778 ( new_n9155 , new_n9057 , new_n9154 );
  xor  g08779 ( new_n9156 , new_n9022 , new_n9054 );
  not  g08780 ( new_n9157 , new_n9156 );
  xor  g08781 ( new_n9158 , new_n9127 , new_n9128 );
  or   g08782 ( new_n9159 , new_n9157 , new_n9158 );
  xor  g08783 ( new_n9160 , new_n9157 , new_n9158 );
  xnor g08784 ( new_n9161 , new_n9081 , new_n9098 );
  xor  g08785 ( new_n9162 , new_n9028 , new_n9046 );
  xor  g08786 ( new_n9163 , new_n9063 , new_n9066 );
  nand g08787 ( new_n9164 , pi160 , pi217 );
  xor  g08788 ( new_n9165 , new_n8757 , new_n9030 );
  nor  g08789 ( new_n9166 , new_n9164 , new_n9165 );
  xor  g08790 ( new_n9167 , new_n9064 , new_n9065 );
  or   g08791 ( new_n9168 , new_n9166 , new_n9167 );
  xor  g08792 ( new_n9169 , new_n9037 , new_n9038 );
  xor  g08793 ( new_n9170 , new_n9166 , new_n9167 );
  nand g08794 ( new_n9171 , new_n9169 , new_n9170 );
  nand g08795 ( new_n9172 , new_n9168 , new_n9171 );
  nand g08796 ( new_n9173 , new_n9163 , new_n9172 );
  xor  g08797 ( new_n9174 , new_n9042 , new_n9044 );
  not  g08798 ( new_n9175 , new_n9174 );
  xor  g08799 ( new_n9176 , new_n9163 , new_n9172 );
  nand g08800 ( new_n9177 , new_n9175 , new_n9176 );
  nand g08801 ( new_n9178 , new_n9173 , new_n9177 );
  nand g08802 ( new_n9179 , new_n9162 , new_n9178 );
  xor  g08803 ( new_n9180 , new_n9069 , new_n9080 );
  not  g08804 ( new_n9181 , new_n9180 );
  xor  g08805 ( new_n9182 , new_n9162 , new_n9178 );
  nand g08806 ( new_n9183 , new_n9181 , new_n9182 );
  nand g08807 ( new_n9184 , new_n9179 , new_n9183 );
  or   g08808 ( new_n9185 , new_n9161 , new_n9184 );
  xor  g08809 ( new_n9186 , new_n9050 , new_n9052 );
  xor  g08810 ( new_n9187 , new_n9161 , new_n9184 );
  nand g08811 ( new_n9188 , new_n9186 , new_n9187 );
  nand g08812 ( new_n9189 , new_n9185 , new_n9188 );
  nand g08813 ( new_n9190 , new_n9160 , new_n9189 );
  nand g08814 ( new_n9191 , new_n9159 , new_n9190 );
  xor  g08815 ( new_n9192 , new_n9057 , new_n9154 );
  nand g08816 ( new_n9193 , new_n9191 , new_n9192 );
  nand g08817 ( new_n9194 , new_n9155 , new_n9193 );
  nand g08818 ( new_n9195 , new_n9131 , new_n9152 );
  nand g08819 ( new_n9196 , new_n9130 , new_n9153 );
  nand g08820 ( new_n9197 , new_n9195 , new_n9196 );
  xor  g08821 ( new_n9198 , new_n9194 , new_n9197 );
  nand g08822 ( new_n9199 , pi111 , pi155 );
  nand g08823 ( new_n9200 , pi023 , pi024 );
  xor  g08824 ( new_n9201 , new_n9199 , new_n9200 );
  nand g08825 ( new_n9202 , pi076 , pi176 );
  or   g08826 ( new_n9203 , new_n8677 , new_n8734 );
  nand g08827 ( new_n9204 , new_n8733 , new_n8735 );
  nand g08828 ( new_n9205 , new_n9203 , new_n9204 );
  xor  g08829 ( new_n9206 , new_n9202 , new_n9205 );
  nand g08830 ( new_n9207 , pi040 , pi216 );
  nand g08831 ( new_n9208 , pi041 , pi174 );
  xor  g08832 ( new_n9209 , new_n9207 , new_n9208 );
  nand g08833 ( new_n9210 , pi079 , pi125 );
  xor  g08834 ( new_n9211 , new_n9209 , new_n9210 );
  nand g08835 ( new_n9212 , pi157 , pi182 );
  nand g08836 ( new_n9213 , new_n8729 , new_n8730 );
  nand g08837 ( new_n9214 , new_n8676 , new_n8731 );
  nand g08838 ( new_n9215 , new_n9213 , new_n9214 );
  nand g08839 ( new_n9216 , new_n8740 , new_n8743 );
  not  g08840 ( new_n9217 , new_n8736 );
  nand g08841 ( new_n9218 , new_n9217 , new_n8744 );
  nand g08842 ( new_n9219 , new_n9216 , new_n9218 );
  xor  g08843 ( new_n9220 , new_n9215 , new_n9219 );
  xor  g08844 ( new_n9221 , new_n9212 , new_n9220 );
  xor  g08845 ( new_n9222 , new_n9211 , new_n9221 );
  xor  g08846 ( new_n9223 , new_n9206 , new_n9222 );
  xor  g08847 ( new_n9224 , new_n9201 , new_n9223 );
  xor  g08848 ( new_n9225 , new_n9198 , new_n9224 );
  nand g08849 ( new_n9226 , pi142 , pi191 );
  nand g08850 ( new_n9227 , new_n8737 , new_n8738 );
  nand g08851 ( new_n9228 , new_n8703 , new_n8739 );
  nand g08852 ( new_n9229 , new_n9227 , new_n9228 );
  xor  g08853 ( new_n9230 , new_n9226 , new_n9229 );
  nand g08854 ( new_n9231 , pi017 , pi138 );
  nand g08855 ( new_n9232 , new_n9142 , new_n9145 );
  nand g08856 ( new_n9233 , new_n9138 , new_n9146 );
  nand g08857 ( new_n9234 , new_n9232 , new_n9233 );
  xor  g08858 ( new_n9235 , new_n9231 , new_n9234 );
  nand g08859 ( new_n9236 , new_n9139 , new_n9140 );
  nand g08860 ( new_n9237 , new_n9116 , new_n9141 );
  nand g08861 ( new_n9238 , new_n9236 , new_n9237 );
  nand g08862 ( new_n9239 , pi192 , pi249 );
  or   g08863 ( new_n9240 , new_n8704 , new_n8748 );
  nand g08864 ( new_n9241 , new_n8745 , new_n8749 );
  nand g08865 ( new_n9242 , new_n9240 , new_n9241 );
  xor  g08866 ( new_n9243 , new_n9239 , new_n9242 );
  nand g08867 ( new_n9244 , pi222 , pi251 );
  xor  g08868 ( new_n9245 , new_n9243 , new_n9244 );
  xor  g08869 ( new_n9246 , new_n9238 , new_n9245 );
  xor  g08870 ( new_n9247 , new_n9235 , new_n9246 );
  nand g08871 ( new_n9248 , new_n9132 , new_n9133 );
  nand g08872 ( new_n9249 , new_n9105 , new_n9134 );
  nand g08873 ( new_n9250 , new_n9248 , new_n9249 );
  or   g08874 ( new_n9251 , new_n9106 , new_n9136 );
  not  g08875 ( new_n9252 , new_n9135 );
  nand g08876 ( new_n9253 , new_n9252 , new_n9137 );
  nand g08877 ( new_n9254 , new_n9251 , new_n9253 );
  xor  g08878 ( new_n9255 , new_n9250 , new_n9254 );
  xor  g08879 ( new_n9256 , new_n9247 , new_n9255 );
  xor  g08880 ( new_n9257 , new_n9230 , new_n9256 );
  or   g08881 ( new_n9258 , new_n8769 , new_n9017 );
  nand g08882 ( new_n9259 , new_n9018 , new_n9056 );
  nand g08883 ( new_n9260 , new_n9258 , new_n9259 );
  nand g08884 ( new_n9261 , pi121 , pi122 );
  nand g08885 ( new_n9262 , pi001 , pi231 );
  xor  g08886 ( new_n9263 , new_n9261 , new_n9262 );
  nand g08887 ( new_n9264 , new_n8838 , new_n8841 );
  nand g08888 ( new_n9265 , new_n8834 , new_n8842 );
  nand g08889 ( new_n9266 , new_n9264 , new_n9265 );
  nand g08890 ( new_n9267 , pi099 , pi224 );
  xor  g08891 ( new_n9268 , new_n9266 , new_n9267 );
  nand g08892 ( new_n9269 , new_n8775 , new_n8829 );
  nand g08893 ( new_n9270 , new_n8828 , new_n8830 );
  nand g08894 ( new_n9271 , new_n9269 , new_n9270 );
  nand g08895 ( new_n9272 , new_n8835 , new_n8836 );
  nand g08896 ( new_n9273 , new_n8790 , new_n8837 );
  nand g08897 ( new_n9274 , new_n9272 , new_n9273 );
  nand g08898 ( new_n9275 , pi123 , pi255 );
  xor  g08899 ( new_n9276 , new_n9274 , new_n9275 );
  xor  g08900 ( new_n9277 , new_n9271 , new_n9276 );
  or   g08901 ( new_n9278 , new_n8776 , new_n8832 );
  not  g08902 ( new_n9279 , new_n8831 );
  nand g08903 ( new_n9280 , new_n9279 , new_n8833 );
  nand g08904 ( new_n9281 , new_n9278 , new_n9280 );
  nand g08905 ( new_n9282 , pi071 , pi232 );
  nand g08906 ( new_n9283 , pi127 , pi169 );
  xor  g08907 ( new_n9284 , new_n9282 , new_n9283 );
  xor  g08908 ( new_n9285 , new_n9281 , new_n9284 );
  xor  g08909 ( new_n9286 , new_n9277 , new_n9285 );
  xor  g08910 ( new_n9287 , new_n9268 , new_n9286 );
  xor  g08911 ( new_n9288 , new_n9263 , new_n9287 );
  xor  g08912 ( new_n9289 , new_n9260 , new_n9288 );
  nand g08913 ( new_n9290 , new_n8905 , new_n8926 );
  nand g08914 ( new_n9291 , new_n8903 , new_n8927 );
  nand g08915 ( new_n9292 , new_n9290 , new_n9291 );
  nand g08916 ( new_n9293 , pi082 , pi087 );
  xor  g08917 ( new_n9294 , new_n9292 , new_n9293 );
  and  g08918 ( new_n9295 , new_n8928 , new_n8972 );
  or   g08919 ( new_n9296 , new_n8971 , new_n9295 );
  nand g08920 ( new_n9297 , pi059 , pi140 );
  nand g08921 ( new_n9298 , pi094 , pi242 );
  xor  g08922 ( new_n9299 , new_n9297 , new_n9298 );
  xor  g08923 ( new_n9300 , new_n9296 , new_n9299 );
  xor  g08924 ( new_n9301 , new_n9294 , new_n9300 );
  nand g08925 ( new_n9302 , pi135 , pi252 );
  nand g08926 ( new_n9303 , pi137 , pi217 );
  nand g08927 ( new_n9304 , pi129 , pi160 );
  xor  g08928 ( new_n9305 , new_n9303 , new_n9304 );
  or   g08929 ( new_n9306 , new_n8885 , new_n8900 );
  nand g08930 ( new_n9307 , new_n8880 , new_n8901 );
  nand g08931 ( new_n9308 , new_n9306 , new_n9307 );
  nand g08932 ( new_n9309 , pi021 , pi219 );
  nand g08933 ( new_n9310 , pi005 , pi102 );
  xor  g08934 ( new_n9311 , new_n9309 , new_n9310 );
  xor  g08935 ( new_n9312 , new_n9308 , new_n9311 );
  xor  g08936 ( new_n9313 , new_n9305 , new_n9312 );
  nand g08937 ( new_n9314 , new_n9117 , new_n9149 );
  not  g08938 ( new_n9315 , new_n9151 );
  nand g08939 ( new_n9316 , new_n9147 , new_n9315 );
  nand g08940 ( new_n9317 , new_n9314 , new_n9316 );
  nand g08941 ( new_n9318 , new_n8871 , new_n8872 );
  nand g08942 ( new_n9319 , new_n8870 , new_n8873 );
  nand g08943 ( new_n9320 , new_n9318 , new_n9319 );
  nand g08944 ( new_n9321 , new_n8882 , new_n8883 );
  nand g08945 ( new_n9322 , new_n8881 , new_n8884 );
  nand g08946 ( new_n9323 , new_n9321 , new_n9322 );
  xnor g08947 ( new_n9324 , new_n9320 , new_n9323 );
  or   g08948 ( new_n9325 , new_n8876 , new_n8878 );
  nand g08949 ( new_n9326 , new_n8875 , new_n8879 );
  nand g08950 ( new_n9327 , new_n9325 , new_n9326 );
  xor  g08951 ( new_n9328 , new_n9324 , new_n9327 );
  xor  g08952 ( new_n9329 , new_n9317 , new_n9328 );
  xor  g08953 ( new_n9330 , new_n9313 , new_n9329 );
  xor  g08954 ( new_n9331 , new_n9302 , new_n9330 );
  xor  g08955 ( new_n9332 , new_n9301 , new_n9331 );
  xor  g08956 ( new_n9333 , new_n9289 , new_n9332 );
  nand g08957 ( new_n9334 , pi100 , pi177 );
  nor  g08958 ( new_n9335 , new_n8728 , new_n8750 );
  nor  g08959 ( new_n9336 , new_n8751 , new_n8768 );
  or   g08960 ( new_n9337 , new_n9335 , new_n9336 );
  nand g08961 ( new_n9338 , pi081 , pi101 );
  nand g08962 ( new_n9339 , pi106 , pi223 );
  xor  g08963 ( new_n9340 , new_n9338 , new_n9339 );
  xor  g08964 ( new_n9341 , new_n9337 , new_n9340 );
  xor  g08965 ( new_n9342 , new_n9334 , new_n9341 );
  nand g08966 ( new_n9343 , pi225 , pi227 );
  nand g08967 ( new_n9344 , pi020 , pi187 );
  nand g08968 ( new_n9345 , pi060 , pi233 );
  xor  g08969 ( new_n9346 , new_n9344 , new_n9345 );
  xor  g08970 ( new_n9347 , new_n9343 , new_n9346 );
  xor  g08971 ( new_n9348 , new_n9342 , new_n9347 );
  xor  g08972 ( new_n9349 , new_n9333 , new_n9348 );
  xor  g08973 ( new_n9350 , new_n9257 , new_n9349 );
  nand g08974 ( new_n9351 , pi086 , pi210 );
  or   g08975 ( new_n9352 , new_n8843 , new_n8849 );
  nand g08976 ( new_n9353 , new_n8848 , new_n9352 );
  nor  g08977 ( new_n9354 , new_n8827 , new_n8850 );
  nor  g08978 ( new_n9355 , new_n8851 , new_n8868 );
  nor  g08979 ( new_n9356 , new_n9354 , new_n9355 );
  nand g08980 ( new_n9357 , new_n8869 , new_n8974 );
  nand g08981 ( new_n9358 , new_n8975 , new_n9016 );
  nand g08982 ( new_n9359 , new_n9357 , new_n9358 );
  xor  g08983 ( new_n9360 , new_n9356 , new_n9359 );
  xor  g08984 ( new_n9361 , new_n9353 , new_n9360 );
  xor  g08985 ( new_n9362 , new_n9351 , new_n9361 );
  xor  g08986 ( new_n9363 , new_n9350 , new_n9362 );
  xor  g08987 ( po051 , new_n9225 , new_n9363 );
  xor  g08988 ( po052 , new_n3234 , new_n3251 );
  xor  g08989 ( po053 , new_n3452 , new_n3492 );
  xor  g08990 ( po054 , new_n846 , new_n872 );
  xor  g08991 ( po055 , new_n7516 , new_n7530 );
  xor  g08992 ( po056 , new_n3937 , new_n3938 );
  xor  g08993 ( po057 , new_n1807 , new_n1809 );
  xor  g08994 ( po058 , new_n3749 , new_n3750 );
  xor  g08995 ( po059 , new_n5354 , new_n5356 );
  xor  g08996 ( po060 , new_n2547 , new_n2571 );
  xor  g08997 ( po061 , new_n2566 , new_n2567 );
  nand g08998 ( new_n9375 , new_n8656 , new_n8659 );
  nand g08999 ( new_n9376 , new_n8655 , new_n8660 );
  nand g09000 ( new_n9377 , new_n9375 , new_n9376 );
  nand g09001 ( new_n9378 , pi133 , pi227 );
  nand g09002 ( new_n9379 , new_n8652 , new_n8653 );
  nand g09003 ( new_n9380 , new_n8651 , new_n8654 );
  nand g09004 ( new_n9381 , new_n9379 , new_n9380 );
  nand g09005 ( new_n9382 , pi100 , pi189 );
  nand g09006 ( new_n9383 , pi064 , pi217 );
  nand g09007 ( new_n9384 , new_n9382 , new_n9383 );
  nand g09008 ( new_n9385 , pi064 , pi100 );
  or   g09009 ( new_n9386 , new_n8653 , new_n9385 );
  nand g09010 ( new_n9387 , new_n9384 , new_n9386 );
  xor  g09011 ( new_n9388 , new_n9381 , new_n9387 );
  xor  g09012 ( new_n9389 , new_n9378 , new_n9388 );
  nand g09013 ( new_n9390 , pi077 , pi081 );
  nand g09014 ( new_n9391 , pi052 , pi106 );
  nand g09015 ( new_n9392 , new_n9390 , new_n9391 );
  nand g09016 ( new_n9393 , pi077 , pi106 );
  or   g09017 ( new_n9394 , new_n8656 , new_n9393 );
  nand g09018 ( new_n9395 , new_n9392 , new_n9394 );
  xor  g09019 ( new_n9396 , new_n9389 , new_n9395 );
  xor  g09020 ( new_n9397 , new_n9377 , new_n9396 );
  not  g09021 ( new_n9398 , new_n9397 );
  or   g09022 ( new_n9399 , new_n8646 , new_n8649 );
  nand g09023 ( new_n9400 , new_n8650 , new_n8661 );
  nand g09024 ( new_n9401 , new_n9399 , new_n9400 );
  nand g09025 ( new_n9402 , new_n9398 , new_n9401 );
  nand g09026 ( new_n9403 , new_n9389 , new_n9395 );
  nand g09027 ( new_n9404 , new_n9377 , new_n9396 );
  nand g09028 ( new_n9405 , new_n9403 , new_n9404 );
  xor  g09029 ( new_n9406 , new_n9394 , new_n9405 );
  nand g09030 ( new_n9407 , pi189 , pi227 );
  nand g09031 ( new_n9408 , pi084 , pi217 );
  xor  g09032 ( new_n9409 , new_n9407 , new_n9408 );
  xor  g09033 ( new_n9410 , new_n9385 , new_n9409 );
  nand g09034 ( new_n9411 , pi081 , pi133 );
  xor  g09035 ( new_n9412 , new_n9386 , new_n9411 );
  xor  g09036 ( new_n9413 , new_n9410 , new_n9412 );
  nand g09037 ( new_n9414 , pi131 , pi187 );
  nand g09038 ( new_n9415 , pi052 , pi233 );
  xor  g09039 ( new_n9416 , new_n9414 , new_n9415 );
  xor  g09040 ( new_n9417 , new_n9393 , new_n9416 );
  nand g09041 ( new_n9418 , new_n9381 , new_n9387 );
  nand g09042 ( new_n9419 , new_n9378 , new_n9388 );
  nand g09043 ( new_n9420 , new_n9418 , new_n9419 );
  xor  g09044 ( new_n9421 , new_n9417 , new_n9420 );
  xor  g09045 ( new_n9422 , new_n9413 , new_n9421 );
  xor  g09046 ( new_n9423 , new_n9406 , new_n9422 );
  nand g09047 ( new_n9424 , new_n8645 , new_n8662 );
  nand g09048 ( new_n9425 , pi131 , pi233 );
  nand g09049 ( new_n9426 , new_n9424 , new_n9425 );
  xor  g09050 ( new_n9427 , new_n9397 , new_n9401 );
  xor  g09051 ( new_n9428 , new_n9424 , new_n9425 );
  nand g09052 ( new_n9429 , new_n9427 , new_n9428 );
  nand g09053 ( new_n9430 , new_n9426 , new_n9429 );
  xnor g09054 ( new_n9431 , new_n9423 , new_n9430 );
  xor  g09055 ( new_n9432 , new_n9402 , new_n9431 );
  nand g09056 ( new_n9433 , pi035 , pi125 );
  nand g09057 ( new_n9434 , new_n8623 , new_n8624 );
  nand g09058 ( new_n9435 , new_n8622 , new_n8625 );
  nand g09059 ( new_n9436 , new_n9434 , new_n9435 );
  nand g09060 ( new_n9437 , pi204 , pi249 );
  nand g09061 ( new_n9438 , pi015 , pi222 );
  nand g09062 ( new_n9439 , new_n9437 , new_n9438 );
  nand g09063 ( new_n9440 , pi204 , pi222 );
  or   g09064 ( new_n9441 , new_n8622 , new_n9440 );
  nand g09065 ( new_n9442 , new_n9439 , new_n9441 );
  xor  g09066 ( new_n9443 , new_n9436 , new_n9442 );
  xor  g09067 ( new_n9444 , new_n9433 , new_n9443 );
  nand g09068 ( new_n9445 , new_n8627 , new_n8630 );
  nand g09069 ( new_n9446 , new_n8626 , new_n8631 );
  nand g09070 ( new_n9447 , new_n9445 , new_n9446 );
  nand g09071 ( new_n9448 , new_n9444 , new_n9447 );
  or   g09072 ( new_n9449 , new_n9444 , new_n9447 );
  and  g09073 ( new_n9450 , new_n9448 , new_n9449 );
  nand g09074 ( new_n9451 , pi139 , pi176 );
  nand g09075 ( new_n9452 , pi040 , pi208 );
  nand g09076 ( new_n9453 , new_n9451 , new_n9452 );
  nand g09077 ( new_n9454 , pi040 , pi139 );
  or   g09078 ( new_n9455 , new_n8627 , new_n9454 );
  nand g09079 ( new_n9456 , new_n9453 , new_n9455 );
  xor  g09080 ( new_n9457 , new_n9450 , new_n9456 );
  not  g09081 ( new_n9458 , new_n9457 );
  or   g09082 ( new_n9459 , new_n8633 , new_n8636 );
  nand g09083 ( new_n9460 , new_n8632 , new_n8637 );
  nand g09084 ( new_n9461 , new_n9459 , new_n9460 );
  nand g09085 ( new_n9462 , new_n9458 , new_n9461 );
  nand g09086 ( new_n9463 , pi146 , pi249 );
  nand g09087 ( new_n9464 , pi015 , pi125 );
  xor  g09088 ( new_n9465 , new_n9463 , new_n9464 );
  xor  g09089 ( new_n9466 , new_n9440 , new_n9465 );
  nand g09090 ( new_n9467 , pi035 , pi176 );
  xor  g09091 ( new_n9468 , new_n9441 , new_n9467 );
  xor  g09092 ( new_n9469 , new_n9466 , new_n9468 );
  nand g09093 ( new_n9470 , pi174 , pi208 );
  nand g09094 ( new_n9471 , pi157 , pi168 );
  xor  g09095 ( new_n9472 , new_n9470 , new_n9471 );
  xor  g09096 ( new_n9473 , new_n9454 , new_n9472 );
  nand g09097 ( new_n9474 , new_n9436 , new_n9442 );
  nand g09098 ( new_n9475 , new_n9433 , new_n9443 );
  nand g09099 ( new_n9476 , new_n9474 , new_n9475 );
  xor  g09100 ( new_n9477 , new_n9473 , new_n9476 );
  xor  g09101 ( new_n9478 , new_n9469 , new_n9477 );
  nand g09102 ( new_n9479 , new_n9450 , new_n9456 );
  nand g09103 ( new_n9480 , new_n9448 , new_n9479 );
  and  g09104 ( new_n9481 , new_n9455 , new_n9480 );
  nor  g09105 ( new_n9482 , new_n9449 , new_n9455 );
  or   g09106 ( new_n9483 , new_n9481 , new_n9482 );
  xnor g09107 ( new_n9484 , new_n9478 , new_n9483 );
  xor  g09108 ( new_n9485 , new_n9462 , new_n9484 );
  nand g09109 ( new_n9486 , pi168 , pi174 );
  xor  g09110 ( new_n9487 , new_n9457 , new_n9461 );
  or   g09111 ( new_n9488 , new_n9486 , new_n9487 );
  nor  g09112 ( new_n9489 , new_n8621 , new_n8638 );
  xor  g09113 ( new_n9490 , new_n9486 , new_n9487 );
  nand g09114 ( new_n9491 , new_n9489 , new_n9490 );
  nand g09115 ( new_n9492 , new_n9488 , new_n9491 );
  xnor g09116 ( new_n9493 , new_n9485 , new_n9492 );
  xor  g09117 ( new_n9494 , new_n9489 , new_n9490 );
  nand g09118 ( new_n9495 , new_n8639 , new_n8642 );
  nand g09119 ( new_n9496 , new_n8620 , new_n8643 );
  nand g09120 ( new_n9497 , new_n9495 , new_n9496 );
  or   g09121 ( new_n9498 , new_n9494 , new_n9497 );
  xor  g09122 ( new_n9499 , new_n9494 , new_n9497 );
  nand g09123 ( new_n9500 , new_n8577 , new_n8594 );
  nand g09124 ( new_n9501 , pi141 , pi252 );
  nand g09125 ( new_n9502 , pi090 , pi140 );
  nand g09126 ( new_n9503 , pi047 , pi242 );
  nand g09127 ( new_n9504 , new_n9502 , new_n9503 );
  nand g09128 ( new_n9505 , pi047 , pi140 );
  or   g09129 ( new_n9506 , new_n8579 , new_n9505 );
  nand g09130 ( new_n9507 , new_n9504 , new_n9506 );
  xor  g09131 ( new_n9508 , new_n9501 , new_n9507 );
  nand g09132 ( new_n9509 , new_n8579 , new_n8580 );
  nand g09133 ( new_n9510 , new_n8578 , new_n8581 );
  nand g09134 ( new_n9511 , new_n9509 , new_n9510 );
  xor  g09135 ( new_n9512 , new_n9508 , new_n9511 );
  nand g09136 ( new_n9513 , pi121 , pi161 );
  nand g09137 ( new_n9514 , pi231 , pi241 );
  and  g09138 ( new_n9515 , new_n9513 , new_n9514 );
  nand g09139 ( new_n9516 , pi161 , pi231 );
  nor  g09140 ( new_n9517 , new_n8583 , new_n9516 );
  or   g09141 ( new_n9518 , new_n9515 , new_n9517 );
  xnor g09142 ( new_n9519 , new_n9512 , new_n9518 );
  nand g09143 ( new_n9520 , new_n8583 , new_n8586 );
  nand g09144 ( new_n9521 , new_n8582 , new_n8587 );
  nand g09145 ( new_n9522 , new_n9520 , new_n9521 );
  xor  g09146 ( new_n9523 , new_n9519 , new_n9522 );
  not  g09147 ( new_n9524 , new_n8589 );
  nand g09148 ( new_n9525 , new_n9524 , new_n8592 );
  or   g09149 ( new_n9526 , new_n8588 , new_n8593 );
  nand g09150 ( new_n9527 , new_n9525 , new_n9526 );
  xnor g09151 ( new_n9528 , new_n9523 , new_n9527 );
  nand g09152 ( new_n9529 , pi005 , pi236 );
  xor  g09153 ( new_n9530 , new_n9528 , new_n9529 );
  xor  g09154 ( new_n9531 , new_n9500 , new_n9530 );
  nand g09155 ( new_n9532 , new_n8602 , new_n8605 );
  nand g09156 ( new_n9533 , new_n8601 , new_n8606 );
  nand g09157 ( new_n9534 , new_n9532 , new_n9533 );
  nand g09158 ( new_n9535 , pi013 , pi024 );
  nand g09159 ( new_n9536 , new_n8598 , new_n8599 );
  nand g09160 ( new_n9537 , new_n8597 , new_n8600 );
  nand g09161 ( new_n9538 , new_n9536 , new_n9537 );
  nand g09162 ( new_n9539 , pi111 , pi112 );
  nand g09163 ( new_n9540 , pi105 , pi210 );
  nand g09164 ( new_n9541 , new_n9539 , new_n9540 );
  nand g09165 ( new_n9542 , pi105 , pi111 );
  or   g09166 ( new_n9543 , new_n8598 , new_n9542 );
  nand g09167 ( new_n9544 , new_n9541 , new_n9543 );
  xor  g09168 ( new_n9545 , new_n9538 , new_n9544 );
  xor  g09169 ( new_n9546 , new_n9535 , new_n9545 );
  nand g09170 ( new_n9547 , pi104 , pi224 );
  nand g09171 ( new_n9548 , pi212 , pi255 );
  nand g09172 ( new_n9549 , new_n9547 , new_n9548 );
  nand g09173 ( new_n9550 , pi104 , pi255 );
  or   g09174 ( new_n9551 , new_n8602 , new_n9550 );
  nand g09175 ( new_n9552 , new_n9549 , new_n9551 );
  xor  g09176 ( new_n9553 , new_n9546 , new_n9552 );
  xor  g09177 ( new_n9554 , new_n9534 , new_n9553 );
  or   g09178 ( new_n9555 , new_n8608 , new_n8611 );
  nand g09179 ( new_n9556 , new_n8607 , new_n8612 );
  nand g09180 ( new_n9557 , new_n9555 , new_n9556 );
  xor  g09181 ( new_n9558 , new_n9554 , new_n9557 );
  nand g09182 ( new_n9559 , new_n8596 , new_n8613 );
  nand g09183 ( new_n9560 , pi127 , pi213 );
  xor  g09184 ( new_n9561 , new_n9559 , new_n9560 );
  xor  g09185 ( new_n9562 , new_n9558 , new_n9561 );
  xor  g09186 ( new_n9563 , new_n9531 , new_n9562 );
  nand g09187 ( new_n9564 , new_n8614 , new_n8618 );
  not  g09188 ( new_n9565 , new_n8595 );
  nand g09189 ( new_n9566 , new_n9565 , new_n8619 );
  nand g09190 ( new_n9567 , new_n9564 , new_n9566 );
  xor  g09191 ( new_n9568 , new_n9563 , new_n9567 );
  nand g09192 ( new_n9569 , new_n9499 , new_n9568 );
  nand g09193 ( new_n9570 , new_n9498 , new_n9569 );
  xor  g09194 ( new_n9571 , new_n9493 , new_n9570 );
  not  g09195 ( new_n9572 , new_n9571 );
  not  g09196 ( new_n9573 , new_n9554 );
  nand g09197 ( new_n9574 , new_n9573 , new_n9557 );
  nand g09198 ( new_n9575 , pi183 , pi210 );
  nand g09199 ( new_n9576 , pi024 , pi112 );
  xor  g09200 ( new_n9577 , new_n9575 , new_n9576 );
  xor  g09201 ( new_n9578 , new_n9542 , new_n9577 );
  not  g09202 ( new_n9579 , new_n9578 );
  nand g09203 ( new_n9580 , pi013 , pi224 );
  xor  g09204 ( new_n9581 , new_n9543 , new_n9580 );
  xor  g09205 ( new_n9582 , new_n9579 , new_n9581 );
  nand g09206 ( new_n9583 , pi127 , pi212 );
  nand g09207 ( new_n9584 , pi213 , pi232 );
  xor  g09208 ( new_n9585 , new_n9583 , new_n9584 );
  xor  g09209 ( new_n9586 , new_n9550 , new_n9585 );
  nand g09210 ( new_n9587 , new_n9538 , new_n9544 );
  nand g09211 ( new_n9588 , new_n9535 , new_n9545 );
  nand g09212 ( new_n9589 , new_n9587 , new_n9588 );
  xor  g09213 ( new_n9590 , new_n9586 , new_n9589 );
  xor  g09214 ( new_n9591 , new_n9582 , new_n9590 );
  nand g09215 ( new_n9592 , new_n9546 , new_n9552 );
  nand g09216 ( new_n9593 , new_n9534 , new_n9553 );
  nand g09217 ( new_n9594 , new_n9592 , new_n9593 );
  xor  g09218 ( new_n9595 , new_n9551 , new_n9594 );
  xnor g09219 ( new_n9596 , new_n9591 , new_n9595 );
  xnor g09220 ( new_n9597 , new_n9574 , new_n9596 );
  nand g09221 ( new_n9598 , new_n9559 , new_n9560 );
  nand g09222 ( new_n9599 , new_n9558 , new_n9561 );
  nand g09223 ( new_n9600 , new_n9598 , new_n9599 );
  xnor g09224 ( new_n9601 , new_n9597 , new_n9600 );
  nand g09225 ( new_n9602 , new_n9523 , new_n9527 );
  nand g09226 ( new_n9603 , pi018 , pi242 );
  nand g09227 ( new_n9604 , pi090 , pi252 );
  xor  g09228 ( new_n9605 , new_n9603 , new_n9604 );
  xor  g09229 ( new_n9606 , new_n9505 , new_n9605 );
  not  g09230 ( new_n9607 , new_n9606 );
  nand g09231 ( new_n9608 , pi121 , pi141 );
  xor  g09232 ( new_n9609 , new_n9506 , new_n9608 );
  xor  g09233 ( new_n9610 , new_n9607 , new_n9609 );
  nand g09234 ( new_n9611 , pi021 , pi236 );
  nand g09235 ( new_n9612 , pi005 , pi241 );
  xor  g09236 ( new_n9613 , new_n9611 , new_n9612 );
  xor  g09237 ( new_n9614 , new_n9516 , new_n9613 );
  nand g09238 ( new_n9615 , new_n9501 , new_n9507 );
  nand g09239 ( new_n9616 , new_n9508 , new_n9511 );
  nand g09240 ( new_n9617 , new_n9615 , new_n9616 );
  xor  g09241 ( new_n9618 , new_n9614 , new_n9617 );
  xor  g09242 ( new_n9619 , new_n9610 , new_n9618 );
  nor  g09243 ( new_n9620 , new_n9519 , new_n9522 );
  nand g09244 ( new_n9621 , new_n9517 , new_n9620 );
  nor  g09245 ( new_n9622 , new_n9512 , new_n9518 );
  or   g09246 ( new_n9623 , new_n9517 , new_n9622 );
  or   g09247 ( new_n9624 , new_n9620 , new_n9623 );
  nand g09248 ( new_n9625 , new_n9621 , new_n9624 );
  xor  g09249 ( new_n9626 , new_n9619 , new_n9625 );
  xor  g09250 ( new_n9627 , new_n9602 , new_n9626 );
  or   g09251 ( new_n9628 , new_n9528 , new_n9529 );
  not  g09252 ( new_n9629 , new_n9500 );
  nand g09253 ( new_n9630 , new_n9629 , new_n9530 );
  nand g09254 ( new_n9631 , new_n9628 , new_n9630 );
  xor  g09255 ( new_n9632 , new_n9627 , new_n9631 );
  not  g09256 ( new_n9633 , new_n9632 );
  xor  g09257 ( new_n9634 , new_n9601 , new_n9633 );
  nand g09258 ( new_n9635 , new_n9531 , new_n9562 );
  nand g09259 ( new_n9636 , new_n9563 , new_n9567 );
  nand g09260 ( new_n9637 , new_n9635 , new_n9636 );
  xor  g09261 ( new_n9638 , new_n9634 , new_n9637 );
  xor  g09262 ( new_n9639 , new_n9572 , new_n9638 );
  xor  g09263 ( new_n9640 , new_n9432 , new_n9639 );
  xor  g09264 ( new_n9641 , new_n9427 , new_n9428 );
  nand g09265 ( new_n9642 , new_n8644 , new_n8664 );
  nand g09266 ( new_n9643 , new_n8665 , new_n8669 );
  nand g09267 ( new_n9644 , new_n9642 , new_n9643 );
  or   g09268 ( new_n9645 , new_n9641 , new_n9644 );
  xnor g09269 ( new_n9646 , new_n9499 , new_n9568 );
  xor  g09270 ( new_n9647 , new_n9641 , new_n9644 );
  nand g09271 ( new_n9648 , new_n9646 , new_n9647 );
  nand g09272 ( new_n9649 , new_n9645 , new_n9648 );
  xor  g09273 ( po062 , new_n9640 , new_n9649 );
  xor  g09274 ( po063 , new_n9164 , new_n9165 );
  nor  g09275 ( new_n9652 , new_n2978 , new_n3080 );
  not  g09276 ( new_n9653 , new_n3081 );
  nor  g09277 ( new_n9654 , new_n9653 , new_n3118 );
  nor  g09278 ( new_n9655 , new_n9652 , new_n9654 );
  nor  g09279 ( new_n9656 , new_n2852 , new_n2875 );
  nor  g09280 ( new_n9657 , new_n2876 , new_n2893 );
  nor  g09281 ( new_n9658 , new_n9656 , new_n9657 );
  nand g09282 ( new_n9659 , pi182 , pi197 );
  nand g09283 ( new_n9660 , new_n2653 , new_n2654 );
  nand g09284 ( new_n9661 , new_n2601 , new_n2655 );
  nand g09285 ( new_n9662 , new_n9660 , new_n9661 );
  or   g09286 ( new_n9663 , new_n2664 , new_n2667 );
  nand g09287 ( new_n9664 , new_n2660 , new_n2668 );
  nand g09288 ( new_n9665 , new_n9663 , new_n9664 );
  xor  g09289 ( new_n9666 , new_n9662 , new_n9665 );
  xor  g09290 ( new_n9667 , new_n9659 , new_n9666 );
  xor  g09291 ( new_n9668 , new_n9658 , new_n9667 );
  xor  g09292 ( new_n9669 , new_n9655 , new_n9668 );
  nand g09293 ( new_n9670 , pi198 , pi216 );
  nand g09294 ( new_n9671 , new_n2794 , new_n2894 );
  nand g09295 ( new_n9672 , new_n2895 , new_n2936 );
  nand g09296 ( new_n9673 , new_n9671 , new_n9672 );
  nand g09297 ( new_n9674 , pi225 , pi229 );
  nand g09298 ( new_n9675 , pi020 , pi030 );
  nand g09299 ( new_n9676 , pi060 , pi185 );
  xor  g09300 ( new_n9677 , new_n9675 , new_n9676 );
  xor  g09301 ( new_n9678 , new_n9674 , new_n9677 );
  xor  g09302 ( new_n9679 , new_n9673 , new_n9678 );
  nand g09303 ( new_n9680 , new_n3051 , new_n3052 );
  nand g09304 ( new_n9681 , new_n3031 , new_n3053 );
  nand g09305 ( new_n9682 , new_n9680 , new_n9681 );
  nand g09306 ( new_n9683 , pi067 , pi101 );
  nand g09307 ( new_n9684 , pi053 , pi223 );
  xor  g09308 ( new_n9685 , new_n9683 , new_n9684 );
  xor  g09309 ( new_n9686 , new_n9682 , new_n9685 );
  nor  g09310 ( new_n9687 , new_n2652 , new_n2676 );
  nor  g09311 ( new_n9688 , new_n2677 , new_n2692 );
  or   g09312 ( new_n9689 , new_n9687 , new_n9688 );
  nand g09313 ( new_n9690 , pi092 , pi177 );
  xor  g09314 ( new_n9691 , new_n9689 , new_n9690 );
  xor  g09315 ( new_n9692 , new_n9686 , new_n9691 );
  nand g09316 ( new_n9693 , new_n3054 , new_n3057 );
  nand g09317 ( new_n9694 , new_n3050 , new_n3058 );
  nand g09318 ( new_n9695 , new_n9693 , new_n9694 );
  nand g09319 ( new_n9696 , pi062 , pi251 );
  nand g09320 ( new_n9697 , pi078 , pi138 );
  xor  g09321 ( new_n9698 , new_n9696 , new_n9697 );
  nand g09322 ( new_n9699 , pi065 , pi192 );
  or   g09323 ( new_n9700 , new_n2669 , new_n2675 );
  nand g09324 ( new_n9701 , new_n2674 , new_n9700 );
  xor  g09325 ( new_n9702 , new_n9699 , new_n9701 );
  xor  g09326 ( new_n9703 , new_n9698 , new_n9702 );
  xor  g09327 ( new_n9704 , new_n9695 , new_n9703 );
  nand g09328 ( new_n9705 , new_n3044 , new_n3045 );
  nand g09329 ( new_n9706 , new_n3019 , new_n3046 );
  nand g09330 ( new_n9707 , new_n9705 , new_n9706 );
  or   g09331 ( new_n9708 , new_n3020 , new_n3048 );
  not  g09332 ( new_n9709 , new_n3047 );
  nand g09333 ( new_n9710 , new_n9709 , new_n3049 );
  nand g09334 ( new_n9711 , new_n9708 , new_n9710 );
  xor  g09335 ( new_n9712 , new_n9707 , new_n9711 );
  xor  g09336 ( new_n9713 , new_n9704 , new_n9712 );
  xor  g09337 ( new_n9714 , new_n9692 , new_n9713 );
  xor  g09338 ( new_n9715 , new_n9679 , new_n9714 );
  xor  g09339 ( new_n9716 , new_n9670 , new_n9715 );
  nor  g09340 ( new_n9717 , new_n2751 , new_n2775 );
  nor  g09341 ( new_n9718 , new_n2776 , new_n2793 );
  nor  g09342 ( new_n9719 , new_n9717 , new_n9718 );
  nor  g09343 ( new_n9720 , new_n3036 , new_n3060 );
  nor  g09344 ( new_n9721 , new_n3061 , new_n3079 );
  nor  g09345 ( new_n9722 , new_n9720 , new_n9721 );
  xor  g09346 ( new_n9723 , new_n9719 , new_n9722 );
  nand g09347 ( new_n9724 , new_n2752 , new_n2753 );
  nand g09348 ( new_n9725 , new_n2706 , new_n2754 );
  nand g09349 ( new_n9726 , new_n9724 , new_n9725 );
  xor  g09350 ( new_n9727 , new_n9723 , new_n9726 );
  nand g09351 ( new_n9728 , pi209 , pi219 );
  nor  g09352 ( new_n9729 , new_n2708 , new_n2756 );
  nor  g09353 ( new_n9730 , new_n2755 , new_n2758 );
  or   g09354 ( new_n9731 , new_n9729 , new_n9730 );
  xor  g09355 ( new_n9732 , new_n9728 , new_n9731 );
  nand g09356 ( new_n9733 , pi123 , pi130 );
  or   g09357 ( new_n9734 , new_n2768 , new_n2774 );
  nand g09358 ( new_n9735 , new_n2773 , new_n9734 );
  nand g09359 ( new_n9736 , pi122 , pi154 );
  nand g09360 ( new_n9737 , pi001 , pi095 );
  xor  g09361 ( new_n9738 , new_n9736 , new_n9737 );
  xor  g09362 ( new_n9739 , new_n9735 , new_n9738 );
  nand g09363 ( new_n9740 , pi089 , pi135 );
  nand g09364 ( new_n9741 , pi087 , pi153 );
  nand g09365 ( new_n9742 , pi059 , pi158 );
  nand g09366 ( new_n9743 , pi094 , pi254 );
  xnor g09367 ( new_n9744 , new_n9742 , new_n9743 );
  xor  g09368 ( new_n9745 , new_n9741 , new_n9744 );
  xor  g09369 ( new_n9746 , new_n9740 , new_n9745 );
  xor  g09370 ( new_n9747 , new_n9739 , new_n9746 );
  xor  g09371 ( new_n9748 , new_n9733 , new_n9747 );
  nand g09372 ( new_n9749 , new_n2853 , new_n2854 );
  nand g09373 ( new_n9750 , new_n2820 , new_n2855 );
  nand g09374 ( new_n9751 , new_n9749 , new_n9750 );
  nand g09375 ( new_n9752 , new_n2861 , new_n2862 );
  nand g09376 ( new_n9753 , new_n2828 , new_n2863 );
  nand g09377 ( new_n9754 , new_n9752 , new_n9753 );
  nor  g09378 ( new_n9755 , new_n2822 , new_n2857 );
  nor  g09379 ( new_n9756 , new_n2856 , new_n2859 );
  or   g09380 ( new_n9757 , new_n9755 , new_n9756 );
  xor  g09381 ( new_n9758 , new_n9754 , new_n9757 );
  xor  g09382 ( new_n9759 , new_n9751 , new_n9758 );
  nand g09383 ( new_n9760 , pi071 , pi215 );
  nand g09384 ( new_n9761 , pi124 , pi169 );
  xor  g09385 ( new_n9762 , new_n9760 , new_n9761 );
  nand g09386 ( new_n9763 , pi003 , pi099 );
  xor  g09387 ( new_n9764 , new_n9762 , new_n9763 );
  xor  g09388 ( new_n9765 , new_n9759 , new_n9764 );
  xor  g09389 ( new_n9766 , new_n9748 , new_n9765 );
  nand g09390 ( new_n9767 , pi006 , pi102 );
  nand g09391 ( new_n9768 , pi137 , pi190 );
  nand g09392 ( new_n9769 , pi160 , pi220 );
  xor  g09393 ( new_n9770 , new_n9768 , new_n9769 );
  or   g09394 ( new_n9771 , new_n3043 , new_n3059 );
  nand g09395 ( new_n9772 , new_n3040 , new_n9771 );
  xor  g09396 ( new_n9773 , new_n9770 , new_n9772 );
  xor  g09397 ( new_n9774 , new_n9767 , new_n9773 );
  xor  g09398 ( new_n9775 , new_n9766 , new_n9774 );
  xor  g09399 ( new_n9776 , new_n9732 , new_n9775 );
  or   g09400 ( new_n9777 , new_n2864 , new_n2867 );
  nand g09401 ( new_n9778 , new_n2860 , new_n2868 );
  nand g09402 ( new_n9779 , new_n9777 , new_n9778 );
  nand g09403 ( new_n9780 , new_n2715 , new_n2761 );
  nand g09404 ( new_n9781 , new_n2760 , new_n2762 );
  nand g09405 ( new_n9782 , new_n9780 , new_n9781 );
  or   g09406 ( new_n9783 , new_n2763 , new_n2766 );
  nand g09407 ( new_n9784 , new_n2759 , new_n2767 );
  nand g09408 ( new_n9785 , new_n9783 , new_n9784 );
  xor  g09409 ( new_n9786 , new_n9782 , new_n9785 );
  xor  g09410 ( new_n9787 , new_n9779 , new_n9786 );
  xor  g09411 ( new_n9788 , new_n9776 , new_n9787 );
  xor  g09412 ( new_n9789 , new_n9727 , new_n9788 );
  nand g09413 ( new_n9790 , pi079 , pi120 );
  nand g09414 ( new_n9791 , pi076 , pi172 );
  xor  g09415 ( new_n9792 , new_n9790 , new_n9791 );
  nand g09416 ( new_n9793 , new_n2829 , new_n2873 );
  nand g09417 ( new_n9794 , new_n2870 , new_n2874 );
  nand g09418 ( new_n9795 , new_n9793 , new_n9794 );
  nand g09419 ( new_n9796 , pi023 , pi073 );
  nand g09420 ( new_n9797 , pi004 , pi155 );
  xor  g09421 ( new_n9798 , new_n9796 , new_n9797 );
  xor  g09422 ( new_n9799 , new_n9795 , new_n9798 );
  nand g09423 ( new_n9800 , pi022 , pi142 );
  nand g09424 ( new_n9801 , new_n2661 , new_n2662 );
  nand g09425 ( new_n9802 , new_n2616 , new_n2663 );
  nand g09426 ( new_n9803 , new_n9801 , new_n9802 );
  xor  g09427 ( new_n9804 , new_n9800 , new_n9803 );
  nand g09428 ( new_n9805 , pi086 , pi170 );
  xor  g09429 ( new_n9806 , new_n9804 , new_n9805 );
  xor  g09430 ( new_n9807 , new_n9799 , new_n9806 );
  xor  g09431 ( new_n9808 , new_n9792 , new_n9807 );
  xor  g09432 ( new_n9809 , new_n9789 , new_n9808 );
  xor  g09433 ( new_n9810 , new_n9716 , new_n9809 );
  or   g09434 ( new_n9811 , new_n2693 , new_n2937 );
  nand g09435 ( new_n9812 , new_n2938 , new_n2977 );
  nand g09436 ( new_n9813 , new_n9811 , new_n9812 );
  nand g09437 ( new_n9814 , pi041 , pi165 );
  or   g09438 ( new_n9815 , new_n2602 , new_n2658 );
  nand g09439 ( new_n9816 , new_n2657 , new_n2659 );
  nand g09440 ( new_n9817 , new_n9815 , new_n9816 );
  xor  g09441 ( new_n9818 , new_n9814 , new_n9817 );
  xor  g09442 ( new_n9819 , new_n9813 , new_n9818 );
  xor  g09443 ( new_n9820 , new_n9810 , new_n9819 );
  xor  g09444 ( po064 , new_n9669 , new_n9820 );
  xor  g09445 ( po065 , new_n9174 , new_n9176 );
  xor  g09446 ( po066 , new_n3101 , new_n3103 );
  xor  g09447 ( po067 , new_n4991 , new_n4992 );
  xor  g09448 ( po068 , new_n6949 , new_n6950 );
  xor  g09449 ( po069 , new_n3822 , new_n3824 );
  xnor g09450 ( po070 , new_n1210 , new_n1211 );
  xor  g09451 ( po071 , new_n9180 , new_n9182 );
  nand g09452 ( new_n9829 , pi007 , pi141 );
  or   g09453 ( new_n9830 , new_n6386 , new_n9829 );
  nand g09454 ( new_n9831 , pi018 , pi051 );
  nand g09455 ( new_n9832 , pi090 , pi108 );
  xor  g09456 ( new_n9833 , new_n9831 , new_n9832 );
  xor  g09457 ( new_n9834 , new_n6385 , new_n9833 );
  not  g09458 ( new_n9835 , new_n9834 );
  xor  g09459 ( new_n9836 , new_n6386 , new_n9829 );
  nand g09460 ( new_n9837 , new_n9835 , new_n9836 );
  nand g09461 ( new_n9838 , new_n9830 , new_n9837 );
  nand g09462 ( new_n9839 , new_n6405 , new_n6406 );
  nand g09463 ( new_n9840 , new_n6404 , new_n6407 );
  nand g09464 ( new_n9841 , new_n9839 , new_n9840 );
  nand g09465 ( new_n9842 , new_n6399 , new_n6403 );
  xor  g09466 ( new_n9843 , new_n9834 , new_n9836 );
  nand g09467 ( new_n9844 , pi113 , pi241 );
  nand g09468 ( new_n9845 , pi038 , pi236 );
  xor  g09469 ( new_n9846 , new_n9844 , new_n9845 );
  xor  g09470 ( new_n9847 , new_n6392 , new_n9846 );
  nor  g09471 ( new_n9848 , new_n6377 , new_n6380 );
  nor  g09472 ( new_n9849 , new_n6381 , new_n6387 );
  nor  g09473 ( new_n9850 , new_n9848 , new_n9849 );
  xor  g09474 ( new_n9851 , new_n9847 , new_n9850 );
  xnor g09475 ( new_n9852 , new_n9843 , new_n9851 );
  nor  g09476 ( new_n9853 , new_n6388 , new_n6394 );
  nor  g09477 ( new_n9854 , new_n6395 , new_n6398 );
  xor  g09478 ( new_n9855 , new_n6393 , new_n9854 );
  nor  g09479 ( new_n9856 , new_n9853 , new_n9855 );
  xor  g09480 ( new_n9857 , new_n9852 , new_n9856 );
  xor  g09481 ( new_n9858 , new_n9842 , new_n9857 );
  xnor g09482 ( new_n9859 , new_n9841 , new_n9858 );
  nand g09483 ( new_n9860 , new_n6432 , new_n6435 );
  nand g09484 ( new_n9861 , pi183 , pi188 );
  nand g09485 ( new_n9862 , pi061 , pi112 );
  xor  g09486 ( new_n9863 , new_n9861 , new_n9862 );
  xor  g09487 ( new_n9864 , new_n6414 , new_n9863 );
  nand g09488 ( new_n9865 , pi012 , pi013 );
  xor  g09489 ( new_n9866 , new_n6415 , new_n9865 );
  xor  g09490 ( new_n9867 , new_n9864 , new_n9866 );
  nand g09491 ( new_n9868 , pi098 , pi212 );
  nand g09492 ( new_n9869 , pi043 , pi213 );
  xor  g09493 ( new_n9870 , new_n9868 , new_n9869 );
  xor  g09494 ( new_n9871 , new_n6425 , new_n9870 );
  nand g09495 ( new_n9872 , new_n6410 , new_n6416 );
  nand g09496 ( new_n9873 , new_n6417 , new_n6420 );
  nand g09497 ( new_n9874 , new_n9872 , new_n9873 );
  xor  g09498 ( new_n9875 , new_n9871 , new_n9874 );
  xnor g09499 ( new_n9876 , new_n9867 , new_n9875 );
  nor  g09500 ( new_n9877 , new_n6421 , new_n6427 );
  nor  g09501 ( new_n9878 , new_n6428 , new_n6431 );
  xor  g09502 ( new_n9879 , new_n6426 , new_n9878 );
  nor  g09503 ( new_n9880 , new_n9877 , new_n9879 );
  not  g09504 ( new_n9881 , new_n9880 );
  xor  g09505 ( new_n9882 , new_n9876 , new_n9881 );
  xor  g09506 ( new_n9883 , new_n9860 , new_n9882 );
  nand g09507 ( new_n9884 , new_n6436 , new_n6437 );
  nand g09508 ( new_n9885 , new_n6409 , new_n6438 );
  nand g09509 ( new_n9886 , new_n9884 , new_n9885 );
  xor  g09510 ( new_n9887 , new_n9883 , new_n9886 );
  xor  g09511 ( new_n9888 , new_n9859 , new_n9887 );
  not  g09512 ( new_n9889 , new_n6439 );
  nor  g09513 ( new_n9890 , new_n6408 , new_n9889 );
  nor  g09514 ( new_n9891 , new_n6440 , new_n6444 );
  nor  g09515 ( new_n9892 , new_n9890 , new_n9891 );
  xor  g09516 ( new_n9893 , new_n9888 , new_n9892 );
  nand g09517 ( new_n9894 , new_n6468 , new_n6472 );
  nand g09518 ( new_n9895 , pi015 , pi179 );
  nand g09519 ( new_n9896 , pi146 , pi162 );
  xor  g09520 ( new_n9897 , new_n9895 , new_n9896 );
  xor  g09521 ( new_n9898 , new_n6450 , new_n9897 );
  not  g09522 ( new_n9899 , new_n9898 );
  nand g09523 ( new_n9900 , pi035 , pi048 );
  xor  g09524 ( new_n9901 , new_n6451 , new_n9900 );
  xor  g09525 ( new_n9902 , new_n9899 , new_n9901 );
  nand g09526 ( new_n9903 , pi168 , pi193 );
  nand g09527 ( new_n9904 , pi208 , pi238 );
  xor  g09528 ( new_n9905 , new_n9903 , new_n9904 );
  xor  g09529 ( new_n9906 , new_n6461 , new_n9905 );
  nand g09530 ( new_n9907 , new_n6446 , new_n6452 );
  nand g09531 ( new_n9908 , new_n6453 , new_n6456 );
  nand g09532 ( new_n9909 , new_n9907 , new_n9908 );
  xor  g09533 ( new_n9910 , new_n9906 , new_n9909 );
  xor  g09534 ( new_n9911 , new_n9902 , new_n9910 );
  nor  g09535 ( new_n9912 , new_n6464 , new_n6467 );
  nand g09536 ( new_n9913 , new_n6462 , new_n9912 );
  nor  g09537 ( new_n9914 , new_n6457 , new_n6463 );
  or   g09538 ( new_n9915 , new_n6462 , new_n9914 );
  or   g09539 ( new_n9916 , new_n9912 , new_n9915 );
  nand g09540 ( new_n9917 , new_n9913 , new_n9916 );
  xor  g09541 ( new_n9918 , new_n9911 , new_n9917 );
  xnor g09542 ( new_n9919 , new_n9894 , new_n9918 );
  nand g09543 ( new_n9920 , new_n6474 , new_n6475 );
  nand g09544 ( new_n9921 , new_n6473 , new_n6476 );
  nand g09545 ( new_n9922 , new_n9920 , new_n9921 );
  xor  g09546 ( new_n9923 , new_n9919 , new_n9922 );
  nor  g09547 ( new_n9924 , new_n9893 , new_n9923 );
  or   g09548 ( new_n9925 , new_n6477 , new_n6480 );
  nand g09549 ( new_n9926 , new_n6445 , new_n6481 );
  nand g09550 ( new_n9927 , new_n9925 , new_n9926 );
  xnor g09551 ( new_n9928 , new_n9893 , new_n9923 );
  nor  g09552 ( new_n9929 , new_n9927 , new_n9928 );
  nor  g09553 ( new_n9930 , new_n9924 , new_n9929 );
  nand g09554 ( new_n9931 , pi064 , pi194 );
  nand g09555 ( new_n9932 , pi052 , pi068 );
  nand g09556 ( new_n9933 , pi036 , pi077 );
  xor  g09557 ( new_n9934 , new_n9932 , new_n9933 );
  xor  g09558 ( new_n9935 , new_n9931 , new_n9934 );
  xor  g09559 ( new_n9936 , new_n9930 , new_n9935 );
  nand g09560 ( new_n9937 , pi068 , pi131 );
  nand g09561 ( new_n9938 , pi036 , pi052 );
  nand g09562 ( new_n9939 , new_n9937 , new_n9938 );
  xor  g09563 ( new_n9940 , new_n9937 , new_n9938 );
  nand g09564 ( new_n9941 , new_n6498 , new_n9940 );
  nand g09565 ( new_n9942 , new_n9939 , new_n9941 );
  xor  g09566 ( new_n9943 , new_n6498 , new_n9940 );
  nand g09567 ( new_n9944 , new_n6483 , new_n6489 );
  nand g09568 ( new_n9945 , new_n6490 , new_n6493 );
  nand g09569 ( new_n9946 , new_n9944 , new_n9945 );
  or   g09570 ( new_n9947 , new_n9943 , new_n9946 );
  nand g09571 ( new_n9948 , pi189 , pi194 );
  nand g09572 ( new_n9949 , pi084 , pi143 );
  xor  g09573 ( new_n9950 , new_n9948 , new_n9949 );
  xor  g09574 ( new_n9951 , new_n6487 , new_n9950 );
  not  g09575 ( new_n9952 , new_n9951 );
  nand g09576 ( new_n9953 , pi085 , pi133 );
  xor  g09577 ( new_n9954 , new_n6488 , new_n9953 );
  xor  g09578 ( new_n9955 , new_n9952 , new_n9954 );
  xor  g09579 ( new_n9956 , new_n9943 , new_n9946 );
  nand g09580 ( new_n9957 , new_n9955 , new_n9956 );
  nand g09581 ( new_n9958 , new_n9947 , new_n9957 );
  xor  g09582 ( new_n9959 , new_n9942 , new_n9958 );
  nand g09583 ( new_n9960 , pi085 , pi189 );
  nand g09584 ( new_n9961 , pi133 , pi180 );
  xor  g09585 ( new_n9962 , new_n9960 , new_n9961 );
  xor  g09586 ( new_n9963 , new_n9959 , new_n9962 );
  nor  g09587 ( new_n9964 , new_n9894 , new_n9918 );
  nor  g09588 ( new_n9965 , new_n9919 , new_n9922 );
  nor  g09589 ( new_n9966 , new_n9964 , new_n9965 );
  nand g09590 ( new_n9967 , pi057 , pi084 );
  xor  g09591 ( new_n9968 , new_n9966 , new_n9967 );
  xor  g09592 ( new_n9969 , new_n9963 , new_n9968 );
  nand g09593 ( new_n9970 , pi159 , pi168 );
  nand g09594 ( new_n9971 , pi033 , pi146 );
  nand g09595 ( new_n9972 , pi152 , pi162 );
  or   g09596 ( new_n9973 , new_n9911 , new_n9917 );
  nand g09597 ( new_n9974 , new_n9916 , new_n9973 );
  xor  g09598 ( new_n9975 , new_n9972 , new_n9974 );
  xor  g09599 ( new_n9976 , new_n9971 , new_n9975 );
  xor  g09600 ( new_n9977 , new_n9970 , new_n9976 );
  nand g09601 ( new_n9978 , new_n9948 , new_n9949 );
  nand g09602 ( new_n9979 , new_n6487 , new_n9950 );
  nand g09603 ( new_n9980 , new_n9978 , new_n9979 );
  or   g09604 ( new_n9981 , new_n6488 , new_n9953 );
  nand g09605 ( new_n9982 , new_n9952 , new_n9954 );
  nand g09606 ( new_n9983 , new_n9981 , new_n9982 );
  xor  g09607 ( new_n9984 , new_n9980 , new_n9983 );
  xor  g09608 ( new_n9985 , new_n9977 , new_n9984 );
  xor  g09609 ( new_n9986 , new_n9969 , new_n9985 );
  xor  g09610 ( new_n9987 , new_n9936 , new_n9986 );
  nand g09611 ( new_n9988 , pi013 , pi144 );
  nand g09612 ( new_n9989 , new_n9871 , new_n9874 );
  nand g09613 ( new_n9990 , new_n9867 , new_n9875 );
  nand g09614 ( new_n9991 , new_n9989 , new_n9990 );
  xor  g09615 ( new_n9992 , new_n9988 , new_n9991 );
  nand g09616 ( new_n9993 , pi012 , pi112 );
  xor  g09617 ( new_n9994 , new_n9992 , new_n9993 );
  xor  g09618 ( new_n9995 , new_n9987 , new_n9994 );
  or   g09619 ( new_n9996 , new_n6451 , new_n9900 );
  nand g09620 ( new_n9997 , new_n9899 , new_n9901 );
  nand g09621 ( new_n9998 , new_n9996 , new_n9997 );
  nand g09622 ( new_n9999 , pi035 , pi237 );
  nand g09623 ( new_n10000 , pi139 , pi238 );
  xor  g09624 ( new_n10001 , new_n9999 , new_n10000 );
  xor  g09625 ( new_n10002 , new_n9998 , new_n10001 );
  nand g09626 ( new_n10003 , new_n6426 , new_n9878 );
  nand g09627 ( new_n10004 , new_n9876 , new_n9881 );
  nand g09628 ( new_n10005 , new_n10003 , new_n10004 );
  nand g09629 ( new_n10006 , pi179 , pi204 );
  xor  g09630 ( new_n10007 , new_n10005 , new_n10006 );
  xor  g09631 ( new_n10008 , new_n10002 , new_n10007 );
  or   g09632 ( new_n10009 , new_n9906 , new_n9909 );
  nand g09633 ( new_n10010 , new_n9902 , new_n9910 );
  nand g09634 ( new_n10011 , new_n10009 , new_n10010 );
  nand g09635 ( new_n10012 , new_n9895 , new_n9896 );
  nand g09636 ( new_n10013 , new_n6450 , new_n9897 );
  nand g09637 ( new_n10014 , new_n10012 , new_n10013 );
  xor  g09638 ( new_n10015 , new_n10011 , new_n10014 );
  xor  g09639 ( new_n10016 , new_n10008 , new_n10015 );
  nand g09640 ( new_n10017 , new_n9861 , new_n9862 );
  nand g09641 ( new_n10018 , new_n6414 , new_n9863 );
  nand g09642 ( new_n10019 , new_n10017 , new_n10018 );
  or   g09643 ( new_n10020 , new_n6415 , new_n9865 );
  not  g09644 ( new_n10021 , new_n9864 );
  nand g09645 ( new_n10022 , new_n10021 , new_n9866 );
  nand g09646 ( new_n10023 , new_n10020 , new_n10022 );
  xor  g09647 ( new_n10024 , new_n10019 , new_n10023 );
  nand g09648 ( new_n10025 , new_n9859 , new_n9887 );
  nand g09649 ( new_n10026 , new_n9888 , new_n9892 );
  nand g09650 ( new_n10027 , new_n10025 , new_n10026 );
  nand g09651 ( new_n10028 , pi126 , pi213 );
  xor  g09652 ( new_n10029 , new_n10027 , new_n10028 );
  nand g09653 ( new_n10030 , new_n9903 , new_n9904 );
  nand g09654 ( new_n10031 , new_n6461 , new_n9905 );
  nand g09655 ( new_n10032 , new_n10030 , new_n10031 );
  nand g09656 ( new_n10033 , pi088 , pi188 );
  not  g09657 ( new_n10034 , new_n9882 );
  nor  g09658 ( new_n10035 , new_n9860 , new_n10034 );
  nor  g09659 ( new_n10036 , new_n9883 , new_n9886 );
  or   g09660 ( new_n10037 , new_n10035 , new_n10036 );
  nand g09661 ( new_n10038 , pi178 , pi183 );
  nand g09662 ( new_n10039 , pi061 , pi105 );
  xor  g09663 ( new_n10040 , new_n10038 , new_n10039 );
  xor  g09664 ( new_n10041 , new_n10037 , new_n10040 );
  xor  g09665 ( new_n10042 , new_n10033 , new_n10041 );
  xor  g09666 ( new_n10043 , new_n10032 , new_n10042 );
  xor  g09667 ( new_n10044 , new_n10029 , new_n10043 );
  nand g09668 ( new_n10045 , pi193 , pi208 );
  nand g09669 ( new_n10046 , pi015 , pi048 );
  xor  g09670 ( new_n10047 , new_n10045 , new_n10046 );
  xor  g09671 ( new_n10048 , new_n10044 , new_n10047 );
  xor  g09672 ( new_n10049 , new_n10024 , new_n10048 );
  xor  g09673 ( new_n10050 , new_n10016 , new_n10049 );
  nand g09674 ( new_n10051 , new_n9868 , new_n9869 );
  nand g09675 ( new_n10052 , new_n6425 , new_n9870 );
  nand g09676 ( new_n10053 , new_n10051 , new_n10052 );
  nand g09677 ( new_n10054 , new_n9842 , new_n9857 );
  nand g09678 ( new_n10055 , new_n9841 , new_n9858 );
  nand g09679 ( new_n10056 , new_n10054 , new_n10055 );
  xor  g09680 ( new_n10057 , new_n10053 , new_n10056 );
  nand g09681 ( new_n10058 , pi043 , pi212 );
  nand g09682 ( new_n10059 , pi098 , pi104 );
  xor  g09683 ( new_n10060 , new_n10058 , new_n10059 );
  nand g09684 ( new_n10061 , new_n6393 , new_n9854 );
  not  g09685 ( new_n10062 , new_n9856 );
  nand g09686 ( new_n10063 , new_n9852 , new_n10062 );
  nand g09687 ( new_n10064 , new_n10061 , new_n10063 );
  nand g09688 ( new_n10065 , pi007 , pi090 );
  nand g09689 ( new_n10066 , pi118 , pi141 );
  xor  g09690 ( new_n10067 , new_n10065 , new_n10066 );
  xor  g09691 ( new_n10068 , new_n10064 , new_n10067 );
  nand g09692 ( new_n10069 , pi047 , pi108 );
  nand g09693 ( new_n10070 , pi028 , pi236 );
  nand g09694 ( new_n10071 , pi018 , pi042 );
  nand g09695 ( new_n10072 , pi051 , pi128 );
  xnor g09696 ( new_n10073 , new_n10071 , new_n10072 );
  xor  g09697 ( new_n10074 , new_n10070 , new_n10073 );
  xor  g09698 ( new_n10075 , new_n10069 , new_n10074 );
  xor  g09699 ( new_n10076 , new_n10068 , new_n10075 );
  xor  g09700 ( new_n10077 , new_n10060 , new_n10076 );
  xor  g09701 ( new_n10078 , new_n10057 , new_n10077 );
  xor  g09702 ( new_n10079 , new_n10050 , new_n10078 );
  xor  g09703 ( new_n10080 , new_n9995 , new_n10079 );
  xor  g09704 ( new_n10081 , new_n9838 , new_n10080 );
  nand g09705 ( new_n10082 , new_n9831 , new_n9832 );
  nand g09706 ( new_n10083 , new_n6385 , new_n9833 );
  nand g09707 ( new_n10084 , new_n10082 , new_n10083 );
  xor  g09708 ( new_n10085 , new_n9927 , new_n9928 );
  nand g09709 ( new_n10086 , new_n6506 , new_n6509 );
  xor  g09710 ( new_n10087 , new_n9955 , new_n9956 );
  nor  g09711 ( new_n10088 , new_n6502 , new_n6505 );
  and  g09712 ( new_n10089 , new_n6499 , new_n10088 );
  or   g09713 ( new_n10090 , new_n6494 , new_n6501 );
  nand g09714 ( new_n10091 , new_n6500 , new_n10090 );
  nor  g09715 ( new_n10092 , new_n10088 , new_n10091 );
  or   g09716 ( new_n10093 , new_n10089 , new_n10092 );
  xor  g09717 ( new_n10094 , new_n10087 , new_n10093 );
  xnor g09718 ( new_n10095 , new_n10086 , new_n10094 );
  nand g09719 ( new_n10096 , new_n6511 , new_n6512 );
  nand g09720 ( new_n10097 , new_n6510 , new_n6513 );
  nand g09721 ( new_n10098 , new_n10096 , new_n10097 );
  xor  g09722 ( new_n10099 , new_n10095 , new_n10098 );
  not  g09723 ( new_n10100 , new_n10099 );
  nor  g09724 ( new_n10101 , new_n10085 , new_n10100 );
  xor  g09725 ( new_n10102 , new_n10085 , new_n10099 );
  nand g09726 ( new_n10103 , new_n6514 , new_n6518 );
  not  g09727 ( new_n10104 , new_n6482 );
  nand g09728 ( new_n10105 , new_n10104 , new_n6519 );
  nand g09729 ( new_n10106 , new_n10103 , new_n10105 );
  nor  g09730 ( new_n10107 , new_n10102 , new_n10106 );
  nor  g09731 ( new_n10108 , new_n10101 , new_n10107 );
  nand g09732 ( new_n10109 , new_n9847 , new_n9850 );
  nand g09733 ( new_n10110 , new_n9843 , new_n9851 );
  nand g09734 ( new_n10111 , new_n10109 , new_n10110 );
  nand g09735 ( new_n10112 , new_n9844 , new_n9845 );
  nand g09736 ( new_n10113 , new_n6392 , new_n9846 );
  nand g09737 ( new_n10114 , new_n10112 , new_n10113 );
  xor  g09738 ( new_n10115 , new_n10111 , new_n10114 );
  xor  g09739 ( new_n10116 , new_n10108 , new_n10115 );
  xor  g09740 ( new_n10117 , new_n10084 , new_n10116 );
  nand g09741 ( new_n10118 , pi038 , pi241 );
  nand g09742 ( new_n10119 , pi113 , pi161 );
  xor  g09743 ( new_n10120 , new_n10118 , new_n10119 );
  nand g09744 ( new_n10121 , pi034 , pi143 );
  nand g09745 ( new_n10122 , pi046 , pi131 );
  xor  g09746 ( new_n10123 , new_n10121 , new_n10122 );
  nor  g09747 ( new_n10124 , new_n10087 , new_n10093 );
  nor  g09748 ( new_n10125 , new_n10092 , new_n10124 );
  nor  g09749 ( new_n10126 , new_n10086 , new_n10094 );
  nor  g09750 ( new_n10127 , new_n10095 , new_n10098 );
  nor  g09751 ( new_n10128 , new_n10126 , new_n10127 );
  xor  g09752 ( new_n10129 , new_n10125 , new_n10128 );
  xor  g09753 ( new_n10130 , new_n10123 , new_n10129 );
  xor  g09754 ( new_n10131 , new_n10120 , new_n10130 );
  xor  g09755 ( new_n10132 , new_n10117 , new_n10131 );
  xor  g09756 ( po072 , new_n10081 , new_n10132 );
  xor  g09757 ( po073 , new_n894 , new_n895 );
  xor  g09758 ( po074 , new_n6198 , new_n6202 );
  xor  g09759 ( po075 , new_n7511 , new_n7532 );
  xor  g09760 ( po076 , new_n6601 , new_n6602 );
  xor  g09761 ( po077 , new_n1190 , new_n1196 );
  xor  g09762 ( po078 , new_n1831 , new_n1832 );
  xor  g09763 ( po079 , new_n5673 , new_n5675 );
  xnor g09764 ( po080 , new_n9169 , new_n9170 );
  xor  g09765 ( po081 , new_n7526 , new_n7528 );
  xor  g09766 ( po082 , new_n6192 , new_n6204 );
  xor  g09767 ( po083 , new_n1202 , new_n1204 );
  not  g09768 ( new_n10145 , new_n722 );
  nand g09769 ( new_n10146 , new_n622 , new_n10145 );
  or   g09770 ( new_n10147 , new_n723 , new_n760 );
  nand g09771 ( new_n10148 , new_n10146 , new_n10147 );
  nand g09772 ( new_n10149 , pi097 , pi167 );
  nand g09773 ( new_n10150 , pi134 , pi166 );
  nand g09774 ( new_n10151 , new_n682 , new_n683 );
  nand g09775 ( new_n10152 , new_n628 , new_n684 );
  nand g09776 ( new_n10153 , new_n10151 , new_n10152 );
  xor  g09777 ( new_n10154 , new_n10150 , new_n10153 );
  xor  g09778 ( new_n10155 , new_n10149 , new_n10154 );
  xor  g09779 ( new_n10156 , new_n10148 , new_n10155 );
  nand g09780 ( new_n10157 , new_n689 , new_n690 );
  nand g09781 ( new_n10158 , new_n643 , new_n691 );
  nand g09782 ( new_n10159 , new_n10157 , new_n10158 );
  nand g09783 ( new_n10160 , pi075 , pi149 );
  nand g09784 ( new_n10161 , pi093 , pi240 );
  xor  g09785 ( new_n10162 , new_n10160 , new_n10161 );
  xor  g09786 ( new_n10163 , new_n10159 , new_n10162 );
  nand g09787 ( new_n10164 , pi019 , pi181 );
  nand g09788 ( new_n10165 , pi000 , pi164 );
  nand g09789 ( new_n10166 , pi115 , pi206 );
  nand g09790 ( new_n10167 , pi032 , pi070 );
  xor  g09791 ( new_n10168 , new_n10166 , new_n10167 );
  nand g09792 ( new_n10169 , pi031 , pi163 );
  nand g09793 ( new_n10170 , new_n483 , new_n580 );
  not  g09794 ( new_n10171 , new_n621 );
  nand g09795 ( new_n10172 , new_n581 , new_n10171 );
  nand g09796 ( new_n10173 , new_n10170 , new_n10172 );
  xor  g09797 ( new_n10174 , new_n10169 , new_n10173 );
  xor  g09798 ( new_n10175 , new_n10168 , new_n10174 );
  xor  g09799 ( new_n10176 , new_n10165 , new_n10175 );
  xor  g09800 ( new_n10177 , new_n10164 , new_n10176 );
  xor  g09801 ( new_n10178 , new_n10163 , new_n10177 );
  nand g09802 ( new_n10179 , new_n505 , new_n558 );
  nand g09803 ( new_n10180 , new_n556 , new_n561 );
  nand g09804 ( new_n10181 , new_n10179 , new_n10180 );
  not  g09805 ( new_n10182 , new_n562 );
  nor  g09806 ( new_n10183 , new_n540 , new_n10182 );
  nor  g09807 ( new_n10184 , new_n563 , new_n579 );
  nor  g09808 ( new_n10185 , new_n10183 , new_n10184 );
  xor  g09809 ( new_n10186 , new_n10181 , new_n10185 );
  or   g09810 ( new_n10187 , new_n629 , new_n686 );
  not  g09811 ( new_n10188 , new_n685 );
  nand g09812 ( new_n10189 , new_n10188 , new_n687 );
  nand g09813 ( new_n10190 , new_n10187 , new_n10189 );
  nand g09814 ( new_n10191 , new_n692 , new_n695 );
  nand g09815 ( new_n10192 , new_n688 , new_n696 );
  nand g09816 ( new_n10193 , new_n10191 , new_n10192 );
  xor  g09817 ( new_n10194 , new_n10190 , new_n10193 );
  xor  g09818 ( new_n10195 , new_n10186 , new_n10194 );
  xor  g09819 ( new_n10196 , new_n10178 , new_n10195 );
  xor  g09820 ( new_n10197 , new_n10156 , new_n10196 );
  nand g09821 ( new_n10198 , pi234 , pi250 );
  nand g09822 ( new_n10199 , new_n820 , new_n821 );
  nand g09823 ( new_n10200 , new_n774 , new_n822 );
  nand g09824 ( new_n10201 , new_n10199 , new_n10200 );
  xor  g09825 ( new_n10202 , new_n10198 , new_n10201 );
  xor  g09826 ( new_n10203 , new_n10197 , new_n10202 );
  nand g09827 ( new_n10204 , new_n783 , new_n829 );
  nand g09828 ( new_n10205 , new_n828 , new_n830 );
  nand g09829 ( new_n10206 , new_n10204 , new_n10205 );
  nand g09830 ( new_n10207 , pi044 , pi247 );
  nand g09831 ( new_n10208 , pi054 , pi080 );
  xor  g09832 ( new_n10209 , new_n10207 , new_n10208 );
  xor  g09833 ( new_n10210 , new_n10206 , new_n10209 );
  or   g09834 ( new_n10211 , new_n681 , new_n702 );
  nand g09835 ( new_n10212 , new_n703 , new_n721 );
  nand g09836 ( new_n10213 , new_n10211 , new_n10212 );
  nand g09837 ( new_n10214 , pi045 , pi214 );
  xor  g09838 ( new_n10215 , new_n10213 , new_n10214 );
  xor  g09839 ( new_n10216 , new_n10210 , new_n10215 );
  nand g09840 ( new_n10217 , pi151 , pi200 );
  nand g09841 ( new_n10218 , pi147 , pi203 );
  nand g09842 ( new_n10219 , new_n644 , new_n699 );
  not  g09843 ( new_n10220 , new_n701 );
  nand g09844 ( new_n10221 , new_n697 , new_n10220 );
  nand g09845 ( new_n10222 , new_n10219 , new_n10221 );
  xor  g09846 ( new_n10223 , new_n10218 , new_n10222 );
  xor  g09847 ( new_n10224 , new_n10217 , new_n10223 );
  nand g09848 ( new_n10225 , pi011 , pi175 );
  or   g09849 ( new_n10226 , new_n831 , new_n834 );
  nand g09850 ( new_n10227 , new_n827 , new_n835 );
  nand g09851 ( new_n10228 , new_n10226 , new_n10227 );
  xor  g09852 ( new_n10229 , new_n10225 , new_n10228 );
  xor  g09853 ( new_n10230 , new_n10224 , new_n10229 );
  nand g09854 ( new_n10231 , pi016 , pi072 );
  nand g09855 ( new_n10232 , pi117 , pi248 );
  nor  g09856 ( new_n10233 , new_n776 , new_n824 );
  nor  g09857 ( new_n10234 , new_n823 , new_n826 );
  or   g09858 ( new_n10235 , new_n10233 , new_n10234 );
  xor  g09859 ( new_n10236 , new_n10232 , new_n10235 );
  xor  g09860 ( new_n10237 , new_n10231 , new_n10236 );
  xor  g09861 ( new_n10238 , new_n10230 , new_n10237 );
  xor  g09862 ( new_n10239 , new_n10216 , new_n10238 );
  xor  g09863 ( new_n10240 , new_n10203 , new_n10239 );
  or   g09864 ( new_n10241 , new_n836 , new_n842 );
  nand g09865 ( new_n10242 , new_n841 , new_n10241 );
  nand g09866 ( new_n10243 , new_n443 , new_n444 );
  nand g09867 ( new_n10244 , new_n389 , new_n445 );
  nand g09868 ( new_n10245 , new_n10243 , new_n10244 );
  xor  g09869 ( new_n10246 , new_n10242 , new_n10245 );
  xor  g09870 ( new_n10247 , new_n10240 , new_n10246 );
  nor  g09871 ( new_n10248 , new_n819 , new_n843 );
  nor  g09872 ( new_n10249 , new_n844 , new_n861 );
  nor  g09873 ( new_n10250 , new_n10248 , new_n10249 );
  nand g09874 ( new_n10251 , new_n451 , new_n452 );
  nand g09875 ( new_n10252 , new_n416 , new_n453 );
  nand g09876 ( new_n10253 , new_n10251 , new_n10252 );
  nand g09877 ( new_n10254 , pi049 , pi096 );
  xor  g09878 ( new_n10255 , new_n10253 , new_n10254 );
  xor  g09879 ( new_n10256 , new_n10250 , new_n10255 );
  nand g09880 ( new_n10257 , new_n761 , new_n863 );
  nand g09881 ( new_n10258 , new_n864 , new_n903 );
  nand g09882 ( new_n10259 , new_n10257 , new_n10258 );
  nand g09883 ( new_n10260 , pi119 , pi202 );
  nand g09884 ( new_n10261 , pi009 , pi103 );
  xor  g09885 ( new_n10262 , new_n10260 , new_n10261 );
  or   g09886 ( new_n10263 , new_n390 , new_n448 );
  nand g09887 ( new_n10264 , new_n447 , new_n449 );
  nand g09888 ( new_n10265 , new_n10263 , new_n10264 );
  xor  g09889 ( new_n10266 , new_n10262 , new_n10265 );
  xor  g09890 ( new_n10267 , new_n10259 , new_n10266 );
  xor  g09891 ( new_n10268 , new_n10256 , new_n10267 );
  nor  g09892 ( new_n10269 , new_n442 , new_n464 );
  nor  g09893 ( new_n10270 , new_n465 , new_n482 );
  nor  g09894 ( new_n10271 , new_n10269 , new_n10270 );
  nand g09895 ( new_n10272 , pi056 , pi201 );
  nand g09896 ( new_n10273 , pi136 , pi245 );
  xor  g09897 ( new_n10274 , new_n10272 , new_n10273 );
  xor  g09898 ( new_n10275 , new_n10271 , new_n10274 );
  nand g09899 ( new_n10276 , pi107 , pi110 );
  nand g09900 ( new_n10277 , pi027 , pi083 );
  nand g09901 ( new_n10278 , pi026 , pi063 );
  nand g09902 ( new_n10279 , pi008 , pi156 );
  xor  g09903 ( new_n10280 , new_n10278 , new_n10279 );
  nand g09904 ( new_n10281 , new_n541 , new_n542 );
  nand g09905 ( new_n10282 , new_n489 , new_n543 );
  nand g09906 ( new_n10283 , new_n10281 , new_n10282 );
  nand g09907 ( new_n10284 , new_n548 , new_n549 );
  nand g09908 ( new_n10285 , new_n504 , new_n550 );
  nand g09909 ( new_n10286 , new_n10284 , new_n10285 );
  xor  g09910 ( new_n10287 , new_n10283 , new_n10286 );
  nand g09911 ( new_n10288 , pi116 , pi145 );
  xor  g09912 ( new_n10289 , new_n10287 , new_n10288 );
  or   g09913 ( new_n10290 , new_n490 , new_n545 );
  not  g09914 ( new_n10291 , new_n544 );
  nand g09915 ( new_n10292 , new_n10291 , new_n546 );
  nand g09916 ( new_n10293 , new_n10290 , new_n10292 );
  or   g09917 ( new_n10294 , new_n417 , new_n462 );
  nand g09918 ( new_n10295 , new_n459 , new_n463 );
  nand g09919 ( new_n10296 , new_n10294 , new_n10295 );
  xor  g09920 ( new_n10297 , new_n10293 , new_n10296 );
  nand g09921 ( new_n10298 , pi091 , pi148 );
  nand g09922 ( new_n10299 , pi114 , pi228 );
  xor  g09923 ( new_n10300 , new_n10298 , new_n10299 );
  nand g09924 ( new_n10301 , pi039 , pi246 );
  nand g09925 ( new_n10302 , new_n551 , new_n554 );
  nand g09926 ( new_n10303 , new_n547 , new_n555 );
  nand g09927 ( new_n10304 , new_n10302 , new_n10303 );
  xnor g09928 ( new_n10305 , new_n10301 , new_n10304 );
  xor  g09929 ( new_n10306 , new_n10300 , new_n10305 );
  xor  g09930 ( new_n10307 , new_n10297 , new_n10306 );
  xor  g09931 ( new_n10308 , new_n10289 , new_n10307 );
  xor  g09932 ( new_n10309 , new_n10280 , new_n10308 );
  xor  g09933 ( new_n10310 , new_n10277 , new_n10309 );
  xor  g09934 ( new_n10311 , new_n10276 , new_n10310 );
  xor  g09935 ( new_n10312 , new_n10275 , new_n10311 );
  nand g09936 ( new_n10313 , pi171 , pi235 );
  nand g09937 ( new_n10314 , new_n454 , new_n457 );
  not  g09938 ( new_n10315 , new_n450 );
  nand g09939 ( new_n10316 , new_n10315 , new_n458 );
  nand g09940 ( new_n10317 , new_n10314 , new_n10316 );
  xor  g09941 ( new_n10318 , new_n10313 , new_n10317 );
  xor  g09942 ( new_n10319 , new_n10312 , new_n10318 );
  xor  g09943 ( new_n10320 , new_n10268 , new_n10319 );
  xor  g09944 ( po084 , new_n10247 , new_n10320 );
  xor  g09945 ( po085 , new_n10102 , new_n10106 );
  nand g09946 ( new_n10323 , new_n9611 , new_n9612 );
  nand g09947 ( new_n10324 , new_n9516 , new_n9613 );
  nand g09948 ( new_n10325 , new_n10323 , new_n10324 );
  or   g09949 ( new_n10326 , new_n9506 , new_n9608 );
  nand g09950 ( new_n10327 , new_n9607 , new_n9609 );
  nand g09951 ( new_n10328 , new_n10326 , new_n10327 );
  xor  g09952 ( new_n10329 , new_n10325 , new_n10328 );
  nor  g09953 ( new_n10330 , new_n9423 , new_n9430 );
  nor  g09954 ( new_n10331 , new_n9402 , new_n9431 );
  nor  g09955 ( new_n10332 , new_n10330 , new_n10331 );
  nand g09956 ( new_n10333 , pi088 , pi210 );
  nand g09957 ( new_n10334 , pi111 , pi183 );
  nand g09958 ( new_n10335 , pi024 , pi105 );
  xor  g09959 ( new_n10336 , new_n10334 , new_n10335 );
  nand g09960 ( new_n10337 , pi191 , pi213 );
  nand g09961 ( new_n10338 , new_n9601 , new_n9633 );
  nand g09962 ( new_n10339 , new_n9634 , new_n9637 );
  nand g09963 ( new_n10340 , new_n10338 , new_n10339 );
  xor  g09964 ( new_n10341 , new_n10337 , new_n10340 );
  xor  g09965 ( new_n10342 , new_n10336 , new_n10341 );
  xor  g09966 ( new_n10343 , new_n10333 , new_n10342 );
  nand g09967 ( new_n10344 , new_n9414 , new_n9415 );
  nand g09968 ( new_n10345 , new_n9393 , new_n9416 );
  nand g09969 ( new_n10346 , new_n10344 , new_n10345 );
  nand g09970 ( new_n10347 , pi106 , pi133 );
  nand g09971 ( new_n10348 , new_n9407 , new_n9408 );
  nand g09972 ( new_n10349 , new_n9385 , new_n9409 );
  nand g09973 ( new_n10350 , new_n10348 , new_n10349 );
  xor  g09974 ( new_n10351 , new_n10347 , new_n10350 );
  xor  g09975 ( new_n10352 , new_n10346 , new_n10351 );
  xor  g09976 ( new_n10353 , new_n10343 , new_n10352 );
  nand g09977 ( new_n10354 , pi017 , pi168 );
  nand g09978 ( new_n10355 , new_n9417 , new_n9420 );
  nand g09979 ( new_n10356 , new_n9413 , new_n9421 );
  nand g09980 ( new_n10357 , new_n10355 , new_n10356 );
  xor  g09981 ( new_n10358 , new_n10354 , new_n10357 );
  or   g09982 ( new_n10359 , new_n9551 , new_n9594 );
  nand g09983 ( new_n10360 , new_n9591 , new_n9595 );
  nand g09984 ( new_n10361 , new_n10359 , new_n10360 );
  nor  g09985 ( new_n10362 , new_n9574 , new_n9596 );
  nor  g09986 ( new_n10363 , new_n9597 , new_n9600 );
  nor  g09987 ( new_n10364 , new_n10362 , new_n10363 );
  xor  g09988 ( new_n10365 , new_n10361 , new_n10364 );
  nand g09989 ( new_n10366 , pi157 , pi208 );
  nand g09990 ( new_n10367 , new_n9463 , new_n9464 );
  nand g09991 ( new_n10368 , new_n9440 , new_n9465 );
  nand g09992 ( new_n10369 , new_n10367 , new_n10368 );
  or   g09993 ( new_n10370 , new_n9441 , new_n9467 );
  not  g09994 ( new_n10371 , new_n9466 );
  nand g09995 ( new_n10372 , new_n10371 , new_n9468 );
  nand g09996 ( new_n10373 , new_n10370 , new_n10372 );
  xor  g09997 ( new_n10374 , new_n10369 , new_n10373 );
  xor  g09998 ( new_n10375 , new_n10366 , new_n10374 );
  xor  g09999 ( new_n10376 , new_n10365 , new_n10375 );
  nand g10000 ( new_n10377 , pi125 , pi204 );
  nand g10001 ( new_n10378 , new_n9470 , new_n9471 );
  nand g10002 ( new_n10379 , new_n9454 , new_n9472 );
  nand g10003 ( new_n10380 , new_n10378 , new_n10379 );
  nand g10004 ( new_n10381 , pi035 , pi040 );
  nand g10005 ( new_n10382 , pi139 , pi174 );
  xor  g10006 ( new_n10383 , new_n10381 , new_n10382 );
  xor  g10007 ( new_n10384 , new_n10380 , new_n10383 );
  xor  g10008 ( new_n10385 , new_n10377 , new_n10384 );
  nand g10009 ( new_n10386 , pi015 , pi176 );
  nand g10010 ( new_n10387 , new_n9473 , new_n9476 );
  nand g10011 ( new_n10388 , new_n9469 , new_n9477 );
  nand g10012 ( new_n10389 , new_n10387 , new_n10388 );
  xor  g10013 ( new_n10390 , new_n10386 , new_n10389 );
  xor  g10014 ( new_n10391 , new_n10385 , new_n10390 );
  xor  g10015 ( new_n10392 , new_n10376 , new_n10391 );
  nand g10016 ( new_n10393 , pi146 , pi222 );
  nand g10017 ( new_n10394 , pi152 , pi249 );
  nor  g10018 ( new_n10395 , new_n9478 , new_n9483 );
  nor  g10019 ( new_n10396 , new_n9482 , new_n10395 );
  xor  g10020 ( new_n10397 , new_n10394 , new_n10396 );
  xor  g10021 ( new_n10398 , new_n10393 , new_n10397 );
  xor  g10022 ( new_n10399 , new_n10392 , new_n10398 );
  xor  g10023 ( new_n10400 , new_n10358 , new_n10399 );
  or   g10024 ( new_n10401 , new_n9462 , new_n9484 );
  nand g10025 ( new_n10402 , new_n9485 , new_n9492 );
  nand g10026 ( new_n10403 , new_n10401 , new_n10402 );
  nand g10027 ( new_n10404 , pi064 , pi227 );
  nand g10028 ( new_n10405 , pi084 , pi100 );
  xor  g10029 ( new_n10406 , new_n10404 , new_n10405 );
  nand g10030 ( new_n10407 , pi081 , pi189 );
  xor  g10031 ( new_n10408 , new_n10406 , new_n10407 );
  nand g10032 ( new_n10409 , pi052 , pi187 );
  or   g10033 ( new_n10410 , new_n9386 , new_n9411 );
  not  g10034 ( new_n10411 , new_n9410 );
  nand g10035 ( new_n10412 , new_n10411 , new_n9412 );
  nand g10036 ( new_n10413 , new_n10410 , new_n10412 );
  xor  g10037 ( new_n10414 , new_n10409 , new_n10413 );
  nand g10038 ( new_n10415 , pi077 , pi233 );
  xor  g10039 ( new_n10416 , new_n10414 , new_n10415 );
  xor  g10040 ( new_n10417 , new_n10408 , new_n10416 );
  xor  g10041 ( new_n10418 , new_n10403 , new_n10417 );
  xor  g10042 ( new_n10419 , new_n10400 , new_n10418 );
  xor  g10043 ( new_n10420 , new_n10353 , new_n10419 );
  xor  g10044 ( new_n10421 , new_n10332 , new_n10420 );
  xor  g10045 ( new_n10422 , new_n10329 , new_n10421 );
  nand g10046 ( new_n10423 , new_n9603 , new_n9604 );
  nand g10047 ( new_n10424 , new_n9505 , new_n9605 );
  nand g10048 ( new_n10425 , new_n10423 , new_n10424 );
  or   g10049 ( new_n10426 , new_n9614 , new_n9617 );
  nand g10050 ( new_n10427 , new_n9610 , new_n9618 );
  nand g10051 ( new_n10428 , new_n10426 , new_n10427 );
  nand g10052 ( new_n10429 , pi021 , pi241 );
  nand g10053 ( new_n10430 , pi005 , pi161 );
  xor  g10054 ( new_n10431 , new_n10429 , new_n10430 );
  xor  g10055 ( new_n10432 , new_n10428 , new_n10431 );
  xor  g10056 ( new_n10433 , new_n10425 , new_n10432 );
  nand g10057 ( new_n10434 , new_n9394 , new_n9405 );
  nand g10058 ( new_n10435 , new_n9406 , new_n9422 );
  nand g10059 ( new_n10436 , new_n10434 , new_n10435 );
  nand g10060 ( new_n10437 , pi047 , pi252 );
  nand g10061 ( new_n10438 , new_n9575 , new_n9576 );
  nand g10062 ( new_n10439 , new_n9542 , new_n9577 );
  nand g10063 ( new_n10440 , new_n10438 , new_n10439 );
  nand g10064 ( new_n10441 , new_n9583 , new_n9584 );
  nand g10065 ( new_n10442 , new_n9550 , new_n9585 );
  nand g10066 ( new_n10443 , new_n10441 , new_n10442 );
  xor  g10067 ( new_n10444 , new_n10440 , new_n10443 );
  nand g10068 ( new_n10445 , pi112 , pi224 );
  xor  g10069 ( new_n10446 , new_n10444 , new_n10445 );
  or   g10070 ( new_n10447 , new_n9543 , new_n9580 );
  nand g10071 ( new_n10448 , new_n9579 , new_n9581 );
  nand g10072 ( new_n10449 , new_n10447 , new_n10448 );
  nand g10073 ( new_n10450 , pi212 , pi232 );
  nand g10074 ( new_n10451 , pi104 , pi127 );
  xor  g10075 ( new_n10452 , new_n10450 , new_n10451 );
  nand g10076 ( new_n10453 , pi013 , pi255 );
  nand g10077 ( new_n10454 , new_n9586 , new_n9589 );
  not  g10078 ( new_n10455 , new_n9582 );
  nand g10079 ( new_n10456 , new_n10455 , new_n9590 );
  nand g10080 ( new_n10457 , new_n10454 , new_n10456 );
  xnor g10081 ( new_n10458 , new_n10453 , new_n10457 );
  xor  g10082 ( new_n10459 , new_n10452 , new_n10458 );
  xor  g10083 ( new_n10460 , new_n10449 , new_n10459 );
  xor  g10084 ( new_n10461 , new_n10446 , new_n10460 );
  xor  g10085 ( new_n10462 , new_n10437 , new_n10461 );
  xor  g10086 ( new_n10463 , new_n10436 , new_n10462 );
  nand g10087 ( new_n10464 , new_n9432 , new_n9639 );
  nand g10088 ( new_n10465 , new_n9640 , new_n9649 );
  nand g10089 ( new_n10466 , new_n10464 , new_n10465 );
  nand g10090 ( new_n10467 , pi018 , pi140 );
  nand g10091 ( new_n10468 , pi128 , pi242 );
  xor  g10092 ( new_n10469 , new_n10467 , new_n10468 );
  or   g10093 ( new_n10470 , new_n9602 , new_n9626 );
  nand g10094 ( new_n10471 , new_n9627 , new_n9631 );
  nand g10095 ( new_n10472 , new_n10470 , new_n10471 );
  nand g10096 ( new_n10473 , pi082 , pi236 );
  xor  g10097 ( new_n10474 , new_n10472 , new_n10473 );
  xor  g10098 ( new_n10475 , new_n10469 , new_n10474 );
  or   g10099 ( new_n10476 , new_n9619 , new_n9625 );
  nand g10100 ( new_n10477 , new_n9624 , new_n10476 );
  nand g10101 ( new_n10478 , pi090 , pi121 );
  nand g10102 ( new_n10479 , pi141 , pi231 );
  xor  g10103 ( new_n10480 , new_n10478 , new_n10479 );
  xor  g10104 ( new_n10481 , new_n10477 , new_n10480 );
  xor  g10105 ( new_n10482 , new_n10475 , new_n10481 );
  xor  g10106 ( new_n10483 , new_n10466 , new_n10482 );
  xor  g10107 ( new_n10484 , new_n10463 , new_n10483 );
  nor  g10108 ( new_n10485 , new_n9493 , new_n9570 );
  nor  g10109 ( new_n10486 , new_n9572 , new_n9638 );
  or   g10110 ( new_n10487 , new_n10485 , new_n10486 );
  nand g10111 ( new_n10488 , pi034 , pi217 );
  nand g10112 ( new_n10489 , pi129 , pi131 );
  xor  g10113 ( new_n10490 , new_n10488 , new_n10489 );
  xor  g10114 ( new_n10491 , new_n10487 , new_n10490 );
  xor  g10115 ( new_n10492 , new_n10484 , new_n10491 );
  xor  g10116 ( new_n10493 , new_n10433 , new_n10492 );
  xor  g10117 ( po086 , new_n10422 , new_n10493 );
  xnor g10118 ( po087 , new_n7521 , new_n7522 );
  xnor g10119 ( po088 , new_n4803 , new_n4804 );
  xor  g10120 ( po089 , new_n3067 , new_n3088 );
  xor  g10121 ( po090 , new_n2561 , new_n2562 );
  xor  g10122 ( po091 , new_n3499 , new_n3501 );
  xnor g10123 ( po092 , new_n5667 , new_n5677 );
  xor  g10124 ( po093 , new_n9160 , new_n9189 );
  xor  g10125 ( po094 , new_n899 , new_n901 );
  xor  g10126 ( po095 , new_n1049 , new_n1050 );
  xor  g10127 ( po096 , new_n3505 , new_n3506 );
  nand g10128 ( new_n10505 , pi213 , pi243 );
  or   g10129 ( new_n10506 , new_n5119 , new_n5142 );
  nand g10130 ( new_n10507 , new_n5143 , new_n5152 );
  nand g10131 ( new_n10508 , new_n10506 , new_n10507 );
  nor  g10132 ( new_n10509 , new_n5135 , new_n5141 );
  nor  g10133 ( new_n10510 , new_n5140 , new_n10509 );
  xor  g10134 ( new_n10511 , new_n10508 , new_n10510 );
  xor  g10135 ( new_n10512 , new_n10505 , new_n10511 );
  nand g10136 ( new_n10513 , pi183 , pi207 );
  nand g10137 ( new_n10514 , pi066 , pi105 );
  xor  g10138 ( new_n10515 , new_n10513 , new_n10514 );
  nand g10139 ( new_n10516 , pi088 , pi226 );
  xor  g10140 ( new_n10517 , new_n10515 , new_n10516 );
  nand g10141 ( new_n10518 , new_n5223 , new_n5224 );
  nand g10142 ( new_n10519 , new_n5193 , new_n5225 );
  nand g10143 ( new_n10520 , new_n10518 , new_n10519 );
  not  g10144 ( new_n10521 , new_n5153 );
  nand g10145 ( new_n10522 , new_n5074 , new_n10521 );
  or   g10146 ( new_n10523 , new_n5154 , new_n5171 );
  nand g10147 ( new_n10524 , new_n10522 , new_n10523 );
  xor  g10148 ( new_n10525 , new_n10520 , new_n10524 );
  xor  g10149 ( new_n10526 , new_n10517 , new_n10525 );
  xor  g10150 ( new_n10527 , new_n10512 , new_n10526 );
  nand g10151 ( new_n10528 , pi208 , pi218 );
  nand g10152 ( new_n10529 , new_n5216 , new_n5217 );
  nand g10153 ( new_n10530 , new_n5178 , new_n5218 );
  nand g10154 ( new_n10531 , new_n10529 , new_n10530 );
  or   g10155 ( new_n10532 , new_n5179 , new_n5220 );
  not  g10156 ( new_n10533 , new_n5219 );
  nand g10157 ( new_n10534 , new_n10533 , new_n5221 );
  nand g10158 ( new_n10535 , new_n10532 , new_n10534 );
  xor  g10159 ( new_n10536 , new_n10531 , new_n10535 );
  xor  g10160 ( new_n10537 , new_n10528 , new_n10536 );
  xor  g10161 ( new_n10538 , new_n10527 , new_n10537 );
  nand g10162 ( new_n10539 , pi058 , pi204 );
  or   g10163 ( new_n10540 , new_n5275 , new_n5316 );
  not  g10164 ( new_n10541 , new_n5315 );
  nand g10165 ( new_n10542 , new_n10541 , new_n5317 );
  nand g10166 ( new_n10543 , new_n10540 , new_n10542 );
  nand g10167 ( new_n10544 , pi035 , pi199 );
  nand g10168 ( new_n10545 , pi139 , pi195 );
  xor  g10169 ( new_n10546 , new_n10544 , new_n10545 );
  xor  g10170 ( new_n10547 , new_n10543 , new_n10546 );
  xor  g10171 ( new_n10548 , new_n10539 , new_n10547 );
  nand g10172 ( new_n10549 , pi015 , pi211 );
  nand g10173 ( new_n10550 , new_n5226 , new_n5229 );
  nand g10174 ( new_n10551 , new_n5222 , new_n5230 );
  nand g10175 ( new_n10552 , new_n10550 , new_n10551 );
  xor  g10176 ( new_n10553 , new_n10549 , new_n10552 );
  xor  g10177 ( new_n10554 , new_n10548 , new_n10553 );
  xor  g10178 ( new_n10555 , new_n10538 , new_n10554 );
  nand g10179 ( new_n10556 , new_n5043 , new_n5044 );
  nand g10180 ( new_n10557 , new_n5005 , new_n5045 );
  nand g10181 ( new_n10558 , new_n10556 , new_n10557 );
  nand g10182 ( new_n10559 , new_n5050 , new_n5051 );
  nand g10183 ( new_n10560 , new_n5020 , new_n5052 );
  nand g10184 ( new_n10561 , new_n10559 , new_n10560 );
  xor  g10185 ( new_n10562 , new_n10558 , new_n10561 );
  or   g10186 ( new_n10563 , new_n5006 , new_n5047 );
  not  g10187 ( new_n10564 , new_n5046 );
  nand g10188 ( new_n10565 , new_n10564 , new_n5048 );
  nand g10189 ( new_n10566 , new_n10563 , new_n10565 );
  xor  g10190 ( new_n10567 , new_n10562 , new_n10566 );
  xor  g10191 ( new_n10568 , new_n10555 , new_n10567 );
  nand g10192 ( new_n10569 , new_n5290 , new_n5329 );
  nand g10193 ( new_n10570 , new_n5327 , new_n5332 );
  nand g10194 ( new_n10571 , new_n10569 , new_n10570 );
  not  g10195 ( new_n10572 , new_n5333 );
  nor  g10196 ( new_n10573 , new_n5311 , new_n10572 );
  nor  g10197 ( new_n10574 , new_n5334 , new_n5345 );
  nor  g10198 ( new_n10575 , new_n10573 , new_n10574 );
  xor  g10199 ( new_n10576 , new_n10571 , new_n10575 );
  nand g10200 ( new_n10577 , pi029 , pi034 );
  nand g10201 ( new_n10578 , pi010 , pi131 );
  xor  g10202 ( new_n10579 , new_n10577 , new_n10578 );
  nand g10203 ( new_n10580 , new_n5053 , new_n5056 );
  nand g10204 ( new_n10581 , new_n5049 , new_n5057 );
  nand g10205 ( new_n10582 , new_n10580 , new_n10581 );
  nand g10206 ( new_n10583 , pi074 , pi241 );
  nand g10207 ( new_n10584 , pi161 , pi253 );
  xor  g10208 ( new_n10585 , new_n10583 , new_n10584 );
  xor  g10209 ( new_n10586 , new_n10582 , new_n10585 );
  xor  g10210 ( new_n10587 , new_n10579 , new_n10586 );
  xor  g10211 ( new_n10588 , new_n10576 , new_n10587 );
  xor  g10212 ( new_n10589 , new_n10568 , new_n10588 );
  nand g10213 ( new_n10590 , pi069 , pi084 );
  nand g10214 ( new_n10591 , new_n5312 , new_n5313 );
  nand g10215 ( new_n10592 , new_n5274 , new_n5314 );
  nand g10216 ( new_n10593 , new_n10591 , new_n10592 );
  xor  g10217 ( new_n10594 , new_n10590 , new_n10593 );
  xor  g10218 ( new_n10595 , new_n10589 , new_n10594 );
  nand g10219 ( new_n10596 , new_n5236 , new_n5245 );
  nand g10220 ( new_n10597 , new_n5215 , new_n5246 );
  nand g10221 ( new_n10598 , new_n10596 , new_n10597 );
  nand g10222 ( new_n10599 , pi150 , pi189 );
  nand g10223 ( new_n10600 , pi133 , pi221 );
  xor  g10224 ( new_n10601 , new_n10599 , new_n10600 );
  xor  g10225 ( new_n10602 , new_n10598 , new_n10601 );
  not  g10226 ( new_n10603 , new_n5247 );
  nor  g10227 ( new_n10604 , new_n5172 , new_n10603 );
  nor  g10228 ( new_n10605 , new_n5248 , new_n5267 );
  nor  g10229 ( new_n10606 , new_n10604 , new_n10605 );
  nand g10230 ( new_n10607 , pi064 , pi244 );
  xor  g10231 ( new_n10608 , new_n10606 , new_n10607 );
  xor  g10232 ( new_n10609 , new_n10602 , new_n10608 );
  nand g10233 ( new_n10610 , pi052 , pi184 );
  nand g10234 ( new_n10611 , pi077 , pi196 );
  xor  g10235 ( new_n10612 , new_n10610 , new_n10611 );
  nand g10236 ( new_n10613 , new_n5322 , new_n5325 );
  nand g10237 ( new_n10614 , new_n5318 , new_n5326 );
  nand g10238 ( new_n10615 , new_n10613 , new_n10614 );
  nand g10239 ( new_n10616 , pi146 , pi186 );
  nand g10240 ( new_n10617 , pi037 , pi168 );
  xor  g10241 ( new_n10618 , new_n10616 , new_n10617 );
  xor  g10242 ( new_n10619 , new_n10615 , new_n10618 );
  nand g10243 ( new_n10620 , pi132 , pi152 );
  nand g10244 ( new_n10621 , new_n5194 , new_n5233 );
  not  g10245 ( new_n10622 , new_n5235 );
  nand g10246 ( new_n10623 , new_n5231 , new_n10622 );
  nand g10247 ( new_n10624 , new_n10621 , new_n10623 );
  xor  g10248 ( new_n10625 , new_n10620 , new_n10624 );
  nand g10249 ( new_n10626 , new_n5319 , new_n5320 );
  nand g10250 ( new_n10627 , new_n5289 , new_n5321 );
  nand g10251 ( new_n10628 , new_n10626 , new_n10627 );
  xor  g10252 ( new_n10629 , new_n10625 , new_n10628 );
  xor  g10253 ( new_n10630 , new_n10619 , new_n10629 );
  xor  g10254 ( new_n10631 , new_n10612 , new_n10630 );
  xor  g10255 ( new_n10632 , new_n10609 , new_n10631 );
  xor  g10256 ( new_n10633 , new_n10595 , new_n10632 );
  nand g10257 ( new_n10634 , new_n5021 , new_n5060 );
  not  g10258 ( new_n10635 , new_n5062 );
  nand g10259 ( new_n10636 , new_n5058 , new_n10635 );
  nand g10260 ( new_n10637 , new_n10634 , new_n10636 );
  nand g10261 ( new_n10638 , pi047 , pi173 );
  nand g10262 ( new_n10639 , pi014 , pi018 );
  xor  g10263 ( new_n10640 , new_n10638 , new_n10639 );
  xor  g10264 ( new_n10641 , new_n10637 , new_n10640 );
  xor  g10265 ( new_n10642 , new_n10633 , new_n10641 );
  nand g10266 ( new_n10643 , pi090 , pi230 );
  nand g10267 ( new_n10644 , pi050 , pi141 );
  xor  g10268 ( new_n10645 , new_n10643 , new_n10644 );
  nand g10269 ( new_n10646 , new_n5130 , new_n5133 );
  nand g10270 ( new_n10647 , new_n5126 , new_n5134 );
  nand g10271 ( new_n10648 , new_n10646 , new_n10647 );
  nand g10272 ( new_n10649 , new_n5127 , new_n5128 );
  nand g10273 ( new_n10650 , new_n5095 , new_n5129 );
  nand g10274 ( new_n10651 , new_n10649 , new_n10650 );
  xor  g10275 ( new_n10652 , new_n10648 , new_n10651 );
  nand g10276 ( new_n10653 , pi055 , pi112 );
  or   g10277 ( new_n10654 , new_n5087 , new_n5124 );
  not  g10278 ( new_n10655 , new_n5123 );
  nand g10279 ( new_n10656 , new_n10655 , new_n5125 );
  nand g10280 ( new_n10657 , new_n10654 , new_n10656 );
  nand g10281 ( new_n10658 , pi212 , pi239 );
  nand g10282 ( new_n10659 , pi025 , pi104 );
  xor  g10283 ( new_n10660 , new_n10658 , new_n10659 );
  xor  g10284 ( new_n10661 , new_n10657 , new_n10660 );
  xor  g10285 ( new_n10662 , new_n10653 , new_n10661 );
  nand g10286 ( new_n10663 , pi002 , pi013 );
  nand g10287 ( new_n10664 , new_n5120 , new_n5121 );
  nand g10288 ( new_n10665 , new_n5086 , new_n5122 );
  nand g10289 ( new_n10666 , new_n10664 , new_n10665 );
  xor  g10290 ( new_n10667 , new_n10663 , new_n10666 );
  xor  g10291 ( new_n10668 , new_n10662 , new_n10667 );
  xor  g10292 ( new_n10669 , new_n10652 , new_n10668 );
  xor  g10293 ( new_n10670 , new_n10645 , new_n10669 );
  nor  g10294 ( new_n10671 , new_n5268 , new_n5346 );
  not  g10295 ( new_n10672 , new_n5347 );
  nor  g10296 ( new_n10673 , new_n10672 , new_n5363 );
  nor  g10297 ( new_n10674 , new_n10671 , new_n10673 );
  nand g10298 ( new_n10675 , pi205 , pi236 );
  xor  g10299 ( new_n10676 , new_n10674 , new_n10675 );
  xor  g10300 ( new_n10677 , new_n10670 , new_n10676 );
  nor  g10301 ( new_n10678 , new_n5042 , new_n5063 );
  nor  g10302 ( new_n10679 , new_n5064 , new_n5073 );
  nor  g10303 ( new_n10680 , new_n10678 , new_n10679 );
  nand g10304 ( new_n10681 , pi109 , pi128 );
  xor  g10305 ( new_n10682 , new_n10680 , new_n10681 );
  xor  g10306 ( new_n10683 , new_n10677 , new_n10682 );
  xor  g10307 ( po097 , new_n10642 , new_n10683 );
  xor  g10308 ( po098 , new_n1801 , new_n1803 );
  xnor g10309 ( po099 , new_n7740 , new_n7741 );
  xnor g10310 ( po100 , new_n889 , new_n890 );
  xor  g10311 ( po101 , new_n885 , new_n887 );
  xor  g10312 ( po102 , new_n1043 , new_n1045 );
  xor  g10313 ( po103 , new_n3115 , new_n3116 );
  xor  g10314 ( po104 , new_n1986 , new_n2554 );
  xnor g10315 ( po105 , new_n3694 , new_n3695 );
  xor  g10316 ( po106 , new_n5762 , new_n5764 );
  xor  g10317 ( po107 , new_n9191 , new_n9192 );
  xor  g10318 ( po108 , new_n3607 , new_n3683 );
  or   g10319 ( new_n10696 , new_n4496 , new_n4530 );
  not  g10320 ( new_n10697 , new_n4529 );
  nand g10321 ( new_n10698 , new_n10697 , new_n4531 );
  nand g10322 ( new_n10699 , new_n10696 , new_n10698 );
  nand g10323 ( new_n10700 , pi046 , pi103 );
  nor  g10324 ( new_n10701 , new_n4525 , new_n4546 );
  not  g10325 ( new_n10702 , new_n4547 );
  nor  g10326 ( new_n10703 , new_n10702 , new_n4556 );
  nor  g10327 ( new_n10704 , new_n10701 , new_n10703 );
  xor  g10328 ( new_n10705 , new_n10700 , new_n10704 );
  xor  g10329 ( new_n10706 , new_n10699 , new_n10705 );
  nand g10330 ( new_n10707 , pi000 , pi188 );
  nand g10331 ( new_n10708 , pi115 , pi178 );
  nand g10332 ( new_n10709 , pi061 , pi070 );
  xor  g10333 ( new_n10710 , new_n10708 , new_n10709 );
  nand g10334 ( new_n10711 , new_n4438 , new_n4439 );
  nand g10335 ( new_n10712 , new_n4407 , new_n4440 );
  nand g10336 ( new_n10713 , new_n10711 , new_n10712 );
  nand g10337 ( new_n10714 , pi048 , pi167 );
  or   g10338 ( new_n10715 , new_n4400 , new_n4435 );
  not  g10339 ( new_n10716 , new_n4434 );
  nand g10340 ( new_n10717 , new_n10716 , new_n4436 );
  nand g10341 ( new_n10718 , new_n10715 , new_n10717 );
  xor  g10342 ( new_n10719 , new_n10714 , new_n10718 );
  xor  g10343 ( new_n10720 , new_n10713 , new_n10719 );
  nand g10344 ( new_n10721 , new_n4313 , new_n4353 );
  nand g10345 ( new_n10722 , new_n4351 , new_n4356 );
  nand g10346 ( new_n10723 , new_n10721 , new_n10722 );
  nand g10347 ( new_n10724 , pi149 , pi237 );
  nand g10348 ( new_n10725 , pi238 , pi240 );
  xor  g10349 ( new_n10726 , new_n10724 , new_n10725 );
  nand g10350 ( new_n10727 , pi179 , pi181 );
  xor  g10351 ( new_n10728 , new_n10726 , new_n10727 );
  nand g10352 ( new_n10729 , pi134 , pi193 );
  nand g10353 ( new_n10730 , new_n4441 , new_n4444 );
  nand g10354 ( new_n10731 , new_n4437 , new_n4445 );
  nand g10355 ( new_n10732 , new_n10730 , new_n10731 );
  xor  g10356 ( new_n10733 , new_n10729 , new_n10732 );
  nand g10357 ( new_n10734 , new_n4431 , new_n4432 );
  nand g10358 ( new_n10735 , new_n4399 , new_n4433 );
  nand g10359 ( new_n10736 , new_n10734 , new_n10735 );
  xor  g10360 ( new_n10737 , new_n10733 , new_n10736 );
  xor  g10361 ( new_n10738 , new_n10728 , new_n10737 );
  xor  g10362 ( new_n10739 , new_n10723 , new_n10738 );
  xor  g10363 ( new_n10740 , new_n10720 , new_n10739 );
  xor  g10364 ( new_n10741 , new_n10710 , new_n10740 );
  xor  g10365 ( new_n10742 , new_n10707 , new_n10741 );
  not  g10366 ( new_n10743 , new_n4452 );
  nor  g10367 ( new_n10744 , new_n4430 , new_n10743 );
  nor  g10368 ( new_n10745 , new_n4453 , new_n4463 );
  nor  g10369 ( new_n10746 , new_n10744 , new_n10745 );
  nand g10370 ( new_n10747 , new_n4526 , new_n4527 );
  nand g10371 ( new_n10748 , new_n4495 , new_n4528 );
  nand g10372 ( new_n10749 , new_n10747 , new_n10748 );
  nand g10373 ( new_n10750 , new_n4536 , new_n4539 );
  nand g10374 ( new_n10751 , new_n4532 , new_n4540 );
  nand g10375 ( new_n10752 , new_n10750 , new_n10751 );
  xor  g10376 ( new_n10753 , new_n10749 , new_n10752 );
  nand g10377 ( new_n10754 , pi068 , pi117 );
  nand g10378 ( new_n10755 , pi016 , pi036 );
  xor  g10379 ( new_n10756 , new_n10754 , new_n10755 );
  nand g10380 ( new_n10757 , pi057 , pi214 );
  xor  g10381 ( new_n10758 , new_n10756 , new_n10757 );
  xor  g10382 ( new_n10759 , new_n10753 , new_n10758 );
  xor  g10383 ( new_n10760 , new_n10746 , new_n10759 );
  xor  g10384 ( new_n10761 , new_n10742 , new_n10760 );
  nand g10385 ( new_n10762 , new_n4386 , new_n4464 );
  nand g10386 ( new_n10763 , new_n4465 , new_n4481 );
  nand g10387 ( new_n10764 , new_n10762 , new_n10763 );
  nand g10388 ( new_n10765 , pi126 , pi163 );
  not  g10389 ( new_n10766 , new_n4357 );
  nor  g10390 ( new_n10767 , new_n4335 , new_n10766 );
  nor  g10391 ( new_n10768 , new_n4358 , new_n4367 );
  or   g10392 ( new_n10769 , new_n10767 , new_n10768 );
  xor  g10393 ( new_n10770 , new_n10765 , new_n10769 );
  nand g10394 ( new_n10771 , new_n4291 , new_n4369 );
  nand g10395 ( new_n10772 , new_n4370 , new_n4385 );
  nand g10396 ( new_n10773 , new_n10771 , new_n10772 );
  nand g10397 ( new_n10774 , pi162 , pi203 );
  nand g10398 ( new_n10775 , new_n4408 , new_n4448 );
  nand g10399 ( new_n10776 , new_n4446 , new_n4451 );
  nand g10400 ( new_n10777 , new_n10775 , new_n10776 );
  xor  g10401 ( new_n10778 , new_n10774 , new_n10777 );
  nand g10402 ( new_n10779 , pi033 , pi200 );
  nand g10403 ( new_n10780 , pi159 , pi175 );
  xor  g10404 ( new_n10781 , new_n10779 , new_n10780 );
  nand g10405 ( new_n10782 , new_n4533 , new_n4534 );
  nand g10406 ( new_n10783 , new_n4503 , new_n4535 );
  nand g10407 ( new_n10784 , new_n10782 , new_n10783 );
  xor  g10408 ( new_n10785 , new_n10781 , new_n10784 );
  xor  g10409 ( new_n10786 , new_n10778 , new_n10785 );
  nand g10410 ( new_n10787 , pi194 , pi234 );
  nand g10411 ( new_n10788 , pi085 , pi247 );
  nand g10412 ( new_n10789 , pi080 , pi180 );
  xor  g10413 ( new_n10790 , new_n10788 , new_n10789 );
  xor  g10414 ( new_n10791 , new_n10787 , new_n10790 );
  xor  g10415 ( new_n10792 , new_n10786 , new_n10791 );
  xor  g10416 ( new_n10793 , new_n10773 , new_n10792 );
  xor  g10417 ( new_n10794 , new_n10770 , new_n10793 );
  xor  g10418 ( new_n10795 , new_n10764 , new_n10794 );
  xor  g10419 ( new_n10796 , new_n10761 , new_n10795 );
  nand g10420 ( new_n10797 , new_n4343 , new_n4344 );
  nand g10421 ( new_n10798 , new_n4312 , new_n4345 );
  nand g10422 ( new_n10799 , new_n10797 , new_n10798 );
  or   g10423 ( new_n10800 , new_n4298 , new_n4340 );
  not  g10424 ( new_n10801 , new_n4339 );
  nand g10425 ( new_n10802 , new_n10801 , new_n4341 );
  nand g10426 ( new_n10803 , new_n10800 , new_n10802 );
  xor  g10427 ( new_n10804 , new_n10799 , new_n10803 );
  nand g10428 ( new_n10805 , new_n4336 , new_n4337 );
  nand g10429 ( new_n10806 , new_n4297 , new_n4338 );
  nand g10430 ( new_n10807 , new_n10805 , new_n10806 );
  nand g10431 ( new_n10808 , pi012 , pi116 );
  xor  g10432 ( new_n10809 , new_n10807 , new_n10808 );
  xor  g10433 ( new_n10810 , new_n10804 , new_n10809 );
  nand g10434 ( new_n10811 , new_n4504 , new_n4543 );
  not  g10435 ( new_n10812 , new_n4545 );
  nand g10436 ( new_n10813 , new_n4541 , new_n10812 );
  nand g10437 ( new_n10814 , new_n10811 , new_n10813 );
  nand g10438 ( new_n10815 , pi108 , pi156 );
  nand g10439 ( new_n10816 , pi051 , pi083 );
  nand g10440 ( new_n10817 , pi028 , pi107 );
  xor  g10441 ( new_n10818 , new_n10816 , new_n10817 );
  xor  g10442 ( new_n10819 , new_n10815 , new_n10818 );
  nand g10443 ( new_n10820 , pi007 , pi201 );
  nand g10444 ( new_n10821 , pi118 , pi245 );
  xor  g10445 ( new_n10822 , new_n10820 , new_n10821 );
  nand g10446 ( new_n10823 , pi042 , pi063 );
  xor  g10447 ( new_n10824 , new_n10822 , new_n10823 );
  nand g10448 ( new_n10825 , new_n4252 , new_n4286 );
  not  g10449 ( new_n10826 , new_n4288 );
  nand g10450 ( new_n10827 , new_n4284 , new_n10826 );
  nand g10451 ( new_n10828 , new_n10825 , new_n10827 );
  nand g10452 ( new_n10829 , new_n4267 , new_n4289 );
  nand g10453 ( new_n10830 , new_n4266 , new_n4290 );
  nand g10454 ( new_n10831 , new_n10829 , new_n10830 );
  xor  g10455 ( new_n10832 , new_n10828 , new_n10831 );
  xor  g10456 ( new_n10833 , new_n10824 , new_n10832 );
  xor  g10457 ( new_n10834 , new_n10819 , new_n10833 );
  nand g10458 ( new_n10835 , pi043 , pi148 );
  nand g10459 ( new_n10836 , pi098 , pi228 );
  xor  g10460 ( new_n10837 , new_n10835 , new_n10836 );
  nand g10461 ( new_n10838 , pi039 , pi144 );
  nand g10462 ( new_n10839 , new_n4346 , new_n4349 );
  nand g10463 ( new_n10840 , new_n4342 , new_n4350 );
  nand g10464 ( new_n10841 , new_n10839 , new_n10840 );
  xor  g10465 ( new_n10842 , new_n10838 , new_n10841 );
  xor  g10466 ( new_n10843 , new_n10837 , new_n10842 );
  xor  g10467 ( new_n10844 , new_n10834 , new_n10843 );
  xor  g10468 ( new_n10845 , new_n10814 , new_n10844 );
  xor  g10469 ( new_n10846 , new_n10810 , new_n10845 );
  nand g10470 ( new_n10847 , pi143 , pi202 );
  nand g10471 ( new_n10848 , new_n4557 , new_n4574 );
  not  g10472 ( new_n10849 , new_n4482 );
  nand g10473 ( new_n10850 , new_n10849 , new_n4575 );
  nand g10474 ( new_n10851 , new_n10848 , new_n10850 );
  nand g10475 ( new_n10852 , pi038 , pi171 );
  nand g10476 ( new_n10853 , pi049 , pi113 );
  xor  g10477 ( new_n10854 , new_n10852 , new_n10853 );
  xor  g10478 ( new_n10855 , new_n10851 , new_n10854 );
  or   g10479 ( new_n10856 , new_n4241 , new_n4273 );
  nand g10480 ( new_n10857 , new_n4272 , new_n4274 );
  nand g10481 ( new_n10858 , new_n10856 , new_n10857 );
  or   g10482 ( new_n10859 , new_n4279 , new_n4282 );
  nand g10483 ( new_n10860 , new_n4275 , new_n4283 );
  nand g10484 ( new_n10861 , new_n10859 , new_n10860 );
  nand g10485 ( new_n10862 , new_n4268 , new_n4269 );
  nand g10486 ( new_n10863 , new_n4240 , new_n4270 );
  nand g10487 ( new_n10864 , new_n10862 , new_n10863 );
  nand g10488 ( new_n10865 , new_n4276 , new_n4277 );
  nand g10489 ( new_n10866 , new_n4251 , new_n4278 );
  nand g10490 ( new_n10867 , new_n10865 , new_n10866 );
  xor  g10491 ( new_n10868 , new_n10864 , new_n10867 );
  xor  g10492 ( new_n10869 , new_n10861 , new_n10868 );
  xor  g10493 ( new_n10870 , new_n10858 , new_n10869 );
  xor  g10494 ( new_n10871 , new_n10855 , new_n10870 );
  xor  g10495 ( new_n10872 , new_n10847 , new_n10871 );
  xor  g10496 ( new_n10873 , new_n10846 , new_n10872 );
  xor  g10497 ( new_n10874 , new_n10796 , new_n10873 );
  xor  g10498 ( po109 , new_n10706 , new_n10874 );
  xor  g10499 ( po110 , new_n4948 , new_n4949 );
  xor  g10500 ( po111 , new_n3107 , new_n3108 );
  xor  g10501 ( po112 , new_n8105 , new_n8106 );
  xor  g10502 ( po113 , new_n8110 , new_n8112 );
  xor  g10503 ( po114 , new_n8421 , new_n8423 );
  xor  g10504 ( po115 , new_n7055 , new_n7057 );
  xor  g10505 ( po116 , new_n9186 , new_n9187 );
  xor  g10506 ( po117 , new_n9646 , new_n9647 );
  xor  g10507 ( po118 , new_n8414 , new_n8425 );
  xor  g10508 ( po119 , new_n4570 , new_n4572 );
endmodule


