// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Fri Aug 16 22:57:15 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604,
    n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112,
    n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288,
    n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558,
    n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738,
    n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088,
    n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272,
    n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479,
    n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816,
    n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136,
    n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349,
    n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618,
    n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952,
    n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319,
    n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722,
    n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031,
    n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213,
    n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443,
    n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822,
    n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379,
    n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590,
    n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790,
    n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305,
    n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566,
    n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731,
    n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963,
    n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305,
    n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614,
    n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827,
    n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251,
    n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493,
    n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926,
    n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117,
    n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514,
    n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763,
    n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220,
    n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479,
    n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667,
    n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121,
    n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398,
    n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650,
    n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900,
    n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263,
    n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494,
    n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783,
    n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230,
    n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603,
    n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899,
    n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271,
    n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546,
    n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918,
    n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247,
    n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524,
    n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968,
    n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095,
    n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954,
    n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227,
    n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496,
    n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880,
    n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107,
    n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327,
    n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531,
    n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770,
    n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040,
    n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259,
    n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478,
    n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946,
    n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287,
    n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674,
    n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898,
    n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068,
    n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309,
    n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492,
    n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764,
    n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068,
    n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333,
    n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657,
    n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912,
    n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129,
    n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485,
    n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023,
    n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240,
    n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435,
    n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643,
    n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926,
    n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191,
    n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512,
    n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752,
    n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089,
    n27104, n27120, n27134, n27188,
    n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194  );
  input  n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583,
    n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099,
    n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279,
    n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536,
    n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689,
    n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035,
    n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210,
    n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421,
    n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809,
    n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030,
    n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324,
    n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582,
    n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945,
    n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306,
    n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665,
    n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026,
    n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211,
    n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438,
    n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752,
    n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369,
    n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556,
    n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785,
    n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149,
    n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524,
    n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721,
    n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949,
    n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285,
    n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581,
    n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806,
    n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246,
    n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460,
    n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872,
    n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096,
    n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411,
    n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739,
    n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201,
    n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473,
    n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630,
    n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113,
    n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384,
    n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626,
    n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892,
    n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190,
    n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490,
    n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781,
    n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148,
    n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576,
    n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826,
    n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258,
    n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539,
    n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884,
    n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223,
    n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521,
    n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911,
    n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090,
    n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911,
    n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171,
    n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483,
    n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745,
    n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081,
    n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282,
    n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515,
    n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701,
    n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036,
    n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250,
    n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470,
    n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929,
    n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276,
    n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654,
    n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839,
    n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043,
    n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290,
    n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470,
    n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660,
    n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065,
    n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304,
    n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586,
    n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895,
    n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093,
    n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374,
    n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937,
    n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168,
    n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381,
    n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629,
    n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923,
    n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180,
    n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510,
    n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748,
    n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037,
    n27089, n27104, n27120, n27134, n27188;
  output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355_1, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361_1, new_n2362, new_n2363_1, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374_1, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387_1, new_n2388_1, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409_1, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416_1, new_n2417, new_n2418, new_n2419, new_n2420_1,
    new_n2421_1, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440_1, new_n2441, new_n2442, new_n2443, new_n2444_1,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479_1, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513_1, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533_1, new_n2534,
    new_n2535_1, new_n2536, new_n2537_1, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547_1, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552,
    new_n2553_1, new_n2554, new_n2555_1, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560_1, new_n2561_1, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570_1,
    new_n2571, new_n2572, new_n2573_1, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578_1, new_n2579, new_n2580, new_n2581, new_n2582_1,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602_1, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619_1,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2646_1, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659_1, new_n2660, new_n2661_1, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680_1, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693_1,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703_1, new_n2704, new_n2705,
    new_n2706_1, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711_1,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731_1, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743_1, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761_1, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774_1, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779_1, new_n2780, new_n2781, new_n2782, new_n2783_1,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809_1, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816_1, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826_1, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853_1, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858_1, new_n2859, new_n2860_1, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886_1, new_n2887_1, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929_1, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944_1, new_n2945,
    new_n2946, new_n2947, new_n2948_1, new_n2949, new_n2950, new_n2951,
    new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961_1, new_n2962, new_n2963,
    new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969,
    new_n2970, new_n2971_1, new_n2972, new_n2973, new_n2974, new_n2975,
    new_n2976, new_n2977, new_n2978_1, new_n2979_1, new_n2980, new_n2981,
    new_n2982, new_n2983, new_n2984, new_n2985_1, new_n2986, new_n2987,
    new_n2988, new_n2989, new_n2990, new_n2991, new_n2992, new_n2993,
    new_n2994, new_n2996, new_n2997, new_n2998, new_n2999_1, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010_1, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017_1, new_n3018_1,
    new_n3019, new_n3020_1, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030_1,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067_1, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076_1, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089_1, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125_1, new_n3126_1,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136_1, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161_1, new_n3162,
    new_n3163, new_n3164_1, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208_1, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219_1, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228_1,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235_1, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244_1, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253_1, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260_1, new_n3261, new_n3262, new_n3263_1, new_n3264,
    new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279_1, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289_1, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301_1, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306_1,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3313,
    new_n3314, new_n3315, new_n3316_1, new_n3317, new_n3318, new_n3319,
    new_n3320_1, new_n3321, new_n3322, new_n3323, new_n3324_1, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332_1, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343_1,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349_1,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366_1, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390_1, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425_1, new_n3426_1, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439,
    new_n3440, new_n3441, new_n3442, new_n3443, new_n3444, new_n3445,
    new_n3446, new_n3447, new_n3448, new_n3449, new_n3450, new_n3451_1,
    new_n3452, new_n3453, new_n3454, new_n3455, new_n3456, new_n3457,
    new_n3458, new_n3459_1, new_n3460_1, new_n3461, new_n3462, new_n3463,
    new_n3464, new_n3465, new_n3466, new_n3467, new_n3468_1, new_n3469,
    new_n3470, new_n3471, new_n3472, new_n3473, new_n3474, new_n3475,
    new_n3476, new_n3477, new_n3478, new_n3479, new_n3480_1, new_n3481,
    new_n3482, new_n3483, new_n3484, new_n3485, new_n3486, new_n3487,
    new_n3488, new_n3489, new_n3490, new_n3491, new_n3492, new_n3493,
    new_n3494, new_n3495, new_n3496, new_n3497, new_n3498, new_n3499,
    new_n3500, new_n3501, new_n3502_1, new_n3503, new_n3504, new_n3505,
    new_n3506_1, new_n3507, new_n3508, new_n3509, new_n3510, new_n3511,
    new_n3512, new_n3513, new_n3514, new_n3515, new_n3516_1, new_n3517,
    new_n3518, new_n3519, new_n3520, new_n3521, new_n3522, new_n3523,
    new_n3524, new_n3525, new_n3526, new_n3527, new_n3528_1, new_n3529,
    new_n3530, new_n3531, new_n3532, new_n3533, new_n3534, new_n3535,
    new_n3536, new_n3537, new_n3538, new_n3539, new_n3540, new_n3541_1,
    new_n3542, new_n3543, new_n3544, new_n3545, new_n3546, new_n3547,
    new_n3548, new_n3549, new_n3550, new_n3551, new_n3552, new_n3553,
    new_n3554, new_n3555_1, new_n3556, new_n3557, new_n3558, new_n3559,
    new_n3560, new_n3561_1, new_n3562, new_n3563_1, new_n3564, new_n3565,
    new_n3566, new_n3567, new_n3568, new_n3569, new_n3570_1, new_n3571,
    new_n3572, new_n3573, new_n3574, new_n3575, new_n3576, new_n3577,
    new_n3578, new_n3579, new_n3580, new_n3581, new_n3582_1, new_n3583,
    new_n3584, new_n3585, new_n3586, new_n3587, new_n3588, new_n3589,
    new_n3590, new_n3591, new_n3592, new_n3593, new_n3594, new_n3595,
    new_n3596, new_n3597, new_n3598, new_n3599, new_n3600, new_n3601,
    new_n3602, new_n3603, new_n3604, new_n3605, new_n3606, new_n3607,
    new_n3608, new_n3609, new_n3610, new_n3611, new_n3612, new_n3613,
    new_n3614, new_n3615, new_n3616, new_n3617_1, new_n3618_1, new_n3619,
    new_n3620, new_n3621, new_n3622, new_n3623, new_n3624, new_n3625,
    new_n3626, new_n3627, new_n3628, new_n3629, new_n3630, new_n3631,
    new_n3632, new_n3633, new_n3634, new_n3635, new_n3636, new_n3637,
    new_n3638, new_n3639, new_n3640, new_n3641, new_n3642_1, new_n3643,
    new_n3644, new_n3645, new_n3646, new_n3647, new_n3648, new_n3649_1,
    new_n3650, new_n3651, new_n3652, new_n3653, new_n3654, new_n3655,
    new_n3656, new_n3657, new_n3658, new_n3659, new_n3660, new_n3661,
    new_n3662, new_n3663, new_n3664, new_n3665_1, new_n3666, new_n3667,
    new_n3668, new_n3669, new_n3670, new_n3671, new_n3672, new_n3673,
    new_n3674, new_n3675, new_n3676, new_n3677, new_n3678, new_n3679_1,
    new_n3680, new_n3681, new_n3682, new_n3683, new_n3684, new_n3685,
    new_n3686, new_n3687, new_n3688, new_n3689, new_n3690, new_n3691,
    new_n3692, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710_1,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725_1, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733_1, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740_1,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755_1, new_n3756, new_n3757, new_n3758_1,
    new_n3759, new_n3760_1, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781_1, new_n3782,
    new_n3783, new_n3784, new_n3785_1, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794_1,
    new_n3795_1, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828_1, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849, new_n3850_1, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860,
    new_n3861, new_n3862, new_n3863, new_n3864, new_n3865, new_n3866,
    new_n3867, new_n3868, new_n3869_1, new_n3870, new_n3871_1, new_n3872,
    new_n3873, new_n3874, new_n3875, new_n3876, new_n3877, new_n3878,
    new_n3879, new_n3880, new_n3881, new_n3882, new_n3883, new_n3884,
    new_n3885, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890,
    new_n3891_1, new_n3892, new_n3893, new_n3894, new_n3895, new_n3896,
    new_n3897, new_n3898, new_n3899, new_n3900, new_n3901, new_n3902,
    new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908,
    new_n3909_1, new_n3910, new_n3911, new_n3912, new_n3913, new_n3914,
    new_n3915, new_n3916, new_n3917, new_n3918_1, new_n3919, new_n3920,
    new_n3921, new_n3922, new_n3923, new_n3924, new_n3925_1, new_n3926,
    new_n3927, new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1,
    new_n3933, new_n3934_1, new_n3935, new_n3936, new_n3937, new_n3938,
    new_n3939, new_n3940, new_n3941, new_n3942, new_n3943, new_n3944,
    new_n3945_1, new_n3946, new_n3947, new_n3948, new_n3949, new_n3950,
    new_n3951, new_n3952_1, new_n3953, new_n3954, new_n3955, new_n3956,
    new_n3957, new_n3958, new_n3959_1, new_n3960, new_n3961, new_n3962_1,
    new_n3963, new_n3964, new_n3965, new_n3966, new_n3967, new_n3968,
    new_n3969, new_n3970, new_n3971_1, new_n3972, new_n3973, new_n3974,
    new_n3975, new_n3976, new_n3977, new_n3978, new_n3979, new_n3980,
    new_n3981, new_n3982, new_n3983_1, new_n3984_1, new_n3985, new_n3986,
    new_n3987, new_n3988, new_n3989, new_n3990, new_n3991, new_n3992,
    new_n3993, new_n3994, new_n3995, new_n3996, new_n3997, new_n3998,
    new_n3999, new_n4000_1, new_n4001, new_n4002, new_n4003, new_n4004,
    new_n4005, new_n4006, new_n4007, new_n4008, new_n4009, new_n4010_1,
    new_n4011, new_n4012, new_n4013, new_n4014_1, new_n4015, new_n4016,
    new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022,
    new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028,
    new_n4029, new_n4030, new_n4031, new_n4032, new_n4033, new_n4034,
    new_n4035, new_n4036, new_n4037, new_n4038, new_n4039, new_n4040,
    new_n4041, new_n4042, new_n4043, new_n4044, new_n4045, new_n4046,
    new_n4047, new_n4048, new_n4049, new_n4050, new_n4051, new_n4052,
    new_n4053, new_n4054, new_n4055, new_n4056, new_n4057, new_n4058,
    new_n4059, new_n4060, new_n4061, new_n4062, new_n4064, new_n4065,
    new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071_1,
    new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083,
    new_n4084, new_n4085_1, new_n4086, new_n4087, new_n4088_1, new_n4089_1,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4094, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100_1, new_n4101,
    new_n4102, new_n4103_1, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119_1,
    new_n4120, new_n4121, new_n4122, new_n4123_1, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134_1, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141, new_n4142, new_n4143,
    new_n4144, new_n4145, new_n4146_1, new_n4147, new_n4148, new_n4149,
    new_n4150_1, new_n4151_1, new_n4152_1, new_n4153_1, new_n4154,
    new_n4155, new_n4156, new_n4157, new_n4158, new_n4159, new_n4160,
    new_n4161, new_n4162, new_n4163, new_n4164, new_n4165_1, new_n4166,
    new_n4167, new_n4168, new_n4169, new_n4170, new_n4171, new_n4172_1,
    new_n4173_1, new_n4174, new_n4175, new_n4176_1, new_n4177, new_n4178,
    new_n4179, new_n4180, new_n4181, new_n4182, new_n4183, new_n4184,
    new_n4185, new_n4186_1, new_n4187, new_n4188, new_n4189, new_n4190,
    new_n4191, new_n4192, new_n4193, new_n4194, new_n4195, new_n4196,
    new_n4197, new_n4198, new_n4199, new_n4200, new_n4201, new_n4202,
    new_n4203, new_n4204_1, new_n4205_1, new_n4206, new_n4207, new_n4208,
    new_n4209, new_n4210, new_n4211, new_n4212, new_n4213, new_n4214,
    new_n4215_1, new_n4216, new_n4217, new_n4218, new_n4219, new_n4220,
    new_n4221_1, new_n4222, new_n4223, new_n4224_1, new_n4225, new_n4226,
    new_n4227, new_n4228, new_n4229, new_n4230, new_n4231_1, new_n4232,
    new_n4233, new_n4234, new_n4235, new_n4236, new_n4237, new_n4238,
    new_n4239, new_n4240, new_n4241, new_n4242, new_n4243, new_n4244,
    new_n4245, new_n4246, new_n4247, new_n4248, new_n4249, new_n4250,
    new_n4251, new_n4252, new_n4253, new_n4254, new_n4255, new_n4256_1,
    new_n4257, new_n4258, new_n4259, new_n4260, new_n4261, new_n4262,
    new_n4263, new_n4264, new_n4265, new_n4266_1, new_n4267, new_n4268,
    new_n4269, new_n4270, new_n4271, new_n4272_1, new_n4273, new_n4274,
    new_n4275, new_n4276, new_n4277, new_n4278, new_n4279, new_n4280,
    new_n4281, new_n4282, new_n4283, new_n4284, new_n4285, new_n4286,
    new_n4287, new_n4288, new_n4289, new_n4290, new_n4291, new_n4292,
    new_n4293, new_n4294, new_n4295, new_n4296, new_n4297, new_n4298,
    new_n4299, new_n4300, new_n4301, new_n4302, new_n4303, new_n4304,
    new_n4305, new_n4306_1, new_n4307, new_n4308, new_n4309, new_n4310,
    new_n4311, new_n4312, new_n4313, new_n4315, new_n4316, new_n4317,
    new_n4318, new_n4319_1, new_n4320, new_n4321, new_n4322, new_n4323,
    new_n4324, new_n4325_1, new_n4326_1, new_n4327, new_n4328, new_n4329,
    new_n4330, new_n4331, new_n4332, new_n4333, new_n4334, new_n4335,
    new_n4336, new_n4337, new_n4338, new_n4339, new_n4340_1, new_n4341,
    new_n4342, new_n4343, new_n4344, new_n4345, new_n4346, new_n4347,
    new_n4348, new_n4349, new_n4350, new_n4351, new_n4352, new_n4353,
    new_n4354, new_n4355, new_n4356, new_n4357, new_n4358, new_n4359,
    new_n4360, new_n4361, new_n4362, new_n4363, new_n4364, new_n4365,
    new_n4366, new_n4367, new_n4368, new_n4369, new_n4370, new_n4371,
    new_n4372, new_n4373, new_n4374_1, new_n4375, new_n4376_1, new_n4377,
    new_n4378, new_n4379, new_n4380, new_n4381, new_n4382, new_n4383,
    new_n4384, new_n4385, new_n4386, new_n4387, new_n4388, new_n4389,
    new_n4390, new_n4391, new_n4392, new_n4393, new_n4394, new_n4395,
    new_n4396, new_n4397, new_n4398, new_n4399, new_n4400, new_n4401_1,
    new_n4402, new_n4403, new_n4404, new_n4405, new_n4406, new_n4407,
    new_n4408, new_n4409_1, new_n4410, new_n4411, new_n4412, new_n4413,
    new_n4414, new_n4415, new_n4416, new_n4417, new_n4418, new_n4419,
    new_n4420, new_n4421, new_n4422, new_n4423, new_n4424_1, new_n4425,
    new_n4426_1, new_n4427, new_n4428, new_n4429, new_n4430, new_n4431,
    new_n4432_1, new_n4433, new_n4434, new_n4435, new_n4436, new_n4437,
    new_n4438, new_n4439, new_n4440, new_n4441_1, new_n4442, new_n4443,
    new_n4444, new_n4445, new_n4446, new_n4447, new_n4448, new_n4449,
    new_n4450, new_n4451_1, new_n4452, new_n4453, new_n4454, new_n4455,
    new_n4456, new_n4457, new_n4458, new_n4459, new_n4460, new_n4461,
    new_n4462, new_n4463, new_n4464, new_n4465, new_n4466, new_n4467,
    new_n4468, new_n4469, new_n4470, new_n4471, new_n4472, new_n4473,
    new_n4474, new_n4475, new_n4476_1, new_n4477, new_n4478_1, new_n4479,
    new_n4480, new_n4481, new_n4482, new_n4483, new_n4484, new_n4485,
    new_n4486, new_n4487, new_n4488, new_n4489, new_n4490, new_n4491,
    new_n4492, new_n4493, new_n4494, new_n4495, new_n4496, new_n4497,
    new_n4498, new_n4499, new_n4500, new_n4501, new_n4502, new_n4503,
    new_n4504, new_n4505, new_n4506, new_n4507, new_n4508, new_n4509,
    new_n4510, new_n4511, new_n4512, new_n4513, new_n4514_1, new_n4515,
    new_n4516, new_n4517, new_n4518, new_n4519, new_n4520, new_n4521,
    new_n4522, new_n4523, new_n4524, new_n4525, new_n4526, new_n4527,
    new_n4528, new_n4529_1, new_n4530, new_n4531, new_n4532, new_n4534,
    new_n4535, new_n4536, new_n4537, new_n4538, new_n4539, new_n4540,
    new_n4541, new_n4542, new_n4543, new_n4544, new_n4545, new_n4546,
    new_n4547, new_n4548, new_n4549, new_n4550, new_n4551, new_n4552_1,
    new_n4553, new_n4554, new_n4555, new_n4556, new_n4557, new_n4558,
    new_n4559, new_n4560, new_n4561, new_n4562, new_n4563, new_n4564,
    new_n4565, new_n4566, new_n4567, new_n4568, new_n4569, new_n4570,
    new_n4571, new_n4572, new_n4573, new_n4574, new_n4575, new_n4576,
    new_n4577, new_n4578, new_n4579, new_n4580, new_n4581, new_n4582,
    new_n4583, new_n4584, new_n4585, new_n4586, new_n4587, new_n4588_1,
    new_n4589, new_n4590_1, new_n4591, new_n4592, new_n4593, new_n4594,
    new_n4595_1, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600,
    new_n4601, new_n4602, new_n4603, new_n4604, new_n4605, new_n4606,
    new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612,
    new_n4613, new_n4614, new_n4615, new_n4616, new_n4617, new_n4618,
    new_n4620, new_n4621, new_n4622, new_n4623, new_n4624_1, new_n4625,
    new_n4626, new_n4627, new_n4628, new_n4629, new_n4630, new_n4631,
    new_n4632, new_n4633, new_n4634, new_n4635, new_n4636, new_n4637,
    new_n4638, new_n4639, new_n4640, new_n4641, new_n4642, new_n4643,
    new_n4644, new_n4645, new_n4646_1, new_n4647, new_n4648, new_n4649,
    new_n4650, new_n4651, new_n4652, new_n4653, new_n4654, new_n4655,
    new_n4656, new_n4657, new_n4658, new_n4659, new_n4660, new_n4661,
    new_n4662, new_n4663, new_n4664, new_n4665_1, new_n4666, new_n4667,
    new_n4668, new_n4669, new_n4670, new_n4671, new_n4672, new_n4673,
    new_n4674_1, new_n4675, new_n4676, new_n4677, new_n4678, new_n4679,
    new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685,
    new_n4686, new_n4687, new_n4688, new_n4689, new_n4690, new_n4691,
    new_n4692, new_n4693_1, new_n4694, new_n4695, new_n4696, new_n4697,
    new_n4698, new_n4699, new_n4700, new_n4701, new_n4702, new_n4703,
    new_n4704, new_n4705, new_n4706, new_n4707, new_n4708, new_n4709,
    new_n4710, new_n4711, new_n4712, new_n4713, new_n4714, new_n4715,
    new_n4716, new_n4717, new_n4718, new_n4719, new_n4720, new_n4721,
    new_n4722_1, new_n4723, new_n4724, new_n4725, new_n4726, new_n4727,
    new_n4728, new_n4729, new_n4730, new_n4731_1, new_n4732, new_n4733,
    new_n4734, new_n4735, new_n4736, new_n4737, new_n4738, new_n4739,
    new_n4740, new_n4741, new_n4742, new_n4743, new_n4744, new_n4745_1,
    new_n4746, new_n4747_1, new_n4748, new_n4749, new_n4750, new_n4751,
    new_n4752, new_n4753, new_n4754, new_n4755, new_n4756, new_n4757,
    new_n4758, new_n4759, new_n4760, new_n4761, new_n4762, new_n4763,
    new_n4764, new_n4765, new_n4766_1, new_n4767, new_n4768, new_n4769,
    new_n4770_1, new_n4771, new_n4772, new_n4773, new_n4774, new_n4775,
    new_n4776, new_n4777_1, new_n4778, new_n4779, new_n4780, new_n4781,
    new_n4782, new_n4783, new_n4784, new_n4785_1, new_n4786, new_n4787,
    new_n4788, new_n4789, new_n4790, new_n4791, new_n4792, new_n4793,
    new_n4794, new_n4795, new_n4796, new_n4797, new_n4798, new_n4799,
    new_n4800, new_n4801, new_n4802, new_n4803, new_n4804_1, new_n4805,
    new_n4806, new_n4807, new_n4808, new_n4809, new_n4810_1, new_n4812_1,
    new_n4813, new_n4814_1, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850_1, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858_1, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891_1, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913_1, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925_1, new_n4926,
    new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932,
    new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938,
    new_n4939_1, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947_1, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952_1, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957_1, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964_1, new_n4965, new_n4966_1, new_n4967_1, new_n4968,
    new_n4969, new_n4970, new_n4971, new_n4972_1, new_n4973, new_n4974,
    new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980,
    new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986,
    new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998,
    new_n4999, new_n5000, new_n5001, new_n5002, new_n5003, new_n5004,
    new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010,
    new_n5011_1, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016,
    new_n5017, new_n5018, new_n5019, new_n5020_1, new_n5021, new_n5022,
    new_n5023, new_n5024_1, new_n5025_1, new_n5026_1, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031_1, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046_1,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060_1, new_n5061, new_n5062_1, new_n5063, new_n5064_1,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077_1, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082_1,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098_1, new_n5099, new_n5100,
    new_n5101_1, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115_1, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120_1, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128_1, new_n5129, new_n5130,
    new_n5131_1, new_n5132, new_n5133, new_n5134, new_n5136, new_n5137,
    new_n5138, new_n5139, new_n5140_1, new_n5141, new_n5142, new_n5143,
    new_n5144, new_n5145, new_n5146, new_n5147, new_n5148, new_n5149,
    new_n5150, new_n5151, new_n5152, new_n5153, new_n5154, new_n5155,
    new_n5156, new_n5157, new_n5158_1, new_n5159, new_n5160, new_n5161,
    new_n5162, new_n5163, new_n5164, new_n5165, new_n5166, new_n5167,
    new_n5168_1, new_n5169, new_n5170, new_n5171, new_n5172, new_n5173,
    new_n5174, new_n5175, new_n5176, new_n5177, new_n5178, new_n5179,
    new_n5180, new_n5181, new_n5182, new_n5183, new_n5184_1, new_n5185,
    new_n5186, new_n5187, new_n5188, new_n5189, new_n5190, new_n5191,
    new_n5192, new_n5193, new_n5194, new_n5195, new_n5196, new_n5197,
    new_n5198, new_n5199, new_n5200, new_n5201, new_n5202, new_n5203,
    new_n5204, new_n5205, new_n5206, new_n5207, new_n5208, new_n5209,
    new_n5210, new_n5211_1, new_n5212, new_n5213_1, new_n5214, new_n5215,
    new_n5216, new_n5217, new_n5218, new_n5219, new_n5220, new_n5221,
    new_n5222, new_n5223, new_n5224, new_n5225, new_n5226_1, new_n5227,
    new_n5228_1, new_n5229, new_n5230, new_n5231, new_n5232, new_n5233,
    new_n5234, new_n5235, new_n5236, new_n5237, new_n5238, new_n5239,
    new_n5240, new_n5241, new_n5242, new_n5243, new_n5244, new_n5245,
    new_n5246, new_n5247, new_n5248, new_n5249, new_n5250, new_n5251,
    new_n5252, new_n5253, new_n5254, new_n5255_1, new_n5256_1, new_n5257,
    new_n5258, new_n5259, new_n5260, new_n5261, new_n5262, new_n5263,
    new_n5264, new_n5265_1, new_n5266, new_n5267, new_n5268, new_n5269,
    new_n5270, new_n5271, new_n5272, new_n5273_1, new_n5274_1, new_n5275,
    new_n5276, new_n5277, new_n5278, new_n5279, new_n5280, new_n5281,
    new_n5282, new_n5283, new_n5284, new_n5285, new_n5286, new_n5287,
    new_n5288, new_n5289, new_n5290, new_n5291, new_n5292, new_n5293,
    new_n5294, new_n5295, new_n5296, new_n5297, new_n5298, new_n5299,
    new_n5300_1, new_n5301, new_n5302_1, new_n5303, new_n5304, new_n5305,
    new_n5306, new_n5307, new_n5308, new_n5309, new_n5310, new_n5311,
    new_n5312, new_n5313, new_n5314, new_n5315, new_n5316, new_n5317,
    new_n5318, new_n5319, new_n5320, new_n5321, new_n5322, new_n5323,
    new_n5324, new_n5326, new_n5327, new_n5328, new_n5329, new_n5330_1,
    new_n5331, new_n5332, new_n5333, new_n5334, new_n5335, new_n5336,
    new_n5337_1, new_n5338, new_n5339, new_n5340, new_n5341, new_n5342,
    new_n5343, new_n5344, new_n5345, new_n5346, new_n5347, new_n5348,
    new_n5349, new_n5350, new_n5351_1, new_n5352, new_n5353_1, new_n5354,
    new_n5355, new_n5356, new_n5357, new_n5358, new_n5359, new_n5360,
    new_n5361, new_n5362, new_n5363, new_n5364, new_n5365, new_n5366,
    new_n5367, new_n5368, new_n5369, new_n5370, new_n5371, new_n5372,
    new_n5373, new_n5374, new_n5375, new_n5376_1, new_n5377, new_n5378,
    new_n5379, new_n5380, new_n5381, new_n5382, new_n5383, new_n5384,
    new_n5385, new_n5386_1, new_n5387, new_n5388, new_n5389, new_n5390,
    new_n5391, new_n5392, new_n5393, new_n5394, new_n5395, new_n5396,
    new_n5397, new_n5398, new_n5399_1, new_n5400_1, new_n5401, new_n5402,
    new_n5403_1, new_n5404, new_n5405, new_n5406, new_n5407, new_n5408,
    new_n5409, new_n5410, new_n5411, new_n5412, new_n5413, new_n5414,
    new_n5415, new_n5416, new_n5417, new_n5418, new_n5419, new_n5420,
    new_n5421, new_n5422, new_n5423, new_n5424, new_n5425, new_n5426,
    new_n5427, new_n5428, new_n5429, new_n5430_1, new_n5431, new_n5432,
    new_n5433, new_n5434, new_n5435, new_n5436, new_n5437, new_n5438_1,
    new_n5439_1, new_n5440, new_n5441, new_n5442, new_n5443_1, new_n5444,
    new_n5445, new_n5446, new_n5447, new_n5448, new_n5449, new_n5450,
    new_n5451_1, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456,
    new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462,
    new_n5463, new_n5464, new_n5465, new_n5466, new_n5467, new_n5468,
    new_n5469, new_n5470, new_n5471, new_n5472_1, new_n5473, new_n5474,
    new_n5475, new_n5476, new_n5477, new_n5478, new_n5479, new_n5480,
    new_n5481, new_n5482, new_n5483, new_n5484, new_n5485_1, new_n5486,
    new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492,
    new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498,
    new_n5499, new_n5500, new_n5501, new_n5502, new_n5503, new_n5504,
    new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510,
    new_n5511, new_n5512, new_n5513, new_n5514, new_n5515, new_n5516,
    new_n5517_1, new_n5518, new_n5519, new_n5520, new_n5521_1, new_n5522,
    new_n5523, new_n5524_1, new_n5525, new_n5526, new_n5527, new_n5528,
    new_n5529, new_n5530, new_n5531, new_n5532_1, new_n5533, new_n5534,
    new_n5535, new_n5536, new_n5537, new_n5538, new_n5539, new_n5540,
    new_n5541, new_n5542, new_n5543, new_n5544, new_n5545, new_n5546,
    new_n5547, new_n5548, new_n5549, new_n5550, new_n5551, new_n5552,
    new_n5553, new_n5554, new_n5555, new_n5556, new_n5557, new_n5558,
    new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564_1,
    new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570,
    new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576,
    new_n5577, new_n5578, new_n5579_1, new_n5580, new_n5581, new_n5582,
    new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588,
    new_n5589, new_n5590, new_n5591, new_n5592, new_n5593_1, new_n5594,
    new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600,
    new_n5601, new_n5602, new_n5603_1, new_n5604, new_n5605_1, new_n5606,
    new_n5607, new_n5608, new_n5609_1, new_n5610, new_n5611, new_n5612,
    new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618,
    new_n5619, new_n5620, new_n5621, new_n5622, new_n5623, new_n5624,
    new_n5625, new_n5626, new_n5627, new_n5628, new_n5629, new_n5630,
    new_n5631, new_n5632, new_n5633, new_n5634_1, new_n5635, new_n5636,
    new_n5637, new_n5638, new_n5639, new_n5640, new_n5641, new_n5642,
    new_n5643_1, new_n5644, new_n5645, new_n5646, new_n5647, new_n5648,
    new_n5649, new_n5650, new_n5651, new_n5652, new_n5653, new_n5654,
    new_n5655, new_n5656, new_n5657, new_n5658, new_n5659, new_n5660,
    new_n5661, new_n5663, new_n5664, new_n5665, new_n5666, new_n5667,
    new_n5668, new_n5669, new_n5670, new_n5671, new_n5672, new_n5673,
    new_n5674, new_n5675, new_n5676, new_n5677, new_n5678, new_n5679,
    new_n5680_1, new_n5681, new_n5682, new_n5683, new_n5684, new_n5685,
    new_n5686, new_n5687_1, new_n5688, new_n5689, new_n5690, new_n5691,
    new_n5692, new_n5693, new_n5694, new_n5695, new_n5696_1, new_n5697,
    new_n5698, new_n5699, new_n5700_1, new_n5701, new_n5702, new_n5703,
    new_n5704_1, new_n5705, new_n5706, new_n5707, new_n5708, new_n5709,
    new_n5710, new_n5711, new_n5712, new_n5713, new_n5714, new_n5715,
    new_n5716, new_n5717, new_n5718, new_n5719, new_n5720, new_n5721,
    new_n5722, new_n5723, new_n5724, new_n5725, new_n5726, new_n5727,
    new_n5728, new_n5729, new_n5730, new_n5731, new_n5732_1, new_n5733,
    new_n5734, new_n5735, new_n5736, new_n5737, new_n5738, new_n5739,
    new_n5740, new_n5742_1, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752_1,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765_1, new_n5766, new_n5767, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776_1,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782_1,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822_1, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833_1, new_n5834_1, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840_1, new_n5841_1, new_n5842_1,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850_1, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857, new_n5858, new_n5859, new_n5860,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882_1, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5889, new_n5890, new_n5891,
    new_n5892, new_n5893, new_n5894, new_n5895, new_n5896, new_n5897,
    new_n5898, new_n5899, new_n5900, new_n5901, new_n5902, new_n5903_1,
    new_n5904_1, new_n5905, new_n5906, new_n5907, new_n5908, new_n5909,
    new_n5910, new_n5911_1, new_n5912, new_n5913, new_n5914, new_n5915,
    new_n5916, new_n5917, new_n5918, new_n5919, new_n5920, new_n5921,
    new_n5922, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927,
    new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933,
    new_n5934, new_n5935, new_n5936_1, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943_1, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980_1, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012_1, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022_1, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031_1, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044_1, new_n6045, new_n6046_1, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084_1, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104_1, new_n6105_1, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160_1, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6168,
    new_n6169, new_n6170, new_n6171_1, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183_1, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189_1, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204_1,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218_1, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223_1, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233_1, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245_1, new_n6246,
    new_n6247, new_n6248_1, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256_1, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271_1, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276_1,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308_1, new_n6309, new_n6310, new_n6311_1, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323_1, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330_1,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339_1, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354_1,
    new_n6355, new_n6356_1, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369_1, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375_1, new_n6376, new_n6377, new_n6378,
    new_n6379_1, new_n6380, new_n6381_1, new_n6382, new_n6383_1, new_n6384,
    new_n6385_1, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397_1, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407_1, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427_1, new_n6428, new_n6429, new_n6430, new_n6431_1, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437_1, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456_1,
    new_n6457_1, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465_1, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470_1, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476_1, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485_1, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502_1, new_n6503, new_n6504,
    new_n6505, new_n6506_1, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513_1, new_n6514_1, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542_1, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556_1, new_n6557, new_n6558_1, new_n6560_1,
    new_n6561, new_n6562, new_n6563, new_n6564, new_n6565, new_n6566,
    new_n6567_1, new_n6568, new_n6569, new_n6570, new_n6571, new_n6573,
    new_n6575, new_n6576_1, new_n6577, new_n6578, new_n6579, new_n6580,
    new_n6581, new_n6582, new_n6583, new_n6584, new_n6585, new_n6586,
    new_n6587_1, new_n6588, new_n6589, new_n6590_1, new_n6591, new_n6592,
    new_n6593, new_n6594, new_n6595, new_n6596_1, new_n6597, new_n6598,
    new_n6599, new_n6600, new_n6601, new_n6602, new_n6603, new_n6604,
    new_n6605, new_n6606, new_n6607, new_n6608, new_n6609, new_n6611_1,
    new_n6612_1, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628_1, new_n6629,
    new_n6630_1, new_n6631_1, new_n6632, new_n6633, new_n6634_1, new_n6635,
    new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641,
    new_n6642, new_n6643, new_n6644, new_n6647, new_n6649, new_n6650,
    new_n6651, new_n6652_1, new_n6653, new_n6654, new_n6655_1, new_n6656,
    new_n6657, new_n6658, new_n6659_1, new_n6660, new_n6661, new_n6662,
    new_n6663, new_n6664, new_n6665, new_n6666, new_n6667, new_n6668,
    new_n6669_1, new_n6670, new_n6671_1, new_n6672, new_n6673_1,
    new_n6674_1, new_n6675, new_n6676, new_n6677, new_n6678, new_n6679,
    new_n6680, new_n6681, new_n6682, new_n6683, new_n6684_1, new_n6685,
    new_n6686, new_n6687, new_n6688, new_n6689, new_n6690, new_n6691_1,
    new_n6692, new_n6693, new_n6694, new_n6695, new_n6696, new_n6697,
    new_n6698, new_n6699, new_n6700, new_n6701, new_n6702, new_n6703,
    new_n6704, new_n6705, new_n6706_1, new_n6707_1, new_n6708, new_n6709,
    new_n6710, new_n6711, new_n6712, new_n6713, new_n6714, new_n6715,
    new_n6716, new_n6717, new_n6718, new_n6719, new_n6720, new_n6721,
    new_n6722, new_n6723, new_n6724, new_n6725, new_n6726, new_n6727,
    new_n6728, new_n6729_1, new_n6730, new_n6731, new_n6732, new_n6733,
    new_n6734, new_n6735, new_n6736_1, new_n6737, new_n6738, new_n6739,
    new_n6740, new_n6741, new_n6742, new_n6743, new_n6744, new_n6745,
    new_n6746, new_n6747, new_n6748, new_n6749, new_n6750, new_n6751,
    new_n6752, new_n6753, new_n6754, new_n6755, new_n6756, new_n6757,
    new_n6758, new_n6759, new_n6760, new_n6761, new_n6762, new_n6763,
    new_n6764, new_n6765, new_n6766, new_n6767, new_n6768, new_n6769,
    new_n6770, new_n6771, new_n6772, new_n6773_1, new_n6774, new_n6775_1,
    new_n6776, new_n6777, new_n6778, new_n6779, new_n6780, new_n6781,
    new_n6782, new_n6783, new_n6784, new_n6785_1, new_n6786, new_n6787,
    new_n6788, new_n6789, new_n6790_1, new_n6791_1, new_n6792, new_n6793,
    new_n6794_1, new_n6795, new_n6796, new_n6797, new_n6798, new_n6799,
    new_n6800, new_n6801, new_n6802_1, new_n6803, new_n6804, new_n6805,
    new_n6806, new_n6807, new_n6808, new_n6809, new_n6810, new_n6811,
    new_n6812, new_n6813, new_n6814_1, new_n6815, new_n6816, new_n6817,
    new_n6818, new_n6819, new_n6820, new_n6821, new_n6822, new_n6823,
    new_n6824, new_n6825, new_n6826_1, new_n6827, new_n6828, new_n6829,
    new_n6830, new_n6831, new_n6832, new_n6833, new_n6834, new_n6835_1,
    new_n6836, new_n6837, new_n6838, new_n6839, new_n6840, new_n6841,
    new_n6842, new_n6843, new_n6844, new_n6845, new_n6846, new_n6847,
    new_n6848, new_n6849, new_n6850, new_n6851, new_n6852, new_n6853_1,
    new_n6854, new_n6855, new_n6856, new_n6857, new_n6858, new_n6859,
    new_n6860, new_n6861_1, new_n6862_1, new_n6863_1, new_n6864, new_n6865,
    new_n6866, new_n6867_1, new_n6868, new_n6869, new_n6870, new_n6871,
    new_n6872, new_n6873, new_n6874, new_n6875, new_n6876, new_n6877,
    new_n6878, new_n6879, new_n6880, new_n6881, new_n6882, new_n6883,
    new_n6884, new_n6885, new_n6886, new_n6887, new_n6888, new_n6889,
    new_n6890, new_n6891, new_n6892, new_n6893, new_n6894, new_n6895,
    new_n6896, new_n6897, new_n6898, new_n6899, new_n6900, new_n6901,
    new_n6902, new_n6903, new_n6904, new_n6905, new_n6906, new_n6907,
    new_n6908, new_n6909, new_n6910, new_n6911, new_n6912, new_n6913,
    new_n6914, new_n6915, new_n6916, new_n6917, new_n6918, new_n6919,
    new_n6920, new_n6921, new_n6922, new_n6923, new_n6924, new_n6925,
    new_n6926, new_n6927, new_n6928, new_n6929, new_n6930, new_n6931,
    new_n6932, new_n6933, new_n6934, new_n6935, new_n6936, new_n6937,
    new_n6938, new_n6939, new_n6940, new_n6941, new_n6942, new_n6943,
    new_n6944, new_n6945, new_n6946, new_n6947, new_n6948, new_n6949,
    new_n6950, new_n6951, new_n6952, new_n6953, new_n6954, new_n6955,
    new_n6956, new_n6957, new_n6958, new_n6959, new_n6960, new_n6961,
    new_n6962, new_n6963, new_n6964, new_n6965_1, new_n6966, new_n6967_1,
    new_n6968, new_n6969, new_n6970, new_n6971_1, new_n6972, new_n6973,
    new_n6974, new_n6975_1, new_n6976, new_n6977, new_n6978, new_n6979,
    new_n6980, new_n6981, new_n6982, new_n6983_1, new_n6984, new_n6985_1,
    new_n6986, new_n6987, new_n6988, new_n6989, new_n6991, new_n6992,
    new_n6993, new_n6994, new_n6995, new_n6996, new_n6997, new_n6998_1,
    new_n6999, new_n7000, new_n7001, new_n7002, new_n7003, new_n7004,
    new_n7005, new_n7006, new_n7007, new_n7008, new_n7009, new_n7010,
    new_n7011, new_n7012, new_n7013, new_n7014, new_n7015, new_n7016,
    new_n7017, new_n7018, new_n7019, new_n7020, new_n7021, new_n7022,
    new_n7023, new_n7024, new_n7025, new_n7026_1, new_n7027, new_n7028,
    new_n7029, new_n7030, new_n7031, new_n7032_1, new_n7033, new_n7034,
    new_n7035, new_n7036, new_n7037, new_n7038_1, new_n7039, new_n7040,
    new_n7041, new_n7042, new_n7043, new_n7044, new_n7045, new_n7046,
    new_n7047, new_n7048, new_n7049, new_n7050, new_n7051, new_n7052,
    new_n7053, new_n7054, new_n7055, new_n7056, new_n7057_1, new_n7058,
    new_n7059, new_n7060, new_n7061, new_n7062, new_n7063, new_n7064,
    new_n7065, new_n7066, new_n7067, new_n7068, new_n7069, new_n7070,
    new_n7071, new_n7072, new_n7073, new_n7074, new_n7075, new_n7076,
    new_n7077, new_n7078, new_n7079_1, new_n7080, new_n7081, new_n7082,
    new_n7083, new_n7084, new_n7085, new_n7086, new_n7087, new_n7088,
    new_n7089, new_n7090, new_n7091, new_n7092, new_n7093, new_n7094,
    new_n7095, new_n7096, new_n7097, new_n7098, new_n7099_1, new_n7100,
    new_n7101, new_n7102, new_n7103, new_n7104, new_n7105, new_n7106,
    new_n7107, new_n7108, new_n7109, new_n7110, new_n7111, new_n7112,
    new_n7113, new_n7114, new_n7115, new_n7116, new_n7117, new_n7118,
    new_n7119, new_n7120, new_n7121, new_n7122, new_n7123, new_n7124,
    new_n7125, new_n7126, new_n7127, new_n7128, new_n7129, new_n7130,
    new_n7131, new_n7132, new_n7133, new_n7134, new_n7135, new_n7136,
    new_n7137, new_n7138, new_n7139_1, new_n7140, new_n7141, new_n7142,
    new_n7143, new_n7144, new_n7145, new_n7146, new_n7147, new_n7148,
    new_n7149_1, new_n7150, new_n7151, new_n7152, new_n7153, new_n7154,
    new_n7155, new_n7156, new_n7157, new_n7158, new_n7159, new_n7160,
    new_n7161, new_n7162, new_n7163, new_n7164, new_n7165, new_n7166,
    new_n7167, new_n7168, new_n7169, new_n7170, new_n7171, new_n7172,
    new_n7173, new_n7174, new_n7175, new_n7176, new_n7177, new_n7178,
    new_n7179, new_n7180, new_n7181, new_n7182, new_n7183, new_n7184,
    new_n7185, new_n7186, new_n7187, new_n7188, new_n7189, new_n7190_1,
    new_n7191, new_n7192, new_n7193, new_n7194, new_n7195, new_n7196,
    new_n7197, new_n7198, new_n7199, new_n7200, new_n7201, new_n7202,
    new_n7203, new_n7204, new_n7205, new_n7206, new_n7207, new_n7208,
    new_n7209, new_n7210, new_n7211, new_n7212, new_n7213, new_n7214,
    new_n7215, new_n7216, new_n7217, new_n7218, new_n7219, new_n7220,
    new_n7221, new_n7222, new_n7223, new_n7224, new_n7225, new_n7226,
    new_n7227, new_n7228, new_n7229_1, new_n7230_1, new_n7231, new_n7232,
    new_n7233_1, new_n7234, new_n7235, new_n7236_1, new_n7237, new_n7238,
    new_n7239, new_n7240, new_n7241, new_n7242, new_n7243, new_n7244,
    new_n7245, new_n7246, new_n7247, new_n7248, new_n7249, new_n7250,
    new_n7251, new_n7252, new_n7253_1, new_n7254, new_n7255, new_n7256_1,
    new_n7257, new_n7258, new_n7259, new_n7260, new_n7261, new_n7262,
    new_n7263, new_n7264, new_n7265, new_n7266, new_n7267, new_n7268_1,
    new_n7269, new_n7270, new_n7271, new_n7272, new_n7273, new_n7274,
    new_n7275, new_n7276, new_n7277_1, new_n7278, new_n7279, new_n7280_1,
    new_n7281, new_n7282, new_n7283, new_n7284, new_n7285, new_n7286,
    new_n7287, new_n7288, new_n7289, new_n7290, new_n7291, new_n7292,
    new_n7293, new_n7294, new_n7295, new_n7296, new_n7297, new_n7298_1,
    new_n7299, new_n7300, new_n7301, new_n7303, new_n7304, new_n7305_1,
    new_n7306, new_n7307, new_n7308_1, new_n7309, new_n7310, new_n7311,
    new_n7312, new_n7313_1, new_n7314, new_n7315, new_n7316, new_n7317,
    new_n7318, new_n7319, new_n7320, new_n7321, new_n7322, new_n7323,
    new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329,
    new_n7330_1, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335_1,
    new_n7336, new_n7337, new_n7338, new_n7339_1, new_n7340, new_n7341,
    new_n7342, new_n7343, new_n7344, new_n7345, new_n7346_1, new_n7347,
    new_n7348, new_n7349_1, new_n7350, new_n7351, new_n7352, new_n7353,
    new_n7354, new_n7355, new_n7356, new_n7357, new_n7358, new_n7359,
    new_n7360, new_n7361, new_n7362, new_n7363_1, new_n7364, new_n7365,
    new_n7366, new_n7367, new_n7368, new_n7369, new_n7370, new_n7371,
    new_n7372, new_n7373, new_n7374, new_n7375, new_n7376, new_n7377_1,
    new_n7378, new_n7379, new_n7380, new_n7381, new_n7382, new_n7383,
    new_n7384, new_n7385, new_n7386, new_n7387, new_n7388, new_n7389,
    new_n7390_1, new_n7391, new_n7392, new_n7393, new_n7394, new_n7395,
    new_n7396, new_n7397, new_n7398, new_n7399, new_n7400, new_n7401,
    new_n7402, new_n7403_1, new_n7404, new_n7405, new_n7406, new_n7407,
    new_n7408_1, new_n7409, new_n7410, new_n7411, new_n7412, new_n7413,
    new_n7414, new_n7415, new_n7416, new_n7417, new_n7418, new_n7419,
    new_n7420, new_n7421_1, new_n7422, new_n7423, new_n7424, new_n7425,
    new_n7426, new_n7427, new_n7428_1, new_n7429, new_n7430, new_n7431,
    new_n7432_1, new_n7433, new_n7434, new_n7435, new_n7436, new_n7437_1,
    new_n7438, new_n7439, new_n7440, new_n7441, new_n7442, new_n7443,
    new_n7444, new_n7445, new_n7446, new_n7447, new_n7448, new_n7449,
    new_n7450, new_n7451, new_n7452, new_n7453, new_n7454, new_n7455,
    new_n7456, new_n7457, new_n7458, new_n7459, new_n7460_1, new_n7461,
    new_n7462, new_n7463, new_n7464, new_n7465, new_n7466, new_n7467,
    new_n7468, new_n7469, new_n7470, new_n7471, new_n7472, new_n7473,
    new_n7474, new_n7475_1, new_n7476, new_n7477_1, new_n7478, new_n7479,
    new_n7480, new_n7481, new_n7482, new_n7483, new_n7484, new_n7485,
    new_n7486, new_n7487, new_n7488, new_n7489, new_n7490, new_n7491,
    new_n7492, new_n7493, new_n7494, new_n7495, new_n7496, new_n7497,
    new_n7498, new_n7499, new_n7500, new_n7501, new_n7502, new_n7503,
    new_n7504, new_n7505, new_n7506, new_n7507_1, new_n7508, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514_1, new_n7515, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523,
    new_n7524_1, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558_1, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566_1, new_n7567, new_n7568, new_n7569_1, new_n7570, new_n7571,
    new_n7572_1, new_n7573, new_n7574, new_n7575_1, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585_1, new_n7586, new_n7587, new_n7588_1, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593_1, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598_1, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607_1,
    new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616_1, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630_1, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643_1, new_n7644,
    new_n7645, new_n7646, new_n7647_1, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657_1, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670_1, new_n7671, new_n7672, new_n7673, new_n7674_1,
    new_n7675, new_n7676, new_n7677, new_n7678_1, new_n7679_1, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686_1,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692_1,
    new_n7693_1, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698_1,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708_1, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721_1, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7729,
    new_n7730, new_n7731_1, new_n7732, new_n7733, new_n7734, new_n7735,
    new_n7736, new_n7737, new_n7738, new_n7739, new_n7740, new_n7741,
    new_n7742, new_n7743, new_n7744, new_n7745, new_n7746, new_n7747,
    new_n7748, new_n7749, new_n7750, new_n7751_1, new_n7752, new_n7753,
    new_n7754, new_n7755, new_n7756, new_n7757, new_n7758, new_n7759_1,
    new_n7760, new_n7761, new_n7762, new_n7763, new_n7764, new_n7765,
    new_n7766, new_n7767, new_n7768, new_n7769_1, new_n7770, new_n7771,
    new_n7772, new_n7773_1, new_n7774, new_n7775, new_n7776, new_n7777,
    new_n7778, new_n7779, new_n7780_1, new_n7781, new_n7782, new_n7783,
    new_n7784, new_n7785, new_n7786, new_n7787, new_n7788_1, new_n7789,
    new_n7790, new_n7791, new_n7792, new_n7793, new_n7794_1, new_n7795,
    new_n7796, new_n7797, new_n7798, new_n7799, new_n7800, new_n7801,
    new_n7802, new_n7803, new_n7804, new_n7805, new_n7806, new_n7807,
    new_n7808, new_n7809, new_n7810, new_n7811_1, new_n7812, new_n7813,
    new_n7814, new_n7815, new_n7816, new_n7817, new_n7818, new_n7819,
    new_n7820, new_n7821, new_n7822, new_n7823, new_n7824, new_n7825,
    new_n7826, new_n7827, new_n7828, new_n7829, new_n7830_1, new_n7831,
    new_n7832, new_n7833, new_n7834_1, new_n7835, new_n7836, new_n7837,
    new_n7838, new_n7839, new_n7840, new_n7841_1, new_n7842, new_n7843,
    new_n7844, new_n7845, new_n7846, new_n7847, new_n7848, new_n7849,
    new_n7850, new_n7851, new_n7852, new_n7853, new_n7854, new_n7855,
    new_n7856, new_n7857, new_n7858, new_n7859, new_n7860, new_n7861,
    new_n7862, new_n7863, new_n7864, new_n7865, new_n7866, new_n7867,
    new_n7868, new_n7869, new_n7870, new_n7871, new_n7872, new_n7873,
    new_n7874, new_n7875, new_n7876_1, new_n7877, new_n7878, new_n7879,
    new_n7880, new_n7881, new_n7882, new_n7883, new_n7884_1, new_n7885,
    new_n7886, new_n7887, new_n7888, new_n7889, new_n7890, new_n7891,
    new_n7892, new_n7893, new_n7894, new_n7895, new_n7896, new_n7897,
    new_n7898, new_n7899, new_n7900, new_n7901, new_n7902, new_n7903,
    new_n7904, new_n7905, new_n7906, new_n7907, new_n7908, new_n7909,
    new_n7910, new_n7911, new_n7912, new_n7913, new_n7914, new_n7915,
    new_n7916, new_n7917_1, new_n7918, new_n7919, new_n7920, new_n7921,
    new_n7922, new_n7923, new_n7924, new_n7925, new_n7926, new_n7927,
    new_n7928, new_n7929, new_n7930, new_n7931, new_n7932, new_n7933,
    new_n7934, new_n7935, new_n7936, new_n7937_1, new_n7938, new_n7939,
    new_n7940, new_n7941, new_n7942, new_n7943_1, new_n7944, new_n7945,
    new_n7946, new_n7947, new_n7948, new_n7949_1, new_n7950_1, new_n7951,
    new_n7952, new_n7953, new_n7954, new_n7955, new_n7956, new_n7957,
    new_n7958, new_n7959_1, new_n7960, new_n7961, new_n7962, new_n7963_1,
    new_n7964, new_n7965, new_n7966, new_n7967, new_n7968_1, new_n7969,
    new_n7970, new_n7971, new_n7972, new_n7973, new_n7974, new_n7975,
    new_n7976, new_n7977, new_n7978, new_n7979, new_n7980, new_n7981,
    new_n7982, new_n7983, new_n7984, new_n7985, new_n7986, new_n7987,
    new_n7988, new_n7990, new_n7991, new_n7992_1, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999_1, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006_1,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027_1, new_n8028, new_n8029, new_n8030,
    new_n8031_1, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042_1,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052_1, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067_1, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095_1, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103_1, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109_1, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127_1, new_n8128, new_n8129, new_n8130_1, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135_1, new_n8136, new_n8137, new_n8138,
    new_n8139_1, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148_1, new_n8149_1, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159_1, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179_1, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194_1, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215_1, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244_1, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255_1, new_n8256_1, new_n8257, new_n8258,
    new_n8259_1, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267_1, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8275, new_n8276_1, new_n8277,
    new_n8278, new_n8279, new_n8280, new_n8281, new_n8282, new_n8283,
    new_n8284, new_n8285_1, new_n8286, new_n8287, new_n8288_1, new_n8289,
    new_n8291, new_n8292, new_n8293, new_n8294, new_n8295, new_n8296,
    new_n8297, new_n8298, new_n8299, new_n8300, new_n8301, new_n8302,
    new_n8303, new_n8304, new_n8305_1, new_n8306_1, new_n8307, new_n8308,
    new_n8309_1, new_n8310, new_n8311, new_n8312, new_n8313, new_n8314,
    new_n8315, new_n8316, new_n8317, new_n8318, new_n8319, new_n8320_1,
    new_n8321_1, new_n8322, new_n8323, new_n8324_1, new_n8325, new_n8326,
    new_n8327, new_n8328, new_n8329, new_n8330, new_n8331, new_n8332,
    new_n8333, new_n8334, new_n8335, new_n8336, new_n8337, new_n8338,
    new_n8339_1, new_n8340, new_n8341, new_n8342, new_n8343, new_n8344,
    new_n8345, new_n8346, new_n8347, new_n8348, new_n8349, new_n8350,
    new_n8351, new_n8352, new_n8353, new_n8354, new_n8355, new_n8356,
    new_n8357, new_n8358, new_n8359, new_n8360, new_n8361, new_n8362,
    new_n8363_1, new_n8364, new_n8365, new_n8366, new_n8367, new_n8368,
    new_n8369, new_n8370, new_n8371, new_n8372, new_n8373, new_n8374,
    new_n8375, new_n8376_1, new_n8377, new_n8378, new_n8379, new_n8380,
    new_n8381_1, new_n8382, new_n8383, new_n8384, new_n8385, new_n8386,
    new_n8387, new_n8388, new_n8389, new_n8390, new_n8391, new_n8392,
    new_n8393, new_n8394, new_n8395, new_n8396, new_n8397, new_n8398,
    new_n8399_1, new_n8400, new_n8401, new_n8402, new_n8403, new_n8404,
    new_n8405_1, new_n8406, new_n8407, new_n8408_1, new_n8409, new_n8410,
    new_n8411, new_n8412, new_n8413, new_n8414, new_n8415, new_n8416,
    new_n8417_1, new_n8418, new_n8419, new_n8420, new_n8421, new_n8422,
    new_n8423, new_n8424, new_n8425, new_n8426, new_n8427, new_n8428,
    new_n8429, new_n8430, new_n8431, new_n8432_1, new_n8433, new_n8434,
    new_n8435, new_n8436, new_n8437, new_n8438, new_n8439_1, new_n8440,
    new_n8441, new_n8442, new_n8443, new_n8444, new_n8445, new_n8446,
    new_n8447, new_n8448, new_n8449, new_n8450, new_n8451, new_n8452,
    new_n8453_1, new_n8454, new_n8455, new_n8456, new_n8457, new_n8458,
    new_n8459, new_n8460, new_n8461, new_n8462, new_n8463, new_n8464,
    new_n8465, new_n8466, new_n8467, new_n8468, new_n8469, new_n8470,
    new_n8471, new_n8472, new_n8473, new_n8474, new_n8475, new_n8476,
    new_n8477, new_n8478, new_n8479, new_n8480_1, new_n8481, new_n8482,
    new_n8483, new_n8484, new_n8485, new_n8486, new_n8487, new_n8488,
    new_n8489_1, new_n8490, new_n8491, new_n8492, new_n8493, new_n8494,
    new_n8495, new_n8496, new_n8497, new_n8498, new_n8499, new_n8500,
    new_n8501, new_n8502, new_n8503, new_n8504, new_n8505_1, new_n8506,
    new_n8507, new_n8508, new_n8509, new_n8510_1, new_n8511, new_n8512,
    new_n8513, new_n8514, new_n8515, new_n8516, new_n8517, new_n8518,
    new_n8519_1, new_n8520, new_n8521, new_n8522, new_n8523, new_n8524,
    new_n8525, new_n8526_1, new_n8527, new_n8528, new_n8529, new_n8530,
    new_n8531, new_n8532, new_n8533, new_n8534, new_n8535_1, new_n8536,
    new_n8537, new_n8538, new_n8539, new_n8540, new_n8541, new_n8542,
    new_n8543, new_n8544, new_n8545, new_n8546, new_n8547, new_n8548,
    new_n8549, new_n8550_1, new_n8551, new_n8552, new_n8553, new_n8554,
    new_n8555, new_n8556, new_n8557, new_n8558, new_n8559, new_n8560,
    new_n8561, new_n8562, new_n8563_1, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581_1, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594_1, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608_1, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614_1, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620_1, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637_1, new_n8638_1, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656_1, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662_1, new_n8663,
    new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678_1, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687_1,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694_1, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716_1, new_n8717,
    new_n8718, new_n8719, new_n8720, new_n8721_1, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744_1, new_n8745_1, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782_1, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803_1, new_n8804, new_n8805, new_n8806_1, new_n8807, new_n8808,
    new_n8809_1, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821_1, new_n8822, new_n8823, new_n8824_1, new_n8825, new_n8826,
    new_n8827_1, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849_1, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856_1,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861_1, new_n8862_1,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869_1, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884_1, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909_1, new_n8910,
    new_n8911_1, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920_1, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943_1, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964_1,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971_1, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982_1,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993_1, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003_1, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012_1,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032_1, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042_1,
    new_n9043, new_n9044, new_n9045, new_n9046_1, new_n9047_1, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090_1,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9104_1, new_n9105, new_n9106, new_n9107, new_n9108, new_n9109,
    new_n9110, new_n9111, new_n9112, new_n9113, new_n9114, new_n9115,
    new_n9116, new_n9117, new_n9118, new_n9119, new_n9120, new_n9121,
    new_n9122, new_n9123, new_n9124, new_n9125, new_n9126, new_n9127,
    new_n9128, new_n9129_1, new_n9130, new_n9131, new_n9132, new_n9133,
    new_n9134, new_n9135, new_n9136, new_n9137, new_n9138, new_n9139,
    new_n9140, new_n9141, new_n9142, new_n9143, new_n9144, new_n9145,
    new_n9146_1, new_n9147, new_n9148, new_n9149, new_n9150, new_n9151,
    new_n9152, new_n9153, new_n9154, new_n9155, new_n9156, new_n9157,
    new_n9158, new_n9159, new_n9160, new_n9161, new_n9162, new_n9163,
    new_n9164_1, new_n9165, new_n9166_1, new_n9167, new_n9168, new_n9169,
    new_n9170, new_n9171, new_n9172_1, new_n9173, new_n9174, new_n9175,
    new_n9176, new_n9177, new_n9178, new_n9179, new_n9180, new_n9181,
    new_n9182_1, new_n9183, new_n9184, new_n9185, new_n9186, new_n9187,
    new_n9188, new_n9189, new_n9190, new_n9191_1, new_n9192, new_n9193,
    new_n9194, new_n9195, new_n9196, new_n9197, new_n9198, new_n9199,
    new_n9200, new_n9201, new_n9202, new_n9203, new_n9204, new_n9205,
    new_n9206, new_n9207, new_n9208, new_n9209, new_n9210, new_n9211,
    new_n9212, new_n9213, new_n9214, new_n9215, new_n9216, new_n9217_1,
    new_n9218, new_n9219, new_n9220_1, new_n9221, new_n9222, new_n9223,
    new_n9224, new_n9225, new_n9226, new_n9227, new_n9228, new_n9229,
    new_n9230, new_n9231, new_n9232, new_n9233, new_n9234, new_n9235,
    new_n9236, new_n9237, new_n9238, new_n9239, new_n9240, new_n9241,
    new_n9242, new_n9243, new_n9244, new_n9245, new_n9246_1, new_n9247,
    new_n9248, new_n9249, new_n9250, new_n9251_1, new_n9252, new_n9253,
    new_n9254, new_n9255, new_n9256, new_n9257, new_n9258, new_n9259_1,
    new_n9260, new_n9261_1, new_n9262, new_n9263, new_n9264, new_n9265,
    new_n9266, new_n9267, new_n9268, new_n9269, new_n9270, new_n9271,
    new_n9272, new_n9273, new_n9274, new_n9275, new_n9276, new_n9277,
    new_n9278, new_n9279, new_n9280, new_n9281, new_n9282, new_n9283,
    new_n9284, new_n9285, new_n9286, new_n9287_1, new_n9288, new_n9289,
    new_n9290, new_n9291, new_n9292, new_n9293, new_n9294, new_n9295,
    new_n9296, new_n9297, new_n9298, new_n9299, new_n9300, new_n9301,
    new_n9302, new_n9303, new_n9304, new_n9305, new_n9306, new_n9307,
    new_n9308_1, new_n9309, new_n9310, new_n9311, new_n9312, new_n9313,
    new_n9314, new_n9315, new_n9316, new_n9317, new_n9318_1, new_n9319,
    new_n9320, new_n9321, new_n9322, new_n9323_1, new_n9324, new_n9325,
    new_n9326, new_n9327, new_n9328, new_n9329, new_n9330, new_n9331,
    new_n9332, new_n9333, new_n9334, new_n9335, new_n9336, new_n9337,
    new_n9338, new_n9339, new_n9340, new_n9341, new_n9342, new_n9343,
    new_n9344_1, new_n9345, new_n9346, new_n9347, new_n9348, new_n9349,
    new_n9350, new_n9351, new_n9352, new_n9353, new_n9354, new_n9355,
    new_n9356, new_n9357, new_n9358, new_n9359, new_n9360, new_n9361,
    new_n9362, new_n9363, new_n9364_1, new_n9365, new_n9366, new_n9367,
    new_n9368, new_n9369, new_n9370, new_n9371_1, new_n9372_1, new_n9373,
    new_n9374, new_n9375, new_n9376, new_n9377, new_n9378, new_n9379,
    new_n9380_1, new_n9381, new_n9382_1, new_n9383, new_n9384, new_n9385,
    new_n9386, new_n9387, new_n9388, new_n9389, new_n9390, new_n9391,
    new_n9392, new_n9393, new_n9394, new_n9395, new_n9396_1, new_n9397,
    new_n9398, new_n9399_1, new_n9400, new_n9401, new_n9402, new_n9403_1,
    new_n9404, new_n9405, new_n9406, new_n9407, new_n9408, new_n9409,
    new_n9410, new_n9411, new_n9412, new_n9413, new_n9414, new_n9415,
    new_n9416, new_n9417, new_n9418, new_n9419_1, new_n9420, new_n9421,
    new_n9422, new_n9423_1, new_n9424, new_n9425, new_n9426, new_n9427,
    new_n9428, new_n9430_1, new_n9432, new_n9433, new_n9434, new_n9435_1,
    new_n9436, new_n9437, new_n9438, new_n9439, new_n9440, new_n9441,
    new_n9442, new_n9443, new_n9444, new_n9445_1, new_n9446, new_n9447,
    new_n9448, new_n9449, new_n9450, new_n9451_1, new_n9452, new_n9453,
    new_n9454, new_n9455, new_n9456, new_n9457, new_n9458_1, new_n9459_1,
    new_n9460_1, new_n9461, new_n9462, new_n9463, new_n9464, new_n9465,
    new_n9466, new_n9467, new_n9468, new_n9469, new_n9470, new_n9471,
    new_n9472, new_n9473, new_n9474, new_n9475, new_n9476, new_n9477,
    new_n9478, new_n9479, new_n9480, new_n9481, new_n9482, new_n9483,
    new_n9484, new_n9485, new_n9486, new_n9487, new_n9488, new_n9489,
    new_n9490, new_n9491, new_n9492, new_n9493_1, new_n9494, new_n9495,
    new_n9496, new_n9497, new_n9498, new_n9499, new_n9500, new_n9501,
    new_n9502, new_n9503, new_n9504, new_n9505, new_n9506, new_n9507_1,
    new_n9508_1, new_n9509, new_n9510, new_n9511, new_n9512_1, new_n9513,
    new_n9514, new_n9515, new_n9516, new_n9517, new_n9518, new_n9519,
    new_n9520, new_n9521, new_n9522, new_n9523, new_n9524, new_n9525,
    new_n9526, new_n9527, new_n9528, new_n9529, new_n9530, new_n9531,
    new_n9532, new_n9533, new_n9534, new_n9535, new_n9536, new_n9537,
    new_n9538, new_n9539, new_n9540, new_n9541, new_n9542, new_n9543,
    new_n9544, new_n9545, new_n9546, new_n9547, new_n9548, new_n9549,
    new_n9550, new_n9551, new_n9552_1, new_n9553, new_n9554_1, new_n9555,
    new_n9556_1, new_n9557_1, new_n9558_1, new_n9559, new_n9560, new_n9561,
    new_n9562, new_n9563, new_n9564, new_n9565, new_n9566, new_n9567,
    new_n9568, new_n9569, new_n9570, new_n9571, new_n9572, new_n9573,
    new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579,
    new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585,
    new_n9586, new_n9587, new_n9588, new_n9589, new_n9590, new_n9591,
    new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597,
    new_n9598_1, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603,
    new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609,
    new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615,
    new_n9616_1, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621,
    new_n9622_1, new_n9623, new_n9624, new_n9625, new_n9626_1, new_n9627,
    new_n9628, new_n9629, new_n9631, new_n9632, new_n9633_1, new_n9634,
    new_n9635_1, new_n9636, new_n9637, new_n9638, new_n9639, new_n9640,
    new_n9641, new_n9642, new_n9643, new_n9644, new_n9645, new_n9646_1,
    new_n9647, new_n9648_1, new_n9649, new_n9650, new_n9651, new_n9652,
    new_n9653, new_n9654, new_n9655_1, new_n9656, new_n9657, new_n9658,
    new_n9659, new_n9660, new_n9661, new_n9662, new_n9663, new_n9664,
    new_n9665, new_n9666, new_n9667, new_n9668, new_n9669, new_n9670,
    new_n9671, new_n9672, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689_1,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695_1,
    new_n9696, new_n9697, new_n9698, new_n9699_1, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725,
    new_n9726_1, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753_1, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761_1, new_n9762,
    new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1, new_n9768,
    new_n9769, new_n9770, new_n9771_1, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778_1, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783_1, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803_1, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832_1, new_n9833_1, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838_1, new_n9839, new_n9840,
    new_n9841, new_n9843, new_n9844, new_n9845, new_n9846, new_n9847,
    new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865,
    new_n9866, new_n9867_1, new_n9868, new_n9869, new_n9870, new_n9871,
    new_n9872_1, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877,
    new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883,
    new_n9884, new_n9885, new_n9886, new_n9887, new_n9888, new_n9889,
    new_n9890_1, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895,
    new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901,
    new_n9902, new_n9903, new_n9904, new_n9905, new_n9906, new_n9907,
    new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915, new_n9916, new_n9917_1, new_n9918, new_n9919_1,
    new_n9920, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926_1, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934_1, new_n9935, new_n9936, new_n9937,
    new_n9938_1, new_n9939, new_n9940, new_n9941, new_n9943, new_n9944,
    new_n9945, new_n9946_1, new_n9947, new_n9948, new_n9949, new_n9950,
    new_n9951, new_n9952, new_n9953, new_n9954, new_n9955, new_n9956,
    new_n9957, new_n9958, new_n9959, new_n9960, new_n9961, new_n9962,
    new_n9963, new_n9964, new_n9965, new_n9966, new_n9967_1, new_n9968_1,
    new_n9969, new_n9970, new_n9971, new_n9972, new_n9973, new_n9974,
    new_n9975, new_n9976, new_n9977, new_n9978, new_n9979, new_n9980,
    new_n9981, new_n9982, new_n9983, new_n9984, new_n9985, new_n9986,
    new_n9987, new_n9988, new_n9989, new_n9990, new_n9991, new_n9992,
    new_n9993, new_n9994, new_n9995, new_n9996, new_n9997, new_n9998,
    new_n9999, new_n10000, new_n10001, new_n10002, new_n10003, new_n10004,
    new_n10005, new_n10006, new_n10007, new_n10008, new_n10009_1,
    new_n10010_1, new_n10011, new_n10012, new_n10013, new_n10014,
    new_n10015, new_n10016, new_n10017_1, new_n10018_1, new_n10019_1,
    new_n10020, new_n10021_1, new_n10022, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053_1,
    new_n10054, new_n10055_1, new_n10056, new_n10057_1, new_n10058,
    new_n10059, new_n10060, new_n10061, new_n10062, new_n10063, new_n10064,
    new_n10065, new_n10066, new_n10067, new_n10068, new_n10069, new_n10070,
    new_n10071, new_n10072, new_n10073, new_n10074, new_n10075, new_n10076,
    new_n10077, new_n10078, new_n10079, new_n10080, new_n10081, new_n10082,
    new_n10083, new_n10084, new_n10085, new_n10086, new_n10087, new_n10088,
    new_n10089, new_n10090, new_n10091, new_n10092, new_n10093, new_n10094,
    new_n10095, new_n10096_1, new_n10097, new_n10098, new_n10099,
    new_n10100, new_n10101_1, new_n10102, new_n10103, new_n10104,
    new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111_1, new_n10112, new_n10113, new_n10114, new_n10115,
    new_n10116, new_n10117_1, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125_1,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10133, new_n10134, new_n10135, new_n10136, new_n10137,
    new_n10138, new_n10139, new_n10140, new_n10141, new_n10142, new_n10143,
    new_n10144, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158_1, new_n10159, new_n10160,
    new_n10161, new_n10162, new_n10163, new_n10164, new_n10165_1,
    new_n10166, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171,
    new_n10172, new_n10173, new_n10174, new_n10175, new_n10176, new_n10177,
    new_n10178, new_n10179, new_n10180, new_n10181, new_n10182, new_n10183,
    new_n10184, new_n10185, new_n10186, new_n10187, new_n10188, new_n10189,
    new_n10190, new_n10191, new_n10192, new_n10193, new_n10194, new_n10195,
    new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201_1, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223,
    new_n10224, new_n10225, new_n10226, new_n10227, new_n10228, new_n10229,
    new_n10230, new_n10231, new_n10232, new_n10233, new_n10234, new_n10235,
    new_n10236_1, new_n10237, new_n10238, new_n10239_1, new_n10240,
    new_n10241, new_n10242, new_n10243, new_n10244_1, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250_1,
    new_n10251, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261_1, new_n10262_1,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275_1, new_n10276, new_n10277, new_n10278, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285,
    new_n10286, new_n10287_1, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295_1,
    new_n10296, new_n10297, new_n10298, new_n10299, new_n10300, new_n10301,
    new_n10302, new_n10303, new_n10304, new_n10305, new_n10306, new_n10307,
    new_n10308, new_n10309, new_n10310, new_n10311, new_n10312, new_n10313,
    new_n10314, new_n10315, new_n10316, new_n10317, new_n10318, new_n10319,
    new_n10320, new_n10321_1, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326_1, new_n10327_1, new_n10328, new_n10329,
    new_n10330_1, new_n10331, new_n10332, new_n10333, new_n10334,
    new_n10335, new_n10336, new_n10337, new_n10338, new_n10339,
    new_n10340_1, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345_1, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356_1, new_n10357, new_n10358, new_n10359, new_n10360,
    new_n10361, new_n10362, new_n10363, new_n10364, new_n10365, new_n10366,
    new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372_1, new_n10373, new_n10374, new_n10375, new_n10376,
    new_n10377, new_n10378, new_n10379, new_n10380, new_n10381, new_n10382,
    new_n10383, new_n10384, new_n10385_1, new_n10386, new_n10387_1,
    new_n10388_1, new_n10389, new_n10390_1, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404_1, new_n10405_1, new_n10406, new_n10407, new_n10408,
    new_n10409_1, new_n10410, new_n10411_1, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420_1, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432_1, new_n10433, new_n10434, new_n10435,
    new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10454,
    new_n10455, new_n10456, new_n10457, new_n10458, new_n10459, new_n10460,
    new_n10461, new_n10462, new_n10463, new_n10464, new_n10465, new_n10466,
    new_n10467, new_n10468, new_n10469, new_n10470, new_n10471, new_n10472,
    new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483,
    new_n10484_1, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489_1, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10504, new_n10505,
    new_n10506, new_n10507, new_n10508, new_n10509, new_n10510, new_n10511,
    new_n10512, new_n10513, new_n10514_1, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525_1, new_n10526, new_n10527,
    new_n10528, new_n10529, new_n10530, new_n10531, new_n10532, new_n10533,
    new_n10534, new_n10535, new_n10536, new_n10537, new_n10538, new_n10539,
    new_n10540_1, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561_1,
    new_n10562, new_n10563, new_n10564_1, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577_1,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588_1,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593_1,
    new_n10594, new_n10595_1, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611_1, new_n10612, new_n10613, new_n10614_1, new_n10615,
    new_n10616, new_n10617_1, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628_1, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647_1, new_n10649,
    new_n10651, new_n10653_1, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692_1,
    new_n10693, new_n10694_1, new_n10695, new_n10696, new_n10697,
    new_n10698, new_n10699, new_n10700, new_n10701_1, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710_1, new_n10711, new_n10712_1, new_n10713,
    new_n10714, new_n10715, new_n10716, new_n10717, new_n10718, new_n10719,
    new_n10720, new_n10721, new_n10722, new_n10723, new_n10724, new_n10725,
    new_n10726, new_n10727, new_n10728, new_n10729, new_n10730, new_n10731,
    new_n10732, new_n10733, new_n10734, new_n10735, new_n10736, new_n10737,
    new_n10738, new_n10739_1, new_n10740, new_n10741, new_n10742,
    new_n10743, new_n10744, new_n10745, new_n10746, new_n10747, new_n10748,
    new_n10749, new_n10750, new_n10751, new_n10752, new_n10753, new_n10754,
    new_n10755, new_n10756_1, new_n10757, new_n10758, new_n10759,
    new_n10760, new_n10761, new_n10762, new_n10763_1, new_n10764,
    new_n10765, new_n10766, new_n10767, new_n10768, new_n10769, new_n10770,
    new_n10771, new_n10772, new_n10773, new_n10774, new_n10775_1,
    new_n10776, new_n10777, new_n10778, new_n10779, new_n10780_1,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791,
    new_n10792_1, new_n10793, new_n10794, new_n10795, new_n10796,
    new_n10797, new_n10798, new_n10799, new_n10800, new_n10801, new_n10802,
    new_n10803, new_n10804, new_n10805, new_n10806, new_n10807, new_n10808,
    new_n10809, new_n10810, new_n10811, new_n10812, new_n10813, new_n10814,
    new_n10815, new_n10816, new_n10817_1, new_n10818, new_n10819,
    new_n10820, new_n10821, new_n10822, new_n10823, new_n10824, new_n10825,
    new_n10826, new_n10827, new_n10828, new_n10829, new_n10830, new_n10831,
    new_n10832, new_n10833, new_n10834_1, new_n10835, new_n10836,
    new_n10837, new_n10838, new_n10839, new_n10840, new_n10841, new_n10842,
    new_n10843, new_n10844, new_n10845, new_n10846, new_n10847, new_n10848,
    new_n10849, new_n10850, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874_1, new_n10875, new_n10876, new_n10877, new_n10878,
    new_n10879, new_n10880, new_n10881, new_n10882, new_n10883, new_n10884,
    new_n10885, new_n10886, new_n10887, new_n10888, new_n10889, new_n10890,
    new_n10891, new_n10892, new_n10893, new_n10894, new_n10895, new_n10896,
    new_n10897, new_n10898, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913, new_n10914,
    new_n10915, new_n10916, new_n10917, new_n10918, new_n10919, new_n10920,
    new_n10921, new_n10922, new_n10923, new_n10924_1, new_n10925,
    new_n10926, new_n10927, new_n10928, new_n10929, new_n10930, new_n10931,
    new_n10932, new_n10933, new_n10934, new_n10935, new_n10936, new_n10937,
    new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943_1, new_n10944, new_n10945, new_n10946, new_n10947,
    new_n10948, new_n10949, new_n10950, new_n10951, new_n10952, new_n10953,
    new_n10954, new_n10955, new_n10956, new_n10957, new_n10958, new_n10959,
    new_n10960, new_n10961_1, new_n10962, new_n10963, new_n10964,
    new_n10965, new_n10967, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990,
    new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996,
    new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002,
    new_n11003, new_n11004, new_n11005_1, new_n11006, new_n11007,
    new_n11008, new_n11009, new_n11010, new_n11011_1, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023_1,
    new_n11024, new_n11025_1, new_n11026, new_n11027, new_n11028,
    new_n11029, new_n11030, new_n11031, new_n11032, new_n11033, new_n11034,
    new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040,
    new_n11041, new_n11042, new_n11043, new_n11044_1, new_n11045,
    new_n11046, new_n11047, new_n11048, new_n11049, new_n11050, new_n11051,
    new_n11052, new_n11053, new_n11054, new_n11055, new_n11056_1,
    new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062,
    new_n11063_1, new_n11064, new_n11065, new_n11066, new_n11067,
    new_n11068, new_n11069, new_n11070, new_n11071, new_n11072, new_n11073,
    new_n11074, new_n11075, new_n11076, new_n11077, new_n11078_1,
    new_n11079, new_n11080_1, new_n11081, new_n11082, new_n11083,
    new_n11084, new_n11085, new_n11086, new_n11087, new_n11088, new_n11090,
    new_n11091, new_n11092, new_n11093, new_n11094_1, new_n11095,
    new_n11096, new_n11097, new_n11098, new_n11099, new_n11100,
    new_n11101_1, new_n11102, new_n11103_1, new_n11104, new_n11105,
    new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111,
    new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117,
    new_n11118, new_n11119, new_n11120_1, new_n11121_1, new_n11122,
    new_n11123, new_n11124, new_n11125, new_n11126, new_n11127_1,
    new_n11128, new_n11129, new_n11130, new_n11131, new_n11132_1,
    new_n11133, new_n11134_1, new_n11135, new_n11136, new_n11137,
    new_n11138_1, new_n11139, new_n11140, new_n11141, new_n11142,
    new_n11143, new_n11144, new_n11145, new_n11146, new_n11147, new_n11148,
    new_n11149, new_n11150, new_n11151, new_n11152, new_n11153, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178,
    new_n11179, new_n11180, new_n11181, new_n11182_1, new_n11183,
    new_n11184_1, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192_1, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201_1, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220_1, new_n11221,
    new_n11222, new_n11223_1, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234_1, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245_1, new_n11246, new_n11247, new_n11249,
    new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257, new_n11258, new_n11259, new_n11260, new_n11261_1,
    new_n11262, new_n11264, new_n11265, new_n11266_1, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272,
    new_n11273_1, new_n11274, new_n11275_1, new_n11276, new_n11277,
    new_n11278, new_n11279, new_n11280, new_n11281, new_n11282, new_n11283,
    new_n11284, new_n11285, new_n11286, new_n11288, new_n11289, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296, new_n11297,
    new_n11298, new_n11299, new_n11300, new_n11301, new_n11302_1,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311, new_n11312, new_n11313_1,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324,
    new_n11325_1, new_n11326_1, new_n11327, new_n11328, new_n11329,
    new_n11330_1, new_n11331, new_n11332, new_n11333, new_n11334,
    new_n11335, new_n11336, new_n11337, new_n11338, new_n11339, new_n11340,
    new_n11341, new_n11342, new_n11343, new_n11344, new_n11345, new_n11346,
    new_n11347_1, new_n11348_1, new_n11349, new_n11350, new_n11351,
    new_n11352_1, new_n11353, new_n11354, new_n11355, new_n11356_1,
    new_n11357, new_n11358, new_n11359, new_n11360, new_n11361, new_n11362,
    new_n11363, new_n11364, new_n11365, new_n11366, new_n11367, new_n11368,
    new_n11369, new_n11370, new_n11371, new_n11372, new_n11373, new_n11374,
    new_n11375_1, new_n11376, new_n11377, new_n11378, new_n11379_1,
    new_n11380, new_n11381, new_n11382, new_n11383, new_n11384, new_n11385,
    new_n11386_1, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391_1, new_n11392, new_n11393, new_n11394, new_n11395,
    new_n11396, new_n11397, new_n11398_1, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403_1, new_n11404, new_n11405,
    new_n11406, new_n11407, new_n11408, new_n11409, new_n11410, new_n11411,
    new_n11412, new_n11413, new_n11414, new_n11415, new_n11416, new_n11417,
    new_n11418, new_n11419_1, new_n11420, new_n11421, new_n11422,
    new_n11423, new_n11424_1, new_n11425, new_n11426, new_n11427,
    new_n11428, new_n11429, new_n11430, new_n11431, new_n11432, new_n11433,
    new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439_1, new_n11440, new_n11441, new_n11442, new_n11443,
    new_n11444, new_n11445, new_n11446, new_n11447, new_n11448, new_n11449,
    new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455_1, new_n11456, new_n11457, new_n11458, new_n11459,
    new_n11460, new_n11461, new_n11462_1, new_n11463, new_n11464,
    new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470_1, new_n11471, new_n11472_1, new_n11473_1, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479_1,
    new_n11480, new_n11481_1, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486_1, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496_1, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503_1, new_n11504, new_n11505,
    new_n11506_1, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515_1,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536, new_n11537, new_n11538_1,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548_1, new_n11549,
    new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555,
    new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561,
    new_n11562, new_n11563, new_n11564_1, new_n11565, new_n11566_1,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579_1, new_n11580_1, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11587, new_n11588, new_n11589,
    new_n11590, new_n11591_1, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607_1, new_n11608, new_n11609, new_n11610, new_n11611,
    new_n11612, new_n11613, new_n11614, new_n11615_1, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11623,
    new_n11624, new_n11625, new_n11626, new_n11627, new_n11628, new_n11629,
    new_n11630_1, new_n11631, new_n11632, new_n11633, new_n11634,
    new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640,
    new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647_1, new_n11648, new_n11649, new_n11650, new_n11651,
    new_n11652, new_n11653, new_n11654, new_n11655, new_n11656, new_n11657,
    new_n11658, new_n11659, new_n11660, new_n11661, new_n11662, new_n11663,
    new_n11664, new_n11665, new_n11666, new_n11667_1, new_n11668,
    new_n11669, new_n11670, new_n11671, new_n11672, new_n11673,
    new_n11674_1, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682_1, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706, new_n11707,
    new_n11708, new_n11709, new_n11710_1, new_n11711, new_n11712_1,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724_1, new_n11725, new_n11726, new_n11727, new_n11728,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736_1, new_n11737, new_n11738, new_n11739,
    new_n11740, new_n11741_1, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749_1,
    new_n11750, new_n11751, new_n11752, new_n11753, new_n11754, new_n11755,
    new_n11756, new_n11757, new_n11758, new_n11759, new_n11760, new_n11761,
    new_n11762, new_n11763, new_n11764, new_n11765, new_n11766, new_n11767,
    new_n11768, new_n11769, new_n11770_1, new_n11771_1, new_n11772,
    new_n11773, new_n11774, new_n11775_1, new_n11776, new_n11777,
    new_n11778, new_n11779, new_n11780, new_n11781, new_n11782, new_n11783,
    new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789,
    new_n11790, new_n11791, new_n11792, new_n11793, new_n11794, new_n11795,
    new_n11796, new_n11797, new_n11798, new_n11799, new_n11800, new_n11801,
    new_n11802, new_n11803, new_n11804, new_n11805, new_n11806, new_n11807,
    new_n11808, new_n11809, new_n11810, new_n11811, new_n11812, new_n11813,
    new_n11814, new_n11815, new_n11816, new_n11817, new_n11818_1,
    new_n11819, new_n11820, new_n11821, new_n11822, new_n11823, new_n11824,
    new_n11825, new_n11826, new_n11827, new_n11828, new_n11829, new_n11830,
    new_n11831, new_n11832, new_n11833, new_n11834, new_n11836,
    new_n11837_1, new_n11838, new_n11839, new_n11840, new_n11841_1,
    new_n11842_1, new_n11843_1, new_n11844, new_n11845, new_n11846,
    new_n11847, new_n11848, new_n11849, new_n11850, new_n11851, new_n11852,
    new_n11853, new_n11854, new_n11855, new_n11856, new_n11857, new_n11858,
    new_n11859, new_n11860, new_n11861, new_n11862, new_n11863, new_n11864,
    new_n11865, new_n11866, new_n11867, new_n11868, new_n11869, new_n11870,
    new_n11871, new_n11872, new_n11873, new_n11874, new_n11875, new_n11876,
    new_n11877, new_n11878, new_n11879, new_n11880, new_n11881, new_n11882,
    new_n11883, new_n11884, new_n11885, new_n11886, new_n11887, new_n11888,
    new_n11889, new_n11890, new_n11891, new_n11892, new_n11893, new_n11894,
    new_n11895, new_n11896, new_n11897, new_n11898_1, new_n11899,
    new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905_1, new_n11906, new_n11907, new_n11908, new_n11909,
    new_n11910, new_n11911, new_n11912, new_n11913, new_n11914, new_n11915,
    new_n11916, new_n11917, new_n11918, new_n11919, new_n11920, new_n11921,
    new_n11922, new_n11923, new_n11924, new_n11925, new_n11926_1,
    new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932,
    new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938,
    new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944,
    new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950,
    new_n11951, new_n11952, new_n11953, new_n11954, new_n11955, new_n11956,
    new_n11957, new_n11958, new_n11959, new_n11960, new_n11961, new_n11962,
    new_n11963, new_n11964, new_n11965_1, new_n11966, new_n11967,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980_1, new_n11981, new_n11982, new_n11983, new_n11984,
    new_n11985, new_n11986, new_n11987, new_n11988, new_n11989, new_n11990,
    new_n11991, new_n11992, new_n11993, new_n11994, new_n11995, new_n11996,
    new_n11997, new_n11998, new_n11999, new_n12000_1, new_n12001,
    new_n12002, new_n12003_1, new_n12004, new_n12005, new_n12006,
    new_n12007, new_n12008, new_n12009, new_n12010, new_n12011_1,
    new_n12012, new_n12013, new_n12014, new_n12015, new_n12016, new_n12017,
    new_n12018, new_n12019, new_n12020, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044, new_n12045, new_n12046, new_n12047,
    new_n12048, new_n12049, new_n12050, new_n12051, new_n12052, new_n12053,
    new_n12054, new_n12055, new_n12056, new_n12057, new_n12058, new_n12059,
    new_n12060, new_n12061, new_n12062, new_n12063, new_n12064, new_n12065,
    new_n12066, new_n12067, new_n12068, new_n12069, new_n12070, new_n12071,
    new_n12072_1, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12109, new_n12110, new_n12111, new_n12112,
    new_n12113_1, new_n12114, new_n12115, new_n12116, new_n12117,
    new_n12118, new_n12119, new_n12120, new_n12121_1, new_n12122,
    new_n12123, new_n12124, new_n12125, new_n12126, new_n12127, new_n12128,
    new_n12129, new_n12130, new_n12131_1, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144, new_n12145,
    new_n12146_1, new_n12147, new_n12148, new_n12149, new_n12150,
    new_n12151, new_n12152_1, new_n12153_1, new_n12154, new_n12155,
    new_n12156, new_n12157_1, new_n12158_1, new_n12159, new_n12160,
    new_n12161_1, new_n12162, new_n12163, new_n12164, new_n12165,
    new_n12166, new_n12167, new_n12168, new_n12169, new_n12170, new_n12171,
    new_n12172, new_n12173, new_n12174, new_n12175, new_n12176, new_n12177,
    new_n12178, new_n12179_1, new_n12180, new_n12181, new_n12182,
    new_n12183, new_n12184, new_n12185, new_n12186, new_n12187, new_n12188,
    new_n12189, new_n12190, new_n12191, new_n12192_1, new_n12193,
    new_n12194, new_n12195, new_n12196, new_n12197, new_n12198, new_n12199,
    new_n12200, new_n12201, new_n12202, new_n12203, new_n12204, new_n12205,
    new_n12206, new_n12207, new_n12208, new_n12209_1, new_n12210,
    new_n12211, new_n12212, new_n12213, new_n12215, new_n12216, new_n12217,
    new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223_1, new_n12224, new_n12225_1, new_n12226, new_n12227,
    new_n12228_1, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235_1, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247, new_n12248, new_n12249,
    new_n12250, new_n12251, new_n12252, new_n12253, new_n12254, new_n12255,
    new_n12256, new_n12257, new_n12258, new_n12259, new_n12260, new_n12261,
    new_n12262, new_n12263, new_n12264, new_n12265, new_n12266, new_n12267,
    new_n12268, new_n12269, new_n12270, new_n12271, new_n12272, new_n12273,
    new_n12274, new_n12275, new_n12276, new_n12277, new_n12278, new_n12279,
    new_n12280, new_n12281, new_n12282, new_n12283, new_n12284, new_n12285,
    new_n12286, new_n12287, new_n12288, new_n12289, new_n12290, new_n12291,
    new_n12292, new_n12293, new_n12294, new_n12295, new_n12296, new_n12297,
    new_n12298, new_n12299, new_n12300, new_n12301, new_n12302_1,
    new_n12303, new_n12304_1, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315_1, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12322, new_n12323,
    new_n12324_1, new_n12325_1, new_n12326, new_n12327, new_n12328,
    new_n12329_1, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341_1, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346_1, new_n12347, new_n12348, new_n12349_1, new_n12350,
    new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364_1, new_n12365, new_n12366, new_n12367,
    new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373,
    new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380_1, new_n12381, new_n12382, new_n12383_1, new_n12384_1,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397_1, new_n12398_1, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408_1, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446_1, new_n12447,
    new_n12448, new_n12449_1, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461_1, new_n12462_1, new_n12463,
    new_n12464, new_n12465, new_n12466, new_n12467_1, new_n12468,
    new_n12469_1, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495_1, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507_1,
    new_n12508, new_n12509, new_n12510, new_n12511, new_n12512, new_n12513,
    new_n12514, new_n12515_1, new_n12516_1, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12525,
    new_n12526, new_n12527, new_n12528, new_n12529, new_n12530, new_n12531,
    new_n12532, new_n12533, new_n12534, new_n12535, new_n12537, new_n12538,
    new_n12539, new_n12540_1, new_n12541, new_n12542, new_n12543,
    new_n12544, new_n12545_1, new_n12546_1, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552_1, new_n12553,
    new_n12554, new_n12555, new_n12556, new_n12557, new_n12558, new_n12559,
    new_n12560, new_n12561, new_n12562_1, new_n12563, new_n12564,
    new_n12565, new_n12566_1, new_n12567, new_n12568, new_n12569_1,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587_1, new_n12588, new_n12589, new_n12590, new_n12591,
    new_n12592, new_n12593_1, new_n12594, new_n12595, new_n12596,
    new_n12597, new_n12598, new_n12599, new_n12600, new_n12601, new_n12602,
    new_n12603, new_n12604, new_n12605, new_n12606, new_n12607_1,
    new_n12608, new_n12609, new_n12610, new_n12611, new_n12612, new_n12613,
    new_n12614, new_n12615, new_n12616, new_n12617, new_n12618, new_n12619,
    new_n12620_1, new_n12621_1, new_n12622, new_n12623, new_n12624,
    new_n12625, new_n12626_1, new_n12627, new_n12628, new_n12629,
    new_n12630, new_n12631, new_n12632, new_n12633, new_n12634, new_n12635,
    new_n12636, new_n12637, new_n12638, new_n12639, new_n12640, new_n12641,
    new_n12642, new_n12643, new_n12644, new_n12645, new_n12646, new_n12647,
    new_n12648, new_n12649, new_n12650_1, new_n12651, new_n12653,
    new_n12654_1, new_n12655, new_n12656, new_n12657_1, new_n12658,
    new_n12659, new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665_1, new_n12666, new_n12667, new_n12668, new_n12669,
    new_n12670_1, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12699, new_n12700, new_n12701, new_n12702_1, new_n12703,
    new_n12704, new_n12705, new_n12706, new_n12707_1, new_n12708,
    new_n12709, new_n12710, new_n12711, new_n12712, new_n12713, new_n12714,
    new_n12715, new_n12716, new_n12717, new_n12718, new_n12719, new_n12720,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725_1,
    new_n12726, new_n12727_1, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12740_1, new_n12741,
    new_n12742_1, new_n12743, new_n12744, new_n12745, new_n12746_1,
    new_n12747, new_n12748, new_n12749, new_n12750, new_n12751, new_n12752,
    new_n12753, new_n12754, new_n12755, new_n12756_1, new_n12757,
    new_n12758, new_n12759, new_n12760, new_n12761, new_n12762, new_n12763,
    new_n12764, new_n12765, new_n12766, new_n12767, new_n12768, new_n12769,
    new_n12770, new_n12771, new_n12772, new_n12773, new_n12774, new_n12775,
    new_n12776, new_n12777, new_n12778, new_n12779, new_n12780, new_n12781,
    new_n12782, new_n12783_1, new_n12784, new_n12785, new_n12786,
    new_n12787, new_n12788, new_n12789, new_n12790, new_n12791, new_n12792,
    new_n12793, new_n12794, new_n12795, new_n12796, new_n12797, new_n12798,
    new_n12799, new_n12800, new_n12801_1, new_n12802, new_n12803,
    new_n12804, new_n12805, new_n12806, new_n12807, new_n12808, new_n12809,
    new_n12810, new_n12811_1, new_n12812_1, new_n12813, new_n12814,
    new_n12815, new_n12816_1, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821_1, new_n12822, new_n12823, new_n12824,
    new_n12825, new_n12826, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843_1, new_n12844, new_n12845, new_n12846, new_n12847,
    new_n12848, new_n12849, new_n12850, new_n12851, new_n12852, new_n12853,
    new_n12854, new_n12855, new_n12856, new_n12857, new_n12858, new_n12859,
    new_n12860, new_n12861_1, new_n12862, new_n12863, new_n12864_1,
    new_n12865_1, new_n12866, new_n12867, new_n12868, new_n12869,
    new_n12870_1, new_n12871_1, new_n12872, new_n12873_1, new_n12874,
    new_n12875_1, new_n12876, new_n12877, new_n12878, new_n12879,
    new_n12880, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12893, new_n12894, new_n12895, new_n12896, new_n12897, new_n12898,
    new_n12899, new_n12900_1, new_n12901, new_n12902, new_n12903,
    new_n12904_1, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917_1, new_n12918, new_n12919,
    new_n12920, new_n12921, new_n12922, new_n12923, new_n12924, new_n12925,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941_1, new_n12942_1,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956_1, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12973,
    new_n12974, new_n12975, new_n12976, new_n12977, new_n12978_1,
    new_n12979, new_n12980_1, new_n12981, new_n12982, new_n12983,
    new_n12984, new_n12985_1, new_n12986, new_n12987_1, new_n12988,
    new_n12989, new_n12990, new_n12991, new_n12992_1, new_n12993,
    new_n12994, new_n12995, new_n12996, new_n12997, new_n12998, new_n12999,
    new_n13000, new_n13001, new_n13002, new_n13003, new_n13004,
    new_n13005_1, new_n13006, new_n13007, new_n13008, new_n13009,
    new_n13010, new_n13011, new_n13012, new_n13013, new_n13014, new_n13015,
    new_n13016, new_n13017, new_n13018, new_n13019, new_n13020, new_n13021,
    new_n13022, new_n13023, new_n13024, new_n13025, new_n13026_1,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043_1,
    new_n13044_1, new_n13045, new_n13046, new_n13047, new_n13048_1,
    new_n13049, new_n13050, new_n13051, new_n13052, new_n13053,
    new_n13054_1, new_n13055, new_n13056, new_n13057, new_n13058,
    new_n13059, new_n13060, new_n13061, new_n13062, new_n13063, new_n13064,
    new_n13065, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070,
    new_n13071, new_n13072, new_n13073, new_n13074_1, new_n13075,
    new_n13076, new_n13077, new_n13078, new_n13079, new_n13080, new_n13081,
    new_n13082_1, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096_1, new_n13097,
    new_n13098, new_n13099, new_n13100, new_n13101, new_n13102, new_n13103,
    new_n13104, new_n13105, new_n13106, new_n13107, new_n13108, new_n13109,
    new_n13110_1, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116_1, new_n13117, new_n13118, new_n13119,
    new_n13120, new_n13121, new_n13123, new_n13125, new_n13127, new_n13129,
    new_n13130, new_n13131, new_n13132, new_n13133, new_n13134, new_n13135,
    new_n13136, new_n13137_1, new_n13138, new_n13139, new_n13140,
    new_n13141_1, new_n13142, new_n13143, new_n13144_1, new_n13145,
    new_n13146, new_n13147, new_n13148, new_n13149, new_n13150, new_n13151,
    new_n13152, new_n13153, new_n13154, new_n13155, new_n13156, new_n13157,
    new_n13158, new_n13159, new_n13160, new_n13161, new_n13162, new_n13163,
    new_n13164, new_n13165, new_n13166, new_n13167, new_n13168_1,
    new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174,
    new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180,
    new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13186,
    new_n13187, new_n13188, new_n13189, new_n13190_1, new_n13191,
    new_n13192, new_n13193, new_n13194, new_n13195, new_n13196, new_n13197,
    new_n13198_1, new_n13199_1, new_n13200, new_n13201, new_n13202,
    new_n13203, new_n13204_1, new_n13205, new_n13206, new_n13207,
    new_n13208, new_n13209_1, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263_1, new_n13264, new_n13265,
    new_n13266, new_n13267, new_n13268, new_n13269, new_n13270_1,
    new_n13271, new_n13272, new_n13273_1, new_n13274, new_n13275,
    new_n13276, new_n13277, new_n13278, new_n13279, new_n13280, new_n13281,
    new_n13282, new_n13284, new_n13285_1, new_n13286, new_n13287,
    new_n13288, new_n13289, new_n13290, new_n13291, new_n13292, new_n13293,
    new_n13294, new_n13295, new_n13296, new_n13297, new_n13298, new_n13299,
    new_n13300, new_n13301, new_n13302, new_n13303, new_n13304, new_n13305,
    new_n13306, new_n13307, new_n13308, new_n13309, new_n13310, new_n13311,
    new_n13312, new_n13313, new_n13314, new_n13315, new_n13316, new_n13317,
    new_n13318, new_n13319_1, new_n13320, new_n13321, new_n13322,
    new_n13323, new_n13324, new_n13325, new_n13326, new_n13327, new_n13328,
    new_n13329, new_n13330, new_n13331, new_n13332, new_n13333_1,
    new_n13334, new_n13335, new_n13336, new_n13337, new_n13338_1,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367_1,
    new_n13368, new_n13369, new_n13370, new_n13371, new_n13372, new_n13373,
    new_n13374, new_n13375, new_n13376, new_n13377, new_n13378, new_n13379,
    new_n13380, new_n13381, new_n13382, new_n13383, new_n13384, new_n13385,
    new_n13386, new_n13387, new_n13388, new_n13389, new_n13390, new_n13391,
    new_n13392, new_n13393, new_n13394, new_n13395, new_n13396, new_n13397,
    new_n13398, new_n13399, new_n13400, new_n13401, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407_1, new_n13408,
    new_n13409_1, new_n13410, new_n13411, new_n13412, new_n13413,
    new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419_1, new_n13420, new_n13421, new_n13422, new_n13423,
    new_n13424_1, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453_1, new_n13454, new_n13455, new_n13456_1, new_n13457_1,
    new_n13458, new_n13459, new_n13460_1, new_n13461, new_n13462,
    new_n13463, new_n13464, new_n13465, new_n13466, new_n13467, new_n13468,
    new_n13469, new_n13470, new_n13471, new_n13472, new_n13473, new_n13474,
    new_n13475, new_n13476, new_n13477_1, new_n13478, new_n13479,
    new_n13480, new_n13481, new_n13482, new_n13483, new_n13484_1,
    new_n13485, new_n13486_1, new_n13487_1, new_n13488, new_n13489,
    new_n13490_1, new_n13491, new_n13492, new_n13493, new_n13494_1,
    new_n13496, new_n13498, new_n13500_1, new_n13501_1, new_n13502,
    new_n13503, new_n13504, new_n13505, new_n13506_1, new_n13507,
    new_n13508, new_n13510, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13532, new_n13533, new_n13534,
    new_n13535, new_n13537, new_n13539, new_n13540, new_n13541, new_n13542,
    new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548_1, new_n13549_1, new_n13550, new_n13551_1, new_n13552,
    new_n13553, new_n13554, new_n13555, new_n13556, new_n13557, new_n13558,
    new_n13559, new_n13560, new_n13561, new_n13562, new_n13563, new_n13564,
    new_n13565, new_n13566, new_n13567, new_n13568, new_n13569, new_n13570,
    new_n13571, new_n13572, new_n13573, new_n13574, new_n13575, new_n13576,
    new_n13577, new_n13578, new_n13579, new_n13580, new_n13581, new_n13582,
    new_n13583, new_n13584, new_n13585, new_n13586, new_n13587, new_n13588,
    new_n13589, new_n13590, new_n13591, new_n13592, new_n13593, new_n13594,
    new_n13595, new_n13596, new_n13597, new_n13598, new_n13599, new_n13600,
    new_n13601, new_n13602_1, new_n13603, new_n13604, new_n13605,
    new_n13606, new_n13607, new_n13608, new_n13609, new_n13610, new_n13611,
    new_n13612, new_n13613, new_n13614, new_n13615, new_n13616, new_n13617,
    new_n13618, new_n13619, new_n13620, new_n13621, new_n13622, new_n13623,
    new_n13624, new_n13625, new_n13626_1, new_n13627, new_n13628,
    new_n13629, new_n13630, new_n13631, new_n13632, new_n13633, new_n13634,
    new_n13635, new_n13636, new_n13637, new_n13638, new_n13639, new_n13640,
    new_n13641, new_n13642, new_n13643, new_n13644, new_n13645, new_n13646,
    new_n13647, new_n13648, new_n13649, new_n13650, new_n13651, new_n13652,
    new_n13653, new_n13654, new_n13655, new_n13656, new_n13657, new_n13658,
    new_n13659, new_n13660, new_n13661, new_n13662, new_n13663, new_n13664,
    new_n13665, new_n13666, new_n13667, new_n13668_1, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677_1, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683_1, new_n13684, new_n13685,
    new_n13686, new_n13687, new_n13688, new_n13689, new_n13690, new_n13691,
    new_n13692, new_n13693, new_n13694, new_n13695, new_n13696, new_n13697,
    new_n13698, new_n13699, new_n13700, new_n13701, new_n13702, new_n13703,
    new_n13704, new_n13705, new_n13706, new_n13707, new_n13708_1,
    new_n13709, new_n13710_1, new_n13711, new_n13712, new_n13713,
    new_n13714_1, new_n13715, new_n13716, new_n13717, new_n13718,
    new_n13719_1, new_n13720, new_n13721, new_n13722_1, new_n13723,
    new_n13724, new_n13725, new_n13726, new_n13727, new_n13728, new_n13729,
    new_n13730, new_n13731, new_n13732, new_n13733, new_n13734, new_n13735,
    new_n13736, new_n13737, new_n13738, new_n13740, new_n13742, new_n13743,
    new_n13744, new_n13745, new_n13746, new_n13747, new_n13748, new_n13749,
    new_n13750, new_n13751, new_n13752, new_n13753, new_n13754_1,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764_1, new_n13765,
    new_n13766, new_n13767, new_n13768, new_n13769, new_n13770, new_n13771,
    new_n13772, new_n13773, new_n13774, new_n13775_1, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781_1,
    new_n13782, new_n13783_1, new_n13784, new_n13785, new_n13786,
    new_n13787, new_n13788, new_n13789, new_n13790, new_n13791, new_n13792,
    new_n13793, new_n13794, new_n13795, new_n13796, new_n13797,
    new_n13798_1, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808,
    new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814,
    new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820,
    new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826,
    new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832,
    new_n13833, new_n13834, new_n13835_1, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843,
    new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850_1, new_n13851_1, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912_1, new_n13913, new_n13914_1,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922_1, new_n13923_1, new_n13924, new_n13925,
    new_n13926, new_n13927, new_n13928, new_n13929, new_n13930, new_n13931,
    new_n13932, new_n13933, new_n13934, new_n13935, new_n13936, new_n13937,
    new_n13938, new_n13939, new_n13940, new_n13941, new_n13942, new_n13943,
    new_n13944, new_n13945, new_n13946, new_n13947, new_n13948, new_n13949,
    new_n13950, new_n13951_1, new_n13952, new_n13953, new_n13954,
    new_n13955, new_n13956, new_n13957, new_n13958, new_n13959, new_n13960,
    new_n13961, new_n13962, new_n13963, new_n13964, new_n13965, new_n13966,
    new_n13967, new_n13968, new_n13969, new_n13970, new_n13971, new_n13972,
    new_n13973, new_n13974, new_n13975, new_n13976, new_n13977, new_n13978,
    new_n13979, new_n13980, new_n13981, new_n13982, new_n13983, new_n13984,
    new_n13985, new_n13986, new_n13987, new_n13988, new_n13989, new_n13990,
    new_n13991, new_n13992, new_n13993, new_n13995, new_n13996, new_n13997,
    new_n13998, new_n13999, new_n14000, new_n14001, new_n14002, new_n14003,
    new_n14004_1, new_n14005, new_n14006, new_n14007, new_n14008,
    new_n14009, new_n14010, new_n14011, new_n14012, new_n14013, new_n14014,
    new_n14015, new_n14016, new_n14017, new_n14018, new_n14019, new_n14020,
    new_n14021, new_n14022, new_n14023, new_n14024, new_n14025, new_n14026,
    new_n14027, new_n14029, new_n14031, new_n14033, new_n14034, new_n14035,
    new_n14036_1, new_n14037, new_n14038, new_n14039, new_n14040,
    new_n14041, new_n14042, new_n14043, new_n14044, new_n14045, new_n14046,
    new_n14047, new_n14048, new_n14049, new_n14050, new_n14051, new_n14052,
    new_n14053, new_n14054, new_n14055, new_n14056, new_n14057, new_n14058,
    new_n14059_1, new_n14060, new_n14061, new_n14062, new_n14063,
    new_n14064, new_n14065, new_n14066, new_n14067, new_n14068, new_n14069,
    new_n14070, new_n14071_1, new_n14072, new_n14073, new_n14074,
    new_n14075, new_n14076, new_n14077, new_n14078, new_n14079, new_n14080,
    new_n14081_1, new_n14082, new_n14083, new_n14084, new_n14085,
    new_n14086, new_n14087, new_n14088, new_n14089, new_n14090_1,
    new_n14091, new_n14092, new_n14093, new_n14095_1, new_n14097,
    new_n14098, new_n14099, new_n14100, new_n14101, new_n14102, new_n14103,
    new_n14104, new_n14105, new_n14106, new_n14107_1, new_n14108,
    new_n14109, new_n14110, new_n14111, new_n14112, new_n14113, new_n14114,
    new_n14115, new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121_1, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126_1, new_n14127, new_n14128, new_n14129, new_n14130_1,
    new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136_1, new_n14137, new_n14138, new_n14139, new_n14140,
    new_n14141, new_n14142, new_n14143, new_n14144, new_n14145, new_n14146,
    new_n14147_1, new_n14148_1, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14163,
    new_n14164, new_n14165, new_n14166, new_n14167, new_n14168, new_n14169,
    new_n14170, new_n14171, new_n14172, new_n14173, new_n14174_1,
    new_n14175, new_n14176, new_n14177, new_n14178, new_n14179, new_n14180,
    new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186,
    new_n14187, new_n14188, new_n14189, new_n14190_1, new_n14191,
    new_n14192, new_n14193, new_n14194, new_n14195, new_n14196, new_n14197,
    new_n14198, new_n14199, new_n14200, new_n14201, new_n14202, new_n14203,
    new_n14204, new_n14205, new_n14206, new_n14207, new_n14208, new_n14209,
    new_n14210, new_n14211_1, new_n14212, new_n14213, new_n14214,
    new_n14215, new_n14216, new_n14217, new_n14218, new_n14219, new_n14220,
    new_n14221, new_n14222_1, new_n14223, new_n14224, new_n14225,
    new_n14226, new_n14227, new_n14228, new_n14229, new_n14230_1,
    new_n14231, new_n14232, new_n14233, new_n14234, new_n14235, new_n14236,
    new_n14237, new_n14238, new_n14239, new_n14240, new_n14241, new_n14242,
    new_n14243, new_n14244, new_n14245, new_n14246, new_n14247, new_n14248,
    new_n14249, new_n14250, new_n14251, new_n14252, new_n14253, new_n14254,
    new_n14255, new_n14256, new_n14257, new_n14258, new_n14259, new_n14260,
    new_n14261, new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267_1, new_n14268, new_n14269, new_n14270, new_n14271_1,
    new_n14272, new_n14273, new_n14274, new_n14275_1, new_n14276,
    new_n14277_1, new_n14278, new_n14279, new_n14280, new_n14281,
    new_n14282, new_n14283, new_n14284, new_n14285, new_n14286, new_n14287,
    new_n14288, new_n14289, new_n14290, new_n14291, new_n14292, new_n14293,
    new_n14294_1, new_n14295, new_n14296, new_n14297, new_n14298,
    new_n14299, new_n14300, new_n14301, new_n14302, new_n14303, new_n14304,
    new_n14305, new_n14306, new_n14307, new_n14308, new_n14309,
    new_n14310_1, new_n14311, new_n14312, new_n14313, new_n14314,
    new_n14315, new_n14316, new_n14317, new_n14318, new_n14319, new_n14320,
    new_n14321, new_n14322, new_n14323_1, new_n14324, new_n14325,
    new_n14326_1, new_n14327, new_n14328, new_n14329, new_n14330,
    new_n14331, new_n14332, new_n14333, new_n14334, new_n14336, new_n14338,
    new_n14339, new_n14340, new_n14341, new_n14342_1, new_n14343,
    new_n14344, new_n14345_1, new_n14346, new_n14347, new_n14348,
    new_n14349, new_n14350, new_n14351, new_n14352, new_n14353_1,
    new_n14354, new_n14355, new_n14356, new_n14357, new_n14358, new_n14359,
    new_n14360, new_n14361, new_n14362, new_n14363, new_n14364_1,
    new_n14365, new_n14366, new_n14367, new_n14368, new_n14369, new_n14371,
    new_n14372, new_n14373, new_n14374, new_n14375_1, new_n14376,
    new_n14377, new_n14378, new_n14379, new_n14380, new_n14381, new_n14382,
    new_n14383, new_n14384, new_n14385, new_n14386, new_n14387, new_n14388,
    new_n14389, new_n14390, new_n14391, new_n14392, new_n14393, new_n14394,
    new_n14395, new_n14396, new_n14397, new_n14398, new_n14399, new_n14400,
    new_n14401, new_n14402, new_n14403, new_n14404, new_n14405, new_n14406,
    new_n14407, new_n14408, new_n14409, new_n14410, new_n14411,
    new_n14412_1, new_n14413, new_n14414_1, new_n14415, new_n14416,
    new_n14417, new_n14418, new_n14419, new_n14420, new_n14421, new_n14422,
    new_n14423, new_n14424, new_n14425, new_n14426, new_n14427, new_n14428,
    new_n14429, new_n14430, new_n14431, new_n14432, new_n14433, new_n14434,
    new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440_1, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457_1, new_n14458, new_n14459, new_n14460, new_n14461,
    new_n14462, new_n14463, new_n14464_1, new_n14465, new_n14466,
    new_n14467, new_n14468, new_n14469, new_n14470, new_n14471_1,
    new_n14472, new_n14473, new_n14474, new_n14475_1, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510_1, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535,
    new_n14536, new_n14537, new_n14538, new_n14539, new_n14540,
    new_n14541_1, new_n14542, new_n14543, new_n14544, new_n14545,
    new_n14546_1, new_n14547_1, new_n14548, new_n14549, new_n14550,
    new_n14551, new_n14552, new_n14553, new_n14554, new_n14555, new_n14556,
    new_n14557, new_n14558, new_n14559, new_n14560, new_n14561, new_n14562,
    new_n14563, new_n14564, new_n14565, new_n14566, new_n14567, new_n14568,
    new_n14569, new_n14570_1, new_n14571, new_n14572, new_n14573,
    new_n14574, new_n14575_1, new_n14576_1, new_n14577, new_n14578,
    new_n14579, new_n14580, new_n14581, new_n14582, new_n14583, new_n14584,
    new_n14585, new_n14586, new_n14587, new_n14588, new_n14589, new_n14590,
    new_n14591, new_n14592, new_n14593_1, new_n14594, new_n14595,
    new_n14596, new_n14597, new_n14598, new_n14599, new_n14600, new_n14601,
    new_n14602, new_n14603_1, new_n14604, new_n14605, new_n14606,
    new_n14607, new_n14608, new_n14609, new_n14610, new_n14611, new_n14612,
    new_n14613, new_n14614, new_n14615, new_n14616, new_n14617, new_n14618,
    new_n14619, new_n14620, new_n14621, new_n14622, new_n14623, new_n14624,
    new_n14625, new_n14626, new_n14627, new_n14628, new_n14629, new_n14630,
    new_n14631, new_n14632, new_n14633_1, new_n14634, new_n14635,
    new_n14636_1, new_n14637, new_n14638, new_n14639, new_n14640,
    new_n14641, new_n14642, new_n14643, new_n14644, new_n14645, new_n14646,
    new_n14647, new_n14648, new_n14649, new_n14650, new_n14651, new_n14652,
    new_n14653, new_n14654, new_n14655, new_n14656, new_n14657, new_n14658,
    new_n14659, new_n14660, new_n14661, new_n14662, new_n14663, new_n14664,
    new_n14665, new_n14666, new_n14667, new_n14668, new_n14669, new_n14670,
    new_n14671, new_n14672, new_n14673, new_n14674, new_n14675, new_n14676,
    new_n14677, new_n14678, new_n14679, new_n14680_1, new_n14681,
    new_n14682, new_n14683, new_n14684_1, new_n14685, new_n14686,
    new_n14687, new_n14688, new_n14689, new_n14690, new_n14691,
    new_n14692_1, new_n14693, new_n14694, new_n14695, new_n14696,
    new_n14697, new_n14698, new_n14699, new_n14700, new_n14701_1,
    new_n14702_1, new_n14703, new_n14704_1, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14721, new_n14723, new_n14724, new_n14725, new_n14726,
    new_n14727, new_n14728, new_n14729, new_n14730, new_n14731, new_n14732,
    new_n14733, new_n14734_1, new_n14735, new_n14736, new_n14737,
    new_n14738, new_n14739, new_n14740, new_n14741, new_n14742, new_n14743,
    new_n14744, new_n14745, new_n14746_1, new_n14747, new_n14748,
    new_n14749, new_n14750, new_n14751, new_n14752, new_n14753, new_n14754,
    new_n14755, new_n14756, new_n14757, new_n14758, new_n14759, new_n14760,
    new_n14761, new_n14762, new_n14763_1, new_n14764, new_n14765,
    new_n14766, new_n14767, new_n14768, new_n14769, new_n14770, new_n14771,
    new_n14772_1, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782,
    new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788,
    new_n14789, new_n14790_1, new_n14791, new_n14792, new_n14793,
    new_n14794, new_n14795, new_n14796, new_n14798, new_n14800, new_n14803,
    new_n14804, new_n14805, new_n14806, new_n14807, new_n14808, new_n14809,
    new_n14810, new_n14811, new_n14812, new_n14813, new_n14814, new_n14815,
    new_n14816, new_n14817, new_n14818, new_n14819_1, new_n14821,
    new_n14823, new_n14825, new_n14826_1, new_n14827_1, new_n14828,
    new_n14829, new_n14830, new_n14831, new_n14832, new_n14833, new_n14834,
    new_n14835, new_n14836, new_n14837, new_n14838, new_n14839_1,
    new_n14840, new_n14841, new_n14842, new_n14843, new_n14844, new_n14845,
    new_n14846, new_n14847, new_n14848, new_n14849_1, new_n14850,
    new_n14851, new_n14854, new_n14856, new_n14857, new_n14858, new_n14859,
    new_n14860, new_n14861, new_n14862, new_n14863, new_n14864, new_n14865,
    new_n14866, new_n14867, new_n14868, new_n14869, new_n14870, new_n14871,
    new_n14872, new_n14873, new_n14874, new_n14875, new_n14876, new_n14877,
    new_n14878, new_n14879, new_n14880, new_n14881, new_n14882, new_n14883,
    new_n14884, new_n14885, new_n14886, new_n14887, new_n14888, new_n14889,
    new_n14890, new_n14891_1, new_n14893, new_n14894, new_n14895,
    new_n14896, new_n14897, new_n14898, new_n14899_1, new_n14900,
    new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906,
    new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912,
    new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918,
    new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924,
    new_n14925, new_n14926, new_n14928, new_n14930, new_n14931_1,
    new_n14932, new_n14934, new_n14935, new_n14936, new_n14937, new_n14938,
    new_n14939, new_n14940, new_n14941, new_n14942, new_n14943,
    new_n14944_1, new_n14945, new_n14946, new_n14947, new_n14948,
    new_n14949, new_n14950, new_n14951, new_n14952, new_n14953,
    new_n14954_1, new_n14955, new_n14956, new_n14957, new_n14958,
    new_n14959, new_n14960, new_n14961, new_n14962, new_n14963, new_n14964,
    new_n14965, new_n14966, new_n14967, new_n14968, new_n14969, new_n14970,
    new_n14971, new_n14972, new_n14973, new_n14974, new_n14975, new_n14976,
    new_n14977_1, new_n14978, new_n14979, new_n14980, new_n14981,
    new_n14982, new_n14983, new_n14984, new_n14985, new_n14986, new_n14987,
    new_n14989_1, new_n14991, new_n14992, new_n14993, new_n14994,
    new_n14995, new_n14996, new_n14997, new_n14998, new_n14999, new_n15000,
    new_n15001, new_n15002_1, new_n15003, new_n15004_1, new_n15005,
    new_n15006, new_n15007, new_n15008, new_n15009, new_n15010,
    new_n15011_1, new_n15012, new_n15013, new_n15014, new_n15015,
    new_n15016, new_n15017, new_n15018, new_n15019_1, new_n15020,
    new_n15021, new_n15022, new_n15023, new_n15024, new_n15025, new_n15026,
    new_n15027, new_n15028, new_n15029, new_n15030, new_n15031_1,
    new_n15032, new_n15033_1, new_n15034, new_n15035, new_n15036,
    new_n15037, new_n15038, new_n15039, new_n15040, new_n15041, new_n15042,
    new_n15043, new_n15044, new_n15045, new_n15046, new_n15047, new_n15048,
    new_n15049, new_n15050, new_n15051, new_n15052_1, new_n15053_1,
    new_n15054, new_n15055, new_n15056, new_n15057, new_n15058, new_n15059,
    new_n15060, new_n15061, new_n15062, new_n15063, new_n15064, new_n15065,
    new_n15066, new_n15067, new_n15068, new_n15069, new_n15070, new_n15071,
    new_n15072, new_n15073, new_n15074, new_n15075, new_n15076,
    new_n15077_1, new_n15078, new_n15079, new_n15080, new_n15081,
    new_n15082_1, new_n15083, new_n15084, new_n15085, new_n15086,
    new_n15087, new_n15088, new_n15089, new_n15090, new_n15091, new_n15092,
    new_n15093, new_n15094_1, new_n15095, new_n15096, new_n15097,
    new_n15098, new_n15099, new_n15100, new_n15101, new_n15102, new_n15103,
    new_n15104, new_n15106, new_n15107, new_n15108, new_n15109, new_n15110,
    new_n15111, new_n15112, new_n15113, new_n15114, new_n15115, new_n15116,
    new_n15117, new_n15118_1, new_n15119, new_n15120, new_n15121,
    new_n15122, new_n15123, new_n15124, new_n15125, new_n15126, new_n15127,
    new_n15128_1, new_n15129, new_n15130, new_n15131, new_n15132,
    new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138,
    new_n15139_1, new_n15140, new_n15141, new_n15142, new_n15143,
    new_n15144, new_n15145_1, new_n15146_1, new_n15147, new_n15148,
    new_n15149, new_n15150, new_n15151, new_n15152, new_n15153, new_n15154,
    new_n15155, new_n15156, new_n15157, new_n15158, new_n15159, new_n15160,
    new_n15161, new_n15162, new_n15163, new_n15164, new_n15165_1,
    new_n15166, new_n15167_1, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175,
    new_n15176_1, new_n15177, new_n15178, new_n15179, new_n15180_1,
    new_n15181, new_n15182_1, new_n15183, new_n15184, new_n15185,
    new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191,
    new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197,
    new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203,
    new_n15204, new_n15205_1, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230_1, new_n15232,
    new_n15233, new_n15234, new_n15235, new_n15236, new_n15237, new_n15238,
    new_n15239, new_n15240, new_n15241_1, new_n15242, new_n15243,
    new_n15244, new_n15245, new_n15246, new_n15247, new_n15248, new_n15249,
    new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15255_1, new_n15256, new_n15257, new_n15258_1, new_n15259,
    new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265,
    new_n15266, new_n15267, new_n15268, new_n15269, new_n15270,
    new_n15271_1, new_n15272, new_n15273, new_n15274, new_n15275_1,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15286, new_n15288,
    new_n15289_1, new_n15290, new_n15291, new_n15292, new_n15293,
    new_n15294, new_n15295, new_n15296, new_n15297, new_n15298, new_n15299,
    new_n15300_1, new_n15301, new_n15303, new_n15304, new_n15305,
    new_n15306, new_n15307_1, new_n15308, new_n15309, new_n15310,
    new_n15311, new_n15312, new_n15313, new_n15314, new_n15315, new_n15316,
    new_n15317, new_n15318, new_n15319, new_n15320, new_n15321, new_n15322,
    new_n15323, new_n15324, new_n15325, new_n15326, new_n15327_1,
    new_n15328, new_n15329, new_n15330, new_n15331, new_n15332_1,
    new_n15333, new_n15334, new_n15335, new_n15336, new_n15337, new_n15338,
    new_n15339, new_n15340, new_n15341, new_n15342, new_n15343, new_n15344,
    new_n15345_1, new_n15346, new_n15347, new_n15348, new_n15349,
    new_n15350, new_n15351, new_n15352, new_n15353_1, new_n15354,
    new_n15355, new_n15356, new_n15357, new_n15358, new_n15359, new_n15360,
    new_n15361, new_n15362, new_n15363, new_n15364, new_n15365,
    new_n15366_1, new_n15367, new_n15368, new_n15369, new_n15370,
    new_n15371, new_n15372, new_n15373, new_n15374, new_n15375, new_n15376,
    new_n15377, new_n15378_1, new_n15379, new_n15380, new_n15381,
    new_n15382_1, new_n15383, new_n15384, new_n15385, new_n15386,
    new_n15387, new_n15388, new_n15389, new_n15390, new_n15391, new_n15392,
    new_n15393, new_n15394, new_n15395, new_n15396, new_n15397, new_n15398,
    new_n15399, new_n15400, new_n15401, new_n15402, new_n15403, new_n15404,
    new_n15405, new_n15406, new_n15407_1, new_n15408, new_n15409,
    new_n15410, new_n15411, new_n15412, new_n15413, new_n15414, new_n15415,
    new_n15416, new_n15417, new_n15418, new_n15419, new_n15420, new_n15421,
    new_n15422, new_n15423, new_n15424_1, new_n15425, new_n15426,
    new_n15427, new_n15428_1, new_n15429, new_n15430, new_n15431,
    new_n15432, new_n15433, new_n15434, new_n15435_1, new_n15436,
    new_n15437, new_n15438_1, new_n15439, new_n15440, new_n15441,
    new_n15442, new_n15443, new_n15444, new_n15445, new_n15446, new_n15447,
    new_n15448, new_n15449, new_n15450, new_n15451, new_n15452, new_n15453,
    new_n15454, new_n15455, new_n15456, new_n15457, new_n15458, new_n15459,
    new_n15460, new_n15461, new_n15462, new_n15463, new_n15464,
    new_n15465_1, new_n15466, new_n15467_1, new_n15468, new_n15469,
    new_n15470_1, new_n15471, new_n15472, new_n15473, new_n15474,
    new_n15475, new_n15476, new_n15477_1, new_n15478, new_n15480,
    new_n15482, new_n15483, new_n15484, new_n15485, new_n15486, new_n15487,
    new_n15488, new_n15489, new_n15490_1, new_n15491, new_n15492,
    new_n15493, new_n15494, new_n15495, new_n15496_1, new_n15497,
    new_n15498, new_n15499, new_n15500, new_n15501_1, new_n15502,
    new_n15503, new_n15504, new_n15505, new_n15506_1, new_n15507,
    new_n15508_1, new_n15509, new_n15510, new_n15511, new_n15512,
    new_n15513, new_n15514, new_n15515, new_n15516, new_n15517, new_n15518,
    new_n15519, new_n15520, new_n15521, new_n15522, new_n15523, new_n15524,
    new_n15525, new_n15526, new_n15527, new_n15528, new_n15529, new_n15530,
    new_n15531, new_n15532, new_n15533, new_n15534, new_n15535, new_n15536,
    new_n15537, new_n15538, new_n15539_1, new_n15540, new_n15541,
    new_n15542, new_n15543, new_n15544, new_n15545, new_n15546_1,
    new_n15547, new_n15548, new_n15549, new_n15550, new_n15551, new_n15552,
    new_n15553, new_n15554, new_n15555_1, new_n15556, new_n15557,
    new_n15558_1, new_n15559_1, new_n15560, new_n15561, new_n15562,
    new_n15563, new_n15564, new_n15565, new_n15566, new_n15567, new_n15568,
    new_n15569, new_n15570_1, new_n15571, new_n15572, new_n15573_1,
    new_n15574, new_n15575, new_n15576, new_n15578, new_n15579, new_n15580,
    new_n15581, new_n15582, new_n15584, new_n15586, new_n15587,
    new_n15588_1, new_n15589, new_n15590_1, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597,
    new_n15598_1, new_n15599, new_n15600, new_n15601, new_n15602_1,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613,
    new_n15614_1, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635,
    new_n15636_1, new_n15637, new_n15638, new_n15639, new_n15640,
    new_n15641, new_n15642, new_n15643, new_n15644, new_n15645, new_n15646,
    new_n15647, new_n15648, new_n15649, new_n15650, new_n15651,
    new_n15652_1, new_n15653, new_n15654, new_n15655, new_n15656,
    new_n15657, new_n15658, new_n15659, new_n15660, new_n15661,
    new_n15662_1, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15684, new_n15685,
    new_n15686, new_n15687, new_n15688, new_n15689, new_n15690, new_n15691,
    new_n15692, new_n15693, new_n15694, new_n15695, new_n15696, new_n15697,
    new_n15698, new_n15699, new_n15700, new_n15701, new_n15702, new_n15703,
    new_n15704, new_n15705, new_n15706, new_n15707, new_n15708, new_n15709,
    new_n15710, new_n15711, new_n15712, new_n15713, new_n15714, new_n15715,
    new_n15716_1, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726,
    new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732,
    new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738,
    new_n15739, new_n15740, new_n15741, new_n15742, new_n15743_1,
    new_n15744, new_n15745, new_n15746, new_n15747, new_n15748,
    new_n15749_1, new_n15750, new_n15751, new_n15752, new_n15753,
    new_n15754, new_n15755, new_n15756, new_n15757, new_n15758, new_n15759,
    new_n15760, new_n15761_1, new_n15762_1, new_n15763, new_n15764,
    new_n15765, new_n15766_1, new_n15767, new_n15768, new_n15769,
    new_n15770, new_n15771, new_n15772, new_n15773, new_n15774, new_n15775,
    new_n15776, new_n15777, new_n15778, new_n15779, new_n15780_1,
    new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786,
    new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793_1, new_n15794, new_n15795, new_n15796, new_n15797,
    new_n15798, new_n15799, new_n15800, new_n15801, new_n15802, new_n15803,
    new_n15804, new_n15805, new_n15806, new_n15807, new_n15808, new_n15809,
    new_n15810, new_n15811, new_n15812_1, new_n15814, new_n15816_1,
    new_n15817, new_n15818, new_n15819, new_n15820, new_n15821, new_n15822,
    new_n15823, new_n15824, new_n15825, new_n15826, new_n15827, new_n15828,
    new_n15829, new_n15830, new_n15831_1, new_n15832, new_n15833,
    new_n15834, new_n15835, new_n15836, new_n15837, new_n15838, new_n15839,
    new_n15840, new_n15841, new_n15842, new_n15843, new_n15844, new_n15845,
    new_n15846_1, new_n15847, new_n15848, new_n15849, new_n15850,
    new_n15851, new_n15852, new_n15853, new_n15854, new_n15855, new_n15856,
    new_n15857, new_n15858, new_n15859_1, new_n15860, new_n15861,
    new_n15862, new_n15863, new_n15864, new_n15865, new_n15866, new_n15867,
    new_n15868, new_n15869_1, new_n15870, new_n15871, new_n15873,
    new_n15875, new_n15876, new_n15877, new_n15878, new_n15879, new_n15880,
    new_n15881, new_n15882, new_n15883, new_n15884_1, new_n15885_1,
    new_n15886, new_n15887, new_n15888, new_n15889_1, new_n15890,
    new_n15891, new_n15892, new_n15893, new_n15894, new_n15895, new_n15896,
    new_n15897, new_n15898, new_n15899, new_n15900, new_n15901, new_n15902,
    new_n15903, new_n15904, new_n15905, new_n15906, new_n15907, new_n15908,
    new_n15909, new_n15910, new_n15911, new_n15912, new_n15913, new_n15914,
    new_n15915, new_n15916, new_n15917_1, new_n15918_1, new_n15919,
    new_n15920, new_n15921, new_n15922_1, new_n15923, new_n15924,
    new_n15925, new_n15926, new_n15927, new_n15928, new_n15929, new_n15930,
    new_n15931, new_n15932, new_n15933, new_n15934, new_n15935,
    new_n15936_1, new_n15937, new_n15938, new_n15939, new_n15940,
    new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946,
    new_n15947_1, new_n15948, new_n15949, new_n15950, new_n15951,
    new_n15952, new_n15953, new_n15954, new_n15955, new_n15956_1,
    new_n15957, new_n15958_1, new_n15959, new_n15960, new_n15961,
    new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967_1, new_n15968, new_n15969, new_n15970, new_n15971,
    new_n15972, new_n15973, new_n15974, new_n15975, new_n15976, new_n15977,
    new_n15978, new_n15979_1, new_n15980, new_n15981, new_n15982,
    new_n15983, new_n15984, new_n15985, new_n15986_1, new_n15987,
    new_n15988, new_n15989, new_n15990, new_n15991, new_n15992, new_n15993,
    new_n15994, new_n15995, new_n15996, new_n15997, new_n15998, new_n15999,
    new_n16000, new_n16001, new_n16002, new_n16003, new_n16004, new_n16005,
    new_n16006, new_n16007, new_n16008, new_n16009, new_n16010, new_n16011,
    new_n16012, new_n16013_1, new_n16014, new_n16015, new_n16016,
    new_n16018, new_n16019, new_n16020, new_n16021, new_n16022, new_n16023,
    new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029_1, new_n16030, new_n16031, new_n16032, new_n16033,
    new_n16034, new_n16035, new_n16036, new_n16037, new_n16038, new_n16039,
    new_n16040, new_n16041, new_n16042, new_n16043, new_n16044, new_n16045,
    new_n16046, new_n16047, new_n16049, new_n16050, new_n16051, new_n16052,
    new_n16053, new_n16054, new_n16055, new_n16056, new_n16057, new_n16058,
    new_n16059, new_n16060_1, new_n16061, new_n16062_1, new_n16063,
    new_n16064, new_n16065, new_n16066, new_n16067, new_n16068_1,
    new_n16069, new_n16070, new_n16071, new_n16072, new_n16073, new_n16074,
    new_n16075, new_n16076, new_n16077, new_n16078, new_n16079,
    new_n16080_1, new_n16081, new_n16082, new_n16083, new_n16084,
    new_n16085, new_n16086, new_n16087, new_n16088, new_n16089, new_n16090,
    new_n16091, new_n16092, new_n16093, new_n16094, new_n16095, new_n16096,
    new_n16097, new_n16098_1, new_n16099, new_n16100, new_n16101,
    new_n16102, new_n16103, new_n16104, new_n16105, new_n16106, new_n16107,
    new_n16108, new_n16109, new_n16110_1, new_n16111, new_n16112,
    new_n16113, new_n16114, new_n16115, new_n16116, new_n16117, new_n16118,
    new_n16119, new_n16120, new_n16121, new_n16122, new_n16123, new_n16124,
    new_n16125, new_n16126, new_n16127, new_n16128, new_n16129, new_n16130,
    new_n16131, new_n16132, new_n16133, new_n16134, new_n16135, new_n16136,
    new_n16137, new_n16138, new_n16139, new_n16140, new_n16141,
    new_n16142_1, new_n16143, new_n16144, new_n16145, new_n16146,
    new_n16147, new_n16148, new_n16149, new_n16150, new_n16151, new_n16152,
    new_n16153, new_n16154, new_n16155, new_n16156, new_n16157,
    new_n16158_1, new_n16159, new_n16160, new_n16161, new_n16162,
    new_n16163, new_n16164, new_n16165, new_n16166, new_n16167_1,
    new_n16168, new_n16169, new_n16170, new_n16171, new_n16172, new_n16173,
    new_n16174, new_n16175, new_n16176, new_n16177, new_n16178, new_n16179,
    new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185_1, new_n16186, new_n16187, new_n16188, new_n16189,
    new_n16190, new_n16191, new_n16192, new_n16193, new_n16194, new_n16195,
    new_n16196_1, new_n16197, new_n16198, new_n16199, new_n16200,
    new_n16201, new_n16202, new_n16203, new_n16204, new_n16205,
    new_n16206_1, new_n16207, new_n16208, new_n16209, new_n16210,
    new_n16211, new_n16212, new_n16213, new_n16214, new_n16215_1,
    new_n16216, new_n16217_1, new_n16218_1, new_n16219_1, new_n16220,
    new_n16221, new_n16222, new_n16223_1, new_n16224, new_n16225,
    new_n16226, new_n16227, new_n16228, new_n16229, new_n16230_1,
    new_n16231, new_n16232, new_n16233, new_n16234, new_n16235, new_n16236,
    new_n16237, new_n16238, new_n16239, new_n16240, new_n16241, new_n16242,
    new_n16243_1, new_n16244, new_n16245, new_n16246, new_n16247_1,
    new_n16248, new_n16249, new_n16250, new_n16251, new_n16252, new_n16253,
    new_n16254, new_n16255, new_n16256, new_n16257, new_n16258, new_n16259,
    new_n16260, new_n16261, new_n16262, new_n16263, new_n16265, new_n16266,
    new_n16267, new_n16268, new_n16269, new_n16270, new_n16271, new_n16272,
    new_n16273, new_n16274, new_n16275_1, new_n16276, new_n16277,
    new_n16278, new_n16279_1, new_n16280, new_n16281, new_n16282,
    new_n16283, new_n16284, new_n16285, new_n16286, new_n16287, new_n16288,
    new_n16289, new_n16290, new_n16291, new_n16292, new_n16293, new_n16294,
    new_n16295, new_n16296, new_n16297, new_n16298, new_n16299, new_n16300,
    new_n16301, new_n16302, new_n16303, new_n16304, new_n16305, new_n16306,
    new_n16307, new_n16308, new_n16309, new_n16310, new_n16311, new_n16312,
    new_n16313, new_n16314, new_n16315, new_n16316, new_n16317, new_n16318,
    new_n16319, new_n16320, new_n16321, new_n16322_1, new_n16323,
    new_n16324, new_n16325, new_n16326, new_n16327_1, new_n16328,
    new_n16329, new_n16330, new_n16331, new_n16332, new_n16333, new_n16334,
    new_n16335, new_n16336, new_n16337, new_n16338, new_n16339, new_n16340,
    new_n16341, new_n16342, new_n16343, new_n16344, new_n16345, new_n16346,
    new_n16347, new_n16348, new_n16349, new_n16350_1, new_n16351,
    new_n16352, new_n16353, new_n16354, new_n16355, new_n16356, new_n16357,
    new_n16358, new_n16359, new_n16360, new_n16361, new_n16362, new_n16363,
    new_n16364, new_n16365, new_n16366, new_n16367_1, new_n16368,
    new_n16369, new_n16370, new_n16371, new_n16372, new_n16373, new_n16374,
    new_n16375, new_n16376_1, new_n16377, new_n16378, new_n16379_1,
    new_n16380, new_n16381, new_n16382, new_n16383, new_n16384, new_n16385,
    new_n16386, new_n16387, new_n16388, new_n16389, new_n16390, new_n16391,
    new_n16392, new_n16393, new_n16394, new_n16395, new_n16396_1,
    new_n16397, new_n16398_1, new_n16399, new_n16400, new_n16401,
    new_n16402, new_n16403, new_n16404, new_n16405, new_n16406_1,
    new_n16407_1, new_n16408, new_n16409, new_n16410, new_n16411,
    new_n16412, new_n16413, new_n16414, new_n16415, new_n16416, new_n16417,
    new_n16418, new_n16419_1, new_n16420, new_n16421, new_n16422,
    new_n16423, new_n16424_1, new_n16425, new_n16426, new_n16427,
    new_n16428_1, new_n16429, new_n16430, new_n16431, new_n16432,
    new_n16433_1, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439_1, new_n16440_1, new_n16441, new_n16442,
    new_n16443, new_n16444, new_n16445_1, new_n16446, new_n16447,
    new_n16448, new_n16449, new_n16450, new_n16451, new_n16452, new_n16453,
    new_n16454, new_n16455, new_n16456, new_n16457, new_n16458, new_n16459,
    new_n16460_1, new_n16461, new_n16462, new_n16463, new_n16464,
    new_n16465, new_n16467, new_n16468, new_n16469, new_n16470, new_n16471,
    new_n16472, new_n16473, new_n16474, new_n16475, new_n16476_1,
    new_n16477, new_n16478, new_n16479, new_n16480, new_n16481_1,
    new_n16482_1, new_n16483, new_n16484, new_n16485, new_n16486,
    new_n16487, new_n16488, new_n16489, new_n16490, new_n16491, new_n16492,
    new_n16493_1, new_n16494, new_n16495, new_n16496, new_n16497,
    new_n16498, new_n16499, new_n16500, new_n16501, new_n16502_1,
    new_n16503, new_n16504, new_n16505, new_n16506_1, new_n16507_1,
    new_n16508, new_n16509, new_n16510, new_n16511, new_n16512, new_n16513,
    new_n16514, new_n16515, new_n16516_1, new_n16517_1, new_n16518,
    new_n16519, new_n16520, new_n16521_1, new_n16522, new_n16523,
    new_n16524_1, new_n16525, new_n16526, new_n16527_1, new_n16528,
    new_n16529, new_n16530, new_n16531, new_n16532, new_n16533, new_n16534,
    new_n16535, new_n16536, new_n16537, new_n16538, new_n16539, new_n16540,
    new_n16541, new_n16542, new_n16543, new_n16544_1, new_n16545,
    new_n16546, new_n16547, new_n16548, new_n16549, new_n16550, new_n16551,
    new_n16552, new_n16553, new_n16554_1, new_n16555, new_n16556,
    new_n16557, new_n16558, new_n16559, new_n16560, new_n16561, new_n16562,
    new_n16563, new_n16564, new_n16565, new_n16566, new_n16567, new_n16568,
    new_n16569, new_n16570, new_n16571, new_n16572, new_n16573, new_n16574,
    new_n16575, new_n16576, new_n16577, new_n16578, new_n16579, new_n16580,
    new_n16581, new_n16582, new_n16583_1, new_n16584_1, new_n16585,
    new_n16586, new_n16587, new_n16588, new_n16589_1, new_n16590,
    new_n16591, new_n16592, new_n16593, new_n16594, new_n16595,
    new_n16596_1, new_n16597, new_n16598, new_n16599, new_n16600,
    new_n16601, new_n16602, new_n16603, new_n16604, new_n16605, new_n16606,
    new_n16607, new_n16608_1, new_n16609, new_n16610, new_n16611,
    new_n16612, new_n16613, new_n16614, new_n16615, new_n16616,
    new_n16617_1, new_n16618, new_n16619, new_n16620, new_n16621,
    new_n16622, new_n16623, new_n16624, new_n16625, new_n16626, new_n16627,
    new_n16628, new_n16629, new_n16630_1, new_n16631, new_n16632,
    new_n16633, new_n16634, new_n16635, new_n16637, new_n16638, new_n16639,
    new_n16640_1, new_n16641, new_n16642, new_n16643, new_n16644,
    new_n16645, new_n16646, new_n16647, new_n16648, new_n16649, new_n16650,
    new_n16651, new_n16652, new_n16653, new_n16654, new_n16655,
    new_n16656_1, new_n16657, new_n16658, new_n16659, new_n16660,
    new_n16661, new_n16662, new_n16663, new_n16664, new_n16665, new_n16666,
    new_n16667, new_n16668, new_n16669, new_n16670, new_n16671, new_n16672,
    new_n16673, new_n16674_1, new_n16675, new_n16676, new_n16677,
    new_n16678, new_n16679, new_n16680, new_n16681, new_n16682_1,
    new_n16683, new_n16684_1, new_n16685, new_n16686, new_n16687,
    new_n16688_1, new_n16689, new_n16690, new_n16691, new_n16692,
    new_n16693, new_n16694, new_n16695, new_n16696, new_n16697, new_n16698,
    new_n16699, new_n16700, new_n16701, new_n16702, new_n16703, new_n16704,
    new_n16705, new_n16706, new_n16707, new_n16708, new_n16709, new_n16710,
    new_n16711, new_n16712, new_n16713, new_n16714, new_n16715, new_n16716,
    new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722_1, new_n16723, new_n16724, new_n16725, new_n16726,
    new_n16727, new_n16728, new_n16729, new_n16730, new_n16731, new_n16732,
    new_n16733_1, new_n16734, new_n16735, new_n16736, new_n16737,
    new_n16738, new_n16739, new_n16740, new_n16741, new_n16742,
    new_n16743_1, new_n16744, new_n16745, new_n16746, new_n16747,
    new_n16748, new_n16749, new_n16750, new_n16751, new_n16752, new_n16753,
    new_n16754, new_n16755, new_n16756, new_n16757, new_n16758, new_n16759,
    new_n16760, new_n16761, new_n16762, new_n16763, new_n16764, new_n16765,
    new_n16766, new_n16768, new_n16769, new_n16770, new_n16771, new_n16772,
    new_n16773, new_n16774, new_n16775, new_n16776, new_n16777, new_n16778,
    new_n16779, new_n16780, new_n16781, new_n16782, new_n16783, new_n16784,
    new_n16785, new_n16786, new_n16787, new_n16788, new_n16789, new_n16790,
    new_n16791, new_n16792, new_n16793, new_n16794, new_n16795, new_n16796,
    new_n16797, new_n16798_1, new_n16799, new_n16800, new_n16801,
    new_n16802, new_n16803, new_n16804, new_n16805, new_n16806, new_n16807,
    new_n16808, new_n16809, new_n16810, new_n16811, new_n16812_1,
    new_n16813, new_n16814, new_n16815, new_n16816, new_n16817,
    new_n16818_1, new_n16819, new_n16820, new_n16821, new_n16822,
    new_n16823, new_n16824_1, new_n16825, new_n16826, new_n16827,
    new_n16828, new_n16829, new_n16830, new_n16831, new_n16832, new_n16833,
    new_n16834_1, new_n16835, new_n16836, new_n16837_1, new_n16839,
    new_n16841_1, new_n16842, new_n16843, new_n16844, new_n16845,
    new_n16846, new_n16847, new_n16848, new_n16849, new_n16850, new_n16851,
    new_n16852, new_n16853, new_n16854, new_n16855, new_n16856, new_n16857,
    new_n16858, new_n16859, new_n16860, new_n16861, new_n16862, new_n16863,
    new_n16864, new_n16865, new_n16866, new_n16867, new_n16868, new_n16869,
    new_n16870, new_n16871, new_n16872, new_n16873, new_n16874, new_n16875,
    new_n16876, new_n16877, new_n16878, new_n16879, new_n16880, new_n16881,
    new_n16882, new_n16883, new_n16884, new_n16885_1, new_n16886,
    new_n16887, new_n16888, new_n16889, new_n16890, new_n16891, new_n16892,
    new_n16893, new_n16894, new_n16895, new_n16896, new_n16897, new_n16898,
    new_n16899, new_n16900, new_n16901, new_n16902, new_n16903, new_n16904,
    new_n16905_1, new_n16906, new_n16907, new_n16908, new_n16909,
    new_n16910, new_n16911_1, new_n16912, new_n16913, new_n16914,
    new_n16915, new_n16916, new_n16917, new_n16918, new_n16919, new_n16920,
    new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926,
    new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951_1, new_n16952, new_n16953, new_n16954_1, new_n16955,
    new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961,
    new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967,
    new_n16968_1, new_n16969, new_n16970, new_n16971_1, new_n16972,
    new_n16973, new_n16974, new_n16975, new_n16976, new_n16977, new_n16978,
    new_n16979, new_n16980, new_n16981, new_n16982, new_n16983, new_n16984,
    new_n16985, new_n16986, new_n16987, new_n16988_1, new_n16989_1,
    new_n16990, new_n16991, new_n16992, new_n16993, new_n16994_1,
    new_n16995, new_n16996, new_n16997, new_n16999, new_n17000, new_n17001,
    new_n17002, new_n17003, new_n17004, new_n17005, new_n17006_1,
    new_n17007, new_n17008, new_n17009, new_n17010, new_n17011, new_n17012,
    new_n17013, new_n17014, new_n17015, new_n17016, new_n17017, new_n17018,
    new_n17019, new_n17020, new_n17021, new_n17022, new_n17023, new_n17024,
    new_n17025, new_n17026, new_n17027, new_n17028, new_n17029, new_n17030,
    new_n17031, new_n17032, new_n17033, new_n17034, new_n17035_1,
    new_n17036, new_n17037_1, new_n17038, new_n17039, new_n17040,
    new_n17041, new_n17042, new_n17043, new_n17044, new_n17045, new_n17046,
    new_n17047, new_n17048, new_n17049, new_n17050, new_n17051, new_n17052,
    new_n17053, new_n17054, new_n17055, new_n17056, new_n17057, new_n17058,
    new_n17059, new_n17060, new_n17061, new_n17062, new_n17063, new_n17064,
    new_n17065, new_n17066, new_n17067, new_n17068_1, new_n17069_1,
    new_n17070_1, new_n17071, new_n17072, new_n17073, new_n17074,
    new_n17075_1, new_n17076, new_n17077_1, new_n17078, new_n17079,
    new_n17080, new_n17081, new_n17082, new_n17083, new_n17084_1,
    new_n17085, new_n17086, new_n17087, new_n17088, new_n17089,
    new_n17090_1, new_n17091, new_n17092, new_n17093, new_n17094,
    new_n17095_1, new_n17096, new_n17097, new_n17098, new_n17099,
    new_n17100, new_n17101, new_n17102, new_n17103, new_n17104_1,
    new_n17105, new_n17106_1, new_n17107, new_n17108, new_n17109,
    new_n17110, new_n17111, new_n17112, new_n17113, new_n17114, new_n17115,
    new_n17116, new_n17117, new_n17118, new_n17119_1, new_n17120,
    new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126,
    new_n17127, new_n17128, new_n17129, new_n17131, new_n17133, new_n17135,
    new_n17137, new_n17139, new_n17141, new_n17143, new_n17144, new_n17145,
    new_n17146, new_n17147, new_n17148, new_n17149, new_n17150, new_n17151,
    new_n17152, new_n17153, new_n17154, new_n17155, new_n17156, new_n17157,
    new_n17158, new_n17160, new_n17161, new_n17162, new_n17163_1,
    new_n17164, new_n17165, new_n17166, new_n17167, new_n17168_1,
    new_n17169, new_n17170, new_n17171, new_n17172, new_n17173, new_n17174,
    new_n17175, new_n17176, new_n17177, new_n17178, new_n17179, new_n17180,
    new_n17181, new_n17182, new_n17183, new_n17184, new_n17185, new_n17186,
    new_n17187, new_n17188, new_n17189, new_n17190, new_n17191, new_n17192,
    new_n17193, new_n17194, new_n17195, new_n17196, new_n17197, new_n17198,
    new_n17199, new_n17200, new_n17201, new_n17202_1, new_n17203,
    new_n17204, new_n17205, new_n17206, new_n17209, new_n17210, new_n17211,
    new_n17212, new_n17213, new_n17214, new_n17215, new_n17216, new_n17217,
    new_n17218, new_n17219_1, new_n17220, new_n17221, new_n17222,
    new_n17223, new_n17224, new_n17225, new_n17226, new_n17227, new_n17228,
    new_n17229, new_n17230, new_n17231, new_n17232_1, new_n17233,
    new_n17234, new_n17235, new_n17236_1, new_n17237, new_n17238,
    new_n17239, new_n17240, new_n17241, new_n17242, new_n17243_1,
    new_n17244, new_n17245, new_n17246, new_n17247, new_n17248, new_n17249,
    new_n17250_1, new_n17251_1, new_n17252, new_n17253, new_n17254,
    new_n17255, new_n17256, new_n17257, new_n17258, new_n17259, new_n17260,
    new_n17261, new_n17262, new_n17263_1, new_n17264, new_n17265,
    new_n17266, new_n17267, new_n17268, new_n17269, new_n17270, new_n17271,
    new_n17272, new_n17273, new_n17274, new_n17275, new_n17276, new_n17277,
    new_n17279, new_n17281, new_n17283, new_n17285_1, new_n17287,
    new_n17288, new_n17289, new_n17290, new_n17291, new_n17292, new_n17293,
    new_n17294, new_n17295, new_n17296, new_n17297, new_n17298, new_n17299,
    new_n17300, new_n17301, new_n17302_1, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320_1, new_n17321,
    new_n17322, new_n17323, new_n17324, new_n17325, new_n17326, new_n17327,
    new_n17328, new_n17329, new_n17330, new_n17331, new_n17332, new_n17333,
    new_n17334, new_n17335, new_n17336, new_n17337_1, new_n17338,
    new_n17339, new_n17340, new_n17341, new_n17342, new_n17343,
    new_n17344_1, new_n17345, new_n17346, new_n17347, new_n17348,
    new_n17349, new_n17350, new_n17351_1, new_n17352, new_n17353,
    new_n17354, new_n17355, new_n17356, new_n17357, new_n17358,
    new_n17359_1, new_n17360, new_n17361, new_n17362, new_n17363,
    new_n17364, new_n17365, new_n17366, new_n17367, new_n17368, new_n17369,
    new_n17370, new_n17371, new_n17372, new_n17373, new_n17374, new_n17375,
    new_n17376, new_n17377, new_n17378, new_n17379, new_n17380, new_n17381,
    new_n17382, new_n17383, new_n17384, new_n17385, new_n17386,
    new_n17387_1, new_n17388, new_n17389, new_n17390, new_n17391_1,
    new_n17392_1, new_n17393, new_n17394, new_n17395, new_n17396,
    new_n17397, new_n17398, new_n17399, new_n17400, new_n17401, new_n17402,
    new_n17403, new_n17404, new_n17405, new_n17406, new_n17407, new_n17408,
    new_n17409, new_n17410, new_n17411, new_n17412, new_n17413, new_n17414,
    new_n17415, new_n17416, new_n17417, new_n17418, new_n17419, new_n17420,
    new_n17421_1, new_n17422, new_n17423, new_n17424, new_n17425,
    new_n17426, new_n17427, new_n17428, new_n17429, new_n17430, new_n17431,
    new_n17432_1, new_n17433, new_n17434, new_n17435, new_n17436_1,
    new_n17437, new_n17438, new_n17439, new_n17440_1, new_n17441,
    new_n17442, new_n17444, new_n17446, new_n17447, new_n17448, new_n17449,
    new_n17450_1, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17458_1, new_n17459,
    new_n17460, new_n17461_1, new_n17462, new_n17463, new_n17464,
    new_n17465, new_n17466_1, new_n17467, new_n17468, new_n17469,
    new_n17470, new_n17471, new_n17472, new_n17473, new_n17474, new_n17475,
    new_n17476, new_n17477, new_n17478, new_n17479, new_n17480, new_n17481,
    new_n17482, new_n17483, new_n17484, new_n17485, new_n17486, new_n17487,
    new_n17488, new_n17489, new_n17490, new_n17491, new_n17492,
    new_n17493_1, new_n17494, new_n17495, new_n17496, new_n17497,
    new_n17498, new_n17499, new_n17500_1, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17508,
    new_n17509, new_n17510, new_n17511, new_n17513, new_n17514, new_n17515,
    new_n17516, new_n17517, new_n17518, new_n17519, new_n17520, new_n17521,
    new_n17522, new_n17523, new_n17524_1, new_n17525, new_n17526,
    new_n17527, new_n17528, new_n17529_1, new_n17530, new_n17531,
    new_n17532, new_n17533, new_n17534, new_n17535, new_n17536, new_n17537,
    new_n17538, new_n17539, new_n17540, new_n17541, new_n17542, new_n17543,
    new_n17544, new_n17545, new_n17546, new_n17547, new_n17549, new_n17551,
    new_n17552, new_n17553, new_n17554, new_n17555, new_n17556,
    new_n17557_1, new_n17558, new_n17559, new_n17560, new_n17561,
    new_n17562, new_n17563, new_n17564, new_n17565, new_n17566, new_n17567,
    new_n17568, new_n17569, new_n17570, new_n17571, new_n17572, new_n17573,
    new_n17574, new_n17575, new_n17576, new_n17577, new_n17578, new_n17579,
    new_n17580, new_n17581, new_n17582, new_n17583_1, new_n17584,
    new_n17585, new_n17586, new_n17587, new_n17588, new_n17589, new_n17590,
    new_n17591, new_n17592_1, new_n17594, new_n17595, new_n17596,
    new_n17597, new_n17598, new_n17599, new_n17600, new_n17601, new_n17602,
    new_n17603, new_n17604, new_n17605, new_n17606, new_n17607, new_n17608,
    new_n17609, new_n17610, new_n17611, new_n17612, new_n17613, new_n17614,
    new_n17615, new_n17616, new_n17617, new_n17618, new_n17619, new_n17620,
    new_n17621, new_n17622, new_n17623, new_n17624, new_n17625, new_n17626,
    new_n17627, new_n17628, new_n17629, new_n17630, new_n17631, new_n17632,
    new_n17633, new_n17634, new_n17635, new_n17636, new_n17637,
    new_n17638_1, new_n17639, new_n17640, new_n17641, new_n17642,
    new_n17644, new_n17645, new_n17646, new_n17647, new_n17648, new_n17649,
    new_n17650, new_n17651, new_n17652, new_n17653, new_n17654, new_n17655,
    new_n17656, new_n17657, new_n17658, new_n17659, new_n17660, new_n17661,
    new_n17662, new_n17663, new_n17664_1, new_n17665, new_n17666,
    new_n17667, new_n17668, new_n17669, new_n17670, new_n17671, new_n17672,
    new_n17673, new_n17674, new_n17675, new_n17676, new_n17677, new_n17678,
    new_n17679, new_n17680, new_n17681, new_n17682, new_n17683, new_n17684,
    new_n17685, new_n17686, new_n17687_1, new_n17688, new_n17689,
    new_n17690, new_n17691, new_n17692, new_n17693, new_n17694, new_n17695,
    new_n17696, new_n17697, new_n17698, new_n17699, new_n17700, new_n17701,
    new_n17702, new_n17703, new_n17704, new_n17705, new_n17706, new_n17707,
    new_n17708, new_n17709, new_n17710, new_n17711, new_n17712, new_n17713,
    new_n17714, new_n17715, new_n17716, new_n17717, new_n17718, new_n17719,
    new_n17720, new_n17721_1, new_n17722, new_n17723, new_n17724,
    new_n17725, new_n17726, new_n17727, new_n17728, new_n17729, new_n17730,
    new_n17731, new_n17732, new_n17733, new_n17734, new_n17735_1,
    new_n17736, new_n17737, new_n17738_1, new_n17739, new_n17740,
    new_n17741, new_n17742, new_n17743, new_n17744, new_n17745,
    new_n17746_1, new_n17747, new_n17748, new_n17749_1, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780,
    new_n17781, new_n17782, new_n17783, new_n17784_1, new_n17785,
    new_n17786, new_n17787, new_n17788, new_n17789, new_n17790, new_n17791,
    new_n17792, new_n17793, new_n17794, new_n17795, new_n17796, new_n17797,
    new_n17798, new_n17799, new_n17800, new_n17801, new_n17802, new_n17803,
    new_n17804, new_n17805, new_n17806, new_n17807, new_n17808, new_n17809,
    new_n17810, new_n17811, new_n17812, new_n17813, new_n17814, new_n17815,
    new_n17816, new_n17817, new_n17818, new_n17819, new_n17820_1,
    new_n17821, new_n17822, new_n17823, new_n17824, new_n17825, new_n17826,
    new_n17827, new_n17828, new_n17829, new_n17830, new_n17831, new_n17832,
    new_n17833, new_n17834, new_n17835, new_n17836, new_n17837, new_n17838,
    new_n17839, new_n17840, new_n17841, new_n17842, new_n17843, new_n17844,
    new_n17845, new_n17847, new_n17849, new_n17851, new_n17853, new_n17854,
    new_n17855_1, new_n17856, new_n17857, new_n17858, new_n17859,
    new_n17860, new_n17861, new_n17862, new_n17863, new_n17864, new_n17865,
    new_n17866, new_n17867, new_n17868, new_n17869, new_n17870, new_n17871,
    new_n17872, new_n17874, new_n17876, new_n17877_1, new_n17878,
    new_n17879, new_n17880, new_n17881, new_n17882, new_n17883, new_n17884,
    new_n17885, new_n17886, new_n17887, new_n17888, new_n17889_1,
    new_n17890, new_n17891, new_n17892, new_n17893, new_n17894, new_n17895,
    new_n17896, new_n17897, new_n17898, new_n17899, new_n17900, new_n17901,
    new_n17902, new_n17903, new_n17904, new_n17905, new_n17906, new_n17907,
    new_n17908, new_n17909, new_n17910, new_n17911_1, new_n17912_1,
    new_n17913, new_n17914, new_n17915, new_n17916, new_n17917, new_n17918,
    new_n17919, new_n17920, new_n17921, new_n17922, new_n17923, new_n17924,
    new_n17925, new_n17926, new_n17927_1, new_n17928, new_n17929,
    new_n17930, new_n17931_1, new_n17932, new_n17933, new_n17934,
    new_n17935, new_n17936, new_n17937, new_n17938, new_n17939, new_n17940,
    new_n17941, new_n17942, new_n17943, new_n17944, new_n17945, new_n17946,
    new_n17947, new_n17948_1, new_n17949, new_n17950, new_n17951,
    new_n17952, new_n17953, new_n17954_1, new_n17955, new_n17956_1,
    new_n17957, new_n17958, new_n17959_1, new_n17960, new_n17961,
    new_n17962, new_n17963_1, new_n17964, new_n17965, new_n17966,
    new_n17967, new_n17968_1, new_n17969, new_n17970, new_n17971,
    new_n17972, new_n17973, new_n17974, new_n17975, new_n17976_1,
    new_n17977, new_n17978, new_n17979, new_n17980, new_n17981, new_n17982,
    new_n17983, new_n17984, new_n17985, new_n17986, new_n17987, new_n17988,
    new_n17989, new_n17990, new_n17991, new_n17992, new_n17993, new_n17994,
    new_n17995, new_n17996, new_n17997, new_n17999, new_n18001, new_n18002,
    new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008,
    new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014,
    new_n18015, new_n18016, new_n18017, new_n18018, new_n18019, new_n18020,
    new_n18021, new_n18022, new_n18024, new_n18025_1, new_n18026,
    new_n18027, new_n18028, new_n18029, new_n18030, new_n18031, new_n18032,
    new_n18033, new_n18034, new_n18035_1, new_n18036, new_n18037,
    new_n18038, new_n18039, new_n18040, new_n18041, new_n18042,
    new_n18043_1, new_n18044, new_n18045_1, new_n18046, new_n18047,
    new_n18048, new_n18049, new_n18050, new_n18051, new_n18053, new_n18055,
    new_n18056, new_n18057, new_n18058, new_n18059_1, new_n18060,
    new_n18061_1, new_n18062, new_n18063, new_n18064, new_n18065,
    new_n18066, new_n18067, new_n18068, new_n18069, new_n18070,
    new_n18071_1, new_n18072, new_n18073, new_n18074, new_n18075,
    new_n18076, new_n18077, new_n18078, new_n18079, new_n18080, new_n18081,
    new_n18082, new_n18083, new_n18084, new_n18085, new_n18086, new_n18087,
    new_n18088, new_n18089, new_n18090, new_n18091, new_n18092, new_n18093,
    new_n18094, new_n18095, new_n18096, new_n18097, new_n18098, new_n18100,
    new_n18101, new_n18102, new_n18103, new_n18104, new_n18105_1,
    new_n18106, new_n18107, new_n18108, new_n18109, new_n18110, new_n18111,
    new_n18112, new_n18113, new_n18114, new_n18115, new_n18116, new_n18117,
    new_n18118, new_n18119, new_n18120, new_n18121, new_n18122, new_n18123,
    new_n18124, new_n18125, new_n18126, new_n18127, new_n18128, new_n18129,
    new_n18130, new_n18131, new_n18132, new_n18133, new_n18134, new_n18135,
    new_n18136, new_n18137, new_n18138, new_n18139, new_n18140, new_n18141,
    new_n18142, new_n18143_1, new_n18144, new_n18145_1, new_n18146,
    new_n18147, new_n18148, new_n18149, new_n18150, new_n18151_1,
    new_n18152_1, new_n18153, new_n18154, new_n18155, new_n18156,
    new_n18157_1, new_n18158, new_n18159, new_n18160, new_n18161,
    new_n18162, new_n18163, new_n18164, new_n18165, new_n18166, new_n18167,
    new_n18168, new_n18169, new_n18170, new_n18171_1, new_n18172,
    new_n18173, new_n18174, new_n18175, new_n18176, new_n18177, new_n18178,
    new_n18179, new_n18180, new_n18181, new_n18182, new_n18183, new_n18184,
    new_n18185, new_n18186, new_n18187, new_n18188, new_n18189, new_n18190,
    new_n18191, new_n18192, new_n18193_1, new_n18194, new_n18195,
    new_n18196, new_n18197, new_n18198, new_n18199, new_n18200, new_n18201,
    new_n18202, new_n18203, new_n18204, new_n18205, new_n18206, new_n18207,
    new_n18208, new_n18209, new_n18210, new_n18211, new_n18212, new_n18213,
    new_n18214, new_n18215, new_n18216, new_n18217, new_n18218, new_n18219,
    new_n18220, new_n18221, new_n18222, new_n18223, new_n18224, new_n18225,
    new_n18226, new_n18227_1, new_n18228, new_n18229, new_n18230,
    new_n18231, new_n18232_1, new_n18233, new_n18234, new_n18235,
    new_n18236, new_n18237, new_n18238_1, new_n18239, new_n18240,
    new_n18241_1, new_n18242, new_n18243, new_n18244, new_n18245,
    new_n18246, new_n18247, new_n18248, new_n18249, new_n18250, new_n18251,
    new_n18252, new_n18253, new_n18254_1, new_n18255, new_n18256,
    new_n18257, new_n18258, new_n18259, new_n18260, new_n18261, new_n18262,
    new_n18263, new_n18264, new_n18265, new_n18266, new_n18267, new_n18268,
    new_n18269, new_n18270, new_n18271, new_n18272, new_n18273,
    new_n18274_1, new_n18275, new_n18276, new_n18277, new_n18278,
    new_n18279, new_n18280, new_n18281, new_n18282, new_n18283, new_n18284,
    new_n18285, new_n18286, new_n18287, new_n18288_1, new_n18289,
    new_n18290_1, new_n18291, new_n18292, new_n18293, new_n18294,
    new_n18295_1, new_n18296, new_n18297, new_n18298, new_n18299,
    new_n18300, new_n18301_1, new_n18302, new_n18303, new_n18304_1,
    new_n18305, new_n18306, new_n18307, new_n18308, new_n18309,
    new_n18310_1, new_n18311_1, new_n18313, new_n18314, new_n18315,
    new_n18316, new_n18317, new_n18318, new_n18319, new_n18320, new_n18321,
    new_n18322, new_n18323_1, new_n18324, new_n18325, new_n18326,
    new_n18327, new_n18328, new_n18329, new_n18330, new_n18331,
    new_n18332_1, new_n18333, new_n18334, new_n18335, new_n18336,
    new_n18337, new_n18338, new_n18339, new_n18340, new_n18341, new_n18342,
    new_n18343_1, new_n18344, new_n18345_1, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18350_1, new_n18351, new_n18352,
    new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358,
    new_n18359, new_n18360, new_n18361, new_n18362_1, new_n18363,
    new_n18364, new_n18365, new_n18366, new_n18367, new_n18368, new_n18369,
    new_n18370, new_n18371, new_n18372, new_n18373, new_n18374, new_n18375,
    new_n18376, new_n18377_1, new_n18378, new_n18379, new_n18380,
    new_n18381, new_n18382, new_n18383, new_n18384, new_n18385, new_n18386,
    new_n18387, new_n18388, new_n18389, new_n18390, new_n18391, new_n18392,
    new_n18393, new_n18394, new_n18395, new_n18396, new_n18397, new_n18398,
    new_n18399, new_n18400, new_n18401, new_n18402, new_n18403, new_n18404,
    new_n18405_1, new_n18406, new_n18407, new_n18408, new_n18409_1,
    new_n18410, new_n18411, new_n18412, new_n18413, new_n18414_1,
    new_n18415, new_n18416, new_n18417, new_n18418_1, new_n18419,
    new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425,
    new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431,
    new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437_1, new_n18438, new_n18439_1, new_n18442, new_n18443,
    new_n18444_1, new_n18445_1, new_n18446, new_n18447, new_n18448,
    new_n18449, new_n18450, new_n18451, new_n18452_1, new_n18453,
    new_n18454, new_n18455, new_n18456, new_n18457, new_n18458, new_n18459,
    new_n18460, new_n18461, new_n18462, new_n18463, new_n18464, new_n18465,
    new_n18466, new_n18467_1, new_n18468, new_n18469, new_n18470,
    new_n18471, new_n18472, new_n18473, new_n18474, new_n18475, new_n18476,
    new_n18477, new_n18478, new_n18479, new_n18480, new_n18481,
    new_n18482_1, new_n18483_1, new_n18484, new_n18485, new_n18486,
    new_n18487, new_n18488, new_n18489, new_n18490, new_n18491, new_n18492,
    new_n18493, new_n18494, new_n18495, new_n18496_1, new_n18497,
    new_n18498, new_n18499, new_n18500, new_n18501, new_n18502, new_n18503,
    new_n18504, new_n18505, new_n18506, new_n18507, new_n18508,
    new_n18509_1, new_n18510, new_n18511, new_n18512, new_n18513_1,
    new_n18514, new_n18515_1, new_n18516, new_n18517, new_n18518,
    new_n18519, new_n18520, new_n18521, new_n18522, new_n18523, new_n18524,
    new_n18525, new_n18526, new_n18527, new_n18528, new_n18529, new_n18530,
    new_n18531, new_n18532, new_n18533, new_n18534, new_n18535, new_n18536,
    new_n18537_1, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18555, new_n18556, new_n18557, new_n18558_1,
    new_n18559, new_n18560, new_n18561, new_n18562, new_n18563, new_n18564,
    new_n18565, new_n18566, new_n18567, new_n18568, new_n18569, new_n18570,
    new_n18571, new_n18572_1, new_n18573, new_n18575, new_n18576_1,
    new_n18577, new_n18578_1, new_n18579, new_n18580, new_n18581,
    new_n18582_1, new_n18583_1, new_n18584_1, new_n18585, new_n18586,
    new_n18587, new_n18588, new_n18589, new_n18590, new_n18591, new_n18592,
    new_n18593, new_n18594, new_n18595, new_n18596, new_n18597, new_n18598,
    new_n18599, new_n18600, new_n18601, new_n18602, new_n18603, new_n18604,
    new_n18605, new_n18606, new_n18607, new_n18608, new_n18609,
    new_n18610_1, new_n18611, new_n18612, new_n18613, new_n18614,
    new_n18615, new_n18616, new_n18617, new_n18618, new_n18619, new_n18620,
    new_n18621, new_n18622, new_n18623, new_n18624, new_n18625, new_n18626,
    new_n18627, new_n18628, new_n18630, new_n18631, new_n18632, new_n18633,
    new_n18634, new_n18635_1, new_n18636, new_n18637, new_n18638,
    new_n18639, new_n18640, new_n18641, new_n18642, new_n18643, new_n18644,
    new_n18645, new_n18646, new_n18647, new_n18648, new_n18649_1,
    new_n18650, new_n18651, new_n18653_1, new_n18655, new_n18656,
    new_n18657, new_n18658, new_n18659, new_n18660, new_n18661, new_n18662,
    new_n18663, new_n18664, new_n18665, new_n18666, new_n18667, new_n18668,
    new_n18669, new_n18670, new_n18671, new_n18672, new_n18673, new_n18674,
    new_n18675, new_n18676, new_n18677, new_n18678, new_n18679_1,
    new_n18680, new_n18681, new_n18682, new_n18683, new_n18684, new_n18685,
    new_n18686, new_n18687, new_n18688, new_n18689, new_n18690_1,
    new_n18691, new_n18692, new_n18693_1, new_n18694, new_n18695,
    new_n18696, new_n18697, new_n18698, new_n18699, new_n18700, new_n18701,
    new_n18702, new_n18703, new_n18704, new_n18705, new_n18706, new_n18707,
    new_n18708_1, new_n18709, new_n18710, new_n18711, new_n18712,
    new_n18713, new_n18714, new_n18715, new_n18716, new_n18717, new_n18718,
    new_n18719, new_n18720, new_n18721_1, new_n18722, new_n18723,
    new_n18724, new_n18725_1, new_n18726, new_n18727, new_n18728,
    new_n18729, new_n18730, new_n18731, new_n18732, new_n18733, new_n18735,
    new_n18737_1, new_n18739, new_n18740, new_n18741, new_n18742,
    new_n18743, new_n18744, new_n18745_1, new_n18746, new_n18747,
    new_n18748, new_n18749, new_n18751_1, new_n18753, new_n18755,
    new_n18756, new_n18757, new_n18758, new_n18759, new_n18760, new_n18761,
    new_n18762, new_n18763, new_n18764, new_n18765, new_n18766, new_n18767,
    new_n18768, new_n18769, new_n18770, new_n18771, new_n18772, new_n18773,
    new_n18774, new_n18775, new_n18776, new_n18777, new_n18778, new_n18779,
    new_n18780_1, new_n18781, new_n18782_1, new_n18783, new_n18784,
    new_n18785, new_n18786, new_n18787, new_n18788, new_n18789, new_n18790,
    new_n18791, new_n18793, new_n18795, new_n18796, new_n18797, new_n18798,
    new_n18799, new_n18800, new_n18801, new_n18802_1, new_n18803,
    new_n18804, new_n18805, new_n18806, new_n18807, new_n18808, new_n18809,
    new_n18810, new_n18811, new_n18812, new_n18813, new_n18814, new_n18815,
    new_n18816, new_n18817, new_n18818, new_n18819, new_n18820, new_n18821,
    new_n18822, new_n18823, new_n18824, new_n18825, new_n18826, new_n18827,
    new_n18828, new_n18829, new_n18830_1, new_n18831_1, new_n18832,
    new_n18833, new_n18834, new_n18835, new_n18836, new_n18837, new_n18838,
    new_n18839, new_n18840, new_n18841, new_n18842, new_n18843_1,
    new_n18844, new_n18845, new_n18846, new_n18847, new_n18848, new_n18849,
    new_n18850, new_n18851, new_n18852, new_n18853, new_n18854, new_n18855,
    new_n18856, new_n18857, new_n18858_1, new_n18859_1, new_n18860,
    new_n18861, new_n18862, new_n18863, new_n18864_1, new_n18865_1,
    new_n18866, new_n18867, new_n18868, new_n18869, new_n18870, new_n18871,
    new_n18872, new_n18873, new_n18874, new_n18875, new_n18876, new_n18877,
    new_n18878, new_n18879, new_n18880_1, new_n18881, new_n18882,
    new_n18883, new_n18884, new_n18885, new_n18886_1, new_n18887_1,
    new_n18888, new_n18889, new_n18890, new_n18891, new_n18892, new_n18893,
    new_n18894, new_n18895, new_n18896, new_n18897, new_n18898, new_n18899,
    new_n18900, new_n18901_1, new_n18902, new_n18903, new_n18904,
    new_n18905, new_n18906, new_n18907_1, new_n18908, new_n18909,
    new_n18910, new_n18911, new_n18912, new_n18913, new_n18914, new_n18915,
    new_n18916, new_n18917, new_n18918, new_n18919_1, new_n18921,
    new_n18923, new_n18925, new_n18926_1, new_n18927, new_n18928,
    new_n18929, new_n18930, new_n18931, new_n18932, new_n18933, new_n18934,
    new_n18935, new_n18936, new_n18937, new_n18938, new_n18939,
    new_n18940_1, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945_1, new_n18946, new_n18947, new_n18948, new_n18949,
    new_n18950, new_n18951, new_n18952, new_n18953, new_n18954, new_n18955,
    new_n18956, new_n18957, new_n18958, new_n18959, new_n18960, new_n18961,
    new_n18962_1, new_n18963, new_n18964, new_n18965, new_n18966,
    new_n18967, new_n18968, new_n18969, new_n18970_1, new_n18971,
    new_n18972, new_n18973, new_n18974, new_n18975, new_n18976,
    new_n18977_1, new_n18978, new_n18979, new_n18980, new_n18981,
    new_n18982_1, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999_1, new_n19000, new_n19001, new_n19002, new_n19003,
    new_n19004, new_n19005_1, new_n19006, new_n19007, new_n19008,
    new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014,
    new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020,
    new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026,
    new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032,
    new_n19033_1, new_n19034, new_n19035, new_n19036, new_n19037,
    new_n19038, new_n19039, new_n19040, new_n19041, new_n19042_1,
    new_n19043, new_n19044_1, new_n19045, new_n19046, new_n19047,
    new_n19048, new_n19049, new_n19050, new_n19051, new_n19052, new_n19053,
    new_n19054, new_n19055, new_n19056, new_n19057, new_n19058, new_n19059,
    new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19065,
    new_n19066, new_n19067, new_n19068, new_n19069, new_n19070, new_n19071,
    new_n19072, new_n19073, new_n19074, new_n19075, new_n19076, new_n19077,
    new_n19078, new_n19079, new_n19080, new_n19081_1, new_n19083,
    new_n19084, new_n19085, new_n19086, new_n19087, new_n19088, new_n19089,
    new_n19090, new_n19091, new_n19092, new_n19093, new_n19094, new_n19095,
    new_n19096, new_n19097, new_n19098, new_n19099, new_n19100, new_n19101,
    new_n19102, new_n19103, new_n19105, new_n19106, new_n19107_1,
    new_n19108, new_n19109, new_n19110, new_n19111, new_n19112, new_n19113,
    new_n19114, new_n19115, new_n19116_1, new_n19117, new_n19118,
    new_n19119, new_n19120, new_n19121, new_n19122, new_n19123, new_n19124,
    new_n19125_1, new_n19126, new_n19127, new_n19128, new_n19129,
    new_n19130, new_n19131, new_n19132, new_n19133, new_n19134, new_n19135,
    new_n19136, new_n19137, new_n19138, new_n19139, new_n19140,
    new_n19141_1, new_n19142, new_n19143, new_n19144_1, new_n19145,
    new_n19146, new_n19147, new_n19149, new_n19150, new_n19151, new_n19152,
    new_n19153, new_n19154, new_n19155, new_n19156, new_n19157, new_n19158,
    new_n19159, new_n19160, new_n19161, new_n19162, new_n19163_1,
    new_n19164_1, new_n19165, new_n19166, new_n19167, new_n19168,
    new_n19169, new_n19170, new_n19171, new_n19172, new_n19173,
    new_n19174_1, new_n19175, new_n19176_1, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19191,
    new_n19192, new_n19193, new_n19194, new_n19195, new_n19196_1,
    new_n19197, new_n19198, new_n19199, new_n19200, new_n19201,
    new_n19202_1, new_n19203, new_n19204, new_n19205, new_n19206,
    new_n19207, new_n19208, new_n19209, new_n19210, new_n19211, new_n19212,
    new_n19213, new_n19214, new_n19215, new_n19216, new_n19217, new_n19218,
    new_n19219, new_n19220_1, new_n19221_1, new_n19222, new_n19223_1,
    new_n19224_1, new_n19225, new_n19227, new_n19229, new_n19230,
    new_n19231, new_n19232, new_n19233_1, new_n19234_1, new_n19235,
    new_n19236, new_n19237, new_n19238, new_n19239, new_n19240, new_n19241,
    new_n19242, new_n19243, new_n19244_1, new_n19245, new_n19246,
    new_n19247, new_n19248, new_n19249, new_n19251, new_n19252, new_n19253,
    new_n19254, new_n19255, new_n19256, new_n19257, new_n19258, new_n19259,
    new_n19260, new_n19261, new_n19262, new_n19263, new_n19264, new_n19265,
    new_n19266, new_n19267, new_n19268, new_n19269, new_n19270_1,
    new_n19271, new_n19272, new_n19273, new_n19274, new_n19275, new_n19276,
    new_n19277, new_n19278, new_n19279, new_n19280, new_n19281,
    new_n19282_1, new_n19283, new_n19284, new_n19285, new_n19286,
    new_n19287, new_n19288, new_n19289, new_n19290, new_n19291, new_n19292,
    new_n19293, new_n19294, new_n19295, new_n19296, new_n19297, new_n19298,
    new_n19299, new_n19300, new_n19301, new_n19302, new_n19303, new_n19304,
    new_n19305, new_n19306, new_n19307, new_n19308, new_n19309, new_n19310,
    new_n19311, new_n19312, new_n19313, new_n19314_1, new_n19315_1,
    new_n19316, new_n19317, new_n19318, new_n19319, new_n19320, new_n19321,
    new_n19322, new_n19323_1, new_n19324, new_n19325, new_n19326,
    new_n19327_1, new_n19329, new_n19330, new_n19331, new_n19332,
    new_n19333_1, new_n19334, new_n19335, new_n19336, new_n19337,
    new_n19338, new_n19339, new_n19340, new_n19341, new_n19342, new_n19343,
    new_n19344, new_n19345, new_n19346, new_n19347, new_n19348_1,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353,
    new_n19354_1, new_n19355, new_n19356, new_n19357_1, new_n19358,
    new_n19359, new_n19360, new_n19361_1, new_n19362, new_n19363,
    new_n19364, new_n19365, new_n19366, new_n19367_1, new_n19368,
    new_n19369, new_n19370, new_n19371, new_n19372, new_n19373, new_n19374,
    new_n19375, new_n19376, new_n19377, new_n19378, new_n19379, new_n19380,
    new_n19381, new_n19382, new_n19383, new_n19384, new_n19385_1,
    new_n19386, new_n19387, new_n19388, new_n19389_1, new_n19390,
    new_n19391, new_n19392, new_n19393, new_n19394, new_n19395, new_n19396,
    new_n19397, new_n19398, new_n19399, new_n19400, new_n19401_1,
    new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407,
    new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414_1, new_n19415, new_n19416, new_n19417, new_n19418,
    new_n19419, new_n19420, new_n19421, new_n19422, new_n19423,
    new_n19424_1, new_n19425, new_n19426, new_n19427, new_n19428,
    new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434,
    new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440,
    new_n19441, new_n19442, new_n19443, new_n19444, new_n19445, new_n19446,
    new_n19447, new_n19448, new_n19449, new_n19450_1, new_n19451,
    new_n19452, new_n19453, new_n19454_1, new_n19455, new_n19456,
    new_n19457, new_n19458_1, new_n19459, new_n19460, new_n19461,
    new_n19462, new_n19463, new_n19464, new_n19465, new_n19466,
    new_n19467_1, new_n19468, new_n19469, new_n19470, new_n19471,
    new_n19472_1, new_n19473, new_n19474, new_n19475, new_n19476,
    new_n19477_1, new_n19478, new_n19479, new_n19480, new_n19481,
    new_n19482, new_n19483, new_n19484, new_n19485, new_n19486, new_n19487,
    new_n19488, new_n19489, new_n19490, new_n19491, new_n19492, new_n19493,
    new_n19494_1, new_n19495, new_n19496_1, new_n19497, new_n19498,
    new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504,
    new_n19505, new_n19506, new_n19507, new_n19508, new_n19509, new_n19510,
    new_n19511, new_n19512, new_n19513, new_n19515_1, new_n19516,
    new_n19517, new_n19518, new_n19519, new_n19520, new_n19521, new_n19522,
    new_n19523_1, new_n19524, new_n19525, new_n19526, new_n19527,
    new_n19528, new_n19529, new_n19530, new_n19532, new_n19534, new_n19535,
    new_n19536, new_n19537, new_n19538, new_n19539_1, new_n19540,
    new_n19541, new_n19542, new_n19543, new_n19544, new_n19545, new_n19547,
    new_n19549, new_n19551, new_n19553, new_n19554, new_n19555, new_n19556,
    new_n19557, new_n19558, new_n19559, new_n19560, new_n19561, new_n19562,
    new_n19564, new_n19566, new_n19568, new_n19570_1, new_n19572,
    new_n19574, new_n19575_1, new_n19576, new_n19577, new_n19578,
    new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584_1, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602_1, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608_1, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617_1, new_n19618_1, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623_1, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641_1, new_n19642, new_n19643,
    new_n19644, new_n19645, new_n19646, new_n19647, new_n19648_1,
    new_n19649, new_n19650, new_n19651, new_n19652_1, new_n19653,
    new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659,
    new_n19660, new_n19661, new_n19662, new_n19663, new_n19664_1,
    new_n19665, new_n19666, new_n19667, new_n19668, new_n19669, new_n19670,
    new_n19671, new_n19672, new_n19673, new_n19674, new_n19675, new_n19677,
    new_n19678, new_n19679, new_n19680_1, new_n19681, new_n19682,
    new_n19683, new_n19684, new_n19685, new_n19686, new_n19687, new_n19688,
    new_n19689, new_n19690, new_n19691, new_n19692, new_n19693, new_n19694,
    new_n19695, new_n19696, new_n19697, new_n19698, new_n19699, new_n19700,
    new_n19701_1, new_n19702, new_n19703, new_n19704, new_n19705,
    new_n19706, new_n19707, new_n19708, new_n19709, new_n19710, new_n19711,
    new_n19712, new_n19713, new_n19714, new_n19715, new_n19716, new_n19717,
    new_n19718, new_n19719, new_n19720, new_n19721, new_n19722, new_n19723,
    new_n19724, new_n19725, new_n19726, new_n19727, new_n19729, new_n19730,
    new_n19731, new_n19732, new_n19733, new_n19734, new_n19735,
    new_n19736_1, new_n19737, new_n19738, new_n19739, new_n19740,
    new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746,
    new_n19747, new_n19748, new_n19749_1, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756_1,
    new_n19757, new_n19758, new_n19759, new_n19760, new_n19761, new_n19762,
    new_n19763, new_n19764, new_n19765, new_n19766, new_n19767_1,
    new_n19768, new_n19769, new_n19770_1, new_n19771, new_n19772,
    new_n19773, new_n19774, new_n19775, new_n19776, new_n19777, new_n19778,
    new_n19779, new_n19780_1, new_n19781, new_n19782, new_n19783,
    new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789_1, new_n19790, new_n19791, new_n19792_1, new_n19793,
    new_n19794, new_n19795, new_n19796, new_n19797, new_n19798_1,
    new_n19799, new_n19800, new_n19801, new_n19802, new_n19803_1,
    new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809,
    new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815,
    new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821,
    new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827,
    new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833,
    new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839,
    new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845,
    new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851,
    new_n19852, new_n19853, new_n19854, new_n19855, new_n19856, new_n19857,
    new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863,
    new_n19864, new_n19865, new_n19866, new_n19867, new_n19868, new_n19869,
    new_n19870, new_n19871, new_n19872, new_n19873_1, new_n19874,
    new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19880,
    new_n19881, new_n19882, new_n19883, new_n19884, new_n19885, new_n19886,
    new_n19887, new_n19888, new_n19889, new_n19890, new_n19891, new_n19892,
    new_n19893, new_n19894, new_n19895, new_n19896, new_n19897, new_n19898,
    new_n19899, new_n19900, new_n19901, new_n19903, new_n19904,
    new_n19905_1, new_n19906, new_n19907, new_n19908, new_n19909_1,
    new_n19910, new_n19911_1, new_n19912, new_n19913, new_n19914,
    new_n19915, new_n19916_1, new_n19917, new_n19918, new_n19919,
    new_n19920, new_n19921, new_n19922_1, new_n19923_1, new_n19924,
    new_n19925, new_n19926, new_n19927, new_n19928, new_n19929,
    new_n19930_1, new_n19931, new_n19932, new_n19933, new_n19934,
    new_n19935, new_n19936, new_n19937, new_n19938, new_n19939, new_n19940,
    new_n19941_1, new_n19942, new_n19943, new_n19944, new_n19945,
    new_n19946, new_n19947, new_n19948, new_n19949, new_n19950, new_n19951,
    new_n19953, new_n19955, new_n19956, new_n19957, new_n19958, new_n19959,
    new_n19960, new_n19961, new_n19962, new_n19963, new_n19964, new_n19965,
    new_n19966, new_n19967, new_n19968_1, new_n19969, new_n19970,
    new_n19971, new_n19972, new_n19974, new_n19976, new_n19977, new_n19978,
    new_n19979, new_n19980, new_n19981, new_n19982, new_n19983, new_n19984,
    new_n19985, new_n19986, new_n19987, new_n19988_1, new_n19990,
    new_n19992, new_n19994, new_n19995, new_n19996, new_n19997, new_n19998,
    new_n19999, new_n20000, new_n20001, new_n20002, new_n20003,
    new_n20004_1, new_n20005, new_n20006, new_n20007, new_n20008,
    new_n20009, new_n20010, new_n20011, new_n20012, new_n20013_1,
    new_n20014, new_n20015, new_n20016, new_n20017_1, new_n20018,
    new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024,
    new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030,
    new_n20031, new_n20032, new_n20033_1, new_n20034, new_n20035,
    new_n20036_1, new_n20037, new_n20038, new_n20039, new_n20040_1,
    new_n20041, new_n20043, new_n20045, new_n20046, new_n20047, new_n20048,
    new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061_1, new_n20062, new_n20063, new_n20064, new_n20065,
    new_n20066, new_n20067, new_n20068, new_n20069_1, new_n20070,
    new_n20071, new_n20072, new_n20073, new_n20074, new_n20075, new_n20076,
    new_n20077_1, new_n20078, new_n20079, new_n20080, new_n20081,
    new_n20082, new_n20083, new_n20084, new_n20085, new_n20086_1,
    new_n20087, new_n20088, new_n20089, new_n20090, new_n20091, new_n20092,
    new_n20093, new_n20094, new_n20095, new_n20096_1, new_n20097,
    new_n20098, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103_1, new_n20104, new_n20105, new_n20106, new_n20107,
    new_n20108, new_n20109, new_n20110, new_n20111, new_n20112, new_n20113,
    new_n20114, new_n20115, new_n20116, new_n20117, new_n20118, new_n20119,
    new_n20120, new_n20121, new_n20122, new_n20123, new_n20124, new_n20125,
    new_n20126_1, new_n20127, new_n20128, new_n20129, new_n20130,
    new_n20131, new_n20132, new_n20133, new_n20134, new_n20135, new_n20137,
    new_n20138_1, new_n20139, new_n20140, new_n20141, new_n20142,
    new_n20143, new_n20144, new_n20145, new_n20146, new_n20147, new_n20148,
    new_n20149_1, new_n20150, new_n20151_1, new_n20152, new_n20153,
    new_n20154, new_n20155, new_n20156, new_n20157, new_n20158, new_n20159,
    new_n20160, new_n20161, new_n20162, new_n20163, new_n20164, new_n20165,
    new_n20166, new_n20167, new_n20168, new_n20169_1, new_n20170,
    new_n20171, new_n20172, new_n20173, new_n20174, new_n20175, new_n20176,
    new_n20177, new_n20178, new_n20179_1, new_n20180, new_n20181,
    new_n20183, new_n20184, new_n20185, new_n20186, new_n20187_1,
    new_n20188, new_n20189, new_n20190, new_n20191, new_n20192, new_n20193,
    new_n20194, new_n20195, new_n20196, new_n20197, new_n20198, new_n20199,
    new_n20200, new_n20201, new_n20202, new_n20203, new_n20204, new_n20205,
    new_n20206, new_n20207, new_n20208, new_n20209, new_n20210, new_n20211,
    new_n20212, new_n20213_1, new_n20214, new_n20215, new_n20216,
    new_n20217, new_n20218, new_n20219, new_n20220, new_n20221, new_n20222,
    new_n20223, new_n20224, new_n20225, new_n20226, new_n20227, new_n20228,
    new_n20229, new_n20230, new_n20231, new_n20232, new_n20233, new_n20234,
    new_n20235_1, new_n20236, new_n20237, new_n20238, new_n20239,
    new_n20240, new_n20241, new_n20242, new_n20244, new_n20246, new_n20248,
    new_n20249, new_n20251, new_n20253, new_n20254, new_n20255, new_n20256,
    new_n20257, new_n20258, new_n20259_1, new_n20260, new_n20261,
    new_n20262, new_n20263, new_n20264, new_n20265, new_n20266, new_n20267,
    new_n20268, new_n20269, new_n20270, new_n20271, new_n20272, new_n20273,
    new_n20274, new_n20275, new_n20276, new_n20277, new_n20278,
    new_n20279_1, new_n20280, new_n20281, new_n20282, new_n20283,
    new_n20284, new_n20285, new_n20286, new_n20287_1, new_n20288,
    new_n20289, new_n20290, new_n20291, new_n20292, new_n20293, new_n20294,
    new_n20295, new_n20296, new_n20297, new_n20298, new_n20299, new_n20300,
    new_n20301_1, new_n20302, new_n20303, new_n20304, new_n20305,
    new_n20306, new_n20307, new_n20308, new_n20309, new_n20310, new_n20311,
    new_n20312, new_n20313, new_n20314, new_n20315, new_n20316, new_n20317,
    new_n20318, new_n20320, new_n20322, new_n20323, new_n20324, new_n20325,
    new_n20326, new_n20327, new_n20328, new_n20329, new_n20330_1,
    new_n20331, new_n20332, new_n20333_1, new_n20334, new_n20335,
    new_n20336, new_n20337, new_n20338, new_n20339, new_n20340, new_n20341,
    new_n20342, new_n20343, new_n20344, new_n20345, new_n20346, new_n20347,
    new_n20348, new_n20349_1, new_n20350, new_n20351, new_n20352,
    new_n20353, new_n20354, new_n20355_1, new_n20356, new_n20358,
    new_n20360, new_n20361, new_n20362, new_n20363, new_n20364, new_n20365,
    new_n20366_1, new_n20367, new_n20368, new_n20369, new_n20370,
    new_n20371, new_n20372, new_n20373, new_n20374, new_n20375, new_n20376,
    new_n20377, new_n20379, new_n20380, new_n20381, new_n20382, new_n20384,
    new_n20386, new_n20389, new_n20390, new_n20391, new_n20392, new_n20393,
    new_n20394, new_n20395, new_n20396, new_n20397, new_n20398, new_n20399,
    new_n20400, new_n20401, new_n20402_1, new_n20403_1, new_n20404,
    new_n20405, new_n20406, new_n20407, new_n20408, new_n20409_1,
    new_n20410, new_n20411_1, new_n20412, new_n20413, new_n20414,
    new_n20415, new_n20416, new_n20417, new_n20418, new_n20419, new_n20420,
    new_n20421, new_n20422, new_n20423, new_n20424_1, new_n20425,
    new_n20426, new_n20427, new_n20428, new_n20429_1, new_n20430,
    new_n20431, new_n20432, new_n20433, new_n20434, new_n20435,
    new_n20436_1, new_n20437, new_n20438, new_n20439, new_n20440,
    new_n20441_1, new_n20442, new_n20443, new_n20444, new_n20445_1,
    new_n20446, new_n20447, new_n20448, new_n20449, new_n20450_1,
    new_n20451, new_n20452, new_n20453, new_n20454, new_n20455_1,
    new_n20456, new_n20457, new_n20458, new_n20459, new_n20460, new_n20461,
    new_n20462, new_n20463, new_n20464, new_n20465, new_n20466, new_n20467,
    new_n20468, new_n20469, new_n20470_1, new_n20471, new_n20472,
    new_n20473, new_n20474, new_n20475, new_n20476, new_n20477,
    new_n20478_1, new_n20479, new_n20480, new_n20481, new_n20482,
    new_n20483, new_n20484, new_n20485, new_n20486, new_n20487, new_n20488,
    new_n20489_1, new_n20490_1, new_n20491, new_n20492, new_n20493,
    new_n20494, new_n20495_1, new_n20496, new_n20497, new_n20498,
    new_n20499, new_n20500, new_n20501, new_n20502, new_n20503, new_n20504,
    new_n20505, new_n20506, new_n20507, new_n20508, new_n20509, new_n20510,
    new_n20511, new_n20512, new_n20513, new_n20514, new_n20515_1,
    new_n20516, new_n20517, new_n20518, new_n20519, new_n20520, new_n20521,
    new_n20522, new_n20523, new_n20524, new_n20526, new_n20528, new_n20530,
    new_n20531, new_n20532, new_n20533_1, new_n20534, new_n20535,
    new_n20536, new_n20537, new_n20538, new_n20539, new_n20540, new_n20541,
    new_n20542, new_n20543, new_n20544, new_n20545, new_n20546, new_n20547,
    new_n20548, new_n20549, new_n20551, new_n20553, new_n20555, new_n20557,
    new_n20559, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565,
    new_n20566, new_n20567, new_n20568, new_n20569, new_n20570, new_n20571,
    new_n20572, new_n20573, new_n20574, new_n20575, new_n20576, new_n20577,
    new_n20578, new_n20579, new_n20580, new_n20581, new_n20582_1,
    new_n20583, new_n20584, new_n20585, new_n20586, new_n20587, new_n20588,
    new_n20589, new_n20590_1, new_n20591, new_n20592, new_n20593,
    new_n20594, new_n20595, new_n20596, new_n20597, new_n20598, new_n20599,
    new_n20600, new_n20601, new_n20602_1, new_n20603, new_n20604_1,
    new_n20605, new_n20606, new_n20607, new_n20608, new_n20609_1,
    new_n20610, new_n20611, new_n20612, new_n20613, new_n20614, new_n20615,
    new_n20616, new_n20617, new_n20618, new_n20619, new_n20620, new_n20621,
    new_n20622, new_n20623_1, new_n20624, new_n20625, new_n20626,
    new_n20627, new_n20628, new_n20629_1, new_n20630, new_n20631,
    new_n20632, new_n20633, new_n20634, new_n20635, new_n20636, new_n20637,
    new_n20638, new_n20639, new_n20641, new_n20643, new_n20644, new_n20645,
    new_n20646, new_n20647, new_n20648, new_n20649, new_n20650, new_n20651,
    new_n20652, new_n20653, new_n20654, new_n20655, new_n20656, new_n20657,
    new_n20658_1, new_n20659, new_n20660, new_n20661_1, new_n20662,
    new_n20663, new_n20664, new_n20665, new_n20666, new_n20667, new_n20668,
    new_n20669, new_n20670, new_n20671, new_n20672, new_n20673_1,
    new_n20674, new_n20675, new_n20676, new_n20677, new_n20678_1,
    new_n20679, new_n20680_1, new_n20681, new_n20682, new_n20683,
    new_n20684, new_n20685_1, new_n20686, new_n20687, new_n20688,
    new_n20689, new_n20690, new_n20691_1, new_n20692, new_n20693,
    new_n20694, new_n20695, new_n20696_1, new_n20697, new_n20698,
    new_n20699, new_n20700_1, new_n20701, new_n20702, new_n20703,
    new_n20704_1, new_n20705_1, new_n20706, new_n20707, new_n20708,
    new_n20709_1, new_n20710, new_n20711, new_n20712, new_n20713_1,
    new_n20714, new_n20715, new_n20716, new_n20717, new_n20718, new_n20719,
    new_n20720, new_n20721, new_n20722_1, new_n20723_1, new_n20725,
    new_n20726, new_n20727, new_n20728, new_n20729, new_n20730, new_n20731,
    new_n20732, new_n20733, new_n20734, new_n20735, new_n20736, new_n20737,
    new_n20738, new_n20739, new_n20740, new_n20741, new_n20742, new_n20743,
    new_n20744, new_n20745, new_n20746, new_n20747, new_n20748_1,
    new_n20749, new_n20750, new_n20751, new_n20752, new_n20753, new_n20754,
    new_n20755, new_n20756, new_n20757, new_n20758, new_n20759, new_n20760,
    new_n20761_1, new_n20762, new_n20763, new_n20764, new_n20765,
    new_n20766, new_n20767, new_n20768, new_n20769, new_n20770, new_n20771,
    new_n20772, new_n20773, new_n20774_1, new_n20776, new_n20777,
    new_n20778, new_n20779, new_n20780, new_n20781, new_n20782, new_n20783,
    new_n20784, new_n20785, new_n20786, new_n20787, new_n20788_1,
    new_n20789, new_n20790, new_n20791, new_n20792, new_n20793,
    new_n20794_1, new_n20795_1, new_n20796, new_n20797, new_n20798,
    new_n20799, new_n20800, new_n20801, new_n20802, new_n20803_1,
    new_n20804, new_n20805, new_n20806, new_n20807, new_n20808, new_n20809,
    new_n20810, new_n20811, new_n20812, new_n20813, new_n20814, new_n20815,
    new_n20816, new_n20817, new_n20818, new_n20819, new_n20820, new_n20821,
    new_n20822, new_n20823, new_n20824, new_n20825, new_n20826_1,
    new_n20827, new_n20828, new_n20829, new_n20830, new_n20831, new_n20832,
    new_n20833, new_n20835, new_n20838, new_n20840, new_n20841, new_n20842,
    new_n20843, new_n20844, new_n20845, new_n20846, new_n20847, new_n20848,
    new_n20849, new_n20850, new_n20851, new_n20852, new_n20853, new_n20854,
    new_n20855, new_n20856, new_n20857, new_n20858, new_n20859, new_n20860,
    new_n20861, new_n20862, new_n20863, new_n20864, new_n20865, new_n20866,
    new_n20869_1, new_n20871, new_n20873, new_n20874, new_n20875,
    new_n20876, new_n20877, new_n20878, new_n20879_1, new_n20880,
    new_n20881, new_n20882, new_n20883, new_n20884, new_n20885, new_n20886,
    new_n20887, new_n20888, new_n20889, new_n20890, new_n20891, new_n20892,
    new_n20893, new_n20894, new_n20895, new_n20896, new_n20897, new_n20898,
    new_n20899, new_n20900, new_n20901, new_n20902, new_n20903, new_n20904,
    new_n20905, new_n20906, new_n20907, new_n20908, new_n20909, new_n20910,
    new_n20911, new_n20912, new_n20913, new_n20914, new_n20915_1,
    new_n20916, new_n20917, new_n20918, new_n20919, new_n20920, new_n20921,
    new_n20922, new_n20923_1, new_n20925, new_n20926, new_n20928,
    new_n20929_1, new_n20930, new_n20931, new_n20932, new_n20933,
    new_n20934, new_n20935_1, new_n20936_1, new_n20937, new_n20938,
    new_n20939, new_n20941, new_n20943, new_n20945, new_n20946_1,
    new_n20947, new_n20948, new_n20949, new_n20950, new_n20951, new_n20952,
    new_n20953, new_n20954, new_n20955, new_n20956, new_n20957, new_n20958,
    new_n20959, new_n20960, new_n20961, new_n20962, new_n20963, new_n20964,
    new_n20965, new_n20966, new_n20967, new_n20968, new_n20969, new_n20971,
    new_n20972, new_n20973, new_n20974, new_n20975, new_n20976, new_n20977,
    new_n20978, new_n20979, new_n20980, new_n20981, new_n20982, new_n20983,
    new_n20984, new_n20985, new_n20986_1, new_n20987, new_n20988,
    new_n20989, new_n20990, new_n20991, new_n20992, new_n20993, new_n20994,
    new_n20995, new_n20996, new_n20997, new_n20998, new_n20999, new_n21000,
    new_n21001, new_n21002, new_n21003, new_n21004, new_n21005, new_n21006,
    new_n21007, new_n21008_1, new_n21009, new_n21010, new_n21011,
    new_n21012, new_n21013, new_n21014, new_n21015, new_n21016,
    new_n21017_1, new_n21018, new_n21019, new_n21020, new_n21021,
    new_n21022, new_n21023, new_n21024, new_n21025, new_n21026, new_n21027,
    new_n21028, new_n21029, new_n21030, new_n21031, new_n21032, new_n21033,
    new_n21034_1, new_n21035, new_n21036, new_n21037, new_n21038,
    new_n21039, new_n21040, new_n21041, new_n21042, new_n21043, new_n21044,
    new_n21045, new_n21046_1, new_n21047, new_n21048, new_n21049,
    new_n21050, new_n21052, new_n21053, new_n21054, new_n21055, new_n21056,
    new_n21057, new_n21058, new_n21060, new_n21061, new_n21062_1,
    new_n21063, new_n21064, new_n21065, new_n21066, new_n21067, new_n21068,
    new_n21069, new_n21070, new_n21071, new_n21072, new_n21073, new_n21074,
    new_n21075, new_n21076, new_n21077, new_n21078_1, new_n21079,
    new_n21080, new_n21081, new_n21082, new_n21083, new_n21084, new_n21085,
    new_n21086, new_n21087, new_n21088, new_n21089, new_n21090, new_n21091,
    new_n21092, new_n21093_1, new_n21094_1, new_n21095_1, new_n21096,
    new_n21097, new_n21098, new_n21099, new_n21100, new_n21101, new_n21102,
    new_n21103, new_n21104, new_n21105, new_n21106, new_n21107, new_n21108,
    new_n21109, new_n21110, new_n21111, new_n21112, new_n21113, new_n21114,
    new_n21115, new_n21116, new_n21117, new_n21118, new_n21119, new_n21120,
    new_n21121, new_n21122, new_n21123_1, new_n21124, new_n21125,
    new_n21126, new_n21127, new_n21128, new_n21129, new_n21130, new_n21131,
    new_n21132, new_n21133, new_n21134_1, new_n21135, new_n21136,
    new_n21137, new_n21138_1, new_n21139, new_n21140, new_n21141,
    new_n21142, new_n21143, new_n21144, new_n21145, new_n21146, new_n21147,
    new_n21148, new_n21149, new_n21150, new_n21151, new_n21152, new_n21153,
    new_n21154_1, new_n21155, new_n21156, new_n21157_1, new_n21158,
    new_n21159, new_n21160, new_n21161, new_n21162, new_n21163, new_n21164,
    new_n21165, new_n21166, new_n21167, new_n21168_1, new_n21169,
    new_n21170, new_n21171, new_n21172, new_n21173_1, new_n21174,
    new_n21175, new_n21176_1, new_n21177, new_n21178, new_n21179,
    new_n21180, new_n21181, new_n21182_1, new_n21183, new_n21184,
    new_n21185, new_n21186, new_n21187, new_n21188, new_n21189, new_n21190,
    new_n21191, new_n21192, new_n21193_1, new_n21194, new_n21195,
    new_n21196, new_n21197, new_n21198, new_n21199, new_n21200, new_n21201,
    new_n21202, new_n21203_1, new_n21204, new_n21205, new_n21206,
    new_n21207, new_n21208, new_n21209, new_n21210, new_n21211, new_n21212,
    new_n21213, new_n21214, new_n21215, new_n21216, new_n21217, new_n21218,
    new_n21219, new_n21220, new_n21221, new_n21222_1, new_n21223,
    new_n21224, new_n21225_1, new_n21226_1, new_n21227, new_n21228,
    new_n21229, new_n21230, new_n21231, new_n21232, new_n21233, new_n21234,
    new_n21235, new_n21236, new_n21237, new_n21238_1, new_n21239,
    new_n21240, new_n21241, new_n21242, new_n21243, new_n21244, new_n21245,
    new_n21246, new_n21247, new_n21248, new_n21249, new_n21250, new_n21251,
    new_n21252, new_n21253, new_n21254_1, new_n21255, new_n21256,
    new_n21257, new_n21258, new_n21259, new_n21260, new_n21261, new_n21262,
    new_n21263, new_n21264, new_n21265, new_n21266, new_n21267, new_n21268,
    new_n21269, new_n21270, new_n21271, new_n21272, new_n21273, new_n21274,
    new_n21275, new_n21276_1, new_n21277, new_n21278, new_n21281,
    new_n21282, new_n21283, new_n21284, new_n21285, new_n21286,
    new_n21287_1, new_n21288, new_n21289, new_n21290, new_n21291,
    new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297,
    new_n21298_1, new_n21299, new_n21300, new_n21301, new_n21302_1,
    new_n21303, new_n21304, new_n21306, new_n21307, new_n21308, new_n21309,
    new_n21310, new_n21311, new_n21312, new_n21313, new_n21314, new_n21315,
    new_n21316, new_n21317_1, new_n21318, new_n21319, new_n21320,
    new_n21321, new_n21322, new_n21323, new_n21324, new_n21326, new_n21328,
    new_n21329, new_n21330, new_n21331, new_n21332, new_n21333, new_n21335,
    new_n21337, new_n21339, new_n21341, new_n21342, new_n21343, new_n21344,
    new_n21345, new_n21346, new_n21347, new_n21348, new_n21349_1,
    new_n21350, new_n21351, new_n21352, new_n21353, new_n21354, new_n21355,
    new_n21356, new_n21357, new_n21358, new_n21359, new_n21360, new_n21361,
    new_n21362, new_n21363, new_n21364, new_n21365_1, new_n21366,
    new_n21367_1, new_n21368, new_n21369, new_n21370, new_n21371,
    new_n21372, new_n21373, new_n21374, new_n21375, new_n21376, new_n21377,
    new_n21378, new_n21379, new_n21380, new_n21381, new_n21382, new_n21383,
    new_n21384, new_n21385, new_n21386, new_n21387, new_n21388, new_n21389,
    new_n21390, new_n21391, new_n21392, new_n21393, new_n21394, new_n21395,
    new_n21396_1, new_n21397, new_n21398_1, new_n21399_1, new_n21400,
    new_n21401, new_n21402, new_n21403, new_n21404_1, new_n21405,
    new_n21406, new_n21407, new_n21408, new_n21409, new_n21410, new_n21411,
    new_n21412, new_n21413, new_n21414, new_n21415, new_n21416, new_n21417,
    new_n21418, new_n21419, new_n21420, new_n21421, new_n21422, new_n21423,
    new_n21424, new_n21425, new_n21426, new_n21427, new_n21428, new_n21429,
    new_n21430, new_n21431, new_n21432, new_n21433, new_n21434, new_n21435,
    new_n21436, new_n21437, new_n21438, new_n21439, new_n21440, new_n21441,
    new_n21442, new_n21443, new_n21444, new_n21445, new_n21446_1,
    new_n21447, new_n21448, new_n21449, new_n21450, new_n21451, new_n21452,
    new_n21453, new_n21454, new_n21455, new_n21456, new_n21457, new_n21458,
    new_n21460, new_n21462, new_n21464, new_n21465, new_n21466, new_n21467,
    new_n21468, new_n21469, new_n21470, new_n21471_1, new_n21472_1,
    new_n21473, new_n21474, new_n21475, new_n21476, new_n21477, new_n21478,
    new_n21479, new_n21480, new_n21481, new_n21483, new_n21484, new_n21485,
    new_n21486, new_n21487, new_n21488, new_n21489_1, new_n21490,
    new_n21491, new_n21492, new_n21493, new_n21494, new_n21495, new_n21496,
    new_n21497, new_n21498, new_n21499, new_n21500, new_n21501, new_n21502,
    new_n21503, new_n21504, new_n21505, new_n21506, new_n21507, new_n21508,
    new_n21509, new_n21510, new_n21511, new_n21512, new_n21513, new_n21514,
    new_n21515, new_n21516, new_n21517, new_n21518, new_n21519, new_n21520,
    new_n21521, new_n21522, new_n21523, new_n21524, new_n21525_1,
    new_n21526, new_n21527, new_n21528, new_n21529, new_n21530, new_n21531,
    new_n21532, new_n21533, new_n21534, new_n21535, new_n21536, new_n21537,
    new_n21538_1, new_n21539, new_n21540, new_n21542, new_n21544,
    new_n21545, new_n21546, new_n21547, new_n21548, new_n21549_1,
    new_n21550, new_n21551, new_n21552, new_n21553, new_n21554, new_n21555,
    new_n21556, new_n21557, new_n21558, new_n21559, new_n21560, new_n21561,
    new_n21562, new_n21563, new_n21564, new_n21565, new_n21566, new_n21567,
    new_n21568, new_n21569, new_n21570, new_n21571, new_n21572, new_n21573,
    new_n21574, new_n21575, new_n21576, new_n21577, new_n21578, new_n21579,
    new_n21581, new_n21582, new_n21583, new_n21584, new_n21585, new_n21586,
    new_n21587, new_n21588, new_n21589, new_n21590, new_n21591, new_n21592,
    new_n21593, new_n21594, new_n21595, new_n21596, new_n21597, new_n21598,
    new_n21599_1, new_n21600, new_n21601, new_n21602, new_n21603,
    new_n21604, new_n21605, new_n21606, new_n21607, new_n21608, new_n21609,
    new_n21610, new_n21611, new_n21612, new_n21613, new_n21614,
    new_n21615_1, new_n21616, new_n21617, new_n21618, new_n21619,
    new_n21620, new_n21621, new_n21622, new_n21624, new_n21625, new_n21627,
    new_n21629, new_n21631, new_n21632, new_n21633, new_n21634, new_n21635,
    new_n21636, new_n21637_1, new_n21638, new_n21639, new_n21640,
    new_n21641, new_n21642, new_n21643, new_n21644, new_n21645_1,
    new_n21646, new_n21647, new_n21648, new_n21649_1, new_n21650,
    new_n21651, new_n21652, new_n21653, new_n21654_1, new_n21655,
    new_n21657, new_n21659, new_n21661, new_n21663, new_n21664,
    new_n21665_1, new_n21666, new_n21667, new_n21668, new_n21669,
    new_n21670, new_n21671, new_n21672, new_n21673, new_n21674_1,
    new_n21675, new_n21676, new_n21677, new_n21678, new_n21679,
    new_n21680_1, new_n21681, new_n21682, new_n21683, new_n21684,
    new_n21685_1, new_n21686, new_n21687_1, new_n21688, new_n21689,
    new_n21690, new_n21691, new_n21692, new_n21693, new_n21694, new_n21695,
    new_n21696, new_n21697, new_n21698, new_n21699, new_n21700, new_n21701,
    new_n21702, new_n21703, new_n21704, new_n21705, new_n21706, new_n21707,
    new_n21708, new_n21709, new_n21710, new_n21711, new_n21712, new_n21713,
    new_n21714, new_n21715, new_n21716, new_n21717_1, new_n21718,
    new_n21719_1, new_n21720, new_n21721, new_n21722, new_n21723,
    new_n21724, new_n21725, new_n21726, new_n21727, new_n21728, new_n21729,
    new_n21730, new_n21731, new_n21732, new_n21733, new_n21734,
    new_n21735_1, new_n21736, new_n21737, new_n21738, new_n21739,
    new_n21740, new_n21741, new_n21742, new_n21743, new_n21744, new_n21745,
    new_n21746, new_n21747, new_n21748, new_n21749_1, new_n21750_1,
    new_n21751, new_n21752, new_n21753_1, new_n21754, new_n21755,
    new_n21756, new_n21757, new_n21758, new_n21760, new_n21762, new_n21764,
    new_n21766, new_n21768, new_n21769, new_n21770, new_n21771, new_n21772,
    new_n21773, new_n21774, new_n21775, new_n21776, new_n21777, new_n21778,
    new_n21779_1, new_n21780, new_n21781, new_n21782, new_n21783,
    new_n21784_1, new_n21785, new_n21786, new_n21787, new_n21788,
    new_n21789, new_n21791, new_n21792, new_n21793, new_n21794, new_n21795,
    new_n21796, new_n21797, new_n21798, new_n21799, new_n21800_1,
    new_n21801, new_n21802, new_n21803, new_n21804, new_n21805, new_n21806,
    new_n21807, new_n21808, new_n21809, new_n21810, new_n21811, new_n21812,
    new_n21813, new_n21814, new_n21815, new_n21816, new_n21817, new_n21818,
    new_n21819, new_n21820_1, new_n21821, new_n21822, new_n21823,
    new_n21824, new_n21825, new_n21826, new_n21827, new_n21828, new_n21829,
    new_n21830, new_n21831, new_n21832_1, new_n21833, new_n21834,
    new_n21835, new_n21836, new_n21837, new_n21838, new_n21839_1,
    new_n21840, new_n21841, new_n21842, new_n21843, new_n21844, new_n21845,
    new_n21846, new_n21847, new_n21848, new_n21849, new_n21850, new_n21851,
    new_n21852, new_n21853, new_n21854, new_n21855, new_n21856, new_n21857,
    new_n21858, new_n21859, new_n21860, new_n21861, new_n21862, new_n21863,
    new_n21864, new_n21865, new_n21866, new_n21867, new_n21868, new_n21869,
    new_n21870, new_n21871, new_n21872, new_n21873, new_n21876, new_n21878,
    new_n21880, new_n21881, new_n21882, new_n21883, new_n21884, new_n21885,
    new_n21886, new_n21887, new_n21888, new_n21889, new_n21890, new_n21891,
    new_n21892, new_n21893, new_n21894, new_n21895, new_n21896, new_n21897,
    new_n21898_1, new_n21899, new_n21900, new_n21901, new_n21902,
    new_n21903, new_n21904, new_n21905_1, new_n21906, new_n21907,
    new_n21908, new_n21909, new_n21910, new_n21911, new_n21912, new_n21913,
    new_n21914, new_n21915_1, new_n21916, new_n21917, new_n21918,
    new_n21919, new_n21920, new_n21921, new_n21922, new_n21923, new_n21924,
    new_n21925, new_n21926, new_n21927, new_n21928, new_n21929, new_n21930,
    new_n21931, new_n21932, new_n21933, new_n21934_1, new_n21935,
    new_n21936, new_n21937, new_n21938, new_n21939, new_n21940, new_n21941,
    new_n21942, new_n21943_1, new_n21944, new_n21945, new_n21946,
    new_n21948, new_n21950, new_n21951, new_n21952, new_n21953, new_n21954,
    new_n21955, new_n21956, new_n21957_1, new_n21958, new_n21959,
    new_n21960_1, new_n21961, new_n21962, new_n21963, new_n21964,
    new_n21965, new_n21966, new_n21967, new_n21968, new_n21969, new_n21970,
    new_n21971, new_n21972, new_n21973, new_n21974, new_n21975,
    new_n21976_1, new_n21977, new_n21978, new_n21979, new_n21980,
    new_n21981_1, new_n21982, new_n21983, new_n21984, new_n21985,
    new_n21986_1, new_n21987, new_n21988, new_n21989, new_n21990,
    new_n21991, new_n21992, new_n21993_1, new_n21994, new_n21995,
    new_n21996, new_n21997_1, new_n21998, new_n21999, new_n22000,
    new_n22001, new_n22002, new_n22003, new_n22004, new_n22005, new_n22006,
    new_n22007, new_n22008, new_n22009, new_n22010, new_n22011, new_n22012,
    new_n22013, new_n22014, new_n22015, new_n22016_1, new_n22017,
    new_n22018, new_n22020, new_n22022, new_n22023, new_n22024, new_n22025,
    new_n22026, new_n22027_1, new_n22028, new_n22029, new_n22030,
    new_n22031, new_n22032, new_n22033, new_n22034, new_n22035, new_n22036,
    new_n22037, new_n22038, new_n22039, new_n22040, new_n22042,
    new_n22043_1, new_n22044, new_n22045, new_n22046, new_n22047,
    new_n22048, new_n22049, new_n22050_1, new_n22051, new_n22052,
    new_n22053, new_n22054, new_n22055, new_n22056, new_n22057, new_n22058,
    new_n22059, new_n22060, new_n22062, new_n22063_1, new_n22064,
    new_n22065, new_n22066, new_n22067, new_n22068_1, new_n22069,
    new_n22070, new_n22071, new_n22072_1, new_n22073, new_n22074,
    new_n22075, new_n22076_1, new_n22077, new_n22078, new_n22079,
    new_n22080, new_n22081, new_n22082, new_n22083, new_n22084, new_n22085,
    new_n22086, new_n22087, new_n22088, new_n22089, new_n22090_1,
    new_n22091, new_n22092, new_n22093, new_n22094, new_n22095, new_n22096,
    new_n22097, new_n22098, new_n22099, new_n22100, new_n22101, new_n22102,
    new_n22103, new_n22104, new_n22105, new_n22106, new_n22107_1,
    new_n22108, new_n22109, new_n22110, new_n22111, new_n22112,
    new_n22113_1, new_n22114, new_n22115, new_n22117, new_n22119,
    new_n22121, new_n22122, new_n22123, new_n22124_1, new_n22125,
    new_n22126_1, new_n22127, new_n22128, new_n22129, new_n22130_1,
    new_n22131, new_n22132, new_n22133, new_n22134, new_n22135, new_n22136,
    new_n22137, new_n22138, new_n22139, new_n22140, new_n22141, new_n22142,
    new_n22143, new_n22144_1, new_n22145, new_n22146, new_n22147,
    new_n22148, new_n22149, new_n22150_1, new_n22151, new_n22152,
    new_n22153, new_n22154, new_n22155, new_n22156, new_n22157_1,
    new_n22158, new_n22159, new_n22160, new_n22161, new_n22162, new_n22163,
    new_n22164, new_n22165, new_n22166, new_n22167, new_n22168, new_n22169,
    new_n22170, new_n22171, new_n22172, new_n22173_1, new_n22174,
    new_n22175, new_n22176, new_n22178, new_n22179, new_n22180, new_n22181,
    new_n22182, new_n22183, new_n22184, new_n22185, new_n22186, new_n22187,
    new_n22188, new_n22189, new_n22190, new_n22191, new_n22192, new_n22193,
    new_n22194, new_n22195, new_n22196, new_n22197, new_n22198_1,
    new_n22199, new_n22200, new_n22201_1, new_n22202, new_n22203,
    new_n22204, new_n22205, new_n22206, new_n22207, new_n22208, new_n22210,
    new_n22211, new_n22212, new_n22213_1, new_n22214, new_n22215,
    new_n22216, new_n22217, new_n22218, new_n22219, new_n22220, new_n22221,
    new_n22222, new_n22223, new_n22224, new_n22225, new_n22226, new_n22227,
    new_n22228, new_n22229, new_n22230, new_n22232, new_n22234, new_n22236,
    new_n22238, new_n22239, new_n22240, new_n22241, new_n22242, new_n22243,
    new_n22244, new_n22245, new_n22246, new_n22247, new_n22248, new_n22249,
    new_n22250, new_n22252, new_n22254, new_n22255, new_n22256, new_n22257,
    new_n22258, new_n22259, new_n22260, new_n22261, new_n22262, new_n22263,
    new_n22264, new_n22265, new_n22266, new_n22267, new_n22268, new_n22269,
    new_n22270_1, new_n22271, new_n22272, new_n22273, new_n22274_1,
    new_n22275, new_n22276, new_n22277, new_n22278, new_n22279, new_n22280,
    new_n22281, new_n22282, new_n22283_1, new_n22284, new_n22285,
    new_n22286, new_n22287, new_n22288, new_n22289, new_n22290_1,
    new_n22291, new_n22292, new_n22293, new_n22294, new_n22295, new_n22296,
    new_n22297, new_n22298, new_n22299, new_n22300, new_n22301, new_n22302,
    new_n22303, new_n22304, new_n22305, new_n22306, new_n22307, new_n22308,
    new_n22309_1, new_n22310, new_n22311_1, new_n22312, new_n22313,
    new_n22314, new_n22315, new_n22316, new_n22317_1, new_n22318,
    new_n22319, new_n22320, new_n22321, new_n22322, new_n22323, new_n22325,
    new_n22327, new_n22329, new_n22331, new_n22332_1, new_n22333,
    new_n22334, new_n22335_1, new_n22336, new_n22337, new_n22338,
    new_n22339, new_n22340, new_n22341_1, new_n22342, new_n22343,
    new_n22344, new_n22345, new_n22346, new_n22347, new_n22348, new_n22349,
    new_n22350, new_n22351, new_n22353_1, new_n22355, new_n22357,
    new_n22358_1, new_n22359_1, new_n22360, new_n22361, new_n22362,
    new_n22363, new_n22364, new_n22365, new_n22366, new_n22367, new_n22368,
    new_n22369, new_n22370, new_n22371, new_n22372, new_n22373, new_n22374,
    new_n22375, new_n22376, new_n22377, new_n22378, new_n22379_1,
    new_n22380, new_n22381, new_n22382, new_n22383, new_n22384, new_n22385,
    new_n22386, new_n22387, new_n22388, new_n22389, new_n22390, new_n22391,
    new_n22392, new_n22393, new_n22394, new_n22395, new_n22396, new_n22397,
    new_n22398, new_n22399, new_n22400, new_n22401, new_n22402, new_n22403,
    new_n22404, new_n22405, new_n22406, new_n22407, new_n22408, new_n22409,
    new_n22410, new_n22411, new_n22412, new_n22413, new_n22414, new_n22415,
    new_n22416, new_n22417, new_n22418, new_n22419, new_n22420, new_n22421,
    new_n22422, new_n22423, new_n22424, new_n22425, new_n22426, new_n22427,
    new_n22428, new_n22429, new_n22430, new_n22431, new_n22432,
    new_n22433_1, new_n22434, new_n22435, new_n22436, new_n22437,
    new_n22438, new_n22439, new_n22440, new_n22441, new_n22442_1,
    new_n22443, new_n22444_1, new_n22445, new_n22446, new_n22447,
    new_n22448, new_n22449, new_n22450, new_n22451, new_n22452, new_n22453,
    new_n22454, new_n22455, new_n22456, new_n22457, new_n22458, new_n22459,
    new_n22460, new_n22461, new_n22462, new_n22463, new_n22464, new_n22465,
    new_n22467_1, new_n22469, new_n22471, new_n22473, new_n22475,
    new_n22477, new_n22479, new_n22480, new_n22481, new_n22482, new_n22483,
    new_n22484_1, new_n22485, new_n22486, new_n22487, new_n22488,
    new_n22489_1, new_n22490, new_n22491, new_n22492_1, new_n22493,
    new_n22494_1, new_n22495, new_n22496, new_n22497, new_n22498,
    new_n22499, new_n22500, new_n22501, new_n22502, new_n22503, new_n22504,
    new_n22505, new_n22506, new_n22507, new_n22508, new_n22509, new_n22510,
    new_n22511, new_n22512, new_n22513, new_n22514, new_n22515, new_n22516,
    new_n22517, new_n22518, new_n22519, new_n22520, new_n22521, new_n22522,
    new_n22523, new_n22525, new_n22527, new_n22529, new_n22530, new_n22531,
    new_n22532, new_n22533_1, new_n22534, new_n22535, new_n22536,
    new_n22537, new_n22538, new_n22539, new_n22540, new_n22541, new_n22542,
    new_n22543, new_n22544, new_n22545, new_n22546, new_n22547, new_n22548,
    new_n22549, new_n22550, new_n22551, new_n22552, new_n22553,
    new_n22554_1, new_n22555, new_n22556, new_n22557, new_n22558,
    new_n22559, new_n22560, new_n22561, new_n22562, new_n22563, new_n22564,
    new_n22565, new_n22566, new_n22567, new_n22568, new_n22569, new_n22570,
    new_n22571, new_n22572, new_n22573, new_n22574, new_n22575, new_n22576,
    new_n22577, new_n22578, new_n22579, new_n22580, new_n22581, new_n22582,
    new_n22583, new_n22584_1, new_n22585, new_n22586, new_n22587,
    new_n22588_1, new_n22589_1, new_n22590, new_n22591_1, new_n22592,
    new_n22593, new_n22594, new_n22595, new_n22596, new_n22597_1,
    new_n22598, new_n22599, new_n22600, new_n22601, new_n22602, new_n22603,
    new_n22604, new_n22605, new_n22606, new_n22607, new_n22608, new_n22609,
    new_n22610, new_n22611, new_n22612, new_n22613, new_n22614, new_n22615,
    new_n22616, new_n22617, new_n22618, new_n22619_1, new_n22620_1,
    new_n22621, new_n22622, new_n22623_1, new_n22624, new_n22625,
    new_n22626_1, new_n22627, new_n22628, new_n22629, new_n22630,
    new_n22631_1, new_n22633, new_n22634, new_n22635, new_n22636,
    new_n22637, new_n22638, new_n22639, new_n22640, new_n22642, new_n22644,
    new_n22646, new_n22647, new_n22648, new_n22649, new_n22650, new_n22651,
    new_n22652, new_n22653, new_n22654, new_n22655, new_n22656, new_n22657,
    new_n22658, new_n22659, new_n22660_1, new_n22661, new_n22662,
    new_n22663, new_n22664, new_n22665, new_n22666, new_n22667, new_n22668,
    new_n22669, new_n22670, new_n22671, new_n22672, new_n22673, new_n22674,
    new_n22676, new_n22677, new_n22678, new_n22679, new_n22680, new_n22681,
    new_n22682, new_n22683, new_n22684, new_n22685, new_n22686, new_n22687,
    new_n22688, new_n22689, new_n22690, new_n22691, new_n22692, new_n22693,
    new_n22694, new_n22695, new_n22696, new_n22697_1, new_n22698,
    new_n22699, new_n22700, new_n22701, new_n22702, new_n22703, new_n22704,
    new_n22705, new_n22706, new_n22707, new_n22708, new_n22709, new_n22710,
    new_n22711, new_n22712, new_n22713, new_n22714_1, new_n22715,
    new_n22716, new_n22717, new_n22718, new_n22719, new_n22720, new_n22721,
    new_n22722, new_n22723, new_n22724, new_n22725, new_n22726, new_n22727,
    new_n22728, new_n22729, new_n22730, new_n22731, new_n22732, new_n22733,
    new_n22734, new_n22735, new_n22736, new_n22737, new_n22738, new_n22739,
    new_n22740, new_n22741, new_n22742, new_n22743, new_n22744, new_n22745,
    new_n22746, new_n22747, new_n22748, new_n22749, new_n22750, new_n22751,
    new_n22753, new_n22755, new_n22757, new_n22758, new_n22759, new_n22760,
    new_n22761_1, new_n22762, new_n22763, new_n22764_1, new_n22765,
    new_n22766, new_n22767, new_n22768, new_n22769, new_n22770, new_n22771,
    new_n22772, new_n22773, new_n22774, new_n22775, new_n22776, new_n22777,
    new_n22778, new_n22779_1, new_n22780, new_n22781, new_n22782,
    new_n22783, new_n22784, new_n22785, new_n22786, new_n22787_1,
    new_n22788, new_n22789, new_n22790, new_n22791, new_n22792,
    new_n22793_1, new_n22794, new_n22795, new_n22796, new_n22797,
    new_n22798, new_n22799, new_n22800, new_n22801, new_n22802, new_n22803,
    new_n22804, new_n22805, new_n22806, new_n22807, new_n22808, new_n22809,
    new_n22810, new_n22811, new_n22812, new_n22813, new_n22814, new_n22815,
    new_n22816, new_n22817, new_n22818, new_n22819_1, new_n22820,
    new_n22821, new_n22822, new_n22823, new_n22824, new_n22825, new_n22826,
    new_n22827, new_n22828, new_n22829, new_n22830, new_n22831, new_n22832,
    new_n22833, new_n22834, new_n22835, new_n22836, new_n22837, new_n22838,
    new_n22839, new_n22840, new_n22841, new_n22842, new_n22843_1,
    new_n22844, new_n22845, new_n22846, new_n22847, new_n22848, new_n22849,
    new_n22850, new_n22851, new_n22852, new_n22853, new_n22854, new_n22855,
    new_n22856, new_n22857, new_n22858_1, new_n22859, new_n22860,
    new_n22861, new_n22862, new_n22863, new_n22864, new_n22865, new_n22866,
    new_n22867, new_n22868, new_n22869, new_n22870_1, new_n22871_1,
    new_n22872, new_n22874, new_n22876, new_n22877, new_n22878,
    new_n22879_1, new_n22880, new_n22881, new_n22882, new_n22883,
    new_n22884, new_n22885, new_n22886, new_n22887, new_n22888, new_n22889,
    new_n22890, new_n22891_1, new_n22892, new_n22893, new_n22894,
    new_n22895, new_n22896, new_n22897_1, new_n22898, new_n22899,
    new_n22900, new_n22901, new_n22902, new_n22903_1, new_n22904,
    new_n22905, new_n22906, new_n22907_1, new_n22908, new_n22909,
    new_n22910_1, new_n22911, new_n22912, new_n22913, new_n22914_1,
    new_n22915, new_n22916, new_n22917, new_n22918_1, new_n22919,
    new_n22920, new_n22921, new_n22922, new_n22923, new_n22924, new_n22925,
    new_n22926, new_n22927, new_n22928, new_n22929, new_n22930, new_n22931,
    new_n22932, new_n22933, new_n22934, new_n22935, new_n22936, new_n22937,
    new_n22938, new_n22939_1, new_n22940, new_n22941, new_n22942,
    new_n22943, new_n22944, new_n22945, new_n22946, new_n22947, new_n22948,
    new_n22949, new_n22950, new_n22951, new_n22952, new_n22954, new_n22956,
    new_n22958, new_n22960, new_n22962, new_n22964, new_n22965, new_n22967,
    new_n22970, new_n22971, new_n22972, new_n22973, new_n22974, new_n22975,
    new_n22976, new_n22977, new_n22978, new_n22979, new_n22980, new_n22981,
    new_n22982, new_n22983, new_n22984, new_n22985, new_n22986, new_n22987,
    new_n22988, new_n22989, new_n22990, new_n22991, new_n22992, new_n22993,
    new_n22994, new_n22995, new_n22996, new_n22997, new_n22998_1,
    new_n22999, new_n23000, new_n23001, new_n23002, new_n23003, new_n23004,
    new_n23005, new_n23006_1, new_n23007_1, new_n23008, new_n23009_1,
    new_n23010, new_n23011, new_n23012, new_n23013, new_n23014_1,
    new_n23015, new_n23016, new_n23017, new_n23018, new_n23019, new_n23020,
    new_n23021, new_n23022, new_n23023, new_n23024, new_n23025, new_n23026,
    new_n23027, new_n23028, new_n23029, new_n23030, new_n23031, new_n23032,
    new_n23033, new_n23034, new_n23035_1, new_n23036, new_n23037,
    new_n23038, new_n23039_1, new_n23040, new_n23041, new_n23042,
    new_n23043, new_n23044, new_n23045, new_n23046, new_n23047_1,
    new_n23048, new_n23049, new_n23050, new_n23051, new_n23052, new_n23053,
    new_n23054, new_n23055, new_n23056, new_n23057, new_n23058_1,
    new_n23059, new_n23060, new_n23061, new_n23062, new_n23063, new_n23064,
    new_n23065_1, new_n23066_1, new_n23067_1, new_n23068_1, new_n23069,
    new_n23070, new_n23071, new_n23072, new_n23073, new_n23074, new_n23075,
    new_n23076, new_n23077, new_n23078, new_n23079, new_n23080, new_n23081,
    new_n23082, new_n23083, new_n23084, new_n23085, new_n23086, new_n23087,
    new_n23088, new_n23089, new_n23090, new_n23091, new_n23092, new_n23093,
    new_n23094, new_n23095, new_n23096, new_n23097, new_n23098, new_n23099,
    new_n23100, new_n23101, new_n23102, new_n23103, new_n23104, new_n23105,
    new_n23106, new_n23107, new_n23108, new_n23109, new_n23110, new_n23111,
    new_n23112, new_n23113, new_n23114, new_n23115, new_n23116, new_n23117,
    new_n23118, new_n23119, new_n23120_1, new_n23121, new_n23122,
    new_n23123, new_n23124, new_n23127, new_n23128, new_n23129, new_n23130,
    new_n23131, new_n23132, new_n23133, new_n23134, new_n23135, new_n23136,
    new_n23137, new_n23138, new_n23139, new_n23140, new_n23141, new_n23142,
    new_n23143, new_n23144, new_n23145, new_n23146_1, new_n23147,
    new_n23148, new_n23149, new_n23150, new_n23151, new_n23152, new_n23153,
    new_n23154, new_n23155, new_n23156, new_n23157, new_n23158, new_n23159,
    new_n23160_1, new_n23161, new_n23162, new_n23163, new_n23164,
    new_n23165, new_n23166_1, new_n23167, new_n23168, new_n23169,
    new_n23170, new_n23171, new_n23172, new_n23173, new_n23174, new_n23175,
    new_n23176, new_n23177, new_n23178, new_n23179, new_n23180, new_n23181,
    new_n23182, new_n23183, new_n23184, new_n23185, new_n23186, new_n23187,
    new_n23188, new_n23189, new_n23190, new_n23191, new_n23192, new_n23193,
    new_n23194, new_n23195, new_n23196, new_n23197, new_n23198, new_n23199,
    new_n23200_1, new_n23201, new_n23202, new_n23203, new_n23204,
    new_n23205, new_n23206, new_n23207, new_n23208, new_n23209, new_n23210,
    new_n23211, new_n23212, new_n23213, new_n23214, new_n23215, new_n23216,
    new_n23217, new_n23218, new_n23219, new_n23220, new_n23221, new_n23222,
    new_n23223, new_n23224, new_n23225, new_n23226, new_n23227, new_n23228,
    new_n23229, new_n23231, new_n23233, new_n23235, new_n23237,
    new_n23238_1, new_n23239, new_n23240, new_n23241, new_n23242,
    new_n23243, new_n23244, new_n23245, new_n23246, new_n23247_1,
    new_n23248_1, new_n23249, new_n23250_1, new_n23251, new_n23252,
    new_n23253, new_n23254, new_n23255, new_n23256, new_n23257, new_n23258,
    new_n23259, new_n23260, new_n23261, new_n23262, new_n23263, new_n23264,
    new_n23265, new_n23266, new_n23267, new_n23268, new_n23269,
    new_n23270_1, new_n23271, new_n23272_1, new_n23273, new_n23274,
    new_n23275, new_n23276, new_n23277, new_n23278, new_n23279, new_n23280,
    new_n23281, new_n23282, new_n23283, new_n23284, new_n23285, new_n23286,
    new_n23287, new_n23288, new_n23289_1, new_n23290, new_n23291,
    new_n23292, new_n23293, new_n23294, new_n23295, new_n23296, new_n23297,
    new_n23298, new_n23299, new_n23300, new_n23301, new_n23302, new_n23303,
    new_n23304_1, new_n23305_1, new_n23306, new_n23307, new_n23308,
    new_n23309, new_n23310, new_n23311, new_n23312, new_n23313, new_n23314,
    new_n23315, new_n23316, new_n23317, new_n23318, new_n23319, new_n23320,
    new_n23321, new_n23322, new_n23323, new_n23324, new_n23325, new_n23326,
    new_n23327, new_n23328, new_n23329, new_n23330, new_n23331, new_n23332,
    new_n23333_1, new_n23334, new_n23335, new_n23336, new_n23337,
    new_n23338, new_n23339, new_n23340, new_n23341_1, new_n23342_1,
    new_n23343, new_n23345, new_n23346, new_n23347, new_n23348, new_n23349,
    new_n23350, new_n23351, new_n23352, new_n23353, new_n23355_1,
    new_n23356, new_n23357, new_n23358, new_n23359, new_n23360, new_n23361,
    new_n23362, new_n23363, new_n23364, new_n23365, new_n23366, new_n23367,
    new_n23368, new_n23369_1, new_n23370, new_n23371_1, new_n23372,
    new_n23373, new_n23374, new_n23375, new_n23376, new_n23377, new_n23378,
    new_n23380, new_n23382, new_n23384, new_n23386, new_n23388, new_n23390,
    new_n23391, new_n23392, new_n23393, new_n23394, new_n23395, new_n23396,
    new_n23397, new_n23398, new_n23399, new_n23400, new_n23401_1,
    new_n23402, new_n23403, new_n23404, new_n23405, new_n23406, new_n23408,
    new_n23411, new_n23413, new_n23415, new_n23417, new_n23419, new_n23421,
    new_n23423, new_n23426, new_n23427, new_n23428, new_n23429_1,
    new_n23430_1, new_n23431, new_n23432, new_n23433_1, new_n23434_1,
    new_n23435, new_n23436, new_n23437, new_n23438, new_n23439, new_n23440,
    new_n23441, new_n23442, new_n23443, new_n23444, new_n23445, new_n23446,
    new_n23447, new_n23448, new_n23449, new_n23450_1, new_n23451,
    new_n23452, new_n23453, new_n23454, new_n23455, new_n23456, new_n23457,
    new_n23458, new_n23459, new_n23460, new_n23461, new_n23462,
    new_n23463_1, new_n23464, new_n23466, new_n23468, new_n23469,
    new_n23470, new_n23471_1, new_n23472, new_n23473, new_n23474,
    new_n23475, new_n23476, new_n23477, new_n23478, new_n23479,
    new_n23480_1, new_n23481, new_n23482, new_n23483, new_n23484,
    new_n23485, new_n23486, new_n23487, new_n23488, new_n23489, new_n23490,
    new_n23491, new_n23492, new_n23493_1, new_n23494, new_n23495,
    new_n23496, new_n23497, new_n23498, new_n23499, new_n23501, new_n23502,
    new_n23503, new_n23504, new_n23505, new_n23506, new_n23507, new_n23508,
    new_n23509, new_n23510, new_n23511, new_n23512, new_n23513_1,
    new_n23514, new_n23515, new_n23516, new_n23517, new_n23518, new_n23519,
    new_n23520, new_n23521, new_n23522, new_n23523, new_n23524, new_n23525,
    new_n23526, new_n23527, new_n23528, new_n23529_1, new_n23530,
    new_n23531, new_n23532, new_n23533, new_n23534, new_n23535, new_n23536,
    new_n23537, new_n23538, new_n23539, new_n23540, new_n23541_1,
    new_n23542, new_n23543, new_n23544, new_n23545, new_n23546_1,
    new_n23547, new_n23548, new_n23549, new_n23550_1, new_n23551,
    new_n23552, new_n23553, new_n23554, new_n23555, new_n23556, new_n23557,
    new_n23558, new_n23559, new_n23560, new_n23561, new_n23562, new_n23563,
    new_n23564, new_n23565, new_n23566, new_n23567, new_n23568, new_n23569,
    new_n23570, new_n23571, new_n23572, new_n23573, new_n23574, new_n23575,
    new_n23576, new_n23577, new_n23578, new_n23579, new_n23580, new_n23581,
    new_n23582, new_n23583, new_n23584, new_n23585_1, new_n23586_1,
    new_n23587, new_n23588_1, new_n23589, new_n23590, new_n23591,
    new_n23592, new_n23593, new_n23594, new_n23595, new_n23596, new_n23597,
    new_n23598, new_n23599, new_n23600, new_n23601, new_n23602, new_n23603,
    new_n23604, new_n23605, new_n23606, new_n23607, new_n23608, new_n23609,
    new_n23610, new_n23611, new_n23612, new_n23613, new_n23614, new_n23615,
    new_n23616, new_n23617, new_n23618, new_n23619_1, new_n23620,
    new_n23621, new_n23622, new_n23623, new_n23624_1, new_n23625,
    new_n23626, new_n23627, new_n23628_1, new_n23629, new_n23630,
    new_n23631, new_n23632, new_n23633, new_n23634, new_n23635, new_n23636,
    new_n23637_1, new_n23638, new_n23639, new_n23640, new_n23641,
    new_n23642, new_n23643, new_n23644, new_n23645, new_n23646, new_n23647,
    new_n23648, new_n23649, new_n23650, new_n23651, new_n23652, new_n23653,
    new_n23654, new_n23655, new_n23656, new_n23657_1, new_n23658,
    new_n23659, new_n23660, new_n23661, new_n23662, new_n23663_1,
    new_n23664, new_n23665, new_n23666, new_n23667, new_n23668,
    new_n23669_1, new_n23670, new_n23671, new_n23672, new_n23673,
    new_n23674, new_n23675, new_n23676, new_n23677, new_n23678, new_n23679,
    new_n23680, new_n23681, new_n23682, new_n23684_1, new_n23686,
    new_n23688, new_n23690_1, new_n23691, new_n23692, new_n23693,
    new_n23694, new_n23695, new_n23696, new_n23697_1, new_n23698,
    new_n23699, new_n23700, new_n23701, new_n23702, new_n23703, new_n23704,
    new_n23705, new_n23706, new_n23707, new_n23708, new_n23709, new_n23710,
    new_n23711, new_n23712, new_n23713, new_n23714_1, new_n23715,
    new_n23716, new_n23718, new_n23720, new_n23721, new_n23722, new_n23723,
    new_n23724, new_n23725, new_n23726, new_n23727, new_n23728, new_n23729,
    new_n23730, new_n23731, new_n23732, new_n23733, new_n23734, new_n23735,
    new_n23736, new_n23737, new_n23738, new_n23740, new_n23742, new_n23743,
    new_n23744, new_n23745, new_n23746, new_n23747, new_n23748_1,
    new_n23749, new_n23751, new_n23753, new_n23755_1, new_n23757,
    new_n23759, new_n23761, new_n23763, new_n23764, new_n23765, new_n23766,
    new_n23767, new_n23768, new_n23769, new_n23770, new_n23771, new_n23772,
    new_n23773, new_n23774, new_n23775_1, new_n23776, new_n23777,
    new_n23778, new_n23779, new_n23780, new_n23781, new_n23783, new_n23785,
    new_n23787, new_n23788, new_n23789, new_n23790, new_n23791, new_n23792,
    new_n23793, new_n23794, new_n23795, new_n23796, new_n23797, new_n23798,
    new_n23800, new_n23801, new_n23802, new_n23803, new_n23804, new_n23805,
    new_n23806, new_n23807, new_n23808, new_n23809, new_n23810, new_n23811,
    new_n23812, new_n23813, new_n23814, new_n23815, new_n23816, new_n23817,
    new_n23818, new_n23819, new_n23820, new_n23821, new_n23822, new_n23823,
    new_n23825, new_n23826, new_n23827, new_n23828, new_n23829, new_n23830,
    new_n23831_1, new_n23832, new_n23833, new_n23834, new_n23835,
    new_n23836, new_n23837, new_n23838, new_n23839, new_n23840, new_n23841,
    new_n23842_1, new_n23843, new_n23844, new_n23845, new_n23846,
    new_n23847, new_n23848, new_n23849_1, new_n23850, new_n23851,
    new_n23852, new_n23853, new_n23854, new_n23855, new_n23856_1,
    new_n23857, new_n23858, new_n23859, new_n23860, new_n23862, new_n23863,
    new_n23864, new_n23865, new_n23866, new_n23867, new_n23868, new_n23869,
    new_n23870, new_n23871, new_n23872, new_n23873, new_n23874, new_n23875,
    new_n23876, new_n23877, new_n23878, new_n23879, new_n23880, new_n23881,
    new_n23882, new_n23883_1, new_n23884, new_n23885, new_n23886,
    new_n23887, new_n23888_1, new_n23889, new_n23890, new_n23891,
    new_n23892, new_n23893, new_n23894, new_n23895_1, new_n23896,
    new_n23897, new_n23898, new_n23899_1, new_n23900, new_n23901,
    new_n23902, new_n23903_1, new_n23904, new_n23905, new_n23906,
    new_n23907, new_n23908, new_n23909, new_n23910, new_n23911,
    new_n23912_1, new_n23913_1, new_n23914, new_n23915, new_n23916,
    new_n23917, new_n23918, new_n23919, new_n23920, new_n23921, new_n23922,
    new_n23923_1, new_n23924_1, new_n23925, new_n23926, new_n23927,
    new_n23928, new_n23929, new_n23930, new_n23931, new_n23932, new_n23933,
    new_n23934, new_n23935_1, new_n23936, new_n23937, new_n23938,
    new_n23939, new_n23940, new_n23941, new_n23942_1, new_n23943,
    new_n23944, new_n23945, new_n23946, new_n23947, new_n23948, new_n23949,
    new_n23950, new_n23951, new_n23952, new_n23953, new_n23954_1,
    new_n23955, new_n23956, new_n23957, new_n23958_1, new_n23960,
    new_n23962, new_n23964, new_n23966, new_n23967, new_n23968, new_n23969,
    new_n23970, new_n23971, new_n23972, new_n23973, new_n23974_1,
    new_n23975, new_n23976, new_n23977, new_n23978, new_n23979, new_n23980,
    new_n23981, new_n23982, new_n23983, new_n23984, new_n23985,
    new_n23986_1, new_n23987, new_n23988, new_n23989, new_n23990,
    new_n23991, new_n23992, new_n23993, new_n23994, new_n23995, new_n23996,
    new_n23997, new_n23998, new_n23999, new_n24000, new_n24001,
    new_n24002_1, new_n24003, new_n24004_1, new_n24005, new_n24006,
    new_n24007, new_n24008, new_n24009, new_n24010, new_n24011, new_n24012,
    new_n24013, new_n24014, new_n24015, new_n24016, new_n24017, new_n24018,
    new_n24019, new_n24020, new_n24021, new_n24022, new_n24023, new_n24024,
    new_n24025, new_n24026, new_n24027, new_n24028, new_n24029, new_n24030,
    new_n24031, new_n24032_1, new_n24033, new_n24034, new_n24035,
    new_n24036, new_n24037, new_n24038, new_n24039_1, new_n24040,
    new_n24041, new_n24042, new_n24043, new_n24044, new_n24045, new_n24046,
    new_n24047, new_n24048_1, new_n24049, new_n24050, new_n24051,
    new_n24052_1, new_n24053, new_n24054, new_n24055, new_n24056,
    new_n24057, new_n24058, new_n24059, new_n24060, new_n24061, new_n24062,
    new_n24063, new_n24064, new_n24065, new_n24066, new_n24067, new_n24068,
    new_n24069, new_n24070, new_n24071, new_n24072, new_n24073, new_n24074,
    new_n24075, new_n24076, new_n24077, new_n24078, new_n24079, new_n24080,
    new_n24081, new_n24082, new_n24083, new_n24084, new_n24085_1,
    new_n24086, new_n24087, new_n24088, new_n24089, new_n24090, new_n24091,
    new_n24092_1, new_n24093_1, new_n24094, new_n24095, new_n24096_1,
    new_n24097_1, new_n24098, new_n24099, new_n24100, new_n24101,
    new_n24102, new_n24103, new_n24104, new_n24106, new_n24108, new_n24110,
    new_n24112, new_n24114, new_n24116, new_n24118, new_n24119_1,
    new_n24120, new_n24121, new_n24122, new_n24123, new_n24124, new_n24125,
    new_n24126, new_n24127, new_n24128, new_n24129_1, new_n24130,
    new_n24131, new_n24132, new_n24133_1, new_n24134, new_n24135,
    new_n24136, new_n24137, new_n24138, new_n24139, new_n24140,
    new_n24141_1, new_n24142, new_n24143, new_n24144, new_n24145_1,
    new_n24146_1, new_n24147, new_n24148, new_n24149, new_n24150_1,
    new_n24151, new_n24152, new_n24153, new_n24154, new_n24155_1,
    new_n24157, new_n24158, new_n24159, new_n24160_1, new_n24161,
    new_n24162, new_n24163, new_n24164, new_n24165, new_n24166,
    new_n24167_1, new_n24168, new_n24169, new_n24170_1, new_n24171,
    new_n24172_1, new_n24173, new_n24174, new_n24175, new_n24176,
    new_n24177_1, new_n24178, new_n24179, new_n24180, new_n24181,
    new_n24182, new_n24183, new_n24184, new_n24185, new_n24186, new_n24187,
    new_n24188, new_n24189, new_n24190, new_n24191, new_n24192, new_n24194,
    new_n24196_1, new_n24198, new_n24200, new_n24202, new_n24204,
    new_n24206, new_n24208, new_n24209, new_n24210, new_n24211, new_n24212,
    new_n24213, new_n24214, new_n24215, new_n24216, new_n24217, new_n24218,
    new_n24219, new_n24220, new_n24222, new_n24224, new_n24226, new_n24227,
    new_n24228_1, new_n24229, new_n24230, new_n24231, new_n24232,
    new_n24233, new_n24234, new_n24235, new_n24236, new_n24237, new_n24238,
    new_n24239, new_n24240, new_n24241, new_n24242, new_n24243, new_n24244,
    new_n24245, new_n24246, new_n24247, new_n24248, new_n24249, new_n24250,
    new_n24251, new_n24252, new_n24253, new_n24254, new_n24255, new_n24256,
    new_n24257, new_n24258_1, new_n24259, new_n24260_1, new_n24262,
    new_n24264, new_n24265, new_n24266, new_n24267, new_n24268, new_n24269,
    new_n24270, new_n24271, new_n24272, new_n24273, new_n24274, new_n24275,
    new_n24276, new_n24277, new_n24278_1, new_n24279, new_n24280,
    new_n24281, new_n24282, new_n24283, new_n24284, new_n24285, new_n24286,
    new_n24287, new_n24288, new_n24289_1, new_n24290, new_n24291,
    new_n24292, new_n24293, new_n24294, new_n24295, new_n24296,
    new_n24297_1, new_n24298, new_n24299, new_n24300, new_n24301,
    new_n24302, new_n24303, new_n24304, new_n24305, new_n24306,
    new_n24307_1, new_n24308, new_n24309, new_n24310, new_n24311,
    new_n24312, new_n24313, new_n24314, new_n24315, new_n24316, new_n24317,
    new_n24318, new_n24319_1, new_n24320, new_n24321, new_n24322,
    new_n24323_1, new_n24324, new_n24325, new_n24326, new_n24327_1,
    new_n24328, new_n24329, new_n24330, new_n24331, new_n24332, new_n24334,
    new_n24335, new_n24336, new_n24337, new_n24338, new_n24339, new_n24340,
    new_n24341, new_n24342_1, new_n24343, new_n24344, new_n24345_1,
    new_n24346, new_n24347_1, new_n24348, new_n24349, new_n24350,
    new_n24351, new_n24352, new_n24353, new_n24354, new_n24355, new_n24356,
    new_n24357, new_n24358, new_n24359, new_n24360, new_n24361, new_n24362,
    new_n24363, new_n24364, new_n24365, new_n24367, new_n24369, new_n24370,
    new_n24371, new_n24372, new_n24373_1, new_n24374_1, new_n24375,
    new_n24376, new_n24377, new_n24378, new_n24379, new_n24380, new_n24381,
    new_n24382, new_n24383, new_n24384, new_n24385, new_n24386, new_n24387,
    new_n24388, new_n24389, new_n24390, new_n24391, new_n24392, new_n24393,
    new_n24394, new_n24395, new_n24396, new_n24397, new_n24398, new_n24399,
    new_n24400, new_n24401, new_n24402, new_n24403, new_n24404, new_n24405,
    new_n24406_1, new_n24408, new_n24410, new_n24412, new_n24414,
    new_n24415_1, new_n24416, new_n24417, new_n24418, new_n24419,
    new_n24420, new_n24421_1, new_n24422, new_n24423, new_n24424,
    new_n24425, new_n24426, new_n24427, new_n24428, new_n24429, new_n24430,
    new_n24431_1, new_n24432, new_n24433, new_n24434, new_n24435,
    new_n24436, new_n24437, new_n24438, new_n24439, new_n24440, new_n24441,
    new_n24442, new_n24443, new_n24444, new_n24445, new_n24446, new_n24447,
    new_n24448, new_n24449, new_n24450, new_n24451, new_n24452, new_n24453,
    new_n24454, new_n24455, new_n24456, new_n24457, new_n24459, new_n24461,
    new_n24462, new_n24463, new_n24464, new_n24465, new_n24466, new_n24467,
    new_n24468, new_n24469, new_n24470, new_n24471, new_n24472_1,
    new_n24473, new_n24474, new_n24475, new_n24476_1, new_n24477,
    new_n24478, new_n24479, new_n24480, new_n24481, new_n24482,
    new_n24483_1, new_n24484, new_n24485_1, new_n24486, new_n24487,
    new_n24488, new_n24489, new_n24491, new_n24493, new_n24496, new_n24498,
    new_n24500, new_n24502, new_n24503, new_n24504, new_n24505, new_n24506,
    new_n24507, new_n24508, new_n24509, new_n24510, new_n24511,
    new_n24512_1, new_n24513, new_n24514, new_n24515, new_n24516,
    new_n24517, new_n24518, new_n24519, new_n24520, new_n24521, new_n24522,
    new_n24523, new_n24524, new_n24525, new_n24526, new_n24527, new_n24528,
    new_n24529, new_n24530, new_n24531, new_n24532, new_n24533, new_n24534,
    new_n24535, new_n24536, new_n24537, new_n24538, new_n24539, new_n24540,
    new_n24541, new_n24542, new_n24543, new_n24544, new_n24545, new_n24546,
    new_n24547, new_n24548, new_n24549, new_n24550, new_n24551, new_n24552,
    new_n24553, new_n24554, new_n24555, new_n24556, new_n24557,
    new_n24558_1, new_n24559, new_n24560, new_n24561, new_n24563,
    new_n24565, new_n24567, new_n24569, new_n24571, new_n24575, new_n24577,
    new_n24578, new_n24579_1, new_n24580, new_n24581, new_n24582,
    new_n24583, new_n24584, new_n24585, new_n24588, new_n24590, new_n24592,
    new_n24595, new_n24597, new_n24599, new_n24601, new_n24603, new_n24606,
    new_n24608, new_n24609, new_n24611, new_n24613, new_n24615, new_n24616,
    new_n24617, new_n24618_1, new_n24619, new_n24620_1, new_n24621,
    new_n24622, new_n24623, new_n24624, new_n24625, new_n24626_1,
    new_n24627, new_n24628, new_n24629_1, new_n24630, new_n24631,
    new_n24632, new_n24633, new_n24634, new_n24635, new_n24636_1,
    new_n24637, new_n24638_1, new_n24639, new_n24640, new_n24641,
    new_n24643, new_n24644, new_n24645, new_n24646, new_n24647, new_n24648,
    new_n24649, new_n24650, new_n24651, new_n24652, new_n24653, new_n24654,
    new_n24655, new_n24656, new_n24657, new_n24658, new_n24659, new_n24660,
    new_n24662, new_n24663, new_n24664, new_n24665, new_n24666, new_n24667,
    new_n24668, new_n24669, new_n24670, new_n24671, new_n24672, new_n24673,
    new_n24674, new_n24676, new_n24678, new_n24680, new_n24682, new_n24683,
    new_n24684, new_n24685, new_n24686, new_n24687, new_n24688, new_n24689,
    new_n24690, new_n24691, new_n24692, new_n24693, new_n24694, new_n24695,
    new_n24696, new_n24697, new_n24698, new_n24699, new_n24700, new_n24701,
    new_n24702, new_n24703, new_n24704, new_n24705, new_n24706, new_n24707,
    new_n24708, new_n24709, new_n24711, new_n24714, new_n24716, new_n24718,
    new_n24720, new_n24722, new_n24724, new_n24725, new_n24726, new_n24727,
    new_n24728, new_n24730, new_n24732_1, new_n24734, new_n24736,
    new_n24738, new_n24739, new_n24740, new_n24741, new_n24742, new_n24743,
    new_n24745, new_n24748, new_n24750, new_n24752, new_n24754, new_n24756,
    new_n24758_1, new_n24760, new_n24761, new_n24762, new_n24763,
    new_n24764, new_n24765, new_n24766, new_n24767, new_n24768_1,
    new_n24769, new_n24770, new_n24771, new_n24772, new_n24773, new_n24774,
    new_n24775, new_n24776, new_n24777, new_n24778, new_n24780, new_n24782,
    new_n24784_1, new_n24786_1, new_n24787, new_n24788, new_n24789,
    new_n24790, new_n24794, new_n24796, new_n24798, new_n24800, new_n24801,
    new_n24802, new_n24803, new_n24804, new_n24805, new_n24806,
    new_n24807_1, new_n24808, new_n24809, new_n24810, new_n24811,
    new_n24812, new_n24813, new_n24814, new_n24815, new_n24816, new_n24817,
    new_n24818, new_n24819, new_n24820, new_n24821, new_n24822, new_n24823,
    new_n24824, new_n24825, new_n24826_1, new_n24827, new_n24828,
    new_n24829, new_n24830, new_n24831, new_n24832, new_n24833, new_n24834,
    new_n24835, new_n24836, new_n24837, new_n24838, new_n24839,
    new_n24840_1, new_n24841_1, new_n24842, new_n24843, new_n24844,
    new_n24845, new_n24846, new_n24847, new_n24848, new_n24849, new_n24850,
    new_n24851, new_n24852, new_n24853_1, new_n24855, new_n24857_1,
    new_n24858, new_n24859, new_n24860, new_n24861, new_n24862, new_n24863,
    new_n24864, new_n24865, new_n24866, new_n24867, new_n24868, new_n24870,
    new_n24871, new_n24872, new_n24873, new_n24874, new_n24875, new_n24876,
    new_n24877, new_n24878, new_n24879_1, new_n24880, new_n24881,
    new_n24882, new_n24883, new_n24884, new_n24885, new_n24886,
    new_n24887_1, new_n24888, new_n24889, new_n24891, new_n24893,
    new_n24895, new_n24899, new_n24901, new_n24903, new_n24905, new_n24906,
    new_n24907, new_n24908, new_n24909, new_n24910, new_n24911, new_n24912,
    new_n24913, new_n24914, new_n24915, new_n24916, new_n24917, new_n24918,
    new_n24919, new_n24920, new_n24921, new_n24922, new_n24923, new_n24924,
    new_n24925, new_n24926, new_n24927, new_n24928, new_n24929, new_n24930,
    new_n24931, new_n24932, new_n24933, new_n24935, new_n24937_1,
    new_n24939, new_n24941, new_n24943, new_n24944, new_n24945, new_n24947,
    new_n24948, new_n24950, new_n24952, new_n24954, new_n24957, new_n24959,
    new_n24961, new_n24963, new_n24964, new_n24965, new_n24966, new_n24967,
    new_n24968, new_n24969, new_n24970, new_n24971, new_n24972, new_n24973,
    new_n24974, new_n24975, new_n24976, new_n24977, new_n24978, new_n24979,
    new_n24980, new_n24981, new_n24982, new_n24983, new_n24984, new_n24985,
    new_n24986, new_n24987, new_n24988, new_n24989, new_n24990, new_n24991,
    new_n24992, new_n24993, new_n24994, new_n24995, new_n24996, new_n24997,
    new_n24998_1, new_n24999, new_n25000, new_n25001, new_n25002,
    new_n25003, new_n25004, new_n25005, new_n25006_1, new_n25007,
    new_n25008, new_n25009, new_n25010, new_n25011, new_n25012, new_n25013,
    new_n25014, new_n25015, new_n25016, new_n25017, new_n25018, new_n25019,
    new_n25020, new_n25021, new_n25022, new_n25023_1, new_n25024,
    new_n25025, new_n25026, new_n25027, new_n25028, new_n25029, new_n25030,
    new_n25031, new_n25032_1, new_n25033, new_n25034, new_n25035,
    new_n25036, new_n25038, new_n25039, new_n25040, new_n25041, new_n25042,
    new_n25043, new_n25044, new_n25045, new_n25046, new_n25047, new_n25048,
    new_n25049, new_n25050, new_n25051, new_n25052, new_n25053, new_n25054,
    new_n25055, new_n25056, new_n25057, new_n25058, new_n25059, new_n25060,
    new_n25061, new_n25062_1, new_n25063, new_n25064, new_n25065,
    new_n25066, new_n25067, new_n25068_1, new_n25069, new_n25070,
    new_n25071, new_n25072, new_n25073_1, new_n25074_1, new_n25075,
    new_n25076, new_n25077, new_n25078, new_n25079, new_n25080, new_n25081,
    new_n25082, new_n25083_1, new_n25084, new_n25085, new_n25086,
    new_n25087, new_n25088, new_n25089, new_n25090, new_n25091, new_n25092,
    new_n25093, new_n25094_1, new_n25095, new_n25096, new_n25097_1,
    new_n25098, new_n25099, new_n25100, new_n25101, new_n25102, new_n25103,
    new_n25104, new_n25105, new_n25106, new_n25107, new_n25108, new_n25109,
    new_n25111, new_n25113, new_n25114, new_n25115, new_n25116, new_n25117,
    new_n25118, new_n25119_1, new_n25120_1, new_n25121, new_n25122,
    new_n25123, new_n25124, new_n25125, new_n25126_1, new_n25128,
    new_n25130, new_n25132, new_n25134, new_n25136, new_n25137, new_n25138,
    new_n25139, new_n25140, new_n25141, new_n25142, new_n25143, new_n25144,
    new_n25145, new_n25146, new_n25147, new_n25148, new_n25149, new_n25150,
    new_n25151, new_n25152, new_n25153, new_n25154, new_n25155_1,
    new_n25156, new_n25157, new_n25158, new_n25159, new_n25160, new_n25161,
    new_n25162, new_n25163, new_n25164, new_n25165, new_n25166, new_n25167,
    new_n25168_1, new_n25169, new_n25170, new_n25171, new_n25172,
    new_n25173, new_n25174, new_n25175, new_n25176, new_n25177, new_n25178,
    new_n25179, new_n25180, new_n25181_1, new_n25182, new_n25183,
    new_n25184, new_n25185, new_n25186, new_n25187, new_n25188, new_n25189,
    new_n25190, new_n25191, new_n25192, new_n25193, new_n25194, new_n25195,
    new_n25196, new_n25197, new_n25198, new_n25199, new_n25200_1,
    new_n25201, new_n25202, new_n25203, new_n25204, new_n25205, new_n25206,
    new_n25207, new_n25208, new_n25209_1, new_n25210, new_n25211,
    new_n25212, new_n25213, new_n25214, new_n25215_1, new_n25216,
    new_n25217, new_n25218, new_n25219, new_n25220, new_n25221, new_n25222,
    new_n25223, new_n25225, new_n25226, new_n25227, new_n25228, new_n25229,
    new_n25230, new_n25231, new_n25232, new_n25233, new_n25235, new_n25237,
    new_n25238, new_n25239, new_n25240_1, new_n25241, new_n25242,
    new_n25244_1, new_n25246, new_n25248, new_n25250, new_n25252,
    new_n25253, new_n25254_1, new_n25255, new_n25256_1, new_n25257,
    new_n25258, new_n25259, new_n25260, new_n25261, new_n25262, new_n25263,
    new_n25264, new_n25265, new_n25266, new_n25267, new_n25268, new_n25269,
    new_n25270, new_n25271, new_n25272, new_n25273, new_n25274, new_n25275,
    new_n25276, new_n25277, new_n25278, new_n25279, new_n25280, new_n25281,
    new_n25282, new_n25283, new_n25284, new_n25285, new_n25286, new_n25287,
    new_n25288, new_n25289, new_n25290, new_n25291, new_n25292,
    new_n25293_1, new_n25294, new_n25295, new_n25296_1, new_n25297,
    new_n25298, new_n25299, new_n25300, new_n25301, new_n25302, new_n25303,
    new_n25304, new_n25305, new_n25306, new_n25307, new_n25308, new_n25309,
    new_n25310, new_n25311, new_n25312, new_n25313, new_n25314, new_n25315,
    new_n25316_1, new_n25317, new_n25318, new_n25319, new_n25320,
    new_n25321, new_n25322, new_n25323, new_n25325, new_n25327, new_n25329,
    new_n25331_1, new_n25333, new_n25335, new_n25337_1, new_n25338,
    new_n25339, new_n25340, new_n25341, new_n25342, new_n25344, new_n25346,
    new_n25348, new_n25350, new_n25351, new_n25353, new_n25355, new_n25357,
    new_n25358, new_n25359, new_n25360, new_n25361, new_n25362_1,
    new_n25363, new_n25364, new_n25365_1, new_n25366, new_n25367,
    new_n25368, new_n25369, new_n25370_1, new_n25371, new_n25372,
    new_n25373, new_n25374, new_n25375, new_n25376, new_n25377, new_n25378,
    new_n25379, new_n25380, new_n25381_1, new_n25382, new_n25383,
    new_n25384, new_n25385, new_n25386, new_n25387, new_n25388, new_n25389,
    new_n25390, new_n25391, new_n25392, new_n25393, new_n25394, new_n25395,
    new_n25396, new_n25397, new_n25398, new_n25399, new_n25400, new_n25401,
    new_n25403, new_n25405, new_n25406, new_n25408, new_n25410, new_n25413,
    new_n25417, new_n25418, new_n25419, new_n25420, new_n25421, new_n25422,
    new_n25423, new_n25424, new_n25425, new_n25426, new_n25427, new_n25429,
    new_n25432, new_n25434, new_n25436, new_n25439, new_n25441, new_n25443,
    new_n25445, new_n25446, new_n25447, new_n25448, new_n25449, new_n25450,
    new_n25451, new_n25452, new_n25453, new_n25454, new_n25455, new_n25456,
    new_n25457, new_n25458, new_n25459, new_n25460_1, new_n25462,
    new_n25463, new_n25464_1, new_n25465, new_n25466, new_n25467,
    new_n25468_1, new_n25469, new_n25470, new_n25471_1, new_n25472,
    new_n25473, new_n25474, new_n25475_1, new_n25476, new_n25477,
    new_n25481, new_n25483, new_n25485, new_n25486, new_n25487, new_n25488,
    new_n25489, new_n25490, new_n25491, new_n25492, new_n25493,
    new_n25494_1, new_n25495, new_n25496, new_n25497, new_n25498,
    new_n25499_1, new_n25500, new_n25501, new_n25502, new_n25503,
    new_n25504, new_n25505, new_n25506, new_n25507, new_n25508, new_n25509,
    new_n25511, new_n25513_1, new_n25514, new_n25515, new_n25516,
    new_n25517, new_n25518_1, new_n25519, new_n25520, new_n25521,
    new_n25522, new_n25523_1, new_n25524, new_n25525, new_n25526,
    new_n25527, new_n25528, new_n25529, new_n25530, new_n25531,
    new_n25532_1, new_n25533, new_n25534, new_n25535, new_n25536,
    new_n25537, new_n25538, new_n25539_1, new_n25540, new_n25541,
    new_n25542, new_n25544, new_n25545, new_n25546, new_n25547, new_n25548,
    new_n25549, new_n25550_1, new_n25551, new_n25552, new_n25553,
    new_n25556, new_n25558, new_n25559, new_n25561, new_n25562, new_n25564,
    new_n25566, new_n25568, new_n25570, new_n25571, new_n25572, new_n25573,
    new_n25574, new_n25575, new_n25576, new_n25577, new_n25578, new_n25579,
    new_n25580, new_n25581, new_n25582, new_n25583, new_n25584, new_n25585,
    new_n25586_1, new_n25587, new_n25588, new_n25589, new_n25590,
    new_n25591, new_n25592, new_n25593, new_n25594, new_n25595, new_n25596,
    new_n25597, new_n25598, new_n25599, new_n25600, new_n25601, new_n25602,
    new_n25603, new_n25604, new_n25605, new_n25606, new_n25607, new_n25608,
    new_n25609, new_n25610, new_n25611_1, new_n25612, new_n25613,
    new_n25614_1, new_n25615, new_n25616, new_n25617, new_n25618,
    new_n25619_1, new_n25621, new_n25622, new_n25623, new_n25624,
    new_n25625, new_n25626, new_n25627, new_n25628, new_n25629_1,
    new_n25630, new_n25631, new_n25632, new_n25633, new_n25634, new_n25635,
    new_n25636, new_n25637, new_n25638, new_n25639, new_n25640, new_n25641,
    new_n25642, new_n25643_1, new_n25644, new_n25645, new_n25646,
    new_n25647, new_n25648, new_n25649, new_n25650, new_n25651, new_n25652,
    new_n25653, new_n25654, new_n25655, new_n25656, new_n25657, new_n25658,
    new_n25659, new_n25660, new_n25661, new_n25662, new_n25663, new_n25664,
    new_n25665_1, new_n25666, new_n25667, new_n25668, new_n25669,
    new_n25670, new_n25671, new_n25672, new_n25673, new_n25674, new_n25675,
    new_n25676, new_n25677, new_n25678, new_n25679, new_n25680, new_n25681,
    new_n25682, new_n25684, new_n25686, new_n25688, new_n25690, new_n25692,
    new_n25694_1, new_n25696, new_n25698, new_n25700, new_n25702,
    new_n25704, new_n25706_1, new_n25708, new_n25709, new_n25710,
    new_n25711, new_n25712, new_n25714, new_n25716, new_n25719_1,
    new_n25721, new_n25723, new_n25725, new_n25727, new_n25729, new_n25731,
    new_n25733, new_n25734, new_n25735, new_n25736, new_n25737,
    new_n25738_1, new_n25739, new_n25740, new_n25741, new_n25742,
    new_n25743, new_n25744, new_n25745, new_n25746, new_n25747, new_n25748,
    new_n25749_1, new_n25750, new_n25751_1, new_n25752, new_n25753,
    new_n25754, new_n25755, new_n25756_1, new_n25757, new_n25758_1,
    new_n25759, new_n25760, new_n25761, new_n25762, new_n25763, new_n25764,
    new_n25765, new_n25766, new_n25767, new_n25768, new_n25769, new_n25770,
    new_n25771, new_n25772, new_n25773_1, new_n25775, new_n25777,
    new_n25778, new_n25779, new_n25780, new_n25781, new_n25782, new_n25783,
    new_n25784_1, new_n25785, new_n25786, new_n25787, new_n25788,
    new_n25789, new_n25790, new_n25792_1, new_n25794, new_n25797_1,
    new_n25799, new_n25801, new_n25802, new_n25803, new_n25804, new_n25805,
    new_n25806, new_n25807, new_n25808, new_n25809, new_n25810, new_n25811,
    new_n25812, new_n25813, new_n25814, new_n25815, new_n25816_1,
    new_n25817, new_n25818, new_n25819, new_n25820, new_n25821, new_n25822,
    new_n25823, new_n25824, new_n25825, new_n25826_1, new_n25827,
    new_n25828, new_n25829, new_n25830, new_n25831, new_n25832, new_n25833,
    new_n25834, new_n25835, new_n25836, new_n25837, new_n25838,
    new_n25839_1, new_n25840_1, new_n25841, new_n25842, new_n25843,
    new_n25844, new_n25845, new_n25846, new_n25847, new_n25848, new_n25849,
    new_n25850, new_n25851, new_n25852, new_n25853, new_n25854, new_n25855,
    new_n25856, new_n25857, new_n25858, new_n25859, new_n25860, new_n25861,
    new_n25862, new_n25863, new_n25864, new_n25865, new_n25866, new_n25867,
    new_n25868, new_n25869, new_n25870, new_n25871, new_n25872_1,
    new_n25873_1, new_n25874, new_n25875, new_n25876, new_n25877_1,
    new_n25878, new_n25879, new_n25880, new_n25881, new_n25882, new_n25883,
    new_n25884, new_n25885, new_n25886, new_n25887, new_n25888, new_n25889,
    new_n25890, new_n25891, new_n25892, new_n25893, new_n25894, new_n25895,
    new_n25896, new_n25897, new_n25898, new_n25899, new_n25900, new_n25901,
    new_n25902, new_n25903, new_n25904, new_n25905, new_n25906, new_n25907,
    new_n25908, new_n25909, new_n25910, new_n25911, new_n25912, new_n25913,
    new_n25914, new_n25915, new_n25916, new_n25917, new_n25918, new_n25919,
    new_n25920, new_n25921, new_n25922, new_n25923_1, new_n25924,
    new_n25925, new_n25926_1, new_n25927, new_n25928, new_n25929,
    new_n25930, new_n25931, new_n25932, new_n25933, new_n25934_1,
    new_n25935, new_n25936, new_n25937, new_n25938_1, new_n25939,
    new_n25941, new_n25943, new_n25945, new_n25947, new_n25949, new_n25950,
    new_n25951, new_n25952, new_n25953, new_n25954, new_n25955, new_n25956,
    new_n25957, new_n25958, new_n25959, new_n25960, new_n25961, new_n25962,
    new_n25963, new_n25964, new_n25965, new_n25967, new_n25969, new_n25971,
    new_n25973, new_n25974_1, new_n25975, new_n25976, new_n25977,
    new_n25978, new_n25979, new_n25980, new_n25981, new_n25982, new_n25983,
    new_n25984, new_n25985_1, new_n25986, new_n25987, new_n25988,
    new_n25989, new_n25990, new_n25991, new_n25992, new_n25993,
    new_n25994_1, new_n25995, new_n25996, new_n25997, new_n25998,
    new_n25999, new_n26001, new_n26002, new_n26003, new_n26004, new_n26006,
    new_n26008, new_n26010, new_n26011, new_n26012, new_n26014, new_n26016,
    new_n26018, new_n26020, new_n26023, new_n26025, new_n26027, new_n26029,
    new_n26030, new_n26031, new_n26032, new_n26033, new_n26034, new_n26035,
    new_n26036_1, new_n26037, new_n26038, new_n26039, new_n26040,
    new_n26041, new_n26042, new_n26043, new_n26044, new_n26045, new_n26046,
    new_n26047, new_n26048, new_n26049, new_n26050, new_n26051, new_n26052,
    new_n26053_1, new_n26054_1, new_n26055, new_n26057, new_n26059,
    new_n26061, new_n26063, new_n26065, new_n26067, new_n26069, new_n26071,
    new_n26073, new_n26075, new_n26077, new_n26079, new_n26081, new_n26083,
    new_n26085, new_n26087, new_n26090, new_n26092, new_n26094, new_n26095,
    new_n26096_1, new_n26097, new_n26098, new_n26099, new_n26100,
    new_n26101, new_n26102, new_n26103, new_n26104, new_n26105, new_n26106,
    new_n26107_1, new_n26108, new_n26109, new_n26110, new_n26111_1,
    new_n26112, new_n26113_1, new_n26114, new_n26115, new_n26116,
    new_n26117, new_n26118, new_n26119, new_n26120, new_n26121, new_n26122,
    new_n26123, new_n26124, new_n26125, new_n26126, new_n26127, new_n26128,
    new_n26129, new_n26130, new_n26131, new_n26132, new_n26133, new_n26134,
    new_n26136, new_n26138, new_n26140, new_n26142, new_n26144, new_n26146,
    new_n26148, new_n26149, new_n26150, new_n26151, new_n26152, new_n26153,
    new_n26154, new_n26155, new_n26156_1, new_n26157, new_n26158,
    new_n26159_1, new_n26160, new_n26163, new_n26165, new_n26166,
    new_n26168, new_n26170, new_n26171, new_n26172, new_n26173, new_n26174,
    new_n26175, new_n26178, new_n26179_1, new_n26180_1, new_n26181,
    new_n26182, new_n26183, new_n26184, new_n26185, new_n26186, new_n26187,
    new_n26188, new_n26189, new_n26190, new_n26191_1, new_n26192,
    new_n26193, new_n26194, new_n26195, new_n26197, new_n26199, new_n26200,
    new_n26201, new_n26202, new_n26203, new_n26204, new_n26205, new_n26206,
    new_n26207, new_n26208, new_n26209, new_n26210, new_n26211, new_n26212,
    new_n26213, new_n26214, new_n26215, new_n26216, new_n26217, new_n26218,
    new_n26219, new_n26220_1, new_n26221, new_n26222, new_n26223,
    new_n26224_1, new_n26225, new_n26226, new_n26227, new_n26228,
    new_n26229_1, new_n26230, new_n26231, new_n26232, new_n26233,
    new_n26234, new_n26235, new_n26236, new_n26237_1, new_n26238,
    new_n26240, new_n26242, new_n26244, new_n26246, new_n26248,
    new_n26250_1, new_n26252, new_n26254, new_n26256, new_n26259,
    new_n26262, new_n26264_1, new_n26266, new_n26268, new_n26271,
    new_n26273, new_n26275, new_n26277, new_n26279, new_n26281, new_n26282,
    new_n26283, new_n26284, new_n26285, new_n26286, new_n26287_1,
    new_n26288, new_n26289, new_n26290, new_n26291, new_n26292, new_n26294,
    new_n26296, new_n26297, new_n26298, new_n26299, new_n26300, new_n26301,
    new_n26302, new_n26303, new_n26304, new_n26305, new_n26306, new_n26307,
    new_n26308, new_n26309, new_n26310, new_n26311, new_n26312, new_n26313,
    new_n26315, new_n26317_1, new_n26319, new_n26320, new_n26321,
    new_n26322, new_n26323, new_n26325, new_n26327, new_n26329, new_n26333,
    new_n26335, new_n26336, new_n26337, new_n26338, new_n26339, new_n26340,
    new_n26341, new_n26342, new_n26344, new_n26345, new_n26346, new_n26347,
    new_n26348, new_n26349, new_n26350, new_n26351, new_n26352,
    new_n26353_1, new_n26354, new_n26355, new_n26356, new_n26357,
    new_n26358, new_n26359, new_n26360, new_n26361, new_n26362, new_n26363,
    new_n26364, new_n26365, new_n26366, new_n26368, new_n26370, new_n26372,
    new_n26374, new_n26376, new_n26378, new_n26380, new_n26382, new_n26384,
    new_n26386, new_n26388, new_n26390, new_n26392, new_n26394,
    new_n26396_1, new_n26398, new_n26400, new_n26402, new_n26404,
    new_n26406, new_n26408_1, new_n26410, new_n26411, new_n26412,
    new_n26413, new_n26414, new_n26415, new_n26416, new_n26417, new_n26418,
    new_n26419, new_n26420, new_n26421, new_n26422, new_n26423, new_n26424,
    new_n26425, new_n26426, new_n26428, new_n26430, new_n26432, new_n26434,
    new_n26435, new_n26436, new_n26437, new_n26438, new_n26440, new_n26442,
    new_n26444, new_n26446, new_n26448, new_n26450, new_n26452_1,
    new_n26454, new_n26456, new_n26458, new_n26460, new_n26462, new_n26464,
    new_n26466, new_n26468, new_n26471, new_n26473, new_n26475, new_n26477,
    new_n26479, new_n26481, new_n26484, new_n26487, new_n26489, new_n26490,
    new_n26491, new_n26492_1, new_n26493, new_n26495, new_n26497,
    new_n26499, new_n26501, new_n26503, new_n26505, new_n26507, new_n26509,
    new_n26511, new_n26513, new_n26515_1, new_n26517, new_n26519,
    new_n26520, new_n26521, new_n26522, new_n26523, new_n26524, new_n26526,
    new_n26528, new_n26530, new_n26531, new_n26532, new_n26533, new_n26534,
    new_n26535, new_n26538_1, new_n26540, new_n26542, new_n26543,
    new_n26544, new_n26545, new_n26546, new_n26547, new_n26548, new_n26549,
    new_n26551, new_n26553_1, new_n26555, new_n26557, new_n26559,
    new_n26561, new_n26563, new_n26565_1, new_n26568, new_n26570,
    new_n26572_1, new_n26574, new_n26576, new_n26578, new_n26580,
    new_n26581, new_n26582, new_n26585, new_n26586, new_n26587,
    new_n26590_1, new_n26592, new_n26594, new_n26596, new_n26598_1,
    new_n26600, new_n26604, new_n26606, new_n26608, new_n26610, new_n26612,
    new_n26614, new_n26616, new_n26619, new_n26621, new_n26624, new_n26626,
    new_n26628, new_n26630, new_n26631, new_n26632, new_n26633, new_n26634,
    new_n26635, new_n26637, new_n26639, new_n26641, new_n26645, new_n26648,
    new_n26649, new_n26650, new_n26651, new_n26652, new_n26653, new_n26654,
    new_n26655, new_n26656_1, new_n26658, new_n26659, new_n26661,
    new_n26664, new_n26666, new_n26668, new_n26670, new_n26672,
    new_n26674_1, new_n26676, new_n26678, new_n26680, new_n26681_1,
    new_n26682, new_n26683, new_n26684, new_n26685, new_n26686, new_n26687,
    new_n26688, new_n26689, new_n26690, new_n26691, new_n26693, new_n26695,
    new_n26697, new_n26699, new_n26701, new_n26703, new_n26705,
    new_n26707_1, new_n26709, new_n26711, new_n26713, new_n26715,
    new_n26717, new_n26719_1, new_n26721, new_n26723, new_n26725_1,
    new_n26726, new_n26727_1, new_n26728, new_n26729_1, new_n26730,
    new_n26731, new_n26732, new_n26733, new_n26734, new_n26735, new_n26736,
    new_n26737, new_n26738, new_n26739, new_n26741, new_n26743,
    new_n26744_1, new_n26746, new_n26750, new_n26751, new_n26752_1,
    new_n26753, new_n26756, new_n26758, new_n26760, new_n26761, new_n26762,
    new_n26763, new_n26764, new_n26766, new_n26767, new_n26768, new_n26769,
    new_n26770, new_n26771, new_n26772, new_n26773, new_n26774,
    new_n26775_1, new_n26776, new_n26777, new_n26778, new_n26779,
    new_n26780_1, new_n26781, new_n26782, new_n26783, new_n26784,
    new_n26785, new_n26786, new_n26787, new_n26788, new_n26789, new_n26790,
    new_n26792, new_n26794_1, new_n26796, new_n26797_1, new_n26798,
    new_n26799, new_n26801_1, new_n26803, new_n26805, new_n26807,
    new_n26809, new_n26811, new_n26813, new_n26815_1, new_n26817,
    new_n26819, new_n26821, new_n26823_1, new_n26825, new_n26827,
    new_n26829, new_n26832, new_n26834, new_n26836, new_n26838, new_n26840,
    new_n26842, new_n26844, new_n26846, new_n26848, new_n26850, new_n26852,
    new_n26854, new_n26856, new_n26857, new_n26858, new_n26859, new_n26860,
    new_n26862, new_n26864, new_n26865, new_n26867, new_n26869, new_n26871,
    new_n26874, new_n26876, new_n26878, new_n26880, new_n26882_1,
    new_n26884, new_n26887, new_n26889, new_n26891, new_n26893, new_n26895,
    new_n26897, new_n26899, new_n26901, new_n26903, new_n26905_1,
    new_n26907, new_n26910, new_n26913_1, new_n26915, new_n26917,
    new_n26919, new_n26921_1, new_n26923_1, new_n26925, new_n26927,
    new_n26929_1, new_n26931, new_n26933, new_n26935, new_n26937,
    new_n26939, new_n26941, new_n26943_1, new_n26945, new_n26947,
    new_n26949, new_n26950, new_n26952, new_n26954, new_n26956, new_n26958,
    new_n26960, new_n26962, new_n26964, new_n26966, new_n26968,
    new_n26970_1, new_n26974, new_n26975, new_n26976, new_n26977,
    new_n26978, new_n26979_1, new_n26980, new_n26982, new_n26984,
    new_n26986_1, new_n26988, new_n26990, new_n26992, new_n26994,
    new_n26996, new_n26998, new_n27000, new_n27002, new_n27004_1,
    new_n27006, new_n27007, new_n27008, new_n27009, new_n27010,
    new_n27011_1, new_n27012, new_n27013, new_n27014, new_n27015,
    new_n27017, new_n27019_1, new_n27021, new_n27023, new_n27025,
    new_n27026, new_n27027, new_n27028, new_n27029, new_n27030, new_n27032,
    new_n27034, new_n27035, new_n27036, new_n27038, new_n27040, new_n27042,
    new_n27044, new_n27046, new_n27048, new_n27049, new_n27050,
    new_n27051_1, new_n27052, new_n27053, new_n27054, new_n27055,
    new_n27056, new_n27057, new_n27058, new_n27059, new_n27060, new_n27062,
    new_n27065, new_n27067, new_n27069, new_n27071, new_n27073, new_n27075,
    new_n27077, new_n27079_1, new_n27081, new_n27083, new_n27085,
    new_n27087, new_n27089_1, new_n27091, new_n27093, new_n27095,
    new_n27097, new_n27099, new_n27101, new_n27103, new_n27105, new_n27107,
    new_n27109, new_n27111, new_n27113, new_n27115, new_n27117, new_n27119,
    new_n27121, new_n27123, new_n27125, new_n27127, new_n27129, new_n27131,
    new_n27133, new_n27135, new_n27137, new_n27139, new_n27141, new_n27143,
    new_n27146, new_n27148, new_n27150, new_n27152, new_n27154, new_n27156,
    new_n27158_1, new_n27160, new_n27162, new_n27164, new_n27165,
    new_n27167, new_n27169, new_n27171, new_n27173, new_n27175, new_n27177,
    new_n27179, new_n27181, new_n27183, new_n27185, new_n27187, new_n27189,
    new_n27191, new_n27193, new_n27195, new_n27197, new_n27199, new_n27201,
    new_n27203, new_n27205, new_n27206, new_n27207, new_n27208, new_n27209,
    new_n27210, new_n27211, new_n27212, new_n27213, new_n27214, new_n27215,
    new_n27216, new_n27218, new_n27220, new_n27222, new_n27224, new_n27226,
    new_n27228, new_n27230, new_n27232, new_n27234, new_n27236, new_n27238,
    new_n27240, new_n27242, new_n27244, new_n27245, new_n27246, new_n27247,
    new_n27248, new_n27249, new_n27251, new_n27252, new_n27254, new_n27256,
    new_n27258, new_n27259, new_n27261, new_n27263, new_n27265, new_n27267,
    new_n27269, new_n27270, new_n27271, new_n27272, new_n27273, new_n27274,
    new_n27275, new_n27276, new_n27277, new_n27278, new_n27279, new_n27280,
    new_n27282, new_n27284, new_n27286, new_n27288, new_n27290, new_n27291,
    new_n27293, new_n27295, new_n27298, new_n27300, new_n27302, new_n27304,
    new_n27305, new_n27306, new_n27308, new_n27310, new_n27312, new_n27314,
    new_n27316, new_n27318, new_n27320, new_n27321, new_n27323, new_n27325,
    new_n27327, new_n27329, new_n27331, new_n27333, new_n27334, new_n27335,
    new_n27336, new_n27337, new_n27338, new_n27339, new_n27341, new_n27343,
    new_n27345, new_n27347, new_n27349, new_n27351, new_n27353, new_n27355,
    new_n27357, new_n27359, new_n27361, new_n27363, new_n27364, new_n27365,
    new_n27367, new_n27369, new_n27371, new_n27373, new_n27374, new_n27375,
    new_n27376, new_n27379, new_n27381, new_n27383, new_n27386, new_n27388,
    new_n27390, new_n27392, new_n27394, new_n27396, new_n27398, new_n27399,
    new_n27401, new_n27403, new_n27405, new_n27407, new_n27409, new_n27411,
    new_n27413, new_n27415, new_n27417, new_n27419, new_n27421, new_n27422,
    new_n27424, new_n27426, new_n27428, new_n27430, new_n27432, new_n27434,
    new_n27436, new_n27438, new_n27440, new_n27441, new_n27442, new_n27443,
    new_n27444, new_n27445, new_n27446, new_n27447, new_n27449, new_n27451,
    new_n27453, new_n27455, new_n27457, new_n27458, new_n27460, new_n27461,
    new_n27462, new_n27463, new_n27465, new_n27467, new_n27469, new_n27471,
    new_n27472, new_n27473, new_n27474, new_n27475, new_n27476, new_n27477,
    new_n27478, new_n27479, new_n27480, new_n27481, new_n27482, new_n27483,
    new_n27484, new_n27485, new_n27486, new_n27487, new_n27488, new_n27489,
    new_n27490, new_n27491, new_n27492, new_n27494, new_n27496, new_n27498,
    new_n27500, new_n27501, new_n27502, new_n27503, new_n27505, new_n27507,
    new_n27509, new_n27510, new_n27511, new_n27513, new_n27515, new_n27517,
    new_n27519, new_n27521, new_n27524, new_n27526, new_n27528, new_n27529,
    new_n27531, new_n27534, new_n27536, new_n27538, new_n27541, new_n27543,
    new_n27545, new_n27547, new_n27549, new_n27552, new_n27554, new_n27556,
    new_n27558, new_n27560, new_n27562, new_n27563, new_n27564, new_n27565,
    new_n27566, new_n27568, new_n27569, new_n27570, new_n27571, new_n27572,
    new_n27574, new_n27577, new_n27579, new_n27581, new_n27583, new_n27585,
    new_n27587, new_n27589, new_n27591, new_n27593, new_n27595, new_n27597,
    new_n27599, new_n27601, new_n27603, new_n27605, new_n27607, new_n27609,
    new_n27611, new_n27613, new_n27614, new_n27616, new_n27618, new_n27620,
    new_n27621, new_n27622, new_n27623, new_n27625, new_n27626, new_n27629,
    new_n27631, new_n27633, new_n27635, new_n27637, new_n27639, new_n27641,
    new_n27643, new_n27645, new_n27646, new_n27647, new_n27648, new_n27650,
    new_n27652, new_n27654, new_n27656, new_n27658, new_n27660, new_n27662,
    new_n27665, new_n27668, new_n27670, new_n27672, new_n27674, new_n27676,
    new_n27678, new_n27681, new_n27683, new_n27685, new_n27687, new_n27689,
    new_n27691, new_n27695, new_n27697, new_n27699, new_n27701, new_n27703,
    new_n27706, new_n27708, new_n27709, new_n27711, new_n27713, new_n27715,
    new_n27717, new_n27719, new_n27721, new_n27723, new_n27726, new_n27727,
    new_n27729, new_n27731, new_n27733, new_n27735, new_n27737, new_n27739,
    new_n27741, new_n27742, new_n27744, new_n27746, new_n27749, new_n27751,
    new_n27753, new_n27755, new_n27757, new_n27759, new_n27761, new_n27763,
    new_n27765, new_n27766, new_n27768, new_n27770, new_n27772, new_n27775,
    new_n27777, new_n27779, new_n27781, new_n27783, new_n27786, new_n27788,
    new_n27790, new_n27792, new_n27794, new_n27796, new_n27798, new_n27800,
    new_n27802, new_n27804, new_n27806, new_n27808, new_n27810, new_n27812,
    new_n27814, new_n27816, new_n27818, new_n27820, new_n27822, new_n27824,
    new_n27826, new_n27828, new_n27831, new_n27833, new_n27835, new_n27837,
    new_n27839, new_n27841, new_n27843, new_n27845, new_n27847, new_n27849,
    new_n27851, new_n27853, new_n27855, new_n27857, new_n27859, new_n27861,
    new_n27864, new_n27866, new_n27869, new_n27871, new_n27873, new_n27875,
    new_n27877, new_n27879, new_n27881, new_n27882, new_n27884, new_n27886,
    new_n27888, new_n27890, new_n27892, new_n27895, new_n27897, new_n27899,
    new_n27901, new_n27903, new_n27905, new_n27907, new_n27909, new_n27911,
    new_n27913, new_n27915, new_n27917, new_n27919, new_n27921, new_n27923,
    new_n27925, new_n27927, new_n27929, new_n27932, new_n27934, new_n27936,
    new_n27938, new_n27941, new_n27943, new_n27945, new_n27947, new_n27949,
    new_n27951, new_n27953, new_n27955, new_n27957, new_n27959, new_n27961,
    new_n27963, new_n27965, new_n27967, new_n27969, new_n27971, new_n27972,
    new_n27973, new_n27975, new_n27977, new_n27979, new_n27981, new_n27982,
    new_n27984, new_n27986, new_n27988, new_n27990, new_n27992, new_n27995,
    new_n27997, new_n28000, new_n28002, new_n28005, new_n28007, new_n28010,
    new_n28012, new_n28014, new_n28016, new_n28019, new_n28020, new_n28022,
    new_n28024, new_n28026, new_n28028, new_n28030, new_n28032, new_n28033,
    new_n28035, new_n28037, new_n28040, new_n28042, new_n28044, new_n28046,
    new_n28048, new_n28050, new_n28052, new_n28054, new_n28056, new_n28058,
    new_n28060, new_n28062, new_n28064, new_n28065, new_n28067, new_n28069,
    new_n28071, new_n28073, new_n28075, new_n28076, new_n28078, new_n28080,
    new_n28082, new_n28085, new_n28087, new_n28089, new_n28091, new_n28093,
    new_n28095, new_n28097, new_n28099, new_n28101, new_n28103, new_n28105,
    new_n28107, new_n28109, new_n28111, new_n28113, new_n28115, new_n28117,
    new_n28119, new_n28121, new_n28123, new_n28126, new_n28128, new_n28131,
    new_n28133, new_n28134, new_n28136, new_n28138;
  not_8  g00000(.A(n8745), .Y(new_n2349));
  not_8  g00001(.A(n24278), .Y(new_n2350));
  nand_5 g00002(.A(new_n2350), .B(new_n2349), .Y(new_n2351));
  nand_5 g00003(.A(n24278), .B(n8745), .Y(new_n2352));
  not_8  g00004(.A(n15636), .Y(new_n2353));
  not_8  g00005(.A(n24618), .Y(new_n2354));
  nand_5 g00006(.A(new_n2354), .B(new_n2353), .Y(new_n2355_1));
  nand_5 g00007(.A(n24618), .B(n15636), .Y(new_n2356));
  not_8  g00008(.A(n3952), .Y(new_n2357));
  not_8  g00009(.A(n20077), .Y(new_n2358));
  nand_5 g00010(.A(new_n2358), .B(new_n2357), .Y(new_n2359));
  nand_5 g00011(.A(n20077), .B(n3952), .Y(new_n2360));
  nand_5 g00012(.A(n12315), .B(n6794), .Y(new_n2361_1));
  nand_5 g00013(.A(new_n2361_1), .B(new_n2360), .Y(new_n2362));
  nand_5 g00014(.A(new_n2362), .B(new_n2359), .Y(new_n2363_1));
  nand_5 g00015(.A(new_n2363_1), .B(new_n2356), .Y(new_n2364));
  nand_5 g00016(.A(new_n2364), .B(new_n2355_1), .Y(new_n2365));
  nand_5 g00017(.A(new_n2365), .B(new_n2352), .Y(new_n2366));
  nand_5 g00018(.A(new_n2366), .B(new_n2351), .Y(new_n2367));
  not_8  g00019(.A(new_n2367), .Y(new_n2368));
  nand_5 g00020(.A(n4812), .B(n1777), .Y(new_n2369));
  not_8  g00021(.A(n1777), .Y(new_n2370));
  not_8  g00022(.A(n4812), .Y(new_n2371));
  nand_5 g00023(.A(new_n2371), .B(new_n2370), .Y(new_n2372));
  nand_5 g00024(.A(new_n2372), .B(new_n2369), .Y(new_n2373));
  xor_4  g00025(.A(new_n2373), .B(new_n2368), .Y(new_n2374_1));
  not_8  g00026(.A(new_n2374_1), .Y(new_n2375));
  nand_5 g00027(.A(n13781), .B(n5704), .Y(new_n2376));
  not_8  g00028(.A(n5704), .Y(new_n2377));
  not_8  g00029(.A(n13781), .Y(new_n2378));
  nand_5 g00030(.A(new_n2378), .B(new_n2377), .Y(new_n2379));
  nand_5 g00031(.A(new_n2379), .B(new_n2376), .Y(new_n2380));
  not_8  g00032(.A(new_n2376), .Y(new_n2381));
  nand_5 g00033(.A(n18409), .B(n11486), .Y(new_n2382));
  not_8  g00034(.A(n11486), .Y(new_n2383));
  not_8  g00035(.A(n18409), .Y(new_n2384));
  nand_5 g00036(.A(new_n2384), .B(new_n2383), .Y(new_n2385));
  nand_5 g00037(.A(new_n2385), .B(new_n2382), .Y(new_n2386));
  xor_4  g00038(.A(new_n2386), .B(new_n2381), .Y(new_n2387_1));
  nand_5 g00039(.A(new_n2387_1), .B(new_n2380), .Y(new_n2388_1));
  nand_5 g00040(.A(new_n2382), .B(new_n2376), .Y(new_n2389));
  nand_5 g00041(.A(new_n2389), .B(new_n2385), .Y(new_n2390));
  not_8  g00042(.A(new_n2390), .Y(new_n2391));
  nand_5 g00043(.A(n16722), .B(n13708), .Y(new_n2392));
  not_8  g00044(.A(n13708), .Y(new_n2393));
  not_8  g00045(.A(n16722), .Y(new_n2394));
  nand_5 g00046(.A(new_n2394), .B(new_n2393), .Y(new_n2395));
  nand_5 g00047(.A(new_n2395), .B(new_n2392), .Y(new_n2396));
  xor_4  g00048(.A(new_n2396), .B(new_n2391), .Y(new_n2397));
  not_8  g00049(.A(new_n2397), .Y(new_n2398));
  nor_5  g00050(.A(new_n2398), .B(new_n2388_1), .Y(new_n2399));
  nand_5 g00051(.A(n19911), .B(n3480), .Y(new_n2400));
  not_8  g00052(.A(n3480), .Y(new_n2401));
  not_8  g00053(.A(n19911), .Y(new_n2402));
  nand_5 g00054(.A(new_n2402), .B(new_n2401), .Y(new_n2403));
  nand_5 g00055(.A(new_n2403), .B(new_n2400), .Y(new_n2404));
  nand_5 g00056(.A(new_n2392), .B(new_n2390), .Y(new_n2405));
  nand_5 g00057(.A(new_n2405), .B(new_n2395), .Y(new_n2406));
  not_8  g00058(.A(new_n2406), .Y(new_n2407));
  xor_4  g00059(.A(new_n2407), .B(new_n2404), .Y(new_n2408));
  nand_5 g00060(.A(new_n2408), .B(new_n2399), .Y(new_n2409_1));
  nand_5 g00061(.A(n3018), .B(n2731), .Y(new_n2410));
  not_8  g00062(.A(n2731), .Y(new_n2411));
  not_8  g00063(.A(n3018), .Y(new_n2412));
  nand_5 g00064(.A(new_n2412), .B(new_n2411), .Y(new_n2413));
  nand_5 g00065(.A(new_n2413), .B(new_n2410), .Y(new_n2414));
  nand_5 g00066(.A(new_n2406), .B(new_n2400), .Y(new_n2415));
  nand_5 g00067(.A(new_n2415), .B(new_n2403), .Y(new_n2416_1));
  not_8  g00068(.A(new_n2416_1), .Y(new_n2417));
  xor_4  g00069(.A(new_n2417), .B(new_n2414), .Y(new_n2418));
  not_8  g00070(.A(new_n2418), .Y(new_n2419));
  nor_5  g00071(.A(new_n2419), .B(new_n2409_1), .Y(new_n2420_1));
  not_8  g00072(.A(new_n2420_1), .Y(new_n2421_1));
  nand_5 g00073(.A(new_n2419), .B(new_n2409_1), .Y(new_n2422));
  and_5  g00074(.A(new_n2422), .B(new_n2421_1), .Y(new_n2423));
  nand_5 g00075(.A(new_n2423), .B(new_n2375), .Y(new_n2424));
  or_5   g00076(.A(new_n2423), .B(new_n2375), .Y(new_n2425));
  not_8  g00077(.A(new_n2399), .Y(new_n2426));
  not_8  g00078(.A(new_n2408), .Y(new_n2427));
  nand_5 g00079(.A(new_n2427), .B(new_n2426), .Y(new_n2428));
  and_5  g00080(.A(new_n2428), .B(new_n2409_1), .Y(new_n2429));
  nand_5 g00081(.A(new_n2352), .B(new_n2351), .Y(new_n2430));
  xor_4  g00082(.A(new_n2430), .B(new_n2365), .Y(new_n2431));
  nand_5 g00083(.A(new_n2431), .B(new_n2429), .Y(new_n2432));
  or_5   g00084(.A(new_n2431), .B(new_n2429), .Y(new_n2433));
  nand_5 g00085(.A(new_n2398), .B(new_n2388_1), .Y(new_n2434));
  nand_5 g00086(.A(new_n2434), .B(new_n2426), .Y(new_n2435));
  nand_5 g00087(.A(new_n2356), .B(new_n2355_1), .Y(new_n2436));
  xor_4  g00088(.A(new_n2436), .B(new_n2363_1), .Y(new_n2437));
  not_8  g00089(.A(new_n2437), .Y(new_n2438));
  or_5   g00090(.A(new_n2438), .B(new_n2435), .Y(new_n2439));
  nand_5 g00091(.A(new_n2438), .B(new_n2435), .Y(new_n2440_1));
  not_8  g00092(.A(new_n2380), .Y(new_n2441));
  not_8  g00093(.A(n6794), .Y(new_n2442));
  not_8  g00094(.A(n12315), .Y(new_n2443));
  nand_5 g00095(.A(new_n2443), .B(new_n2442), .Y(new_n2444_1));
  and_5  g00096(.A(new_n2444_1), .B(new_n2361_1), .Y(new_n2445));
  nand_5 g00097(.A(new_n2445), .B(new_n2441), .Y(new_n2446));
  nand_5 g00098(.A(new_n2360), .B(new_n2359), .Y(new_n2447));
  nor_5  g00099(.A(new_n2447), .B(new_n2446), .Y(new_n2448));
  not_8  g00100(.A(new_n2448), .Y(new_n2449));
  xor_4  g00101(.A(new_n2447), .B(new_n2361_1), .Y(new_n2450));
  not_8  g00102(.A(new_n2450), .Y(new_n2451));
  nand_5 g00103(.A(new_n2451), .B(new_n2446), .Y(new_n2452));
  xor_4  g00104(.A(new_n2387_1), .B(new_n2441), .Y(new_n2453));
  not_8  g00105(.A(new_n2453), .Y(new_n2454));
  nand_5 g00106(.A(new_n2454), .B(new_n2452), .Y(new_n2455));
  nand_5 g00107(.A(new_n2455), .B(new_n2449), .Y(new_n2456));
  nand_5 g00108(.A(new_n2456), .B(new_n2440_1), .Y(new_n2457));
  nand_5 g00109(.A(new_n2457), .B(new_n2439), .Y(new_n2458));
  nand_5 g00110(.A(new_n2458), .B(new_n2433), .Y(new_n2459));
  nand_5 g00111(.A(new_n2459), .B(new_n2432), .Y(new_n2460));
  nand_5 g00112(.A(new_n2460), .B(new_n2425), .Y(new_n2461));
  nand_5 g00113(.A(new_n2461), .B(new_n2424), .Y(new_n2462));
  nand_5 g00114(.A(new_n2369), .B(new_n2367), .Y(new_n2463));
  nand_5 g00115(.A(new_n2463), .B(new_n2372), .Y(new_n2464));
  not_8  g00116(.A(new_n2464), .Y(new_n2465));
  nand_5 g00117(.A(n26823), .B(n22660), .Y(new_n2466));
  not_8  g00118(.A(n22660), .Y(new_n2467));
  not_8  g00119(.A(n26823), .Y(new_n2468));
  nand_5 g00120(.A(new_n2468), .B(new_n2467), .Y(new_n2469));
  nand_5 g00121(.A(new_n2469), .B(new_n2466), .Y(new_n2470));
  xor_4  g00122(.A(new_n2470), .B(new_n2465), .Y(new_n2471));
  not_8  g00123(.A(new_n2471), .Y(new_n2472));
  nand_5 g00124(.A(n26660), .B(n18907), .Y(new_n2473));
  not_8  g00125(.A(n18907), .Y(new_n2474));
  not_8  g00126(.A(n26660), .Y(new_n2475));
  nand_5 g00127(.A(new_n2475), .B(new_n2474), .Y(new_n2476));
  nand_5 g00128(.A(new_n2476), .B(new_n2473), .Y(new_n2477));
  nand_5 g00129(.A(new_n2416_1), .B(new_n2410), .Y(new_n2478));
  nand_5 g00130(.A(new_n2478), .B(new_n2413), .Y(new_n2479_1));
  not_8  g00131(.A(new_n2479_1), .Y(new_n2480));
  xor_4  g00132(.A(new_n2480), .B(new_n2477), .Y(new_n2481));
  nand_5 g00133(.A(new_n2481), .B(new_n2420_1), .Y(new_n2482));
  not_8  g00134(.A(new_n2481), .Y(new_n2483));
  nand_5 g00135(.A(new_n2483), .B(new_n2421_1), .Y(new_n2484));
  and_5  g00136(.A(new_n2484), .B(new_n2482), .Y(new_n2485));
  nand_5 g00137(.A(new_n2485), .B(new_n2472), .Y(new_n2486));
  or_5   g00138(.A(new_n2485), .B(new_n2472), .Y(new_n2487));
  nand_5 g00139(.A(new_n2487), .B(new_n2486), .Y(new_n2488));
  xor_4  g00140(.A(new_n2488), .B(new_n2462), .Y(new_n2489));
  not_8  g00141(.A(n9557), .Y(new_n2490));
  nand_5 g00142(.A(n21832), .B(new_n2490), .Y(new_n2491));
  not_8  g00143(.A(n21832), .Y(new_n2492));
  nand_5 g00144(.A(new_n2492), .B(n9557), .Y(new_n2493));
  not_8  g00145(.A(n3136), .Y(new_n2494));
  nand_5 g00146(.A(n26913), .B(new_n2494), .Y(new_n2495));
  not_8  g00147(.A(n26913), .Y(new_n2496));
  nand_5 g00148(.A(new_n2496), .B(n3136), .Y(new_n2497));
  not_8  g00149(.A(n6385), .Y(new_n2498));
  nand_5 g00150(.A(n16223), .B(new_n2498), .Y(new_n2499));
  not_8  g00151(.A(n16223), .Y(new_n2500));
  nand_5 g00152(.A(new_n2500), .B(n6385), .Y(new_n2501));
  not_8  g00153(.A(n20138), .Y(new_n2502));
  nand_5 g00154(.A(new_n2502), .B(n19494), .Y(new_n2503));
  not_8  g00155(.A(n19494), .Y(new_n2504));
  nand_5 g00156(.A(n20138), .B(new_n2504), .Y(new_n2505));
  not_8  g00157(.A(n2387), .Y(new_n2506));
  nand_5 g00158(.A(n9251), .B(new_n2506), .Y(new_n2507));
  nand_5 g00159(.A(new_n2507), .B(new_n2505), .Y(new_n2508));
  nand_5 g00160(.A(new_n2508), .B(new_n2503), .Y(new_n2509));
  nand_5 g00161(.A(new_n2509), .B(new_n2501), .Y(new_n2510));
  nand_5 g00162(.A(new_n2510), .B(new_n2499), .Y(new_n2511));
  nand_5 g00163(.A(new_n2511), .B(new_n2497), .Y(new_n2512));
  nand_5 g00164(.A(new_n2512), .B(new_n2495), .Y(new_n2513_1));
  nand_5 g00165(.A(new_n2513_1), .B(new_n2493), .Y(new_n2514));
  nand_5 g00166(.A(new_n2514), .B(new_n2491), .Y(new_n2515_1));
  not_8  g00167(.A(n25643), .Y(new_n2516));
  nand_5 g00168(.A(new_n2516), .B(n21753), .Y(new_n2517));
  not_8  g00169(.A(n21753), .Y(new_n2518));
  nand_5 g00170(.A(n25643), .B(new_n2518), .Y(new_n2519));
  nand_5 g00171(.A(new_n2519), .B(new_n2517), .Y(new_n2520));
  xor_4  g00172(.A(new_n2520), .B(new_n2515_1), .Y(new_n2521));
  nand_5 g00173(.A(new_n2521), .B(new_n2489), .Y(new_n2522));
  not_8  g00174(.A(new_n2522), .Y(new_n2523));
  nor_5  g00175(.A(new_n2521), .B(new_n2489), .Y(new_n2524));
  nand_5 g00176(.A(new_n2425), .B(new_n2424), .Y(new_n2525));
  xor_4  g00177(.A(new_n2525), .B(new_n2460), .Y(new_n2526));
  nand_5 g00178(.A(new_n2493), .B(new_n2491), .Y(new_n2527));
  xor_4  g00179(.A(new_n2527), .B(new_n2513_1), .Y(new_n2528));
  or_5   g00180(.A(new_n2528), .B(new_n2526), .Y(new_n2529));
  nand_5 g00181(.A(new_n2528), .B(new_n2526), .Y(new_n2530));
  nand_5 g00182(.A(new_n2433), .B(new_n2432), .Y(new_n2531));
  xor_4  g00183(.A(new_n2531), .B(new_n2458), .Y(new_n2532));
  nand_5 g00184(.A(new_n2497), .B(new_n2495), .Y(new_n2533_1));
  xor_4  g00185(.A(new_n2533_1), .B(new_n2511), .Y(new_n2534));
  or_5   g00186(.A(new_n2534), .B(new_n2532), .Y(new_n2535_1));
  nand_5 g00187(.A(new_n2534), .B(new_n2532), .Y(new_n2536));
  nand_5 g00188(.A(new_n2440_1), .B(new_n2439), .Y(new_n2537_1));
  xor_4  g00189(.A(new_n2537_1), .B(new_n2456), .Y(new_n2538));
  nand_5 g00190(.A(new_n2501), .B(new_n2499), .Y(new_n2539));
  xor_4  g00191(.A(new_n2539), .B(new_n2509), .Y(new_n2540));
  or_5   g00192(.A(new_n2540), .B(new_n2538), .Y(new_n2541));
  nand_5 g00193(.A(new_n2540), .B(new_n2538), .Y(new_n2542));
  xor_4  g00194(.A(new_n2445), .B(new_n2441), .Y(new_n2543));
  not_8  g00195(.A(new_n2543), .Y(new_n2544));
  xor_4  g00196(.A(n9251), .B(new_n2506), .Y(new_n2545));
  nor_5  g00197(.A(new_n2545), .B(new_n2544), .Y(new_n2546));
  nand_5 g00198(.A(new_n2505), .B(new_n2503), .Y(new_n2547_1));
  xnor_4 g00199(.A(new_n2547_1), .B(new_n2507), .Y(new_n2548));
  nand_5 g00200(.A(new_n2548), .B(new_n2546), .Y(new_n2549));
  not_8  g00201(.A(new_n2549), .Y(new_n2550));
  nand_5 g00202(.A(new_n2452), .B(new_n2449), .Y(new_n2551));
  xor_4  g00203(.A(new_n2551), .B(new_n2453), .Y(new_n2552));
  not_8  g00204(.A(new_n2552), .Y(new_n2553_1));
  nor_5  g00205(.A(new_n2548), .B(new_n2546), .Y(new_n2554));
  nor_5  g00206(.A(new_n2554), .B(new_n2553_1), .Y(new_n2555_1));
  nor_5  g00207(.A(new_n2555_1), .B(new_n2550), .Y(new_n2556));
  not_8  g00208(.A(new_n2556), .Y(new_n2557));
  nand_5 g00209(.A(new_n2557), .B(new_n2542), .Y(new_n2558));
  nand_5 g00210(.A(new_n2558), .B(new_n2541), .Y(new_n2559));
  nand_5 g00211(.A(new_n2559), .B(new_n2536), .Y(new_n2560_1));
  nand_5 g00212(.A(new_n2560_1), .B(new_n2535_1), .Y(new_n2561_1));
  nand_5 g00213(.A(new_n2561_1), .B(new_n2530), .Y(new_n2562));
  nand_5 g00214(.A(new_n2562), .B(new_n2529), .Y(new_n2563));
  nor_5  g00215(.A(new_n2563), .B(new_n2524), .Y(new_n2564));
  nor_5  g00216(.A(new_n2564), .B(new_n2523), .Y(new_n2565));
  nand_5 g00217(.A(new_n2487), .B(new_n2462), .Y(new_n2566));
  nand_5 g00218(.A(new_n2566), .B(new_n2486), .Y(new_n2567));
  not_8  g00219(.A(n13783), .Y(new_n2568));
  not_8  g00220(.A(n22332), .Y(new_n2569));
  nand_5 g00221(.A(new_n2569), .B(new_n2568), .Y(new_n2570_1));
  nand_5 g00222(.A(n22332), .B(n13783), .Y(new_n2571));
  nand_5 g00223(.A(new_n2571), .B(new_n2570_1), .Y(new_n2572));
  nand_5 g00224(.A(new_n2479_1), .B(new_n2473), .Y(new_n2573_1));
  nand_5 g00225(.A(new_n2573_1), .B(new_n2476), .Y(new_n2574));
  xnor_4 g00226(.A(new_n2574), .B(new_n2572), .Y(new_n2575));
  not_8  g00227(.A(new_n2575), .Y(new_n2576));
  nor_5  g00228(.A(new_n2576), .B(new_n2482), .Y(new_n2577));
  not_8  g00229(.A(new_n2577), .Y(new_n2578_1));
  nand_5 g00230(.A(new_n2576), .B(new_n2482), .Y(new_n2579));
  and_5  g00231(.A(new_n2579), .B(new_n2578_1), .Y(new_n2580));
  nand_5 g00232(.A(new_n2466), .B(new_n2464), .Y(new_n2581));
  nand_5 g00233(.A(new_n2581), .B(new_n2469), .Y(new_n2582_1));
  not_8  g00234(.A(new_n2582_1), .Y(new_n2583));
  not_8  g00235(.A(n7751), .Y(new_n2584));
  not_8  g00236(.A(n13490), .Y(new_n2585));
  nand_5 g00237(.A(new_n2585), .B(new_n2584), .Y(new_n2586));
  nand_5 g00238(.A(n13490), .B(n7751), .Y(new_n2587));
  nand_5 g00239(.A(new_n2587), .B(new_n2586), .Y(new_n2588));
  xor_4  g00240(.A(new_n2588), .B(new_n2583), .Y(new_n2589));
  not_8  g00241(.A(new_n2589), .Y(new_n2590));
  nand_5 g00242(.A(new_n2590), .B(new_n2580), .Y(new_n2591));
  or_5   g00243(.A(new_n2590), .B(new_n2580), .Y(new_n2592));
  nand_5 g00244(.A(new_n2592), .B(new_n2591), .Y(new_n2593));
  xor_4  g00245(.A(new_n2593), .B(new_n2567), .Y(new_n2594));
  not_8  g00246(.A(new_n2594), .Y(new_n2595));
  nand_5 g00247(.A(new_n2519), .B(new_n2515_1), .Y(new_n2596));
  nand_5 g00248(.A(new_n2596), .B(new_n2517), .Y(new_n2597));
  not_8  g00249(.A(new_n2597), .Y(new_n2598));
  not_8  g00250(.A(n9942), .Y(new_n2599));
  nand_5 g00251(.A(n10739), .B(new_n2599), .Y(new_n2600));
  not_8  g00252(.A(n10739), .Y(new_n2601));
  nand_5 g00253(.A(new_n2601), .B(n9942), .Y(new_n2602_1));
  nand_5 g00254(.A(new_n2602_1), .B(new_n2600), .Y(new_n2603));
  xor_4  g00255(.A(new_n2603), .B(new_n2598), .Y(new_n2604));
  or_5   g00256(.A(new_n2604), .B(new_n2595), .Y(new_n2605));
  not_8  g00257(.A(new_n2605), .Y(new_n2606));
  nand_5 g00258(.A(new_n2604), .B(new_n2595), .Y(new_n2607));
  not_8  g00259(.A(new_n2607), .Y(new_n2608));
  nor_5  g00260(.A(new_n2608), .B(new_n2606), .Y(new_n2609));
  xor_4  g00261(.A(new_n2609), .B(new_n2565), .Y(n7));
  not_8  g00262(.A(n4588), .Y(new_n2611));
  nand_5 g00263(.A(n3618), .B(n1681), .Y(new_n2612));
  not_8  g00264(.A(n1681), .Y(new_n2613));
  not_8  g00265(.A(n3618), .Y(new_n2614));
  nand_5 g00266(.A(new_n2614), .B(new_n2613), .Y(new_n2615));
  and_5  g00267(.A(new_n2615), .B(new_n2612), .Y(new_n2616));
  xor_4  g00268(.A(new_n2616), .B(new_n2611), .Y(new_n2617));
  not_8  g00269(.A(new_n2617), .Y(new_n2618));
  not_8  g00270(.A(n22201), .Y(new_n2619_1));
  not_8  g00271(.A(n583), .Y(new_n2620));
  nand_5 g00272(.A(n22843), .B(new_n2620), .Y(new_n2621));
  not_8  g00273(.A(n22843), .Y(new_n2622));
  nand_5 g00274(.A(new_n2622), .B(n583), .Y(new_n2623));
  and_5  g00275(.A(new_n2623), .B(new_n2621), .Y(new_n2624));
  xor_4  g00276(.A(new_n2624), .B(new_n2619_1), .Y(new_n2625));
  nand_5 g00277(.A(new_n2625), .B(new_n2618), .Y(new_n2626));
  not_8  g00278(.A(new_n2626), .Y(new_n2627));
  nor_5  g00279(.A(new_n2625), .B(new_n2618), .Y(new_n2628));
  nor_5  g00280(.A(new_n2628), .B(new_n2627), .Y(n50));
  nand_5 g00281(.A(n21398), .B(n14090), .Y(new_n2630));
  not_8  g00282(.A(n14090), .Y(new_n2631));
  not_8  g00283(.A(n21398), .Y(new_n2632));
  nand_5 g00284(.A(new_n2632), .B(new_n2631), .Y(new_n2633));
  and_5  g00285(.A(new_n2633), .B(new_n2630), .Y(new_n2634));
  xor_4  g00286(.A(new_n2634), .B(n25926), .Y(new_n2635));
  not_8  g00287(.A(n21687), .Y(new_n2636));
  nand_5 g00288(.A(n19922), .B(n6773), .Y(new_n2637));
  not_8  g00289(.A(new_n2637), .Y(new_n2638));
  nor_5  g00290(.A(n19922), .B(n6773), .Y(new_n2639));
  or_5   g00291(.A(new_n2639), .B(new_n2638), .Y(new_n2640));
  xor_4  g00292(.A(new_n2640), .B(new_n2636), .Y(new_n2641));
  nand_5 g00293(.A(new_n2641), .B(new_n2635), .Y(new_n2642));
  not_8  g00294(.A(new_n2642), .Y(new_n2643));
  nor_5  g00295(.A(new_n2641), .B(new_n2635), .Y(new_n2644));
  nor_5  g00296(.A(new_n2644), .B(new_n2643), .Y(n55));
  nand_5 g00297(.A(n20040), .B(n9396), .Y(new_n2646_1));
  not_8  g00298(.A(n9396), .Y(new_n2647));
  not_8  g00299(.A(n20040), .Y(new_n2648));
  nand_5 g00300(.A(new_n2648), .B(new_n2647), .Y(new_n2649));
  nand_5 g00301(.A(new_n2649), .B(new_n2646_1), .Y(new_n2650));
  not_8  g00302(.A(n1999), .Y(new_n2651));
  not_8  g00303(.A(n19531), .Y(new_n2652));
  nand_5 g00304(.A(new_n2652), .B(new_n2651), .Y(new_n2653));
  nand_5 g00305(.A(n19531), .B(n1999), .Y(new_n2654));
  or_5   g00306(.A(n25168), .B(n18345), .Y(new_n2655));
  nand_5 g00307(.A(n25168), .B(n18345), .Y(new_n2656));
  not_8  g00308(.A(n9318), .Y(new_n2657));
  not_8  g00309(.A(n13190), .Y(new_n2658));
  nand_5 g00310(.A(new_n2658), .B(new_n2657), .Y(new_n2659_1));
  nand_5 g00311(.A(n13190), .B(n9318), .Y(new_n2660));
  or_5   g00312(.A(n19477), .B(n3460), .Y(new_n2661_1));
  nand_5 g00313(.A(n19477), .B(n3460), .Y(new_n2662));
  not_8  g00314(.A(n5226), .Y(new_n2663));
  not_8  g00315(.A(n11223), .Y(new_n2664));
  nand_5 g00316(.A(new_n2664), .B(new_n2663), .Y(new_n2665));
  nand_5 g00317(.A(n11223), .B(n5226), .Y(new_n2666));
  or_5   g00318(.A(n17664), .B(n5115), .Y(new_n2667));
  nand_5 g00319(.A(n17664), .B(n5115), .Y(new_n2668));
  not_8  g00320(.A(n23369), .Y(new_n2669));
  not_8  g00321(.A(n26572), .Y(new_n2670));
  nand_5 g00322(.A(new_n2670), .B(new_n2669), .Y(new_n2671));
  nand_5 g00323(.A(n26572), .B(n23369), .Y(new_n2672));
  not_8  g00324(.A(n1136), .Y(new_n2673));
  not_8  g00325(.A(n11667), .Y(new_n2674));
  nand_5 g00326(.A(new_n2674), .B(new_n2673), .Y(new_n2675));
  nand_5 g00327(.A(n11667), .B(n1136), .Y(new_n2676));
  nand_5 g00328(.A(n21398), .B(n19234), .Y(new_n2677));
  nand_5 g00329(.A(new_n2677), .B(new_n2676), .Y(new_n2678));
  nand_5 g00330(.A(new_n2678), .B(new_n2675), .Y(new_n2679));
  nand_5 g00331(.A(new_n2679), .B(new_n2672), .Y(new_n2680_1));
  nand_5 g00332(.A(new_n2680_1), .B(new_n2671), .Y(new_n2681));
  nand_5 g00333(.A(new_n2681), .B(new_n2668), .Y(new_n2682));
  nand_5 g00334(.A(new_n2682), .B(new_n2667), .Y(new_n2683));
  nand_5 g00335(.A(new_n2683), .B(new_n2666), .Y(new_n2684));
  nand_5 g00336(.A(new_n2684), .B(new_n2665), .Y(new_n2685));
  nand_5 g00337(.A(new_n2685), .B(new_n2662), .Y(new_n2686));
  nand_5 g00338(.A(new_n2686), .B(new_n2661_1), .Y(new_n2687));
  nand_5 g00339(.A(new_n2687), .B(new_n2660), .Y(new_n2688));
  nand_5 g00340(.A(new_n2688), .B(new_n2659_1), .Y(new_n2689));
  nand_5 g00341(.A(new_n2689), .B(new_n2656), .Y(new_n2690));
  nand_5 g00342(.A(new_n2690), .B(new_n2655), .Y(new_n2691));
  nand_5 g00343(.A(new_n2691), .B(new_n2654), .Y(new_n2692));
  nand_5 g00344(.A(new_n2692), .B(new_n2653), .Y(new_n2693_1));
  not_8  g00345(.A(new_n2693_1), .Y(new_n2694));
  xor_4  g00346(.A(new_n2694), .B(new_n2650), .Y(new_n2695));
  not_8  g00347(.A(new_n2695), .Y(new_n2696));
  nand_5 g00348(.A(new_n2696), .B(n25365), .Y(new_n2697));
  or_5   g00349(.A(new_n2696), .B(n25365), .Y(new_n2698));
  nand_5 g00350(.A(new_n2698), .B(new_n2697), .Y(new_n2699));
  nand_5 g00351(.A(new_n2654), .B(new_n2653), .Y(new_n2700));
  xor_4  g00352(.A(new_n2700), .B(new_n2691), .Y(new_n2701));
  nand_5 g00353(.A(new_n2701), .B(n14704), .Y(new_n2702));
  not_8  g00354(.A(n14704), .Y(new_n2703_1));
  not_8  g00355(.A(new_n2701), .Y(new_n2704));
  nand_5 g00356(.A(new_n2704), .B(new_n2703_1), .Y(new_n2705));
  nand_5 g00357(.A(new_n2656), .B(new_n2655), .Y(new_n2706_1));
  xor_4  g00358(.A(new_n2706_1), .B(new_n2689), .Y(new_n2707));
  nand_5 g00359(.A(new_n2707), .B(n19270), .Y(new_n2708));
  not_8  g00360(.A(n19270), .Y(new_n2709));
  not_8  g00361(.A(new_n2707), .Y(new_n2710));
  nand_5 g00362(.A(new_n2710), .B(new_n2709), .Y(new_n2711_1));
  nand_5 g00363(.A(new_n2660), .B(new_n2659_1), .Y(new_n2712));
  xor_4  g00364(.A(new_n2712), .B(new_n2687), .Y(new_n2713));
  nand_5 g00365(.A(new_n2713), .B(n8687), .Y(new_n2714));
  not_8  g00366(.A(n8687), .Y(new_n2715));
  not_8  g00367(.A(new_n2713), .Y(new_n2716));
  nand_5 g00368(.A(new_n2716), .B(new_n2715), .Y(new_n2717));
  nand_5 g00369(.A(new_n2662), .B(new_n2661_1), .Y(new_n2718));
  xor_4  g00370(.A(new_n2718), .B(new_n2685), .Y(new_n2719));
  nand_5 g00371(.A(new_n2719), .B(n24768), .Y(new_n2720));
  or_5   g00372(.A(new_n2719), .B(n24768), .Y(new_n2721));
  nand_5 g00373(.A(new_n2666), .B(new_n2665), .Y(new_n2722));
  xor_4  g00374(.A(new_n2722), .B(new_n2683), .Y(new_n2723));
  nand_5 g00375(.A(new_n2723), .B(n26483), .Y(new_n2724));
  not_8  g00376(.A(n26483), .Y(new_n2725));
  not_8  g00377(.A(new_n2723), .Y(new_n2726));
  nand_5 g00378(.A(new_n2726), .B(new_n2725), .Y(new_n2727));
  nand_5 g00379(.A(new_n2668), .B(new_n2667), .Y(new_n2728));
  xor_4  g00380(.A(new_n2728), .B(new_n2681), .Y(new_n2729));
  nand_5 g00381(.A(new_n2729), .B(n15979), .Y(new_n2730));
  or_5   g00382(.A(new_n2729), .B(n15979), .Y(new_n2731_1));
  nand_5 g00383(.A(new_n2672), .B(new_n2671), .Y(new_n2732));
  xor_4  g00384(.A(new_n2732), .B(new_n2679), .Y(new_n2733));
  nand_5 g00385(.A(new_n2733), .B(n8638), .Y(new_n2734));
  not_8  g00386(.A(n8638), .Y(new_n2735));
  not_8  g00387(.A(new_n2733), .Y(new_n2736));
  nand_5 g00388(.A(new_n2736), .B(new_n2735), .Y(new_n2737));
  nand_5 g00389(.A(new_n2676), .B(new_n2675), .Y(new_n2738));
  xor_4  g00390(.A(new_n2738), .B(new_n2677), .Y(new_n2739));
  nand_5 g00391(.A(new_n2739), .B(n16247), .Y(new_n2740));
  not_8  g00392(.A(n16247), .Y(new_n2741));
  not_8  g00393(.A(new_n2739), .Y(new_n2742));
  nand_5 g00394(.A(new_n2742), .B(new_n2741), .Y(new_n2743_1));
  not_8  g00395(.A(n19234), .Y(new_n2744));
  nand_5 g00396(.A(new_n2632), .B(new_n2744), .Y(new_n2745));
  and_5  g00397(.A(new_n2745), .B(new_n2677), .Y(new_n2746));
  nand_5 g00398(.A(new_n2746), .B(n23541), .Y(new_n2747));
  not_8  g00399(.A(new_n2747), .Y(new_n2748));
  nand_5 g00400(.A(new_n2748), .B(new_n2743_1), .Y(new_n2749));
  nand_5 g00401(.A(new_n2749), .B(new_n2740), .Y(new_n2750));
  nand_5 g00402(.A(new_n2750), .B(new_n2737), .Y(new_n2751));
  nand_5 g00403(.A(new_n2751), .B(new_n2734), .Y(new_n2752));
  nand_5 g00404(.A(new_n2752), .B(new_n2731_1), .Y(new_n2753));
  nand_5 g00405(.A(new_n2753), .B(new_n2730), .Y(new_n2754));
  nand_5 g00406(.A(new_n2754), .B(new_n2727), .Y(new_n2755));
  nand_5 g00407(.A(new_n2755), .B(new_n2724), .Y(new_n2756));
  nand_5 g00408(.A(new_n2756), .B(new_n2721), .Y(new_n2757));
  nand_5 g00409(.A(new_n2757), .B(new_n2720), .Y(new_n2758));
  nand_5 g00410(.A(new_n2758), .B(new_n2717), .Y(new_n2759));
  nand_5 g00411(.A(new_n2759), .B(new_n2714), .Y(new_n2760));
  nand_5 g00412(.A(new_n2760), .B(new_n2711_1), .Y(new_n2761_1));
  nand_5 g00413(.A(new_n2761_1), .B(new_n2708), .Y(new_n2762));
  nand_5 g00414(.A(new_n2762), .B(new_n2705), .Y(new_n2763));
  nand_5 g00415(.A(new_n2763), .B(new_n2702), .Y(new_n2764));
  xor_4  g00416(.A(new_n2764), .B(new_n2699), .Y(new_n2765));
  not_8  g00417(.A(n22793), .Y(new_n2766));
  not_8  g00418(.A(n25523), .Y(new_n2767));
  not_8  g00419(.A(n23430), .Y(new_n2768));
  not_8  g00420(.A(n11503), .Y(new_n2769));
  not_8  g00421(.A(n18151), .Y(new_n2770));
  nand_5 g00422(.A(new_n2770), .B(new_n2769), .Y(new_n2771));
  or_5   g00423(.A(new_n2771), .B(n16971), .Y(new_n2772));
  nor_5  g00424(.A(new_n2772), .B(n10411), .Y(new_n2773));
  nand_5 g00425(.A(new_n2773), .B(new_n2768), .Y(new_n2774_1));
  nor_5  g00426(.A(new_n2774_1), .B(n5579), .Y(new_n2775));
  nand_5 g00427(.A(new_n2775), .B(new_n2767), .Y(new_n2776));
  nor_5  g00428(.A(new_n2776), .B(n8439), .Y(new_n2777));
  nand_5 g00429(.A(new_n2777), .B(new_n2766), .Y(new_n2778));
  xor_4  g00430(.A(new_n2778), .B(n13951), .Y(new_n2779_1));
  nand_5 g00431(.A(n22270), .B(n2944), .Y(new_n2780));
  not_8  g00432(.A(n2944), .Y(new_n2781));
  not_8  g00433(.A(n22270), .Y(new_n2782));
  nand_5 g00434(.A(new_n2782), .B(new_n2781), .Y(new_n2783_1));
  nand_5 g00435(.A(new_n2783_1), .B(new_n2780), .Y(new_n2784));
  not_8  g00436(.A(n767), .Y(new_n2785));
  not_8  g00437(.A(n8806), .Y(new_n2786));
  nand_5 g00438(.A(new_n2786), .B(new_n2785), .Y(new_n2787));
  not_8  g00439(.A(new_n2787), .Y(new_n2788));
  nand_5 g00440(.A(n8806), .B(n767), .Y(new_n2789));
  not_8  g00441(.A(new_n2789), .Y(new_n2790));
  not_8  g00442(.A(n2479), .Y(new_n2791));
  not_8  g00443(.A(n7330), .Y(new_n2792));
  nand_5 g00444(.A(new_n2792), .B(new_n2791), .Y(new_n2793));
  not_8  g00445(.A(new_n2793), .Y(new_n2794));
  nand_5 g00446(.A(n7330), .B(n2479), .Y(new_n2795));
  not_8  g00447(.A(new_n2795), .Y(new_n2796));
  not_8  g00448(.A(n9372), .Y(new_n2797));
  not_8  g00449(.A(n22492), .Y(new_n2798));
  nand_5 g00450(.A(new_n2798), .B(new_n2797), .Y(new_n2799));
  not_8  g00451(.A(new_n2799), .Y(new_n2800));
  nand_5 g00452(.A(n22492), .B(n9372), .Y(new_n2801));
  not_8  g00453(.A(new_n2801), .Y(new_n2802));
  not_8  g00454(.A(n6596), .Y(new_n2803));
  not_8  g00455(.A(n6556), .Y(new_n2804));
  not_8  g00456(.A(n7149), .Y(new_n2805));
  not_8  g00457(.A(n22871), .Y(new_n2806));
  nand_5 g00458(.A(new_n2806), .B(new_n2805), .Y(new_n2807));
  nand_5 g00459(.A(n22871), .B(n7149), .Y(new_n2808));
  not_8  g00460(.A(n14148), .Y(new_n2809_1));
  not_8  g00461(.A(n14275), .Y(new_n2810));
  nand_5 g00462(.A(new_n2810), .B(new_n2809_1), .Y(new_n2811));
  nand_5 g00463(.A(n14275), .B(n14148), .Y(new_n2812));
  nand_5 g00464(.A(n25023), .B(n1152), .Y(new_n2813));
  nand_5 g00465(.A(new_n2813), .B(new_n2812), .Y(new_n2814));
  nand_5 g00466(.A(new_n2814), .B(new_n2811), .Y(new_n2815));
  nand_5 g00467(.A(new_n2815), .B(new_n2808), .Y(new_n2816_1));
  nand_5 g00468(.A(new_n2816_1), .B(new_n2807), .Y(new_n2817));
  nand_5 g00469(.A(new_n2817), .B(new_n2804), .Y(new_n2818));
  not_8  g00470(.A(new_n2818), .Y(new_n2819));
  nor_5  g00471(.A(new_n2817), .B(new_n2804), .Y(new_n2820));
  nor_5  g00472(.A(new_n2820), .B(n18558), .Y(new_n2821));
  nor_5  g00473(.A(new_n2821), .B(new_n2819), .Y(new_n2822));
  or_5   g00474(.A(new_n2822), .B(n3468), .Y(new_n2823));
  not_8  g00475(.A(n15289), .Y(new_n2824));
  nand_5 g00476(.A(new_n2822), .B(n3468), .Y(new_n2825));
  nand_5 g00477(.A(new_n2825), .B(new_n2824), .Y(new_n2826_1));
  nand_5 g00478(.A(new_n2826_1), .B(new_n2823), .Y(new_n2827));
  nand_5 g00479(.A(new_n2827), .B(new_n2803), .Y(new_n2828));
  not_8  g00480(.A(new_n2828), .Y(new_n2829));
  nor_5  g00481(.A(new_n2827), .B(new_n2803), .Y(new_n2830));
  nor_5  g00482(.A(new_n2830), .B(n12821), .Y(new_n2831));
  nor_5  g00483(.A(new_n2831), .B(new_n2829), .Y(new_n2832));
  nor_5  g00484(.A(new_n2832), .B(new_n2802), .Y(new_n2833));
  nor_5  g00485(.A(new_n2833), .B(new_n2800), .Y(new_n2834));
  nor_5  g00486(.A(new_n2834), .B(new_n2796), .Y(new_n2835));
  nor_5  g00487(.A(new_n2835), .B(new_n2794), .Y(new_n2836));
  nor_5  g00488(.A(new_n2836), .B(new_n2790), .Y(new_n2837));
  nor_5  g00489(.A(new_n2837), .B(new_n2788), .Y(new_n2838));
  not_8  g00490(.A(new_n2838), .Y(new_n2839));
  xor_4  g00491(.A(new_n2839), .B(new_n2784), .Y(new_n2840));
  not_8  g00492(.A(new_n2840), .Y(new_n2841));
  nand_5 g00493(.A(new_n2841), .B(new_n2779_1), .Y(new_n2842));
  not_8  g00494(.A(new_n2842), .Y(new_n2843));
  nor_5  g00495(.A(new_n2841), .B(new_n2779_1), .Y(new_n2844));
  nor_5  g00496(.A(new_n2844), .B(new_n2843), .Y(new_n2845));
  xor_4  g00497(.A(new_n2777), .B(new_n2766), .Y(new_n2846));
  nand_5 g00498(.A(new_n2789), .B(new_n2787), .Y(new_n2847));
  xor_4  g00499(.A(new_n2847), .B(new_n2836), .Y(new_n2848));
  or_5   g00500(.A(new_n2848), .B(new_n2846), .Y(new_n2849));
  nand_5 g00501(.A(new_n2848), .B(new_n2846), .Y(new_n2850));
  xor_4  g00502(.A(new_n2776), .B(n8439), .Y(new_n2851));
  nand_5 g00503(.A(new_n2795), .B(new_n2793), .Y(new_n2852));
  xor_4  g00504(.A(new_n2852), .B(new_n2834), .Y(new_n2853_1));
  or_5   g00505(.A(new_n2853_1), .B(new_n2851), .Y(new_n2854));
  nand_5 g00506(.A(new_n2853_1), .B(new_n2851), .Y(new_n2855));
  xor_4  g00507(.A(new_n2775), .B(new_n2767), .Y(new_n2856));
  nand_5 g00508(.A(new_n2801), .B(new_n2799), .Y(new_n2857));
  xor_4  g00509(.A(new_n2857), .B(new_n2832), .Y(new_n2858_1));
  or_5   g00510(.A(new_n2858_1), .B(new_n2856), .Y(new_n2859));
  nand_5 g00511(.A(new_n2858_1), .B(new_n2856), .Y(new_n2860_1));
  xor_4  g00512(.A(new_n2774_1), .B(n5579), .Y(new_n2861));
  not_8  g00513(.A(n12821), .Y(new_n2862));
  nor_5  g00514(.A(new_n2830), .B(new_n2829), .Y(new_n2863));
  xor_4  g00515(.A(new_n2863), .B(new_n2862), .Y(new_n2864));
  or_5   g00516(.A(new_n2864), .B(new_n2861), .Y(new_n2865));
  nand_5 g00517(.A(new_n2864), .B(new_n2861), .Y(new_n2866));
  xor_4  g00518(.A(new_n2773), .B(new_n2768), .Y(new_n2867));
  and_5  g00519(.A(new_n2825), .B(new_n2823), .Y(new_n2868));
  xor_4  g00520(.A(new_n2868), .B(new_n2824), .Y(new_n2869));
  or_5   g00521(.A(new_n2869), .B(new_n2867), .Y(new_n2870));
  nand_5 g00522(.A(new_n2869), .B(new_n2867), .Y(new_n2871));
  not_8  g00523(.A(n18558), .Y(new_n2872));
  nor_5  g00524(.A(new_n2820), .B(new_n2819), .Y(new_n2873));
  xor_4  g00525(.A(new_n2873), .B(new_n2872), .Y(new_n2874));
  not_8  g00526(.A(new_n2874), .Y(new_n2875));
  not_8  g00527(.A(n10411), .Y(new_n2876));
  xor_4  g00528(.A(new_n2772), .B(new_n2876), .Y(new_n2877));
  nand_5 g00529(.A(new_n2877), .B(new_n2875), .Y(new_n2878));
  or_5   g00530(.A(new_n2877), .B(new_n2875), .Y(new_n2879));
  nand_5 g00531(.A(new_n2771), .B(n16971), .Y(new_n2880));
  and_5  g00532(.A(new_n2880), .B(new_n2772), .Y(new_n2881));
  nand_5 g00533(.A(new_n2808), .B(new_n2807), .Y(new_n2882));
  xor_4  g00534(.A(new_n2882), .B(new_n2815), .Y(new_n2883));
  not_8  g00535(.A(new_n2883), .Y(new_n2884));
  or_5   g00536(.A(new_n2884), .B(new_n2881), .Y(new_n2885));
  nand_5 g00537(.A(new_n2884), .B(new_n2881), .Y(new_n2886_1));
  xor_4  g00538(.A(n18151), .B(n11503), .Y(new_n2887_1));
  nand_5 g00539(.A(new_n2812), .B(new_n2811), .Y(new_n2888));
  xor_4  g00540(.A(new_n2888), .B(new_n2813), .Y(new_n2889));
  not_8  g00541(.A(new_n2889), .Y(new_n2890));
  or_5   g00542(.A(new_n2890), .B(new_n2887_1), .Y(new_n2891));
  nand_5 g00543(.A(new_n2890), .B(new_n2887_1), .Y(new_n2892));
  xor_4  g00544(.A(n25023), .B(n1152), .Y(new_n2893));
  nand_5 g00545(.A(new_n2893), .B(new_n2770), .Y(new_n2894));
  not_8  g00546(.A(new_n2894), .Y(new_n2895));
  nand_5 g00547(.A(new_n2895), .B(new_n2892), .Y(new_n2896));
  nand_5 g00548(.A(new_n2896), .B(new_n2891), .Y(new_n2897));
  nand_5 g00549(.A(new_n2897), .B(new_n2886_1), .Y(new_n2898));
  nand_5 g00550(.A(new_n2898), .B(new_n2885), .Y(new_n2899));
  nand_5 g00551(.A(new_n2899), .B(new_n2879), .Y(new_n2900));
  nand_5 g00552(.A(new_n2900), .B(new_n2878), .Y(new_n2901));
  nand_5 g00553(.A(new_n2901), .B(new_n2871), .Y(new_n2902));
  nand_5 g00554(.A(new_n2902), .B(new_n2870), .Y(new_n2903));
  nand_5 g00555(.A(new_n2903), .B(new_n2866), .Y(new_n2904));
  nand_5 g00556(.A(new_n2904), .B(new_n2865), .Y(new_n2905));
  nand_5 g00557(.A(new_n2905), .B(new_n2860_1), .Y(new_n2906));
  nand_5 g00558(.A(new_n2906), .B(new_n2859), .Y(new_n2907));
  nand_5 g00559(.A(new_n2907), .B(new_n2855), .Y(new_n2908));
  nand_5 g00560(.A(new_n2908), .B(new_n2854), .Y(new_n2909));
  nand_5 g00561(.A(new_n2909), .B(new_n2850), .Y(new_n2910));
  nand_5 g00562(.A(new_n2910), .B(new_n2849), .Y(new_n2911));
  xor_4  g00563(.A(new_n2911), .B(new_n2845), .Y(new_n2912));
  or_5   g00564(.A(new_n2912), .B(new_n2765), .Y(new_n2913));
  nand_5 g00565(.A(new_n2912), .B(new_n2765), .Y(new_n2914));
  nand_5 g00566(.A(new_n2914), .B(new_n2913), .Y(new_n2915));
  nand_5 g00567(.A(new_n2702), .B(new_n2705), .Y(new_n2916));
  xor_4  g00568(.A(new_n2916), .B(new_n2762), .Y(new_n2917));
  not_8  g00569(.A(new_n2917), .Y(new_n2918));
  nand_5 g00570(.A(new_n2850), .B(new_n2849), .Y(new_n2919));
  xor_4  g00571(.A(new_n2919), .B(new_n2909), .Y(new_n2920));
  nand_5 g00572(.A(new_n2920), .B(new_n2918), .Y(new_n2921));
  or_5   g00573(.A(new_n2920), .B(new_n2918), .Y(new_n2922));
  nand_5 g00574(.A(new_n2708), .B(new_n2711_1), .Y(new_n2923));
  xor_4  g00575(.A(new_n2923), .B(new_n2760), .Y(new_n2924));
  not_8  g00576(.A(new_n2924), .Y(new_n2925));
  nand_5 g00577(.A(new_n2855), .B(new_n2854), .Y(new_n2926));
  xor_4  g00578(.A(new_n2926), .B(new_n2907), .Y(new_n2927));
  nand_5 g00579(.A(new_n2927), .B(new_n2925), .Y(new_n2928));
  or_5   g00580(.A(new_n2927), .B(new_n2925), .Y(new_n2929_1));
  nand_5 g00581(.A(new_n2714), .B(new_n2717), .Y(new_n2930));
  xor_4  g00582(.A(new_n2930), .B(new_n2758), .Y(new_n2931));
  not_8  g00583(.A(new_n2931), .Y(new_n2932));
  nand_5 g00584(.A(new_n2860_1), .B(new_n2859), .Y(new_n2933));
  xor_4  g00585(.A(new_n2933), .B(new_n2905), .Y(new_n2934));
  nand_5 g00586(.A(new_n2934), .B(new_n2932), .Y(new_n2935));
  or_5   g00587(.A(new_n2934), .B(new_n2932), .Y(new_n2936));
  nand_5 g00588(.A(new_n2720), .B(new_n2721), .Y(new_n2937));
  xor_4  g00589(.A(new_n2937), .B(new_n2756), .Y(new_n2938));
  not_8  g00590(.A(new_n2938), .Y(new_n2939));
  nand_5 g00591(.A(new_n2866), .B(new_n2865), .Y(new_n2940));
  xor_4  g00592(.A(new_n2940), .B(new_n2903), .Y(new_n2941));
  nand_5 g00593(.A(new_n2941), .B(new_n2939), .Y(new_n2942));
  or_5   g00594(.A(new_n2941), .B(new_n2939), .Y(new_n2943));
  nand_5 g00595(.A(new_n2724), .B(new_n2727), .Y(new_n2944_1));
  xor_4  g00596(.A(new_n2944_1), .B(new_n2754), .Y(new_n2945));
  not_8  g00597(.A(new_n2945), .Y(new_n2946));
  nand_5 g00598(.A(new_n2871), .B(new_n2870), .Y(new_n2947));
  xor_4  g00599(.A(new_n2947), .B(new_n2901), .Y(new_n2948_1));
  nand_5 g00600(.A(new_n2948_1), .B(new_n2946), .Y(new_n2949));
  or_5   g00601(.A(new_n2948_1), .B(new_n2946), .Y(new_n2950));
  nand_5 g00602(.A(new_n2730), .B(new_n2731_1), .Y(new_n2951));
  xor_4  g00603(.A(new_n2951), .B(new_n2752), .Y(new_n2952));
  not_8  g00604(.A(new_n2952), .Y(new_n2953));
  nand_5 g00605(.A(new_n2879), .B(new_n2878), .Y(new_n2954));
  xor_4  g00606(.A(new_n2954), .B(new_n2899), .Y(new_n2955));
  nand_5 g00607(.A(new_n2955), .B(new_n2953), .Y(new_n2956));
  or_5   g00608(.A(new_n2955), .B(new_n2953), .Y(new_n2957));
  nand_5 g00609(.A(new_n2734), .B(new_n2737), .Y(new_n2958));
  xor_4  g00610(.A(new_n2958), .B(new_n2750), .Y(new_n2959));
  not_8  g00611(.A(new_n2959), .Y(new_n2960));
  nand_5 g00612(.A(new_n2886_1), .B(new_n2885), .Y(new_n2961_1));
  xor_4  g00613(.A(new_n2961_1), .B(new_n2897), .Y(new_n2962));
  nand_5 g00614(.A(new_n2962), .B(new_n2960), .Y(new_n2963));
  or_5   g00615(.A(new_n2962), .B(new_n2960), .Y(new_n2964));
  nand_5 g00616(.A(new_n2892), .B(new_n2891), .Y(new_n2965));
  xor_4  g00617(.A(new_n2965), .B(new_n2895), .Y(new_n2966));
  nand_5 g00618(.A(new_n2740), .B(new_n2743_1), .Y(new_n2967));
  xor_4  g00619(.A(new_n2967), .B(new_n2748), .Y(new_n2968));
  not_8  g00620(.A(new_n2968), .Y(new_n2969));
  nand_5 g00621(.A(new_n2969), .B(new_n2966), .Y(new_n2970));
  not_8  g00622(.A(new_n2967), .Y(new_n2971_1));
  nor_5  g00623(.A(new_n2971_1), .B(new_n2966), .Y(new_n2972));
  not_8  g00624(.A(n23541), .Y(new_n2973));
  not_8  g00625(.A(new_n2746), .Y(new_n2974));
  nand_5 g00626(.A(new_n2974), .B(new_n2973), .Y(new_n2975));
  and_5  g00627(.A(new_n2975), .B(new_n2747), .Y(new_n2976));
  xor_4  g00628(.A(new_n2893), .B(n18151), .Y(new_n2977));
  nand_5 g00629(.A(new_n2977), .B(new_n2976), .Y(new_n2978_1));
  or_5   g00630(.A(new_n2978_1), .B(new_n2972), .Y(new_n2979_1));
  nand_5 g00631(.A(new_n2979_1), .B(new_n2970), .Y(new_n2980));
  nand_5 g00632(.A(new_n2980), .B(new_n2964), .Y(new_n2981));
  nand_5 g00633(.A(new_n2981), .B(new_n2963), .Y(new_n2982));
  nand_5 g00634(.A(new_n2982), .B(new_n2957), .Y(new_n2983));
  nand_5 g00635(.A(new_n2983), .B(new_n2956), .Y(new_n2984));
  nand_5 g00636(.A(new_n2984), .B(new_n2950), .Y(new_n2985_1));
  nand_5 g00637(.A(new_n2985_1), .B(new_n2949), .Y(new_n2986));
  nand_5 g00638(.A(new_n2986), .B(new_n2943), .Y(new_n2987));
  nand_5 g00639(.A(new_n2987), .B(new_n2942), .Y(new_n2988));
  nand_5 g00640(.A(new_n2988), .B(new_n2936), .Y(new_n2989));
  nand_5 g00641(.A(new_n2989), .B(new_n2935), .Y(new_n2990));
  nand_5 g00642(.A(new_n2990), .B(new_n2929_1), .Y(new_n2991));
  nand_5 g00643(.A(new_n2991), .B(new_n2928), .Y(new_n2992));
  nand_5 g00644(.A(new_n2992), .B(new_n2922), .Y(new_n2993));
  nand_5 g00645(.A(new_n2993), .B(new_n2921), .Y(new_n2994));
  xnor_4 g00646(.A(new_n2994), .B(new_n2915), .Y(n108));
  nand_5 g00647(.A(new_n2798), .B(n12875), .Y(new_n2996));
  not_8  g00648(.A(n12875), .Y(new_n2997));
  nand_5 g00649(.A(n22492), .B(new_n2997), .Y(new_n2998));
  nand_5 g00650(.A(new_n2862), .B(n2035), .Y(new_n2999_1));
  not_8  g00651(.A(n2035), .Y(new_n3000));
  nand_5 g00652(.A(n12821), .B(new_n3000), .Y(new_n3001));
  not_8  g00653(.A(n3468), .Y(new_n3002));
  nand_5 g00654(.A(n5213), .B(new_n3002), .Y(new_n3003));
  not_8  g00655(.A(n5213), .Y(new_n3004));
  nand_5 g00656(.A(new_n3004), .B(n3468), .Y(new_n3005));
  nand_5 g00657(.A(new_n2872), .B(n4665), .Y(new_n3006));
  not_8  g00658(.A(n4665), .Y(new_n3007));
  nand_5 g00659(.A(n18558), .B(new_n3007), .Y(new_n3008));
  nand_5 g00660(.A(n19005), .B(new_n2805), .Y(new_n3009));
  not_8  g00661(.A(n19005), .Y(new_n3010_1));
  nand_5 g00662(.A(new_n3010_1), .B(n7149), .Y(new_n3011));
  nand_5 g00663(.A(new_n2809_1), .B(n4326), .Y(new_n3012));
  not_8  g00664(.A(n4326), .Y(new_n3013));
  nand_5 g00665(.A(n14148), .B(new_n3013), .Y(new_n3014));
  not_8  g00666(.A(n5438), .Y(new_n3015));
  nand_5 g00667(.A(new_n3015), .B(n1152), .Y(new_n3016));
  nand_5 g00668(.A(new_n3016), .B(new_n3014), .Y(new_n3017_1));
  nand_5 g00669(.A(new_n3017_1), .B(new_n3012), .Y(new_n3018_1));
  nand_5 g00670(.A(new_n3018_1), .B(new_n3011), .Y(new_n3019));
  nand_5 g00671(.A(new_n3019), .B(new_n3009), .Y(new_n3020_1));
  nand_5 g00672(.A(new_n3020_1), .B(new_n3008), .Y(new_n3021));
  nand_5 g00673(.A(new_n3021), .B(new_n3006), .Y(new_n3022));
  nand_5 g00674(.A(new_n3022), .B(new_n3005), .Y(new_n3023));
  nand_5 g00675(.A(new_n3023), .B(new_n3003), .Y(new_n3024));
  nand_5 g00676(.A(new_n3024), .B(new_n3001), .Y(new_n3025));
  nand_5 g00677(.A(new_n3025), .B(new_n2999_1), .Y(new_n3026));
  nand_5 g00678(.A(new_n3026), .B(new_n2998), .Y(new_n3027));
  nand_5 g00679(.A(new_n3027), .B(new_n2996), .Y(new_n3028));
  nand_5 g00680(.A(new_n2792), .B(n1662), .Y(new_n3029));
  not_8  g00681(.A(n1662), .Y(new_n3030_1));
  nand_5 g00682(.A(n7330), .B(new_n3030_1), .Y(new_n3031));
  nand_5 g00683(.A(new_n3031), .B(new_n3029), .Y(new_n3032));
  xor_4  g00684(.A(new_n3032), .B(new_n3028), .Y(new_n3033));
  not_8  g00685(.A(n7099), .Y(new_n3034));
  not_8  g00686(.A(n24620), .Y(new_n3035));
  nand_5 g00687(.A(new_n3035), .B(new_n3034), .Y(new_n3036));
  nand_5 g00688(.A(n24620), .B(n7099), .Y(new_n3037));
  not_8  g00689(.A(n5211), .Y(new_n3038));
  not_8  g00690(.A(n12811), .Y(new_n3039));
  nand_5 g00691(.A(new_n3039), .B(new_n3038), .Y(new_n3040));
  nand_5 g00692(.A(n12811), .B(n5211), .Y(new_n3041));
  not_8  g00693(.A(n1118), .Y(new_n3042));
  not_8  g00694(.A(n12956), .Y(new_n3043));
  nand_5 g00695(.A(new_n3043), .B(new_n3042), .Y(new_n3044));
  nand_5 g00696(.A(n12956), .B(n1118), .Y(new_n3045));
  not_8  g00697(.A(n18295), .Y(new_n3046));
  not_8  g00698(.A(n25974), .Y(new_n3047));
  nand_5 g00699(.A(new_n3047), .B(new_n3046), .Y(new_n3048));
  nand_5 g00700(.A(n25974), .B(n18295), .Y(new_n3049));
  not_8  g00701(.A(n1630), .Y(new_n3050));
  not_8  g00702(.A(n6502), .Y(new_n3051));
  nand_5 g00703(.A(new_n3051), .B(new_n3050), .Y(new_n3052));
  nand_5 g00704(.A(n6502), .B(n1630), .Y(new_n3053));
  nand_5 g00705(.A(n15780), .B(n1451), .Y(new_n3054));
  nand_5 g00706(.A(new_n3054), .B(new_n3053), .Y(new_n3055));
  nand_5 g00707(.A(new_n3055), .B(new_n3052), .Y(new_n3056));
  nand_5 g00708(.A(new_n3056), .B(new_n3049), .Y(new_n3057));
  nand_5 g00709(.A(new_n3057), .B(new_n3048), .Y(new_n3058));
  nand_5 g00710(.A(new_n3058), .B(new_n3045), .Y(new_n3059));
  nand_5 g00711(.A(new_n3059), .B(new_n3044), .Y(new_n3060));
  nand_5 g00712(.A(new_n3060), .B(new_n3041), .Y(new_n3061));
  nand_5 g00713(.A(new_n3061), .B(new_n3040), .Y(new_n3062));
  nand_5 g00714(.A(new_n3062), .B(new_n3037), .Y(new_n3063));
  nand_5 g00715(.A(new_n3063), .B(new_n3036), .Y(new_n3064));
  not_8  g00716(.A(new_n3064), .Y(new_n3065));
  nand_5 g00717(.A(n23529), .B(n20700), .Y(new_n3066));
  not_8  g00718(.A(n20700), .Y(new_n3067_1));
  not_8  g00719(.A(n23529), .Y(new_n3068));
  nand_5 g00720(.A(new_n3068), .B(new_n3067_1), .Y(new_n3069));
  nand_5 g00721(.A(new_n3069), .B(new_n3066), .Y(new_n3070));
  xor_4  g00722(.A(new_n3070), .B(new_n3065), .Y(new_n3071));
  not_8  g00723(.A(n20929), .Y(new_n3072));
  not_8  g00724(.A(n23068), .Y(new_n3073));
  nand_5 g00725(.A(new_n3073), .B(new_n3072), .Y(new_n3074));
  not_8  g00726(.A(new_n3074), .Y(new_n3075));
  nand_5 g00727(.A(n23068), .B(n20929), .Y(new_n3076_1));
  not_8  g00728(.A(new_n3076_1), .Y(new_n3077));
  not_8  g00729(.A(n8006), .Y(new_n3078));
  not_8  g00730(.A(n19514), .Y(new_n3079));
  nand_5 g00731(.A(new_n3079), .B(new_n3078), .Y(new_n3080));
  not_8  g00732(.A(new_n3080), .Y(new_n3081));
  nand_5 g00733(.A(n19514), .B(n8006), .Y(new_n3082));
  not_8  g00734(.A(new_n3082), .Y(new_n3083));
  not_8  g00735(.A(n10053), .Y(new_n3084));
  not_8  g00736(.A(n8399), .Y(new_n3085));
  not_8  g00737(.A(n16396), .Y(new_n3086));
  nand_5 g00738(.A(new_n3086), .B(new_n3085), .Y(new_n3087));
  nand_5 g00739(.A(n16396), .B(n8399), .Y(new_n3088));
  not_8  g00740(.A(n9399), .Y(new_n3089_1));
  not_8  g00741(.A(n9507), .Y(new_n3090));
  nand_5 g00742(.A(new_n3090), .B(new_n3089_1), .Y(new_n3091));
  nand_5 g00743(.A(n9507), .B(n9399), .Y(new_n3092));
  nand_5 g00744(.A(n26979), .B(n2088), .Y(new_n3093));
  nand_5 g00745(.A(new_n3093), .B(new_n3092), .Y(new_n3094));
  nand_5 g00746(.A(new_n3094), .B(new_n3091), .Y(new_n3095));
  nand_5 g00747(.A(new_n3095), .B(new_n3088), .Y(new_n3096));
  nand_5 g00748(.A(new_n3096), .B(new_n3087), .Y(new_n3097));
  nand_5 g00749(.A(new_n3097), .B(new_n3084), .Y(new_n3098));
  not_8  g00750(.A(new_n3098), .Y(new_n3099));
  nor_5  g00751(.A(new_n3097), .B(new_n3084), .Y(new_n3100));
  nor_5  g00752(.A(new_n3100), .B(n25074), .Y(new_n3101));
  nor_5  g00753(.A(new_n3101), .B(new_n3099), .Y(new_n3102));
  nor_5  g00754(.A(new_n3102), .B(new_n3083), .Y(new_n3103));
  nor_5  g00755(.A(new_n3103), .B(new_n3081), .Y(new_n3104));
  nor_5  g00756(.A(new_n3104), .B(new_n3077), .Y(new_n3105));
  nor_5  g00757(.A(new_n3105), .B(new_n3075), .Y(new_n3106));
  nand_5 g00758(.A(n26510), .B(n10710), .Y(new_n3107));
  not_8  g00759(.A(n10710), .Y(new_n3108));
  not_8  g00760(.A(n26510), .Y(new_n3109));
  nand_5 g00761(.A(new_n3109), .B(new_n3108), .Y(new_n3110));
  nand_5 g00762(.A(new_n3110), .B(new_n3107), .Y(new_n3111));
  xor_4  g00763(.A(new_n3111), .B(new_n3106), .Y(new_n3112));
  not_8  g00764(.A(new_n3112), .Y(new_n3113));
  nand_5 g00765(.A(new_n3113), .B(new_n3071), .Y(new_n3114));
  not_8  g00766(.A(new_n3071), .Y(new_n3115));
  nand_5 g00767(.A(new_n3112), .B(new_n3115), .Y(new_n3116));
  nand_5 g00768(.A(new_n3037), .B(new_n3036), .Y(new_n3117));
  xor_4  g00769(.A(new_n3117), .B(new_n3062), .Y(new_n3118));
  not_8  g00770(.A(new_n3118), .Y(new_n3119));
  nand_5 g00771(.A(new_n3076_1), .B(new_n3074), .Y(new_n3120));
  xor_4  g00772(.A(new_n3120), .B(new_n3104), .Y(new_n3121));
  not_8  g00773(.A(new_n3121), .Y(new_n3122));
  nand_5 g00774(.A(new_n3122), .B(new_n3119), .Y(new_n3123));
  nand_5 g00775(.A(new_n3121), .B(new_n3118), .Y(new_n3124));
  nand_5 g00776(.A(new_n3041), .B(new_n3040), .Y(new_n3125_1));
  xor_4  g00777(.A(new_n3125_1), .B(new_n3060), .Y(new_n3126_1));
  not_8  g00778(.A(new_n3126_1), .Y(new_n3127));
  nand_5 g00779(.A(new_n3082), .B(new_n3080), .Y(new_n3128));
  xor_4  g00780(.A(new_n3128), .B(new_n3102), .Y(new_n3129));
  not_8  g00781(.A(new_n3129), .Y(new_n3130));
  nand_5 g00782(.A(new_n3130), .B(new_n3127), .Y(new_n3131));
  nand_5 g00783(.A(new_n3129), .B(new_n3126_1), .Y(new_n3132));
  nand_5 g00784(.A(new_n3045), .B(new_n3044), .Y(new_n3133));
  xor_4  g00785(.A(new_n3133), .B(new_n3058), .Y(new_n3134));
  not_8  g00786(.A(new_n3134), .Y(new_n3135));
  not_8  g00787(.A(n25074), .Y(new_n3136_1));
  nor_5  g00788(.A(new_n3100), .B(new_n3099), .Y(new_n3137));
  xor_4  g00789(.A(new_n3137), .B(new_n3136_1), .Y(new_n3138));
  not_8  g00790(.A(new_n3138), .Y(new_n3139));
  nand_5 g00791(.A(new_n3139), .B(new_n3135), .Y(new_n3140));
  nand_5 g00792(.A(new_n3138), .B(new_n3134), .Y(new_n3141));
  nand_5 g00793(.A(new_n3049), .B(new_n3048), .Y(new_n3142));
  xor_4  g00794(.A(new_n3142), .B(new_n3056), .Y(new_n3143));
  not_8  g00795(.A(new_n3143), .Y(new_n3144));
  nand_5 g00796(.A(new_n3088), .B(new_n3087), .Y(new_n3145));
  xor_4  g00797(.A(new_n3145), .B(new_n3095), .Y(new_n3146));
  nand_5 g00798(.A(new_n3146), .B(new_n3144), .Y(new_n3147));
  not_8  g00799(.A(new_n3146), .Y(new_n3148));
  nand_5 g00800(.A(new_n3148), .B(new_n3143), .Y(new_n3149));
  nand_5 g00801(.A(new_n3053), .B(new_n3052), .Y(new_n3150));
  xor_4  g00802(.A(new_n3150), .B(new_n3054), .Y(new_n3151));
  not_8  g00803(.A(new_n3151), .Y(new_n3152));
  nand_5 g00804(.A(new_n3092), .B(new_n3091), .Y(new_n3153));
  xor_4  g00805(.A(new_n3153), .B(new_n3093), .Y(new_n3154));
  nand_5 g00806(.A(new_n3154), .B(new_n3152), .Y(new_n3155));
  not_8  g00807(.A(new_n3154), .Y(new_n3156));
  nand_5 g00808(.A(new_n3156), .B(new_n3151), .Y(new_n3157));
  not_8  g00809(.A(n1451), .Y(new_n3158));
  not_8  g00810(.A(n15780), .Y(new_n3159));
  nand_5 g00811(.A(new_n3159), .B(new_n3158), .Y(new_n3160));
  and_5  g00812(.A(new_n3160), .B(new_n3054), .Y(new_n3161_1));
  not_8  g00813(.A(new_n3161_1), .Y(new_n3162));
  not_8  g00814(.A(n2088), .Y(new_n3163));
  not_8  g00815(.A(n26979), .Y(new_n3164_1));
  nand_5 g00816(.A(new_n3164_1), .B(new_n3163), .Y(new_n3165));
  and_5  g00817(.A(new_n3165), .B(new_n3093), .Y(new_n3166));
  nand_5 g00818(.A(new_n3166), .B(new_n3162), .Y(new_n3167));
  not_8  g00819(.A(new_n3167), .Y(new_n3168));
  nand_5 g00820(.A(new_n3168), .B(new_n3157), .Y(new_n3169));
  nand_5 g00821(.A(new_n3169), .B(new_n3155), .Y(new_n3170));
  nand_5 g00822(.A(new_n3170), .B(new_n3149), .Y(new_n3171));
  nand_5 g00823(.A(new_n3171), .B(new_n3147), .Y(new_n3172));
  nand_5 g00824(.A(new_n3172), .B(new_n3141), .Y(new_n3173));
  nand_5 g00825(.A(new_n3173), .B(new_n3140), .Y(new_n3174));
  nand_5 g00826(.A(new_n3174), .B(new_n3132), .Y(new_n3175));
  nand_5 g00827(.A(new_n3175), .B(new_n3131), .Y(new_n3176));
  nand_5 g00828(.A(new_n3176), .B(new_n3124), .Y(new_n3177));
  nand_5 g00829(.A(new_n3177), .B(new_n3123), .Y(new_n3178));
  nand_5 g00830(.A(new_n3178), .B(new_n3116), .Y(new_n3179));
  nand_5 g00831(.A(new_n3179), .B(new_n3114), .Y(new_n3180));
  nand_5 g00832(.A(new_n3066), .B(new_n3064), .Y(new_n3181));
  nand_5 g00833(.A(new_n3181), .B(new_n3069), .Y(new_n3182));
  not_8  g00834(.A(new_n3182), .Y(new_n3183));
  nand_5 g00835(.A(n19701), .B(n7437), .Y(new_n3184));
  not_8  g00836(.A(n7437), .Y(new_n3185));
  not_8  g00837(.A(n19701), .Y(new_n3186));
  nand_5 g00838(.A(new_n3186), .B(new_n3185), .Y(new_n3187));
  nand_5 g00839(.A(new_n3187), .B(new_n3184), .Y(new_n3188));
  xor_4  g00840(.A(new_n3188), .B(new_n3183), .Y(new_n3189));
  not_8  g00841(.A(new_n3110), .Y(new_n3190));
  not_8  g00842(.A(new_n3107), .Y(new_n3191));
  nor_5  g00843(.A(new_n3191), .B(new_n3106), .Y(new_n3192));
  nor_5  g00844(.A(new_n3192), .B(new_n3190), .Y(new_n3193));
  not_8  g00845(.A(n11841), .Y(new_n3194));
  not_8  g00846(.A(n17077), .Y(new_n3195));
  nand_5 g00847(.A(new_n3195), .B(new_n3194), .Y(new_n3196));
  nand_5 g00848(.A(n17077), .B(n11841), .Y(new_n3197));
  nand_5 g00849(.A(new_n3197), .B(new_n3196), .Y(new_n3198));
  xor_4  g00850(.A(new_n3198), .B(new_n3193), .Y(new_n3199));
  not_8  g00851(.A(new_n3199), .Y(new_n3200));
  nand_5 g00852(.A(new_n3200), .B(new_n3189), .Y(new_n3201));
  not_8  g00853(.A(new_n3189), .Y(new_n3202));
  nand_5 g00854(.A(new_n3199), .B(new_n3202), .Y(new_n3203));
  nand_5 g00855(.A(new_n3203), .B(new_n3201), .Y(new_n3204));
  xor_4  g00856(.A(new_n3204), .B(new_n3180), .Y(new_n3205));
  not_8  g00857(.A(new_n3205), .Y(new_n3206));
  or_5   g00858(.A(new_n3206), .B(new_n3033), .Y(new_n3207));
  nand_5 g00859(.A(new_n3206), .B(new_n3033), .Y(new_n3208_1));
  nand_5 g00860(.A(new_n2998), .B(new_n2996), .Y(new_n3209));
  xor_4  g00861(.A(new_n3209), .B(new_n3026), .Y(new_n3210));
  nand_5 g00862(.A(new_n3114), .B(new_n3116), .Y(new_n3211));
  xor_4  g00863(.A(new_n3211), .B(new_n3178), .Y(new_n3212));
  not_8  g00864(.A(new_n3212), .Y(new_n3213));
  or_5   g00865(.A(new_n3213), .B(new_n3210), .Y(new_n3214));
  nand_5 g00866(.A(new_n3213), .B(new_n3210), .Y(new_n3215));
  nand_5 g00867(.A(new_n3001), .B(new_n2999_1), .Y(new_n3216));
  xor_4  g00868(.A(new_n3216), .B(new_n3024), .Y(new_n3217));
  nand_5 g00869(.A(new_n3123), .B(new_n3124), .Y(new_n3218));
  xor_4  g00870(.A(new_n3218), .B(new_n3176), .Y(new_n3219_1));
  not_8  g00871(.A(new_n3219_1), .Y(new_n3220));
  or_5   g00872(.A(new_n3220), .B(new_n3217), .Y(new_n3221));
  nand_5 g00873(.A(new_n3220), .B(new_n3217), .Y(new_n3222));
  nand_5 g00874(.A(new_n3005), .B(new_n3003), .Y(new_n3223));
  xor_4  g00875(.A(new_n3223), .B(new_n3022), .Y(new_n3224));
  nand_5 g00876(.A(new_n3131), .B(new_n3132), .Y(new_n3225));
  xor_4  g00877(.A(new_n3225), .B(new_n3174), .Y(new_n3226));
  not_8  g00878(.A(new_n3226), .Y(new_n3227));
  or_5   g00879(.A(new_n3227), .B(new_n3224), .Y(new_n3228_1));
  nand_5 g00880(.A(new_n3227), .B(new_n3224), .Y(new_n3229));
  nand_5 g00881(.A(new_n3008), .B(new_n3006), .Y(new_n3230));
  xor_4  g00882(.A(new_n3230), .B(new_n3020_1), .Y(new_n3231));
  nand_5 g00883(.A(new_n3140), .B(new_n3141), .Y(new_n3232));
  xor_4  g00884(.A(new_n3232), .B(new_n3172), .Y(new_n3233));
  not_8  g00885(.A(new_n3233), .Y(new_n3234));
  or_5   g00886(.A(new_n3234), .B(new_n3231), .Y(new_n3235_1));
  nand_5 g00887(.A(new_n3234), .B(new_n3231), .Y(new_n3236));
  nand_5 g00888(.A(new_n3011), .B(new_n3009), .Y(new_n3237));
  xor_4  g00889(.A(new_n3237), .B(new_n3018_1), .Y(new_n3238));
  nand_5 g00890(.A(new_n3147), .B(new_n3149), .Y(new_n3239));
  xor_4  g00891(.A(new_n3239), .B(new_n3170), .Y(new_n3240));
  not_8  g00892(.A(new_n3240), .Y(new_n3241));
  or_5   g00893(.A(new_n3241), .B(new_n3238), .Y(new_n3242));
  nand_5 g00894(.A(new_n3241), .B(new_n3238), .Y(new_n3243));
  not_8  g00895(.A(new_n3166), .Y(new_n3244_1));
  nand_5 g00896(.A(new_n3244_1), .B(new_n3161_1), .Y(new_n3245));
  and_5  g00897(.A(new_n3245), .B(new_n3167), .Y(new_n3246));
  not_8  g00898(.A(new_n3246), .Y(new_n3247));
  not_8  g00899(.A(n1152), .Y(new_n3248));
  nand_5 g00900(.A(n5438), .B(new_n3248), .Y(new_n3249));
  nand_5 g00901(.A(new_n3249), .B(new_n3016), .Y(new_n3250));
  nand_5 g00902(.A(new_n3250), .B(new_n3247), .Y(new_n3251));
  not_8  g00903(.A(new_n3016), .Y(new_n3252));
  and_5  g00904(.A(new_n3014), .B(new_n3012), .Y(new_n3253_1));
  xor_4  g00905(.A(new_n3253_1), .B(new_n3252), .Y(new_n3254));
  or_5   g00906(.A(new_n3254), .B(new_n3251), .Y(new_n3255));
  nand_5 g00907(.A(new_n3254), .B(new_n3251), .Y(new_n3256));
  nand_5 g00908(.A(new_n3155), .B(new_n3157), .Y(new_n3257));
  xor_4  g00909(.A(new_n3257), .B(new_n3168), .Y(new_n3258));
  nand_5 g00910(.A(new_n3258), .B(new_n3256), .Y(new_n3259));
  nand_5 g00911(.A(new_n3259), .B(new_n3255), .Y(new_n3260_1));
  nand_5 g00912(.A(new_n3260_1), .B(new_n3243), .Y(new_n3261));
  nand_5 g00913(.A(new_n3261), .B(new_n3242), .Y(new_n3262));
  nand_5 g00914(.A(new_n3262), .B(new_n3236), .Y(new_n3263_1));
  nand_5 g00915(.A(new_n3263_1), .B(new_n3235_1), .Y(new_n3264));
  nand_5 g00916(.A(new_n3264), .B(new_n3229), .Y(new_n3265));
  nand_5 g00917(.A(new_n3265), .B(new_n3228_1), .Y(new_n3266));
  nand_5 g00918(.A(new_n3266), .B(new_n3222), .Y(new_n3267));
  nand_5 g00919(.A(new_n3267), .B(new_n3221), .Y(new_n3268));
  nand_5 g00920(.A(new_n3268), .B(new_n3215), .Y(new_n3269));
  nand_5 g00921(.A(new_n3269), .B(new_n3214), .Y(new_n3270));
  nand_5 g00922(.A(new_n3270), .B(new_n3208_1), .Y(new_n3271));
  nand_5 g00923(.A(new_n3271), .B(new_n3207), .Y(new_n3272));
  nand_5 g00924(.A(new_n3031), .B(new_n3028), .Y(new_n3273));
  nand_5 g00925(.A(new_n3273), .B(new_n3029), .Y(new_n3274));
  nand_5 g00926(.A(n22379), .B(new_n2785), .Y(new_n3275));
  not_8  g00927(.A(n22379), .Y(new_n3276));
  nand_5 g00928(.A(new_n3276), .B(n767), .Y(new_n3277));
  nand_5 g00929(.A(new_n3277), .B(new_n3275), .Y(new_n3278));
  xnor_4 g00930(.A(new_n3278), .B(new_n3274), .Y(new_n3279_1));
  nand_5 g00931(.A(new_n3203), .B(new_n3180), .Y(new_n3280));
  nand_5 g00932(.A(new_n3280), .B(new_n3201), .Y(new_n3281));
  not_8  g00933(.A(new_n3281), .Y(new_n3282));
  nand_5 g00934(.A(new_n3184), .B(new_n3182), .Y(new_n3283));
  nand_5 g00935(.A(new_n3283), .B(new_n3187), .Y(new_n3284));
  not_8  g00936(.A(new_n3284), .Y(new_n3285));
  not_8  g00937(.A(n6814), .Y(new_n3286));
  not_8  g00938(.A(n10763), .Y(new_n3287));
  nand_5 g00939(.A(new_n3287), .B(new_n3286), .Y(new_n3288));
  nand_5 g00940(.A(n10763), .B(n6814), .Y(new_n3289_1));
  nand_5 g00941(.A(new_n3289_1), .B(new_n3288), .Y(new_n3290));
  xor_4  g00942(.A(new_n3290), .B(new_n3285), .Y(new_n3291));
  not_8  g00943(.A(new_n3193), .Y(new_n3292));
  nand_5 g00944(.A(new_n3197), .B(new_n3292), .Y(new_n3293));
  nand_5 g00945(.A(new_n3293), .B(new_n3196), .Y(new_n3294));
  not_8  g00946(.A(n12657), .Y(new_n3295));
  not_8  g00947(.A(n27089), .Y(new_n3296));
  nand_5 g00948(.A(new_n3296), .B(new_n3295), .Y(new_n3297));
  nand_5 g00949(.A(n27089), .B(n12657), .Y(new_n3298));
  nand_5 g00950(.A(new_n3298), .B(new_n3297), .Y(new_n3299));
  xor_4  g00951(.A(new_n3299), .B(new_n3294), .Y(new_n3300));
  nand_5 g00952(.A(new_n3300), .B(new_n3291), .Y(new_n3301_1));
  not_8  g00953(.A(new_n3291), .Y(new_n3302));
  not_8  g00954(.A(new_n3300), .Y(new_n3303));
  nand_5 g00955(.A(new_n3303), .B(new_n3302), .Y(new_n3304));
  nand_5 g00956(.A(new_n3304), .B(new_n3301_1), .Y(new_n3305));
  xor_4  g00957(.A(new_n3305), .B(new_n3282), .Y(new_n3306_1));
  not_8  g00958(.A(new_n3306_1), .Y(new_n3307));
  nand_5 g00959(.A(new_n3307), .B(new_n3279_1), .Y(new_n3308));
  not_8  g00960(.A(new_n3308), .Y(new_n3309));
  nor_5  g00961(.A(new_n3307), .B(new_n3279_1), .Y(new_n3310));
  nor_5  g00962(.A(new_n3310), .B(new_n3309), .Y(new_n3311));
  xor_4  g00963(.A(new_n3311), .B(new_n3272), .Y(n142));
  not_8  g00964(.A(n4319), .Y(new_n3313));
  not_8  g00965(.A(n7335), .Y(new_n3314));
  nand_5 g00966(.A(new_n3314), .B(new_n3313), .Y(new_n3315));
  nand_5 g00967(.A(n7335), .B(n4319), .Y(new_n3316_1));
  not_8  g00968(.A(n5696), .Y(new_n3317));
  not_8  g00969(.A(n23463), .Y(new_n3318));
  nand_5 g00970(.A(new_n3318), .B(new_n3317), .Y(new_n3319));
  nand_5 g00971(.A(n23463), .B(n5696), .Y(new_n3320_1));
  not_8  g00972(.A(n13074), .Y(new_n3321));
  not_8  g00973(.A(n13367), .Y(new_n3322));
  nand_5 g00974(.A(new_n3322), .B(new_n3321), .Y(new_n3323));
  nand_5 g00975(.A(n13367), .B(n13074), .Y(new_n3324_1));
  not_8  g00976(.A(n932), .Y(new_n3325));
  nand_5 g00977(.A(new_n2601), .B(new_n3325), .Y(new_n3326));
  nand_5 g00978(.A(n10739), .B(n932), .Y(new_n3327));
  not_8  g00979(.A(n6691), .Y(new_n3328));
  nand_5 g00980(.A(new_n2518), .B(new_n3328), .Y(new_n3329));
  nand_5 g00981(.A(n21753), .B(n6691), .Y(new_n3330));
  not_8  g00982(.A(n3260), .Y(new_n3331));
  nand_5 g00983(.A(new_n2492), .B(new_n3331), .Y(new_n3332_1));
  nand_5 g00984(.A(n21832), .B(n3260), .Y(new_n3333));
  not_8  g00985(.A(n20489), .Y(new_n3334));
  nand_5 g00986(.A(new_n2496), .B(new_n3334), .Y(new_n3335));
  nand_5 g00987(.A(n26913), .B(n20489), .Y(new_n3336));
  not_8  g00988(.A(n2355), .Y(new_n3337));
  nand_5 g00989(.A(new_n2500), .B(new_n3337), .Y(new_n3338));
  nand_5 g00990(.A(n16223), .B(n2355), .Y(new_n3339));
  not_8  g00991(.A(n11121), .Y(new_n3340_1));
  nand_5 g00992(.A(new_n2504), .B(new_n3340_1), .Y(new_n3341));
  nand_5 g00993(.A(n19494), .B(n11121), .Y(new_n3342));
  nand_5 g00994(.A(n16217), .B(n2387), .Y(new_n3343_1));
  nand_5 g00995(.A(new_n3343_1), .B(new_n3342), .Y(new_n3344));
  nand_5 g00996(.A(new_n3344), .B(new_n3341), .Y(new_n3345));
  nand_5 g00997(.A(new_n3345), .B(new_n3339), .Y(new_n3346));
  nand_5 g00998(.A(new_n3346), .B(new_n3338), .Y(new_n3347));
  nand_5 g00999(.A(new_n3347), .B(new_n3336), .Y(new_n3348));
  nand_5 g01000(.A(new_n3348), .B(new_n3335), .Y(new_n3349_1));
  nand_5 g01001(.A(new_n3349_1), .B(new_n3333), .Y(new_n3350));
  nand_5 g01002(.A(new_n3350), .B(new_n3332_1), .Y(new_n3351));
  nand_5 g01003(.A(new_n3351), .B(new_n3330), .Y(new_n3352));
  nand_5 g01004(.A(new_n3352), .B(new_n3329), .Y(new_n3353));
  nand_5 g01005(.A(new_n3353), .B(new_n3327), .Y(new_n3354));
  nand_5 g01006(.A(new_n3354), .B(new_n3326), .Y(new_n3355));
  nand_5 g01007(.A(new_n3355), .B(new_n3324_1), .Y(new_n3356));
  nand_5 g01008(.A(new_n3356), .B(new_n3323), .Y(new_n3357));
  nand_5 g01009(.A(new_n3357), .B(new_n3320_1), .Y(new_n3358));
  nand_5 g01010(.A(new_n3358), .B(new_n3319), .Y(new_n3359));
  nand_5 g01011(.A(new_n3359), .B(new_n3316_1), .Y(new_n3360));
  nand_5 g01012(.A(new_n3360), .B(new_n3315), .Y(new_n3361));
  nand_5 g01013(.A(new_n3316_1), .B(new_n3315), .Y(new_n3362));
  xor_4  g01014(.A(new_n3362), .B(new_n3359), .Y(new_n3363));
  not_8  g01015(.A(new_n3363), .Y(new_n3364));
  or_5   g01016(.A(new_n3364), .B(n5025), .Y(new_n3365));
  nand_5 g01017(.A(new_n3364), .B(n5025), .Y(new_n3366_1));
  not_8  g01018(.A(n6485), .Y(new_n3367));
  nand_5 g01019(.A(new_n3320_1), .B(new_n3319), .Y(new_n3368));
  xor_4  g01020(.A(new_n3368), .B(new_n3357), .Y(new_n3369));
  nand_5 g01021(.A(new_n3369), .B(new_n3367), .Y(new_n3370));
  not_8  g01022(.A(new_n3369), .Y(new_n3371));
  nand_5 g01023(.A(new_n3371), .B(n6485), .Y(new_n3372));
  not_8  g01024(.A(n26036), .Y(new_n3373));
  nand_5 g01025(.A(new_n3324_1), .B(new_n3323), .Y(new_n3374));
  xor_4  g01026(.A(new_n3374), .B(new_n3355), .Y(new_n3375));
  nand_5 g01027(.A(new_n3375), .B(new_n3373), .Y(new_n3376));
  not_8  g01028(.A(new_n3375), .Y(new_n3377));
  nand_5 g01029(.A(new_n3377), .B(n26036), .Y(new_n3378));
  not_8  g01030(.A(n19770), .Y(new_n3379));
  nand_5 g01031(.A(new_n3327), .B(new_n3326), .Y(new_n3380));
  xor_4  g01032(.A(new_n3380), .B(new_n3353), .Y(new_n3381));
  nand_5 g01033(.A(new_n3381), .B(new_n3379), .Y(new_n3382));
  not_8  g01034(.A(new_n3381), .Y(new_n3383));
  nand_5 g01035(.A(new_n3383), .B(n19770), .Y(new_n3384));
  not_8  g01036(.A(n8782), .Y(new_n3385));
  nand_5 g01037(.A(new_n3330), .B(new_n3329), .Y(new_n3386));
  xor_4  g01038(.A(new_n3386), .B(new_n3351), .Y(new_n3387));
  nand_5 g01039(.A(new_n3387), .B(new_n3385), .Y(new_n3388));
  not_8  g01040(.A(new_n3387), .Y(new_n3389));
  nand_5 g01041(.A(new_n3389), .B(n8782), .Y(new_n3390_1));
  not_8  g01042(.A(n8678), .Y(new_n3391));
  nand_5 g01043(.A(new_n3333), .B(new_n3332_1), .Y(new_n3392));
  xor_4  g01044(.A(new_n3392), .B(new_n3349_1), .Y(new_n3393));
  nand_5 g01045(.A(new_n3393), .B(new_n3391), .Y(new_n3394));
  not_8  g01046(.A(new_n3393), .Y(new_n3395));
  nand_5 g01047(.A(new_n3395), .B(n8678), .Y(new_n3396));
  not_8  g01048(.A(n1432), .Y(new_n3397));
  nand_5 g01049(.A(new_n3336), .B(new_n3335), .Y(new_n3398));
  xor_4  g01050(.A(new_n3398), .B(new_n3347), .Y(new_n3399));
  nand_5 g01051(.A(new_n3399), .B(new_n3397), .Y(new_n3400));
  not_8  g01052(.A(new_n3399), .Y(new_n3401));
  nand_5 g01053(.A(new_n3401), .B(n1432), .Y(new_n3402));
  not_8  g01054(.A(n21599), .Y(new_n3403));
  nand_5 g01055(.A(new_n3339), .B(new_n3338), .Y(new_n3404));
  xor_4  g01056(.A(new_n3404), .B(new_n3345), .Y(new_n3405));
  nand_5 g01057(.A(new_n3405), .B(new_n3403), .Y(new_n3406));
  not_8  g01058(.A(new_n3405), .Y(new_n3407));
  nand_5 g01059(.A(new_n3407), .B(n21599), .Y(new_n3408));
  not_8  g01060(.A(n11424), .Y(new_n3409));
  not_8  g01061(.A(n16217), .Y(new_n3410));
  nand_5 g01062(.A(new_n3410), .B(new_n2506), .Y(new_n3411));
  and_5  g01063(.A(new_n3411), .B(new_n3343_1), .Y(new_n3412));
  nand_5 g01064(.A(new_n3412), .B(new_n3409), .Y(new_n3413));
  nor_5  g01065(.A(new_n3413), .B(n25336), .Y(new_n3414));
  not_8  g01066(.A(new_n3414), .Y(new_n3415));
  nand_5 g01067(.A(new_n3413), .B(n25336), .Y(new_n3416));
  nand_5 g01068(.A(new_n3342), .B(new_n3341), .Y(new_n3417));
  not_8  g01069(.A(new_n3417), .Y(new_n3418));
  xor_4  g01070(.A(new_n3418), .B(new_n3343_1), .Y(new_n3419));
  not_8  g01071(.A(new_n3419), .Y(new_n3420));
  nand_5 g01072(.A(new_n3420), .B(new_n3416), .Y(new_n3421));
  nand_5 g01073(.A(new_n3421), .B(new_n3415), .Y(new_n3422));
  nand_5 g01074(.A(new_n3422), .B(new_n3408), .Y(new_n3423));
  nand_5 g01075(.A(new_n3423), .B(new_n3406), .Y(new_n3424));
  nand_5 g01076(.A(new_n3424), .B(new_n3402), .Y(new_n3425_1));
  nand_5 g01077(.A(new_n3425_1), .B(new_n3400), .Y(new_n3426_1));
  nand_5 g01078(.A(new_n3426_1), .B(new_n3396), .Y(new_n3427));
  nand_5 g01079(.A(new_n3427), .B(new_n3394), .Y(new_n3428));
  nand_5 g01080(.A(new_n3428), .B(new_n3390_1), .Y(new_n3429));
  nand_5 g01081(.A(new_n3429), .B(new_n3388), .Y(new_n3430));
  nand_5 g01082(.A(new_n3430), .B(new_n3384), .Y(new_n3431));
  nand_5 g01083(.A(new_n3431), .B(new_n3382), .Y(new_n3432));
  nand_5 g01084(.A(new_n3432), .B(new_n3378), .Y(new_n3433));
  nand_5 g01085(.A(new_n3433), .B(new_n3376), .Y(new_n3434));
  nand_5 g01086(.A(new_n3434), .B(new_n3372), .Y(new_n3435));
  nand_5 g01087(.A(new_n3435), .B(new_n3370), .Y(new_n3436));
  nand_5 g01088(.A(new_n3436), .B(new_n3366_1), .Y(new_n3437));
  nand_5 g01089(.A(new_n3437), .B(new_n3365), .Y(new_n3438));
  not_8  g01090(.A(new_n3438), .Y(new_n3439));
  nand_5 g01091(.A(new_n3439), .B(new_n3361), .Y(new_n3440));
  not_8  g01092(.A(new_n3440), .Y(new_n3441));
  not_8  g01093(.A(n9967), .Y(new_n3442));
  nand_5 g01094(.A(new_n2443), .B(new_n2357), .Y(new_n3443));
  or_5   g01095(.A(new_n3443), .B(n24618), .Y(new_n3444));
  nor_5  g01096(.A(new_n3444), .B(n24278), .Y(new_n3445));
  nand_5 g01097(.A(new_n3445), .B(new_n2371), .Y(new_n3446));
  nor_5  g01098(.A(new_n3446), .B(n26823), .Y(new_n3447));
  nand_5 g01099(.A(new_n3447), .B(new_n2584), .Y(new_n3448));
  nor_5  g01100(.A(new_n3448), .B(n20946), .Y(new_n3449));
  nand_5 g01101(.A(new_n3449), .B(new_n3442), .Y(new_n3450));
  nor_5  g01102(.A(new_n3450), .B(n3425), .Y(new_n3451_1));
  not_8  g01103(.A(new_n3451_1), .Y(new_n3452));
  nand_5 g01104(.A(new_n3450), .B(n3425), .Y(new_n3453));
  and_5  g01105(.A(new_n3453), .B(new_n3452), .Y(new_n3454));
  not_8  g01106(.A(new_n3454), .Y(new_n3455));
  nand_5 g01107(.A(new_n3365), .B(new_n3366_1), .Y(new_n3456));
  xor_4  g01108(.A(new_n3456), .B(new_n3436), .Y(new_n3457));
  not_8  g01109(.A(new_n3457), .Y(new_n3458));
  nand_5 g01110(.A(new_n3458), .B(new_n3455), .Y(new_n3459_1));
  xor_4  g01111(.A(new_n3449), .B(new_n3442), .Y(new_n3460_1));
  nand_5 g01112(.A(new_n3370), .B(new_n3372), .Y(new_n3461));
  xor_4  g01113(.A(new_n3461), .B(new_n3434), .Y(new_n3462));
  nand_5 g01114(.A(new_n3462), .B(new_n3460_1), .Y(new_n3463));
  not_8  g01115(.A(new_n3460_1), .Y(new_n3464));
  not_8  g01116(.A(new_n3462), .Y(new_n3465));
  nand_5 g01117(.A(new_n3465), .B(new_n3464), .Y(new_n3466));
  xor_4  g01118(.A(new_n3448), .B(n20946), .Y(new_n3467));
  nand_5 g01119(.A(new_n3376), .B(new_n3378), .Y(new_n3468_1));
  xor_4  g01120(.A(new_n3468_1), .B(new_n3432), .Y(new_n3469));
  nand_5 g01121(.A(new_n3469), .B(new_n3467), .Y(new_n3470));
  not_8  g01122(.A(new_n3467), .Y(new_n3471));
  not_8  g01123(.A(new_n3469), .Y(new_n3472));
  nand_5 g01124(.A(new_n3472), .B(new_n3471), .Y(new_n3473));
  xor_4  g01125(.A(new_n3447), .B(new_n2584), .Y(new_n3474));
  nand_5 g01126(.A(new_n3382), .B(new_n3384), .Y(new_n3475));
  xor_4  g01127(.A(new_n3475), .B(new_n3430), .Y(new_n3476));
  nand_5 g01128(.A(new_n3476), .B(new_n3474), .Y(new_n3477));
  not_8  g01129(.A(new_n3474), .Y(new_n3478));
  not_8  g01130(.A(new_n3476), .Y(new_n3479));
  nand_5 g01131(.A(new_n3479), .B(new_n3478), .Y(new_n3480_1));
  xor_4  g01132(.A(new_n3446), .B(n26823), .Y(new_n3481));
  nand_5 g01133(.A(new_n3388), .B(new_n3390_1), .Y(new_n3482));
  xor_4  g01134(.A(new_n3482), .B(new_n3428), .Y(new_n3483));
  nand_5 g01135(.A(new_n3483), .B(new_n3481), .Y(new_n3484));
  not_8  g01136(.A(new_n3481), .Y(new_n3485));
  not_8  g01137(.A(new_n3483), .Y(new_n3486));
  nand_5 g01138(.A(new_n3486), .B(new_n3485), .Y(new_n3487));
  xor_4  g01139(.A(new_n3445), .B(new_n2371), .Y(new_n3488));
  nand_5 g01140(.A(new_n3394), .B(new_n3396), .Y(new_n3489));
  xor_4  g01141(.A(new_n3489), .B(new_n3426_1), .Y(new_n3490));
  nand_5 g01142(.A(new_n3490), .B(new_n3488), .Y(new_n3491));
  not_8  g01143(.A(new_n3488), .Y(new_n3492));
  not_8  g01144(.A(new_n3490), .Y(new_n3493));
  nand_5 g01145(.A(new_n3493), .B(new_n3492), .Y(new_n3494));
  xor_4  g01146(.A(new_n3444), .B(n24278), .Y(new_n3495));
  nand_5 g01147(.A(new_n3400), .B(new_n3402), .Y(new_n3496));
  xor_4  g01148(.A(new_n3496), .B(new_n3424), .Y(new_n3497));
  nand_5 g01149(.A(new_n3497), .B(new_n3495), .Y(new_n3498));
  or_5   g01150(.A(new_n3497), .B(new_n3495), .Y(new_n3499));
  nand_5 g01151(.A(new_n3443), .B(n24618), .Y(new_n3500));
  and_5  g01152(.A(new_n3500), .B(new_n3444), .Y(new_n3501));
  nand_5 g01153(.A(new_n3406), .B(new_n3408), .Y(new_n3502_1));
  xor_4  g01154(.A(new_n3502_1), .B(new_n3422), .Y(new_n3503));
  nand_5 g01155(.A(new_n3503), .B(new_n3501), .Y(new_n3504));
  or_5   g01156(.A(new_n3503), .B(new_n3501), .Y(new_n3505));
  or_5   g01157(.A(new_n3412), .B(new_n3409), .Y(new_n3506_1));
  and_5  g01158(.A(new_n3506_1), .B(new_n3413), .Y(new_n3507));
  not_8  g01159(.A(new_n3507), .Y(new_n3508));
  nand_5 g01160(.A(new_n3508), .B(n12315), .Y(new_n3509));
  nand_5 g01161(.A(n12315), .B(n3952), .Y(new_n3510));
  and_5  g01162(.A(new_n3510), .B(new_n3443), .Y(new_n3511));
  not_8  g01163(.A(new_n3511), .Y(new_n3512));
  nand_5 g01164(.A(new_n3512), .B(new_n3509), .Y(new_n3513));
  nor_5  g01165(.A(new_n3509), .B(n3952), .Y(new_n3514));
  not_8  g01166(.A(new_n3514), .Y(new_n3515));
  nand_5 g01167(.A(new_n3415), .B(new_n3416), .Y(new_n3516_1));
  xor_4  g01168(.A(new_n3516_1), .B(new_n3419), .Y(new_n3517));
  nand_5 g01169(.A(new_n3517), .B(new_n3515), .Y(new_n3518));
  nand_5 g01170(.A(new_n3518), .B(new_n3513), .Y(new_n3519));
  not_8  g01171(.A(new_n3519), .Y(new_n3520));
  nand_5 g01172(.A(new_n3520), .B(new_n3505), .Y(new_n3521));
  nand_5 g01173(.A(new_n3521), .B(new_n3504), .Y(new_n3522));
  nand_5 g01174(.A(new_n3522), .B(new_n3499), .Y(new_n3523));
  nand_5 g01175(.A(new_n3523), .B(new_n3498), .Y(new_n3524));
  nand_5 g01176(.A(new_n3524), .B(new_n3494), .Y(new_n3525));
  nand_5 g01177(.A(new_n3525), .B(new_n3491), .Y(new_n3526));
  nand_5 g01178(.A(new_n3526), .B(new_n3487), .Y(new_n3527));
  nand_5 g01179(.A(new_n3527), .B(new_n3484), .Y(new_n3528_1));
  nand_5 g01180(.A(new_n3528_1), .B(new_n3480_1), .Y(new_n3529));
  nand_5 g01181(.A(new_n3529), .B(new_n3477), .Y(new_n3530));
  nand_5 g01182(.A(new_n3530), .B(new_n3473), .Y(new_n3531));
  nand_5 g01183(.A(new_n3531), .B(new_n3470), .Y(new_n3532));
  nand_5 g01184(.A(new_n3532), .B(new_n3466), .Y(new_n3533));
  nand_5 g01185(.A(new_n3533), .B(new_n3463), .Y(new_n3534));
  nand_5 g01186(.A(new_n3534), .B(new_n3459_1), .Y(new_n3535));
  not_8  g01187(.A(new_n3535), .Y(new_n3536));
  nand_5 g01188(.A(new_n3457), .B(new_n3454), .Y(new_n3537));
  nand_5 g01189(.A(new_n3537), .B(new_n3452), .Y(new_n3538));
  nor_5  g01190(.A(new_n3538), .B(new_n3536), .Y(new_n3539));
  nand_5 g01191(.A(new_n3539), .B(new_n3441), .Y(new_n3540));
  not_8  g01192(.A(n5101), .Y(new_n3541_1));
  not_8  g01193(.A(n7593), .Y(new_n3542));
  nand_5 g01194(.A(new_n3542), .B(new_n3541_1), .Y(new_n3543));
  nand_5 g01195(.A(n7593), .B(n5101), .Y(new_n3544));
  not_8  g01196(.A(n3228), .Y(new_n3545));
  not_8  g01197(.A(n6861), .Y(new_n3546));
  not_8  g01198(.A(n2328), .Y(new_n3547));
  not_8  g01199(.A(n14603), .Y(new_n3548));
  not_8  g01200(.A(n15053), .Y(new_n3549));
  nand_5 g01201(.A(new_n3549), .B(new_n3548), .Y(new_n3550));
  nand_5 g01202(.A(n15053), .B(n14603), .Y(new_n3551));
  not_8  g01203(.A(n20794), .Y(new_n3552));
  not_8  g01204(.A(n25471), .Y(new_n3553));
  nand_5 g01205(.A(new_n3553), .B(new_n3552), .Y(new_n3554));
  nand_5 g01206(.A(n25471), .B(n20794), .Y(new_n3555_1));
  nand_5 g01207(.A(n23333), .B(n16502), .Y(new_n3556));
  nand_5 g01208(.A(new_n3556), .B(new_n3555_1), .Y(new_n3557));
  nand_5 g01209(.A(new_n3557), .B(new_n3554), .Y(new_n3558));
  nand_5 g01210(.A(new_n3558), .B(new_n3551), .Y(new_n3559));
  nand_5 g01211(.A(new_n3559), .B(new_n3550), .Y(new_n3560));
  nand_5 g01212(.A(new_n3560), .B(new_n3547), .Y(new_n3561_1));
  not_8  g01213(.A(new_n3561_1), .Y(new_n3562));
  nor_5  g01214(.A(new_n3560), .B(new_n3547), .Y(new_n3563_1));
  nor_5  g01215(.A(new_n3563_1), .B(n18737), .Y(new_n3564));
  nor_5  g01216(.A(new_n3564), .B(new_n3562), .Y(new_n3565));
  or_5   g01217(.A(new_n3565), .B(n19357), .Y(new_n3566));
  not_8  g01218(.A(n21471), .Y(new_n3567));
  nand_5 g01219(.A(new_n3565), .B(n19357), .Y(new_n3568));
  nand_5 g01220(.A(new_n3568), .B(new_n3567), .Y(new_n3569));
  nand_5 g01221(.A(new_n3569), .B(new_n3566), .Y(new_n3570_1));
  nand_5 g01222(.A(new_n3570_1), .B(new_n3546), .Y(new_n3571));
  not_8  g01223(.A(new_n3571), .Y(new_n3572));
  nor_5  g01224(.A(new_n3570_1), .B(new_n3546), .Y(new_n3573));
  nor_5  g01225(.A(new_n3573), .B(n25738), .Y(new_n3574));
  nor_5  g01226(.A(new_n3574), .B(new_n3572), .Y(new_n3575));
  or_5   g01227(.A(new_n3575), .B(n5302), .Y(new_n3576));
  not_8  g01228(.A(n19116), .Y(new_n3577));
  nand_5 g01229(.A(new_n3575), .B(n5302), .Y(new_n3578));
  nand_5 g01230(.A(new_n3578), .B(new_n3577), .Y(new_n3579));
  nand_5 g01231(.A(new_n3579), .B(new_n3576), .Y(new_n3580));
  nand_5 g01232(.A(new_n3580), .B(new_n3545), .Y(new_n3581));
  not_8  g01233(.A(new_n3581), .Y(new_n3582_1));
  nor_5  g01234(.A(new_n3580), .B(new_n3545), .Y(new_n3583));
  nor_5  g01235(.A(new_n3583), .B(n22470), .Y(new_n3584));
  nor_5  g01236(.A(new_n3584), .B(new_n3582_1), .Y(new_n3585));
  or_5   g01237(.A(new_n3585), .B(n337), .Y(new_n3586));
  not_8  g01238(.A(n16507), .Y(new_n3587));
  nand_5 g01239(.A(new_n3585), .B(n337), .Y(new_n3588));
  nand_5 g01240(.A(new_n3588), .B(new_n3587), .Y(new_n3589));
  nand_5 g01241(.A(new_n3589), .B(new_n3586), .Y(new_n3590));
  nand_5 g01242(.A(new_n3590), .B(new_n3544), .Y(new_n3591));
  nand_5 g01243(.A(new_n3591), .B(new_n3543), .Y(new_n3592));
  not_8  g01244(.A(new_n3361), .Y(new_n3593));
  nand_5 g01245(.A(new_n3438), .B(new_n3593), .Y(new_n3594));
  and_5  g01246(.A(new_n3594), .B(new_n3440), .Y(new_n3595));
  not_8  g01247(.A(new_n3595), .Y(new_n3596));
  xor_4  g01248(.A(new_n3596), .B(new_n3539), .Y(new_n3597));
  or_5   g01249(.A(new_n3597), .B(new_n3592), .Y(new_n3598));
  nand_5 g01250(.A(new_n3597), .B(new_n3592), .Y(new_n3599));
  nand_5 g01251(.A(new_n3544), .B(new_n3543), .Y(new_n3600));
  xor_4  g01252(.A(new_n3600), .B(new_n3590), .Y(new_n3601));
  not_8  g01253(.A(new_n3601), .Y(new_n3602));
  nand_5 g01254(.A(new_n3537), .B(new_n3459_1), .Y(new_n3603));
  xor_4  g01255(.A(new_n3603), .B(new_n3534), .Y(new_n3604));
  or_5   g01256(.A(new_n3604), .B(new_n3602), .Y(new_n3605));
  nand_5 g01257(.A(new_n3604), .B(new_n3602), .Y(new_n3606));
  nand_5 g01258(.A(new_n3588), .B(new_n3586), .Y(new_n3607));
  xor_4  g01259(.A(new_n3607), .B(n16507), .Y(new_n3608));
  nand_5 g01260(.A(new_n3463), .B(new_n3466), .Y(new_n3609));
  xor_4  g01261(.A(new_n3609), .B(new_n3532), .Y(new_n3610));
  or_5   g01262(.A(new_n3610), .B(new_n3608), .Y(new_n3611));
  nand_5 g01263(.A(new_n3610), .B(new_n3608), .Y(new_n3612));
  not_8  g01264(.A(n22470), .Y(new_n3613));
  nor_5  g01265(.A(new_n3583), .B(new_n3582_1), .Y(new_n3614));
  xor_4  g01266(.A(new_n3614), .B(new_n3613), .Y(new_n3615));
  nand_5 g01267(.A(new_n3470), .B(new_n3473), .Y(new_n3616));
  xor_4  g01268(.A(new_n3616), .B(new_n3530), .Y(new_n3617_1));
  or_5   g01269(.A(new_n3617_1), .B(new_n3615), .Y(new_n3618_1));
  nand_5 g01270(.A(new_n3617_1), .B(new_n3615), .Y(new_n3619));
  nand_5 g01271(.A(new_n3578), .B(new_n3576), .Y(new_n3620));
  xor_4  g01272(.A(new_n3620), .B(n19116), .Y(new_n3621));
  nand_5 g01273(.A(new_n3477), .B(new_n3480_1), .Y(new_n3622));
  xor_4  g01274(.A(new_n3622), .B(new_n3528_1), .Y(new_n3623));
  or_5   g01275(.A(new_n3623), .B(new_n3621), .Y(new_n3624));
  nand_5 g01276(.A(new_n3623), .B(new_n3621), .Y(new_n3625));
  not_8  g01277(.A(n25738), .Y(new_n3626));
  nor_5  g01278(.A(new_n3573), .B(new_n3572), .Y(new_n3627));
  xor_4  g01279(.A(new_n3627), .B(new_n3626), .Y(new_n3628));
  nand_5 g01280(.A(new_n3484), .B(new_n3487), .Y(new_n3629));
  xor_4  g01281(.A(new_n3629), .B(new_n3526), .Y(new_n3630));
  or_5   g01282(.A(new_n3630), .B(new_n3628), .Y(new_n3631));
  nand_5 g01283(.A(new_n3630), .B(new_n3628), .Y(new_n3632));
  nand_5 g01284(.A(new_n3568), .B(new_n3566), .Y(new_n3633));
  xor_4  g01285(.A(new_n3633), .B(n21471), .Y(new_n3634));
  nand_5 g01286(.A(new_n3491), .B(new_n3494), .Y(new_n3635));
  xor_4  g01287(.A(new_n3635), .B(new_n3524), .Y(new_n3636));
  or_5   g01288(.A(new_n3636), .B(new_n3634), .Y(new_n3637));
  nand_5 g01289(.A(new_n3636), .B(new_n3634), .Y(new_n3638));
  not_8  g01290(.A(n18737), .Y(new_n3639));
  nor_5  g01291(.A(new_n3563_1), .B(new_n3562), .Y(new_n3640));
  xor_4  g01292(.A(new_n3640), .B(new_n3639), .Y(new_n3641));
  nand_5 g01293(.A(new_n3498), .B(new_n3499), .Y(new_n3642_1));
  xor_4  g01294(.A(new_n3642_1), .B(new_n3522), .Y(new_n3643));
  or_5   g01295(.A(new_n3643), .B(new_n3641), .Y(new_n3644));
  nand_5 g01296(.A(new_n3643), .B(new_n3641), .Y(new_n3645));
  nand_5 g01297(.A(new_n3551), .B(new_n3550), .Y(new_n3646));
  xor_4  g01298(.A(new_n3646), .B(new_n3558), .Y(new_n3647));
  not_8  g01299(.A(new_n3647), .Y(new_n3648));
  nand_5 g01300(.A(new_n3504), .B(new_n3505), .Y(new_n3649_1));
  xor_4  g01301(.A(new_n3649_1), .B(new_n3520), .Y(new_n3650));
  or_5   g01302(.A(new_n3650), .B(new_n3648), .Y(new_n3651));
  nand_5 g01303(.A(new_n3650), .B(new_n3648), .Y(new_n3652));
  not_8  g01304(.A(n16502), .Y(new_n3653));
  not_8  g01305(.A(n23333), .Y(new_n3654));
  nand_5 g01306(.A(new_n3654), .B(new_n3653), .Y(new_n3655));
  nand_5 g01307(.A(new_n3655), .B(new_n3556), .Y(new_n3656));
  nand_5 g01308(.A(new_n3507), .B(new_n2443), .Y(new_n3657));
  nand_5 g01309(.A(new_n3657), .B(new_n3509), .Y(new_n3658));
  nor_5  g01310(.A(new_n3658), .B(new_n3656), .Y(new_n3659));
  nand_5 g01311(.A(new_n3555_1), .B(new_n3554), .Y(new_n3660));
  not_8  g01312(.A(new_n3660), .Y(new_n3661));
  nand_5 g01313(.A(new_n3661), .B(new_n3659), .Y(new_n3662));
  xor_4  g01314(.A(new_n3660), .B(new_n3556), .Y(new_n3663));
  nor_5  g01315(.A(new_n3663), .B(new_n3659), .Y(new_n3664));
  not_8  g01316(.A(new_n3664), .Y(new_n3665_1));
  nand_5 g01317(.A(new_n3515), .B(new_n3513), .Y(new_n3666));
  xor_4  g01318(.A(new_n3666), .B(new_n3517), .Y(new_n3667));
  nand_5 g01319(.A(new_n3667), .B(new_n3665_1), .Y(new_n3668));
  nand_5 g01320(.A(new_n3668), .B(new_n3662), .Y(new_n3669));
  nand_5 g01321(.A(new_n3669), .B(new_n3652), .Y(new_n3670));
  nand_5 g01322(.A(new_n3670), .B(new_n3651), .Y(new_n3671));
  nand_5 g01323(.A(new_n3671), .B(new_n3645), .Y(new_n3672));
  nand_5 g01324(.A(new_n3672), .B(new_n3644), .Y(new_n3673));
  nand_5 g01325(.A(new_n3673), .B(new_n3638), .Y(new_n3674));
  nand_5 g01326(.A(new_n3674), .B(new_n3637), .Y(new_n3675));
  nand_5 g01327(.A(new_n3675), .B(new_n3632), .Y(new_n3676));
  nand_5 g01328(.A(new_n3676), .B(new_n3631), .Y(new_n3677));
  nand_5 g01329(.A(new_n3677), .B(new_n3625), .Y(new_n3678));
  nand_5 g01330(.A(new_n3678), .B(new_n3624), .Y(new_n3679_1));
  nand_5 g01331(.A(new_n3679_1), .B(new_n3619), .Y(new_n3680));
  nand_5 g01332(.A(new_n3680), .B(new_n3618_1), .Y(new_n3681));
  nand_5 g01333(.A(new_n3681), .B(new_n3612), .Y(new_n3682));
  nand_5 g01334(.A(new_n3682), .B(new_n3611), .Y(new_n3683));
  nand_5 g01335(.A(new_n3683), .B(new_n3606), .Y(new_n3684));
  nand_5 g01336(.A(new_n3684), .B(new_n3605), .Y(new_n3685));
  nand_5 g01337(.A(new_n3685), .B(new_n3599), .Y(new_n3686));
  nand_5 g01338(.A(new_n3686), .B(new_n3598), .Y(new_n3687));
  nor_5  g01339(.A(new_n3539), .B(new_n3441), .Y(new_n3688));
  nand_5 g01340(.A(new_n3596), .B(new_n3540), .Y(new_n3689));
  nor_5  g01341(.A(new_n3689), .B(new_n3688), .Y(new_n3690));
  not_8  g01342(.A(new_n3690), .Y(new_n3691));
  nand_5 g01343(.A(new_n3691), .B(new_n3687), .Y(new_n3692));
  xor_4  g01344(.A(new_n3692), .B(new_n3540), .Y(n175));
  not_8  g01345(.A(n21489), .Y(new_n3694));
  not_8  g01346(.A(n13912), .Y(new_n3695));
  not_8  g01347(.A(n9598), .Y(new_n3696));
  not_8  g01348(.A(n21993), .Y(new_n3697));
  not_8  g01349(.A(n25565), .Y(new_n3698));
  nand_5 g01350(.A(new_n3698), .B(new_n3697), .Y(new_n3699));
  or_5   g01351(.A(new_n3699), .B(n11273), .Y(new_n3700));
  nor_5  g01352(.A(new_n3700), .B(n22290), .Y(new_n3701));
  nand_5 g01353(.A(new_n3701), .B(new_n3696), .Y(new_n3702));
  nor_5  g01354(.A(new_n3702), .B(n7670), .Y(new_n3703));
  nand_5 g01355(.A(new_n3703), .B(new_n3695), .Y(new_n3704));
  nor_5  g01356(.A(new_n3704), .B(n20213), .Y(new_n3705));
  nand_5 g01357(.A(new_n3705), .B(new_n3694), .Y(new_n3706));
  nor_5  g01358(.A(new_n3706), .B(n9259), .Y(new_n3707));
  not_8  g01359(.A(new_n3707), .Y(new_n3708));
  nand_5 g01360(.A(new_n3706), .B(n9259), .Y(new_n3709));
  and_5  g01361(.A(new_n3709), .B(new_n3708), .Y(new_n3710_1));
  not_8  g01362(.A(n3506), .Y(new_n3711));
  nand_5 g01363(.A(new_n3711), .B(n2743), .Y(new_n3712));
  not_8  g01364(.A(n2743), .Y(new_n3713));
  nand_5 g01365(.A(n3506), .B(new_n3713), .Y(new_n3714));
  nand_5 g01366(.A(new_n3714), .B(new_n3712), .Y(new_n3715));
  not_8  g01367(.A(n14899), .Y(new_n3716));
  nand_5 g01368(.A(new_n3716), .B(n7026), .Y(new_n3717));
  not_8  g01369(.A(n7026), .Y(new_n3718));
  nand_5 g01370(.A(n14899), .B(new_n3718), .Y(new_n3719));
  not_8  g01371(.A(n18444), .Y(new_n3720));
  nand_5 g01372(.A(new_n3720), .B(n13719), .Y(new_n3721));
  not_8  g01373(.A(n13719), .Y(new_n3722));
  nand_5 g01374(.A(n18444), .B(new_n3722), .Y(new_n3723));
  not_8  g01375(.A(n24638), .Y(new_n3724));
  nand_5 g01376(.A(new_n3724), .B(n442), .Y(new_n3725_1));
  not_8  g01377(.A(n442), .Y(new_n3726));
  nand_5 g01378(.A(n24638), .B(new_n3726), .Y(new_n3727));
  not_8  g01379(.A(n21674), .Y(new_n3728));
  nand_5 g01380(.A(new_n3728), .B(n9172), .Y(new_n3729));
  not_8  g01381(.A(n9172), .Y(new_n3730));
  nand_5 g01382(.A(n21674), .B(new_n3730), .Y(new_n3731));
  not_8  g01383(.A(n17251), .Y(new_n3732));
  nand_5 g01384(.A(new_n3732), .B(n4913), .Y(new_n3733_1));
  not_8  g01385(.A(n4913), .Y(new_n3734));
  nand_5 g01386(.A(n17251), .B(new_n3734), .Y(new_n3735));
  not_8  g01387(.A(n14790), .Y(new_n3736));
  nand_5 g01388(.A(new_n3736), .B(n604), .Y(new_n3737));
  not_8  g01389(.A(n604), .Y(new_n3738));
  nand_5 g01390(.A(n14790), .B(new_n3738), .Y(new_n3739));
  not_8  g01391(.A(n10096), .Y(new_n3740_1));
  nand_5 g01392(.A(n16824), .B(new_n3740_1), .Y(new_n3741));
  not_8  g01393(.A(n16824), .Y(new_n3742));
  nand_5 g01394(.A(new_n3742), .B(n10096), .Y(new_n3743));
  not_8  g01395(.A(n16994), .Y(new_n3744));
  nand_5 g01396(.A(new_n3744), .B(n16521), .Y(new_n3745));
  not_8  g01397(.A(n16521), .Y(new_n3746));
  nand_5 g01398(.A(n16994), .B(new_n3746), .Y(new_n3747));
  not_8  g01399(.A(n7139), .Y(new_n3748));
  nand_5 g01400(.A(n9246), .B(new_n3748), .Y(new_n3749));
  nand_5 g01401(.A(new_n3749), .B(new_n3747), .Y(new_n3750));
  nand_5 g01402(.A(new_n3750), .B(new_n3745), .Y(new_n3751));
  nand_5 g01403(.A(new_n3751), .B(new_n3743), .Y(new_n3752));
  nand_5 g01404(.A(new_n3752), .B(new_n3741), .Y(new_n3753));
  nand_5 g01405(.A(new_n3753), .B(new_n3739), .Y(new_n3754));
  nand_5 g01406(.A(new_n3754), .B(new_n3737), .Y(new_n3755_1));
  nand_5 g01407(.A(new_n3755_1), .B(new_n3735), .Y(new_n3756));
  nand_5 g01408(.A(new_n3756), .B(new_n3733_1), .Y(new_n3757));
  nand_5 g01409(.A(new_n3757), .B(new_n3731), .Y(new_n3758_1));
  nand_5 g01410(.A(new_n3758_1), .B(new_n3729), .Y(new_n3759));
  nand_5 g01411(.A(new_n3759), .B(new_n3727), .Y(new_n3760_1));
  nand_5 g01412(.A(new_n3760_1), .B(new_n3725_1), .Y(new_n3761));
  nand_5 g01413(.A(new_n3761), .B(new_n3723), .Y(new_n3762));
  nand_5 g01414(.A(new_n3762), .B(new_n3721), .Y(new_n3763));
  nand_5 g01415(.A(new_n3763), .B(new_n3719), .Y(new_n3764));
  nand_5 g01416(.A(new_n3764), .B(new_n3717), .Y(new_n3765));
  not_8  g01417(.A(new_n3765), .Y(new_n3766));
  xor_4  g01418(.A(new_n3766), .B(new_n3715), .Y(new_n3767));
  nand_5 g01419(.A(new_n3767), .B(new_n3710_1), .Y(new_n3768));
  not_8  g01420(.A(new_n3710_1), .Y(new_n3769));
  not_8  g01421(.A(new_n3767), .Y(new_n3770));
  nand_5 g01422(.A(new_n3770), .B(new_n3769), .Y(new_n3771));
  nand_5 g01423(.A(new_n3771), .B(new_n3768), .Y(new_n3772));
  xor_4  g01424(.A(new_n3705), .B(n21489), .Y(new_n3773));
  nand_5 g01425(.A(new_n3719), .B(new_n3717), .Y(new_n3774));
  xor_4  g01426(.A(new_n3774), .B(new_n3763), .Y(new_n3775));
  nand_5 g01427(.A(new_n3775), .B(new_n3773), .Y(new_n3776));
  or_5   g01428(.A(new_n3775), .B(new_n3773), .Y(new_n3777));
  not_8  g01429(.A(n20213), .Y(new_n3778));
  xor_4  g01430(.A(new_n3704), .B(new_n3778), .Y(new_n3779));
  nand_5 g01431(.A(new_n3723), .B(new_n3721), .Y(new_n3780));
  xor_4  g01432(.A(new_n3780), .B(new_n3761), .Y(new_n3781_1));
  nand_5 g01433(.A(new_n3781_1), .B(new_n3779), .Y(new_n3782));
  not_8  g01434(.A(new_n3779), .Y(new_n3783));
  not_8  g01435(.A(new_n3781_1), .Y(new_n3784));
  nand_5 g01436(.A(new_n3784), .B(new_n3783), .Y(new_n3785_1));
  xor_4  g01437(.A(new_n3703), .B(n13912), .Y(new_n3786));
  nand_5 g01438(.A(new_n3727), .B(new_n3725_1), .Y(new_n3787));
  xor_4  g01439(.A(new_n3787), .B(new_n3759), .Y(new_n3788));
  nand_5 g01440(.A(new_n3788), .B(new_n3786), .Y(new_n3789));
  not_8  g01441(.A(new_n3786), .Y(new_n3790));
  not_8  g01442(.A(new_n3788), .Y(new_n3791));
  nand_5 g01443(.A(new_n3791), .B(new_n3790), .Y(new_n3792));
  not_8  g01444(.A(n7670), .Y(new_n3793));
  xor_4  g01445(.A(new_n3702), .B(new_n3793), .Y(new_n3794_1));
  nand_5 g01446(.A(new_n3731), .B(new_n3729), .Y(new_n3795_1));
  xor_4  g01447(.A(new_n3795_1), .B(new_n3757), .Y(new_n3796));
  nand_5 g01448(.A(new_n3796), .B(new_n3794_1), .Y(new_n3797));
  or_5   g01449(.A(new_n3796), .B(new_n3794_1), .Y(new_n3798));
  xor_4  g01450(.A(new_n3701), .B(new_n3696), .Y(new_n3799));
  not_8  g01451(.A(new_n3799), .Y(new_n3800));
  nand_5 g01452(.A(new_n3735), .B(new_n3733_1), .Y(new_n3801));
  xor_4  g01453(.A(new_n3801), .B(new_n3755_1), .Y(new_n3802));
  nand_5 g01454(.A(new_n3802), .B(new_n3800), .Y(new_n3803));
  or_5   g01455(.A(new_n3802), .B(new_n3800), .Y(new_n3804));
  xor_4  g01456(.A(new_n3700), .B(n22290), .Y(new_n3805));
  not_8  g01457(.A(new_n3805), .Y(new_n3806));
  nand_5 g01458(.A(new_n3739), .B(new_n3737), .Y(new_n3807));
  xor_4  g01459(.A(new_n3807), .B(new_n3753), .Y(new_n3808));
  nand_5 g01460(.A(new_n3808), .B(new_n3806), .Y(new_n3809));
  or_5   g01461(.A(new_n3808), .B(new_n3806), .Y(new_n3810));
  nand_5 g01462(.A(new_n3699), .B(n11273), .Y(new_n3811));
  and_5  g01463(.A(new_n3811), .B(new_n3700), .Y(new_n3812));
  not_8  g01464(.A(new_n3812), .Y(new_n3813));
  nand_5 g01465(.A(new_n3743), .B(new_n3741), .Y(new_n3814));
  xor_4  g01466(.A(new_n3814), .B(new_n3751), .Y(new_n3815));
  nand_5 g01467(.A(new_n3815), .B(new_n3813), .Y(new_n3816));
  nor_5  g01468(.A(new_n3815), .B(new_n3813), .Y(new_n3817));
  not_8  g01469(.A(new_n3817), .Y(new_n3818));
  nand_5 g01470(.A(n25565), .B(n21993), .Y(new_n3819));
  and_5  g01471(.A(new_n3819), .B(new_n3699), .Y(new_n3820));
  not_8  g01472(.A(new_n3820), .Y(new_n3821));
  and_5  g01473(.A(new_n3747), .B(new_n3745), .Y(new_n3822));
  xor_4  g01474(.A(new_n3822), .B(new_n3749), .Y(new_n3823));
  not_8  g01475(.A(new_n3823), .Y(new_n3824));
  nand_5 g01476(.A(new_n3824), .B(new_n3821), .Y(new_n3825));
  nand_5 g01477(.A(new_n3823), .B(new_n3820), .Y(new_n3826));
  not_8  g01478(.A(n9246), .Y(new_n3827));
  nand_5 g01479(.A(new_n3827), .B(n7139), .Y(new_n3828_1));
  and_5  g01480(.A(new_n3828_1), .B(new_n3749), .Y(new_n3829));
  not_8  g01481(.A(new_n3829), .Y(new_n3830));
  nand_5 g01482(.A(new_n3830), .B(n21993), .Y(new_n3831));
  nand_5 g01483(.A(new_n3831), .B(new_n3826), .Y(new_n3832));
  nand_5 g01484(.A(new_n3832), .B(new_n3825), .Y(new_n3833));
  nand_5 g01485(.A(new_n3833), .B(new_n3818), .Y(new_n3834));
  nand_5 g01486(.A(new_n3834), .B(new_n3816), .Y(new_n3835));
  nand_5 g01487(.A(new_n3835), .B(new_n3810), .Y(new_n3836));
  nand_5 g01488(.A(new_n3836), .B(new_n3809), .Y(new_n3837));
  nand_5 g01489(.A(new_n3837), .B(new_n3804), .Y(new_n3838));
  nand_5 g01490(.A(new_n3838), .B(new_n3803), .Y(new_n3839));
  nand_5 g01491(.A(new_n3839), .B(new_n3798), .Y(new_n3840));
  nand_5 g01492(.A(new_n3840), .B(new_n3797), .Y(new_n3841));
  nand_5 g01493(.A(new_n3841), .B(new_n3792), .Y(new_n3842_1));
  nand_5 g01494(.A(new_n3842_1), .B(new_n3789), .Y(new_n3843));
  nand_5 g01495(.A(new_n3843), .B(new_n3785_1), .Y(new_n3844));
  nand_5 g01496(.A(new_n3844), .B(new_n3782), .Y(new_n3845));
  nand_5 g01497(.A(new_n3845), .B(new_n3777), .Y(new_n3846));
  nand_5 g01498(.A(new_n3846), .B(new_n3776), .Y(new_n3847));
  xor_4  g01499(.A(new_n3847), .B(new_n3772), .Y(new_n3848));
  not_8  g01500(.A(n14130), .Y(new_n3849));
  not_8  g01501(.A(n9251), .Y(new_n3850_1));
  nand_5 g01502(.A(new_n2502), .B(new_n3850_1), .Y(new_n3851));
  or_5   g01503(.A(new_n3851), .B(n6385), .Y(new_n3852));
  nor_5  g01504(.A(new_n3852), .B(n3136), .Y(new_n3853));
  nand_5 g01505(.A(new_n3853), .B(new_n2490), .Y(new_n3854));
  nor_5  g01506(.A(new_n3854), .B(n25643), .Y(new_n3855));
  nand_5 g01507(.A(new_n3855), .B(new_n2599), .Y(new_n3856));
  nor_5  g01508(.A(new_n3856), .B(n16482), .Y(new_n3857));
  nand_5 g01509(.A(new_n3857), .B(new_n3849), .Y(new_n3858));
  not_8  g01510(.A(new_n3858), .Y(new_n3859));
  nor_5  g01511(.A(new_n3857), .B(new_n3849), .Y(new_n3860));
  nor_5  g01512(.A(new_n3860), .B(new_n3859), .Y(new_n3861));
  or_5   g01513(.A(new_n3861), .B(n10117), .Y(new_n3862));
  nand_5 g01514(.A(new_n3861), .B(n10117), .Y(new_n3863));
  xor_4  g01515(.A(new_n3856), .B(n16482), .Y(new_n3864));
  or_5   g01516(.A(new_n3864), .B(n13460), .Y(new_n3865));
  nand_5 g01517(.A(new_n3864), .B(n13460), .Y(new_n3866));
  xor_4  g01518(.A(new_n3855), .B(new_n2599), .Y(new_n3867));
  or_5   g01519(.A(new_n3867), .B(n6104), .Y(new_n3868));
  nand_5 g01520(.A(new_n3867), .B(n6104), .Y(new_n3869_1));
  xor_4  g01521(.A(new_n3854), .B(n25643), .Y(new_n3870));
  or_5   g01522(.A(new_n3870), .B(n4119), .Y(new_n3871_1));
  nand_5 g01523(.A(new_n3870), .B(n4119), .Y(new_n3872));
  xor_4  g01524(.A(new_n3853), .B(new_n2490), .Y(new_n3873));
  or_5   g01525(.A(new_n3873), .B(n14510), .Y(new_n3874));
  nand_5 g01526(.A(new_n3873), .B(n14510), .Y(new_n3875));
  xor_4  g01527(.A(new_n3852), .B(n3136), .Y(new_n3876));
  or_5   g01528(.A(new_n3876), .B(n13263), .Y(new_n3877));
  nand_5 g01529(.A(new_n3876), .B(n13263), .Y(new_n3878));
  nand_5 g01530(.A(new_n3851), .B(n6385), .Y(new_n3879));
  and_5  g01531(.A(new_n3879), .B(new_n3852), .Y(new_n3880));
  or_5   g01532(.A(new_n3880), .B(n20455), .Y(new_n3881));
  nand_5 g01533(.A(new_n3880), .B(n20455), .Y(new_n3882));
  nand_5 g01534(.A(n20138), .B(n9251), .Y(new_n3883));
  and_5  g01535(.A(new_n3883), .B(new_n3851), .Y(new_n3884));
  or_5   g01536(.A(new_n3884), .B(n1639), .Y(new_n3885));
  nand_5 g01537(.A(n16968), .B(n9251), .Y(new_n3886));
  nand_5 g01538(.A(new_n3884), .B(n1639), .Y(new_n3887));
  nand_5 g01539(.A(new_n3887), .B(new_n3886), .Y(new_n3888));
  nand_5 g01540(.A(new_n3888), .B(new_n3885), .Y(new_n3889));
  nand_5 g01541(.A(new_n3889), .B(new_n3882), .Y(new_n3890));
  nand_5 g01542(.A(new_n3890), .B(new_n3881), .Y(new_n3891_1));
  nand_5 g01543(.A(new_n3891_1), .B(new_n3878), .Y(new_n3892));
  nand_5 g01544(.A(new_n3892), .B(new_n3877), .Y(new_n3893));
  nand_5 g01545(.A(new_n3893), .B(new_n3875), .Y(new_n3894));
  nand_5 g01546(.A(new_n3894), .B(new_n3874), .Y(new_n3895));
  nand_5 g01547(.A(new_n3895), .B(new_n3872), .Y(new_n3896));
  nand_5 g01548(.A(new_n3896), .B(new_n3871_1), .Y(new_n3897));
  nand_5 g01549(.A(new_n3897), .B(new_n3869_1), .Y(new_n3898));
  nand_5 g01550(.A(new_n3898), .B(new_n3868), .Y(new_n3899));
  nand_5 g01551(.A(new_n3899), .B(new_n3866), .Y(new_n3900));
  nand_5 g01552(.A(new_n3900), .B(new_n3865), .Y(new_n3901));
  nand_5 g01553(.A(new_n3901), .B(new_n3863), .Y(new_n3902));
  nand_5 g01554(.A(new_n3902), .B(new_n3862), .Y(new_n3903));
  xor_4  g01555(.A(new_n3858), .B(n8856), .Y(new_n3904));
  xor_4  g01556(.A(new_n3904), .B(n25494), .Y(new_n3905));
  xor_4  g01557(.A(new_n3905), .B(new_n3903), .Y(new_n3906));
  not_8  g01558(.A(new_n3906), .Y(new_n3907));
  nand_5 g01559(.A(new_n3907), .B(n26180), .Y(new_n3908));
  not_8  g01560(.A(n26180), .Y(new_n3909_1));
  nand_5 g01561(.A(new_n3906), .B(new_n3909_1), .Y(new_n3910));
  nand_5 g01562(.A(new_n3910), .B(new_n3908), .Y(new_n3911));
  nand_5 g01563(.A(new_n3863), .B(new_n3862), .Y(new_n3912));
  xor_4  g01564(.A(new_n3912), .B(new_n3901), .Y(new_n3913));
  nand_5 g01565(.A(new_n3913), .B(n24004), .Y(new_n3914));
  not_8  g01566(.A(n24004), .Y(new_n3915));
  not_8  g01567(.A(new_n3913), .Y(new_n3916));
  nand_5 g01568(.A(new_n3916), .B(new_n3915), .Y(new_n3917));
  nand_5 g01569(.A(new_n3866), .B(new_n3865), .Y(new_n3918_1));
  xor_4  g01570(.A(new_n3918_1), .B(new_n3899), .Y(new_n3919));
  nand_5 g01571(.A(new_n3919), .B(n12871), .Y(new_n3920));
  not_8  g01572(.A(n12871), .Y(new_n3921));
  not_8  g01573(.A(new_n3919), .Y(new_n3922));
  nand_5 g01574(.A(new_n3922), .B(new_n3921), .Y(new_n3923));
  nand_5 g01575(.A(new_n3869_1), .B(new_n3868), .Y(new_n3924));
  xor_4  g01576(.A(new_n3924), .B(new_n3897), .Y(new_n3925_1));
  nand_5 g01577(.A(new_n3925_1), .B(n23304), .Y(new_n3926));
  not_8  g01578(.A(n23304), .Y(new_n3927));
  not_8  g01579(.A(new_n3925_1), .Y(new_n3928));
  nand_5 g01580(.A(new_n3928), .B(new_n3927), .Y(new_n3929));
  nand_5 g01581(.A(new_n3872), .B(new_n3871_1), .Y(new_n3930));
  xor_4  g01582(.A(new_n3930), .B(new_n3895), .Y(new_n3931));
  nand_5 g01583(.A(new_n3931), .B(n19361), .Y(new_n3932_1));
  not_8  g01584(.A(n19361), .Y(new_n3933));
  not_8  g01585(.A(new_n3931), .Y(new_n3934_1));
  nand_5 g01586(.A(new_n3934_1), .B(new_n3933), .Y(new_n3935));
  nand_5 g01587(.A(new_n3875), .B(new_n3874), .Y(new_n3936));
  xor_4  g01588(.A(new_n3936), .B(new_n3893), .Y(new_n3937));
  nand_5 g01589(.A(new_n3937), .B(n1437), .Y(new_n3938));
  not_8  g01590(.A(n1437), .Y(new_n3939));
  not_8  g01591(.A(new_n3937), .Y(new_n3940));
  nand_5 g01592(.A(new_n3940), .B(new_n3939), .Y(new_n3941));
  nand_5 g01593(.A(new_n3878), .B(new_n3877), .Y(new_n3942));
  xor_4  g01594(.A(new_n3942), .B(new_n3891_1), .Y(new_n3943));
  nand_5 g01595(.A(new_n3943), .B(n4722), .Y(new_n3944));
  not_8  g01596(.A(n4722), .Y(new_n3945_1));
  not_8  g01597(.A(new_n3943), .Y(new_n3946));
  nand_5 g01598(.A(new_n3946), .B(new_n3945_1), .Y(new_n3947));
  nand_5 g01599(.A(new_n3882), .B(new_n3881), .Y(new_n3948));
  xor_4  g01600(.A(new_n3948), .B(new_n3889), .Y(new_n3949));
  nand_5 g01601(.A(new_n3949), .B(n14633), .Y(new_n3950));
  not_8  g01602(.A(n14633), .Y(new_n3951));
  not_8  g01603(.A(new_n3949), .Y(new_n3952_1));
  nand_5 g01604(.A(new_n3952_1), .B(new_n3951), .Y(new_n3953));
  nand_5 g01605(.A(new_n3887), .B(new_n3885), .Y(new_n3954));
  xor_4  g01606(.A(new_n3954), .B(new_n3886), .Y(new_n3955));
  nand_5 g01607(.A(new_n3955), .B(n8721), .Y(new_n3956));
  not_8  g01608(.A(n8721), .Y(new_n3957));
  not_8  g01609(.A(new_n3955), .Y(new_n3958));
  nand_5 g01610(.A(new_n3958), .B(new_n3957), .Y(new_n3959_1));
  not_8  g01611(.A(n16968), .Y(new_n3960));
  nand_5 g01612(.A(new_n3960), .B(new_n3850_1), .Y(new_n3961));
  and_5  g01613(.A(new_n3961), .B(new_n3886), .Y(new_n3962_1));
  nand_5 g01614(.A(new_n3962_1), .B(n18578), .Y(new_n3963));
  not_8  g01615(.A(new_n3963), .Y(new_n3964));
  nand_5 g01616(.A(new_n3964), .B(new_n3959_1), .Y(new_n3965));
  nand_5 g01617(.A(new_n3965), .B(new_n3956), .Y(new_n3966));
  nand_5 g01618(.A(new_n3966), .B(new_n3953), .Y(new_n3967));
  nand_5 g01619(.A(new_n3967), .B(new_n3950), .Y(new_n3968));
  nand_5 g01620(.A(new_n3968), .B(new_n3947), .Y(new_n3969));
  nand_5 g01621(.A(new_n3969), .B(new_n3944), .Y(new_n3970));
  nand_5 g01622(.A(new_n3970), .B(new_n3941), .Y(new_n3971_1));
  nand_5 g01623(.A(new_n3971_1), .B(new_n3938), .Y(new_n3972));
  nand_5 g01624(.A(new_n3972), .B(new_n3935), .Y(new_n3973));
  nand_5 g01625(.A(new_n3973), .B(new_n3932_1), .Y(new_n3974));
  nand_5 g01626(.A(new_n3974), .B(new_n3929), .Y(new_n3975));
  nand_5 g01627(.A(new_n3975), .B(new_n3926), .Y(new_n3976));
  nand_5 g01628(.A(new_n3976), .B(new_n3923), .Y(new_n3977));
  nand_5 g01629(.A(new_n3977), .B(new_n3920), .Y(new_n3978));
  nand_5 g01630(.A(new_n3978), .B(new_n3917), .Y(new_n3979));
  nand_5 g01631(.A(new_n3979), .B(new_n3914), .Y(new_n3980));
  xor_4  g01632(.A(new_n3980), .B(new_n3911), .Y(new_n3981));
  not_8  g01633(.A(new_n3981), .Y(new_n3982));
  nand_5 g01634(.A(new_n3982), .B(new_n3848), .Y(new_n3983_1));
  or_5   g01635(.A(new_n3982), .B(new_n3848), .Y(new_n3984_1));
  nand_5 g01636(.A(new_n3984_1), .B(new_n3983_1), .Y(new_n3985));
  nand_5 g01637(.A(new_n3914), .B(new_n3917), .Y(new_n3986));
  xor_4  g01638(.A(new_n3986), .B(new_n3978), .Y(new_n3987));
  not_8  g01639(.A(new_n3987), .Y(new_n3988));
  nand_5 g01640(.A(new_n3777), .B(new_n3776), .Y(new_n3989));
  xor_4  g01641(.A(new_n3989), .B(new_n3845), .Y(new_n3990));
  nand_5 g01642(.A(new_n3990), .B(new_n3988), .Y(new_n3991));
  or_5   g01643(.A(new_n3990), .B(new_n3988), .Y(new_n3992));
  nand_5 g01644(.A(new_n3785_1), .B(new_n3782), .Y(new_n3993));
  xor_4  g01645(.A(new_n3993), .B(new_n3843), .Y(new_n3994));
  nand_5 g01646(.A(new_n3920), .B(new_n3923), .Y(new_n3995));
  xor_4  g01647(.A(new_n3995), .B(new_n3976), .Y(new_n3996));
  not_8  g01648(.A(new_n3996), .Y(new_n3997));
  nand_5 g01649(.A(new_n3997), .B(new_n3994), .Y(new_n3998));
  or_5   g01650(.A(new_n3997), .B(new_n3994), .Y(new_n3999));
  nand_5 g01651(.A(new_n3926), .B(new_n3929), .Y(new_n4000_1));
  xor_4  g01652(.A(new_n4000_1), .B(new_n3974), .Y(new_n4001));
  not_8  g01653(.A(new_n4001), .Y(new_n4002));
  nand_5 g01654(.A(new_n3792), .B(new_n3789), .Y(new_n4003));
  xor_4  g01655(.A(new_n4003), .B(new_n3841), .Y(new_n4004));
  nand_5 g01656(.A(new_n4004), .B(new_n4002), .Y(new_n4005));
  or_5   g01657(.A(new_n4004), .B(new_n4002), .Y(new_n4006));
  nand_5 g01658(.A(new_n3932_1), .B(new_n3935), .Y(new_n4007));
  xor_4  g01659(.A(new_n4007), .B(new_n3972), .Y(new_n4008));
  not_8  g01660(.A(new_n4008), .Y(new_n4009));
  nand_5 g01661(.A(new_n3798), .B(new_n3797), .Y(new_n4010_1));
  xor_4  g01662(.A(new_n4010_1), .B(new_n3839), .Y(new_n4011));
  nand_5 g01663(.A(new_n4011), .B(new_n4009), .Y(new_n4012));
  or_5   g01664(.A(new_n4011), .B(new_n4009), .Y(new_n4013));
  nand_5 g01665(.A(new_n3804), .B(new_n3803), .Y(new_n4014_1));
  xor_4  g01666(.A(new_n4014_1), .B(new_n3837), .Y(new_n4015));
  nand_5 g01667(.A(new_n3938), .B(new_n3941), .Y(new_n4016));
  xor_4  g01668(.A(new_n4016), .B(new_n3970), .Y(new_n4017));
  not_8  g01669(.A(new_n4017), .Y(new_n4018));
  nand_5 g01670(.A(new_n4018), .B(new_n4015), .Y(new_n4019));
  or_5   g01671(.A(new_n4018), .B(new_n4015), .Y(new_n4020));
  nand_5 g01672(.A(new_n3810), .B(new_n3809), .Y(new_n4021));
  xor_4  g01673(.A(new_n4021), .B(new_n3835), .Y(new_n4022));
  nand_5 g01674(.A(new_n3944), .B(new_n3947), .Y(new_n4023));
  xor_4  g01675(.A(new_n4023), .B(new_n3968), .Y(new_n4024));
  not_8  g01676(.A(new_n4024), .Y(new_n4025));
  nand_5 g01677(.A(new_n4025), .B(new_n4022), .Y(new_n4026));
  or_5   g01678(.A(new_n4025), .B(new_n4022), .Y(new_n4027));
  nand_5 g01679(.A(new_n3950), .B(new_n3953), .Y(new_n4028));
  xor_4  g01680(.A(new_n4028), .B(new_n3966), .Y(new_n4029));
  not_8  g01681(.A(new_n4029), .Y(new_n4030));
  nand_5 g01682(.A(new_n3818), .B(new_n3816), .Y(new_n4031));
  xor_4  g01683(.A(new_n4031), .B(new_n3833), .Y(new_n4032));
  nand_5 g01684(.A(new_n4032), .B(new_n4030), .Y(new_n4033));
  or_5   g01685(.A(new_n4032), .B(new_n4030), .Y(new_n4034));
  nand_5 g01686(.A(new_n3826), .B(new_n3825), .Y(new_n4035));
  xor_4  g01687(.A(new_n4035), .B(new_n3831), .Y(new_n4036));
  nand_5 g01688(.A(new_n3956), .B(new_n3959_1), .Y(new_n4037));
  xor_4  g01689(.A(new_n4037), .B(new_n3964), .Y(new_n4038));
  not_8  g01690(.A(new_n4038), .Y(new_n4039));
  nand_5 g01691(.A(new_n4039), .B(new_n4036), .Y(new_n4040));
  or_5   g01692(.A(new_n4039), .B(new_n4036), .Y(new_n4041));
  or_5   g01693(.A(new_n3962_1), .B(n18578), .Y(new_n4042));
  nand_5 g01694(.A(new_n4042), .B(new_n3963), .Y(new_n4043));
  nand_5 g01695(.A(new_n3829), .B(new_n3697), .Y(new_n4044));
  nand_5 g01696(.A(new_n4044), .B(new_n3831), .Y(new_n4045));
  nor_5  g01697(.A(new_n4045), .B(new_n4043), .Y(new_n4046));
  nand_5 g01698(.A(new_n4046), .B(new_n4041), .Y(new_n4047));
  nand_5 g01699(.A(new_n4047), .B(new_n4040), .Y(new_n4048));
  nand_5 g01700(.A(new_n4048), .B(new_n4034), .Y(new_n4049));
  nand_5 g01701(.A(new_n4049), .B(new_n4033), .Y(new_n4050));
  nand_5 g01702(.A(new_n4050), .B(new_n4027), .Y(new_n4051));
  nand_5 g01703(.A(new_n4051), .B(new_n4026), .Y(new_n4052));
  nand_5 g01704(.A(new_n4052), .B(new_n4020), .Y(new_n4053));
  nand_5 g01705(.A(new_n4053), .B(new_n4019), .Y(new_n4054));
  nand_5 g01706(.A(new_n4054), .B(new_n4013), .Y(new_n4055));
  nand_5 g01707(.A(new_n4055), .B(new_n4012), .Y(new_n4056));
  nand_5 g01708(.A(new_n4056), .B(new_n4006), .Y(new_n4057));
  nand_5 g01709(.A(new_n4057), .B(new_n4005), .Y(new_n4058));
  nand_5 g01710(.A(new_n4058), .B(new_n3999), .Y(new_n4059));
  nand_5 g01711(.A(new_n4059), .B(new_n3998), .Y(new_n4060));
  nand_5 g01712(.A(new_n4060), .B(new_n3992), .Y(new_n4061));
  nand_5 g01713(.A(new_n4061), .B(new_n3991), .Y(new_n4062));
  xnor_4 g01714(.A(new_n4062), .B(new_n3985), .Y(n235));
  nand_5 g01715(.A(n19911), .B(new_n3084), .Y(new_n4064));
  nand_5 g01716(.A(new_n2402), .B(n10053), .Y(new_n4065));
  nand_5 g01717(.A(n13708), .B(new_n3085), .Y(new_n4066));
  nand_5 g01718(.A(new_n2393), .B(n8399), .Y(new_n4067));
  nand_5 g01719(.A(n18409), .B(new_n3090), .Y(new_n4068));
  nand_5 g01720(.A(new_n2384), .B(n9507), .Y(new_n4069));
  nand_5 g01721(.A(n26979), .B(new_n2377), .Y(new_n4070));
  nand_5 g01722(.A(new_n4070), .B(new_n4069), .Y(new_n4071_1));
  nand_5 g01723(.A(new_n4071_1), .B(new_n4068), .Y(new_n4072));
  nand_5 g01724(.A(new_n4072), .B(new_n4067), .Y(new_n4073));
  nand_5 g01725(.A(new_n4073), .B(new_n4066), .Y(new_n4074));
  nand_5 g01726(.A(new_n4074), .B(new_n4065), .Y(new_n4075));
  nand_5 g01727(.A(new_n4075), .B(new_n4064), .Y(new_n4076));
  nand_5 g01728(.A(new_n3079), .B(n2731), .Y(new_n4077));
  nand_5 g01729(.A(n19514), .B(new_n2411), .Y(new_n4078));
  nand_5 g01730(.A(new_n4078), .B(new_n4077), .Y(new_n4079));
  xor_4  g01731(.A(new_n4079), .B(new_n4076), .Y(new_n4080));
  not_8  g01732(.A(new_n4080), .Y(new_n4081));
  not_8  g01733(.A(n626), .Y(new_n4082));
  not_8  g01734(.A(n19618), .Y(new_n4083));
  not_8  g01735(.A(n12121), .Y(new_n4084));
  not_8  g01736(.A(n22043), .Y(new_n4085_1));
  nand_5 g01737(.A(new_n4085_1), .B(new_n4084), .Y(new_n4086));
  not_8  g01738(.A(new_n4086), .Y(new_n4087));
  nand_5 g01739(.A(new_n4087), .B(new_n4083), .Y(new_n4088_1));
  nor_5  g01740(.A(new_n4088_1), .B(n1204), .Y(new_n4089_1));
  nand_5 g01741(.A(new_n4089_1), .B(new_n4082), .Y(new_n4090));
  not_8  g01742(.A(new_n4090), .Y(new_n4091));
  nor_5  g01743(.A(new_n4089_1), .B(new_n4082), .Y(new_n4092));
  nor_5  g01744(.A(new_n4092), .B(new_n4091), .Y(new_n4093));
  or_5   g01745(.A(new_n4093), .B(new_n4081), .Y(new_n4094));
  nand_5 g01746(.A(new_n4093), .B(new_n4081), .Y(new_n4095));
  nand_5 g01747(.A(new_n4065), .B(new_n4064), .Y(new_n4096));
  xor_4  g01748(.A(new_n4096), .B(new_n4074), .Y(new_n4097));
  not_8  g01749(.A(n1204), .Y(new_n4098));
  xor_4  g01750(.A(new_n4088_1), .B(new_n4098), .Y(new_n4099));
  nand_5 g01751(.A(new_n4099), .B(new_n4097), .Y(new_n4100_1));
  nor_5  g01752(.A(new_n4099), .B(new_n4097), .Y(new_n4101));
  not_8  g01753(.A(new_n4101), .Y(new_n4102));
  and_5  g01754(.A(new_n4069), .B(new_n4068), .Y(new_n4103_1));
  xor_4  g01755(.A(new_n4103_1), .B(new_n4070), .Y(new_n4104));
  not_8  g01756(.A(new_n4104), .Y(new_n4105));
  nand_5 g01757(.A(n22043), .B(n12121), .Y(new_n4106));
  nand_5 g01758(.A(new_n4106), .B(new_n4086), .Y(new_n4107));
  nand_5 g01759(.A(new_n4107), .B(new_n4105), .Y(new_n4108));
  nor_5  g01760(.A(new_n4107), .B(new_n4105), .Y(new_n4109));
  not_8  g01761(.A(new_n4109), .Y(new_n4110));
  nand_5 g01762(.A(new_n3164_1), .B(n5704), .Y(new_n4111));
  and_5  g01763(.A(new_n4111), .B(new_n4070), .Y(new_n4112));
  not_8  g01764(.A(new_n4112), .Y(new_n4113));
  nand_5 g01765(.A(new_n4113), .B(n12121), .Y(new_n4114));
  nand_5 g01766(.A(new_n4114), .B(new_n4110), .Y(new_n4115));
  nand_5 g01767(.A(new_n4115), .B(new_n4108), .Y(new_n4116));
  nand_5 g01768(.A(new_n4067), .B(new_n4066), .Y(new_n4117));
  xor_4  g01769(.A(new_n4117), .B(new_n4072), .Y(new_n4118));
  not_8  g01770(.A(new_n4118), .Y(new_n4119_1));
  xor_4  g01771(.A(new_n4086), .B(n19618), .Y(new_n4120));
  nand_5 g01772(.A(new_n4120), .B(new_n4119_1), .Y(new_n4121));
  nand_5 g01773(.A(new_n4121), .B(new_n4116), .Y(new_n4122));
  nor_5  g01774(.A(new_n4120), .B(new_n4119_1), .Y(new_n4123_1));
  not_8  g01775(.A(new_n4123_1), .Y(new_n4124));
  nand_5 g01776(.A(new_n4124), .B(new_n4122), .Y(new_n4125));
  nand_5 g01777(.A(new_n4125), .B(new_n4102), .Y(new_n4126));
  nand_5 g01778(.A(new_n4126), .B(new_n4100_1), .Y(new_n4127));
  nand_5 g01779(.A(new_n4127), .B(new_n4095), .Y(new_n4128));
  nand_5 g01780(.A(new_n4128), .B(new_n4094), .Y(new_n4129));
  nand_5 g01781(.A(new_n4078), .B(new_n4076), .Y(new_n4130));
  nand_5 g01782(.A(new_n4130), .B(new_n4077), .Y(new_n4131));
  nand_5 g01783(.A(new_n3073), .B(n18907), .Y(new_n4132));
  nand_5 g01784(.A(n23068), .B(new_n2474), .Y(new_n4133));
  nand_5 g01785(.A(new_n4133), .B(new_n4132), .Y(new_n4134_1));
  xor_4  g01786(.A(new_n4134_1), .B(new_n4131), .Y(new_n4135));
  not_8  g01787(.A(new_n4135), .Y(new_n4136));
  not_8  g01788(.A(n5337), .Y(new_n4137));
  nand_5 g01789(.A(new_n4091), .B(new_n4137), .Y(new_n4138));
  not_8  g01790(.A(new_n4138), .Y(new_n4139));
  nor_5  g01791(.A(new_n4091), .B(new_n4137), .Y(new_n4140));
  nor_5  g01792(.A(new_n4140), .B(new_n4139), .Y(new_n4141));
  or_5   g01793(.A(new_n4141), .B(new_n4136), .Y(new_n4142));
  nand_5 g01794(.A(new_n4141), .B(new_n4136), .Y(new_n4143));
  nand_5 g01795(.A(new_n4143), .B(new_n4142), .Y(new_n4144));
  xor_4  g01796(.A(new_n4144), .B(new_n4129), .Y(new_n4145));
  not_8  g01797(.A(n342), .Y(new_n4146_1));
  not_8  g01798(.A(n15967), .Y(new_n4147));
  not_8  g01799(.A(n13319), .Y(new_n4148));
  not_8  g01800(.A(n25435), .Y(new_n4149));
  nand_5 g01801(.A(new_n4149), .B(new_n4148), .Y(new_n4150_1));
  not_8  g01802(.A(new_n4150_1), .Y(new_n4151_1));
  nand_5 g01803(.A(new_n4151_1), .B(new_n4147), .Y(new_n4152_1));
  nor_5  g01804(.A(new_n4152_1), .B(n25797), .Y(new_n4153_1));
  not_8  g01805(.A(new_n4153_1), .Y(new_n4154));
  nand_5 g01806(.A(new_n4152_1), .B(n25797), .Y(new_n4155));
  and_5  g01807(.A(new_n4155), .B(new_n4154), .Y(new_n4156));
  not_8  g01808(.A(new_n4156), .Y(new_n4157));
  nand_5 g01809(.A(new_n4157), .B(new_n4146_1), .Y(new_n4158));
  nand_5 g01810(.A(new_n4156), .B(n342), .Y(new_n4159));
  not_8  g01811(.A(n26553), .Y(new_n4160));
  nand_5 g01812(.A(new_n4150_1), .B(n15967), .Y(new_n4161));
  and_5  g01813(.A(new_n4161), .B(new_n4152_1), .Y(new_n4162));
  not_8  g01814(.A(new_n4162), .Y(new_n4163));
  nand_5 g01815(.A(new_n4163), .B(new_n4160), .Y(new_n4164));
  nand_5 g01816(.A(new_n4162), .B(n26553), .Y(new_n4165_1));
  nand_5 g01817(.A(n25435), .B(n13319), .Y(new_n4166));
  and_5  g01818(.A(new_n4166), .B(new_n4150_1), .Y(new_n4167));
  or_5   g01819(.A(new_n4167), .B(n4964), .Y(new_n4168));
  nand_5 g01820(.A(new_n4167), .B(n4964), .Y(new_n4169));
  nand_5 g01821(.A(n25435), .B(n7876), .Y(new_n4170));
  nand_5 g01822(.A(new_n4170), .B(new_n4169), .Y(new_n4171));
  nand_5 g01823(.A(new_n4171), .B(new_n4168), .Y(new_n4172_1));
  nand_5 g01824(.A(new_n4172_1), .B(new_n4165_1), .Y(new_n4173_1));
  nand_5 g01825(.A(new_n4173_1), .B(new_n4164), .Y(new_n4174));
  nand_5 g01826(.A(new_n4174), .B(new_n4159), .Y(new_n4175));
  nand_5 g01827(.A(new_n4175), .B(new_n4158), .Y(new_n4176_1));
  not_8  g01828(.A(n26107), .Y(new_n4177));
  not_8  g01829(.A(n6369), .Y(new_n4178));
  nand_5 g01830(.A(new_n4153_1), .B(new_n4178), .Y(new_n4179));
  nand_5 g01831(.A(new_n4154), .B(n6369), .Y(new_n4180));
  and_5  g01832(.A(new_n4180), .B(new_n4179), .Y(new_n4181));
  not_8  g01833(.A(new_n4181), .Y(new_n4182));
  nand_5 g01834(.A(new_n4182), .B(new_n4177), .Y(new_n4183));
  nand_5 g01835(.A(new_n4181), .B(n26107), .Y(new_n4184));
  nand_5 g01836(.A(new_n4184), .B(new_n4183), .Y(new_n4185));
  xor_4  g01837(.A(new_n4185), .B(new_n4176_1), .Y(new_n4186_1));
  or_5   g01838(.A(new_n4186_1), .B(n9003), .Y(new_n4187));
  nand_5 g01839(.A(new_n4186_1), .B(n9003), .Y(new_n4188));
  not_8  g01840(.A(n4957), .Y(new_n4189));
  nand_5 g01841(.A(new_n4159), .B(new_n4158), .Y(new_n4190));
  xor_4  g01842(.A(new_n4190), .B(new_n4174), .Y(new_n4191));
  not_8  g01843(.A(new_n4191), .Y(new_n4192));
  nand_5 g01844(.A(new_n4192), .B(new_n4189), .Y(new_n4193));
  nand_5 g01845(.A(new_n4191), .B(n4957), .Y(new_n4194));
  not_8  g01846(.A(n7524), .Y(new_n4195));
  nand_5 g01847(.A(new_n4165_1), .B(new_n4164), .Y(new_n4196));
  xor_4  g01848(.A(new_n4196), .B(new_n4172_1), .Y(new_n4197));
  not_8  g01849(.A(new_n4197), .Y(new_n4198));
  nand_5 g01850(.A(new_n4198), .B(new_n4195), .Y(new_n4199));
  nand_5 g01851(.A(new_n4197), .B(n7524), .Y(new_n4200));
  not_8  g01852(.A(n15743), .Y(new_n4201));
  nand_5 g01853(.A(new_n4169), .B(new_n4168), .Y(new_n4202));
  xor_4  g01854(.A(new_n4202), .B(new_n4170), .Y(new_n4203));
  not_8  g01855(.A(new_n4203), .Y(new_n4204_1));
  nand_5 g01856(.A(new_n4204_1), .B(new_n4201), .Y(new_n4205_1));
  nand_5 g01857(.A(new_n4203), .B(n15743), .Y(new_n4206));
  not_8  g01858(.A(n7876), .Y(new_n4207));
  nand_5 g01859(.A(new_n4149), .B(new_n4207), .Y(new_n4208));
  and_5  g01860(.A(new_n4208), .B(new_n4170), .Y(new_n4209));
  nand_5 g01861(.A(new_n4209), .B(n20658), .Y(new_n4210));
  nand_5 g01862(.A(new_n4210), .B(new_n4206), .Y(new_n4211));
  nand_5 g01863(.A(new_n4211), .B(new_n4205_1), .Y(new_n4212));
  nand_5 g01864(.A(new_n4212), .B(new_n4200), .Y(new_n4213));
  nand_5 g01865(.A(new_n4213), .B(new_n4199), .Y(new_n4214));
  nand_5 g01866(.A(new_n4214), .B(new_n4194), .Y(new_n4215_1));
  nand_5 g01867(.A(new_n4215_1), .B(new_n4193), .Y(new_n4216));
  nand_5 g01868(.A(new_n4216), .B(new_n4188), .Y(new_n4217));
  nand_5 g01869(.A(new_n4217), .B(new_n4187), .Y(new_n4218));
  not_8  g01870(.A(n3161), .Y(new_n4219));
  nand_5 g01871(.A(new_n4184), .B(new_n4176_1), .Y(new_n4220));
  nand_5 g01872(.A(new_n4220), .B(new_n4183), .Y(new_n4221_1));
  not_8  g01873(.A(n22597), .Y(new_n4222));
  nor_5  g01874(.A(new_n4179), .B(n21134), .Y(new_n4223));
  not_8  g01875(.A(new_n4223), .Y(new_n4224_1));
  nand_5 g01876(.A(new_n4179), .B(n21134), .Y(new_n4225));
  and_5  g01877(.A(new_n4225), .B(new_n4224_1), .Y(new_n4226));
  not_8  g01878(.A(new_n4226), .Y(new_n4227));
  nand_5 g01879(.A(new_n4227), .B(new_n4222), .Y(new_n4228));
  nand_5 g01880(.A(new_n4226), .B(n22597), .Y(new_n4229));
  nand_5 g01881(.A(new_n4229), .B(new_n4228), .Y(new_n4230));
  xor_4  g01882(.A(new_n4230), .B(new_n4221_1), .Y(new_n4231_1));
  not_8  g01883(.A(new_n4231_1), .Y(new_n4232));
  nand_5 g01884(.A(new_n4232), .B(new_n4219), .Y(new_n4233));
  nand_5 g01885(.A(new_n4231_1), .B(n3161), .Y(new_n4234));
  nand_5 g01886(.A(new_n4234), .B(new_n4233), .Y(new_n4235));
  xor_4  g01887(.A(new_n4235), .B(new_n4218), .Y(new_n4236));
  nand_5 g01888(.A(new_n4236), .B(new_n4145), .Y(new_n4237));
  or_5   g01889(.A(new_n4236), .B(new_n4145), .Y(new_n4238));
  nand_5 g01890(.A(new_n4094), .B(new_n4095), .Y(new_n4239));
  xor_4  g01891(.A(new_n4239), .B(new_n4127), .Y(new_n4240));
  nand_5 g01892(.A(new_n4187), .B(new_n4188), .Y(new_n4241));
  xor_4  g01893(.A(new_n4241), .B(new_n4216), .Y(new_n4242));
  nand_5 g01894(.A(new_n4242), .B(new_n4240), .Y(new_n4243));
  or_5   g01895(.A(new_n4242), .B(new_n4240), .Y(new_n4244));
  nand_5 g01896(.A(new_n4102), .B(new_n4100_1), .Y(new_n4245));
  xor_4  g01897(.A(new_n4245), .B(new_n4125), .Y(new_n4246));
  nand_5 g01898(.A(new_n4193), .B(new_n4194), .Y(new_n4247));
  xor_4  g01899(.A(new_n4247), .B(new_n4214), .Y(new_n4248));
  nand_5 g01900(.A(new_n4248), .B(new_n4246), .Y(new_n4249));
  or_5   g01901(.A(new_n4248), .B(new_n4246), .Y(new_n4250));
  nand_5 g01902(.A(new_n4124), .B(new_n4121), .Y(new_n4251));
  xor_4  g01903(.A(new_n4251), .B(new_n4116), .Y(new_n4252));
  nand_5 g01904(.A(new_n4199), .B(new_n4200), .Y(new_n4253));
  xor_4  g01905(.A(new_n4253), .B(new_n4212), .Y(new_n4254));
  nand_5 g01906(.A(new_n4254), .B(new_n4252), .Y(new_n4255));
  or_5   g01907(.A(new_n4254), .B(new_n4252), .Y(new_n4256_1));
  nand_5 g01908(.A(new_n4110), .B(new_n4108), .Y(new_n4257));
  xor_4  g01909(.A(new_n4257), .B(new_n4114), .Y(new_n4258));
  nand_5 g01910(.A(new_n4205_1), .B(new_n4206), .Y(new_n4259));
  xor_4  g01911(.A(new_n4259), .B(new_n4210), .Y(new_n4260));
  nand_5 g01912(.A(new_n4260), .B(new_n4258), .Y(new_n4261));
  or_5   g01913(.A(new_n4260), .B(new_n4258), .Y(new_n4262));
  nand_5 g01914(.A(new_n4112), .B(new_n4084), .Y(new_n4263));
  and_5  g01915(.A(new_n4263), .B(new_n4114), .Y(new_n4264));
  xor_4  g01916(.A(new_n4209), .B(n20658), .Y(new_n4265));
  and_5  g01917(.A(new_n4265), .B(new_n4264), .Y(new_n4266_1));
  nand_5 g01918(.A(new_n4266_1), .B(new_n4262), .Y(new_n4267));
  nand_5 g01919(.A(new_n4267), .B(new_n4261), .Y(new_n4268));
  nand_5 g01920(.A(new_n4268), .B(new_n4256_1), .Y(new_n4269));
  nand_5 g01921(.A(new_n4269), .B(new_n4255), .Y(new_n4270));
  nand_5 g01922(.A(new_n4270), .B(new_n4250), .Y(new_n4271));
  nand_5 g01923(.A(new_n4271), .B(new_n4249), .Y(new_n4272_1));
  nand_5 g01924(.A(new_n4272_1), .B(new_n4244), .Y(new_n4273));
  nand_5 g01925(.A(new_n4273), .B(new_n4243), .Y(new_n4274));
  nand_5 g01926(.A(new_n4274), .B(new_n4238), .Y(new_n4275));
  nand_5 g01927(.A(new_n4275), .B(new_n4237), .Y(new_n4276));
  nand_5 g01928(.A(new_n4143), .B(new_n4129), .Y(new_n4277));
  nand_5 g01929(.A(new_n4277), .B(new_n4142), .Y(new_n4278));
  nand_5 g01930(.A(new_n4133), .B(new_n4131), .Y(new_n4279));
  nand_5 g01931(.A(new_n4279), .B(new_n4132), .Y(new_n4280));
  not_8  g01932(.A(new_n4280), .Y(new_n4281));
  nand_5 g01933(.A(new_n3109), .B(n22332), .Y(new_n4282));
  nand_5 g01934(.A(n26510), .B(new_n2569), .Y(new_n4283));
  nand_5 g01935(.A(new_n4283), .B(new_n4282), .Y(new_n4284));
  xor_4  g01936(.A(new_n4284), .B(new_n4281), .Y(new_n4285));
  xor_4  g01937(.A(new_n4138), .B(n4325), .Y(new_n4286));
  nand_5 g01938(.A(new_n4286), .B(new_n4285), .Y(new_n4287));
  or_5   g01939(.A(new_n4286), .B(new_n4285), .Y(new_n4288));
  nand_5 g01940(.A(new_n4288), .B(new_n4287), .Y(new_n4289));
  xor_4  g01941(.A(new_n4289), .B(new_n4278), .Y(new_n4290));
  nand_5 g01942(.A(new_n4234), .B(new_n4218), .Y(new_n4291));
  nand_5 g01943(.A(new_n4291), .B(new_n4233), .Y(new_n4292));
  not_8  g01944(.A(n25749), .Y(new_n4293));
  nand_5 g01945(.A(new_n4229), .B(new_n4221_1), .Y(new_n4294));
  nand_5 g01946(.A(new_n4294), .B(new_n4228), .Y(new_n4295));
  not_8  g01947(.A(new_n4295), .Y(new_n4296));
  not_8  g01948(.A(n19327), .Y(new_n4297));
  not_8  g01949(.A(n2113), .Y(new_n4298));
  nand_5 g01950(.A(new_n4223), .B(new_n4298), .Y(new_n4299));
  nand_5 g01951(.A(new_n4224_1), .B(n2113), .Y(new_n4300));
  and_5  g01952(.A(new_n4300), .B(new_n4299), .Y(new_n4301));
  not_8  g01953(.A(new_n4301), .Y(new_n4302));
  nand_5 g01954(.A(new_n4302), .B(new_n4297), .Y(new_n4303));
  nand_5 g01955(.A(new_n4301), .B(n19327), .Y(new_n4304));
  nand_5 g01956(.A(new_n4304), .B(new_n4303), .Y(new_n4305));
  xor_4  g01957(.A(new_n4305), .B(new_n4296), .Y(new_n4306_1));
  nand_5 g01958(.A(new_n4306_1), .B(new_n4293), .Y(new_n4307));
  or_5   g01959(.A(new_n4306_1), .B(new_n4293), .Y(new_n4308));
  nand_5 g01960(.A(new_n4308), .B(new_n4307), .Y(new_n4309));
  xor_4  g01961(.A(new_n4309), .B(new_n4292), .Y(new_n4310));
  or_5   g01962(.A(new_n4310), .B(new_n4290), .Y(new_n4311));
  nand_5 g01963(.A(new_n4310), .B(new_n4290), .Y(new_n4312));
  nand_5 g01964(.A(new_n4312), .B(new_n4311), .Y(new_n4313));
  xnor_4 g01965(.A(new_n4313), .B(new_n4276), .Y(n242));
  not_8  g01966(.A(n5451), .Y(new_n4315));
  nand_5 g01967(.A(new_n2632), .B(new_n2674), .Y(new_n4316));
  nand_5 g01968(.A(n21398), .B(n11667), .Y(new_n4317));
  and_5  g01969(.A(new_n4317), .B(new_n4316), .Y(new_n4318));
  nand_5 g01970(.A(new_n4318), .B(n22433), .Y(new_n4319_1));
  nand_5 g01971(.A(new_n4319_1), .B(new_n2630), .Y(new_n4320));
  or_5   g01972(.A(new_n4318), .B(n22433), .Y(new_n4321));
  nand_5 g01973(.A(new_n4321), .B(new_n4320), .Y(new_n4322));
  xor_4  g01974(.A(new_n4316), .B(n26572), .Y(new_n4323));
  nand_5 g01975(.A(new_n4323), .B(n11615), .Y(new_n4324));
  nand_5 g01976(.A(new_n4324), .B(new_n4322), .Y(new_n4325_1));
  nor_5  g01977(.A(new_n4323), .B(n11615), .Y(new_n4326_1));
  not_8  g01978(.A(new_n4326_1), .Y(new_n4327));
  nand_5 g01979(.A(new_n4327), .B(new_n4325_1), .Y(new_n4328));
  not_8  g01980(.A(new_n4328), .Y(new_n4329));
  or_5   g01981(.A(new_n4316), .B(n26572), .Y(new_n4330));
  xor_4  g01982(.A(new_n4330), .B(n5115), .Y(new_n4331));
  nand_5 g01983(.A(new_n4331), .B(n16476), .Y(new_n4332));
  nor_5  g01984(.A(new_n4331), .B(n16476), .Y(new_n4333));
  not_8  g01985(.A(new_n4333), .Y(new_n4334));
  nand_5 g01986(.A(new_n4334), .B(new_n4332), .Y(new_n4335));
  xor_4  g01987(.A(new_n4335), .B(new_n4329), .Y(new_n4336));
  nand_5 g01988(.A(new_n4336), .B(new_n4315), .Y(new_n4337));
  not_8  g01989(.A(new_n4336), .Y(new_n4338));
  nand_5 g01990(.A(new_n4338), .B(n5451), .Y(new_n4339));
  not_8  g01991(.A(n5330), .Y(new_n4340_1));
  nand_5 g01992(.A(new_n4327), .B(new_n4324), .Y(new_n4341));
  xor_4  g01993(.A(new_n4341), .B(new_n4322), .Y(new_n4342));
  not_8  g01994(.A(new_n4342), .Y(new_n4343));
  nand_5 g01995(.A(new_n4343), .B(new_n4340_1), .Y(new_n4344));
  nand_5 g01996(.A(new_n4342), .B(n5330), .Y(new_n4345));
  not_8  g01997(.A(n7657), .Y(new_n4346));
  and_5  g01998(.A(new_n4321), .B(new_n4319_1), .Y(new_n4347));
  xor_4  g01999(.A(new_n4347), .B(new_n2630), .Y(new_n4348));
  nand_5 g02000(.A(new_n4348), .B(new_n4346), .Y(new_n4349));
  nand_5 g02001(.A(new_n2634), .B(n25926), .Y(new_n4350));
  not_8  g02002(.A(new_n4348), .Y(new_n4351));
  nand_5 g02003(.A(new_n4351), .B(n7657), .Y(new_n4352));
  nand_5 g02004(.A(new_n4352), .B(new_n4350), .Y(new_n4353));
  nand_5 g02005(.A(new_n4353), .B(new_n4349), .Y(new_n4354));
  nand_5 g02006(.A(new_n4354), .B(new_n4345), .Y(new_n4355));
  nand_5 g02007(.A(new_n4355), .B(new_n4344), .Y(new_n4356));
  nand_5 g02008(.A(new_n4356), .B(new_n4339), .Y(new_n4357));
  nand_5 g02009(.A(new_n4357), .B(new_n4337), .Y(new_n4358));
  not_8  g02010(.A(n18926), .Y(new_n4359));
  nand_5 g02011(.A(new_n4332), .B(new_n4328), .Y(new_n4360));
  nand_5 g02012(.A(new_n4360), .B(new_n4334), .Y(new_n4361));
  not_8  g02013(.A(new_n4361), .Y(new_n4362));
  nor_5  g02014(.A(new_n4330), .B(n5115), .Y(new_n4363));
  xor_4  g02015(.A(new_n4363), .B(new_n2664), .Y(new_n4364));
  nand_5 g02016(.A(new_n4364), .B(n16029), .Y(new_n4365));
  nor_5  g02017(.A(new_n4364), .B(n16029), .Y(new_n4366));
  not_8  g02018(.A(new_n4366), .Y(new_n4367));
  nand_5 g02019(.A(new_n4367), .B(new_n4365), .Y(new_n4368));
  xor_4  g02020(.A(new_n4368), .B(new_n4362), .Y(new_n4369));
  nand_5 g02021(.A(new_n4369), .B(new_n4359), .Y(new_n4370));
  not_8  g02022(.A(new_n4369), .Y(new_n4371));
  nand_5 g02023(.A(new_n4371), .B(n18926), .Y(new_n4372));
  nand_5 g02024(.A(new_n4372), .B(new_n4370), .Y(new_n4373));
  xor_4  g02025(.A(new_n4373), .B(new_n4358), .Y(new_n4374_1));
  not_8  g02026(.A(new_n4374_1), .Y(new_n4375));
  not_8  g02027(.A(n11302), .Y(new_n4376_1));
  not_8  g02028(.A(n10792), .Y(new_n4377));
  not_8  g02029(.A(n19922), .Y(new_n4378));
  nand_5 g02030(.A(new_n4378), .B(new_n4377), .Y(new_n4379));
  or_5   g02031(.A(new_n4379), .B(n9323), .Y(new_n4380));
  nand_5 g02032(.A(new_n4379), .B(n9323), .Y(new_n4381));
  and_5  g02033(.A(new_n4381), .B(new_n4380), .Y(new_n4382));
  not_8  g02034(.A(new_n4382), .Y(new_n4383));
  nand_5 g02035(.A(new_n4383), .B(new_n4376_1), .Y(new_n4384));
  nand_5 g02036(.A(new_n4382), .B(n11302), .Y(new_n4385));
  not_8  g02037(.A(n17090), .Y(new_n4386));
  nand_5 g02038(.A(n19922), .B(n10792), .Y(new_n4387));
  and_5  g02039(.A(new_n4387), .B(new_n4379), .Y(new_n4388));
  not_8  g02040(.A(new_n4388), .Y(new_n4389));
  nand_5 g02041(.A(new_n4389), .B(new_n4386), .Y(new_n4390));
  nand_5 g02042(.A(new_n4388), .B(n17090), .Y(new_n4391));
  nand_5 g02043(.A(new_n4391), .B(new_n2637), .Y(new_n4392));
  nand_5 g02044(.A(new_n4392), .B(new_n4390), .Y(new_n4393));
  nand_5 g02045(.A(new_n4393), .B(new_n4385), .Y(new_n4394));
  nand_5 g02046(.A(new_n4394), .B(new_n4384), .Y(new_n4395));
  not_8  g02047(.A(n10405), .Y(new_n4396));
  nor_5  g02048(.A(new_n4380), .B(n1949), .Y(new_n4397));
  not_8  g02049(.A(new_n4397), .Y(new_n4398));
  nand_5 g02050(.A(new_n4380), .B(n1949), .Y(new_n4399));
  and_5  g02051(.A(new_n4399), .B(new_n4398), .Y(new_n4400));
  not_8  g02052(.A(new_n4400), .Y(new_n4401_1));
  nand_5 g02053(.A(new_n4401_1), .B(new_n4396), .Y(new_n4402));
  nand_5 g02054(.A(new_n4400), .B(n10405), .Y(new_n4403));
  nand_5 g02055(.A(new_n4403), .B(new_n4402), .Y(new_n4404));
  xor_4  g02056(.A(new_n4404), .B(new_n4395), .Y(new_n4405));
  not_8  g02057(.A(new_n4405), .Y(new_n4406));
  not_8  g02058(.A(n20169), .Y(new_n4407));
  not_8  g02059(.A(n8285), .Y(new_n4408));
  nor_5  g02060(.A(n21687), .B(n6729), .Y(new_n4409_1));
  nand_5 g02061(.A(new_n4409_1), .B(new_n4408), .Y(new_n4410));
  xor_4  g02062(.A(new_n4410), .B(new_n4407), .Y(new_n4411));
  or_5   g02063(.A(new_n4411), .B(new_n4406), .Y(new_n4412));
  nand_5 g02064(.A(new_n4411), .B(new_n4406), .Y(new_n4413));
  nand_5 g02065(.A(new_n4385), .B(new_n4384), .Y(new_n4414));
  xor_4  g02066(.A(new_n4414), .B(new_n4393), .Y(new_n4415));
  xor_4  g02067(.A(new_n4409_1), .B(new_n4408), .Y(new_n4416));
  nand_5 g02068(.A(new_n4416), .B(new_n4415), .Y(new_n4417));
  nor_5  g02069(.A(new_n4416), .B(new_n4415), .Y(new_n4418));
  not_8  g02070(.A(new_n4418), .Y(new_n4419));
  and_5  g02071(.A(new_n4391), .B(new_n4390), .Y(new_n4420));
  xor_4  g02072(.A(new_n4420), .B(new_n2638), .Y(new_n4421));
  not_8  g02073(.A(n6729), .Y(new_n4422));
  nor_5  g02074(.A(new_n2636), .B(new_n4422), .Y(new_n4423));
  nor_5  g02075(.A(new_n4423), .B(new_n4409_1), .Y(new_n4424_1));
  or_5   g02076(.A(new_n4424_1), .B(new_n4421), .Y(new_n4425));
  not_8  g02077(.A(new_n2640), .Y(new_n4426_1));
  nand_5 g02078(.A(new_n4426_1), .B(n21687), .Y(new_n4427));
  nand_5 g02079(.A(new_n4424_1), .B(new_n4421), .Y(new_n4428));
  nand_5 g02080(.A(new_n4428), .B(new_n4427), .Y(new_n4429));
  nand_5 g02081(.A(new_n4429), .B(new_n4425), .Y(new_n4430));
  not_8  g02082(.A(new_n4430), .Y(new_n4431));
  nand_5 g02083(.A(new_n4431), .B(new_n4419), .Y(new_n4432_1));
  nand_5 g02084(.A(new_n4432_1), .B(new_n4417), .Y(new_n4433));
  nand_5 g02085(.A(new_n4433), .B(new_n4413), .Y(new_n4434));
  nand_5 g02086(.A(new_n4434), .B(new_n4412), .Y(new_n4435));
  nand_5 g02087(.A(new_n4403), .B(new_n4395), .Y(new_n4436));
  nand_5 g02088(.A(new_n4436), .B(new_n4402), .Y(new_n4437));
  not_8  g02089(.A(n7693), .Y(new_n4438));
  not_8  g02090(.A(n15424), .Y(new_n4439));
  nand_5 g02091(.A(new_n4397), .B(new_n4439), .Y(new_n4440));
  nand_5 g02092(.A(new_n4398), .B(n15424), .Y(new_n4441_1));
  and_5  g02093(.A(new_n4441_1), .B(new_n4440), .Y(new_n4442));
  not_8  g02094(.A(new_n4442), .Y(new_n4443));
  nand_5 g02095(.A(new_n4443), .B(new_n4438), .Y(new_n4444));
  nand_5 g02096(.A(new_n4442), .B(n7693), .Y(new_n4445));
  nand_5 g02097(.A(new_n4445), .B(new_n4444), .Y(new_n4446));
  xor_4  g02098(.A(new_n4446), .B(new_n4437), .Y(new_n4447));
  not_8  g02099(.A(new_n4447), .Y(new_n4448));
  nor_5  g02100(.A(new_n4410), .B(n20169), .Y(new_n4449));
  xor_4  g02101(.A(new_n4449), .B(n19789), .Y(new_n4450));
  or_5   g02102(.A(new_n4450), .B(new_n4448), .Y(new_n4451_1));
  nand_5 g02103(.A(new_n4450), .B(new_n4448), .Y(new_n4452));
  nand_5 g02104(.A(new_n4452), .B(new_n4451_1), .Y(new_n4453));
  xor_4  g02105(.A(new_n4453), .B(new_n4435), .Y(new_n4454));
  or_5   g02106(.A(new_n4454), .B(new_n4375), .Y(new_n4455));
  nand_5 g02107(.A(new_n4454), .B(new_n4375), .Y(new_n4456));
  nand_5 g02108(.A(new_n4337), .B(new_n4339), .Y(new_n4457));
  xor_4  g02109(.A(new_n4457), .B(new_n4356), .Y(new_n4458));
  not_8  g02110(.A(new_n4458), .Y(new_n4459));
  nand_5 g02111(.A(new_n4413), .B(new_n4412), .Y(new_n4460));
  xor_4  g02112(.A(new_n4460), .B(new_n4433), .Y(new_n4461));
  or_5   g02113(.A(new_n4461), .B(new_n4459), .Y(new_n4462));
  nand_5 g02114(.A(new_n4461), .B(new_n4459), .Y(new_n4463));
  nand_5 g02115(.A(new_n4344), .B(new_n4345), .Y(new_n4464));
  xor_4  g02116(.A(new_n4464), .B(new_n4354), .Y(new_n4465));
  not_8  g02117(.A(new_n4465), .Y(new_n4466));
  nand_5 g02118(.A(new_n4419), .B(new_n4417), .Y(new_n4467));
  xor_4  g02119(.A(new_n4467), .B(new_n4431), .Y(new_n4468));
  or_5   g02120(.A(new_n4468), .B(new_n4466), .Y(new_n4469));
  nand_5 g02121(.A(new_n4468), .B(new_n4466), .Y(new_n4470));
  nand_5 g02122(.A(new_n4349), .B(new_n4352), .Y(new_n4471));
  xor_4  g02123(.A(new_n4471), .B(new_n4350), .Y(new_n4472));
  nand_5 g02124(.A(new_n4428), .B(new_n4425), .Y(new_n4473));
  xor_4  g02125(.A(new_n4473), .B(new_n4427), .Y(new_n4474));
  nand_5 g02126(.A(new_n4474), .B(new_n4472), .Y(new_n4475));
  nor_5  g02127(.A(new_n4474), .B(new_n4472), .Y(new_n4476_1));
  not_8  g02128(.A(new_n4476_1), .Y(new_n4477));
  nand_5 g02129(.A(new_n4477), .B(new_n2643), .Y(new_n4478_1));
  nand_5 g02130(.A(new_n4478_1), .B(new_n4475), .Y(new_n4479));
  nand_5 g02131(.A(new_n4479), .B(new_n4470), .Y(new_n4480));
  nand_5 g02132(.A(new_n4480), .B(new_n4469), .Y(new_n4481));
  nand_5 g02133(.A(new_n4481), .B(new_n4463), .Y(new_n4482));
  nand_5 g02134(.A(new_n4482), .B(new_n4462), .Y(new_n4483));
  nand_5 g02135(.A(new_n4483), .B(new_n4456), .Y(new_n4484));
  nand_5 g02136(.A(new_n4484), .B(new_n4455), .Y(new_n4485));
  not_8  g02137(.A(new_n4485), .Y(new_n4486));
  nand_5 g02138(.A(new_n4372), .B(new_n4358), .Y(new_n4487));
  nand_5 g02139(.A(new_n4487), .B(new_n4370), .Y(new_n4488));
  not_8  g02140(.A(n13677), .Y(new_n4489));
  nand_5 g02141(.A(new_n4365), .B(new_n4361), .Y(new_n4490));
  nand_5 g02142(.A(new_n4490), .B(new_n4367), .Y(new_n4491));
  not_8  g02143(.A(new_n4491), .Y(new_n4492));
  nand_5 g02144(.A(new_n4363), .B(new_n2664), .Y(new_n4493));
  nor_5  g02145(.A(new_n4493), .B(n19477), .Y(new_n4494));
  not_8  g02146(.A(new_n4494), .Y(new_n4495));
  nand_5 g02147(.A(new_n4493), .B(n19477), .Y(new_n4496));
  and_5  g02148(.A(new_n4496), .B(new_n4495), .Y(new_n4497));
  or_5   g02149(.A(new_n4497), .B(n11011), .Y(new_n4498));
  nand_5 g02150(.A(new_n4497), .B(n11011), .Y(new_n4499));
  nand_5 g02151(.A(new_n4499), .B(new_n4498), .Y(new_n4500));
  xor_4  g02152(.A(new_n4500), .B(new_n4492), .Y(new_n4501));
  nand_5 g02153(.A(new_n4501), .B(new_n4489), .Y(new_n4502));
  not_8  g02154(.A(new_n4501), .Y(new_n4503));
  nand_5 g02155(.A(new_n4503), .B(n13677), .Y(new_n4504));
  nand_5 g02156(.A(new_n4504), .B(new_n4502), .Y(new_n4505));
  xor_4  g02157(.A(new_n4505), .B(new_n4488), .Y(new_n4506));
  not_8  g02158(.A(new_n4506), .Y(new_n4507));
  nand_5 g02159(.A(new_n4452), .B(new_n4435), .Y(new_n4508));
  nand_5 g02160(.A(new_n4508), .B(new_n4451_1), .Y(new_n4509));
  nand_5 g02161(.A(new_n4445), .B(new_n4437), .Y(new_n4510));
  nand_5 g02162(.A(new_n4510), .B(new_n4444), .Y(new_n4511));
  not_8  g02163(.A(n20151), .Y(new_n4512));
  nor_5  g02164(.A(new_n4440), .B(n25694), .Y(new_n4513));
  not_8  g02165(.A(new_n4513), .Y(new_n4514_1));
  nand_5 g02166(.A(new_n4440), .B(n25694), .Y(new_n4515));
  and_5  g02167(.A(new_n4515), .B(new_n4514_1), .Y(new_n4516));
  not_8  g02168(.A(new_n4516), .Y(new_n4517));
  nand_5 g02169(.A(new_n4517), .B(new_n4512), .Y(new_n4518));
  nand_5 g02170(.A(new_n4516), .B(n20151), .Y(new_n4519));
  nand_5 g02171(.A(new_n4519), .B(new_n4518), .Y(new_n4520));
  xnor_4 g02172(.A(new_n4520), .B(new_n4511), .Y(new_n4521));
  not_8  g02173(.A(n12398), .Y(new_n4522));
  not_8  g02174(.A(n19789), .Y(new_n4523));
  nand_5 g02175(.A(new_n4449), .B(new_n4523), .Y(new_n4524));
  xor_4  g02176(.A(new_n4524), .B(new_n4522), .Y(new_n4525));
  or_5   g02177(.A(new_n4525), .B(new_n4521), .Y(new_n4526));
  nand_5 g02178(.A(new_n4525), .B(new_n4521), .Y(new_n4527));
  nand_5 g02179(.A(new_n4527), .B(new_n4526), .Y(new_n4528));
  xor_4  g02180(.A(new_n4528), .B(new_n4509), .Y(new_n4529_1));
  nand_5 g02181(.A(new_n4529_1), .B(new_n4507), .Y(new_n4530));
  or_5   g02182(.A(new_n4529_1), .B(new_n4507), .Y(new_n4531));
  nand_5 g02183(.A(new_n4531), .B(new_n4530), .Y(new_n4532));
  xor_4  g02184(.A(new_n4532), .B(new_n4486), .Y(n243));
  nand_5 g02185(.A(n25926), .B(n20385), .Y(new_n4534));
  not_8  g02186(.A(n25316), .Y(new_n4535));
  nand_5 g02187(.A(new_n4535), .B(new_n4346), .Y(new_n4536));
  nand_5 g02188(.A(n25316), .B(n7657), .Y(new_n4537));
  nand_5 g02189(.A(new_n4537), .B(new_n4536), .Y(new_n4538));
  xnor_4 g02190(.A(new_n4538), .B(new_n4534), .Y(new_n4539));
  nand_5 g02191(.A(n23065), .B(n6773), .Y(new_n4540));
  not_8  g02192(.A(n6773), .Y(new_n4541));
  not_8  g02193(.A(n23065), .Y(new_n4542));
  nand_5 g02194(.A(new_n4542), .B(new_n4541), .Y(new_n4543));
  and_5  g02195(.A(new_n4543), .B(new_n4540), .Y(new_n4544));
  not_8  g02196(.A(n9380), .Y(new_n4545));
  nand_5 g02197(.A(n24129), .B(new_n4545), .Y(new_n4546));
  not_8  g02198(.A(n24129), .Y(new_n4547));
  nand_5 g02199(.A(new_n4547), .B(n9380), .Y(new_n4548));
  and_5  g02200(.A(new_n4548), .B(new_n4546), .Y(new_n4549));
  not_8  g02201(.A(new_n4549), .Y(new_n4550));
  nand_5 g02202(.A(new_n4550), .B(new_n4544), .Y(new_n4551));
  not_8  g02203(.A(new_n4540), .Y(new_n4552_1));
  not_8  g02204(.A(n27120), .Y(new_n4553));
  nand_5 g02205(.A(new_n4553), .B(new_n4386), .Y(new_n4554));
  nand_5 g02206(.A(n27120), .B(n17090), .Y(new_n4555));
  nand_5 g02207(.A(new_n4555), .B(new_n4554), .Y(new_n4556));
  xor_4  g02208(.A(new_n4556), .B(new_n4552_1), .Y(new_n4557));
  not_8  g02209(.A(new_n4546), .Y(new_n4558));
  not_8  g02210(.A(n22274), .Y(new_n4559));
  nand_5 g02211(.A(new_n4559), .B(n11192), .Y(new_n4560));
  not_8  g02212(.A(n11192), .Y(new_n4561));
  nand_5 g02213(.A(n22274), .B(new_n4561), .Y(new_n4562));
  and_5  g02214(.A(new_n4562), .B(new_n4560), .Y(new_n4563));
  xor_4  g02215(.A(new_n4563), .B(new_n4558), .Y(new_n4564));
  nand_5 g02216(.A(new_n4564), .B(new_n4557), .Y(new_n4565));
  not_8  g02217(.A(new_n4557), .Y(new_n4566));
  not_8  g02218(.A(new_n4564), .Y(new_n4567));
  nand_5 g02219(.A(new_n4567), .B(new_n4566), .Y(new_n4568));
  nand_5 g02220(.A(new_n4568), .B(new_n4565), .Y(new_n4569));
  xor_4  g02221(.A(new_n4569), .B(new_n4551), .Y(new_n4570));
  nand_5 g02222(.A(new_n4570), .B(new_n4539), .Y(new_n4571));
  or_5   g02223(.A(new_n4570), .B(new_n4539), .Y(new_n4572));
  not_8  g02224(.A(n20385), .Y(new_n4573));
  not_8  g02225(.A(n25926), .Y(new_n4574));
  nand_5 g02226(.A(new_n4574), .B(new_n4573), .Y(new_n4575));
  and_5  g02227(.A(new_n4575), .B(new_n4534), .Y(new_n4576));
  not_8  g02228(.A(new_n4576), .Y(new_n4577));
  not_8  g02229(.A(new_n4544), .Y(new_n4578));
  nand_5 g02230(.A(new_n4549), .B(new_n4578), .Y(new_n4579));
  and_5  g02231(.A(new_n4579), .B(new_n4551), .Y(new_n4580));
  or_5   g02232(.A(new_n4580), .B(new_n4577), .Y(new_n4581));
  nand_5 g02233(.A(new_n4581), .B(new_n4572), .Y(new_n4582));
  nand_5 g02234(.A(new_n4582), .B(new_n4571), .Y(new_n4583));
  nand_5 g02235(.A(new_n4537), .B(new_n4534), .Y(new_n4584));
  nand_5 g02236(.A(new_n4584), .B(new_n4536), .Y(new_n4585));
  not_8  g02237(.A(n919), .Y(new_n4586));
  nand_5 g02238(.A(new_n4340_1), .B(new_n4586), .Y(new_n4587));
  nand_5 g02239(.A(n5330), .B(n919), .Y(new_n4588_1));
  nand_5 g02240(.A(new_n4588_1), .B(new_n4587), .Y(new_n4589));
  xnor_4 g02241(.A(new_n4589), .B(new_n4585), .Y(new_n4590_1));
  nand_5 g02242(.A(new_n4568), .B(new_n4551), .Y(new_n4591));
  nand_5 g02243(.A(new_n4591), .B(new_n4565), .Y(new_n4592));
  nand_5 g02244(.A(new_n4555), .B(new_n4540), .Y(new_n4593));
  nand_5 g02245(.A(new_n4593), .B(new_n4554), .Y(new_n4594));
  not_8  g02246(.A(new_n4594), .Y(new_n4595_1));
  not_8  g02247(.A(n24786), .Y(new_n4596));
  nand_5 g02248(.A(new_n4596), .B(new_n4376_1), .Y(new_n4597));
  nand_5 g02249(.A(n24786), .B(n11302), .Y(new_n4598));
  nand_5 g02250(.A(new_n4598), .B(new_n4597), .Y(new_n4599));
  xor_4  g02251(.A(new_n4599), .B(new_n4595_1), .Y(new_n4600));
  nand_5 g02252(.A(new_n4562), .B(new_n4546), .Y(new_n4601));
  nand_5 g02253(.A(new_n4601), .B(new_n4560), .Y(new_n4602));
  not_8  g02254(.A(new_n4602), .Y(new_n4603));
  not_8  g02255(.A(n1689), .Y(new_n4604));
  nand_5 g02256(.A(n20036), .B(new_n4604), .Y(new_n4605));
  not_8  g02257(.A(n20036), .Y(new_n4606));
  nand_5 g02258(.A(new_n4606), .B(n1689), .Y(new_n4607));
  nand_5 g02259(.A(new_n4607), .B(new_n4605), .Y(new_n4608));
  xor_4  g02260(.A(new_n4608), .B(new_n4603), .Y(new_n4609));
  not_8  g02261(.A(new_n4609), .Y(new_n4610));
  nand_5 g02262(.A(new_n4610), .B(new_n4600), .Y(new_n4611));
  not_8  g02263(.A(new_n4600), .Y(new_n4612));
  nand_5 g02264(.A(new_n4609), .B(new_n4612), .Y(new_n4613));
  nand_5 g02265(.A(new_n4613), .B(new_n4611), .Y(new_n4614));
  xor_4  g02266(.A(new_n4614), .B(new_n4592), .Y(new_n4615));
  nand_5 g02267(.A(new_n4615), .B(new_n4590_1), .Y(new_n4616));
  or_5   g02268(.A(new_n4615), .B(new_n4590_1), .Y(new_n4617));
  nand_5 g02269(.A(new_n4617), .B(new_n4616), .Y(new_n4618));
  xnor_4 g02270(.A(new_n4618), .B(new_n4583), .Y(n248));
  not_8  g02271(.A(n14684), .Y(new_n4620));
  not_8  g02272(.A(n6631), .Y(new_n4621));
  not_8  g02273(.A(n24732), .Y(new_n4622));
  nand_5 g02274(.A(new_n4622), .B(new_n4621), .Y(new_n4623));
  not_8  g02275(.A(new_n4623), .Y(new_n4624_1));
  nand_5 g02276(.A(new_n4624_1), .B(new_n4620), .Y(new_n4625));
  nand_5 g02277(.A(new_n4623), .B(n14684), .Y(new_n4626));
  nand_5 g02278(.A(new_n4626), .B(new_n4625), .Y(new_n4627));
  nand_5 g02279(.A(new_n4627), .B(new_n4147), .Y(new_n4628));
  nor_5  g02280(.A(new_n4627), .B(new_n4147), .Y(new_n4629));
  not_8  g02281(.A(new_n4629), .Y(new_n4630));
  nand_5 g02282(.A(n24732), .B(n6631), .Y(new_n4631));
  and_5  g02283(.A(new_n4631), .B(new_n4623), .Y(new_n4632));
  or_5   g02284(.A(new_n4632), .B(n13319), .Y(new_n4633));
  nand_5 g02285(.A(new_n4632), .B(n13319), .Y(new_n4634));
  nand_5 g02286(.A(n25435), .B(n24732), .Y(new_n4635));
  nand_5 g02287(.A(new_n4635), .B(new_n4634), .Y(new_n4636));
  nand_5 g02288(.A(new_n4636), .B(new_n4633), .Y(new_n4637));
  nand_5 g02289(.A(new_n4637), .B(new_n4630), .Y(new_n4638));
  nand_5 g02290(.A(new_n4638), .B(new_n4628), .Y(new_n4639));
  not_8  g02291(.A(new_n4639), .Y(new_n4640));
  not_8  g02292(.A(n25797), .Y(new_n4641));
  not_8  g02293(.A(n17035), .Y(new_n4642));
  not_8  g02294(.A(new_n4625), .Y(new_n4643));
  nand_5 g02295(.A(new_n4643), .B(new_n4642), .Y(new_n4644));
  nand_5 g02296(.A(new_n4625), .B(n17035), .Y(new_n4645));
  nand_5 g02297(.A(new_n4645), .B(new_n4644), .Y(new_n4646_1));
  nand_5 g02298(.A(new_n4646_1), .B(new_n4641), .Y(new_n4647));
  nor_5  g02299(.A(new_n4646_1), .B(new_n4641), .Y(new_n4648));
  not_8  g02300(.A(new_n4648), .Y(new_n4649));
  nand_5 g02301(.A(new_n4649), .B(new_n4647), .Y(new_n4650));
  xor_4  g02302(.A(new_n4650), .B(new_n4640), .Y(new_n4651));
  nand_5 g02303(.A(n12121), .B(n8920), .Y(new_n4652));
  not_8  g02304(.A(n8920), .Y(new_n4653));
  not_8  g02305(.A(n10057), .Y(new_n4654));
  nand_5 g02306(.A(new_n4654), .B(new_n4653), .Y(new_n4655));
  nand_5 g02307(.A(n10057), .B(n8920), .Y(new_n4656));
  and_5  g02308(.A(new_n4656), .B(new_n4655), .Y(new_n4657));
  nand_5 g02309(.A(new_n4657), .B(n22043), .Y(new_n4658));
  nand_5 g02310(.A(new_n4658), .B(new_n4652), .Y(new_n4659));
  or_5   g02311(.A(new_n4657), .B(n22043), .Y(new_n4660));
  nand_5 g02312(.A(new_n4660), .B(new_n4659), .Y(new_n4661));
  not_8  g02313(.A(new_n4661), .Y(new_n4662));
  xor_4  g02314(.A(new_n4655), .B(n26748), .Y(new_n4663));
  nand_5 g02315(.A(new_n4663), .B(n19618), .Y(new_n4664));
  nor_5  g02316(.A(new_n4663), .B(n19618), .Y(new_n4665_1));
  not_8  g02317(.A(new_n4665_1), .Y(new_n4666));
  nand_5 g02318(.A(new_n4666), .B(new_n4664), .Y(new_n4667));
  xor_4  g02319(.A(new_n4667), .B(new_n4662), .Y(new_n4668));
  not_8  g02320(.A(new_n4668), .Y(new_n4669));
  nand_5 g02321(.A(new_n2809_1), .B(new_n3248), .Y(new_n4670));
  nand_5 g02322(.A(n14148), .B(n1152), .Y(new_n4671));
  and_5  g02323(.A(new_n4671), .B(new_n4670), .Y(new_n4672));
  not_8  g02324(.A(new_n4672), .Y(new_n4673));
  nand_5 g02325(.A(new_n4673), .B(new_n3090), .Y(new_n4674_1));
  nand_5 g02326(.A(new_n4672), .B(n9507), .Y(new_n4675));
  nand_5 g02327(.A(n26979), .B(n1152), .Y(new_n4676));
  nand_5 g02328(.A(new_n4676), .B(new_n4675), .Y(new_n4677));
  nand_5 g02329(.A(new_n4677), .B(new_n4674_1), .Y(new_n4678));
  not_8  g02330(.A(new_n4678), .Y(new_n4679));
  or_5   g02331(.A(new_n4670), .B(n7149), .Y(new_n4680));
  nand_5 g02332(.A(new_n4670), .B(n7149), .Y(new_n4681));
  and_5  g02333(.A(new_n4681), .B(new_n4680), .Y(new_n4682));
  not_8  g02334(.A(new_n4682), .Y(new_n4683));
  nand_5 g02335(.A(new_n4683), .B(new_n3085), .Y(new_n4684));
  nand_5 g02336(.A(new_n4682), .B(n8399), .Y(new_n4685));
  nand_5 g02337(.A(new_n4685), .B(new_n4684), .Y(new_n4686));
  xor_4  g02338(.A(new_n4686), .B(new_n4679), .Y(new_n4687));
  not_8  g02339(.A(new_n4687), .Y(new_n4688));
  nand_5 g02340(.A(new_n4688), .B(new_n4669), .Y(new_n4689));
  nand_5 g02341(.A(new_n4687), .B(new_n4668), .Y(new_n4690));
  nand_5 g02342(.A(new_n4660), .B(new_n4658), .Y(new_n4691));
  xor_4  g02343(.A(new_n4691), .B(new_n4652), .Y(new_n4692));
  and_5  g02344(.A(new_n4675), .B(new_n4674_1), .Y(new_n4693_1));
  xor_4  g02345(.A(new_n4693_1), .B(new_n4676), .Y(new_n4694));
  not_8  g02346(.A(new_n4694), .Y(new_n4695));
  nand_5 g02347(.A(new_n4695), .B(new_n4692), .Y(new_n4696));
  nand_5 g02348(.A(new_n4694), .B(new_n4691), .Y(new_n4697));
  nand_5 g02349(.A(new_n4084), .B(new_n4653), .Y(new_n4698));
  and_5  g02350(.A(new_n4698), .B(new_n4652), .Y(new_n4699));
  nand_5 g02351(.A(new_n3164_1), .B(new_n3248), .Y(new_n4700));
  and_5  g02352(.A(new_n4700), .B(new_n4676), .Y(new_n4701));
  nand_5 g02353(.A(new_n4701), .B(new_n4699), .Y(new_n4702));
  not_8  g02354(.A(new_n4702), .Y(new_n4703));
  nand_5 g02355(.A(new_n4703), .B(new_n4697), .Y(new_n4704));
  nand_5 g02356(.A(new_n4704), .B(new_n4696), .Y(new_n4705));
  nand_5 g02357(.A(new_n4705), .B(new_n4690), .Y(new_n4706));
  nand_5 g02358(.A(new_n4706), .B(new_n4689), .Y(new_n4707));
  not_8  g02359(.A(new_n4707), .Y(new_n4708));
  nand_5 g02360(.A(new_n4664), .B(new_n4661), .Y(new_n4709));
  nand_5 g02361(.A(new_n4709), .B(new_n4666), .Y(new_n4710));
  or_5   g02362(.A(new_n4655), .B(n26748), .Y(new_n4711));
  xor_4  g02363(.A(new_n4711), .B(n21276), .Y(new_n4712));
  nand_5 g02364(.A(new_n4712), .B(n1204), .Y(new_n4713));
  or_5   g02365(.A(new_n4712), .B(n1204), .Y(new_n4714));
  nand_5 g02366(.A(new_n4714), .B(new_n4713), .Y(new_n4715));
  xor_4  g02367(.A(new_n4715), .B(new_n4710), .Y(new_n4716));
  not_8  g02368(.A(new_n4716), .Y(new_n4717));
  nand_5 g02369(.A(new_n4685), .B(new_n4678), .Y(new_n4718));
  nand_5 g02370(.A(new_n4718), .B(new_n4684), .Y(new_n4719));
  nor_5  g02371(.A(new_n4680), .B(n18558), .Y(new_n4720));
  not_8  g02372(.A(new_n4720), .Y(new_n4721));
  nand_5 g02373(.A(new_n4680), .B(n18558), .Y(new_n4722_1));
  and_5  g02374(.A(new_n4722_1), .B(new_n4721), .Y(new_n4723));
  not_8  g02375(.A(new_n4723), .Y(new_n4724));
  nand_5 g02376(.A(new_n4724), .B(new_n3084), .Y(new_n4725));
  nand_5 g02377(.A(new_n4723), .B(n10053), .Y(new_n4726));
  nand_5 g02378(.A(new_n4726), .B(new_n4725), .Y(new_n4727));
  xor_4  g02379(.A(new_n4727), .B(new_n4719), .Y(new_n4728));
  not_8  g02380(.A(new_n4728), .Y(new_n4729));
  nand_5 g02381(.A(new_n4729), .B(new_n4717), .Y(new_n4730));
  nand_5 g02382(.A(new_n4728), .B(new_n4716), .Y(new_n4731_1));
  nand_5 g02383(.A(new_n4731_1), .B(new_n4730), .Y(new_n4732));
  xor_4  g02384(.A(new_n4732), .B(new_n4708), .Y(new_n4733));
  not_8  g02385(.A(new_n4733), .Y(new_n4734));
  nand_5 g02386(.A(new_n4734), .B(new_n4651), .Y(new_n4735));
  not_8  g02387(.A(new_n4651), .Y(new_n4736));
  nand_5 g02388(.A(new_n4733), .B(new_n4736), .Y(new_n4737));
  nand_5 g02389(.A(new_n4690), .B(new_n4689), .Y(new_n4738));
  xor_4  g02390(.A(new_n4738), .B(new_n4705), .Y(new_n4739));
  nand_5 g02391(.A(new_n4630), .B(new_n4628), .Y(new_n4740));
  xor_4  g02392(.A(new_n4740), .B(new_n4637), .Y(new_n4741));
  not_8  g02393(.A(new_n4741), .Y(new_n4742));
  nand_5 g02394(.A(new_n4742), .B(new_n4739), .Y(new_n4743));
  or_5   g02395(.A(new_n4742), .B(new_n4739), .Y(new_n4744));
  and_5  g02396(.A(new_n4634), .B(new_n4633), .Y(new_n4745_1));
  xor_4  g02397(.A(new_n4745_1), .B(new_n4635), .Y(new_n4746));
  not_8  g02398(.A(new_n4692), .Y(new_n4747_1));
  nand_5 g02399(.A(new_n4694), .B(new_n4747_1), .Y(new_n4748));
  nand_5 g02400(.A(new_n4748), .B(new_n4696), .Y(new_n4749));
  xor_4  g02401(.A(new_n4749), .B(new_n4703), .Y(new_n4750));
  nand_5 g02402(.A(new_n4750), .B(new_n4746), .Y(new_n4751));
  or_5   g02403(.A(new_n4750), .B(new_n4746), .Y(new_n4752));
  nor_5  g02404(.A(new_n4701), .B(new_n4699), .Y(new_n4753));
  nor_5  g02405(.A(new_n4753), .B(new_n4703), .Y(new_n4754));
  nand_5 g02406(.A(new_n4149), .B(new_n4622), .Y(new_n4755));
  nand_5 g02407(.A(new_n4755), .B(new_n4635), .Y(new_n4756));
  not_8  g02408(.A(new_n4756), .Y(new_n4757));
  nand_5 g02409(.A(new_n4757), .B(new_n4754), .Y(new_n4758));
  nand_5 g02410(.A(new_n4758), .B(new_n4752), .Y(new_n4759));
  nand_5 g02411(.A(new_n4759), .B(new_n4751), .Y(new_n4760));
  nand_5 g02412(.A(new_n4760), .B(new_n4744), .Y(new_n4761));
  nand_5 g02413(.A(new_n4761), .B(new_n4743), .Y(new_n4762));
  nand_5 g02414(.A(new_n4762), .B(new_n4737), .Y(new_n4763));
  nand_5 g02415(.A(new_n4763), .B(new_n4735), .Y(new_n4764));
  nand_5 g02416(.A(new_n4649), .B(new_n4639), .Y(new_n4765));
  nand_5 g02417(.A(new_n4765), .B(new_n4647), .Y(new_n4766_1));
  not_8  g02418(.A(new_n4766_1), .Y(new_n4767));
  not_8  g02419(.A(n19905), .Y(new_n4768));
  not_8  g02420(.A(new_n4644), .Y(new_n4769));
  nand_5 g02421(.A(new_n4769), .B(new_n4768), .Y(new_n4770_1));
  nand_5 g02422(.A(new_n4644), .B(n19905), .Y(new_n4771));
  nand_5 g02423(.A(new_n4771), .B(new_n4770_1), .Y(new_n4772));
  nand_5 g02424(.A(new_n4772), .B(new_n4178), .Y(new_n4773));
  nor_5  g02425(.A(new_n4772), .B(new_n4178), .Y(new_n4774));
  not_8  g02426(.A(new_n4774), .Y(new_n4775));
  nand_5 g02427(.A(new_n4775), .B(new_n4773), .Y(new_n4776));
  xor_4  g02428(.A(new_n4776), .B(new_n4767), .Y(new_n4777_1));
  nand_5 g02429(.A(new_n4731_1), .B(new_n4708), .Y(new_n4778));
  nand_5 g02430(.A(new_n4778), .B(new_n4730), .Y(new_n4779));
  nand_5 g02431(.A(new_n4713), .B(new_n4710), .Y(new_n4780));
  nand_5 g02432(.A(new_n4780), .B(new_n4714), .Y(new_n4781));
  not_8  g02433(.A(n13668), .Y(new_n4782));
  nor_5  g02434(.A(new_n4711), .B(n21276), .Y(new_n4783));
  xor_4  g02435(.A(new_n4783), .B(new_n4782), .Y(new_n4784));
  or_5   g02436(.A(new_n4784), .B(n626), .Y(new_n4785_1));
  nand_5 g02437(.A(new_n4784), .B(n626), .Y(new_n4786));
  nand_5 g02438(.A(new_n4786), .B(new_n4785_1), .Y(new_n4787));
  xor_4  g02439(.A(new_n4787), .B(new_n4781), .Y(new_n4788));
  not_8  g02440(.A(new_n4788), .Y(new_n4789));
  nand_5 g02441(.A(new_n4726), .B(new_n4719), .Y(new_n4790));
  nand_5 g02442(.A(new_n4790), .B(new_n4725), .Y(new_n4791));
  not_8  g02443(.A(new_n4791), .Y(new_n4792));
  nand_5 g02444(.A(new_n4720), .B(new_n3002), .Y(new_n4793));
  nand_5 g02445(.A(new_n4721), .B(n3468), .Y(new_n4794));
  and_5  g02446(.A(new_n4794), .B(new_n4793), .Y(new_n4795));
  not_8  g02447(.A(new_n4795), .Y(new_n4796));
  nand_5 g02448(.A(new_n4796), .B(new_n3079), .Y(new_n4797));
  nand_5 g02449(.A(new_n4795), .B(n19514), .Y(new_n4798));
  nand_5 g02450(.A(new_n4798), .B(new_n4797), .Y(new_n4799));
  xor_4  g02451(.A(new_n4799), .B(new_n4792), .Y(new_n4800));
  nand_5 g02452(.A(new_n4800), .B(new_n4789), .Y(new_n4801));
  not_8  g02453(.A(new_n4800), .Y(new_n4802));
  nand_5 g02454(.A(new_n4802), .B(new_n4788), .Y(new_n4803));
  nand_5 g02455(.A(new_n4803), .B(new_n4801), .Y(new_n4804_1));
  xor_4  g02456(.A(new_n4804_1), .B(new_n4779), .Y(new_n4805));
  not_8  g02457(.A(new_n4805), .Y(new_n4806));
  nand_5 g02458(.A(new_n4806), .B(new_n4777_1), .Y(new_n4807));
  not_8  g02459(.A(new_n4777_1), .Y(new_n4808));
  nand_5 g02460(.A(new_n4805), .B(new_n4808), .Y(new_n4809));
  nand_5 g02461(.A(new_n4809), .B(new_n4807), .Y(new_n4810_1));
  xor_4  g02462(.A(new_n4810_1), .B(new_n4764), .Y(n266));
  nand_5 g02463(.A(new_n2782), .B(n21839), .Y(new_n4812_1));
  not_8  g02464(.A(n21839), .Y(new_n4813));
  nand_5 g02465(.A(n22270), .B(new_n4813), .Y(new_n4814_1));
  nand_5 g02466(.A(n27089), .B(new_n2786), .Y(new_n4815));
  nand_5 g02467(.A(new_n3296), .B(n8806), .Y(new_n4816));
  nand_5 g02468(.A(n11841), .B(new_n2791), .Y(new_n4817));
  nand_5 g02469(.A(new_n3194), .B(n2479), .Y(new_n4818));
  nand_5 g02470(.A(n10710), .B(new_n2797), .Y(new_n4819));
  nand_5 g02471(.A(new_n3108), .B(n9372), .Y(new_n4820));
  nand_5 g02472(.A(n20929), .B(new_n2803), .Y(new_n4821));
  nand_5 g02473(.A(new_n3072), .B(n6596), .Y(new_n4822));
  nand_5 g02474(.A(new_n2824), .B(n8006), .Y(new_n4823));
  nand_5 g02475(.A(n15289), .B(new_n3078), .Y(new_n4824));
  nand_5 g02476(.A(n25074), .B(new_n2804), .Y(new_n4825));
  nand_5 g02477(.A(new_n3136_1), .B(n6556), .Y(new_n4826));
  nand_5 g02478(.A(new_n2806), .B(n16396), .Y(new_n4827));
  nand_5 g02479(.A(n22871), .B(new_n3086), .Y(new_n4828));
  nand_5 g02480(.A(new_n2810), .B(n9399), .Y(new_n4829));
  nand_5 g02481(.A(n14275), .B(new_n3089_1), .Y(new_n4830));
  nand_5 g02482(.A(n25023), .B(new_n3163), .Y(new_n4831));
  nand_5 g02483(.A(new_n4831), .B(new_n4830), .Y(new_n4832));
  nand_5 g02484(.A(new_n4832), .B(new_n4829), .Y(new_n4833));
  nand_5 g02485(.A(new_n4833), .B(new_n4828), .Y(new_n4834));
  nand_5 g02486(.A(new_n4834), .B(new_n4827), .Y(new_n4835));
  nand_5 g02487(.A(new_n4835), .B(new_n4826), .Y(new_n4836));
  nand_5 g02488(.A(new_n4836), .B(new_n4825), .Y(new_n4837));
  nand_5 g02489(.A(new_n4837), .B(new_n4824), .Y(new_n4838));
  nand_5 g02490(.A(new_n4838), .B(new_n4823), .Y(new_n4839));
  nand_5 g02491(.A(new_n4839), .B(new_n4822), .Y(new_n4840));
  nand_5 g02492(.A(new_n4840), .B(new_n4821), .Y(new_n4841));
  nand_5 g02493(.A(new_n4841), .B(new_n4820), .Y(new_n4842));
  nand_5 g02494(.A(new_n4842), .B(new_n4819), .Y(new_n4843));
  nand_5 g02495(.A(new_n4843), .B(new_n4818), .Y(new_n4844));
  nand_5 g02496(.A(new_n4844), .B(new_n4817), .Y(new_n4845));
  nand_5 g02497(.A(new_n4845), .B(new_n4816), .Y(new_n4846));
  nand_5 g02498(.A(new_n4846), .B(new_n4815), .Y(new_n4847));
  nand_5 g02499(.A(new_n4847), .B(new_n4814_1), .Y(new_n4848));
  nand_5 g02500(.A(new_n4848), .B(new_n4812_1), .Y(new_n4849));
  not_8  g02501(.A(n23272), .Y(new_n4850_1));
  nand_5 g02502(.A(new_n4814_1), .B(new_n4812_1), .Y(new_n4851));
  xor_4  g02503(.A(new_n4851), .B(new_n4847), .Y(new_n4852));
  nand_5 g02504(.A(new_n4852), .B(new_n4850_1), .Y(new_n4853));
  not_8  g02505(.A(new_n4852), .Y(new_n4854));
  nand_5 g02506(.A(new_n4854), .B(n23272), .Y(new_n4855));
  not_8  g02507(.A(n11481), .Y(new_n4856));
  nand_5 g02508(.A(new_n4816), .B(new_n4815), .Y(new_n4857));
  xor_4  g02509(.A(new_n4857), .B(new_n4845), .Y(new_n4858_1));
  nand_5 g02510(.A(new_n4858_1), .B(new_n4856), .Y(new_n4859));
  not_8  g02511(.A(new_n4858_1), .Y(new_n4860));
  nand_5 g02512(.A(new_n4860), .B(n11481), .Y(new_n4861));
  not_8  g02513(.A(n16439), .Y(new_n4862));
  nand_5 g02514(.A(new_n4818), .B(new_n4817), .Y(new_n4863));
  xor_4  g02515(.A(new_n4863), .B(new_n4843), .Y(new_n4864));
  nand_5 g02516(.A(new_n4864), .B(new_n4862), .Y(new_n4865));
  not_8  g02517(.A(new_n4864), .Y(new_n4866));
  nand_5 g02518(.A(new_n4866), .B(n16439), .Y(new_n4867));
  not_8  g02519(.A(n15241), .Y(new_n4868));
  nand_5 g02520(.A(new_n4820), .B(new_n4819), .Y(new_n4869));
  xor_4  g02521(.A(new_n4869), .B(new_n4841), .Y(new_n4870));
  nand_5 g02522(.A(new_n4870), .B(new_n4868), .Y(new_n4871));
  not_8  g02523(.A(new_n4870), .Y(new_n4872));
  nand_5 g02524(.A(new_n4872), .B(n15241), .Y(new_n4873));
  not_8  g02525(.A(n7678), .Y(new_n4874));
  nand_5 g02526(.A(new_n4822), .B(new_n4821), .Y(new_n4875));
  xor_4  g02527(.A(new_n4875), .B(new_n4839), .Y(new_n4876));
  nand_5 g02528(.A(new_n4876), .B(new_n4874), .Y(new_n4877));
  not_8  g02529(.A(new_n4876), .Y(new_n4878));
  nand_5 g02530(.A(new_n4878), .B(n7678), .Y(new_n4879));
  not_8  g02531(.A(n3785), .Y(new_n4880));
  nand_5 g02532(.A(new_n4824), .B(new_n4823), .Y(new_n4881));
  xor_4  g02533(.A(new_n4881), .B(new_n4837), .Y(new_n4882));
  nand_5 g02534(.A(new_n4882), .B(new_n4880), .Y(new_n4883));
  not_8  g02535(.A(new_n4882), .Y(new_n4884));
  nand_5 g02536(.A(new_n4884), .B(n3785), .Y(new_n4885));
  not_8  g02537(.A(n20250), .Y(new_n4886));
  nand_5 g02538(.A(new_n4826), .B(new_n4825), .Y(new_n4887));
  xor_4  g02539(.A(new_n4887), .B(new_n4835), .Y(new_n4888));
  nand_5 g02540(.A(new_n4888), .B(new_n4886), .Y(new_n4889));
  not_8  g02541(.A(new_n4888), .Y(new_n4890));
  nand_5 g02542(.A(new_n4890), .B(n20250), .Y(new_n4891_1));
  not_8  g02543(.A(n5822), .Y(new_n4892));
  nand_5 g02544(.A(new_n4828), .B(new_n4827), .Y(new_n4893));
  xor_4  g02545(.A(new_n4893), .B(new_n4833), .Y(new_n4894));
  nand_5 g02546(.A(new_n4894), .B(new_n4892), .Y(new_n4895));
  not_8  g02547(.A(new_n4894), .Y(new_n4896));
  nand_5 g02548(.A(new_n4896), .B(n5822), .Y(new_n4897));
  not_8  g02549(.A(n26443), .Y(new_n4898));
  and_5  g02550(.A(new_n4830), .B(new_n4829), .Y(new_n4899));
  xor_4  g02551(.A(new_n4899), .B(new_n4831), .Y(new_n4900));
  not_8  g02552(.A(new_n4900), .Y(new_n4901));
  nand_5 g02553(.A(new_n4901), .B(new_n4898), .Y(new_n4902));
  nand_5 g02554(.A(new_n4900), .B(n26443), .Y(new_n4903));
  or_5   g02555(.A(n25023), .B(new_n3163), .Y(new_n4904));
  and_5  g02556(.A(new_n4904), .B(new_n4831), .Y(new_n4905));
  not_8  g02557(.A(new_n4905), .Y(new_n4906));
  nand_5 g02558(.A(new_n4906), .B(n1681), .Y(new_n4907));
  nand_5 g02559(.A(new_n4907), .B(new_n4903), .Y(new_n4908));
  nand_5 g02560(.A(new_n4908), .B(new_n4902), .Y(new_n4909));
  nand_5 g02561(.A(new_n4909), .B(new_n4897), .Y(new_n4910));
  nand_5 g02562(.A(new_n4910), .B(new_n4895), .Y(new_n4911));
  nand_5 g02563(.A(new_n4911), .B(new_n4891_1), .Y(new_n4912));
  nand_5 g02564(.A(new_n4912), .B(new_n4889), .Y(new_n4913_1));
  nand_5 g02565(.A(new_n4913_1), .B(new_n4885), .Y(new_n4914));
  nand_5 g02566(.A(new_n4914), .B(new_n4883), .Y(new_n4915));
  nand_5 g02567(.A(new_n4915), .B(new_n4879), .Y(new_n4916));
  nand_5 g02568(.A(new_n4916), .B(new_n4877), .Y(new_n4917));
  nand_5 g02569(.A(new_n4917), .B(new_n4873), .Y(new_n4918));
  nand_5 g02570(.A(new_n4918), .B(new_n4871), .Y(new_n4919));
  nand_5 g02571(.A(new_n4919), .B(new_n4867), .Y(new_n4920));
  nand_5 g02572(.A(new_n4920), .B(new_n4865), .Y(new_n4921));
  nand_5 g02573(.A(new_n4921), .B(new_n4861), .Y(new_n4922));
  nand_5 g02574(.A(new_n4922), .B(new_n4859), .Y(new_n4923));
  nand_5 g02575(.A(new_n4923), .B(new_n4855), .Y(new_n4924));
  nand_5 g02576(.A(new_n4924), .B(new_n4853), .Y(new_n4925_1));
  nor_5  g02577(.A(new_n4925_1), .B(new_n4849), .Y(new_n4926));
  not_8  g02578(.A(new_n4926), .Y(new_n4927));
  not_8  g02579(.A(n24196), .Y(new_n4928));
  not_8  g02580(.A(n25381), .Y(new_n4929));
  not_8  g02581(.A(n268), .Y(new_n4930));
  not_8  g02582(.A(n24032), .Y(new_n4931));
  nand_5 g02583(.A(new_n4931), .B(new_n2622), .Y(new_n4932));
  or_5   g02584(.A(new_n4932), .B(n6785), .Y(new_n4933));
  nor_5  g02585(.A(new_n4933), .B(n24879), .Y(new_n4934));
  nand_5 g02586(.A(new_n4934), .B(new_n4930), .Y(new_n4935));
  nor_5  g02587(.A(new_n4935), .B(n12587), .Y(new_n4936));
  nand_5 g02588(.A(new_n4936), .B(new_n4929), .Y(new_n4937));
  nor_5  g02589(.A(new_n4937), .B(n16376), .Y(new_n4938));
  nand_5 g02590(.A(new_n4938), .B(new_n4928), .Y(new_n4939_1));
  nor_5  g02591(.A(new_n4939_1), .B(n18105), .Y(new_n4940));
  not_8  g02592(.A(new_n4940), .Y(new_n4941));
  not_8  g02593(.A(n25475), .Y(new_n4942));
  nand_5 g02594(.A(new_n4494), .B(new_n2657), .Y(new_n4943));
  nor_5  g02595(.A(new_n4943), .B(n25168), .Y(new_n4944));
  xor_4  g02596(.A(new_n4944), .B(n1999), .Y(new_n4945));
  nand_5 g02597(.A(new_n4945), .B(new_n4942), .Y(new_n4946));
  nor_5  g02598(.A(new_n4945), .B(new_n4942), .Y(new_n4947_1));
  not_8  g02599(.A(new_n4947_1), .Y(new_n4948));
  xor_4  g02600(.A(new_n4943), .B(n25168), .Y(new_n4949));
  or_5   g02601(.A(new_n4949), .B(n23849), .Y(new_n4950));
  nand_5 g02602(.A(new_n4949), .B(n23849), .Y(new_n4951));
  not_8  g02603(.A(n12446), .Y(new_n4952_1));
  nand_5 g02604(.A(new_n4495), .B(n9318), .Y(new_n4953));
  nand_5 g02605(.A(new_n4953), .B(new_n4943), .Y(new_n4954));
  nand_5 g02606(.A(new_n4954), .B(new_n4952_1), .Y(new_n4955));
  nor_5  g02607(.A(new_n4954), .B(new_n4952_1), .Y(new_n4956));
  not_8  g02608(.A(new_n4956), .Y(new_n4957_1));
  nand_5 g02609(.A(new_n4499), .B(new_n4491), .Y(new_n4958));
  nand_5 g02610(.A(new_n4958), .B(new_n4498), .Y(new_n4959));
  nand_5 g02611(.A(new_n4959), .B(new_n4957_1), .Y(new_n4960));
  nand_5 g02612(.A(new_n4960), .B(new_n4955), .Y(new_n4961));
  nand_5 g02613(.A(new_n4961), .B(new_n4951), .Y(new_n4962));
  nand_5 g02614(.A(new_n4962), .B(new_n4950), .Y(new_n4963));
  nand_5 g02615(.A(new_n4963), .B(new_n4948), .Y(new_n4964_1));
  nand_5 g02616(.A(new_n4964_1), .B(new_n4946), .Y(new_n4965));
  not_8  g02617(.A(n18880), .Y(new_n4966_1));
  nand_5 g02618(.A(new_n4944), .B(new_n2651), .Y(new_n4967_1));
  not_8  g02619(.A(new_n4967_1), .Y(new_n4968));
  nand_5 g02620(.A(new_n4968), .B(new_n2647), .Y(new_n4969));
  nand_5 g02621(.A(new_n4967_1), .B(n9396), .Y(new_n4970));
  nand_5 g02622(.A(new_n4970), .B(new_n4969), .Y(new_n4971));
  nand_5 g02623(.A(new_n4971), .B(new_n4966_1), .Y(new_n4972_1));
  not_8  g02624(.A(new_n4972_1), .Y(new_n4973));
  nor_5  g02625(.A(new_n4973), .B(new_n4965), .Y(new_n4974));
  nor_5  g02626(.A(new_n4971), .B(new_n4966_1), .Y(new_n4975));
  not_8  g02627(.A(new_n4975), .Y(new_n4976));
  nand_5 g02628(.A(new_n4976), .B(new_n4969), .Y(new_n4977));
  nor_5  g02629(.A(new_n4977), .B(new_n4974), .Y(new_n4978));
  not_8  g02630(.A(new_n4978), .Y(new_n4979));
  nand_5 g02631(.A(new_n4979), .B(new_n4941), .Y(new_n4980));
  nand_5 g02632(.A(new_n4939_1), .B(n18105), .Y(new_n4981));
  and_5  g02633(.A(new_n4981), .B(new_n4941), .Y(new_n4982));
  nand_5 g02634(.A(new_n4976), .B(new_n4972_1), .Y(new_n4983));
  xor_4  g02635(.A(new_n4983), .B(new_n4965), .Y(new_n4984));
  or_5   g02636(.A(new_n4984), .B(new_n4982), .Y(new_n4985));
  nand_5 g02637(.A(new_n4984), .B(new_n4982), .Y(new_n4986));
  xor_4  g02638(.A(new_n4938), .B(new_n4928), .Y(new_n4987));
  nand_5 g02639(.A(new_n4948), .B(new_n4946), .Y(new_n4988));
  xor_4  g02640(.A(new_n4988), .B(new_n4963), .Y(new_n4989));
  or_5   g02641(.A(new_n4989), .B(new_n4987), .Y(new_n4990));
  nand_5 g02642(.A(new_n4989), .B(new_n4987), .Y(new_n4991));
  xor_4  g02643(.A(new_n4937), .B(n16376), .Y(new_n4992));
  nand_5 g02644(.A(new_n4951), .B(new_n4950), .Y(new_n4993));
  xor_4  g02645(.A(new_n4993), .B(new_n4961), .Y(new_n4994));
  or_5   g02646(.A(new_n4994), .B(new_n4992), .Y(new_n4995));
  nand_5 g02647(.A(new_n4994), .B(new_n4992), .Y(new_n4996));
  xor_4  g02648(.A(new_n4936), .B(new_n4929), .Y(new_n4997));
  nand_5 g02649(.A(new_n4957_1), .B(new_n4955), .Y(new_n4998));
  xor_4  g02650(.A(new_n4998), .B(new_n4959), .Y(new_n4999));
  or_5   g02651(.A(new_n4999), .B(new_n4997), .Y(new_n5000));
  nand_5 g02652(.A(new_n4999), .B(new_n4997), .Y(new_n5001));
  xor_4  g02653(.A(new_n4935), .B(n12587), .Y(new_n5002));
  or_5   g02654(.A(new_n5002), .B(new_n4503), .Y(new_n5003));
  nand_5 g02655(.A(new_n5002), .B(new_n4503), .Y(new_n5004));
  xor_4  g02656(.A(new_n4934), .B(new_n4930), .Y(new_n5005));
  or_5   g02657(.A(new_n5005), .B(new_n4371), .Y(new_n5006));
  nand_5 g02658(.A(new_n5005), .B(new_n4371), .Y(new_n5007));
  xor_4  g02659(.A(new_n4933), .B(n24879), .Y(new_n5008));
  or_5   g02660(.A(new_n5008), .B(new_n4338), .Y(new_n5009));
  nand_5 g02661(.A(new_n5008), .B(new_n4338), .Y(new_n5010));
  nand_5 g02662(.A(new_n4932), .B(n6785), .Y(new_n5011_1));
  and_5  g02663(.A(new_n5011_1), .B(new_n4933), .Y(new_n5012));
  or_5   g02664(.A(new_n5012), .B(new_n4342), .Y(new_n5013));
  nand_5 g02665(.A(new_n5012), .B(new_n4342), .Y(new_n5014));
  nand_5 g02666(.A(n24032), .B(n22843), .Y(new_n5015));
  and_5  g02667(.A(new_n5015), .B(new_n4932), .Y(new_n5016));
  or_5   g02668(.A(new_n5016), .B(new_n4351), .Y(new_n5017));
  nand_5 g02669(.A(new_n5016), .B(new_n4351), .Y(new_n5018));
  nand_5 g02670(.A(new_n2634), .B(n22843), .Y(new_n5019));
  nand_5 g02671(.A(new_n5019), .B(new_n5018), .Y(new_n5020_1));
  nand_5 g02672(.A(new_n5020_1), .B(new_n5017), .Y(new_n5021));
  nand_5 g02673(.A(new_n5021), .B(new_n5014), .Y(new_n5022));
  nand_5 g02674(.A(new_n5022), .B(new_n5013), .Y(new_n5023));
  nand_5 g02675(.A(new_n5023), .B(new_n5010), .Y(new_n5024_1));
  nand_5 g02676(.A(new_n5024_1), .B(new_n5009), .Y(new_n5025_1));
  nand_5 g02677(.A(new_n5025_1), .B(new_n5007), .Y(new_n5026_1));
  nand_5 g02678(.A(new_n5026_1), .B(new_n5006), .Y(new_n5027));
  nand_5 g02679(.A(new_n5027), .B(new_n5004), .Y(new_n5028));
  nand_5 g02680(.A(new_n5028), .B(new_n5003), .Y(new_n5029));
  nand_5 g02681(.A(new_n5029), .B(new_n5001), .Y(new_n5030));
  nand_5 g02682(.A(new_n5030), .B(new_n5000), .Y(new_n5031_1));
  nand_5 g02683(.A(new_n5031_1), .B(new_n4996), .Y(new_n5032));
  nand_5 g02684(.A(new_n5032), .B(new_n4995), .Y(new_n5033));
  nand_5 g02685(.A(new_n5033), .B(new_n4991), .Y(new_n5034));
  nand_5 g02686(.A(new_n5034), .B(new_n4990), .Y(new_n5035));
  nand_5 g02687(.A(new_n5035), .B(new_n4986), .Y(new_n5036));
  nand_5 g02688(.A(new_n5036), .B(new_n4985), .Y(new_n5037));
  not_8  g02689(.A(new_n5037), .Y(new_n5038));
  nor_5  g02690(.A(new_n5038), .B(new_n4980), .Y(new_n5039));
  nor_5  g02691(.A(new_n5039), .B(new_n4927), .Y(new_n5040));
  and_5  g02692(.A(new_n5039), .B(new_n4927), .Y(new_n5041));
  nor_5  g02693(.A(new_n5041), .B(new_n5040), .Y(new_n5042));
  nand_5 g02694(.A(new_n4925_1), .B(new_n4849), .Y(new_n5043));
  and_5  g02695(.A(new_n5043), .B(new_n4927), .Y(new_n5044));
  nand_5 g02696(.A(new_n4978), .B(new_n4940), .Y(new_n5045));
  nand_5 g02697(.A(new_n5045), .B(new_n4980), .Y(new_n5046_1));
  xor_4  g02698(.A(new_n5046_1), .B(new_n5038), .Y(new_n5047));
  nand_5 g02699(.A(new_n5047), .B(new_n5044), .Y(new_n5048));
  nor_5  g02700(.A(new_n5047), .B(new_n5044), .Y(new_n5049));
  not_8  g02701(.A(new_n5049), .Y(new_n5050));
  nand_5 g02702(.A(new_n4855), .B(new_n4853), .Y(new_n5051));
  xor_4  g02703(.A(new_n5051), .B(new_n4923), .Y(new_n5052));
  nand_5 g02704(.A(new_n4986), .B(new_n4985), .Y(new_n5053));
  xor_4  g02705(.A(new_n5053), .B(new_n5035), .Y(new_n5054));
  nand_5 g02706(.A(new_n5054), .B(new_n5052), .Y(new_n5055));
  nor_5  g02707(.A(new_n5054), .B(new_n5052), .Y(new_n5056));
  not_8  g02708(.A(new_n5056), .Y(new_n5057));
  nand_5 g02709(.A(new_n4861), .B(new_n4859), .Y(new_n5058));
  xor_4  g02710(.A(new_n5058), .B(new_n4921), .Y(new_n5059));
  nand_5 g02711(.A(new_n4991), .B(new_n4990), .Y(new_n5060_1));
  xor_4  g02712(.A(new_n5060_1), .B(new_n5033), .Y(new_n5061));
  nand_5 g02713(.A(new_n5061), .B(new_n5059), .Y(new_n5062_1));
  nor_5  g02714(.A(new_n5061), .B(new_n5059), .Y(new_n5063));
  not_8  g02715(.A(new_n5063), .Y(new_n5064_1));
  nand_5 g02716(.A(new_n4867), .B(new_n4865), .Y(new_n5065));
  xor_4  g02717(.A(new_n5065), .B(new_n4919), .Y(new_n5066));
  nand_5 g02718(.A(new_n4996), .B(new_n4995), .Y(new_n5067));
  xor_4  g02719(.A(new_n5067), .B(new_n5031_1), .Y(new_n5068));
  nand_5 g02720(.A(new_n5068), .B(new_n5066), .Y(new_n5069));
  nor_5  g02721(.A(new_n5068), .B(new_n5066), .Y(new_n5070));
  not_8  g02722(.A(new_n5070), .Y(new_n5071));
  nand_5 g02723(.A(new_n4873), .B(new_n4871), .Y(new_n5072));
  xor_4  g02724(.A(new_n5072), .B(new_n4917), .Y(new_n5073));
  nand_5 g02725(.A(new_n5001), .B(new_n5000), .Y(new_n5074));
  xor_4  g02726(.A(new_n5074), .B(new_n5029), .Y(new_n5075));
  nand_5 g02727(.A(new_n5075), .B(new_n5073), .Y(new_n5076));
  or_5   g02728(.A(new_n5075), .B(new_n5073), .Y(new_n5077_1));
  nand_5 g02729(.A(new_n4879), .B(new_n4877), .Y(new_n5078));
  xor_4  g02730(.A(new_n5078), .B(new_n4915), .Y(new_n5079));
  nand_5 g02731(.A(new_n5004), .B(new_n5003), .Y(new_n5080));
  xor_4  g02732(.A(new_n5080), .B(new_n5027), .Y(new_n5081));
  nand_5 g02733(.A(new_n5081), .B(new_n5079), .Y(new_n5082_1));
  or_5   g02734(.A(new_n5081), .B(new_n5079), .Y(new_n5083));
  nand_5 g02735(.A(new_n4885), .B(new_n4883), .Y(new_n5084));
  xor_4  g02736(.A(new_n5084), .B(new_n4913_1), .Y(new_n5085));
  nand_5 g02737(.A(new_n5007), .B(new_n5006), .Y(new_n5086));
  xor_4  g02738(.A(new_n5086), .B(new_n5025_1), .Y(new_n5087));
  nand_5 g02739(.A(new_n5087), .B(new_n5085), .Y(new_n5088));
  or_5   g02740(.A(new_n5087), .B(new_n5085), .Y(new_n5089));
  nand_5 g02741(.A(new_n4891_1), .B(new_n4889), .Y(new_n5090));
  xor_4  g02742(.A(new_n5090), .B(new_n4911), .Y(new_n5091));
  nand_5 g02743(.A(new_n5010), .B(new_n5009), .Y(new_n5092));
  xor_4  g02744(.A(new_n5092), .B(new_n5023), .Y(new_n5093));
  nand_5 g02745(.A(new_n5093), .B(new_n5091), .Y(new_n5094));
  or_5   g02746(.A(new_n5093), .B(new_n5091), .Y(new_n5095));
  nand_5 g02747(.A(new_n4897), .B(new_n4895), .Y(new_n5096));
  xor_4  g02748(.A(new_n5096), .B(new_n4909), .Y(new_n5097));
  nand_5 g02749(.A(new_n5014), .B(new_n5013), .Y(new_n5098_1));
  xor_4  g02750(.A(new_n5098_1), .B(new_n5021), .Y(new_n5099));
  nand_5 g02751(.A(new_n5099), .B(new_n5097), .Y(new_n5100));
  or_5   g02752(.A(new_n5099), .B(new_n5097), .Y(new_n5101_1));
  nand_5 g02753(.A(new_n5018), .B(new_n5017), .Y(new_n5102));
  xor_4  g02754(.A(new_n5102), .B(new_n5019), .Y(new_n5103));
  nand_5 g02755(.A(new_n4903), .B(new_n4902), .Y(new_n5104));
  xor_4  g02756(.A(new_n5104), .B(new_n4907), .Y(new_n5105));
  or_5   g02757(.A(new_n5105), .B(new_n5103), .Y(new_n5106));
  nand_5 g02758(.A(new_n5105), .B(new_n5103), .Y(new_n5107));
  not_8  g02759(.A(new_n2634), .Y(new_n5108));
  nand_5 g02760(.A(new_n5108), .B(new_n2622), .Y(new_n5109));
  nand_5 g02761(.A(new_n5109), .B(new_n5019), .Y(new_n5110));
  nand_5 g02762(.A(new_n4905), .B(new_n2613), .Y(new_n5111));
  nand_5 g02763(.A(new_n5111), .B(new_n4907), .Y(new_n5112));
  or_5   g02764(.A(new_n5112), .B(new_n5110), .Y(new_n5113));
  nand_5 g02765(.A(new_n5113), .B(new_n5107), .Y(new_n5114));
  and_5  g02766(.A(new_n5114), .B(new_n5106), .Y(new_n5115_1));
  nand_5 g02767(.A(new_n5115_1), .B(new_n5101_1), .Y(new_n5116));
  nand_5 g02768(.A(new_n5116), .B(new_n5100), .Y(new_n5117));
  nand_5 g02769(.A(new_n5117), .B(new_n5095), .Y(new_n5118));
  nand_5 g02770(.A(new_n5118), .B(new_n5094), .Y(new_n5119));
  nand_5 g02771(.A(new_n5119), .B(new_n5089), .Y(new_n5120_1));
  nand_5 g02772(.A(new_n5120_1), .B(new_n5088), .Y(new_n5121));
  nand_5 g02773(.A(new_n5121), .B(new_n5083), .Y(new_n5122));
  nand_5 g02774(.A(new_n5122), .B(new_n5082_1), .Y(new_n5123));
  nand_5 g02775(.A(new_n5123), .B(new_n5077_1), .Y(new_n5124));
  nand_5 g02776(.A(new_n5124), .B(new_n5076), .Y(new_n5125));
  nand_5 g02777(.A(new_n5125), .B(new_n5071), .Y(new_n5126));
  nand_5 g02778(.A(new_n5126), .B(new_n5069), .Y(new_n5127));
  nand_5 g02779(.A(new_n5127), .B(new_n5064_1), .Y(new_n5128_1));
  nand_5 g02780(.A(new_n5128_1), .B(new_n5062_1), .Y(new_n5129));
  nand_5 g02781(.A(new_n5129), .B(new_n5057), .Y(new_n5130));
  nand_5 g02782(.A(new_n5130), .B(new_n5055), .Y(new_n5131_1));
  nand_5 g02783(.A(new_n5131_1), .B(new_n5050), .Y(new_n5132));
  nand_5 g02784(.A(new_n5132), .B(new_n5048), .Y(new_n5133));
  not_8  g02785(.A(new_n5133), .Y(new_n5134));
  xor_4  g02786(.A(new_n5134), .B(new_n5042), .Y(n298));
  not_8  g02787(.A(n20455), .Y(new_n5136));
  nand_5 g02788(.A(new_n5136), .B(n5376), .Y(new_n5137));
  not_8  g02789(.A(n5376), .Y(new_n5138));
  nand_5 g02790(.A(n20455), .B(new_n5138), .Y(new_n5139));
  not_8  g02791(.A(n1639), .Y(new_n5140_1));
  nand_5 g02792(.A(n5128), .B(new_n5140_1), .Y(new_n5141));
  not_8  g02793(.A(n5128), .Y(new_n5142));
  nand_5 g02794(.A(new_n5142), .B(n1639), .Y(new_n5143));
  not_8  g02795(.A(n23120), .Y(new_n5144));
  nand_5 g02796(.A(new_n5144), .B(n16968), .Y(new_n5145));
  nand_5 g02797(.A(new_n5145), .B(new_n5143), .Y(new_n5146));
  nand_5 g02798(.A(new_n5146), .B(new_n5141), .Y(new_n5147));
  nand_5 g02799(.A(new_n5147), .B(new_n5139), .Y(new_n5148));
  nand_5 g02800(.A(new_n5148), .B(new_n5137), .Y(new_n5149));
  not_8  g02801(.A(n13263), .Y(new_n5150));
  nand_5 g02802(.A(n21779), .B(new_n5150), .Y(new_n5151));
  or_5   g02803(.A(n21779), .B(new_n5150), .Y(new_n5152));
  nand_5 g02804(.A(new_n5152), .B(new_n5151), .Y(new_n5153));
  xor_4  g02805(.A(new_n5153), .B(new_n5149), .Y(new_n5154));
  not_8  g02806(.A(n196), .Y(new_n5155));
  or_5   g02807(.A(n9460), .B(new_n5155), .Y(new_n5156));
  nand_5 g02808(.A(n9460), .B(new_n5155), .Y(new_n5157));
  not_8  g02809(.A(n11749), .Y(new_n5158_1));
  or_5   g02810(.A(n14954), .B(new_n5158_1), .Y(new_n5159));
  nand_5 g02811(.A(n14954), .B(new_n5158_1), .Y(new_n5160));
  not_8  g02812(.A(n13424), .Y(new_n5161));
  nand_5 g02813(.A(n23831), .B(new_n5161), .Y(new_n5162));
  nand_5 g02814(.A(new_n5162), .B(new_n5160), .Y(new_n5163));
  nand_5 g02815(.A(new_n5163), .B(new_n5159), .Y(new_n5164));
  nand_5 g02816(.A(new_n5164), .B(new_n5157), .Y(new_n5165));
  nand_5 g02817(.A(new_n5165), .B(new_n5156), .Y(new_n5166));
  not_8  g02818(.A(n7460), .Y(new_n5167));
  or_5   g02819(.A(n22068), .B(new_n5167), .Y(new_n5168_1));
  nand_5 g02820(.A(n22068), .B(new_n5167), .Y(new_n5169));
  nand_5 g02821(.A(new_n5169), .B(new_n5168_1), .Y(new_n5170));
  xor_4  g02822(.A(new_n5170), .B(new_n5166), .Y(new_n5171));
  nand_5 g02823(.A(new_n5171), .B(new_n5154), .Y(new_n5172));
  not_8  g02824(.A(new_n5154), .Y(new_n5173));
  not_8  g02825(.A(new_n5171), .Y(new_n5174));
  nand_5 g02826(.A(new_n5174), .B(new_n5173), .Y(new_n5175));
  nand_5 g02827(.A(new_n5139), .B(new_n5137), .Y(new_n5176));
  xor_4  g02828(.A(new_n5176), .B(new_n5147), .Y(new_n5177));
  nand_5 g02829(.A(new_n5157), .B(new_n5156), .Y(new_n5178));
  xor_4  g02830(.A(new_n5178), .B(new_n5164), .Y(new_n5179));
  nand_5 g02831(.A(new_n5179), .B(new_n5177), .Y(new_n5180));
  or_5   g02832(.A(new_n5179), .B(new_n5177), .Y(new_n5181));
  and_5  g02833(.A(new_n5143), .B(new_n5141), .Y(new_n5182));
  xor_4  g02834(.A(new_n5182), .B(new_n5145), .Y(new_n5183));
  not_8  g02835(.A(new_n5183), .Y(new_n5184_1));
  and_5  g02836(.A(new_n5160), .B(new_n5159), .Y(new_n5185));
  xor_4  g02837(.A(new_n5185), .B(new_n5162), .Y(new_n5186));
  not_8  g02838(.A(new_n5186), .Y(new_n5187));
  nand_5 g02839(.A(new_n5187), .B(new_n5184_1), .Y(new_n5188));
  nand_5 g02840(.A(new_n5186), .B(new_n5183), .Y(new_n5189));
  nand_5 g02841(.A(n23120), .B(new_n3960), .Y(new_n5190));
  and_5  g02842(.A(new_n5190), .B(new_n5145), .Y(new_n5191));
  not_8  g02843(.A(new_n5191), .Y(new_n5192));
  xor_4  g02844(.A(n23831), .B(new_n5161), .Y(new_n5193));
  not_8  g02845(.A(new_n5193), .Y(new_n5194));
  nand_5 g02846(.A(new_n5194), .B(new_n5192), .Y(new_n5195));
  nand_5 g02847(.A(new_n5195), .B(new_n5189), .Y(new_n5196));
  nand_5 g02848(.A(new_n5196), .B(new_n5188), .Y(new_n5197));
  nand_5 g02849(.A(new_n5197), .B(new_n5181), .Y(new_n5198));
  nand_5 g02850(.A(new_n5198), .B(new_n5180), .Y(new_n5199));
  nand_5 g02851(.A(new_n5199), .B(new_n5175), .Y(new_n5200));
  nand_5 g02852(.A(new_n5200), .B(new_n5172), .Y(new_n5201));
  nand_5 g02853(.A(new_n5152), .B(new_n5149), .Y(new_n5202));
  nand_5 g02854(.A(new_n5202), .B(new_n5151), .Y(new_n5203));
  not_8  g02855(.A(n14510), .Y(new_n5204));
  nand_5 g02856(.A(n16988), .B(new_n5204), .Y(new_n5205));
  or_5   g02857(.A(n16988), .B(new_n5204), .Y(new_n5206));
  nand_5 g02858(.A(new_n5206), .B(new_n5205), .Y(new_n5207));
  xor_4  g02859(.A(new_n5207), .B(new_n5203), .Y(new_n5208));
  nand_5 g02860(.A(new_n5169), .B(new_n5166), .Y(new_n5209));
  nand_5 g02861(.A(new_n5209), .B(new_n5168_1), .Y(new_n5210));
  not_8  g02862(.A(n6971), .Y(new_n5211_1));
  nand_5 g02863(.A(n24319), .B(new_n5211_1), .Y(new_n5212));
  nor_5  g02864(.A(n24319), .B(new_n5211_1), .Y(new_n5213_1));
  not_8  g02865(.A(new_n5213_1), .Y(new_n5214));
  nand_5 g02866(.A(new_n5214), .B(new_n5212), .Y(new_n5215));
  xor_4  g02867(.A(new_n5215), .B(new_n5210), .Y(new_n5216));
  nand_5 g02868(.A(new_n5216), .B(new_n5208), .Y(new_n5217));
  not_8  g02869(.A(new_n5208), .Y(new_n5218));
  not_8  g02870(.A(new_n5216), .Y(new_n5219));
  nand_5 g02871(.A(new_n5219), .B(new_n5218), .Y(new_n5220));
  nand_5 g02872(.A(new_n5220), .B(new_n5217), .Y(new_n5221));
  xor_4  g02873(.A(new_n5221), .B(new_n5201), .Y(new_n5222));
  not_8  g02874(.A(new_n5222), .Y(new_n5223));
  not_8  g02875(.A(n5752), .Y(new_n5224));
  nand_5 g02876(.A(n14071), .B(new_n5224), .Y(new_n5225));
  not_8  g02877(.A(n14071), .Y(new_n5226_1));
  nand_5 g02878(.A(new_n5226_1), .B(n5752), .Y(new_n5227));
  not_8  g02879(.A(n18171), .Y(new_n5228_1));
  nand_5 g02880(.A(new_n5228_1), .B(n1738), .Y(new_n5229));
  not_8  g02881(.A(n1738), .Y(new_n5230));
  nand_5 g02882(.A(n18171), .B(new_n5230), .Y(new_n5231));
  not_8  g02883(.A(n25073), .Y(new_n5232));
  nand_5 g02884(.A(new_n5232), .B(n12152), .Y(new_n5233));
  not_8  g02885(.A(n12152), .Y(new_n5234));
  nand_5 g02886(.A(n25073), .B(new_n5234), .Y(new_n5235));
  not_8  g02887(.A(n19107), .Y(new_n5236));
  nand_5 g02888(.A(n22309), .B(new_n5236), .Y(new_n5237));
  nand_5 g02889(.A(new_n5237), .B(new_n5235), .Y(new_n5238));
  nand_5 g02890(.A(new_n5238), .B(new_n5233), .Y(new_n5239));
  nand_5 g02891(.A(new_n5239), .B(new_n5231), .Y(new_n5240));
  nand_5 g02892(.A(new_n5240), .B(new_n5229), .Y(new_n5241));
  nand_5 g02893(.A(new_n5241), .B(new_n5227), .Y(new_n5242));
  nand_5 g02894(.A(new_n5242), .B(new_n5225), .Y(new_n5243));
  not_8  g02895(.A(n16158), .Y(new_n5244));
  nand_5 g02896(.A(n24085), .B(new_n5244), .Y(new_n5245));
  not_8  g02897(.A(n24085), .Y(new_n5246));
  nand_5 g02898(.A(new_n5246), .B(n16158), .Y(new_n5247));
  nand_5 g02899(.A(new_n5247), .B(new_n5245), .Y(new_n5248));
  xor_4  g02900(.A(new_n5248), .B(new_n5243), .Y(new_n5249));
  or_5   g02901(.A(new_n5249), .B(new_n5223), .Y(new_n5250));
  nand_5 g02902(.A(new_n5249), .B(new_n5223), .Y(new_n5251));
  nand_5 g02903(.A(new_n5172), .B(new_n5175), .Y(new_n5252));
  xor_4  g02904(.A(new_n5252), .B(new_n5199), .Y(new_n5253));
  not_8  g02905(.A(new_n5253), .Y(new_n5254));
  nand_5 g02906(.A(new_n5227), .B(new_n5225), .Y(new_n5255_1));
  xor_4  g02907(.A(new_n5255_1), .B(new_n5241), .Y(new_n5256_1));
  or_5   g02908(.A(new_n5256_1), .B(new_n5254), .Y(new_n5257));
  nand_5 g02909(.A(new_n5256_1), .B(new_n5254), .Y(new_n5258));
  nand_5 g02910(.A(new_n5181), .B(new_n5180), .Y(new_n5259));
  xor_4  g02911(.A(new_n5259), .B(new_n5197), .Y(new_n5260));
  not_8  g02912(.A(new_n5260), .Y(new_n5261));
  nand_5 g02913(.A(new_n5231), .B(new_n5229), .Y(new_n5262));
  xor_4  g02914(.A(new_n5262), .B(new_n5239), .Y(new_n5263));
  or_5   g02915(.A(new_n5263), .B(new_n5261), .Y(new_n5264));
  nand_5 g02916(.A(new_n5263), .B(new_n5261), .Y(new_n5265_1));
  xor_4  g02917(.A(new_n5193), .B(new_n5191), .Y(new_n5266));
  xor_4  g02918(.A(n22309), .B(new_n5236), .Y(new_n5267));
  not_8  g02919(.A(new_n5267), .Y(new_n5268));
  nand_5 g02920(.A(new_n5268), .B(new_n5266), .Y(new_n5269));
  not_8  g02921(.A(new_n5269), .Y(new_n5270));
  nand_5 g02922(.A(new_n5235), .B(new_n5233), .Y(new_n5271));
  xnor_4 g02923(.A(new_n5271), .B(new_n5237), .Y(new_n5272));
  nand_5 g02924(.A(new_n5272), .B(new_n5270), .Y(new_n5273_1));
  not_8  g02925(.A(new_n5273_1), .Y(new_n5274_1));
  nand_5 g02926(.A(new_n5189), .B(new_n5188), .Y(new_n5275));
  xor_4  g02927(.A(new_n5275), .B(new_n5195), .Y(new_n5276));
  not_8  g02928(.A(new_n5276), .Y(new_n5277));
  nor_5  g02929(.A(new_n5272), .B(new_n5270), .Y(new_n5278));
  nor_5  g02930(.A(new_n5278), .B(new_n5277), .Y(new_n5279));
  nor_5  g02931(.A(new_n5279), .B(new_n5274_1), .Y(new_n5280));
  not_8  g02932(.A(new_n5280), .Y(new_n5281));
  nand_5 g02933(.A(new_n5281), .B(new_n5265_1), .Y(new_n5282));
  nand_5 g02934(.A(new_n5282), .B(new_n5264), .Y(new_n5283));
  nand_5 g02935(.A(new_n5283), .B(new_n5258), .Y(new_n5284));
  nand_5 g02936(.A(new_n5284), .B(new_n5257), .Y(new_n5285));
  nand_5 g02937(.A(new_n5285), .B(new_n5251), .Y(new_n5286));
  nand_5 g02938(.A(new_n5286), .B(new_n5250), .Y(new_n5287));
  nand_5 g02939(.A(new_n5220), .B(new_n5201), .Y(new_n5288));
  nand_5 g02940(.A(new_n5288), .B(new_n5217), .Y(new_n5289));
  nand_5 g02941(.A(new_n5206), .B(new_n5203), .Y(new_n5290));
  nand_5 g02942(.A(new_n5290), .B(new_n5205), .Y(new_n5291));
  not_8  g02943(.A(new_n5291), .Y(new_n5292));
  not_8  g02944(.A(n4119), .Y(new_n5293));
  nand_5 g02945(.A(new_n5293), .B(n1525), .Y(new_n5294));
  or_5   g02946(.A(new_n5293), .B(n1525), .Y(new_n5295));
  nand_5 g02947(.A(new_n5295), .B(new_n5294), .Y(new_n5296));
  xor_4  g02948(.A(new_n5296), .B(new_n5292), .Y(new_n5297));
  not_8  g02949(.A(new_n5297), .Y(new_n5298));
  nand_5 g02950(.A(new_n5214), .B(new_n5210), .Y(new_n5299));
  nand_5 g02951(.A(new_n5299), .B(new_n5212), .Y(new_n5300_1));
  not_8  g02952(.A(new_n5300_1), .Y(new_n5301));
  not_8  g02953(.A(n4272), .Y(new_n5302_1));
  nand_5 g02954(.A(n12626), .B(new_n5302_1), .Y(new_n5303));
  nor_5  g02955(.A(n12626), .B(new_n5302_1), .Y(new_n5304));
  not_8  g02956(.A(new_n5304), .Y(new_n5305));
  nand_5 g02957(.A(new_n5305), .B(new_n5303), .Y(new_n5306));
  xor_4  g02958(.A(new_n5306), .B(new_n5301), .Y(new_n5307));
  not_8  g02959(.A(new_n5307), .Y(new_n5308));
  nand_5 g02960(.A(new_n5308), .B(new_n5298), .Y(new_n5309));
  nand_5 g02961(.A(new_n5307), .B(new_n5297), .Y(new_n5310));
  nand_5 g02962(.A(new_n5310), .B(new_n5309), .Y(new_n5311));
  xor_4  g02963(.A(new_n5311), .B(new_n5289), .Y(new_n5312));
  nand_5 g02964(.A(new_n5247), .B(new_n5243), .Y(new_n5313));
  nand_5 g02965(.A(new_n5313), .B(new_n5245), .Y(new_n5314));
  not_8  g02966(.A(n20604), .Y(new_n5315));
  nand_5 g02967(.A(n21735), .B(new_n5315), .Y(new_n5316));
  not_8  g02968(.A(n21735), .Y(new_n5317));
  nand_5 g02969(.A(new_n5317), .B(n20604), .Y(new_n5318));
  nand_5 g02970(.A(new_n5318), .B(new_n5316), .Y(new_n5319));
  xnor_4 g02971(.A(new_n5319), .B(new_n5314), .Y(new_n5320));
  nand_5 g02972(.A(new_n5320), .B(new_n5312), .Y(new_n5321));
  not_8  g02973(.A(new_n5321), .Y(new_n5322));
  nor_5  g02974(.A(new_n5320), .B(new_n5312), .Y(new_n5323));
  nor_5  g02975(.A(new_n5323), .B(new_n5322), .Y(new_n5324));
  xor_4  g02976(.A(new_n5324), .B(new_n5287), .Y(n317));
  not_8  g02977(.A(n9934), .Y(new_n5326));
  nand_5 g02978(.A(new_n5326), .B(new_n3711), .Y(new_n5327));
  nand_5 g02979(.A(n9934), .B(n3506), .Y(new_n5328));
  nand_5 g02980(.A(new_n4160), .B(new_n3740_1), .Y(new_n5329));
  nand_5 g02981(.A(n26553), .B(n10096), .Y(new_n5330_1));
  not_8  g02982(.A(n4964), .Y(new_n5331));
  nand_5 g02983(.A(new_n3744), .B(new_n5331), .Y(new_n5332));
  nand_5 g02984(.A(n16994), .B(n4964), .Y(new_n5333));
  nand_5 g02985(.A(n9246), .B(n7876), .Y(new_n5334));
  nand_5 g02986(.A(new_n5334), .B(new_n5333), .Y(new_n5335));
  nand_5 g02987(.A(new_n5335), .B(new_n5332), .Y(new_n5336));
  nand_5 g02988(.A(new_n5336), .B(new_n5330_1), .Y(new_n5337_1));
  nand_5 g02989(.A(new_n5337_1), .B(new_n5329), .Y(new_n5338));
  nand_5 g02990(.A(new_n5338), .B(new_n4146_1), .Y(new_n5339));
  not_8  g02991(.A(new_n5339), .Y(new_n5340));
  nor_5  g02992(.A(new_n5338), .B(new_n4146_1), .Y(new_n5341));
  nor_5  g02993(.A(new_n5341), .B(n14790), .Y(new_n5342));
  nor_5  g02994(.A(new_n5342), .B(new_n5340), .Y(new_n5343));
  or_5   g02995(.A(new_n5343), .B(n17251), .Y(new_n5344));
  nand_5 g02996(.A(new_n5343), .B(n17251), .Y(new_n5345));
  nand_5 g02997(.A(new_n5345), .B(new_n4177), .Y(new_n5346));
  nand_5 g02998(.A(new_n5346), .B(new_n5344), .Y(new_n5347));
  nand_5 g02999(.A(new_n5347), .B(new_n3728), .Y(new_n5348));
  not_8  g03000(.A(new_n5348), .Y(new_n5349));
  nor_5  g03001(.A(new_n5347), .B(new_n3728), .Y(new_n5350));
  nor_5  g03002(.A(new_n5350), .B(n22597), .Y(new_n5351_1));
  nor_5  g03003(.A(new_n5351_1), .B(new_n5349), .Y(new_n5352));
  or_5   g03004(.A(new_n5352), .B(n19327), .Y(new_n5353_1));
  nand_5 g03005(.A(new_n5352), .B(n19327), .Y(new_n5354));
  nand_5 g03006(.A(new_n5354), .B(new_n3724), .Y(new_n5355));
  nand_5 g03007(.A(new_n5355), .B(new_n5353_1), .Y(new_n5356));
  nand_5 g03008(.A(new_n5356), .B(new_n3720), .Y(new_n5357));
  not_8  g03009(.A(new_n5357), .Y(new_n5358));
  nor_5  g03010(.A(new_n5356), .B(new_n3720), .Y(new_n5359));
  nor_5  g03011(.A(new_n5359), .B(n26224), .Y(new_n5360));
  nor_5  g03012(.A(new_n5360), .B(new_n5358), .Y(new_n5361));
  or_5   g03013(.A(new_n5361), .B(n14899), .Y(new_n5362));
  not_8  g03014(.A(n18496), .Y(new_n5363));
  nand_5 g03015(.A(new_n5361), .B(n14899), .Y(new_n5364));
  nand_5 g03016(.A(new_n5364), .B(new_n5363), .Y(new_n5365));
  nand_5 g03017(.A(new_n5365), .B(new_n5362), .Y(new_n5366));
  nand_5 g03018(.A(new_n5366), .B(new_n5328), .Y(new_n5367));
  nand_5 g03019(.A(new_n5367), .B(new_n5327), .Y(new_n5368));
  not_8  g03020(.A(n2979), .Y(new_n5369));
  not_8  g03021(.A(n647), .Y(new_n5370));
  not_8  g03022(.A(n26408), .Y(new_n5371));
  nand_5 g03023(.A(new_n5371), .B(new_n5370), .Y(new_n5372));
  nand_5 g03024(.A(n26408), .B(n647), .Y(new_n5373));
  not_8  g03025(.A(n18227), .Y(new_n5374));
  not_8  g03026(.A(n20409), .Y(new_n5375));
  nand_5 g03027(.A(new_n5375), .B(new_n5374), .Y(new_n5376_1));
  nand_5 g03028(.A(n20409), .B(n18227), .Y(new_n5377));
  not_8  g03029(.A(n7377), .Y(new_n5378));
  nand_5 g03030(.A(new_n4293), .B(new_n5378), .Y(new_n5379));
  nand_5 g03031(.A(n25749), .B(n7377), .Y(new_n5380));
  not_8  g03032(.A(n11630), .Y(new_n5381));
  nand_5 g03033(.A(new_n5381), .B(new_n4219), .Y(new_n5382));
  nand_5 g03034(.A(n11630), .B(n3161), .Y(new_n5383));
  not_8  g03035(.A(n9003), .Y(new_n5384));
  not_8  g03036(.A(n13453), .Y(new_n5385));
  nand_5 g03037(.A(new_n5385), .B(new_n5384), .Y(new_n5386_1));
  nand_5 g03038(.A(n13453), .B(n9003), .Y(new_n5387));
  not_8  g03039(.A(n7421), .Y(new_n5388));
  nand_5 g03040(.A(new_n5388), .B(new_n4189), .Y(new_n5389));
  nand_5 g03041(.A(n7421), .B(n4957), .Y(new_n5390));
  not_8  g03042(.A(n19680), .Y(new_n5391));
  nand_5 g03043(.A(new_n5391), .B(new_n4195), .Y(new_n5392));
  nand_5 g03044(.A(n19680), .B(n7524), .Y(new_n5393));
  not_8  g03045(.A(n2809), .Y(new_n5394));
  nand_5 g03046(.A(new_n4201), .B(new_n5394), .Y(new_n5395));
  nand_5 g03047(.A(n15743), .B(n2809), .Y(new_n5396));
  nand_5 g03048(.A(n20658), .B(n15508), .Y(new_n5397));
  nand_5 g03049(.A(new_n5397), .B(new_n5396), .Y(new_n5398));
  nand_5 g03050(.A(new_n5398), .B(new_n5395), .Y(new_n5399_1));
  nand_5 g03051(.A(new_n5399_1), .B(new_n5393), .Y(new_n5400_1));
  nand_5 g03052(.A(new_n5400_1), .B(new_n5392), .Y(new_n5401));
  nand_5 g03053(.A(new_n5401), .B(new_n5390), .Y(new_n5402));
  nand_5 g03054(.A(new_n5402), .B(new_n5389), .Y(new_n5403_1));
  nand_5 g03055(.A(new_n5403_1), .B(new_n5387), .Y(new_n5404));
  nand_5 g03056(.A(new_n5404), .B(new_n5386_1), .Y(new_n5405));
  nand_5 g03057(.A(new_n5405), .B(new_n5383), .Y(new_n5406));
  nand_5 g03058(.A(new_n5406), .B(new_n5382), .Y(new_n5407));
  nand_5 g03059(.A(new_n5407), .B(new_n5380), .Y(new_n5408));
  nand_5 g03060(.A(new_n5408), .B(new_n5379), .Y(new_n5409));
  nand_5 g03061(.A(new_n5409), .B(new_n5377), .Y(new_n5410));
  nand_5 g03062(.A(new_n5410), .B(new_n5376_1), .Y(new_n5411));
  nand_5 g03063(.A(new_n5411), .B(new_n5373), .Y(new_n5412));
  nand_5 g03064(.A(new_n5412), .B(new_n5372), .Y(new_n5413));
  nand_5 g03065(.A(new_n5413), .B(new_n5369), .Y(new_n5414));
  not_8  g03066(.A(new_n5414), .Y(new_n5415));
  nor_5  g03067(.A(new_n5413), .B(new_n5369), .Y(new_n5416));
  nor_5  g03068(.A(new_n5416), .B(n9554), .Y(new_n5417));
  nor_5  g03069(.A(new_n5417), .B(new_n5415), .Y(new_n5418));
  not_8  g03070(.A(n9259), .Y(new_n5419));
  not_8  g03071(.A(n9554), .Y(new_n5420));
  nor_5  g03072(.A(new_n5416), .B(new_n5415), .Y(new_n5421));
  xor_4  g03073(.A(new_n5421), .B(new_n5420), .Y(new_n5422));
  nand_5 g03074(.A(new_n5422), .B(new_n5419), .Y(new_n5423));
  not_8  g03075(.A(new_n5422), .Y(new_n5424));
  nand_5 g03076(.A(new_n5424), .B(n9259), .Y(new_n5425));
  nand_5 g03077(.A(new_n5373), .B(new_n5372), .Y(new_n5426));
  xor_4  g03078(.A(new_n5426), .B(new_n5411), .Y(new_n5427));
  not_8  g03079(.A(new_n5427), .Y(new_n5428));
  nand_5 g03080(.A(new_n5428), .B(new_n3694), .Y(new_n5429));
  nand_5 g03081(.A(new_n5427), .B(n21489), .Y(new_n5430_1));
  nand_5 g03082(.A(new_n5377), .B(new_n5376_1), .Y(new_n5431));
  xor_4  g03083(.A(new_n5431), .B(new_n5409), .Y(new_n5432));
  not_8  g03084(.A(new_n5432), .Y(new_n5433));
  nand_5 g03085(.A(new_n5433), .B(new_n3778), .Y(new_n5434));
  nand_5 g03086(.A(new_n5432), .B(n20213), .Y(new_n5435));
  nand_5 g03087(.A(new_n5380), .B(new_n5379), .Y(new_n5436));
  xor_4  g03088(.A(new_n5436), .B(new_n5407), .Y(new_n5437));
  not_8  g03089(.A(new_n5437), .Y(new_n5438_1));
  nand_5 g03090(.A(new_n5438_1), .B(new_n3695), .Y(new_n5439_1));
  nand_5 g03091(.A(new_n5437), .B(n13912), .Y(new_n5440));
  nand_5 g03092(.A(new_n5383), .B(new_n5382), .Y(new_n5441));
  xor_4  g03093(.A(new_n5441), .B(new_n5405), .Y(new_n5442));
  not_8  g03094(.A(new_n5442), .Y(new_n5443_1));
  nand_5 g03095(.A(new_n5443_1), .B(new_n3793), .Y(new_n5444));
  nand_5 g03096(.A(new_n5442), .B(n7670), .Y(new_n5445));
  nand_5 g03097(.A(new_n5387), .B(new_n5386_1), .Y(new_n5446));
  xor_4  g03098(.A(new_n5446), .B(new_n5403_1), .Y(new_n5447));
  not_8  g03099(.A(new_n5447), .Y(new_n5448));
  nand_5 g03100(.A(new_n5448), .B(new_n3696), .Y(new_n5449));
  nand_5 g03101(.A(new_n5447), .B(n9598), .Y(new_n5450));
  not_8  g03102(.A(n22290), .Y(new_n5451_1));
  nand_5 g03103(.A(new_n5390), .B(new_n5389), .Y(new_n5452));
  xor_4  g03104(.A(new_n5452), .B(new_n5401), .Y(new_n5453));
  not_8  g03105(.A(new_n5453), .Y(new_n5454));
  nand_5 g03106(.A(new_n5454), .B(new_n5451_1), .Y(new_n5455));
  nand_5 g03107(.A(new_n5453), .B(n22290), .Y(new_n5456));
  not_8  g03108(.A(n11273), .Y(new_n5457));
  nand_5 g03109(.A(new_n5393), .B(new_n5392), .Y(new_n5458));
  xor_4  g03110(.A(new_n5458), .B(new_n5399_1), .Y(new_n5459));
  not_8  g03111(.A(new_n5459), .Y(new_n5460));
  nand_5 g03112(.A(new_n5460), .B(new_n5457), .Y(new_n5461));
  nand_5 g03113(.A(new_n5459), .B(n11273), .Y(new_n5462));
  nand_5 g03114(.A(new_n5396), .B(new_n5395), .Y(new_n5463));
  xor_4  g03115(.A(new_n5463), .B(new_n5397), .Y(new_n5464));
  not_8  g03116(.A(new_n5464), .Y(new_n5465));
  nand_5 g03117(.A(new_n5465), .B(new_n3698), .Y(new_n5466));
  nand_5 g03118(.A(new_n5464), .B(n25565), .Y(new_n5467));
  not_8  g03119(.A(n15508), .Y(new_n5468));
  not_8  g03120(.A(n20658), .Y(new_n5469));
  nand_5 g03121(.A(new_n5469), .B(new_n5468), .Y(new_n5470));
  and_5  g03122(.A(new_n5470), .B(new_n5397), .Y(new_n5471));
  nand_5 g03123(.A(new_n5471), .B(n21993), .Y(new_n5472_1));
  nand_5 g03124(.A(new_n5472_1), .B(new_n5467), .Y(new_n5473));
  nand_5 g03125(.A(new_n5473), .B(new_n5466), .Y(new_n5474));
  nand_5 g03126(.A(new_n5474), .B(new_n5462), .Y(new_n5475));
  nand_5 g03127(.A(new_n5475), .B(new_n5461), .Y(new_n5476));
  nand_5 g03128(.A(new_n5476), .B(new_n5456), .Y(new_n5477));
  nand_5 g03129(.A(new_n5477), .B(new_n5455), .Y(new_n5478));
  nand_5 g03130(.A(new_n5478), .B(new_n5450), .Y(new_n5479));
  nand_5 g03131(.A(new_n5479), .B(new_n5449), .Y(new_n5480));
  nand_5 g03132(.A(new_n5480), .B(new_n5445), .Y(new_n5481));
  nand_5 g03133(.A(new_n5481), .B(new_n5444), .Y(new_n5482));
  nand_5 g03134(.A(new_n5482), .B(new_n5440), .Y(new_n5483));
  nand_5 g03135(.A(new_n5483), .B(new_n5439_1), .Y(new_n5484));
  nand_5 g03136(.A(new_n5484), .B(new_n5435), .Y(new_n5485_1));
  nand_5 g03137(.A(new_n5485_1), .B(new_n5434), .Y(new_n5486));
  nand_5 g03138(.A(new_n5486), .B(new_n5430_1), .Y(new_n5487));
  nand_5 g03139(.A(new_n5487), .B(new_n5429), .Y(new_n5488));
  nand_5 g03140(.A(new_n5488), .B(new_n5425), .Y(new_n5489));
  nand_5 g03141(.A(new_n5489), .B(new_n5423), .Y(new_n5490));
  not_8  g03142(.A(new_n5490), .Y(new_n5491));
  nand_5 g03143(.A(new_n5491), .B(new_n5418), .Y(new_n5492));
  not_8  g03144(.A(new_n5418), .Y(new_n5493));
  nand_5 g03145(.A(new_n5490), .B(new_n5493), .Y(new_n5494));
  nand_5 g03146(.A(new_n5494), .B(new_n5492), .Y(new_n5495));
  not_8  g03147(.A(n3740), .Y(new_n5496));
  nand_5 g03148(.A(new_n5423), .B(new_n5425), .Y(new_n5497));
  xor_4  g03149(.A(new_n5497), .B(new_n5488), .Y(new_n5498));
  nand_5 g03150(.A(new_n5498), .B(new_n5496), .Y(new_n5499));
  not_8  g03151(.A(new_n5498), .Y(new_n5500));
  nand_5 g03152(.A(new_n5500), .B(n3740), .Y(new_n5501));
  not_8  g03153(.A(n2858), .Y(new_n5502));
  nand_5 g03154(.A(new_n5429), .B(new_n5430_1), .Y(new_n5503));
  xor_4  g03155(.A(new_n5503), .B(new_n5486), .Y(new_n5504));
  nand_5 g03156(.A(new_n5504), .B(new_n5502), .Y(new_n5505));
  not_8  g03157(.A(new_n5504), .Y(new_n5506));
  nand_5 g03158(.A(new_n5506), .B(n2858), .Y(new_n5507));
  not_8  g03159(.A(n2659), .Y(new_n5508));
  nand_5 g03160(.A(new_n5434), .B(new_n5435), .Y(new_n5509));
  xor_4  g03161(.A(new_n5509), .B(new_n5484), .Y(new_n5510));
  nand_5 g03162(.A(new_n5510), .B(new_n5508), .Y(new_n5511));
  not_8  g03163(.A(new_n5510), .Y(new_n5512));
  nand_5 g03164(.A(new_n5512), .B(n2659), .Y(new_n5513));
  not_8  g03165(.A(n24327), .Y(new_n5514));
  nand_5 g03166(.A(new_n5439_1), .B(new_n5440), .Y(new_n5515));
  xor_4  g03167(.A(new_n5515), .B(new_n5482), .Y(new_n5516));
  nand_5 g03168(.A(new_n5516), .B(new_n5514), .Y(new_n5517_1));
  not_8  g03169(.A(new_n5516), .Y(new_n5518));
  nand_5 g03170(.A(new_n5518), .B(n24327), .Y(new_n5519));
  not_8  g03171(.A(n22198), .Y(new_n5520));
  nand_5 g03172(.A(new_n5444), .B(new_n5445), .Y(new_n5521_1));
  xor_4  g03173(.A(new_n5521_1), .B(new_n5480), .Y(new_n5522));
  nand_5 g03174(.A(new_n5522), .B(new_n5520), .Y(new_n5523));
  not_8  g03175(.A(new_n5522), .Y(new_n5524_1));
  nand_5 g03176(.A(new_n5524_1), .B(n22198), .Y(new_n5525));
  not_8  g03177(.A(n20826), .Y(new_n5526));
  nand_5 g03178(.A(new_n5449), .B(new_n5450), .Y(new_n5527));
  xor_4  g03179(.A(new_n5527), .B(new_n5478), .Y(new_n5528));
  nand_5 g03180(.A(new_n5528), .B(new_n5526), .Y(new_n5529));
  not_8  g03181(.A(new_n5528), .Y(new_n5530));
  nand_5 g03182(.A(new_n5530), .B(n20826), .Y(new_n5531));
  not_8  g03183(.A(n7305), .Y(new_n5532_1));
  nand_5 g03184(.A(new_n5455), .B(new_n5456), .Y(new_n5533));
  xor_4  g03185(.A(new_n5533), .B(new_n5476), .Y(new_n5534));
  nand_5 g03186(.A(new_n5534), .B(new_n5532_1), .Y(new_n5535));
  not_8  g03187(.A(new_n5534), .Y(new_n5536));
  nand_5 g03188(.A(new_n5536), .B(n7305), .Y(new_n5537));
  not_8  g03189(.A(n25872), .Y(new_n5538));
  nand_5 g03190(.A(new_n5461), .B(new_n5462), .Y(new_n5539));
  xor_4  g03191(.A(new_n5539), .B(new_n5474), .Y(new_n5540));
  nand_5 g03192(.A(new_n5540), .B(new_n5538), .Y(new_n5541));
  not_8  g03193(.A(new_n5540), .Y(new_n5542));
  nand_5 g03194(.A(new_n5542), .B(n25872), .Y(new_n5543));
  not_8  g03195(.A(n20259), .Y(new_n5544));
  nand_5 g03196(.A(new_n5466), .B(new_n5467), .Y(new_n5545));
  xor_4  g03197(.A(new_n5545), .B(new_n5472_1), .Y(new_n5546));
  or_5   g03198(.A(new_n5546), .B(new_n5544), .Y(new_n5547));
  nand_5 g03199(.A(new_n5546), .B(new_n5544), .Y(new_n5548));
  not_8  g03200(.A(n3925), .Y(new_n5549));
  xor_4  g03201(.A(new_n5471), .B(n21993), .Y(new_n5550));
  nand_5 g03202(.A(new_n5550), .B(new_n5549), .Y(new_n5551));
  nand_5 g03203(.A(new_n5551), .B(new_n5548), .Y(new_n5552));
  nand_5 g03204(.A(new_n5552), .B(new_n5547), .Y(new_n5553));
  not_8  g03205(.A(new_n5553), .Y(new_n5554));
  nand_5 g03206(.A(new_n5554), .B(new_n5543), .Y(new_n5555));
  nand_5 g03207(.A(new_n5555), .B(new_n5541), .Y(new_n5556));
  nand_5 g03208(.A(new_n5556), .B(new_n5537), .Y(new_n5557));
  nand_5 g03209(.A(new_n5557), .B(new_n5535), .Y(new_n5558));
  nand_5 g03210(.A(new_n5558), .B(new_n5531), .Y(new_n5559));
  nand_5 g03211(.A(new_n5559), .B(new_n5529), .Y(new_n5560));
  nand_5 g03212(.A(new_n5560), .B(new_n5525), .Y(new_n5561));
  nand_5 g03213(.A(new_n5561), .B(new_n5523), .Y(new_n5562));
  nand_5 g03214(.A(new_n5562), .B(new_n5519), .Y(new_n5563));
  nand_5 g03215(.A(new_n5563), .B(new_n5517_1), .Y(new_n5564_1));
  nand_5 g03216(.A(new_n5564_1), .B(new_n5513), .Y(new_n5565));
  nand_5 g03217(.A(new_n5565), .B(new_n5511), .Y(new_n5566));
  nand_5 g03218(.A(new_n5566), .B(new_n5507), .Y(new_n5567));
  nand_5 g03219(.A(new_n5567), .B(new_n5505), .Y(new_n5568));
  nand_5 g03220(.A(new_n5568), .B(new_n5501), .Y(new_n5569));
  nand_5 g03221(.A(new_n5569), .B(new_n5499), .Y(new_n5570));
  xor_4  g03222(.A(new_n5570), .B(new_n5495), .Y(new_n5571));
  or_5   g03223(.A(new_n5571), .B(new_n5368), .Y(new_n5572));
  nand_5 g03224(.A(new_n5571), .B(new_n5368), .Y(new_n5573));
  nand_5 g03225(.A(new_n5573), .B(new_n5572), .Y(new_n5574));
  nand_5 g03226(.A(new_n5328), .B(new_n5327), .Y(new_n5575));
  xor_4  g03227(.A(new_n5575), .B(new_n5366), .Y(new_n5576));
  nand_5 g03228(.A(new_n5499), .B(new_n5501), .Y(new_n5577));
  xor_4  g03229(.A(new_n5577), .B(new_n5568), .Y(new_n5578));
  or_5   g03230(.A(new_n5578), .B(new_n5576), .Y(new_n5579_1));
  nand_5 g03231(.A(new_n5578), .B(new_n5576), .Y(new_n5580));
  and_5  g03232(.A(new_n5364), .B(new_n5362), .Y(new_n5581));
  xor_4  g03233(.A(new_n5581), .B(new_n5363), .Y(new_n5582));
  not_8  g03234(.A(new_n5582), .Y(new_n5583));
  nand_5 g03235(.A(new_n5505), .B(new_n5507), .Y(new_n5584));
  xor_4  g03236(.A(new_n5584), .B(new_n5566), .Y(new_n5585));
  or_5   g03237(.A(new_n5585), .B(new_n5583), .Y(new_n5586));
  nand_5 g03238(.A(new_n5585), .B(new_n5583), .Y(new_n5587));
  not_8  g03239(.A(n26224), .Y(new_n5588));
  nor_5  g03240(.A(new_n5359), .B(new_n5358), .Y(new_n5589));
  xor_4  g03241(.A(new_n5589), .B(new_n5588), .Y(new_n5590));
  not_8  g03242(.A(new_n5590), .Y(new_n5591));
  nand_5 g03243(.A(new_n5511), .B(new_n5513), .Y(new_n5592));
  xor_4  g03244(.A(new_n5592), .B(new_n5564_1), .Y(new_n5593_1));
  or_5   g03245(.A(new_n5593_1), .B(new_n5591), .Y(new_n5594));
  nand_5 g03246(.A(new_n5593_1), .B(new_n5591), .Y(new_n5595));
  and_5  g03247(.A(new_n5354), .B(new_n5353_1), .Y(new_n5596));
  xor_4  g03248(.A(new_n5596), .B(new_n3724), .Y(new_n5597));
  not_8  g03249(.A(new_n5597), .Y(new_n5598));
  nand_5 g03250(.A(new_n5517_1), .B(new_n5519), .Y(new_n5599));
  xor_4  g03251(.A(new_n5599), .B(new_n5562), .Y(new_n5600));
  or_5   g03252(.A(new_n5600), .B(new_n5598), .Y(new_n5601));
  nand_5 g03253(.A(new_n5600), .B(new_n5598), .Y(new_n5602));
  nor_5  g03254(.A(new_n5350), .B(new_n5349), .Y(new_n5603_1));
  xor_4  g03255(.A(new_n5603_1), .B(new_n4222), .Y(new_n5604));
  not_8  g03256(.A(new_n5604), .Y(new_n5605_1));
  nand_5 g03257(.A(new_n5523), .B(new_n5525), .Y(new_n5606));
  xor_4  g03258(.A(new_n5606), .B(new_n5560), .Y(new_n5607));
  or_5   g03259(.A(new_n5607), .B(new_n5605_1), .Y(new_n5608));
  nand_5 g03260(.A(new_n5607), .B(new_n5605_1), .Y(new_n5609_1));
  and_5  g03261(.A(new_n5345), .B(new_n5344), .Y(new_n5610));
  xor_4  g03262(.A(new_n5610), .B(new_n4177), .Y(new_n5611));
  not_8  g03263(.A(new_n5611), .Y(new_n5612));
  nand_5 g03264(.A(new_n5529), .B(new_n5531), .Y(new_n5613));
  xor_4  g03265(.A(new_n5613), .B(new_n5558), .Y(new_n5614));
  or_5   g03266(.A(new_n5614), .B(new_n5612), .Y(new_n5615));
  nand_5 g03267(.A(new_n5614), .B(new_n5612), .Y(new_n5616));
  nor_5  g03268(.A(new_n5341), .B(new_n5340), .Y(new_n5617));
  xor_4  g03269(.A(new_n5617), .B(new_n3736), .Y(new_n5618));
  not_8  g03270(.A(new_n5618), .Y(new_n5619));
  nand_5 g03271(.A(new_n5535), .B(new_n5537), .Y(new_n5620));
  xor_4  g03272(.A(new_n5620), .B(new_n5556), .Y(new_n5621));
  or_5   g03273(.A(new_n5621), .B(new_n5619), .Y(new_n5622));
  nand_5 g03274(.A(new_n5621), .B(new_n5619), .Y(new_n5623));
  nand_5 g03275(.A(new_n5330_1), .B(new_n5329), .Y(new_n5624));
  xor_4  g03276(.A(new_n5624), .B(new_n5336), .Y(new_n5625));
  nand_5 g03277(.A(new_n5541), .B(new_n5543), .Y(new_n5626));
  xor_4  g03278(.A(new_n5626), .B(new_n5554), .Y(new_n5627));
  or_5   g03279(.A(new_n5627), .B(new_n5625), .Y(new_n5628));
  nand_5 g03280(.A(new_n5627), .B(new_n5625), .Y(new_n5629));
  xor_4  g03281(.A(new_n5550), .B(n3925), .Y(new_n5630));
  nand_5 g03282(.A(new_n3827), .B(new_n4207), .Y(new_n5631));
  nand_5 g03283(.A(new_n5631), .B(new_n5334), .Y(new_n5632));
  not_8  g03284(.A(new_n5632), .Y(new_n5633));
  nand_5 g03285(.A(new_n5633), .B(new_n5630), .Y(new_n5634_1));
  not_8  g03286(.A(new_n5634_1), .Y(new_n5635));
  nand_5 g03287(.A(new_n5333), .B(new_n5332), .Y(new_n5636));
  not_8  g03288(.A(new_n5636), .Y(new_n5637));
  nand_5 g03289(.A(new_n5637), .B(new_n5635), .Y(new_n5638));
  xor_4  g03290(.A(new_n5637), .B(new_n5334), .Y(new_n5639));
  nand_5 g03291(.A(new_n5639), .B(new_n5634_1), .Y(new_n5640));
  nand_5 g03292(.A(new_n5548), .B(new_n5547), .Y(new_n5641));
  xnor_4 g03293(.A(new_n5641), .B(new_n5551), .Y(new_n5642));
  nand_5 g03294(.A(new_n5642), .B(new_n5640), .Y(new_n5643_1));
  nand_5 g03295(.A(new_n5643_1), .B(new_n5638), .Y(new_n5644));
  not_8  g03296(.A(new_n5644), .Y(new_n5645));
  nand_5 g03297(.A(new_n5645), .B(new_n5629), .Y(new_n5646));
  nand_5 g03298(.A(new_n5646), .B(new_n5628), .Y(new_n5647));
  nand_5 g03299(.A(new_n5647), .B(new_n5623), .Y(new_n5648));
  nand_5 g03300(.A(new_n5648), .B(new_n5622), .Y(new_n5649));
  nand_5 g03301(.A(new_n5649), .B(new_n5616), .Y(new_n5650));
  nand_5 g03302(.A(new_n5650), .B(new_n5615), .Y(new_n5651));
  nand_5 g03303(.A(new_n5651), .B(new_n5609_1), .Y(new_n5652));
  nand_5 g03304(.A(new_n5652), .B(new_n5608), .Y(new_n5653));
  nand_5 g03305(.A(new_n5653), .B(new_n5602), .Y(new_n5654));
  nand_5 g03306(.A(new_n5654), .B(new_n5601), .Y(new_n5655));
  nand_5 g03307(.A(new_n5655), .B(new_n5595), .Y(new_n5656));
  nand_5 g03308(.A(new_n5656), .B(new_n5594), .Y(new_n5657));
  nand_5 g03309(.A(new_n5657), .B(new_n5587), .Y(new_n5658));
  nand_5 g03310(.A(new_n5658), .B(new_n5586), .Y(new_n5659));
  nand_5 g03311(.A(new_n5659), .B(new_n5580), .Y(new_n5660));
  nand_5 g03312(.A(new_n5660), .B(new_n5579_1), .Y(new_n5661));
  xor_4  g03313(.A(new_n5661), .B(new_n5574), .Y(n332));
  nand_5 g03314(.A(n15780), .B(n2387), .Y(new_n5663));
  nand_5 g03315(.A(new_n2504), .B(new_n3051), .Y(new_n5664));
  nand_5 g03316(.A(n19494), .B(n6502), .Y(new_n5665));
  nand_5 g03317(.A(new_n5665), .B(new_n5664), .Y(new_n5666));
  xnor_4 g03318(.A(new_n5666), .B(new_n5663), .Y(new_n5667));
  not_8  g03319(.A(new_n5667), .Y(new_n5668));
  not_8  g03320(.A(n12495), .Y(new_n5669));
  nand_5 g03321(.A(new_n3159), .B(new_n2506), .Y(new_n5670));
  and_5  g03322(.A(new_n5670), .B(new_n5663), .Y(new_n5671));
  nand_5 g03323(.A(new_n5671), .B(new_n5669), .Y(new_n5672));
  or_5   g03324(.A(new_n5672), .B(n20235), .Y(new_n5673));
  nand_5 g03325(.A(new_n5672), .B(n20235), .Y(new_n5674));
  nand_5 g03326(.A(new_n5674), .B(new_n5673), .Y(new_n5675));
  xor_4  g03327(.A(new_n5675), .B(new_n5668), .Y(new_n5676));
  not_8  g03328(.A(new_n5676), .Y(new_n5677));
  not_8  g03329(.A(n21654), .Y(new_n5678));
  nand_5 g03330(.A(new_n5678), .B(n16502), .Y(new_n5679));
  nand_5 g03331(.A(n21654), .B(new_n3653), .Y(new_n5680_1));
  and_5  g03332(.A(new_n5680_1), .B(new_n5679), .Y(new_n5681));
  not_8  g03333(.A(new_n5681), .Y(new_n5682));
  nand_5 g03334(.A(new_n5682), .B(n17968), .Y(new_n5683));
  not_8  g03335(.A(n23146), .Y(new_n5684));
  not_8  g03336(.A(new_n5679), .Y(new_n5685));
  nand_5 g03337(.A(new_n3553), .B(n23842), .Y(new_n5686));
  not_8  g03338(.A(n23842), .Y(new_n5687_1));
  nand_5 g03339(.A(n25471), .B(new_n5687_1), .Y(new_n5688));
  and_5  g03340(.A(new_n5688), .B(new_n5686), .Y(new_n5689));
  xor_4  g03341(.A(new_n5689), .B(new_n5685), .Y(new_n5690));
  nand_5 g03342(.A(new_n5690), .B(new_n5684), .Y(new_n5691));
  or_5   g03343(.A(new_n5690), .B(new_n5684), .Y(new_n5692));
  nand_5 g03344(.A(new_n5692), .B(new_n5691), .Y(new_n5693));
  xnor_4 g03345(.A(new_n5693), .B(new_n5683), .Y(new_n5694));
  or_5   g03346(.A(new_n5694), .B(new_n5677), .Y(new_n5695));
  nand_5 g03347(.A(new_n5694), .B(new_n5677), .Y(new_n5696_1));
  xor_4  g03348(.A(new_n5671), .B(new_n5669), .Y(new_n5697));
  not_8  g03349(.A(new_n5697), .Y(new_n5698));
  not_8  g03350(.A(n17968), .Y(new_n5699));
  nand_5 g03351(.A(new_n5682), .B(new_n5699), .Y(new_n5700_1));
  nand_5 g03352(.A(new_n5681), .B(n17968), .Y(new_n5701));
  nand_5 g03353(.A(new_n5701), .B(new_n5700_1), .Y(new_n5702));
  nand_5 g03354(.A(new_n5702), .B(new_n5698), .Y(new_n5703));
  not_8  g03355(.A(new_n5703), .Y(new_n5704_1));
  nand_5 g03356(.A(new_n5704_1), .B(new_n5696_1), .Y(new_n5705));
  nand_5 g03357(.A(new_n5705), .B(new_n5695), .Y(new_n5706));
  nand_5 g03358(.A(new_n5674), .B(new_n5668), .Y(new_n5707));
  nand_5 g03359(.A(new_n5707), .B(new_n5673), .Y(new_n5708));
  not_8  g03360(.A(n8381), .Y(new_n5709));
  nand_5 g03361(.A(new_n5665), .B(new_n5663), .Y(new_n5710));
  nand_5 g03362(.A(new_n5710), .B(new_n5664), .Y(new_n5711));
  not_8  g03363(.A(new_n5711), .Y(new_n5712));
  nand_5 g03364(.A(new_n3046), .B(new_n2500), .Y(new_n5713));
  nand_5 g03365(.A(n18295), .B(n16223), .Y(new_n5714));
  nand_5 g03366(.A(new_n5714), .B(new_n5713), .Y(new_n5715));
  xor_4  g03367(.A(new_n5715), .B(new_n5712), .Y(new_n5716));
  not_8  g03368(.A(new_n5716), .Y(new_n5717));
  nand_5 g03369(.A(new_n5717), .B(new_n5709), .Y(new_n5718));
  nand_5 g03370(.A(new_n5716), .B(n8381), .Y(new_n5719));
  nand_5 g03371(.A(new_n5719), .B(new_n5718), .Y(new_n5720));
  xor_4  g03372(.A(new_n5720), .B(new_n5708), .Y(new_n5721));
  nand_5 g03373(.A(new_n5692), .B(new_n5683), .Y(new_n5722));
  nand_5 g03374(.A(new_n5722), .B(new_n5691), .Y(new_n5723));
  not_8  g03375(.A(n11184), .Y(new_n5724));
  nand_5 g03376(.A(new_n5688), .B(new_n5679), .Y(new_n5725));
  nand_5 g03377(.A(new_n5725), .B(new_n5686), .Y(new_n5726));
  not_8  g03378(.A(new_n5726), .Y(new_n5727));
  nand_5 g03379(.A(new_n3549), .B(n3828), .Y(new_n5728));
  not_8  g03380(.A(n3828), .Y(new_n5729));
  nand_5 g03381(.A(n15053), .B(new_n5729), .Y(new_n5730));
  nand_5 g03382(.A(new_n5730), .B(new_n5728), .Y(new_n5731));
  xor_4  g03383(.A(new_n5731), .B(new_n5727), .Y(new_n5732_1));
  not_8  g03384(.A(new_n5732_1), .Y(new_n5733));
  nand_5 g03385(.A(new_n5733), .B(new_n5724), .Y(new_n5734));
  nand_5 g03386(.A(new_n5732_1), .B(n11184), .Y(new_n5735));
  nand_5 g03387(.A(new_n5735), .B(new_n5734), .Y(new_n5736));
  xor_4  g03388(.A(new_n5736), .B(new_n5723), .Y(new_n5737));
  nand_5 g03389(.A(new_n5737), .B(new_n5721), .Y(new_n5738));
  or_5   g03390(.A(new_n5737), .B(new_n5721), .Y(new_n5739));
  nand_5 g03391(.A(new_n5739), .B(new_n5738), .Y(new_n5740));
  xnor_4 g03392(.A(new_n5740), .B(new_n5706), .Y(n357));
  nand_5 g03393(.A(n22309), .B(n9251), .Y(new_n5742_1));
  not_8  g03394(.A(n22309), .Y(new_n5743));
  nand_5 g03395(.A(new_n5743), .B(new_n3850_1), .Y(new_n5744));
  nand_5 g03396(.A(new_n5744), .B(new_n5742_1), .Y(new_n5745));
  nand_5 g03397(.A(new_n5232), .B(new_n2502), .Y(new_n5746));
  nand_5 g03398(.A(n25073), .B(n20138), .Y(new_n5747));
  nand_5 g03399(.A(new_n5747), .B(new_n5746), .Y(new_n5748));
  xnor_4 g03400(.A(new_n5748), .B(new_n5742_1), .Y(new_n5749));
  nand_5 g03401(.A(new_n5749), .B(new_n5745), .Y(new_n5750));
  nand_5 g03402(.A(new_n5747), .B(new_n5742_1), .Y(new_n5751));
  nand_5 g03403(.A(new_n5751), .B(new_n5746), .Y(new_n5752_1));
  not_8  g03404(.A(new_n5752_1), .Y(new_n5753));
  nand_5 g03405(.A(new_n5228_1), .B(new_n2498), .Y(new_n5754));
  nand_5 g03406(.A(n18171), .B(n6385), .Y(new_n5755));
  nand_5 g03407(.A(new_n5755), .B(new_n5754), .Y(new_n5756));
  xor_4  g03408(.A(new_n5756), .B(new_n5753), .Y(new_n5757));
  not_8  g03409(.A(new_n5757), .Y(new_n5758));
  nor_5  g03410(.A(new_n5758), .B(new_n5750), .Y(new_n5759));
  nand_5 g03411(.A(new_n5755), .B(new_n5752_1), .Y(new_n5760));
  nand_5 g03412(.A(new_n5760), .B(new_n5754), .Y(new_n5761));
  nand_5 g03413(.A(new_n5224), .B(new_n2494), .Y(new_n5762));
  nand_5 g03414(.A(n5752), .B(n3136), .Y(new_n5763));
  nand_5 g03415(.A(new_n5763), .B(new_n5762), .Y(new_n5764));
  xor_4  g03416(.A(new_n5764), .B(new_n5761), .Y(new_n5765_1));
  not_8  g03417(.A(new_n5765_1), .Y(new_n5766));
  nand_5 g03418(.A(new_n5766), .B(new_n5759), .Y(new_n5767));
  not_8  g03419(.A(new_n5759), .Y(new_n5768));
  nand_5 g03420(.A(new_n5765_1), .B(new_n5768), .Y(new_n5769));
  and_5  g03421(.A(new_n5769), .B(new_n5767), .Y(new_n5770));
  nand_5 g03422(.A(new_n5770), .B(new_n3399), .Y(new_n5771));
  or_5   g03423(.A(new_n5770), .B(new_n3399), .Y(new_n5772));
  nand_5 g03424(.A(new_n5758), .B(new_n5750), .Y(new_n5773));
  nand_5 g03425(.A(new_n5773), .B(new_n5768), .Y(new_n5774));
  or_5   g03426(.A(new_n5774), .B(new_n3407), .Y(new_n5775));
  nand_5 g03427(.A(new_n5774), .B(new_n3407), .Y(new_n5776_1));
  not_8  g03428(.A(new_n5745), .Y(new_n5777));
  nand_5 g03429(.A(new_n5777), .B(new_n3412), .Y(new_n5778));
  not_8  g03430(.A(new_n5778), .Y(new_n5779));
  nand_5 g03431(.A(new_n5779), .B(new_n3418), .Y(new_n5780));
  nand_5 g03432(.A(new_n5778), .B(new_n3419), .Y(new_n5781));
  xor_4  g03433(.A(new_n5749), .B(new_n5777), .Y(new_n5782_1));
  not_8  g03434(.A(new_n5782_1), .Y(new_n5783));
  nand_5 g03435(.A(new_n5783), .B(new_n5781), .Y(new_n5784));
  nand_5 g03436(.A(new_n5784), .B(new_n5780), .Y(new_n5785));
  nand_5 g03437(.A(new_n5785), .B(new_n5776_1), .Y(new_n5786));
  nand_5 g03438(.A(new_n5786), .B(new_n5775), .Y(new_n5787));
  nand_5 g03439(.A(new_n5787), .B(new_n5772), .Y(new_n5788));
  nand_5 g03440(.A(new_n5788), .B(new_n5771), .Y(new_n5789));
  not_8  g03441(.A(new_n5767), .Y(new_n5790));
  nand_5 g03442(.A(new_n5763), .B(new_n5761), .Y(new_n5791));
  nand_5 g03443(.A(new_n5791), .B(new_n5762), .Y(new_n5792));
  nand_5 g03444(.A(new_n5244), .B(new_n2490), .Y(new_n5793));
  nand_5 g03445(.A(n16158), .B(n9557), .Y(new_n5794));
  nand_5 g03446(.A(new_n5794), .B(new_n5793), .Y(new_n5795));
  xor_4  g03447(.A(new_n5795), .B(new_n5792), .Y(new_n5796));
  not_8  g03448(.A(new_n5796), .Y(new_n5797));
  nand_5 g03449(.A(new_n5797), .B(new_n5790), .Y(new_n5798));
  nand_5 g03450(.A(new_n5796), .B(new_n5767), .Y(new_n5799));
  and_5  g03451(.A(new_n5799), .B(new_n5798), .Y(new_n5800));
  nand_5 g03452(.A(new_n5800), .B(new_n3393), .Y(new_n5801));
  or_5   g03453(.A(new_n5800), .B(new_n3393), .Y(new_n5802));
  nand_5 g03454(.A(new_n5802), .B(new_n5801), .Y(new_n5803));
  xor_4  g03455(.A(new_n5803), .B(new_n5789), .Y(new_n5804));
  nand_5 g03456(.A(n18274), .B(new_n5150), .Y(new_n5805));
  not_8  g03457(.A(n18274), .Y(new_n5806));
  nand_5 g03458(.A(new_n5806), .B(n13263), .Y(new_n5807));
  nand_5 g03459(.A(new_n5136), .B(n3828), .Y(new_n5808));
  nand_5 g03460(.A(n20455), .B(new_n5729), .Y(new_n5809));
  nand_5 g03461(.A(n23842), .B(new_n5140_1), .Y(new_n5810));
  nand_5 g03462(.A(new_n5687_1), .B(n1639), .Y(new_n5811));
  nand_5 g03463(.A(new_n5678), .B(n16968), .Y(new_n5812));
  nand_5 g03464(.A(new_n5812), .B(new_n5811), .Y(new_n5813));
  nand_5 g03465(.A(new_n5813), .B(new_n5810), .Y(new_n5814));
  nand_5 g03466(.A(new_n5814), .B(new_n5809), .Y(new_n5815));
  nand_5 g03467(.A(new_n5815), .B(new_n5808), .Y(new_n5816));
  nand_5 g03468(.A(new_n5816), .B(new_n5807), .Y(new_n5817));
  nand_5 g03469(.A(new_n5817), .B(new_n5805), .Y(new_n5818));
  nand_5 g03470(.A(n21649), .B(new_n5204), .Y(new_n5819));
  not_8  g03471(.A(n21649), .Y(new_n5820));
  nand_5 g03472(.A(new_n5820), .B(n14510), .Y(new_n5821));
  nand_5 g03473(.A(new_n5821), .B(new_n5819), .Y(new_n5822_1));
  xor_4  g03474(.A(new_n5822_1), .B(new_n5818), .Y(new_n5823));
  nand_5 g03475(.A(new_n5823), .B(new_n5804), .Y(new_n5824));
  not_8  g03476(.A(new_n5824), .Y(new_n5825));
  nor_5  g03477(.A(new_n5823), .B(new_n5804), .Y(new_n5826));
  nand_5 g03478(.A(new_n5772), .B(new_n5771), .Y(new_n5827));
  xor_4  g03479(.A(new_n5827), .B(new_n5787), .Y(new_n5828));
  nand_5 g03480(.A(new_n5807), .B(new_n5805), .Y(new_n5829));
  xor_4  g03481(.A(new_n5829), .B(new_n5816), .Y(new_n5830));
  or_5   g03482(.A(new_n5830), .B(new_n5828), .Y(new_n5831));
  nand_5 g03483(.A(new_n5830), .B(new_n5828), .Y(new_n5832));
  nand_5 g03484(.A(new_n5776_1), .B(new_n5775), .Y(new_n5833_1));
  xor_4  g03485(.A(new_n5833_1), .B(new_n5785), .Y(new_n5834_1));
  nand_5 g03486(.A(new_n5809), .B(new_n5808), .Y(new_n5835));
  xor_4  g03487(.A(new_n5835), .B(new_n5814), .Y(new_n5836));
  or_5   g03488(.A(new_n5836), .B(new_n5834_1), .Y(new_n5837));
  nand_5 g03489(.A(new_n5836), .B(new_n5834_1), .Y(new_n5838));
  xor_4  g03490(.A(new_n5745), .B(new_n3412), .Y(new_n5839));
  xor_4  g03491(.A(n21654), .B(new_n3960), .Y(new_n5840_1));
  nor_5  g03492(.A(new_n5840_1), .B(new_n5839), .Y(new_n5841_1));
  nand_5 g03493(.A(new_n5811), .B(new_n5810), .Y(new_n5842_1));
  xnor_4 g03494(.A(new_n5842_1), .B(new_n5812), .Y(new_n5843));
  nand_5 g03495(.A(new_n5843), .B(new_n5841_1), .Y(new_n5844));
  not_8  g03496(.A(new_n5844), .Y(new_n5845));
  nand_5 g03497(.A(new_n5781), .B(new_n5780), .Y(new_n5846));
  xor_4  g03498(.A(new_n5846), .B(new_n5782_1), .Y(new_n5847));
  not_8  g03499(.A(new_n5847), .Y(new_n5848));
  nor_5  g03500(.A(new_n5843), .B(new_n5841_1), .Y(new_n5849));
  nor_5  g03501(.A(new_n5849), .B(new_n5848), .Y(new_n5850_1));
  nor_5  g03502(.A(new_n5850_1), .B(new_n5845), .Y(new_n5851));
  not_8  g03503(.A(new_n5851), .Y(new_n5852));
  nand_5 g03504(.A(new_n5852), .B(new_n5838), .Y(new_n5853));
  nand_5 g03505(.A(new_n5853), .B(new_n5837), .Y(new_n5854));
  nand_5 g03506(.A(new_n5854), .B(new_n5832), .Y(new_n5855));
  nand_5 g03507(.A(new_n5855), .B(new_n5831), .Y(new_n5856));
  nor_5  g03508(.A(new_n5856), .B(new_n5826), .Y(new_n5857));
  nor_5  g03509(.A(new_n5857), .B(new_n5825), .Y(new_n5858));
  nand_5 g03510(.A(new_n5802), .B(new_n5789), .Y(new_n5859));
  nand_5 g03511(.A(new_n5859), .B(new_n5801), .Y(new_n5860));
  nand_5 g03512(.A(new_n5794), .B(new_n5792), .Y(new_n5861));
  nand_5 g03513(.A(new_n5861), .B(new_n5793), .Y(new_n5862));
  nand_5 g03514(.A(new_n2516), .B(new_n5315), .Y(new_n5863));
  nand_5 g03515(.A(n25643), .B(n20604), .Y(new_n5864));
  nand_5 g03516(.A(new_n5864), .B(new_n5863), .Y(new_n5865));
  xor_4  g03517(.A(new_n5865), .B(new_n5862), .Y(new_n5866));
  or_5   g03518(.A(new_n5866), .B(new_n5798), .Y(new_n5867));
  nand_5 g03519(.A(new_n5866), .B(new_n5798), .Y(new_n5868));
  and_5  g03520(.A(new_n5868), .B(new_n5867), .Y(new_n5869));
  nand_5 g03521(.A(new_n5869), .B(new_n3387), .Y(new_n5870));
  or_5   g03522(.A(new_n5869), .B(new_n3387), .Y(new_n5871));
  nand_5 g03523(.A(new_n5871), .B(new_n5870), .Y(new_n5872));
  xor_4  g03524(.A(new_n5872), .B(new_n5860), .Y(new_n5873));
  not_8  g03525(.A(new_n5873), .Y(new_n5874));
  nand_5 g03526(.A(new_n5821), .B(new_n5818), .Y(new_n5875));
  nand_5 g03527(.A(new_n5875), .B(new_n5819), .Y(new_n5876));
  not_8  g03528(.A(new_n5876), .Y(new_n5877));
  nand_5 g03529(.A(n5255), .B(new_n5293), .Y(new_n5878));
  not_8  g03530(.A(n5255), .Y(new_n5879));
  nand_5 g03531(.A(new_n5879), .B(n4119), .Y(new_n5880));
  nand_5 g03532(.A(new_n5880), .B(new_n5878), .Y(new_n5881));
  xor_4  g03533(.A(new_n5881), .B(new_n5877), .Y(new_n5882_1));
  or_5   g03534(.A(new_n5882_1), .B(new_n5874), .Y(new_n5883));
  not_8  g03535(.A(new_n5883), .Y(new_n5884));
  nand_5 g03536(.A(new_n5882_1), .B(new_n5874), .Y(new_n5885));
  not_8  g03537(.A(new_n5885), .Y(new_n5886));
  nor_5  g03538(.A(new_n5886), .B(new_n5884), .Y(new_n5887));
  xor_4  g03539(.A(new_n5887), .B(new_n5858), .Y(n422));
  not_8  g03540(.A(n5302), .Y(new_n5889));
  nand_5 g03541(.A(new_n3654), .B(new_n3552), .Y(new_n5890));
  or_5   g03542(.A(new_n5890), .B(n14603), .Y(new_n5891));
  nor_5  g03543(.A(new_n5891), .B(n18737), .Y(new_n5892));
  nand_5 g03544(.A(new_n5892), .B(new_n3567), .Y(new_n5893));
  nor_5  g03545(.A(new_n5893), .B(n25738), .Y(new_n5894));
  nand_5 g03546(.A(new_n5894), .B(new_n5889), .Y(new_n5895));
  not_8  g03547(.A(new_n5895), .Y(new_n5896));
  nor_5  g03548(.A(new_n5894), .B(new_n5889), .Y(new_n5897));
  nor_5  g03549(.A(new_n5897), .B(new_n5896), .Y(new_n5898));
  or_5   g03550(.A(new_n5898), .B(n19770), .Y(new_n5899));
  nand_5 g03551(.A(new_n5898), .B(n19770), .Y(new_n5900));
  xor_4  g03552(.A(new_n5893), .B(n25738), .Y(new_n5901));
  or_5   g03553(.A(new_n5901), .B(n8782), .Y(new_n5902));
  nand_5 g03554(.A(new_n5901), .B(n8782), .Y(new_n5903_1));
  xor_4  g03555(.A(new_n5892), .B(new_n3567), .Y(new_n5904_1));
  or_5   g03556(.A(new_n5904_1), .B(n8678), .Y(new_n5905));
  nand_5 g03557(.A(new_n5904_1), .B(n8678), .Y(new_n5906));
  xor_4  g03558(.A(new_n5891), .B(n18737), .Y(new_n5907));
  or_5   g03559(.A(new_n5907), .B(n1432), .Y(new_n5908));
  nand_5 g03560(.A(new_n5907), .B(n1432), .Y(new_n5909));
  nand_5 g03561(.A(new_n5890), .B(n14603), .Y(new_n5910));
  nand_5 g03562(.A(new_n5910), .B(new_n5891), .Y(new_n5911_1));
  nand_5 g03563(.A(new_n5911_1), .B(new_n3403), .Y(new_n5912));
  nor_5  g03564(.A(new_n5911_1), .B(new_n3403), .Y(new_n5913));
  not_8  g03565(.A(new_n5913), .Y(new_n5914));
  nand_5 g03566(.A(n23333), .B(n20794), .Y(new_n5915));
  and_5  g03567(.A(new_n5915), .B(new_n5890), .Y(new_n5916));
  or_5   g03568(.A(new_n5916), .B(n25336), .Y(new_n5917));
  nand_5 g03569(.A(new_n5916), .B(n25336), .Y(new_n5918));
  nand_5 g03570(.A(n23333), .B(n11424), .Y(new_n5919));
  nand_5 g03571(.A(new_n5919), .B(new_n5918), .Y(new_n5920));
  nand_5 g03572(.A(new_n5920), .B(new_n5917), .Y(new_n5921));
  nand_5 g03573(.A(new_n5921), .B(new_n5914), .Y(new_n5922));
  nand_5 g03574(.A(new_n5922), .B(new_n5912), .Y(new_n5923));
  nand_5 g03575(.A(new_n5923), .B(new_n5909), .Y(new_n5924));
  nand_5 g03576(.A(new_n5924), .B(new_n5908), .Y(new_n5925));
  nand_5 g03577(.A(new_n5925), .B(new_n5906), .Y(new_n5926));
  nand_5 g03578(.A(new_n5926), .B(new_n5905), .Y(new_n5927));
  nand_5 g03579(.A(new_n5927), .B(new_n5903_1), .Y(new_n5928));
  nand_5 g03580(.A(new_n5928), .B(new_n5902), .Y(new_n5929));
  nand_5 g03581(.A(new_n5929), .B(new_n5900), .Y(new_n5930));
  nand_5 g03582(.A(new_n5930), .B(new_n5899), .Y(new_n5931));
  nand_5 g03583(.A(new_n5896), .B(new_n3545), .Y(new_n5932));
  nand_5 g03584(.A(new_n5895), .B(n3228), .Y(new_n5933));
  and_5  g03585(.A(new_n5933), .B(new_n5932), .Y(new_n5934));
  or_5   g03586(.A(new_n5934), .B(n26036), .Y(new_n5935));
  nand_5 g03587(.A(new_n5934), .B(n26036), .Y(new_n5936_1));
  nand_5 g03588(.A(new_n5936_1), .B(new_n5935), .Y(new_n5937));
  xor_4  g03589(.A(new_n5937), .B(new_n5931), .Y(new_n5938));
  nand_5 g03590(.A(new_n3034), .B(new_n3328), .Y(new_n5939));
  nand_5 g03591(.A(n7099), .B(n6691), .Y(new_n5940));
  nand_5 g03592(.A(new_n3039), .B(new_n3331), .Y(new_n5941));
  nand_5 g03593(.A(n12811), .B(n3260), .Y(new_n5942));
  nand_5 g03594(.A(new_n3334), .B(new_n3042), .Y(new_n5943_1));
  nand_5 g03595(.A(n20489), .B(n1118), .Y(new_n5944));
  nand_5 g03596(.A(new_n3047), .B(new_n3337), .Y(new_n5945));
  nand_5 g03597(.A(n25974), .B(n2355), .Y(new_n5946));
  nand_5 g03598(.A(new_n3340_1), .B(new_n3050), .Y(new_n5947));
  nand_5 g03599(.A(n11121), .B(n1630), .Y(new_n5948));
  nand_5 g03600(.A(n16217), .B(n1451), .Y(new_n5949));
  nand_5 g03601(.A(new_n5949), .B(new_n5948), .Y(new_n5950));
  nand_5 g03602(.A(new_n5950), .B(new_n5947), .Y(new_n5951));
  nand_5 g03603(.A(new_n5951), .B(new_n5946), .Y(new_n5952));
  nand_5 g03604(.A(new_n5952), .B(new_n5945), .Y(new_n5953));
  nand_5 g03605(.A(new_n5953), .B(new_n5944), .Y(new_n5954));
  nand_5 g03606(.A(new_n5954), .B(new_n5943_1), .Y(new_n5955));
  nand_5 g03607(.A(new_n5955), .B(new_n5942), .Y(new_n5956));
  nand_5 g03608(.A(new_n5956), .B(new_n5941), .Y(new_n5957));
  nand_5 g03609(.A(new_n5957), .B(new_n5940), .Y(new_n5958));
  nand_5 g03610(.A(new_n5958), .B(new_n5939), .Y(new_n5959));
  not_8  g03611(.A(new_n5959), .Y(new_n5960));
  nand_5 g03612(.A(n20700), .B(n932), .Y(new_n5961));
  nand_5 g03613(.A(new_n3067_1), .B(new_n3325), .Y(new_n5962));
  nand_5 g03614(.A(new_n5962), .B(new_n5961), .Y(new_n5963));
  xor_4  g03615(.A(new_n5963), .B(new_n5960), .Y(new_n5964_1));
  not_8  g03616(.A(new_n5964_1), .Y(new_n5965));
  nand_5 g03617(.A(new_n2468), .B(new_n3000), .Y(new_n5966));
  nand_5 g03618(.A(n26823), .B(n2035), .Y(new_n5967));
  nand_5 g03619(.A(n5213), .B(n4812), .Y(new_n5968));
  nand_5 g03620(.A(new_n2350), .B(new_n3007), .Y(new_n5969));
  nand_5 g03621(.A(n24278), .B(n4665), .Y(new_n5970));
  nand_5 g03622(.A(new_n2354), .B(new_n3010_1), .Y(new_n5971));
  nand_5 g03623(.A(n24618), .B(n19005), .Y(new_n5972));
  nand_5 g03624(.A(new_n3013), .B(new_n2357), .Y(new_n5973));
  nand_5 g03625(.A(n4326), .B(n3952), .Y(new_n5974));
  nand_5 g03626(.A(n12315), .B(n5438), .Y(new_n5975));
  nand_5 g03627(.A(new_n5975), .B(new_n5974), .Y(new_n5976));
  nand_5 g03628(.A(new_n5976), .B(new_n5973), .Y(new_n5977));
  nand_5 g03629(.A(new_n5977), .B(new_n5972), .Y(new_n5978));
  nand_5 g03630(.A(new_n5978), .B(new_n5971), .Y(new_n5979));
  nand_5 g03631(.A(new_n5979), .B(new_n5970), .Y(new_n5980_1));
  nand_5 g03632(.A(new_n5980_1), .B(new_n5969), .Y(new_n5981));
  nand_5 g03633(.A(new_n5981), .B(new_n5968), .Y(new_n5982));
  nand_5 g03634(.A(new_n3004), .B(new_n2371), .Y(new_n5983));
  nand_5 g03635(.A(new_n5983), .B(new_n5982), .Y(new_n5984));
  nand_5 g03636(.A(new_n5984), .B(new_n5967), .Y(new_n5985));
  nand_5 g03637(.A(new_n5985), .B(new_n5966), .Y(new_n5986));
  nand_5 g03638(.A(new_n2997), .B(new_n2584), .Y(new_n5987));
  nand_5 g03639(.A(n12875), .B(n7751), .Y(new_n5988));
  nand_5 g03640(.A(new_n5988), .B(new_n5987), .Y(new_n5989));
  xor_4  g03641(.A(new_n5989), .B(new_n5986), .Y(new_n5990));
  not_8  g03642(.A(new_n5990), .Y(new_n5991));
  nand_5 g03643(.A(new_n5991), .B(new_n5965), .Y(new_n5992));
  not_8  g03644(.A(new_n5992), .Y(new_n5993));
  nand_5 g03645(.A(new_n5990), .B(new_n5964_1), .Y(new_n5994));
  not_8  g03646(.A(new_n5994), .Y(new_n5995));
  nand_5 g03647(.A(new_n5967), .B(new_n5966), .Y(new_n5996));
  xor_4  g03648(.A(new_n5996), .B(new_n5984), .Y(new_n5997));
  not_8  g03649(.A(new_n5997), .Y(new_n5998));
  nand_5 g03650(.A(new_n5940), .B(new_n5939), .Y(new_n5999));
  xor_4  g03651(.A(new_n5999), .B(new_n5957), .Y(new_n6000));
  nand_5 g03652(.A(new_n6000), .B(new_n5998), .Y(new_n6001));
  not_8  g03653(.A(new_n6001), .Y(new_n6002));
  not_8  g03654(.A(new_n6000), .Y(new_n6003));
  nand_5 g03655(.A(new_n6003), .B(new_n5997), .Y(new_n6004));
  not_8  g03656(.A(new_n6004), .Y(new_n6005));
  nand_5 g03657(.A(new_n5942), .B(new_n5941), .Y(new_n6006));
  xor_4  g03658(.A(new_n6006), .B(new_n5955), .Y(new_n6007));
  nand_5 g03659(.A(new_n5944), .B(new_n5943_1), .Y(new_n6008));
  xor_4  g03660(.A(new_n6008), .B(new_n5953), .Y(new_n6009));
  nand_5 g03661(.A(new_n5970), .B(new_n5969), .Y(new_n6010));
  xor_4  g03662(.A(new_n6010), .B(new_n5979), .Y(new_n6011));
  not_8  g03663(.A(new_n6011), .Y(new_n6012_1));
  nand_5 g03664(.A(new_n6012_1), .B(new_n6009), .Y(new_n6013));
  or_5   g03665(.A(new_n6012_1), .B(new_n6009), .Y(new_n6014));
  nand_5 g03666(.A(new_n5946), .B(new_n5945), .Y(new_n6015));
  xor_4  g03667(.A(new_n6015), .B(new_n5951), .Y(new_n6016));
  nand_5 g03668(.A(new_n5972), .B(new_n5971), .Y(new_n6017));
  xor_4  g03669(.A(new_n6017), .B(new_n5977), .Y(new_n6018));
  not_8  g03670(.A(new_n6018), .Y(new_n6019));
  nand_5 g03671(.A(new_n6019), .B(new_n6016), .Y(new_n6020));
  or_5   g03672(.A(new_n6019), .B(new_n6016), .Y(new_n6021));
  nand_5 g03673(.A(new_n5974), .B(new_n5973), .Y(new_n6022_1));
  xor_4  g03674(.A(new_n6022_1), .B(new_n5975), .Y(new_n6023));
  not_8  g03675(.A(new_n6023), .Y(new_n6024));
  nand_5 g03676(.A(new_n5948), .B(new_n5947), .Y(new_n6025));
  xor_4  g03677(.A(new_n6025), .B(new_n5949), .Y(new_n6026));
  nand_5 g03678(.A(new_n6026), .B(new_n6024), .Y(new_n6027));
  or_5   g03679(.A(new_n6026), .B(new_n6024), .Y(new_n6028));
  nand_5 g03680(.A(new_n2443), .B(new_n3015), .Y(new_n6029));
  and_5  g03681(.A(new_n6029), .B(new_n5975), .Y(new_n6030));
  not_8  g03682(.A(new_n6030), .Y(new_n6031_1));
  nand_5 g03683(.A(new_n3410), .B(new_n3158), .Y(new_n6032));
  and_5  g03684(.A(new_n6032), .B(new_n5949), .Y(new_n6033));
  or_5   g03685(.A(new_n6033), .B(new_n6031_1), .Y(new_n6034));
  nand_5 g03686(.A(new_n6034), .B(new_n6028), .Y(new_n6035));
  nand_5 g03687(.A(new_n6035), .B(new_n6027), .Y(new_n6036));
  nand_5 g03688(.A(new_n6036), .B(new_n6021), .Y(new_n6037));
  nand_5 g03689(.A(new_n6037), .B(new_n6020), .Y(new_n6038));
  nand_5 g03690(.A(new_n6038), .B(new_n6014), .Y(new_n6039));
  nand_5 g03691(.A(new_n6039), .B(new_n6013), .Y(new_n6040));
  nand_5 g03692(.A(new_n6040), .B(new_n6007), .Y(new_n6041));
  not_8  g03693(.A(new_n6041), .Y(new_n6042));
  nor_5  g03694(.A(new_n6040), .B(new_n6007), .Y(new_n6043));
  nand_5 g03695(.A(new_n5983), .B(new_n5968), .Y(new_n6044_1));
  xor_4  g03696(.A(new_n6044_1), .B(new_n5981), .Y(new_n6045));
  nor_5  g03697(.A(new_n6045), .B(new_n6043), .Y(new_n6046_1));
  nor_5  g03698(.A(new_n6046_1), .B(new_n6042), .Y(new_n6047));
  nor_5  g03699(.A(new_n6047), .B(new_n6005), .Y(new_n6048));
  nor_5  g03700(.A(new_n6048), .B(new_n6002), .Y(new_n6049));
  nor_5  g03701(.A(new_n6049), .B(new_n5995), .Y(new_n6050));
  nor_5  g03702(.A(new_n6050), .B(new_n5993), .Y(new_n6051));
  not_8  g03703(.A(new_n6051), .Y(new_n6052));
  nand_5 g03704(.A(new_n5961), .B(new_n5959), .Y(new_n6053));
  nand_5 g03705(.A(new_n6053), .B(new_n5962), .Y(new_n6054));
  not_8  g03706(.A(new_n6054), .Y(new_n6055));
  nand_5 g03707(.A(n13367), .B(n7437), .Y(new_n6056));
  nand_5 g03708(.A(new_n3322), .B(new_n3185), .Y(new_n6057));
  nand_5 g03709(.A(new_n6057), .B(new_n6056), .Y(new_n6058));
  xor_4  g03710(.A(new_n6058), .B(new_n6055), .Y(new_n6059));
  nand_5 g03711(.A(new_n5988), .B(new_n5986), .Y(new_n6060));
  nand_5 g03712(.A(new_n6060), .B(new_n5987), .Y(new_n6061));
  not_8  g03713(.A(n20946), .Y(new_n6062));
  nand_5 g03714(.A(new_n6062), .B(new_n3030_1), .Y(new_n6063));
  nand_5 g03715(.A(n20946), .B(n1662), .Y(new_n6064));
  nand_5 g03716(.A(new_n6064), .B(new_n6063), .Y(new_n6065));
  xor_4  g03717(.A(new_n6065), .B(new_n6061), .Y(new_n6066));
  or_5   g03718(.A(new_n6066), .B(new_n6059), .Y(new_n6067));
  nand_5 g03719(.A(new_n6066), .B(new_n6059), .Y(new_n6068));
  nand_5 g03720(.A(new_n6068), .B(new_n6067), .Y(new_n6069));
  xor_4  g03721(.A(new_n6069), .B(new_n6052), .Y(new_n6070));
  not_8  g03722(.A(new_n6070), .Y(new_n6071));
  or_5   g03723(.A(new_n6071), .B(new_n5938), .Y(new_n6072));
  nand_5 g03724(.A(new_n6071), .B(new_n5938), .Y(new_n6073));
  nand_5 g03725(.A(new_n5900), .B(new_n5899), .Y(new_n6074));
  xor_4  g03726(.A(new_n6074), .B(new_n5929), .Y(new_n6075));
  nand_5 g03727(.A(new_n5994), .B(new_n5992), .Y(new_n6076));
  xor_4  g03728(.A(new_n6076), .B(new_n6049), .Y(new_n6077));
  or_5   g03729(.A(new_n6077), .B(new_n6075), .Y(new_n6078));
  nand_5 g03730(.A(new_n6077), .B(new_n6075), .Y(new_n6079));
  nand_5 g03731(.A(new_n5903_1), .B(new_n5902), .Y(new_n6080));
  xor_4  g03732(.A(new_n6080), .B(new_n5927), .Y(new_n6081));
  nand_5 g03733(.A(new_n6004), .B(new_n6001), .Y(new_n6082));
  xor_4  g03734(.A(new_n6082), .B(new_n6047), .Y(new_n6083));
  or_5   g03735(.A(new_n6083), .B(new_n6081), .Y(new_n6084_1));
  nand_5 g03736(.A(new_n6083), .B(new_n6081), .Y(new_n6085));
  nand_5 g03737(.A(new_n5906), .B(new_n5905), .Y(new_n6086));
  xor_4  g03738(.A(new_n6086), .B(new_n5925), .Y(new_n6087));
  not_8  g03739(.A(new_n6045), .Y(new_n6088));
  nor_5  g03740(.A(new_n6043), .B(new_n6042), .Y(new_n6089));
  xor_4  g03741(.A(new_n6089), .B(new_n6088), .Y(new_n6090));
  or_5   g03742(.A(new_n6090), .B(new_n6087), .Y(new_n6091));
  nand_5 g03743(.A(new_n6090), .B(new_n6087), .Y(new_n6092));
  nand_5 g03744(.A(new_n5909), .B(new_n5908), .Y(new_n6093));
  xor_4  g03745(.A(new_n6093), .B(new_n5923), .Y(new_n6094));
  nand_5 g03746(.A(new_n6014), .B(new_n6013), .Y(new_n6095));
  xor_4  g03747(.A(new_n6095), .B(new_n6038), .Y(new_n6096));
  not_8  g03748(.A(new_n6096), .Y(new_n6097));
  or_5   g03749(.A(new_n6097), .B(new_n6094), .Y(new_n6098));
  nand_5 g03750(.A(new_n6097), .B(new_n6094), .Y(new_n6099));
  nand_5 g03751(.A(new_n6021), .B(new_n6020), .Y(new_n6100));
  xor_4  g03752(.A(new_n6100), .B(new_n6036), .Y(new_n6101));
  not_8  g03753(.A(new_n6101), .Y(new_n6102));
  nand_5 g03754(.A(new_n5914), .B(new_n5912), .Y(new_n6103));
  xor_4  g03755(.A(new_n6103), .B(new_n5921), .Y(new_n6104_1));
  or_5   g03756(.A(new_n6104_1), .B(new_n6102), .Y(new_n6105_1));
  nand_5 g03757(.A(new_n6104_1), .B(new_n6102), .Y(new_n6106));
  nand_5 g03758(.A(new_n5918), .B(new_n5917), .Y(new_n6107));
  xnor_4 g03759(.A(new_n6107), .B(new_n5919), .Y(new_n6108));
  nand_5 g03760(.A(new_n6028), .B(new_n6027), .Y(new_n6109));
  xor_4  g03761(.A(new_n6109), .B(new_n6034), .Y(new_n6110));
  nand_5 g03762(.A(new_n6110), .B(new_n6108), .Y(new_n6111));
  nor_5  g03763(.A(new_n6110), .B(new_n6108), .Y(new_n6112));
  not_8  g03764(.A(new_n6112), .Y(new_n6113));
  xor_4  g03765(.A(new_n6033), .B(new_n6031_1), .Y(new_n6114));
  nand_5 g03766(.A(new_n3654), .B(new_n3409), .Y(new_n6115));
  nand_5 g03767(.A(new_n6115), .B(new_n5919), .Y(new_n6116));
  nor_5  g03768(.A(new_n6116), .B(new_n6114), .Y(new_n6117));
  not_8  g03769(.A(new_n6117), .Y(new_n6118));
  nand_5 g03770(.A(new_n6118), .B(new_n6113), .Y(new_n6119));
  nand_5 g03771(.A(new_n6119), .B(new_n6111), .Y(new_n6120));
  nand_5 g03772(.A(new_n6120), .B(new_n6106), .Y(new_n6121));
  nand_5 g03773(.A(new_n6121), .B(new_n6105_1), .Y(new_n6122));
  nand_5 g03774(.A(new_n6122), .B(new_n6099), .Y(new_n6123));
  nand_5 g03775(.A(new_n6123), .B(new_n6098), .Y(new_n6124));
  nand_5 g03776(.A(new_n6124), .B(new_n6092), .Y(new_n6125));
  nand_5 g03777(.A(new_n6125), .B(new_n6091), .Y(new_n6126));
  nand_5 g03778(.A(new_n6126), .B(new_n6085), .Y(new_n6127));
  nand_5 g03779(.A(new_n6127), .B(new_n6084_1), .Y(new_n6128));
  nand_5 g03780(.A(new_n6128), .B(new_n6079), .Y(new_n6129));
  nand_5 g03781(.A(new_n6129), .B(new_n6078), .Y(new_n6130));
  nand_5 g03782(.A(new_n6130), .B(new_n6073), .Y(new_n6131));
  nand_5 g03783(.A(new_n6131), .B(new_n6072), .Y(new_n6132));
  nand_5 g03784(.A(new_n6068), .B(new_n6052), .Y(new_n6133));
  nand_5 g03785(.A(new_n6133), .B(new_n6067), .Y(new_n6134));
  nand_5 g03786(.A(new_n6064), .B(new_n6061), .Y(new_n6135));
  nand_5 g03787(.A(new_n6135), .B(new_n6063), .Y(new_n6136));
  not_8  g03788(.A(new_n6136), .Y(new_n6137));
  nand_5 g03789(.A(new_n3276), .B(new_n3442), .Y(new_n6138));
  nand_5 g03790(.A(n22379), .B(n9967), .Y(new_n6139));
  nand_5 g03791(.A(new_n6139), .B(new_n6138), .Y(new_n6140));
  xor_4  g03792(.A(new_n6140), .B(new_n6137), .Y(new_n6141));
  not_8  g03793(.A(new_n6141), .Y(new_n6142));
  nand_5 g03794(.A(new_n6056), .B(new_n6054), .Y(new_n6143));
  nand_5 g03795(.A(new_n6143), .B(new_n6057), .Y(new_n6144));
  not_8  g03796(.A(new_n6144), .Y(new_n6145));
  nand_5 g03797(.A(new_n3287), .B(new_n3317), .Y(new_n6146));
  nand_5 g03798(.A(n10763), .B(n5696), .Y(new_n6147));
  nand_5 g03799(.A(new_n6147), .B(new_n6146), .Y(new_n6148));
  xor_4  g03800(.A(new_n6148), .B(new_n6145), .Y(new_n6149));
  or_5   g03801(.A(new_n6149), .B(new_n6142), .Y(new_n6150));
  nand_5 g03802(.A(new_n6149), .B(new_n6142), .Y(new_n6151));
  nand_5 g03803(.A(new_n6151), .B(new_n6150), .Y(new_n6152));
  xor_4  g03804(.A(new_n6152), .B(new_n6134), .Y(new_n6153));
  not_8  g03805(.A(new_n6153), .Y(new_n6154));
  nand_5 g03806(.A(new_n5936_1), .B(new_n5931), .Y(new_n6155));
  nand_5 g03807(.A(new_n6155), .B(new_n5935), .Y(new_n6156));
  or_5   g03808(.A(new_n5932), .B(n337), .Y(new_n6157));
  nand_5 g03809(.A(new_n5932), .B(n337), .Y(new_n6158));
  and_5  g03810(.A(new_n6158), .B(new_n6157), .Y(new_n6159));
  or_5   g03811(.A(new_n6159), .B(n6485), .Y(new_n6160_1));
  nand_5 g03812(.A(new_n6159), .B(n6485), .Y(new_n6161));
  nand_5 g03813(.A(new_n6161), .B(new_n6160_1), .Y(new_n6162));
  xor_4  g03814(.A(new_n6162), .B(new_n6156), .Y(new_n6163));
  nand_5 g03815(.A(new_n6163), .B(new_n6154), .Y(new_n6164));
  or_5   g03816(.A(new_n6163), .B(new_n6154), .Y(new_n6165));
  nand_5 g03817(.A(new_n6165), .B(new_n6164), .Y(new_n6166));
  xor_4  g03818(.A(new_n6166), .B(new_n6132), .Y(n431));
  not_8  g03819(.A(n26797), .Y(new_n6168));
  not_8  g03820(.A(n22554), .Y(new_n6169));
  not_8  g03821(.A(n3909), .Y(new_n6170));
  not_8  g03822(.A(n22173), .Y(new_n6171_1));
  nand_5 g03823(.A(new_n6171_1), .B(new_n2620), .Y(new_n6172));
  or_5   g03824(.A(new_n6172), .B(n2146), .Y(new_n6173));
  nor_5  g03825(.A(new_n6173), .B(n23974), .Y(new_n6174));
  nand_5 g03826(.A(new_n6174), .B(new_n6170), .Y(new_n6175));
  nor_5  g03827(.A(new_n6175), .B(n20429), .Y(new_n6176));
  nand_5 g03828(.A(new_n6176), .B(new_n6169), .Y(new_n6177));
  nor_5  g03829(.A(new_n6177), .B(n23913), .Y(new_n6178));
  nand_5 g03830(.A(new_n6178), .B(new_n6168), .Y(new_n6179));
  nor_5  g03831(.A(new_n6179), .B(n12702), .Y(new_n6180));
  not_8  g03832(.A(new_n6180), .Y(new_n6181));
  nand_5 g03833(.A(new_n6179), .B(n12702), .Y(new_n6182));
  and_5  g03834(.A(new_n6182), .B(new_n6181), .Y(new_n6183_1));
  or_5   g03835(.A(new_n6183_1), .B(n12650), .Y(new_n6184));
  nand_5 g03836(.A(new_n6183_1), .B(n12650), .Y(new_n6185));
  nand_5 g03837(.A(new_n6185), .B(new_n6184), .Y(new_n6186));
  xor_4  g03838(.A(new_n6178), .B(new_n6168), .Y(new_n6187));
  or_5   g03839(.A(new_n6187), .B(n10201), .Y(new_n6188));
  nand_5 g03840(.A(new_n6187), .B(n10201), .Y(new_n6189_1));
  xor_4  g03841(.A(new_n6177), .B(n23913), .Y(new_n6190));
  or_5   g03842(.A(new_n6190), .B(n10593), .Y(new_n6191));
  nand_5 g03843(.A(new_n6190), .B(n10593), .Y(new_n6192));
  xor_4  g03844(.A(new_n6176), .B(new_n6169), .Y(new_n6193));
  or_5   g03845(.A(new_n6193), .B(n18290), .Y(new_n6194));
  nand_5 g03846(.A(new_n6193), .B(n18290), .Y(new_n6195));
  xor_4  g03847(.A(new_n6175), .B(n20429), .Y(new_n6196));
  or_5   g03848(.A(new_n6196), .B(n11580), .Y(new_n6197));
  nand_5 g03849(.A(new_n6196), .B(n11580), .Y(new_n6198));
  xor_4  g03850(.A(new_n6174), .B(new_n6170), .Y(new_n6199));
  or_5   g03851(.A(new_n6199), .B(n15884), .Y(new_n6200));
  nand_5 g03852(.A(new_n6199), .B(n15884), .Y(new_n6201));
  xor_4  g03853(.A(new_n6173), .B(n23974), .Y(new_n6202));
  or_5   g03854(.A(new_n6202), .B(n6356), .Y(new_n6203));
  nand_5 g03855(.A(new_n6202), .B(n6356), .Y(new_n6204_1));
  not_8  g03856(.A(n27104), .Y(new_n6205));
  nand_5 g03857(.A(new_n6172), .B(n2146), .Y(new_n6206));
  nand_5 g03858(.A(new_n6206), .B(new_n6173), .Y(new_n6207));
  nand_5 g03859(.A(new_n6207), .B(new_n6205), .Y(new_n6208));
  nor_5  g03860(.A(new_n6207), .B(new_n6205), .Y(new_n6209));
  not_8  g03861(.A(new_n6209), .Y(new_n6210));
  nand_5 g03862(.A(n22173), .B(n583), .Y(new_n6211));
  and_5  g03863(.A(new_n6211), .B(new_n6172), .Y(new_n6212));
  or_5   g03864(.A(new_n6212), .B(n27188), .Y(new_n6213));
  nand_5 g03865(.A(new_n6212), .B(n27188), .Y(new_n6214));
  nand_5 g03866(.A(n6611), .B(n583), .Y(new_n6215));
  nand_5 g03867(.A(new_n6215), .B(new_n6214), .Y(new_n6216));
  nand_5 g03868(.A(new_n6216), .B(new_n6213), .Y(new_n6217));
  nand_5 g03869(.A(new_n6217), .B(new_n6210), .Y(new_n6218_1));
  nand_5 g03870(.A(new_n6218_1), .B(new_n6208), .Y(new_n6219));
  nand_5 g03871(.A(new_n6219), .B(new_n6204_1), .Y(new_n6220));
  nand_5 g03872(.A(new_n6220), .B(new_n6203), .Y(new_n6221));
  nand_5 g03873(.A(new_n6221), .B(new_n6201), .Y(new_n6222));
  nand_5 g03874(.A(new_n6222), .B(new_n6200), .Y(new_n6223_1));
  nand_5 g03875(.A(new_n6223_1), .B(new_n6198), .Y(new_n6224));
  nand_5 g03876(.A(new_n6224), .B(new_n6197), .Y(new_n6225));
  nand_5 g03877(.A(new_n6225), .B(new_n6195), .Y(new_n6226));
  nand_5 g03878(.A(new_n6226), .B(new_n6194), .Y(new_n6227));
  nand_5 g03879(.A(new_n6227), .B(new_n6192), .Y(new_n6228));
  nand_5 g03880(.A(new_n6228), .B(new_n6191), .Y(new_n6229));
  nand_5 g03881(.A(new_n6229), .B(new_n6189_1), .Y(new_n6230));
  nand_5 g03882(.A(new_n6230), .B(new_n6188), .Y(new_n6231));
  xnor_4 g03883(.A(new_n6231), .B(new_n6186), .Y(new_n6232));
  not_8  g03884(.A(n13494), .Y(new_n6233_1));
  nand_5 g03885(.A(n18880), .B(new_n6233_1), .Y(new_n6234));
  nand_5 g03886(.A(new_n4966_1), .B(n13494), .Y(new_n6235));
  nand_5 g03887(.A(new_n6235), .B(new_n6234), .Y(new_n6236));
  nand_5 g03888(.A(new_n4942), .B(n25345), .Y(new_n6237));
  not_8  g03889(.A(n25345), .Y(new_n6238));
  nand_5 g03890(.A(n25475), .B(new_n6238), .Y(new_n6239));
  not_8  g03891(.A(n23849), .Y(new_n6240));
  nand_5 g03892(.A(new_n6240), .B(n9655), .Y(new_n6241));
  not_8  g03893(.A(n9655), .Y(new_n6242));
  nand_5 g03894(.A(n23849), .B(new_n6242), .Y(new_n6243));
  nand_5 g03895(.A(n13490), .B(new_n4952_1), .Y(new_n6244));
  nand_5 g03896(.A(new_n2585), .B(n12446), .Y(new_n6245_1));
  not_8  g03897(.A(n11011), .Y(new_n6246));
  nand_5 g03898(.A(n22660), .B(new_n6246), .Y(new_n6247));
  nand_5 g03899(.A(new_n2467), .B(n11011), .Y(new_n6248_1));
  not_8  g03900(.A(n16029), .Y(new_n6249));
  nand_5 g03901(.A(new_n6249), .B(n1777), .Y(new_n6250));
  nand_5 g03902(.A(n16029), .B(new_n2370), .Y(new_n6251));
  not_8  g03903(.A(n16476), .Y(new_n6252));
  nand_5 g03904(.A(new_n6252), .B(n8745), .Y(new_n6253));
  nand_5 g03905(.A(n16476), .B(new_n2349), .Y(new_n6254));
  not_8  g03906(.A(n11615), .Y(new_n6255));
  nand_5 g03907(.A(n15636), .B(new_n6255), .Y(new_n6256_1));
  nand_5 g03908(.A(new_n2353), .B(n11615), .Y(new_n6257));
  not_8  g03909(.A(n22433), .Y(new_n6258));
  nand_5 g03910(.A(new_n6258), .B(n20077), .Y(new_n6259));
  nand_5 g03911(.A(n22433), .B(new_n2358), .Y(new_n6260));
  nand_5 g03912(.A(n14090), .B(new_n2442), .Y(new_n6261));
  nand_5 g03913(.A(new_n6261), .B(new_n6260), .Y(new_n6262));
  nand_5 g03914(.A(new_n6262), .B(new_n6259), .Y(new_n6263));
  nand_5 g03915(.A(new_n6263), .B(new_n6257), .Y(new_n6264));
  nand_5 g03916(.A(new_n6264), .B(new_n6256_1), .Y(new_n6265));
  nand_5 g03917(.A(new_n6265), .B(new_n6254), .Y(new_n6266));
  nand_5 g03918(.A(new_n6266), .B(new_n6253), .Y(new_n6267));
  nand_5 g03919(.A(new_n6267), .B(new_n6251), .Y(new_n6268));
  nand_5 g03920(.A(new_n6268), .B(new_n6250), .Y(new_n6269));
  nand_5 g03921(.A(new_n6269), .B(new_n6248_1), .Y(new_n6270));
  nand_5 g03922(.A(new_n6270), .B(new_n6247), .Y(new_n6271_1));
  nand_5 g03923(.A(new_n6271_1), .B(new_n6245_1), .Y(new_n6272));
  nand_5 g03924(.A(new_n6272), .B(new_n6244), .Y(new_n6273));
  nand_5 g03925(.A(new_n6273), .B(new_n6243), .Y(new_n6274));
  nand_5 g03926(.A(new_n6274), .B(new_n6241), .Y(new_n6275));
  nand_5 g03927(.A(new_n6275), .B(new_n6239), .Y(new_n6276_1));
  nand_5 g03928(.A(new_n6276_1), .B(new_n6237), .Y(new_n6277));
  not_8  g03929(.A(new_n6277), .Y(new_n6278));
  xor_4  g03930(.A(new_n6278), .B(new_n6236), .Y(new_n6279));
  not_8  g03931(.A(new_n6279), .Y(new_n6280));
  or_5   g03932(.A(new_n6280), .B(new_n6232), .Y(new_n6281));
  nand_5 g03933(.A(new_n6280), .B(new_n6232), .Y(new_n6282));
  nand_5 g03934(.A(new_n6239), .B(new_n6237), .Y(new_n6283));
  xor_4  g03935(.A(new_n6283), .B(new_n6275), .Y(new_n6284));
  not_8  g03936(.A(new_n6284), .Y(new_n6285));
  nand_5 g03937(.A(new_n6189_1), .B(new_n6188), .Y(new_n6286));
  xor_4  g03938(.A(new_n6286), .B(new_n6229), .Y(new_n6287));
  nand_5 g03939(.A(new_n6287), .B(new_n6285), .Y(new_n6288));
  or_5   g03940(.A(new_n6287), .B(new_n6285), .Y(new_n6289));
  nand_5 g03941(.A(new_n6243), .B(new_n6241), .Y(new_n6290));
  xor_4  g03942(.A(new_n6290), .B(new_n6273), .Y(new_n6291));
  not_8  g03943(.A(new_n6291), .Y(new_n6292));
  nand_5 g03944(.A(new_n6192), .B(new_n6191), .Y(new_n6293));
  xor_4  g03945(.A(new_n6293), .B(new_n6227), .Y(new_n6294));
  nand_5 g03946(.A(new_n6294), .B(new_n6292), .Y(new_n6295));
  nor_5  g03947(.A(new_n6294), .B(new_n6292), .Y(new_n6296));
  not_8  g03948(.A(new_n6296), .Y(new_n6297));
  nand_5 g03949(.A(new_n6245_1), .B(new_n6244), .Y(new_n6298));
  xor_4  g03950(.A(new_n6298), .B(new_n6271_1), .Y(new_n6299));
  not_8  g03951(.A(new_n6299), .Y(new_n6300));
  nand_5 g03952(.A(new_n6195), .B(new_n6194), .Y(new_n6301));
  xor_4  g03953(.A(new_n6301), .B(new_n6225), .Y(new_n6302));
  nand_5 g03954(.A(new_n6302), .B(new_n6300), .Y(new_n6303));
  nor_5  g03955(.A(new_n6302), .B(new_n6300), .Y(new_n6304));
  not_8  g03956(.A(new_n6304), .Y(new_n6305));
  nand_5 g03957(.A(new_n6248_1), .B(new_n6247), .Y(new_n6306));
  xor_4  g03958(.A(new_n6306), .B(new_n6269), .Y(new_n6307));
  not_8  g03959(.A(new_n6307), .Y(new_n6308_1));
  nand_5 g03960(.A(new_n6198), .B(new_n6197), .Y(new_n6309));
  xor_4  g03961(.A(new_n6309), .B(new_n6223_1), .Y(new_n6310));
  nand_5 g03962(.A(new_n6310), .B(new_n6308_1), .Y(new_n6311_1));
  nor_5  g03963(.A(new_n6310), .B(new_n6308_1), .Y(new_n6312));
  not_8  g03964(.A(new_n6312), .Y(new_n6313));
  nand_5 g03965(.A(new_n6251), .B(new_n6250), .Y(new_n6314));
  xor_4  g03966(.A(new_n6314), .B(new_n6267), .Y(new_n6315));
  not_8  g03967(.A(new_n6315), .Y(new_n6316));
  nand_5 g03968(.A(new_n6201), .B(new_n6200), .Y(new_n6317));
  xor_4  g03969(.A(new_n6317), .B(new_n6221), .Y(new_n6318));
  nand_5 g03970(.A(new_n6318), .B(new_n6316), .Y(new_n6319));
  nor_5  g03971(.A(new_n6318), .B(new_n6316), .Y(new_n6320));
  not_8  g03972(.A(new_n6320), .Y(new_n6321));
  nand_5 g03973(.A(new_n6254), .B(new_n6253), .Y(new_n6322));
  xor_4  g03974(.A(new_n6322), .B(new_n6265), .Y(new_n6323_1));
  not_8  g03975(.A(new_n6323_1), .Y(new_n6324));
  nand_5 g03976(.A(new_n6204_1), .B(new_n6203), .Y(new_n6325));
  xor_4  g03977(.A(new_n6325), .B(new_n6219), .Y(new_n6326));
  nand_5 g03978(.A(new_n6326), .B(new_n6324), .Y(new_n6327));
  or_5   g03979(.A(new_n6326), .B(new_n6324), .Y(new_n6328));
  nand_5 g03980(.A(new_n6257), .B(new_n6256_1), .Y(new_n6329));
  xor_4  g03981(.A(new_n6329), .B(new_n6263), .Y(new_n6330_1));
  not_8  g03982(.A(new_n6330_1), .Y(new_n6331));
  nand_5 g03983(.A(new_n6210), .B(new_n6208), .Y(new_n6332));
  xor_4  g03984(.A(new_n6332), .B(new_n6217), .Y(new_n6333));
  nand_5 g03985(.A(new_n6333), .B(new_n6331), .Y(new_n6334));
  or_5   g03986(.A(new_n6333), .B(new_n6331), .Y(new_n6335));
  nand_5 g03987(.A(new_n2631), .B(n6794), .Y(new_n6336));
  and_5  g03988(.A(new_n6336), .B(new_n6261), .Y(new_n6337));
  not_8  g03989(.A(new_n6337), .Y(new_n6338));
  not_8  g03990(.A(n6611), .Y(new_n6339_1));
  nand_5 g03991(.A(new_n6339_1), .B(new_n2620), .Y(new_n6340));
  and_5  g03992(.A(new_n6340), .B(new_n6215), .Y(new_n6341));
  nand_5 g03993(.A(new_n6341), .B(new_n6338), .Y(new_n6342));
  and_5  g03994(.A(new_n6260), .B(new_n6259), .Y(new_n6343));
  xor_4  g03995(.A(new_n6343), .B(new_n6261), .Y(new_n6344));
  not_8  g03996(.A(new_n6344), .Y(new_n6345));
  or_5   g03997(.A(new_n6345), .B(new_n6342), .Y(new_n6346));
  nand_5 g03998(.A(new_n6345), .B(new_n6342), .Y(new_n6347));
  nand_5 g03999(.A(new_n6214), .B(new_n6213), .Y(new_n6348));
  xnor_4 g04000(.A(new_n6348), .B(new_n6215), .Y(new_n6349));
  not_8  g04001(.A(new_n6349), .Y(new_n6350));
  nand_5 g04002(.A(new_n6350), .B(new_n6347), .Y(new_n6351));
  nand_5 g04003(.A(new_n6351), .B(new_n6346), .Y(new_n6352));
  nand_5 g04004(.A(new_n6352), .B(new_n6335), .Y(new_n6353));
  nand_5 g04005(.A(new_n6353), .B(new_n6334), .Y(new_n6354_1));
  nand_5 g04006(.A(new_n6354_1), .B(new_n6328), .Y(new_n6355));
  nand_5 g04007(.A(new_n6355), .B(new_n6327), .Y(new_n6356_1));
  nand_5 g04008(.A(new_n6356_1), .B(new_n6321), .Y(new_n6357));
  nand_5 g04009(.A(new_n6357), .B(new_n6319), .Y(new_n6358));
  nand_5 g04010(.A(new_n6358), .B(new_n6313), .Y(new_n6359));
  nand_5 g04011(.A(new_n6359), .B(new_n6311_1), .Y(new_n6360));
  nand_5 g04012(.A(new_n6360), .B(new_n6305), .Y(new_n6361));
  nand_5 g04013(.A(new_n6361), .B(new_n6303), .Y(new_n6362));
  nand_5 g04014(.A(new_n6362), .B(new_n6297), .Y(new_n6363));
  nand_5 g04015(.A(new_n6363), .B(new_n6295), .Y(new_n6364));
  nand_5 g04016(.A(new_n6364), .B(new_n6289), .Y(new_n6365));
  nand_5 g04017(.A(new_n6365), .B(new_n6288), .Y(new_n6366));
  nand_5 g04018(.A(new_n6366), .B(new_n6282), .Y(new_n6367));
  nand_5 g04019(.A(new_n6367), .B(new_n6281), .Y(new_n6368));
  not_8  g04020(.A(new_n6184), .Y(new_n6369_1));
  nor_5  g04021(.A(new_n6231), .B(new_n6369_1), .Y(new_n6370));
  nand_5 g04022(.A(new_n6185), .B(new_n6181), .Y(new_n6371));
  nor_5  g04023(.A(new_n6371), .B(new_n6370), .Y(new_n6372));
  not_8  g04024(.A(new_n6372), .Y(new_n6373));
  nand_5 g04025(.A(new_n6373), .B(new_n6368), .Y(new_n6374));
  nor_5  g04026(.A(new_n6373), .B(new_n6368), .Y(new_n6375_1));
  not_8  g04027(.A(new_n6375_1), .Y(new_n6376));
  nand_5 g04028(.A(new_n6376), .B(new_n6374), .Y(new_n6377));
  nand_5 g04029(.A(new_n6277), .B(new_n6234), .Y(new_n6378));
  nand_5 g04030(.A(new_n6378), .B(new_n6235), .Y(new_n6379_1));
  xor_4  g04031(.A(new_n6379_1), .B(new_n6377), .Y(new_n6380));
  not_8  g04032(.A(new_n6380), .Y(new_n6381_1));
  not_8  g04033(.A(n8614), .Y(new_n6382));
  nand_5 g04034(.A(n23895), .B(new_n6382), .Y(new_n6383_1));
  not_8  g04035(.A(n23895), .Y(new_n6384));
  nand_5 g04036(.A(new_n6384), .B(n8614), .Y(new_n6385_1));
  not_8  g04037(.A(n15182), .Y(new_n6386));
  nand_5 g04038(.A(n17351), .B(new_n6386), .Y(new_n6387));
  not_8  g04039(.A(n17351), .Y(new_n6388));
  nand_5 g04040(.A(new_n6388), .B(n15182), .Y(new_n6389));
  not_8  g04041(.A(n27037), .Y(new_n6390));
  nand_5 g04042(.A(new_n6390), .B(n11736), .Y(new_n6391));
  not_8  g04043(.A(n11736), .Y(new_n6392));
  nand_5 g04044(.A(n27037), .B(new_n6392), .Y(new_n6393));
  not_8  g04045(.A(n8964), .Y(new_n6394));
  nand_5 g04046(.A(n23200), .B(new_n6394), .Y(new_n6395));
  not_8  g04047(.A(n23200), .Y(new_n6396));
  nand_5 g04048(.A(new_n6396), .B(n8964), .Y(new_n6397_1));
  nand_5 g04049(.A(new_n4512), .B(n17959), .Y(new_n6398));
  not_8  g04050(.A(n17959), .Y(new_n6399));
  nand_5 g04051(.A(n20151), .B(new_n6399), .Y(new_n6400));
  nand_5 g04052(.A(new_n4438), .B(n7566), .Y(new_n6401));
  not_8  g04053(.A(n7566), .Y(new_n6402));
  nand_5 g04054(.A(n7693), .B(new_n6402), .Y(new_n6403));
  nand_5 g04055(.A(new_n4396), .B(n7731), .Y(new_n6404));
  not_8  g04056(.A(n7731), .Y(new_n6405));
  nand_5 g04057(.A(n10405), .B(new_n6405), .Y(new_n6406));
  nand_5 g04058(.A(n12341), .B(new_n4376_1), .Y(new_n6407_1));
  not_8  g04059(.A(n12341), .Y(new_n6408));
  nand_5 g04060(.A(new_n6408), .B(n11302), .Y(new_n6409));
  nand_5 g04061(.A(n20986), .B(new_n4386), .Y(new_n6410));
  not_8  g04062(.A(n20986), .Y(new_n6411));
  nand_5 g04063(.A(new_n6411), .B(n17090), .Y(new_n6412));
  not_8  g04064(.A(n12384), .Y(new_n6413));
  nand_5 g04065(.A(new_n6413), .B(n6773), .Y(new_n6414));
  nand_5 g04066(.A(new_n6414), .B(new_n6412), .Y(new_n6415));
  nand_5 g04067(.A(new_n6415), .B(new_n6410), .Y(new_n6416));
  nand_5 g04068(.A(new_n6416), .B(new_n6409), .Y(new_n6417));
  nand_5 g04069(.A(new_n6417), .B(new_n6407_1), .Y(new_n6418));
  nand_5 g04070(.A(new_n6418), .B(new_n6406), .Y(new_n6419));
  nand_5 g04071(.A(new_n6419), .B(new_n6404), .Y(new_n6420));
  nand_5 g04072(.A(new_n6420), .B(new_n6403), .Y(new_n6421));
  nand_5 g04073(.A(new_n6421), .B(new_n6401), .Y(new_n6422));
  nand_5 g04074(.A(new_n6422), .B(new_n6400), .Y(new_n6423));
  nand_5 g04075(.A(new_n6423), .B(new_n6398), .Y(new_n6424));
  nand_5 g04076(.A(new_n6424), .B(new_n6397_1), .Y(new_n6425));
  nand_5 g04077(.A(new_n6425), .B(new_n6395), .Y(new_n6426));
  nand_5 g04078(.A(new_n6426), .B(new_n6393), .Y(new_n6427_1));
  nand_5 g04079(.A(new_n6427_1), .B(new_n6391), .Y(new_n6428));
  nand_5 g04080(.A(new_n6428), .B(new_n6389), .Y(new_n6429));
  nand_5 g04081(.A(new_n6429), .B(new_n6387), .Y(new_n6430));
  nand_5 g04082(.A(new_n6430), .B(new_n6385_1), .Y(new_n6431_1));
  nand_5 g04083(.A(new_n6431_1), .B(new_n6383_1), .Y(new_n6432));
  nand_5 g04084(.A(new_n6432), .B(new_n6381_1), .Y(new_n6433));
  nand_5 g04085(.A(new_n6385_1), .B(new_n6383_1), .Y(new_n6434));
  xor_4  g04086(.A(new_n6434), .B(new_n6430), .Y(new_n6435));
  nand_5 g04087(.A(new_n6281), .B(new_n6282), .Y(new_n6436));
  xor_4  g04088(.A(new_n6436), .B(new_n6366), .Y(new_n6437_1));
  nand_5 g04089(.A(new_n6437_1), .B(new_n6435), .Y(new_n6438));
  or_5   g04090(.A(new_n6437_1), .B(new_n6435), .Y(new_n6439));
  nand_5 g04091(.A(new_n6389), .B(new_n6387), .Y(new_n6440));
  xor_4  g04092(.A(new_n6440), .B(new_n6428), .Y(new_n6441));
  nand_5 g04093(.A(new_n6289), .B(new_n6288), .Y(new_n6442));
  xor_4  g04094(.A(new_n6442), .B(new_n6364), .Y(new_n6443));
  or_5   g04095(.A(new_n6443), .B(new_n6441), .Y(new_n6444));
  nand_5 g04096(.A(new_n6443), .B(new_n6441), .Y(new_n6445));
  nand_5 g04097(.A(new_n6393), .B(new_n6391), .Y(new_n6446));
  xor_4  g04098(.A(new_n6446), .B(new_n6426), .Y(new_n6447));
  nand_5 g04099(.A(new_n6297), .B(new_n6295), .Y(new_n6448));
  xor_4  g04100(.A(new_n6448), .B(new_n6362), .Y(new_n6449));
  or_5   g04101(.A(new_n6449), .B(new_n6447), .Y(new_n6450));
  nand_5 g04102(.A(new_n6449), .B(new_n6447), .Y(new_n6451));
  nand_5 g04103(.A(new_n6397_1), .B(new_n6395), .Y(new_n6452));
  xor_4  g04104(.A(new_n6452), .B(new_n6424), .Y(new_n6453));
  nand_5 g04105(.A(new_n6305), .B(new_n6303), .Y(new_n6454));
  xor_4  g04106(.A(new_n6454), .B(new_n6360), .Y(new_n6455));
  or_5   g04107(.A(new_n6455), .B(new_n6453), .Y(new_n6456_1));
  nand_5 g04108(.A(new_n6455), .B(new_n6453), .Y(new_n6457_1));
  nand_5 g04109(.A(new_n6400), .B(new_n6398), .Y(new_n6458));
  xor_4  g04110(.A(new_n6458), .B(new_n6422), .Y(new_n6459));
  nand_5 g04111(.A(new_n6313), .B(new_n6311_1), .Y(new_n6460));
  xor_4  g04112(.A(new_n6460), .B(new_n6358), .Y(new_n6461));
  or_5   g04113(.A(new_n6461), .B(new_n6459), .Y(new_n6462));
  nand_5 g04114(.A(new_n6461), .B(new_n6459), .Y(new_n6463));
  nand_5 g04115(.A(new_n6403), .B(new_n6401), .Y(new_n6464));
  xor_4  g04116(.A(new_n6464), .B(new_n6420), .Y(new_n6465_1));
  nand_5 g04117(.A(new_n6321), .B(new_n6319), .Y(new_n6466));
  xor_4  g04118(.A(new_n6466), .B(new_n6356_1), .Y(new_n6467));
  or_5   g04119(.A(new_n6467), .B(new_n6465_1), .Y(new_n6468));
  nand_5 g04120(.A(new_n6467), .B(new_n6465_1), .Y(new_n6469));
  nand_5 g04121(.A(new_n6406), .B(new_n6404), .Y(new_n6470_1));
  xor_4  g04122(.A(new_n6470_1), .B(new_n6418), .Y(new_n6471));
  nand_5 g04123(.A(new_n6327), .B(new_n6328), .Y(new_n6472));
  xor_4  g04124(.A(new_n6472), .B(new_n6354_1), .Y(new_n6473));
  or_5   g04125(.A(new_n6473), .B(new_n6471), .Y(new_n6474));
  nand_5 g04126(.A(new_n6473), .B(new_n6471), .Y(new_n6475));
  nand_5 g04127(.A(new_n6409), .B(new_n6407_1), .Y(new_n6476_1));
  xor_4  g04128(.A(new_n6476_1), .B(new_n6416), .Y(new_n6477));
  nand_5 g04129(.A(new_n6334), .B(new_n6335), .Y(new_n6478));
  xor_4  g04130(.A(new_n6478), .B(new_n6352), .Y(new_n6479));
  or_5   g04131(.A(new_n6479), .B(new_n6477), .Y(new_n6480));
  nand_5 g04132(.A(new_n6479), .B(new_n6477), .Y(new_n6481));
  not_8  g04133(.A(new_n6342), .Y(new_n6482));
  nor_5  g04134(.A(new_n6341), .B(new_n6338), .Y(new_n6483));
  nor_5  g04135(.A(new_n6483), .B(new_n6482), .Y(new_n6484));
  nand_5 g04136(.A(n12384), .B(new_n4541), .Y(new_n6485_1));
  nand_5 g04137(.A(new_n6485_1), .B(new_n6414), .Y(new_n6486));
  nand_5 g04138(.A(new_n6486), .B(new_n6484), .Y(new_n6487));
  not_8  g04139(.A(new_n6414), .Y(new_n6488));
  and_5  g04140(.A(new_n6412), .B(new_n6410), .Y(new_n6489));
  xor_4  g04141(.A(new_n6489), .B(new_n6488), .Y(new_n6490));
  or_5   g04142(.A(new_n6490), .B(new_n6487), .Y(new_n6491));
  nand_5 g04143(.A(new_n6490), .B(new_n6487), .Y(new_n6492));
  nand_5 g04144(.A(new_n6346), .B(new_n6347), .Y(new_n6493));
  xor_4  g04145(.A(new_n6493), .B(new_n6350), .Y(new_n6494));
  not_8  g04146(.A(new_n6494), .Y(new_n6495));
  nand_5 g04147(.A(new_n6495), .B(new_n6492), .Y(new_n6496));
  nand_5 g04148(.A(new_n6496), .B(new_n6491), .Y(new_n6497));
  nand_5 g04149(.A(new_n6497), .B(new_n6481), .Y(new_n6498));
  nand_5 g04150(.A(new_n6498), .B(new_n6480), .Y(new_n6499));
  nand_5 g04151(.A(new_n6499), .B(new_n6475), .Y(new_n6500));
  nand_5 g04152(.A(new_n6500), .B(new_n6474), .Y(new_n6501));
  nand_5 g04153(.A(new_n6501), .B(new_n6469), .Y(new_n6502_1));
  nand_5 g04154(.A(new_n6502_1), .B(new_n6468), .Y(new_n6503));
  nand_5 g04155(.A(new_n6503), .B(new_n6463), .Y(new_n6504));
  nand_5 g04156(.A(new_n6504), .B(new_n6462), .Y(new_n6505));
  nand_5 g04157(.A(new_n6505), .B(new_n6457_1), .Y(new_n6506_1));
  nand_5 g04158(.A(new_n6506_1), .B(new_n6456_1), .Y(new_n6507));
  nand_5 g04159(.A(new_n6507), .B(new_n6451), .Y(new_n6508));
  nand_5 g04160(.A(new_n6508), .B(new_n6450), .Y(new_n6509));
  nand_5 g04161(.A(new_n6509), .B(new_n6445), .Y(new_n6510));
  nand_5 g04162(.A(new_n6510), .B(new_n6444), .Y(new_n6511));
  not_8  g04163(.A(new_n6511), .Y(new_n6512));
  nand_5 g04164(.A(new_n6512), .B(new_n6439), .Y(new_n6513_1));
  nand_5 g04165(.A(new_n6513_1), .B(new_n6438), .Y(new_n6514_1));
  nor_5  g04166(.A(new_n6514_1), .B(new_n6433), .Y(new_n6515));
  nor_5  g04167(.A(new_n6432), .B(new_n6381_1), .Y(new_n6516));
  nand_5 g04168(.A(new_n6516), .B(new_n6514_1), .Y(new_n6517));
  not_8  g04169(.A(new_n6517), .Y(new_n6518));
  nor_5  g04170(.A(new_n6518), .B(new_n6515), .Y(new_n6519));
  nand_5 g04171(.A(new_n6379_1), .B(new_n6375_1), .Y(new_n6520));
  or_5   g04172(.A(new_n6379_1), .B(new_n6374), .Y(new_n6521));
  nand_5 g04173(.A(new_n6521), .B(new_n6520), .Y(new_n6522));
  not_8  g04174(.A(new_n6522), .Y(new_n6523));
  xor_4  g04175(.A(new_n6523), .B(new_n6519), .Y(n457));
  nand_5 g04176(.A(n13781), .B(n2088), .Y(new_n6525));
  nand_5 g04177(.A(new_n3089_1), .B(new_n3163), .Y(new_n6526));
  nand_5 g04178(.A(n9399), .B(n2088), .Y(new_n6527));
  and_5  g04179(.A(new_n6527), .B(new_n6526), .Y(new_n6528));
  not_8  g04180(.A(new_n6528), .Y(new_n6529));
  nand_5 g04181(.A(new_n6529), .B(new_n2383), .Y(new_n6530));
  nand_5 g04182(.A(new_n6528), .B(n11486), .Y(new_n6531));
  and_5  g04183(.A(new_n6531), .B(new_n6530), .Y(new_n6532));
  xor_4  g04184(.A(new_n6532), .B(new_n6525), .Y(new_n6533));
  not_8  g04185(.A(new_n6533), .Y(new_n6534));
  nand_5 g04186(.A(new_n2378), .B(new_n3163), .Y(new_n6535));
  and_5  g04187(.A(new_n6535), .B(new_n6525), .Y(new_n6536));
  not_8  g04188(.A(n24323), .Y(new_n6537));
  nand_5 g04189(.A(new_n6537), .B(n1681), .Y(new_n6538));
  nand_5 g04190(.A(n24323), .B(new_n2613), .Y(new_n6539));
  and_5  g04191(.A(new_n6539), .B(new_n6538), .Y(new_n6540));
  not_8  g04192(.A(new_n6540), .Y(new_n6541));
  nand_5 g04193(.A(new_n6541), .B(new_n6536), .Y(new_n6542_1));
  nand_5 g04194(.A(new_n4898), .B(n25877), .Y(new_n6543));
  not_8  g04195(.A(n25877), .Y(new_n6544));
  nand_5 g04196(.A(n26443), .B(new_n6544), .Y(new_n6545));
  nand_5 g04197(.A(new_n6545), .B(new_n6543), .Y(new_n6546));
  xnor_4 g04198(.A(new_n6546), .B(new_n6538), .Y(new_n6547));
  not_8  g04199(.A(new_n6547), .Y(new_n6548));
  nand_5 g04200(.A(new_n6548), .B(new_n6542_1), .Y(new_n6549));
  or_5   g04201(.A(new_n6548), .B(new_n6542_1), .Y(new_n6550));
  nand_5 g04202(.A(new_n6550), .B(new_n6549), .Y(new_n6551));
  xor_4  g04203(.A(new_n6551), .B(new_n6534), .Y(new_n6552));
  not_8  g04204(.A(new_n6536), .Y(new_n6553));
  xor_4  g04205(.A(new_n6540), .B(new_n6553), .Y(new_n6554));
  nand_5 g04206(.A(new_n6554), .B(new_n6338), .Y(new_n6555));
  nand_5 g04207(.A(new_n6555), .B(new_n6345), .Y(new_n6556_1));
  or_5   g04208(.A(new_n6555), .B(new_n6345), .Y(new_n6557));
  nand_5 g04209(.A(new_n6557), .B(new_n6556_1), .Y(new_n6558_1));
  xor_4  g04210(.A(new_n6558_1), .B(new_n6552), .Y(n463));
  nand_5 g04211(.A(n12121), .B(n6775), .Y(new_n6560_1));
  not_8  g04212(.A(n6775), .Y(new_n6561));
  nand_5 g04213(.A(new_n4084), .B(new_n6561), .Y(new_n6562));
  and_5  g04214(.A(new_n6562), .B(new_n6560_1), .Y(new_n6563));
  nand_5 g04215(.A(new_n6563), .B(n8920), .Y(new_n6564));
  not_8  g04216(.A(new_n6563), .Y(new_n6565));
  nand_5 g04217(.A(new_n6565), .B(new_n4653), .Y(new_n6566));
  and_5  g04218(.A(new_n6566), .B(new_n6564), .Y(new_n6567_1));
  not_8  g04219(.A(new_n6567_1), .Y(new_n6568));
  nand_5 g04220(.A(new_n3161_1), .B(n5438), .Y(new_n6569));
  nand_5 g04221(.A(new_n3162), .B(new_n3015), .Y(new_n6570));
  nand_5 g04222(.A(new_n6570), .B(new_n6569), .Y(new_n6571));
  xor_4  g04223(.A(new_n6571), .B(new_n6568), .Y(n491));
  nand_5 g04224(.A(new_n6475), .B(new_n6474), .Y(new_n6573));
  xnor_4 g04225(.A(new_n6573), .B(new_n6499), .Y(n496));
  not_8  g04226(.A(n16167), .Y(new_n6575));
  xor_4  g04227(.A(new_n6337), .B(new_n6575), .Y(new_n6576_1));
  nand_5 g04228(.A(n25926), .B(n12384), .Y(new_n6577));
  nand_5 g04229(.A(new_n4574), .B(new_n6413), .Y(new_n6578));
  and_5  g04230(.A(new_n6578), .B(new_n6577), .Y(new_n6579));
  nand_5 g04231(.A(new_n6579), .B(n6773), .Y(new_n6580));
  not_8  g04232(.A(new_n6580), .Y(new_n6581));
  nor_5  g04233(.A(new_n6579), .B(n6773), .Y(new_n6582));
  nor_5  g04234(.A(new_n6582), .B(new_n6581), .Y(new_n6583));
  nand_5 g04235(.A(new_n6583), .B(new_n6576_1), .Y(new_n6584));
  nand_5 g04236(.A(new_n4574), .B(new_n4346), .Y(new_n6585));
  nand_5 g04237(.A(n25926), .B(n7657), .Y(new_n6586));
  and_5  g04238(.A(new_n6586), .B(new_n6585), .Y(new_n6587_1));
  not_8  g04239(.A(new_n6587_1), .Y(new_n6588));
  nand_5 g04240(.A(new_n6588), .B(new_n6411), .Y(new_n6589));
  nand_5 g04241(.A(new_n6587_1), .B(n20986), .Y(new_n6590_1));
  nand_5 g04242(.A(new_n6590_1), .B(new_n6589), .Y(new_n6591));
  xor_4  g04243(.A(new_n6591), .B(new_n6577), .Y(new_n6592));
  nor_5  g04244(.A(n17090), .B(n6773), .Y(new_n6593));
  nor_5  g04245(.A(new_n4386), .B(new_n4541), .Y(new_n6594));
  nor_5  g04246(.A(new_n6594), .B(new_n6593), .Y(new_n6595));
  nor_5  g04247(.A(new_n6595), .B(new_n6581), .Y(new_n6596_1));
  nand_5 g04248(.A(new_n6581), .B(new_n4386), .Y(new_n6597));
  not_8  g04249(.A(new_n6597), .Y(new_n6598));
  nor_5  g04250(.A(new_n6598), .B(new_n6596_1), .Y(new_n6599));
  xor_4  g04251(.A(new_n6599), .B(new_n6592), .Y(new_n6600));
  nand_5 g04252(.A(new_n6338), .B(n16167), .Y(new_n6601));
  not_8  g04253(.A(n18745), .Y(new_n6602));
  nand_5 g04254(.A(new_n6345), .B(new_n6602), .Y(new_n6603));
  nand_5 g04255(.A(new_n6344), .B(n18745), .Y(new_n6604));
  nand_5 g04256(.A(new_n6604), .B(new_n6603), .Y(new_n6605));
  xor_4  g04257(.A(new_n6605), .B(new_n6601), .Y(new_n6606));
  or_5   g04258(.A(new_n6606), .B(new_n6600), .Y(new_n6607));
  nand_5 g04259(.A(new_n6606), .B(new_n6600), .Y(new_n6608));
  nand_5 g04260(.A(new_n6608), .B(new_n6607), .Y(new_n6609));
  xor_4  g04261(.A(new_n6609), .B(new_n6584), .Y(n498));
  nand_5 g04262(.A(n12121), .B(n3925), .Y(new_n6611_1));
  nand_5 g04263(.A(new_n4084), .B(new_n5549), .Y(new_n6612_1));
  nand_5 g04264(.A(new_n6612_1), .B(new_n6611_1), .Y(new_n6613));
  nand_5 g04265(.A(new_n6613), .B(new_n5471), .Y(new_n6614));
  nand_5 g04266(.A(new_n4085_1), .B(new_n5544), .Y(new_n6615));
  nand_5 g04267(.A(n22043), .B(n20259), .Y(new_n6616));
  nand_5 g04268(.A(new_n6616), .B(new_n6615), .Y(new_n6617));
  xnor_4 g04269(.A(new_n6617), .B(new_n6611_1), .Y(new_n6618));
  or_5   g04270(.A(new_n6618), .B(new_n5464), .Y(new_n6619));
  nand_5 g04271(.A(new_n6618), .B(new_n5464), .Y(new_n6620));
  nand_5 g04272(.A(new_n6620), .B(new_n6619), .Y(new_n6621));
  xor_4  g04273(.A(new_n6621), .B(new_n6614), .Y(new_n6622));
  or_5   g04274(.A(new_n6622), .B(new_n4204_1), .Y(new_n6623));
  nand_5 g04275(.A(new_n6622), .B(new_n4202), .Y(new_n6624));
  not_8  g04276(.A(new_n4209), .Y(new_n6625));
  xor_4  g04277(.A(new_n6613), .B(new_n5471), .Y(new_n6626));
  nor_5  g04278(.A(new_n6626), .B(new_n6625), .Y(new_n6627));
  nand_5 g04279(.A(new_n6627), .B(new_n6624), .Y(new_n6628_1));
  nand_5 g04280(.A(new_n6628_1), .B(new_n6623), .Y(new_n6629));
  nand_5 g04281(.A(new_n6620), .B(new_n6614), .Y(new_n6630_1));
  nand_5 g04282(.A(new_n6630_1), .B(new_n6619), .Y(new_n6631_1));
  nand_5 g04283(.A(new_n6616), .B(new_n6611_1), .Y(new_n6632));
  nand_5 g04284(.A(new_n6632), .B(new_n6615), .Y(new_n6633));
  nand_5 g04285(.A(new_n5538), .B(new_n4083), .Y(new_n6634_1));
  nand_5 g04286(.A(n25872), .B(n19618), .Y(new_n6635));
  nand_5 g04287(.A(new_n6635), .B(new_n6634_1), .Y(new_n6636));
  xor_4  g04288(.A(new_n6636), .B(new_n6633), .Y(new_n6637));
  nand_5 g04289(.A(new_n6637), .B(new_n5460), .Y(new_n6638));
  or_5   g04290(.A(new_n6637), .B(new_n5460), .Y(new_n6639));
  nand_5 g04291(.A(new_n6639), .B(new_n6638), .Y(new_n6640));
  xor_4  g04292(.A(new_n6640), .B(new_n6631_1), .Y(new_n6641));
  or_5   g04293(.A(new_n6641), .B(new_n4198), .Y(new_n6642));
  nand_5 g04294(.A(new_n6641), .B(new_n4198), .Y(new_n6643));
  nand_5 g04295(.A(new_n6643), .B(new_n6642), .Y(new_n6644));
  xnor_4 g04296(.A(new_n6644), .B(new_n6629), .Y(n521));
  xor_4  g04297(.A(new_n6486), .B(new_n6484), .Y(n548));
  nand_5 g04298(.A(new_n4735), .B(new_n4737), .Y(new_n6647));
  xor_4  g04299(.A(new_n6647), .B(new_n4762), .Y(n554));
  nand_5 g04300(.A(new_n5469), .B(new_n4201), .Y(new_n6649));
  not_8  g04301(.A(new_n6649), .Y(new_n6650));
  nand_5 g04302(.A(new_n6650), .B(new_n4195), .Y(new_n6651));
  nor_5  g04303(.A(new_n6651), .B(n4957), .Y(new_n6652_1));
  nand_5 g04304(.A(new_n6652_1), .B(new_n5384), .Y(new_n6653));
  nor_5  g04305(.A(new_n6653), .B(n3161), .Y(new_n6654));
  nand_5 g04306(.A(new_n6654), .B(new_n4293), .Y(new_n6655_1));
  nor_5  g04307(.A(new_n6655_1), .B(n20409), .Y(new_n6656));
  nand_5 g04308(.A(new_n6656), .B(new_n5370), .Y(new_n6657));
  nand_5 g04309(.A(new_n6657), .B(n2979), .Y(new_n6658));
  nor_5  g04310(.A(new_n6657), .B(n2979), .Y(new_n6659_1));
  not_8  g04311(.A(new_n6659_1), .Y(new_n6660));
  and_5  g04312(.A(new_n6660), .B(new_n6658), .Y(new_n6661));
  nand_5 g04313(.A(n9259), .B(n6456), .Y(new_n6662));
  not_8  g04314(.A(n6456), .Y(new_n6663));
  nand_5 g04315(.A(new_n5419), .B(new_n6663), .Y(new_n6664));
  nand_5 g04316(.A(new_n6664), .B(new_n6662), .Y(new_n6665));
  not_8  g04317(.A(n4085), .Y(new_n6666));
  nand_5 g04318(.A(new_n3694), .B(new_n6666), .Y(new_n6667));
  nand_5 g04319(.A(n21489), .B(n4085), .Y(new_n6668));
  not_8  g04320(.A(n26725), .Y(new_n6669_1));
  nand_5 g04321(.A(new_n6669_1), .B(new_n3778), .Y(new_n6670));
  nand_5 g04322(.A(n26725), .B(n20213), .Y(new_n6671_1));
  not_8  g04323(.A(n11980), .Y(new_n6672));
  nand_5 g04324(.A(new_n3695), .B(new_n6672), .Y(new_n6673_1));
  nand_5 g04325(.A(n13912), .B(n11980), .Y(new_n6674_1));
  not_8  g04326(.A(n3253), .Y(new_n6675));
  nand_5 g04327(.A(new_n3793), .B(new_n6675), .Y(new_n6676));
  nand_5 g04328(.A(n7670), .B(n3253), .Y(new_n6677));
  nand_5 g04329(.A(n9598), .B(n7759), .Y(new_n6678));
  not_8  g04330(.A(n7759), .Y(new_n6679));
  nand_5 g04331(.A(new_n3696), .B(new_n6679), .Y(new_n6680));
  not_8  g04332(.A(n12562), .Y(new_n6681));
  not_8  g04333(.A(n7949), .Y(new_n6682));
  nand_5 g04334(.A(new_n5457), .B(new_n6682), .Y(new_n6683));
  nand_5 g04335(.A(n11273), .B(n7949), .Y(new_n6684_1));
  not_8  g04336(.A(n24374), .Y(new_n6685));
  nand_5 g04337(.A(new_n3698), .B(new_n6685), .Y(new_n6686));
  nand_5 g04338(.A(n25565), .B(n24374), .Y(new_n6687));
  nand_5 g04339(.A(n21993), .B(n14575), .Y(new_n6688));
  nand_5 g04340(.A(new_n6688), .B(new_n6687), .Y(new_n6689));
  nand_5 g04341(.A(new_n6689), .B(new_n6686), .Y(new_n6690));
  nand_5 g04342(.A(new_n6690), .B(new_n6684_1), .Y(new_n6691_1));
  nand_5 g04343(.A(new_n6691_1), .B(new_n6683), .Y(new_n6692));
  nand_5 g04344(.A(new_n6692), .B(new_n6681), .Y(new_n6693));
  not_8  g04345(.A(new_n6693), .Y(new_n6694));
  nor_5  g04346(.A(new_n6692), .B(new_n6681), .Y(new_n6695));
  nor_5  g04347(.A(new_n6695), .B(n22290), .Y(new_n6696));
  nor_5  g04348(.A(new_n6696), .B(new_n6694), .Y(new_n6697));
  nand_5 g04349(.A(new_n6697), .B(new_n6680), .Y(new_n6698));
  and_5  g04350(.A(new_n6698), .B(new_n6678), .Y(new_n6699));
  nand_5 g04351(.A(new_n6699), .B(new_n6677), .Y(new_n6700));
  nand_5 g04352(.A(new_n6700), .B(new_n6676), .Y(new_n6701));
  nand_5 g04353(.A(new_n6701), .B(new_n6674_1), .Y(new_n6702));
  nand_5 g04354(.A(new_n6702), .B(new_n6673_1), .Y(new_n6703));
  nand_5 g04355(.A(new_n6703), .B(new_n6671_1), .Y(new_n6704));
  nand_5 g04356(.A(new_n6704), .B(new_n6670), .Y(new_n6705));
  nand_5 g04357(.A(new_n6705), .B(new_n6668), .Y(new_n6706_1));
  nand_5 g04358(.A(new_n6706_1), .B(new_n6667), .Y(new_n6707_1));
  xor_4  g04359(.A(new_n6707_1), .B(new_n6665), .Y(new_n6708));
  not_8  g04360(.A(new_n6708), .Y(new_n6709));
  nand_5 g04361(.A(new_n6709), .B(new_n6661), .Y(new_n6710));
  not_8  g04362(.A(new_n6661), .Y(new_n6711));
  nand_5 g04363(.A(new_n6708), .B(new_n6711), .Y(new_n6712));
  nand_5 g04364(.A(new_n6712), .B(new_n6710), .Y(new_n6713));
  xor_4  g04365(.A(new_n6656), .B(new_n5370), .Y(new_n6714));
  not_8  g04366(.A(new_n6714), .Y(new_n6715));
  nand_5 g04367(.A(new_n6668), .B(new_n6667), .Y(new_n6716));
  xor_4  g04368(.A(new_n6716), .B(new_n6705), .Y(new_n6717));
  nand_5 g04369(.A(new_n6717), .B(new_n6715), .Y(new_n6718));
  not_8  g04370(.A(new_n6717), .Y(new_n6719));
  nand_5 g04371(.A(new_n6719), .B(new_n6714), .Y(new_n6720));
  xor_4  g04372(.A(new_n6655_1), .B(n20409), .Y(new_n6721));
  not_8  g04373(.A(new_n6721), .Y(new_n6722));
  nand_5 g04374(.A(new_n6671_1), .B(new_n6670), .Y(new_n6723));
  xor_4  g04375(.A(new_n6723), .B(new_n6703), .Y(new_n6724));
  nand_5 g04376(.A(new_n6724), .B(new_n6722), .Y(new_n6725));
  not_8  g04377(.A(new_n6724), .Y(new_n6726));
  nand_5 g04378(.A(new_n6726), .B(new_n6721), .Y(new_n6727));
  xor_4  g04379(.A(new_n6654), .B(new_n4293), .Y(new_n6728));
  not_8  g04380(.A(new_n6728), .Y(new_n6729_1));
  nand_5 g04381(.A(new_n6674_1), .B(new_n6673_1), .Y(new_n6730));
  xor_4  g04382(.A(new_n6730), .B(new_n6701), .Y(new_n6731));
  nand_5 g04383(.A(new_n6731), .B(new_n6729_1), .Y(new_n6732));
  not_8  g04384(.A(new_n6731), .Y(new_n6733));
  nand_5 g04385(.A(new_n6733), .B(new_n6728), .Y(new_n6734));
  xor_4  g04386(.A(new_n6653), .B(n3161), .Y(new_n6735));
  not_8  g04387(.A(new_n6735), .Y(new_n6736_1));
  nand_5 g04388(.A(new_n6677), .B(new_n6676), .Y(new_n6737));
  xor_4  g04389(.A(new_n6737), .B(new_n6699), .Y(new_n6738));
  nand_5 g04390(.A(new_n6738), .B(new_n6736_1), .Y(new_n6739));
  not_8  g04391(.A(new_n6738), .Y(new_n6740));
  nand_5 g04392(.A(new_n6740), .B(new_n6735), .Y(new_n6741));
  xor_4  g04393(.A(new_n6652_1), .B(new_n5384), .Y(new_n6742));
  not_8  g04394(.A(new_n6742), .Y(new_n6743));
  nand_5 g04395(.A(new_n6680), .B(new_n6678), .Y(new_n6744));
  xor_4  g04396(.A(new_n6744), .B(new_n6697), .Y(new_n6745));
  not_8  g04397(.A(new_n6745), .Y(new_n6746));
  nand_5 g04398(.A(new_n6746), .B(new_n6743), .Y(new_n6747));
  nand_5 g04399(.A(new_n6745), .B(new_n6742), .Y(new_n6748));
  xor_4  g04400(.A(new_n6651), .B(n4957), .Y(new_n6749));
  not_8  g04401(.A(new_n6749), .Y(new_n6750));
  nor_5  g04402(.A(new_n6695), .B(new_n6694), .Y(new_n6751));
  xor_4  g04403(.A(new_n6751), .B(new_n5451_1), .Y(new_n6752));
  not_8  g04404(.A(new_n6752), .Y(new_n6753));
  nand_5 g04405(.A(new_n6753), .B(new_n6750), .Y(new_n6754));
  nand_5 g04406(.A(new_n6752), .B(new_n6749), .Y(new_n6755));
  nand_5 g04407(.A(new_n6649), .B(n7524), .Y(new_n6756));
  and_5  g04408(.A(new_n6756), .B(new_n6651), .Y(new_n6757));
  not_8  g04409(.A(new_n6757), .Y(new_n6758));
  nand_5 g04410(.A(new_n6684_1), .B(new_n6683), .Y(new_n6759));
  xor_4  g04411(.A(new_n6759), .B(new_n6690), .Y(new_n6760));
  nand_5 g04412(.A(new_n6760), .B(new_n6758), .Y(new_n6761));
  not_8  g04413(.A(new_n6760), .Y(new_n6762));
  nand_5 g04414(.A(new_n6762), .B(new_n6757), .Y(new_n6763));
  not_8  g04415(.A(n14575), .Y(new_n6764));
  nand_5 g04416(.A(new_n3697), .B(new_n6764), .Y(new_n6765));
  nand_5 g04417(.A(new_n6765), .B(new_n6688), .Y(new_n6766));
  not_8  g04418(.A(new_n6766), .Y(new_n6767));
  nand_5 g04419(.A(new_n6767), .B(new_n5469), .Y(new_n6768));
  nand_5 g04420(.A(n20658), .B(n15743), .Y(new_n6769));
  and_5  g04421(.A(new_n6769), .B(new_n6649), .Y(new_n6770));
  nand_5 g04422(.A(new_n6770), .B(new_n6768), .Y(new_n6771));
  nand_5 g04423(.A(new_n6687), .B(new_n6686), .Y(new_n6772));
  not_8  g04424(.A(new_n6772), .Y(new_n6773_1));
  xor_4  g04425(.A(new_n6773_1), .B(new_n6688), .Y(new_n6774));
  nand_5 g04426(.A(new_n6767), .B(new_n6650), .Y(new_n6775_1));
  nand_5 g04427(.A(new_n6775_1), .B(new_n6774), .Y(new_n6776));
  nand_5 g04428(.A(new_n6776), .B(new_n6771), .Y(new_n6777));
  not_8  g04429(.A(new_n6777), .Y(new_n6778));
  nand_5 g04430(.A(new_n6778), .B(new_n6763), .Y(new_n6779));
  nand_5 g04431(.A(new_n6779), .B(new_n6761), .Y(new_n6780));
  nand_5 g04432(.A(new_n6780), .B(new_n6755), .Y(new_n6781));
  nand_5 g04433(.A(new_n6781), .B(new_n6754), .Y(new_n6782));
  nand_5 g04434(.A(new_n6782), .B(new_n6748), .Y(new_n6783));
  nand_5 g04435(.A(new_n6783), .B(new_n6747), .Y(new_n6784));
  nand_5 g04436(.A(new_n6784), .B(new_n6741), .Y(new_n6785_1));
  nand_5 g04437(.A(new_n6785_1), .B(new_n6739), .Y(new_n6786));
  nand_5 g04438(.A(new_n6786), .B(new_n6734), .Y(new_n6787));
  nand_5 g04439(.A(new_n6787), .B(new_n6732), .Y(new_n6788));
  nand_5 g04440(.A(new_n6788), .B(new_n6727), .Y(new_n6789));
  nand_5 g04441(.A(new_n6789), .B(new_n6725), .Y(new_n6790_1));
  nand_5 g04442(.A(new_n6790_1), .B(new_n6720), .Y(new_n6791_1));
  nand_5 g04443(.A(new_n6791_1), .B(new_n6718), .Y(new_n6792));
  xor_4  g04444(.A(new_n6792), .B(new_n6713), .Y(new_n6793));
  nand_5 g04445(.A(n21784), .B(n3582), .Y(new_n6794_1));
  not_8  g04446(.A(n3582), .Y(new_n6795));
  not_8  g04447(.A(n21784), .Y(new_n6796));
  nand_5 g04448(.A(new_n6796), .B(new_n6795), .Y(new_n6797));
  nand_5 g04449(.A(new_n6797), .B(new_n6794_1), .Y(new_n6798));
  not_8  g04450(.A(n2145), .Y(new_n6799));
  not_8  g04451(.A(n5521), .Y(new_n6800));
  nand_5 g04452(.A(new_n6800), .B(new_n6799), .Y(new_n6801));
  nand_5 g04453(.A(n5521), .B(n2145), .Y(new_n6802_1));
  not_8  g04454(.A(n5031), .Y(new_n6803));
  not_8  g04455(.A(n11926), .Y(new_n6804));
  nand_5 g04456(.A(new_n6804), .B(new_n6803), .Y(new_n6805));
  nand_5 g04457(.A(n11926), .B(n5031), .Y(new_n6806));
  not_8  g04458(.A(n4325), .Y(new_n6807));
  not_8  g04459(.A(n11044), .Y(new_n6808));
  nand_5 g04460(.A(new_n6808), .B(new_n6807), .Y(new_n6809));
  nand_5 g04461(.A(n11044), .B(n4325), .Y(new_n6810));
  not_8  g04462(.A(n2421), .Y(new_n6811));
  nand_5 g04463(.A(new_n4137), .B(new_n6811), .Y(new_n6812));
  nand_5 g04464(.A(n5337), .B(n2421), .Y(new_n6813));
  not_8  g04465(.A(n987), .Y(new_n6814_1));
  nand_5 g04466(.A(new_n6814_1), .B(new_n4082), .Y(new_n6815));
  nand_5 g04467(.A(n987), .B(n626), .Y(new_n6816));
  not_8  g04468(.A(n20478), .Y(new_n6817));
  nand_5 g04469(.A(new_n6817), .B(new_n4098), .Y(new_n6818));
  nand_5 g04470(.A(n20478), .B(n1204), .Y(new_n6819));
  not_8  g04471(.A(n26882), .Y(new_n6820));
  nand_5 g04472(.A(new_n6820), .B(new_n4083), .Y(new_n6821));
  nand_5 g04473(.A(n26882), .B(n19618), .Y(new_n6822));
  not_8  g04474(.A(n22619), .Y(new_n6823));
  nand_5 g04475(.A(new_n6823), .B(new_n4085_1), .Y(new_n6824));
  nand_5 g04476(.A(n22619), .B(n22043), .Y(new_n6825));
  nand_5 g04477(.A(new_n6825), .B(new_n6560_1), .Y(new_n6826_1));
  nand_5 g04478(.A(new_n6826_1), .B(new_n6824), .Y(new_n6827));
  nand_5 g04479(.A(new_n6827), .B(new_n6822), .Y(new_n6828));
  nand_5 g04480(.A(new_n6828), .B(new_n6821), .Y(new_n6829));
  nand_5 g04481(.A(new_n6829), .B(new_n6819), .Y(new_n6830));
  nand_5 g04482(.A(new_n6830), .B(new_n6818), .Y(new_n6831));
  nand_5 g04483(.A(new_n6831), .B(new_n6816), .Y(new_n6832));
  nand_5 g04484(.A(new_n6832), .B(new_n6815), .Y(new_n6833));
  nand_5 g04485(.A(new_n6833), .B(new_n6813), .Y(new_n6834));
  nand_5 g04486(.A(new_n6834), .B(new_n6812), .Y(new_n6835_1));
  nand_5 g04487(.A(new_n6835_1), .B(new_n6810), .Y(new_n6836));
  nand_5 g04488(.A(new_n6836), .B(new_n6809), .Y(new_n6837));
  nand_5 g04489(.A(new_n6837), .B(new_n6806), .Y(new_n6838));
  nand_5 g04490(.A(new_n6838), .B(new_n6805), .Y(new_n6839));
  nand_5 g04491(.A(new_n6839), .B(new_n6802_1), .Y(new_n6840));
  nand_5 g04492(.A(new_n6840), .B(new_n6801), .Y(new_n6841));
  not_8  g04493(.A(new_n6841), .Y(new_n6842));
  xor_4  g04494(.A(new_n6842), .B(new_n6798), .Y(new_n6843));
  not_8  g04495(.A(new_n6843), .Y(new_n6844));
  nand_5 g04496(.A(new_n6844), .B(n8526), .Y(new_n6845));
  not_8  g04497(.A(n8526), .Y(new_n6846));
  nand_5 g04498(.A(new_n6843), .B(new_n6846), .Y(new_n6847));
  nand_5 g04499(.A(new_n6847), .B(new_n6845), .Y(new_n6848));
  not_8  g04500(.A(n2816), .Y(new_n6849));
  nand_5 g04501(.A(new_n6802_1), .B(new_n6801), .Y(new_n6850));
  xor_4  g04502(.A(new_n6850), .B(new_n6839), .Y(new_n6851));
  not_8  g04503(.A(new_n6851), .Y(new_n6852));
  nand_5 g04504(.A(new_n6852), .B(new_n6849), .Y(new_n6853_1));
  nand_5 g04505(.A(new_n6851), .B(n2816), .Y(new_n6854));
  not_8  g04506(.A(n20359), .Y(new_n6855));
  nand_5 g04507(.A(new_n6806), .B(new_n6805), .Y(new_n6856));
  xor_4  g04508(.A(new_n6856), .B(new_n6837), .Y(new_n6857));
  not_8  g04509(.A(new_n6857), .Y(new_n6858));
  nand_5 g04510(.A(new_n6858), .B(new_n6855), .Y(new_n6859));
  nand_5 g04511(.A(new_n6857), .B(n20359), .Y(new_n6860));
  not_8  g04512(.A(n4409), .Y(new_n6861_1));
  nand_5 g04513(.A(new_n6810), .B(new_n6809), .Y(new_n6862_1));
  xor_4  g04514(.A(new_n6862_1), .B(new_n6835_1), .Y(new_n6863_1));
  not_8  g04515(.A(new_n6863_1), .Y(new_n6864));
  nand_5 g04516(.A(new_n6864), .B(new_n6861_1), .Y(new_n6865));
  nand_5 g04517(.A(new_n6863_1), .B(n4409), .Y(new_n6866));
  not_8  g04518(.A(n3570), .Y(new_n6867_1));
  nand_5 g04519(.A(new_n6813), .B(new_n6812), .Y(new_n6868));
  xor_4  g04520(.A(new_n6868), .B(new_n6833), .Y(new_n6869));
  not_8  g04521(.A(new_n6869), .Y(new_n6870));
  nand_5 g04522(.A(new_n6870), .B(new_n6867_1), .Y(new_n6871));
  nand_5 g04523(.A(new_n6869), .B(n3570), .Y(new_n6872));
  nand_5 g04524(.A(new_n6816), .B(new_n6815), .Y(new_n6873));
  xor_4  g04525(.A(new_n6873), .B(new_n6831), .Y(new_n6874));
  not_8  g04526(.A(new_n6874), .Y(new_n6875));
  nand_5 g04527(.A(new_n6875), .B(new_n4782), .Y(new_n6876));
  nand_5 g04528(.A(new_n6874), .B(n13668), .Y(new_n6877));
  not_8  g04529(.A(n21276), .Y(new_n6878));
  nand_5 g04530(.A(new_n6819), .B(new_n6818), .Y(new_n6879));
  xor_4  g04531(.A(new_n6879), .B(new_n6829), .Y(new_n6880));
  not_8  g04532(.A(new_n6880), .Y(new_n6881));
  nand_5 g04533(.A(new_n6881), .B(new_n6878), .Y(new_n6882));
  nand_5 g04534(.A(new_n6880), .B(n21276), .Y(new_n6883));
  not_8  g04535(.A(n26748), .Y(new_n6884));
  nand_5 g04536(.A(new_n6822), .B(new_n6821), .Y(new_n6885));
  xor_4  g04537(.A(new_n6885), .B(new_n6827), .Y(new_n6886));
  not_8  g04538(.A(new_n6886), .Y(new_n6887));
  nand_5 g04539(.A(new_n6887), .B(new_n6884), .Y(new_n6888));
  nand_5 g04540(.A(new_n6886), .B(n26748), .Y(new_n6889));
  nand_5 g04541(.A(new_n6825), .B(new_n6824), .Y(new_n6890));
  xor_4  g04542(.A(new_n6890), .B(new_n6560_1), .Y(new_n6891));
  not_8  g04543(.A(new_n6891), .Y(new_n6892));
  nand_5 g04544(.A(new_n6892), .B(new_n4654), .Y(new_n6893));
  nand_5 g04545(.A(new_n6891), .B(n10057), .Y(new_n6894));
  nand_5 g04546(.A(new_n6894), .B(new_n6564), .Y(new_n6895));
  nand_5 g04547(.A(new_n6895), .B(new_n6893), .Y(new_n6896));
  nand_5 g04548(.A(new_n6896), .B(new_n6889), .Y(new_n6897));
  nand_5 g04549(.A(new_n6897), .B(new_n6888), .Y(new_n6898));
  nand_5 g04550(.A(new_n6898), .B(new_n6883), .Y(new_n6899));
  nand_5 g04551(.A(new_n6899), .B(new_n6882), .Y(new_n6900));
  nand_5 g04552(.A(new_n6900), .B(new_n6877), .Y(new_n6901));
  nand_5 g04553(.A(new_n6901), .B(new_n6876), .Y(new_n6902));
  nand_5 g04554(.A(new_n6902), .B(new_n6872), .Y(new_n6903));
  nand_5 g04555(.A(new_n6903), .B(new_n6871), .Y(new_n6904));
  nand_5 g04556(.A(new_n6904), .B(new_n6866), .Y(new_n6905));
  nand_5 g04557(.A(new_n6905), .B(new_n6865), .Y(new_n6906));
  nand_5 g04558(.A(new_n6906), .B(new_n6860), .Y(new_n6907));
  nand_5 g04559(.A(new_n6907), .B(new_n6859), .Y(new_n6908));
  nand_5 g04560(.A(new_n6908), .B(new_n6854), .Y(new_n6909));
  nand_5 g04561(.A(new_n6909), .B(new_n6853_1), .Y(new_n6910));
  xor_4  g04562(.A(new_n6910), .B(new_n6848), .Y(new_n6911));
  nand_5 g04563(.A(new_n6911), .B(new_n6793), .Y(new_n6912));
  or_5   g04564(.A(new_n6911), .B(new_n6793), .Y(new_n6913));
  nand_5 g04565(.A(new_n6913), .B(new_n6912), .Y(new_n6914));
  nand_5 g04566(.A(new_n6853_1), .B(new_n6854), .Y(new_n6915));
  xor_4  g04567(.A(new_n6915), .B(new_n6908), .Y(new_n6916));
  nand_5 g04568(.A(new_n6720), .B(new_n6718), .Y(new_n6917));
  xor_4  g04569(.A(new_n6917), .B(new_n6790_1), .Y(new_n6918));
  nand_5 g04570(.A(new_n6918), .B(new_n6916), .Y(new_n6919));
  nor_5  g04571(.A(new_n6918), .B(new_n6916), .Y(new_n6920));
  not_8  g04572(.A(new_n6920), .Y(new_n6921));
  nand_5 g04573(.A(new_n6859), .B(new_n6860), .Y(new_n6922));
  xor_4  g04574(.A(new_n6922), .B(new_n6906), .Y(new_n6923));
  nand_5 g04575(.A(new_n6727), .B(new_n6725), .Y(new_n6924));
  xor_4  g04576(.A(new_n6924), .B(new_n6788), .Y(new_n6925));
  nand_5 g04577(.A(new_n6925), .B(new_n6923), .Y(new_n6926));
  nor_5  g04578(.A(new_n6925), .B(new_n6923), .Y(new_n6927));
  not_8  g04579(.A(new_n6927), .Y(new_n6928));
  nand_5 g04580(.A(new_n6865), .B(new_n6866), .Y(new_n6929));
  xor_4  g04581(.A(new_n6929), .B(new_n6904), .Y(new_n6930));
  nand_5 g04582(.A(new_n6734), .B(new_n6732), .Y(new_n6931));
  xor_4  g04583(.A(new_n6931), .B(new_n6786), .Y(new_n6932));
  nand_5 g04584(.A(new_n6932), .B(new_n6930), .Y(new_n6933));
  nor_5  g04585(.A(new_n6932), .B(new_n6930), .Y(new_n6934));
  not_8  g04586(.A(new_n6934), .Y(new_n6935));
  nand_5 g04587(.A(new_n6871), .B(new_n6872), .Y(new_n6936));
  xor_4  g04588(.A(new_n6936), .B(new_n6902), .Y(new_n6937));
  nand_5 g04589(.A(new_n6741), .B(new_n6739), .Y(new_n6938));
  xor_4  g04590(.A(new_n6938), .B(new_n6784), .Y(new_n6939));
  nand_5 g04591(.A(new_n6939), .B(new_n6937), .Y(new_n6940));
  nor_5  g04592(.A(new_n6939), .B(new_n6937), .Y(new_n6941));
  nand_5 g04593(.A(new_n6876), .B(new_n6877), .Y(new_n6942));
  xor_4  g04594(.A(new_n6942), .B(new_n6900), .Y(new_n6943));
  nand_5 g04595(.A(new_n6748), .B(new_n6747), .Y(new_n6944));
  xor_4  g04596(.A(new_n6944), .B(new_n6782), .Y(new_n6945));
  nand_5 g04597(.A(new_n6945), .B(new_n6943), .Y(new_n6946));
  not_8  g04598(.A(new_n6946), .Y(new_n6947));
  nor_5  g04599(.A(new_n6945), .B(new_n6943), .Y(new_n6948));
  nand_5 g04600(.A(new_n6882), .B(new_n6883), .Y(new_n6949));
  xor_4  g04601(.A(new_n6949), .B(new_n6898), .Y(new_n6950));
  nand_5 g04602(.A(new_n6755), .B(new_n6754), .Y(new_n6951));
  xor_4  g04603(.A(new_n6951), .B(new_n6780), .Y(new_n6952));
  nand_5 g04604(.A(new_n6952), .B(new_n6950), .Y(new_n6953));
  or_5   g04605(.A(new_n6952), .B(new_n6950), .Y(new_n6954));
  nand_5 g04606(.A(new_n6888), .B(new_n6889), .Y(new_n6955));
  xor_4  g04607(.A(new_n6955), .B(new_n6896), .Y(new_n6956));
  nand_5 g04608(.A(new_n6763), .B(new_n6761), .Y(new_n6957));
  xor_4  g04609(.A(new_n6957), .B(new_n6778), .Y(new_n6958));
  or_5   g04610(.A(new_n6958), .B(new_n6956), .Y(new_n6959));
  nand_5 g04611(.A(new_n6958), .B(new_n6956), .Y(new_n6960));
  nand_5 g04612(.A(new_n6893), .B(new_n6894), .Y(new_n6961));
  xor_4  g04613(.A(new_n6961), .B(new_n6564), .Y(new_n6962));
  not_8  g04614(.A(new_n6962), .Y(new_n6963));
  not_8  g04615(.A(new_n6774), .Y(new_n6964));
  and_5  g04616(.A(new_n6775_1), .B(new_n6771), .Y(new_n6965_1));
  xor_4  g04617(.A(new_n6965_1), .B(new_n6964), .Y(new_n6966));
  or_5   g04618(.A(new_n6966), .B(new_n6963), .Y(new_n6967_1));
  nand_5 g04619(.A(new_n6966), .B(new_n6963), .Y(new_n6968));
  xor_4  g04620(.A(new_n6766), .B(n20658), .Y(new_n6969));
  nor_5  g04621(.A(new_n6969), .B(new_n6568), .Y(new_n6970));
  nand_5 g04622(.A(new_n6970), .B(new_n6968), .Y(new_n6971_1));
  nand_5 g04623(.A(new_n6971_1), .B(new_n6967_1), .Y(new_n6972));
  not_8  g04624(.A(new_n6972), .Y(new_n6973));
  nand_5 g04625(.A(new_n6973), .B(new_n6960), .Y(new_n6974));
  and_5  g04626(.A(new_n6974), .B(new_n6959), .Y(new_n6975_1));
  nand_5 g04627(.A(new_n6975_1), .B(new_n6954), .Y(new_n6976));
  nand_5 g04628(.A(new_n6976), .B(new_n6953), .Y(new_n6977));
  not_8  g04629(.A(new_n6977), .Y(new_n6978));
  nor_5  g04630(.A(new_n6978), .B(new_n6948), .Y(new_n6979));
  nor_5  g04631(.A(new_n6979), .B(new_n6947), .Y(new_n6980));
  or_5   g04632(.A(new_n6980), .B(new_n6941), .Y(new_n6981));
  nand_5 g04633(.A(new_n6981), .B(new_n6940), .Y(new_n6982));
  nand_5 g04634(.A(new_n6982), .B(new_n6935), .Y(new_n6983_1));
  nand_5 g04635(.A(new_n6983_1), .B(new_n6933), .Y(new_n6984));
  nand_5 g04636(.A(new_n6984), .B(new_n6928), .Y(new_n6985_1));
  nand_5 g04637(.A(new_n6985_1), .B(new_n6926), .Y(new_n6986));
  nand_5 g04638(.A(new_n6986), .B(new_n6921), .Y(new_n6987));
  nand_5 g04639(.A(new_n6987), .B(new_n6919), .Y(new_n6988));
  not_8  g04640(.A(new_n6988), .Y(new_n6989));
  xor_4  g04641(.A(new_n6989), .B(new_n6914), .Y(n567));
  not_8  g04642(.A(n7674), .Y(new_n6991));
  not_8  g04643(.A(n13137), .Y(new_n6992));
  nand_5 g04644(.A(new_n6992), .B(new_n6991), .Y(new_n6993));
  not_8  g04645(.A(new_n6993), .Y(new_n6994));
  nand_5 g04646(.A(n13137), .B(n7674), .Y(new_n6995));
  not_8  g04647(.A(new_n6995), .Y(new_n6996));
  not_8  g04648(.A(n6397), .Y(new_n6997));
  not_8  g04649(.A(n18452), .Y(new_n6998_1));
  nand_5 g04650(.A(new_n6998_1), .B(new_n6997), .Y(new_n6999));
  not_8  g04651(.A(new_n6999), .Y(new_n7000));
  nand_5 g04652(.A(n18452), .B(n6397), .Y(new_n7001));
  not_8  g04653(.A(new_n7001), .Y(new_n7002));
  not_8  g04654(.A(n19196), .Y(new_n7003));
  not_8  g04655(.A(n21317), .Y(new_n7004));
  nand_5 g04656(.A(new_n7004), .B(new_n7003), .Y(new_n7005));
  not_8  g04657(.A(new_n7005), .Y(new_n7006));
  nand_5 g04658(.A(n21317), .B(n19196), .Y(new_n7007));
  not_8  g04659(.A(new_n7007), .Y(new_n7008));
  not_8  g04660(.A(n21226), .Y(new_n7009));
  nand_5 g04661(.A(new_n7009), .B(new_n4523), .Y(new_n7010));
  nand_5 g04662(.A(n21226), .B(n19789), .Y(new_n7011));
  not_8  g04663(.A(n4426), .Y(new_n7012));
  nand_5 g04664(.A(new_n4407), .B(new_n7012), .Y(new_n7013));
  nand_5 g04665(.A(n20169), .B(n4426), .Y(new_n7014));
  nand_5 g04666(.A(new_n4606), .B(new_n4408), .Y(new_n7015));
  nand_5 g04667(.A(n20036), .B(n8285), .Y(new_n7016));
  nand_5 g04668(.A(new_n4561), .B(new_n4422), .Y(new_n7017));
  nand_5 g04669(.A(n11192), .B(n6729), .Y(new_n7018));
  nand_5 g04670(.A(n21687), .B(n9380), .Y(new_n7019));
  nand_5 g04671(.A(new_n7019), .B(new_n7018), .Y(new_n7020));
  nand_5 g04672(.A(new_n7020), .B(new_n7017), .Y(new_n7021));
  nand_5 g04673(.A(new_n7021), .B(new_n7016), .Y(new_n7022));
  nand_5 g04674(.A(new_n7022), .B(new_n7015), .Y(new_n7023));
  nand_5 g04675(.A(new_n7023), .B(new_n7014), .Y(new_n7024));
  nand_5 g04676(.A(new_n7024), .B(new_n7013), .Y(new_n7025));
  nand_5 g04677(.A(new_n7025), .B(new_n7011), .Y(new_n7026_1));
  nand_5 g04678(.A(new_n7026_1), .B(new_n7010), .Y(new_n7027));
  nand_5 g04679(.A(new_n7027), .B(new_n4522), .Y(new_n7028));
  not_8  g04680(.A(new_n7028), .Y(new_n7029));
  nor_5  g04681(.A(new_n7027), .B(new_n4522), .Y(new_n7030));
  nor_5  g04682(.A(new_n7030), .B(n23586), .Y(new_n7031));
  nor_5  g04683(.A(new_n7031), .B(new_n7029), .Y(new_n7032_1));
  nor_5  g04684(.A(new_n7032_1), .B(new_n7008), .Y(new_n7033));
  nor_5  g04685(.A(new_n7033), .B(new_n7006), .Y(new_n7034));
  nor_5  g04686(.A(new_n7034), .B(new_n7002), .Y(new_n7035));
  nor_5  g04687(.A(new_n7035), .B(new_n7000), .Y(new_n7036));
  nor_5  g04688(.A(new_n7036), .B(new_n6996), .Y(new_n7037));
  nor_5  g04689(.A(new_n7037), .B(new_n6994), .Y(new_n7038_1));
  or_5   g04690(.A(new_n7038_1), .B(n1831), .Y(new_n7039));
  not_8  g04691(.A(n10250), .Y(new_n7040));
  nand_5 g04692(.A(new_n7038_1), .B(n1831), .Y(new_n7041));
  nand_5 g04693(.A(new_n7041), .B(new_n7040), .Y(new_n7042));
  nand_5 g04694(.A(new_n7042), .B(new_n7039), .Y(new_n7043));
  not_8  g04695(.A(new_n7043), .Y(new_n7044));
  not_8  g04696(.A(n1288), .Y(new_n7045));
  not_8  g04697(.A(n13110), .Y(new_n7046));
  nand_5 g04698(.A(new_n4513), .B(new_n7046), .Y(new_n7047));
  nor_5  g04699(.A(new_n7047), .B(n1752), .Y(new_n7048));
  nand_5 g04700(.A(new_n7048), .B(new_n7045), .Y(new_n7049));
  nand_5 g04701(.A(new_n7049), .B(n3320), .Y(new_n7050));
  nor_5  g04702(.A(new_n7049), .B(n3320), .Y(new_n7051));
  not_8  g04703(.A(new_n7051), .Y(new_n7052));
  and_5  g04704(.A(new_n7052), .B(new_n7050), .Y(new_n7053));
  not_8  g04705(.A(new_n7053), .Y(new_n7054));
  nand_5 g04706(.A(new_n7054), .B(new_n6382), .Y(new_n7055));
  not_8  g04707(.A(new_n7055), .Y(new_n7056));
  xor_4  g04708(.A(new_n7048), .B(n1288), .Y(new_n7057_1));
  nand_5 g04709(.A(new_n7057_1), .B(new_n6386), .Y(new_n7058));
  not_8  g04710(.A(new_n7057_1), .Y(new_n7059));
  nand_5 g04711(.A(new_n7059), .B(n15182), .Y(new_n7060));
  not_8  g04712(.A(n1752), .Y(new_n7061));
  xor_4  g04713(.A(new_n7047), .B(new_n7061), .Y(new_n7062));
  nand_5 g04714(.A(new_n7062), .B(new_n6390), .Y(new_n7063));
  not_8  g04715(.A(new_n7062), .Y(new_n7064));
  nand_5 g04716(.A(new_n7064), .B(n27037), .Y(new_n7065));
  nand_5 g04717(.A(new_n4514_1), .B(n13110), .Y(new_n7066));
  and_5  g04718(.A(new_n7066), .B(new_n7047), .Y(new_n7067));
  not_8  g04719(.A(new_n7067), .Y(new_n7068));
  nand_5 g04720(.A(new_n7068), .B(new_n6394), .Y(new_n7069));
  nand_5 g04721(.A(new_n7067), .B(n8964), .Y(new_n7070));
  nand_5 g04722(.A(new_n4519), .B(new_n4511), .Y(new_n7071));
  nand_5 g04723(.A(new_n7071), .B(new_n4518), .Y(new_n7072));
  nand_5 g04724(.A(new_n7072), .B(new_n7070), .Y(new_n7073));
  nand_5 g04725(.A(new_n7073), .B(new_n7069), .Y(new_n7074));
  nand_5 g04726(.A(new_n7074), .B(new_n7065), .Y(new_n7075));
  nand_5 g04727(.A(new_n7075), .B(new_n7063), .Y(new_n7076));
  nand_5 g04728(.A(new_n7076), .B(new_n7060), .Y(new_n7077));
  nand_5 g04729(.A(new_n7077), .B(new_n7058), .Y(new_n7078));
  nor_5  g04730(.A(new_n7078), .B(new_n7056), .Y(new_n7079_1));
  nand_5 g04731(.A(new_n7053), .B(n8614), .Y(new_n7080));
  nand_5 g04732(.A(new_n7080), .B(new_n7052), .Y(new_n7081));
  nor_5  g04733(.A(new_n7081), .B(new_n7079_1), .Y(new_n7082));
  or_5   g04734(.A(new_n7082), .B(new_n7044), .Y(new_n7083));
  nand_5 g04735(.A(new_n7082), .B(new_n7044), .Y(new_n7084));
  nand_5 g04736(.A(new_n7084), .B(new_n7083), .Y(new_n7085));
  nand_5 g04737(.A(new_n7041), .B(new_n7039), .Y(new_n7086));
  xor_4  g04738(.A(new_n7086), .B(n10250), .Y(new_n7087));
  nand_5 g04739(.A(new_n7080), .B(new_n7055), .Y(new_n7088));
  xor_4  g04740(.A(new_n7088), .B(new_n7078), .Y(new_n7089));
  not_8  g04741(.A(new_n7089), .Y(new_n7090));
  nand_5 g04742(.A(new_n7090), .B(new_n7087), .Y(new_n7091));
  not_8  g04743(.A(new_n7087), .Y(new_n7092));
  nand_5 g04744(.A(new_n7089), .B(new_n7092), .Y(new_n7093));
  nand_5 g04745(.A(new_n6995), .B(new_n6993), .Y(new_n7094));
  xor_4  g04746(.A(new_n7094), .B(new_n7036), .Y(new_n7095));
  nand_5 g04747(.A(new_n7060), .B(new_n7058), .Y(new_n7096));
  xor_4  g04748(.A(new_n7096), .B(new_n7076), .Y(new_n7097));
  not_8  g04749(.A(new_n7097), .Y(new_n7098));
  nand_5 g04750(.A(new_n7098), .B(new_n7095), .Y(new_n7099_1));
  not_8  g04751(.A(new_n7095), .Y(new_n7100));
  nand_5 g04752(.A(new_n7097), .B(new_n7100), .Y(new_n7101));
  nand_5 g04753(.A(new_n7001), .B(new_n6999), .Y(new_n7102));
  xor_4  g04754(.A(new_n7102), .B(new_n7034), .Y(new_n7103));
  nand_5 g04755(.A(new_n7065), .B(new_n7063), .Y(new_n7104));
  xor_4  g04756(.A(new_n7104), .B(new_n7074), .Y(new_n7105));
  not_8  g04757(.A(new_n7105), .Y(new_n7106));
  nand_5 g04758(.A(new_n7106), .B(new_n7103), .Y(new_n7107));
  not_8  g04759(.A(new_n7103), .Y(new_n7108));
  nand_5 g04760(.A(new_n7105), .B(new_n7108), .Y(new_n7109));
  nand_5 g04761(.A(new_n7007), .B(new_n7005), .Y(new_n7110));
  xor_4  g04762(.A(new_n7110), .B(new_n7032_1), .Y(new_n7111));
  nand_5 g04763(.A(new_n7070), .B(new_n7069), .Y(new_n7112));
  xor_4  g04764(.A(new_n7112), .B(new_n7072), .Y(new_n7113));
  not_8  g04765(.A(new_n7113), .Y(new_n7114));
  nand_5 g04766(.A(new_n7114), .B(new_n7111), .Y(new_n7115));
  not_8  g04767(.A(new_n7111), .Y(new_n7116));
  nand_5 g04768(.A(new_n7113), .B(new_n7116), .Y(new_n7117));
  not_8  g04769(.A(n23586), .Y(new_n7118));
  nor_5  g04770(.A(new_n7030), .B(new_n7029), .Y(new_n7119));
  xor_4  g04771(.A(new_n7119), .B(new_n7118), .Y(new_n7120));
  nand_5 g04772(.A(new_n7120), .B(new_n4521), .Y(new_n7121));
  or_5   g04773(.A(new_n7120), .B(new_n4521), .Y(new_n7122));
  nand_5 g04774(.A(new_n7011), .B(new_n7010), .Y(new_n7123));
  xor_4  g04775(.A(new_n7123), .B(new_n7025), .Y(new_n7124));
  not_8  g04776(.A(new_n7124), .Y(new_n7125));
  nand_5 g04777(.A(new_n7014), .B(new_n7013), .Y(new_n7126));
  xor_4  g04778(.A(new_n7126), .B(new_n7023), .Y(new_n7127));
  not_8  g04779(.A(new_n7127), .Y(new_n7128));
  nand_5 g04780(.A(new_n7128), .B(new_n4406), .Y(new_n7129));
  nand_5 g04781(.A(new_n7127), .B(new_n4405), .Y(new_n7130));
  nand_5 g04782(.A(new_n7016), .B(new_n7015), .Y(new_n7131));
  xor_4  g04783(.A(new_n7131), .B(new_n7021), .Y(new_n7132));
  or_5   g04784(.A(new_n7132), .B(new_n4415), .Y(new_n7133));
  nand_5 g04785(.A(new_n7132), .B(new_n4415), .Y(new_n7134));
  nand_5 g04786(.A(new_n7018), .B(new_n7017), .Y(new_n7135));
  not_8  g04787(.A(new_n7135), .Y(new_n7136));
  xor_4  g04788(.A(new_n7136), .B(new_n7019), .Y(new_n7137));
  not_8  g04789(.A(new_n7137), .Y(new_n7138));
  or_5   g04790(.A(new_n7138), .B(new_n4421), .Y(new_n7139_1));
  nand_5 g04791(.A(new_n7138), .B(new_n4421), .Y(new_n7140));
  nand_5 g04792(.A(new_n2636), .B(new_n4545), .Y(new_n7141));
  and_5  g04793(.A(new_n7141), .B(new_n7019), .Y(new_n7142));
  nand_5 g04794(.A(new_n7142), .B(new_n4426_1), .Y(new_n7143));
  nand_5 g04795(.A(new_n7143), .B(new_n7140), .Y(new_n7144));
  nand_5 g04796(.A(new_n7144), .B(new_n7139_1), .Y(new_n7145));
  nand_5 g04797(.A(new_n7145), .B(new_n7134), .Y(new_n7146));
  nand_5 g04798(.A(new_n7146), .B(new_n7133), .Y(new_n7147));
  nand_5 g04799(.A(new_n7147), .B(new_n7130), .Y(new_n7148));
  nand_5 g04800(.A(new_n7148), .B(new_n7129), .Y(new_n7149_1));
  or_5   g04801(.A(new_n7149_1), .B(new_n7125), .Y(new_n7150));
  nand_5 g04802(.A(new_n7149_1), .B(new_n7125), .Y(new_n7151));
  nand_5 g04803(.A(new_n7151), .B(new_n4447), .Y(new_n7152));
  nand_5 g04804(.A(new_n7152), .B(new_n7150), .Y(new_n7153));
  not_8  g04805(.A(new_n7153), .Y(new_n7154));
  nand_5 g04806(.A(new_n7154), .B(new_n7122), .Y(new_n7155));
  nand_5 g04807(.A(new_n7155), .B(new_n7121), .Y(new_n7156));
  nand_5 g04808(.A(new_n7156), .B(new_n7117), .Y(new_n7157));
  nand_5 g04809(.A(new_n7157), .B(new_n7115), .Y(new_n7158));
  nand_5 g04810(.A(new_n7158), .B(new_n7109), .Y(new_n7159));
  nand_5 g04811(.A(new_n7159), .B(new_n7107), .Y(new_n7160));
  nand_5 g04812(.A(new_n7160), .B(new_n7101), .Y(new_n7161));
  nand_5 g04813(.A(new_n7161), .B(new_n7099_1), .Y(new_n7162));
  nand_5 g04814(.A(new_n7162), .B(new_n7093), .Y(new_n7163));
  nand_5 g04815(.A(new_n7163), .B(new_n7091), .Y(new_n7164));
  xor_4  g04816(.A(new_n7164), .B(new_n7085), .Y(new_n7165));
  not_8  g04817(.A(n6105), .Y(new_n7166));
  not_8  g04818(.A(n15766), .Y(new_n7167));
  nand_5 g04819(.A(new_n7167), .B(new_n7166), .Y(new_n7168));
  nand_5 g04820(.A(n15766), .B(n6105), .Y(new_n7169));
  not_8  g04821(.A(n3795), .Y(new_n7170));
  not_8  g04822(.A(n25629), .Y(new_n7171));
  nand_5 g04823(.A(new_n7171), .B(new_n7170), .Y(new_n7172));
  nand_5 g04824(.A(n25629), .B(n3795), .Y(new_n7173));
  not_8  g04825(.A(n7692), .Y(new_n7174));
  not_8  g04826(.A(n25464), .Y(new_n7175));
  nand_5 g04827(.A(new_n7175), .B(new_n7174), .Y(new_n7176));
  nand_5 g04828(.A(n25464), .B(n7692), .Y(new_n7177));
  not_8  g04829(.A(n4590), .Y(new_n7178));
  not_8  g04830(.A(n23039), .Y(new_n7179));
  nand_5 g04831(.A(new_n7179), .B(new_n7178), .Y(new_n7180));
  nand_5 g04832(.A(n23039), .B(n4590), .Y(new_n7181));
  not_8  g04833(.A(n26752), .Y(new_n7182));
  nand_5 g04834(.A(new_n7182), .B(new_n4489), .Y(new_n7183));
  nand_5 g04835(.A(n26752), .B(n13677), .Y(new_n7184));
  not_8  g04836(.A(n6513), .Y(new_n7185));
  nand_5 g04837(.A(new_n4359), .B(new_n7185), .Y(new_n7186));
  nand_5 g04838(.A(n18926), .B(n6513), .Y(new_n7187));
  not_8  g04839(.A(n3918), .Y(new_n7188));
  nand_5 g04840(.A(new_n4315), .B(new_n7188), .Y(new_n7189));
  nand_5 g04841(.A(n5451), .B(n3918), .Y(new_n7190_1));
  nand_5 g04842(.A(new_n4588_1), .B(new_n4585), .Y(new_n7191));
  nand_5 g04843(.A(new_n7191), .B(new_n4587), .Y(new_n7192));
  nand_5 g04844(.A(new_n7192), .B(new_n7190_1), .Y(new_n7193));
  nand_5 g04845(.A(new_n7193), .B(new_n7189), .Y(new_n7194));
  nand_5 g04846(.A(new_n7194), .B(new_n7187), .Y(new_n7195));
  nand_5 g04847(.A(new_n7195), .B(new_n7186), .Y(new_n7196));
  nand_5 g04848(.A(new_n7196), .B(new_n7184), .Y(new_n7197));
  nand_5 g04849(.A(new_n7197), .B(new_n7183), .Y(new_n7198));
  nand_5 g04850(.A(new_n7198), .B(new_n7181), .Y(new_n7199));
  nand_5 g04851(.A(new_n7199), .B(new_n7180), .Y(new_n7200));
  nand_5 g04852(.A(new_n7200), .B(new_n7177), .Y(new_n7201));
  nand_5 g04853(.A(new_n7201), .B(new_n7176), .Y(new_n7202));
  nand_5 g04854(.A(new_n7202), .B(new_n7173), .Y(new_n7203));
  nand_5 g04855(.A(new_n7203), .B(new_n7172), .Y(new_n7204));
  nand_5 g04856(.A(new_n7204), .B(new_n7169), .Y(new_n7205));
  nand_5 g04857(.A(new_n7205), .B(new_n7168), .Y(new_n7206));
  or_5   g04858(.A(new_n7206), .B(new_n7165), .Y(new_n7207));
  nand_5 g04859(.A(new_n7206), .B(new_n7165), .Y(new_n7208));
  nand_5 g04860(.A(new_n7169), .B(new_n7168), .Y(new_n7209));
  xor_4  g04861(.A(new_n7209), .B(new_n7204), .Y(new_n7210));
  not_8  g04862(.A(new_n7210), .Y(new_n7211));
  nand_5 g04863(.A(new_n7091), .B(new_n7093), .Y(new_n7212));
  xor_4  g04864(.A(new_n7212), .B(new_n7162), .Y(new_n7213));
  or_5   g04865(.A(new_n7213), .B(new_n7211), .Y(new_n7214));
  nand_5 g04866(.A(new_n7213), .B(new_n7211), .Y(new_n7215));
  nand_5 g04867(.A(new_n7173), .B(new_n7172), .Y(new_n7216));
  xor_4  g04868(.A(new_n7216), .B(new_n7202), .Y(new_n7217));
  not_8  g04869(.A(new_n7217), .Y(new_n7218));
  nand_5 g04870(.A(new_n7099_1), .B(new_n7101), .Y(new_n7219));
  xor_4  g04871(.A(new_n7219), .B(new_n7160), .Y(new_n7220));
  or_5   g04872(.A(new_n7220), .B(new_n7218), .Y(new_n7221));
  not_8  g04873(.A(new_n7221), .Y(new_n7222));
  nand_5 g04874(.A(new_n7220), .B(new_n7218), .Y(new_n7223));
  not_8  g04875(.A(new_n7223), .Y(new_n7224));
  nand_5 g04876(.A(new_n7177), .B(new_n7176), .Y(new_n7225));
  xor_4  g04877(.A(new_n7225), .B(new_n7200), .Y(new_n7226));
  not_8  g04878(.A(new_n7226), .Y(new_n7227));
  nand_5 g04879(.A(new_n7107), .B(new_n7109), .Y(new_n7228));
  xor_4  g04880(.A(new_n7228), .B(new_n7158), .Y(new_n7229_1));
  or_5   g04881(.A(new_n7229_1), .B(new_n7227), .Y(new_n7230_1));
  not_8  g04882(.A(new_n7230_1), .Y(new_n7231));
  nand_5 g04883(.A(new_n7229_1), .B(new_n7227), .Y(new_n7232));
  not_8  g04884(.A(new_n7232), .Y(new_n7233_1));
  nand_5 g04885(.A(new_n7181), .B(new_n7180), .Y(new_n7234));
  xor_4  g04886(.A(new_n7234), .B(new_n7198), .Y(new_n7235));
  not_8  g04887(.A(new_n7235), .Y(new_n7236_1));
  nand_5 g04888(.A(new_n7115), .B(new_n7117), .Y(new_n7237));
  xor_4  g04889(.A(new_n7237), .B(new_n7156), .Y(new_n7238));
  nand_5 g04890(.A(new_n7238), .B(new_n7236_1), .Y(new_n7239));
  or_5   g04891(.A(new_n7238), .B(new_n7236_1), .Y(new_n7240));
  nand_5 g04892(.A(new_n7184), .B(new_n7183), .Y(new_n7241));
  xor_4  g04893(.A(new_n7241), .B(new_n7196), .Y(new_n7242));
  not_8  g04894(.A(new_n7242), .Y(new_n7243));
  nand_5 g04895(.A(new_n7121), .B(new_n7122), .Y(new_n7244));
  xor_4  g04896(.A(new_n7244), .B(new_n7154), .Y(new_n7245));
  nand_5 g04897(.A(new_n7245), .B(new_n7243), .Y(new_n7246));
  nor_5  g04898(.A(new_n7245), .B(new_n7243), .Y(new_n7247));
  not_8  g04899(.A(new_n7247), .Y(new_n7248));
  nand_5 g04900(.A(new_n7187), .B(new_n7186), .Y(new_n7249));
  xor_4  g04901(.A(new_n7249), .B(new_n7194), .Y(new_n7250));
  not_8  g04902(.A(new_n7250), .Y(new_n7251));
  nand_5 g04903(.A(new_n7151), .B(new_n7150), .Y(new_n7252));
  xor_4  g04904(.A(new_n7252), .B(new_n4448), .Y(new_n7253_1));
  nand_5 g04905(.A(new_n7253_1), .B(new_n7251), .Y(new_n7254));
  nor_5  g04906(.A(new_n7253_1), .B(new_n7251), .Y(new_n7255));
  not_8  g04907(.A(new_n7255), .Y(new_n7256_1));
  nand_5 g04908(.A(new_n7190_1), .B(new_n7189), .Y(new_n7257));
  xor_4  g04909(.A(new_n7257), .B(new_n7192), .Y(new_n7258));
  not_8  g04910(.A(new_n7258), .Y(new_n7259));
  nand_5 g04911(.A(new_n7129), .B(new_n7130), .Y(new_n7260));
  xor_4  g04912(.A(new_n7260), .B(new_n7147), .Y(new_n7261));
  nand_5 g04913(.A(new_n7261), .B(new_n7259), .Y(new_n7262));
  nor_5  g04914(.A(new_n7261), .B(new_n7259), .Y(new_n7263));
  not_8  g04915(.A(new_n7263), .Y(new_n7264));
  nand_5 g04916(.A(new_n7133), .B(new_n7134), .Y(new_n7265));
  xor_4  g04917(.A(new_n7265), .B(new_n7145), .Y(new_n7266));
  nand_5 g04918(.A(new_n7266), .B(new_n4590_1), .Y(new_n7267));
  nor_5  g04919(.A(new_n7266), .B(new_n4590_1), .Y(new_n7268_1));
  not_8  g04920(.A(new_n7268_1), .Y(new_n7269));
  nand_5 g04921(.A(new_n7139_1), .B(new_n7140), .Y(new_n7270));
  xor_4  g04922(.A(new_n7270), .B(new_n7143), .Y(new_n7271));
  nand_5 g04923(.A(new_n7271), .B(new_n4539), .Y(new_n7272));
  nor_5  g04924(.A(new_n7271), .B(new_n4539), .Y(new_n7273));
  not_8  g04925(.A(new_n7273), .Y(new_n7274));
  not_8  g04926(.A(new_n7142), .Y(new_n7275));
  nand_5 g04927(.A(new_n7275), .B(new_n2640), .Y(new_n7276));
  and_5  g04928(.A(new_n7276), .B(new_n7143), .Y(new_n7277_1));
  or_5   g04929(.A(new_n7277_1), .B(new_n4577), .Y(new_n7278));
  nand_5 g04930(.A(new_n7278), .B(new_n7274), .Y(new_n7279));
  nand_5 g04931(.A(new_n7279), .B(new_n7272), .Y(new_n7280_1));
  nand_5 g04932(.A(new_n7280_1), .B(new_n7269), .Y(new_n7281));
  nand_5 g04933(.A(new_n7281), .B(new_n7267), .Y(new_n7282));
  nand_5 g04934(.A(new_n7282), .B(new_n7264), .Y(new_n7283));
  nand_5 g04935(.A(new_n7283), .B(new_n7262), .Y(new_n7284));
  nand_5 g04936(.A(new_n7284), .B(new_n7256_1), .Y(new_n7285));
  nand_5 g04937(.A(new_n7285), .B(new_n7254), .Y(new_n7286));
  nand_5 g04938(.A(new_n7286), .B(new_n7248), .Y(new_n7287));
  nand_5 g04939(.A(new_n7287), .B(new_n7246), .Y(new_n7288));
  nand_5 g04940(.A(new_n7288), .B(new_n7240), .Y(new_n7289));
  nand_5 g04941(.A(new_n7289), .B(new_n7239), .Y(new_n7290));
  nor_5  g04942(.A(new_n7290), .B(new_n7233_1), .Y(new_n7291));
  nor_5  g04943(.A(new_n7291), .B(new_n7231), .Y(new_n7292));
  nor_5  g04944(.A(new_n7292), .B(new_n7224), .Y(new_n7293));
  nor_5  g04945(.A(new_n7293), .B(new_n7222), .Y(new_n7294));
  not_8  g04946(.A(new_n7294), .Y(new_n7295));
  nand_5 g04947(.A(new_n7295), .B(new_n7215), .Y(new_n7296));
  nand_5 g04948(.A(new_n7296), .B(new_n7214), .Y(new_n7297));
  nand_5 g04949(.A(new_n7297), .B(new_n7208), .Y(new_n7298_1));
  nand_5 g04950(.A(new_n7298_1), .B(new_n7207), .Y(new_n7299));
  nand_5 g04951(.A(new_n7164), .B(new_n7084), .Y(new_n7300));
  nand_5 g04952(.A(new_n7300), .B(new_n7083), .Y(new_n7301));
  and_5  g04953(.A(new_n7301), .B(new_n7299), .Y(n588));
  not_8  g04954(.A(n12113), .Y(new_n7303));
  or_5   g04955(.A(n12917), .B(new_n7303), .Y(new_n7304));
  nand_5 g04956(.A(n12917), .B(new_n7303), .Y(new_n7305_1));
  not_8  g04957(.A(n10614), .Y(new_n7306));
  or_5   g04958(.A(n21898), .B(new_n7306), .Y(new_n7307));
  nand_5 g04959(.A(n21898), .B(new_n7306), .Y(new_n7308_1));
  not_8  g04960(.A(n9926), .Y(new_n7309));
  nand_5 g04961(.A(n11266), .B(new_n7309), .Y(new_n7310));
  not_8  g04962(.A(new_n7310), .Y(new_n7311));
  nor_5  g04963(.A(n11266), .B(new_n7309), .Y(new_n7312));
  not_8  g04964(.A(n2646), .Y(new_n7313_1));
  nand_5 g04965(.A(n22072), .B(new_n7313_1), .Y(new_n7314));
  not_8  g04966(.A(new_n7314), .Y(new_n7315));
  nor_5  g04967(.A(new_n7315), .B(new_n7312), .Y(new_n7316));
  nor_5  g04968(.A(new_n7316), .B(new_n7311), .Y(new_n7317));
  not_8  g04969(.A(new_n7317), .Y(new_n7318));
  nand_5 g04970(.A(new_n7318), .B(new_n7308_1), .Y(new_n7319));
  nand_5 g04971(.A(new_n7319), .B(new_n7307), .Y(new_n7320));
  nand_5 g04972(.A(new_n7320), .B(new_n7305_1), .Y(new_n7321));
  nand_5 g04973(.A(new_n7321), .B(new_n7304), .Y(new_n7322));
  not_8  g04974(.A(n5517), .Y(new_n7323));
  or_5   g04975(.A(n21981), .B(new_n7323), .Y(new_n7324));
  nand_5 g04976(.A(n21981), .B(new_n7323), .Y(new_n7325));
  nand_5 g04977(.A(new_n7325), .B(new_n7324), .Y(new_n7326));
  xor_4  g04978(.A(new_n7326), .B(new_n7322), .Y(new_n7327));
  not_8  g04979(.A(new_n7327), .Y(new_n7328));
  not_8  g04980(.A(n9493), .Y(new_n7329));
  not_8  g04981(.A(n4939), .Y(new_n7330_1));
  not_8  g04982(.A(n15652), .Y(new_n7331));
  nand_5 g04983(.A(new_n7331), .B(new_n7330_1), .Y(new_n7332));
  or_5   g04984(.A(new_n7332), .B(n5605), .Y(new_n7333));
  nor_5  g04985(.A(new_n7333), .B(n2985), .Y(new_n7334));
  not_8  g04986(.A(new_n7334), .Y(new_n7335_1));
  nand_5 g04987(.A(new_n7333), .B(n2985), .Y(new_n7336));
  and_5  g04988(.A(new_n7336), .B(new_n7335_1), .Y(new_n7337));
  not_8  g04989(.A(new_n7337), .Y(new_n7338));
  nand_5 g04990(.A(new_n7338), .B(new_n7329), .Y(new_n7339_1));
  nand_5 g04991(.A(new_n7337), .B(n9493), .Y(new_n7340));
  not_8  g04992(.A(n15167), .Y(new_n7341));
  nand_5 g04993(.A(new_n7332), .B(n5605), .Y(new_n7342));
  and_5  g04994(.A(new_n7342), .B(new_n7333), .Y(new_n7343));
  not_8  g04995(.A(new_n7343), .Y(new_n7344));
  nand_5 g04996(.A(new_n7344), .B(new_n7341), .Y(new_n7345));
  nand_5 g04997(.A(new_n7343), .B(n15167), .Y(new_n7346_1));
  not_8  g04998(.A(n21095), .Y(new_n7347));
  nand_5 g04999(.A(n15652), .B(n4939), .Y(new_n7348));
  and_5  g05000(.A(new_n7348), .B(new_n7332), .Y(new_n7349_1));
  not_8  g05001(.A(new_n7349_1), .Y(new_n7350));
  nand_5 g05002(.A(new_n7350), .B(new_n7347), .Y(new_n7351));
  nand_5 g05003(.A(new_n7349_1), .B(n21095), .Y(new_n7352));
  nand_5 g05004(.A(n8656), .B(n4939), .Y(new_n7353));
  nand_5 g05005(.A(new_n7353), .B(new_n7352), .Y(new_n7354));
  nand_5 g05006(.A(new_n7354), .B(new_n7351), .Y(new_n7355));
  nand_5 g05007(.A(new_n7355), .B(new_n7346_1), .Y(new_n7356));
  nand_5 g05008(.A(new_n7356), .B(new_n7345), .Y(new_n7357));
  nand_5 g05009(.A(new_n7357), .B(new_n7340), .Y(new_n7358));
  nand_5 g05010(.A(new_n7358), .B(new_n7339_1), .Y(new_n7359));
  not_8  g05011(.A(n8244), .Y(new_n7360));
  not_8  g05012(.A(n14576), .Y(new_n7361));
  nand_5 g05013(.A(new_n7334), .B(new_n7361), .Y(new_n7362));
  nand_5 g05014(.A(new_n7335_1), .B(n14576), .Y(new_n7363_1));
  and_5  g05015(.A(new_n7363_1), .B(new_n7362), .Y(new_n7364));
  not_8  g05016(.A(new_n7364), .Y(new_n7365));
  nand_5 g05017(.A(new_n7365), .B(new_n7360), .Y(new_n7366));
  nand_5 g05018(.A(new_n7364), .B(n8244), .Y(new_n7367));
  nand_5 g05019(.A(new_n7367), .B(new_n7366), .Y(new_n7368));
  xor_4  g05020(.A(new_n7368), .B(new_n7359), .Y(new_n7369));
  nand_5 g05021(.A(new_n7369), .B(new_n7328), .Y(new_n7370));
  nor_5  g05022(.A(new_n7369), .B(new_n7328), .Y(new_n7371));
  not_8  g05023(.A(new_n7371), .Y(new_n7372));
  nand_5 g05024(.A(new_n7305_1), .B(new_n7304), .Y(new_n7373));
  xor_4  g05025(.A(new_n7373), .B(new_n7320), .Y(new_n7374));
  not_8  g05026(.A(new_n7374), .Y(new_n7375));
  nand_5 g05027(.A(new_n7340), .B(new_n7339_1), .Y(new_n7376));
  xor_4  g05028(.A(new_n7376), .B(new_n7357), .Y(new_n7377_1));
  nand_5 g05029(.A(new_n7377_1), .B(new_n7375), .Y(new_n7378));
  or_5   g05030(.A(new_n7377_1), .B(new_n7375), .Y(new_n7379));
  nand_5 g05031(.A(new_n7308_1), .B(new_n7307), .Y(new_n7380));
  xor_4  g05032(.A(new_n7380), .B(new_n7317), .Y(new_n7381));
  nand_5 g05033(.A(new_n7346_1), .B(new_n7345), .Y(new_n7382));
  xor_4  g05034(.A(new_n7382), .B(new_n7355), .Y(new_n7383));
  or_5   g05035(.A(new_n7383), .B(new_n7381), .Y(new_n7384));
  nand_5 g05036(.A(new_n7383), .B(new_n7381), .Y(new_n7385));
  nor_5  g05037(.A(new_n7312), .B(new_n7311), .Y(new_n7386));
  xor_4  g05038(.A(new_n7386), .B(new_n7315), .Y(new_n7387));
  nor_5  g05039(.A(n22072), .B(new_n7313_1), .Y(new_n7388));
  nor_5  g05040(.A(new_n7388), .B(new_n7315), .Y(new_n7389));
  not_8  g05041(.A(new_n7389), .Y(new_n7390_1));
  xor_4  g05042(.A(n8656), .B(n4939), .Y(new_n7391));
  nand_5 g05043(.A(new_n7391), .B(new_n7390_1), .Y(new_n7392));
  nand_5 g05044(.A(new_n7392), .B(new_n7387), .Y(new_n7393));
  or_5   g05045(.A(new_n7392), .B(new_n7387), .Y(new_n7394));
  nand_5 g05046(.A(new_n7352), .B(new_n7351), .Y(new_n7395));
  xnor_4 g05047(.A(new_n7395), .B(new_n7353), .Y(new_n7396));
  nand_5 g05048(.A(new_n7396), .B(new_n7394), .Y(new_n7397));
  nand_5 g05049(.A(new_n7397), .B(new_n7393), .Y(new_n7398));
  nand_5 g05050(.A(new_n7398), .B(new_n7385), .Y(new_n7399));
  nand_5 g05051(.A(new_n7399), .B(new_n7384), .Y(new_n7400));
  not_8  g05052(.A(new_n7400), .Y(new_n7401));
  nand_5 g05053(.A(new_n7401), .B(new_n7379), .Y(new_n7402));
  nand_5 g05054(.A(new_n7402), .B(new_n7378), .Y(new_n7403_1));
  nand_5 g05055(.A(new_n7403_1), .B(new_n7372), .Y(new_n7404));
  nand_5 g05056(.A(new_n7404), .B(new_n7370), .Y(new_n7405));
  nand_5 g05057(.A(new_n7325), .B(new_n7322), .Y(new_n7406));
  nand_5 g05058(.A(new_n7406), .B(new_n7324), .Y(new_n7407));
  not_8  g05059(.A(n376), .Y(new_n7408_1));
  or_5   g05060(.A(n7721), .B(new_n7408_1), .Y(new_n7409));
  nand_5 g05061(.A(n7721), .B(new_n7408_1), .Y(new_n7410));
  nand_5 g05062(.A(new_n7410), .B(new_n7409), .Y(new_n7411));
  xor_4  g05063(.A(new_n7411), .B(new_n7407), .Y(new_n7412));
  not_8  g05064(.A(new_n7412), .Y(new_n7413));
  nand_5 g05065(.A(new_n7367), .B(new_n7359), .Y(new_n7414));
  nand_5 g05066(.A(new_n7414), .B(new_n7366), .Y(new_n7415));
  not_8  g05067(.A(n4858), .Y(new_n7416));
  nor_5  g05068(.A(new_n7362), .B(n1269), .Y(new_n7417));
  not_8  g05069(.A(new_n7417), .Y(new_n7418));
  nand_5 g05070(.A(new_n7362), .B(n1269), .Y(new_n7419));
  and_5  g05071(.A(new_n7419), .B(new_n7418), .Y(new_n7420));
  not_8  g05072(.A(new_n7420), .Y(new_n7421_1));
  nand_5 g05073(.A(new_n7421_1), .B(new_n7416), .Y(new_n7422));
  nand_5 g05074(.A(new_n7420), .B(n4858), .Y(new_n7423));
  nand_5 g05075(.A(new_n7423), .B(new_n7422), .Y(new_n7424));
  xor_4  g05076(.A(new_n7424), .B(new_n7415), .Y(new_n7425));
  nand_5 g05077(.A(new_n7425), .B(new_n7413), .Y(new_n7426));
  nor_5  g05078(.A(new_n7425), .B(new_n7413), .Y(new_n7427));
  not_8  g05079(.A(new_n7427), .Y(new_n7428_1));
  nand_5 g05080(.A(new_n7428_1), .B(new_n7426), .Y(new_n7429));
  xor_4  g05081(.A(new_n7429), .B(new_n7405), .Y(new_n7430));
  nand_5 g05082(.A(new_n7430), .B(new_n5308), .Y(new_n7431));
  not_8  g05083(.A(new_n7430), .Y(new_n7432_1));
  nand_5 g05084(.A(new_n7432_1), .B(new_n5307), .Y(new_n7433));
  nand_5 g05085(.A(new_n7372), .B(new_n7370), .Y(new_n7434));
  xor_4  g05086(.A(new_n7434), .B(new_n7403_1), .Y(new_n7435));
  nand_5 g05087(.A(new_n7435), .B(new_n5216), .Y(new_n7436));
  not_8  g05088(.A(new_n7435), .Y(new_n7437_1));
  nand_5 g05089(.A(new_n7437_1), .B(new_n5219), .Y(new_n7438));
  nand_5 g05090(.A(new_n7378), .B(new_n7379), .Y(new_n7439));
  xor_4  g05091(.A(new_n7439), .B(new_n7401), .Y(new_n7440));
  nand_5 g05092(.A(new_n7440), .B(new_n5171), .Y(new_n7441));
  not_8  g05093(.A(new_n7440), .Y(new_n7442));
  nand_5 g05094(.A(new_n7442), .B(new_n5174), .Y(new_n7443));
  nand_5 g05095(.A(new_n7384), .B(new_n7385), .Y(new_n7444));
  xor_4  g05096(.A(new_n7444), .B(new_n7398), .Y(new_n7445));
  not_8  g05097(.A(new_n7445), .Y(new_n7446));
  nand_5 g05098(.A(new_n7446), .B(new_n5179), .Y(new_n7447));
  or_5   g05099(.A(new_n7446), .B(new_n5179), .Y(new_n7448));
  xor_4  g05100(.A(new_n7391), .B(new_n7389), .Y(new_n7449));
  or_5   g05101(.A(new_n7449), .B(new_n5193), .Y(new_n7450));
  nand_5 g05102(.A(new_n7450), .B(new_n5187), .Y(new_n7451));
  or_5   g05103(.A(new_n7450), .B(new_n5187), .Y(new_n7452));
  nand_5 g05104(.A(new_n7393), .B(new_n7394), .Y(new_n7453));
  xor_4  g05105(.A(new_n7453), .B(new_n7396), .Y(new_n7454));
  not_8  g05106(.A(new_n7454), .Y(new_n7455));
  nand_5 g05107(.A(new_n7455), .B(new_n7452), .Y(new_n7456));
  nand_5 g05108(.A(new_n7456), .B(new_n7451), .Y(new_n7457));
  nand_5 g05109(.A(new_n7457), .B(new_n7448), .Y(new_n7458));
  nand_5 g05110(.A(new_n7458), .B(new_n7447), .Y(new_n7459));
  nand_5 g05111(.A(new_n7459), .B(new_n7443), .Y(new_n7460_1));
  nand_5 g05112(.A(new_n7460_1), .B(new_n7441), .Y(new_n7461));
  nand_5 g05113(.A(new_n7461), .B(new_n7438), .Y(new_n7462));
  nand_5 g05114(.A(new_n7462), .B(new_n7436), .Y(new_n7463));
  nand_5 g05115(.A(new_n7463), .B(new_n7433), .Y(new_n7464));
  nand_5 g05116(.A(new_n7464), .B(new_n7431), .Y(new_n7465));
  nand_5 g05117(.A(new_n5305), .B(new_n5300_1), .Y(new_n7466));
  nand_5 g05118(.A(new_n7466), .B(new_n5303), .Y(new_n7467));
  not_8  g05119(.A(new_n7467), .Y(new_n7468));
  not_8  g05120(.A(n18584), .Y(new_n7469));
  or_5   g05121(.A(n19803), .B(new_n7469), .Y(new_n7470));
  nand_5 g05122(.A(n19803), .B(new_n7469), .Y(new_n7471));
  nand_5 g05123(.A(new_n7471), .B(new_n7470), .Y(new_n7472));
  xor_4  g05124(.A(new_n7472), .B(new_n7468), .Y(new_n7473));
  not_8  g05125(.A(new_n7473), .Y(new_n7474));
  nand_5 g05126(.A(new_n7428_1), .B(new_n7405), .Y(new_n7475_1));
  nand_5 g05127(.A(new_n7475_1), .B(new_n7426), .Y(new_n7476));
  not_8  g05128(.A(new_n7476), .Y(new_n7477_1));
  nand_5 g05129(.A(new_n7410), .B(new_n7407), .Y(new_n7478));
  nand_5 g05130(.A(new_n7478), .B(new_n7409), .Y(new_n7479));
  not_8  g05131(.A(new_n7479), .Y(new_n7480));
  not_8  g05132(.A(n7773), .Y(new_n7481));
  nand_5 g05133(.A(n16911), .B(new_n7481), .Y(new_n7482));
  nor_5  g05134(.A(n16911), .B(new_n7481), .Y(new_n7483));
  not_8  g05135(.A(new_n7483), .Y(new_n7484));
  nand_5 g05136(.A(new_n7484), .B(new_n7482), .Y(new_n7485));
  xor_4  g05137(.A(new_n7485), .B(new_n7480), .Y(new_n7486));
  not_8  g05138(.A(new_n7486), .Y(new_n7487));
  nand_5 g05139(.A(new_n7423), .B(new_n7415), .Y(new_n7488));
  nand_5 g05140(.A(new_n7488), .B(new_n7422), .Y(new_n7489));
  not_8  g05141(.A(new_n7489), .Y(new_n7490));
  not_8  g05142(.A(n1742), .Y(new_n7491));
  not_8  g05143(.A(n16818), .Y(new_n7492));
  nand_5 g05144(.A(new_n7417), .B(new_n7492), .Y(new_n7493));
  nand_5 g05145(.A(new_n7418), .B(n16818), .Y(new_n7494));
  and_5  g05146(.A(new_n7494), .B(new_n7493), .Y(new_n7495));
  not_8  g05147(.A(new_n7495), .Y(new_n7496));
  nand_5 g05148(.A(new_n7496), .B(new_n7491), .Y(new_n7497));
  nand_5 g05149(.A(new_n7495), .B(n1742), .Y(new_n7498));
  nand_5 g05150(.A(new_n7498), .B(new_n7497), .Y(new_n7499));
  xor_4  g05151(.A(new_n7499), .B(new_n7490), .Y(new_n7500));
  or_5   g05152(.A(new_n7500), .B(new_n7487), .Y(new_n7501));
  nand_5 g05153(.A(new_n7500), .B(new_n7487), .Y(new_n7502));
  nand_5 g05154(.A(new_n7502), .B(new_n7501), .Y(new_n7503));
  xor_4  g05155(.A(new_n7503), .B(new_n7477_1), .Y(new_n7504));
  not_8  g05156(.A(new_n7504), .Y(new_n7505));
  nand_5 g05157(.A(new_n7505), .B(new_n7474), .Y(new_n7506));
  nand_5 g05158(.A(new_n7504), .B(new_n7473), .Y(new_n7507_1));
  nand_5 g05159(.A(new_n7507_1), .B(new_n7506), .Y(new_n7508));
  xor_4  g05160(.A(new_n7508), .B(new_n7465), .Y(n597));
  xor_4  g05161(.A(n25926), .B(n9646), .Y(new_n7510));
  not_8  g05162(.A(new_n7510), .Y(new_n7511));
  nand_5 g05163(.A(new_n7511), .B(n14230), .Y(new_n7512));
  not_8  g05164(.A(n14230), .Y(new_n7513));
  nand_5 g05165(.A(new_n7510), .B(new_n7513), .Y(new_n7514_1));
  nand_5 g05166(.A(new_n7514_1), .B(new_n7512), .Y(new_n7515));
  xor_4  g05167(.A(new_n7515), .B(new_n6576_1), .Y(n637));
  nand_5 g05168(.A(n24323), .B(n8581), .Y(new_n7517));
  not_8  g05169(.A(new_n7517), .Y(new_n7518));
  not_8  g05170(.A(n5026), .Y(new_n7519));
  nand_5 g05171(.A(new_n6544), .B(new_n7519), .Y(new_n7520));
  nand_5 g05172(.A(n25877), .B(n5026), .Y(new_n7521));
  nand_5 g05173(.A(new_n7521), .B(new_n7520), .Y(new_n7522));
  xor_4  g05174(.A(new_n7522), .B(new_n7518), .Y(new_n7523));
  or_5   g05175(.A(new_n7523), .B(new_n4898), .Y(new_n7524_1));
  nand_5 g05176(.A(new_n7523), .B(new_n4898), .Y(new_n7525));
  not_8  g05177(.A(n8581), .Y(new_n7526));
  nand_5 g05178(.A(new_n6537), .B(new_n7526), .Y(new_n7527));
  and_5  g05179(.A(new_n7527), .B(new_n7517), .Y(new_n7528));
  nand_5 g05180(.A(new_n7528), .B(n1681), .Y(new_n7529));
  not_8  g05181(.A(new_n7529), .Y(new_n7530));
  nand_5 g05182(.A(new_n7530), .B(new_n7525), .Y(new_n7531));
  nand_5 g05183(.A(new_n7531), .B(new_n7524_1), .Y(new_n7532));
  not_8  g05184(.A(new_n7532), .Y(new_n7533));
  nand_5 g05185(.A(new_n7521), .B(new_n7517), .Y(new_n7534));
  nand_5 g05186(.A(new_n7534), .B(new_n7520), .Y(new_n7535));
  not_8  g05187(.A(new_n7535), .Y(new_n7536));
  nand_5 g05188(.A(n15271), .B(n12161), .Y(new_n7537));
  not_8  g05189(.A(n12161), .Y(new_n7538));
  not_8  g05190(.A(n15271), .Y(new_n7539));
  nand_5 g05191(.A(new_n7539), .B(new_n7538), .Y(new_n7540));
  nand_5 g05192(.A(new_n7540), .B(new_n7537), .Y(new_n7541));
  xor_4  g05193(.A(new_n7541), .B(new_n7536), .Y(new_n7542));
  or_5   g05194(.A(new_n7542), .B(new_n4892), .Y(new_n7543));
  nand_5 g05195(.A(new_n7542), .B(new_n4892), .Y(new_n7544));
  nand_5 g05196(.A(new_n7544), .B(new_n7543), .Y(new_n7545));
  xor_4  g05197(.A(new_n7545), .B(new_n7533), .Y(new_n7546));
  not_8  g05198(.A(new_n7546), .Y(new_n7547));
  nand_5 g05199(.A(n25435), .B(n18), .Y(new_n7548));
  not_8  g05200(.A(new_n7548), .Y(new_n7549));
  not_8  g05201(.A(n15490), .Y(new_n7550));
  nand_5 g05202(.A(new_n7550), .B(new_n4148), .Y(new_n7551));
  nand_5 g05203(.A(n15490), .B(n13319), .Y(new_n7552));
  nand_5 g05204(.A(new_n7552), .B(new_n7551), .Y(new_n7553));
  xor_4  g05205(.A(new_n7553), .B(new_n7549), .Y(new_n7554));
  not_8  g05206(.A(new_n7554), .Y(new_n7555));
  nand_5 g05207(.A(new_n7555), .B(n2809), .Y(new_n7556));
  nand_5 g05208(.A(new_n7554), .B(new_n5394), .Y(new_n7557));
  not_8  g05209(.A(n18), .Y(new_n7558_1));
  nand_5 g05210(.A(new_n4149), .B(new_n7558_1), .Y(new_n7559));
  and_5  g05211(.A(new_n7559), .B(new_n7548), .Y(new_n7560));
  nand_5 g05212(.A(new_n7560), .B(n15508), .Y(new_n7561));
  not_8  g05213(.A(new_n7561), .Y(new_n7562));
  nand_5 g05214(.A(new_n7562), .B(new_n7557), .Y(new_n7563));
  nand_5 g05215(.A(new_n7563), .B(new_n7556), .Y(new_n7564));
  nand_5 g05216(.A(new_n7552), .B(new_n7548), .Y(new_n7565));
  nand_5 g05217(.A(new_n7565), .B(new_n7551), .Y(new_n7566_1));
  not_8  g05218(.A(new_n7566_1), .Y(new_n7567));
  nand_5 g05219(.A(n15967), .B(n2783), .Y(new_n7568));
  not_8  g05220(.A(n2783), .Y(new_n7569_1));
  nand_5 g05221(.A(new_n4147), .B(new_n7569_1), .Y(new_n7570));
  nand_5 g05222(.A(new_n7570), .B(new_n7568), .Y(new_n7571));
  xor_4  g05223(.A(new_n7571), .B(new_n7567), .Y(new_n7572_1));
  not_8  g05224(.A(new_n7572_1), .Y(new_n7573));
  nand_5 g05225(.A(new_n7573), .B(n19680), .Y(new_n7574));
  nand_5 g05226(.A(new_n7572_1), .B(new_n5391), .Y(new_n7575_1));
  nand_5 g05227(.A(new_n7575_1), .B(new_n7574), .Y(new_n7576));
  xor_4  g05228(.A(new_n7576), .B(new_n7564), .Y(new_n7577));
  not_8  g05229(.A(new_n7577), .Y(new_n7578));
  nand_5 g05230(.A(new_n7578), .B(new_n7547), .Y(new_n7579));
  nand_5 g05231(.A(new_n7577), .B(new_n7546), .Y(new_n7580));
  nand_5 g05232(.A(new_n7525), .B(new_n7524_1), .Y(new_n7581));
  xor_4  g05233(.A(new_n7581), .B(new_n7529), .Y(new_n7582));
  not_8  g05234(.A(new_n7582), .Y(new_n7583));
  nand_5 g05235(.A(new_n7556), .B(new_n7557), .Y(new_n7584));
  xor_4  g05236(.A(new_n7584), .B(new_n7562), .Y(new_n7585_1));
  not_8  g05237(.A(new_n7585_1), .Y(new_n7586));
  nand_5 g05238(.A(new_n7586), .B(new_n7583), .Y(new_n7587));
  nand_5 g05239(.A(new_n7585_1), .B(new_n7582), .Y(new_n7588_1));
  or_5   g05240(.A(new_n7528), .B(n1681), .Y(new_n7589));
  and_5  g05241(.A(new_n7589), .B(new_n7529), .Y(new_n7590));
  not_8  g05242(.A(new_n7560), .Y(new_n7591));
  nand_5 g05243(.A(new_n7591), .B(new_n5468), .Y(new_n7592));
  nand_5 g05244(.A(new_n7592), .B(new_n7561), .Y(new_n7593_1));
  nor_5  g05245(.A(new_n7593_1), .B(new_n7590), .Y(new_n7594));
  nand_5 g05246(.A(new_n7594), .B(new_n7588_1), .Y(new_n7595));
  nand_5 g05247(.A(new_n7595), .B(new_n7587), .Y(new_n7596));
  nand_5 g05248(.A(new_n7596), .B(new_n7580), .Y(new_n7597));
  nand_5 g05249(.A(new_n7597), .B(new_n7579), .Y(new_n7598_1));
  nand_5 g05250(.A(new_n7544), .B(new_n7532), .Y(new_n7599));
  nand_5 g05251(.A(new_n7599), .B(new_n7543), .Y(new_n7600));
  not_8  g05252(.A(new_n7600), .Y(new_n7601));
  nand_5 g05253(.A(new_n7537), .B(new_n7535), .Y(new_n7602));
  nand_5 g05254(.A(new_n7602), .B(new_n7540), .Y(new_n7603));
  not_8  g05255(.A(new_n7603), .Y(new_n7604));
  not_8  g05256(.A(n11056), .Y(new_n7605));
  not_8  g05257(.A(n18157), .Y(new_n7606));
  nand_5 g05258(.A(new_n7606), .B(new_n7605), .Y(new_n7607_1));
  nand_5 g05259(.A(n18157), .B(n11056), .Y(new_n7608));
  nand_5 g05260(.A(new_n7608), .B(new_n7607_1), .Y(new_n7609));
  xor_4  g05261(.A(new_n7609), .B(new_n7604), .Y(new_n7610_1));
  or_5   g05262(.A(new_n7610_1), .B(new_n4886), .Y(new_n7611));
  nand_5 g05263(.A(new_n7610_1), .B(new_n4886), .Y(new_n7612));
  nand_5 g05264(.A(new_n7612), .B(new_n7611), .Y(new_n7613));
  xor_4  g05265(.A(new_n7613), .B(new_n7601), .Y(new_n7614));
  nand_5 g05266(.A(new_n7575_1), .B(new_n7564), .Y(new_n7615));
  nand_5 g05267(.A(new_n7615), .B(new_n7574), .Y(new_n7616_1));
  nand_5 g05268(.A(new_n7568), .B(new_n7566_1), .Y(new_n7617));
  nand_5 g05269(.A(new_n7617), .B(new_n7570), .Y(new_n7618));
  not_8  g05270(.A(new_n7618), .Y(new_n7619));
  not_8  g05271(.A(n10611), .Y(new_n7620));
  nand_5 g05272(.A(new_n4641), .B(new_n7620), .Y(new_n7621));
  nand_5 g05273(.A(n25797), .B(n10611), .Y(new_n7622));
  nand_5 g05274(.A(new_n7622), .B(new_n7621), .Y(new_n7623));
  xor_4  g05275(.A(new_n7623), .B(new_n7619), .Y(new_n7624));
  not_8  g05276(.A(new_n7624), .Y(new_n7625));
  nand_5 g05277(.A(new_n7625), .B(n7421), .Y(new_n7626));
  nand_5 g05278(.A(new_n7624), .B(new_n5388), .Y(new_n7627));
  nand_5 g05279(.A(new_n7627), .B(new_n7626), .Y(new_n7628));
  xor_4  g05280(.A(new_n7628), .B(new_n7616_1), .Y(new_n7629));
  nand_5 g05281(.A(new_n7629), .B(new_n7614), .Y(new_n7630_1));
  not_8  g05282(.A(new_n7614), .Y(new_n7631));
  not_8  g05283(.A(new_n7629), .Y(new_n7632));
  nand_5 g05284(.A(new_n7632), .B(new_n7631), .Y(new_n7633));
  nand_5 g05285(.A(new_n7633), .B(new_n7630_1), .Y(new_n7634));
  xor_4  g05286(.A(new_n7634), .B(new_n7598_1), .Y(n646));
  nand_5 g05287(.A(new_n2445), .B(new_n6413), .Y(new_n7636));
  nor_5  g05288(.A(new_n7636), .B(n20986), .Y(new_n7637));
  not_8  g05289(.A(new_n7637), .Y(new_n7638));
  nand_5 g05290(.A(new_n7636), .B(n20986), .Y(new_n7639));
  nand_5 g05291(.A(new_n7639), .B(new_n2450), .Y(new_n7640));
  nand_5 g05292(.A(new_n7640), .B(new_n7638), .Y(new_n7641));
  nand_5 g05293(.A(new_n2437), .B(new_n6408), .Y(new_n7642));
  nand_5 g05294(.A(new_n2438), .B(n12341), .Y(new_n7643_1));
  nand_5 g05295(.A(new_n7643_1), .B(new_n7642), .Y(new_n7644));
  xor_4  g05296(.A(new_n7644), .B(new_n7641), .Y(new_n7645));
  nand_5 g05297(.A(new_n2504), .B(new_n2506), .Y(new_n7646));
  or_5   g05298(.A(new_n7646), .B(n16223), .Y(new_n7647_1));
  nand_5 g05299(.A(new_n7646), .B(n16223), .Y(new_n7648));
  and_5  g05300(.A(new_n7648), .B(new_n7647_1), .Y(new_n7649));
  nand_5 g05301(.A(new_n7649), .B(new_n7645), .Y(new_n7650));
  not_8  g05302(.A(new_n7645), .Y(new_n7651));
  not_8  g05303(.A(new_n7649), .Y(new_n7652));
  nand_5 g05304(.A(new_n7652), .B(new_n7651), .Y(new_n7653));
  or_5   g05305(.A(new_n2445), .B(new_n6413), .Y(new_n7654));
  and_5  g05306(.A(new_n7654), .B(new_n7636), .Y(new_n7655));
  not_8  g05307(.A(new_n7655), .Y(new_n7656));
  nand_5 g05308(.A(new_n7656), .B(n2387), .Y(new_n7657_1));
  nand_5 g05309(.A(n19494), .B(n2387), .Y(new_n7658));
  and_5  g05310(.A(new_n7658), .B(new_n7646), .Y(new_n7659));
  not_8  g05311(.A(new_n7659), .Y(new_n7660));
  nand_5 g05312(.A(new_n7660), .B(new_n7657_1), .Y(new_n7661));
  or_5   g05313(.A(new_n7657_1), .B(n19494), .Y(new_n7662));
  and_5  g05314(.A(new_n7638), .B(new_n7639), .Y(new_n7663));
  xor_4  g05315(.A(new_n7663), .B(new_n2450), .Y(new_n7664));
  nand_5 g05316(.A(new_n7664), .B(new_n7662), .Y(new_n7665));
  nand_5 g05317(.A(new_n7665), .B(new_n7661), .Y(new_n7666));
  not_8  g05318(.A(new_n7666), .Y(new_n7667));
  nand_5 g05319(.A(new_n7667), .B(new_n7653), .Y(new_n7668));
  nand_5 g05320(.A(new_n7668), .B(new_n7650), .Y(new_n7669));
  nand_5 g05321(.A(new_n7643_1), .B(new_n7641), .Y(new_n7670_1));
  nand_5 g05322(.A(new_n7670_1), .B(new_n7642), .Y(new_n7671));
  nand_5 g05323(.A(new_n2431), .B(new_n6405), .Y(new_n7672));
  or_5   g05324(.A(new_n2431), .B(new_n6405), .Y(new_n7673));
  nand_5 g05325(.A(new_n7673), .B(new_n7672), .Y(new_n7674_1));
  xor_4  g05326(.A(new_n7674_1), .B(new_n7671), .Y(new_n7675));
  nor_5  g05327(.A(new_n7647_1), .B(n26913), .Y(new_n7676));
  not_8  g05328(.A(new_n7676), .Y(new_n7677));
  nand_5 g05329(.A(new_n7647_1), .B(n26913), .Y(new_n7678_1));
  and_5  g05330(.A(new_n7678_1), .B(new_n7677), .Y(new_n7679_1));
  nand_5 g05331(.A(new_n7679_1), .B(new_n7675), .Y(new_n7680));
  not_8  g05332(.A(new_n7675), .Y(new_n7681));
  not_8  g05333(.A(new_n7679_1), .Y(new_n7682));
  nand_5 g05334(.A(new_n7682), .B(new_n7681), .Y(new_n7683));
  nand_5 g05335(.A(new_n7683), .B(new_n7680), .Y(new_n7684));
  xor_4  g05336(.A(new_n7684), .B(new_n7669), .Y(new_n7685));
  or_5   g05337(.A(new_n7685), .B(new_n3641), .Y(new_n7686_1));
  nand_5 g05338(.A(new_n7685), .B(new_n3641), .Y(new_n7687));
  nand_5 g05339(.A(new_n7650), .B(new_n7653), .Y(new_n7688));
  xor_4  g05340(.A(new_n7688), .B(new_n7667), .Y(new_n7689));
  nand_5 g05341(.A(new_n7689), .B(new_n3648), .Y(new_n7690));
  or_5   g05342(.A(new_n7689), .B(new_n3648), .Y(new_n7691));
  nand_5 g05343(.A(new_n7655), .B(new_n2506), .Y(new_n7692_1));
  nand_5 g05344(.A(new_n7692_1), .B(new_n7657_1), .Y(new_n7693_1));
  nor_5  g05345(.A(new_n7693_1), .B(new_n3656), .Y(new_n7694));
  nand_5 g05346(.A(new_n7694), .B(new_n3661), .Y(new_n7695));
  not_8  g05347(.A(new_n7695), .Y(new_n7696));
  nor_5  g05348(.A(new_n7694), .B(new_n3663), .Y(new_n7697));
  not_8  g05349(.A(new_n7664), .Y(new_n7698_1));
  nand_5 g05350(.A(new_n7661), .B(new_n7662), .Y(new_n7699));
  xor_4  g05351(.A(new_n7699), .B(new_n7698_1), .Y(new_n7700));
  nor_5  g05352(.A(new_n7700), .B(new_n7697), .Y(new_n7701));
  nor_5  g05353(.A(new_n7701), .B(new_n7696), .Y(new_n7702));
  nand_5 g05354(.A(new_n7702), .B(new_n7691), .Y(new_n7703));
  and_5  g05355(.A(new_n7703), .B(new_n7690), .Y(new_n7704));
  nand_5 g05356(.A(new_n7704), .B(new_n7687), .Y(new_n7705));
  nand_5 g05357(.A(new_n7705), .B(new_n7686_1), .Y(new_n7706));
  nand_5 g05358(.A(new_n7683), .B(new_n7669), .Y(new_n7707));
  nand_5 g05359(.A(new_n7707), .B(new_n7680), .Y(new_n7708_1));
  nand_5 g05360(.A(new_n7673), .B(new_n7671), .Y(new_n7709));
  nand_5 g05361(.A(new_n7709), .B(new_n7672), .Y(new_n7710));
  not_8  g05362(.A(new_n7710), .Y(new_n7711));
  nand_5 g05363(.A(new_n2375), .B(new_n6402), .Y(new_n7712));
  nand_5 g05364(.A(new_n2374_1), .B(n7566), .Y(new_n7713));
  nand_5 g05365(.A(new_n7713), .B(new_n7712), .Y(new_n7714));
  xor_4  g05366(.A(new_n7714), .B(new_n7711), .Y(new_n7715));
  not_8  g05367(.A(new_n7715), .Y(new_n7716));
  nand_5 g05368(.A(new_n7676), .B(new_n2492), .Y(new_n7717));
  nand_5 g05369(.A(new_n7677), .B(n21832), .Y(new_n7718));
  and_5  g05370(.A(new_n7718), .B(new_n7717), .Y(new_n7719));
  nand_5 g05371(.A(new_n7719), .B(new_n7716), .Y(new_n7720));
  not_8  g05372(.A(new_n7719), .Y(new_n7721_1));
  nand_5 g05373(.A(new_n7721_1), .B(new_n7715), .Y(new_n7722));
  nand_5 g05374(.A(new_n7722), .B(new_n7720), .Y(new_n7723));
  xor_4  g05375(.A(new_n7723), .B(new_n7708_1), .Y(new_n7724));
  or_5   g05376(.A(new_n7724), .B(new_n3634), .Y(new_n7725));
  nand_5 g05377(.A(new_n7724), .B(new_n3634), .Y(new_n7726));
  nand_5 g05378(.A(new_n7726), .B(new_n7725), .Y(new_n7727));
  xnor_4 g05379(.A(new_n7727), .B(new_n7706), .Y(n696));
  not_8  g05380(.A(n20179), .Y(new_n7729));
  nand_5 g05381(.A(new_n7729), .B(new_n6246), .Y(new_n7730));
  nand_5 g05382(.A(n20179), .B(n11011), .Y(new_n7731_1));
  not_8  g05383(.A(n19228), .Y(new_n7732));
  nand_5 g05384(.A(new_n7732), .B(new_n6249), .Y(new_n7733));
  nand_5 g05385(.A(n19228), .B(n16029), .Y(new_n7734));
  not_8  g05386(.A(n15539), .Y(new_n7735));
  nand_5 g05387(.A(new_n6252), .B(new_n7735), .Y(new_n7736));
  nand_5 g05388(.A(n16476), .B(n15539), .Y(new_n7737));
  not_8  g05389(.A(n8052), .Y(new_n7738));
  nand_5 g05390(.A(new_n6255), .B(new_n7738), .Y(new_n7739));
  nand_5 g05391(.A(n11615), .B(n8052), .Y(new_n7740));
  not_8  g05392(.A(n10158), .Y(new_n7741));
  nand_5 g05393(.A(new_n6258), .B(new_n7741), .Y(new_n7742));
  nand_5 g05394(.A(n22433), .B(n10158), .Y(new_n7743));
  nand_5 g05395(.A(n18962), .B(n14090), .Y(new_n7744));
  nand_5 g05396(.A(new_n7744), .B(new_n7743), .Y(new_n7745));
  nand_5 g05397(.A(new_n7745), .B(new_n7742), .Y(new_n7746));
  nand_5 g05398(.A(new_n7746), .B(new_n7740), .Y(new_n7747));
  nand_5 g05399(.A(new_n7747), .B(new_n7739), .Y(new_n7748));
  nand_5 g05400(.A(new_n7748), .B(new_n7737), .Y(new_n7749));
  nand_5 g05401(.A(new_n7749), .B(new_n7736), .Y(new_n7750));
  nand_5 g05402(.A(new_n7750), .B(new_n7734), .Y(new_n7751_1));
  nand_5 g05403(.A(new_n7751_1), .B(new_n7733), .Y(new_n7752));
  nand_5 g05404(.A(new_n7752), .B(new_n7731_1), .Y(new_n7753));
  nand_5 g05405(.A(new_n7753), .B(new_n7730), .Y(new_n7754));
  not_8  g05406(.A(new_n7754), .Y(new_n7755));
  nand_5 g05407(.A(n12446), .B(n1112), .Y(new_n7756));
  not_8  g05408(.A(n1112), .Y(new_n7757));
  nand_5 g05409(.A(new_n4952_1), .B(new_n7757), .Y(new_n7758));
  nand_5 g05410(.A(new_n7758), .B(new_n7756), .Y(new_n7759_1));
  xor_4  g05411(.A(new_n7759_1), .B(new_n7755), .Y(new_n7760));
  not_8  g05412(.A(new_n7760), .Y(new_n7761));
  nand_5 g05413(.A(new_n7761), .B(n13490), .Y(new_n7762));
  nand_5 g05414(.A(new_n7760), .B(new_n2585), .Y(new_n7763));
  nand_5 g05415(.A(new_n7731_1), .B(new_n7730), .Y(new_n7764));
  xor_4  g05416(.A(new_n7764), .B(new_n7752), .Y(new_n7765));
  nand_5 g05417(.A(new_n7765), .B(n22660), .Y(new_n7766));
  not_8  g05418(.A(new_n7765), .Y(new_n7767));
  nand_5 g05419(.A(new_n7767), .B(new_n2467), .Y(new_n7768));
  nand_5 g05420(.A(new_n7734), .B(new_n7733), .Y(new_n7769_1));
  xor_4  g05421(.A(new_n7769_1), .B(new_n7750), .Y(new_n7770));
  nand_5 g05422(.A(new_n7770), .B(n1777), .Y(new_n7771));
  not_8  g05423(.A(new_n7770), .Y(new_n7772));
  nand_5 g05424(.A(new_n7772), .B(new_n2370), .Y(new_n7773_1));
  nand_5 g05425(.A(new_n7737), .B(new_n7736), .Y(new_n7774));
  xor_4  g05426(.A(new_n7774), .B(new_n7748), .Y(new_n7775));
  nand_5 g05427(.A(new_n7775), .B(n8745), .Y(new_n7776));
  not_8  g05428(.A(new_n7775), .Y(new_n7777));
  nand_5 g05429(.A(new_n7777), .B(new_n2349), .Y(new_n7778));
  nand_5 g05430(.A(new_n7740), .B(new_n7739), .Y(new_n7779));
  xor_4  g05431(.A(new_n7779), .B(new_n7746), .Y(new_n7780_1));
  nand_5 g05432(.A(new_n7780_1), .B(n15636), .Y(new_n7781));
  not_8  g05433(.A(new_n7780_1), .Y(new_n7782));
  nand_5 g05434(.A(new_n7782), .B(new_n2353), .Y(new_n7783));
  not_8  g05435(.A(n18962), .Y(new_n7784));
  nand_5 g05436(.A(new_n7784), .B(new_n2631), .Y(new_n7785));
  and_5  g05437(.A(new_n7785), .B(new_n7744), .Y(new_n7786));
  nand_5 g05438(.A(new_n7786), .B(n6794), .Y(new_n7787));
  nand_5 g05439(.A(new_n7787), .B(new_n2358), .Y(new_n7788_1));
  or_5   g05440(.A(new_n7787), .B(new_n2358), .Y(new_n7789));
  nand_5 g05441(.A(new_n7743), .B(new_n7742), .Y(new_n7790));
  xor_4  g05442(.A(new_n7790), .B(new_n7744), .Y(new_n7791));
  not_8  g05443(.A(new_n7791), .Y(new_n7792));
  nand_5 g05444(.A(new_n7792), .B(new_n7789), .Y(new_n7793));
  nand_5 g05445(.A(new_n7793), .B(new_n7788_1), .Y(new_n7794_1));
  not_8  g05446(.A(new_n7794_1), .Y(new_n7795));
  nand_5 g05447(.A(new_n7795), .B(new_n7783), .Y(new_n7796));
  nand_5 g05448(.A(new_n7796), .B(new_n7781), .Y(new_n7797));
  nand_5 g05449(.A(new_n7797), .B(new_n7778), .Y(new_n7798));
  nand_5 g05450(.A(new_n7798), .B(new_n7776), .Y(new_n7799));
  nand_5 g05451(.A(new_n7799), .B(new_n7773_1), .Y(new_n7800));
  nand_5 g05452(.A(new_n7800), .B(new_n7771), .Y(new_n7801));
  nand_5 g05453(.A(new_n7801), .B(new_n7768), .Y(new_n7802));
  nand_5 g05454(.A(new_n7802), .B(new_n7766), .Y(new_n7803));
  nand_5 g05455(.A(new_n7803), .B(new_n7763), .Y(new_n7804));
  nand_5 g05456(.A(new_n7804), .B(new_n7762), .Y(new_n7805));
  nand_5 g05457(.A(new_n7756), .B(new_n7754), .Y(new_n7806));
  nand_5 g05458(.A(new_n7806), .B(new_n7758), .Y(new_n7807));
  not_8  g05459(.A(new_n7807), .Y(new_n7808));
  nand_5 g05460(.A(n23849), .B(n2289), .Y(new_n7809));
  not_8  g05461(.A(n2289), .Y(new_n7810));
  nand_5 g05462(.A(new_n6240), .B(new_n7810), .Y(new_n7811_1));
  nand_5 g05463(.A(new_n7811_1), .B(new_n7809), .Y(new_n7812));
  xor_4  g05464(.A(new_n7812), .B(new_n7808), .Y(new_n7813));
  not_8  g05465(.A(new_n7813), .Y(new_n7814));
  nand_5 g05466(.A(new_n7814), .B(n9655), .Y(new_n7815));
  nand_5 g05467(.A(new_n7813), .B(new_n6242), .Y(new_n7816));
  nand_5 g05468(.A(new_n7816), .B(new_n7815), .Y(new_n7817));
  xnor_4 g05469(.A(new_n7817), .B(new_n7805), .Y(new_n7818));
  not_8  g05470(.A(n19042), .Y(new_n7819));
  nand_5 g05471(.A(new_n4512), .B(new_n7819), .Y(new_n7820));
  nand_5 g05472(.A(n20151), .B(n19042), .Y(new_n7821));
  not_8  g05473(.A(n19472), .Y(new_n7822));
  nand_5 g05474(.A(new_n7822), .B(new_n4438), .Y(new_n7823));
  nand_5 g05475(.A(n19472), .B(n7693), .Y(new_n7824));
  not_8  g05476(.A(n25370), .Y(new_n7825));
  nand_5 g05477(.A(new_n7825), .B(new_n4396), .Y(new_n7826));
  nand_5 g05478(.A(n25370), .B(n10405), .Y(new_n7827));
  nand_5 g05479(.A(new_n4598), .B(new_n4594), .Y(new_n7828));
  nand_5 g05480(.A(new_n7828), .B(new_n4597), .Y(new_n7829));
  nand_5 g05481(.A(new_n7829), .B(new_n7827), .Y(new_n7830_1));
  nand_5 g05482(.A(new_n7830_1), .B(new_n7826), .Y(new_n7831));
  nand_5 g05483(.A(new_n7831), .B(new_n7824), .Y(new_n7832));
  nand_5 g05484(.A(new_n7832), .B(new_n7823), .Y(new_n7833));
  nand_5 g05485(.A(new_n7833), .B(new_n7821), .Y(new_n7834_1));
  nand_5 g05486(.A(new_n7834_1), .B(new_n7820), .Y(new_n7835));
  not_8  g05487(.A(new_n7835), .Y(new_n7836));
  nand_5 g05488(.A(n8964), .B(n1293), .Y(new_n7837));
  not_8  g05489(.A(n1293), .Y(new_n7838));
  nand_5 g05490(.A(new_n6394), .B(new_n7838), .Y(new_n7839));
  nand_5 g05491(.A(new_n7839), .B(new_n7837), .Y(new_n7840));
  xor_4  g05492(.A(new_n7840), .B(new_n7836), .Y(new_n7841_1));
  not_8  g05493(.A(new_n7841_1), .Y(new_n7842));
  nand_5 g05494(.A(new_n7842), .B(n23200), .Y(new_n7843));
  nand_5 g05495(.A(new_n7841_1), .B(new_n6396), .Y(new_n7844));
  nand_5 g05496(.A(new_n7821), .B(new_n7820), .Y(new_n7845));
  xor_4  g05497(.A(new_n7845), .B(new_n7833), .Y(new_n7846));
  nand_5 g05498(.A(new_n7846), .B(n17959), .Y(new_n7847));
  not_8  g05499(.A(new_n7846), .Y(new_n7848));
  nand_5 g05500(.A(new_n7848), .B(new_n6399), .Y(new_n7849));
  nand_5 g05501(.A(new_n7824), .B(new_n7823), .Y(new_n7850));
  xor_4  g05502(.A(new_n7850), .B(new_n7831), .Y(new_n7851));
  nand_5 g05503(.A(new_n7851), .B(n7566), .Y(new_n7852));
  not_8  g05504(.A(new_n7851), .Y(new_n7853));
  nand_5 g05505(.A(new_n7853), .B(new_n6402), .Y(new_n7854));
  nand_5 g05506(.A(new_n7827), .B(new_n7826), .Y(new_n7855));
  xor_4  g05507(.A(new_n7855), .B(new_n7829), .Y(new_n7856));
  nand_5 g05508(.A(new_n7856), .B(n7731), .Y(new_n7857));
  not_8  g05509(.A(new_n7856), .Y(new_n7858));
  nand_5 g05510(.A(new_n7858), .B(new_n6405), .Y(new_n7859));
  nand_5 g05511(.A(new_n4612), .B(n12341), .Y(new_n7860));
  nand_5 g05512(.A(new_n4600), .B(new_n6408), .Y(new_n7861));
  nand_5 g05513(.A(new_n4566), .B(n20986), .Y(new_n7862));
  nand_5 g05514(.A(new_n4557), .B(new_n6411), .Y(new_n7863));
  nand_5 g05515(.A(new_n4544), .B(n12384), .Y(new_n7864));
  not_8  g05516(.A(new_n7864), .Y(new_n7865));
  nand_5 g05517(.A(new_n7865), .B(new_n7863), .Y(new_n7866));
  nand_5 g05518(.A(new_n7866), .B(new_n7862), .Y(new_n7867));
  nand_5 g05519(.A(new_n7867), .B(new_n7861), .Y(new_n7868));
  nand_5 g05520(.A(new_n7868), .B(new_n7860), .Y(new_n7869));
  nand_5 g05521(.A(new_n7869), .B(new_n7859), .Y(new_n7870));
  nand_5 g05522(.A(new_n7870), .B(new_n7857), .Y(new_n7871));
  nand_5 g05523(.A(new_n7871), .B(new_n7854), .Y(new_n7872));
  nand_5 g05524(.A(new_n7872), .B(new_n7852), .Y(new_n7873));
  nand_5 g05525(.A(new_n7873), .B(new_n7849), .Y(new_n7874));
  nand_5 g05526(.A(new_n7874), .B(new_n7847), .Y(new_n7875));
  nand_5 g05527(.A(new_n7875), .B(new_n7844), .Y(new_n7876_1));
  nand_5 g05528(.A(new_n7876_1), .B(new_n7843), .Y(new_n7877));
  nand_5 g05529(.A(new_n7837), .B(new_n7835), .Y(new_n7878));
  nand_5 g05530(.A(new_n7878), .B(new_n7839), .Y(new_n7879));
  not_8  g05531(.A(new_n7879), .Y(new_n7880));
  nand_5 g05532(.A(n27037), .B(n13775), .Y(new_n7881));
  not_8  g05533(.A(n13775), .Y(new_n7882));
  nand_5 g05534(.A(new_n6390), .B(new_n7882), .Y(new_n7883));
  nand_5 g05535(.A(new_n7883), .B(new_n7881), .Y(new_n7884_1));
  xor_4  g05536(.A(new_n7884_1), .B(new_n7880), .Y(new_n7885));
  not_8  g05537(.A(new_n7885), .Y(new_n7886));
  nand_5 g05538(.A(new_n7886), .B(n11736), .Y(new_n7887));
  nand_5 g05539(.A(new_n7885), .B(new_n6392), .Y(new_n7888));
  nand_5 g05540(.A(new_n7888), .B(new_n7887), .Y(new_n7889));
  xor_4  g05541(.A(new_n7889), .B(new_n7877), .Y(new_n7890));
  or_5   g05542(.A(new_n7890), .B(new_n7818), .Y(new_n7891));
  nand_5 g05543(.A(new_n7890), .B(new_n7818), .Y(new_n7892));
  nand_5 g05544(.A(new_n7763), .B(new_n7762), .Y(new_n7893));
  xor_4  g05545(.A(new_n7893), .B(new_n7803), .Y(new_n7894));
  not_8  g05546(.A(new_n7894), .Y(new_n7895));
  nand_5 g05547(.A(new_n7843), .B(new_n7844), .Y(new_n7896));
  xor_4  g05548(.A(new_n7896), .B(new_n7875), .Y(new_n7897));
  or_5   g05549(.A(new_n7897), .B(new_n7895), .Y(new_n7898));
  nand_5 g05550(.A(new_n7897), .B(new_n7895), .Y(new_n7899));
  nand_5 g05551(.A(new_n7768), .B(new_n7766), .Y(new_n7900));
  xor_4  g05552(.A(new_n7900), .B(new_n7801), .Y(new_n7901));
  not_8  g05553(.A(new_n7901), .Y(new_n7902));
  nand_5 g05554(.A(new_n7847), .B(new_n7849), .Y(new_n7903));
  xor_4  g05555(.A(new_n7903), .B(new_n7873), .Y(new_n7904));
  or_5   g05556(.A(new_n7904), .B(new_n7902), .Y(new_n7905));
  nand_5 g05557(.A(new_n7904), .B(new_n7902), .Y(new_n7906));
  nand_5 g05558(.A(new_n7773_1), .B(new_n7771), .Y(new_n7907));
  xor_4  g05559(.A(new_n7907), .B(new_n7799), .Y(new_n7908));
  not_8  g05560(.A(new_n7908), .Y(new_n7909));
  nand_5 g05561(.A(new_n7852), .B(new_n7854), .Y(new_n7910));
  xor_4  g05562(.A(new_n7910), .B(new_n7871), .Y(new_n7911));
  or_5   g05563(.A(new_n7911), .B(new_n7909), .Y(new_n7912));
  nand_5 g05564(.A(new_n7911), .B(new_n7909), .Y(new_n7913));
  nand_5 g05565(.A(new_n7778), .B(new_n7776), .Y(new_n7914));
  xor_4  g05566(.A(new_n7914), .B(new_n7797), .Y(new_n7915));
  not_8  g05567(.A(new_n7915), .Y(new_n7916));
  nand_5 g05568(.A(new_n7857), .B(new_n7859), .Y(new_n7917_1));
  xor_4  g05569(.A(new_n7917_1), .B(new_n7869), .Y(new_n7918));
  or_5   g05570(.A(new_n7918), .B(new_n7916), .Y(new_n7919));
  nand_5 g05571(.A(new_n7918), .B(new_n7916), .Y(new_n7920));
  nand_5 g05572(.A(new_n7783), .B(new_n7781), .Y(new_n7921));
  xor_4  g05573(.A(new_n7921), .B(new_n7794_1), .Y(new_n7922));
  nand_5 g05574(.A(new_n7860), .B(new_n7861), .Y(new_n7923));
  xor_4  g05575(.A(new_n7923), .B(new_n7867), .Y(new_n7924));
  or_5   g05576(.A(new_n7924), .B(new_n7922), .Y(new_n7925));
  nand_5 g05577(.A(new_n7924), .B(new_n7922), .Y(new_n7926));
  nand_5 g05578(.A(new_n7788_1), .B(new_n7789), .Y(new_n7927));
  xor_4  g05579(.A(new_n7927), .B(new_n7792), .Y(new_n7928));
  nand_5 g05580(.A(new_n7862), .B(new_n7863), .Y(new_n7929));
  xor_4  g05581(.A(new_n7929), .B(new_n7865), .Y(new_n7930));
  or_5   g05582(.A(new_n7930), .B(new_n7928), .Y(new_n7931));
  nand_5 g05583(.A(new_n7930), .B(new_n7928), .Y(new_n7932));
  not_8  g05584(.A(new_n7786), .Y(new_n7933));
  nand_5 g05585(.A(new_n7933), .B(new_n2442), .Y(new_n7934));
  and_5  g05586(.A(new_n7934), .B(new_n7787), .Y(new_n7935));
  nand_5 g05587(.A(new_n4578), .B(new_n6413), .Y(new_n7936));
  nand_5 g05588(.A(new_n7936), .B(new_n7864), .Y(new_n7937_1));
  nand_5 g05589(.A(new_n7937_1), .B(new_n7935), .Y(new_n7938));
  nand_5 g05590(.A(new_n7938), .B(new_n7932), .Y(new_n7939));
  nand_5 g05591(.A(new_n7939), .B(new_n7931), .Y(new_n7940));
  nand_5 g05592(.A(new_n7940), .B(new_n7926), .Y(new_n7941));
  nand_5 g05593(.A(new_n7941), .B(new_n7925), .Y(new_n7942));
  nand_5 g05594(.A(new_n7942), .B(new_n7920), .Y(new_n7943_1));
  nand_5 g05595(.A(new_n7943_1), .B(new_n7919), .Y(new_n7944));
  nand_5 g05596(.A(new_n7944), .B(new_n7913), .Y(new_n7945));
  nand_5 g05597(.A(new_n7945), .B(new_n7912), .Y(new_n7946));
  nand_5 g05598(.A(new_n7946), .B(new_n7906), .Y(new_n7947));
  nand_5 g05599(.A(new_n7947), .B(new_n7905), .Y(new_n7948));
  nand_5 g05600(.A(new_n7948), .B(new_n7899), .Y(new_n7949_1));
  nand_5 g05601(.A(new_n7949_1), .B(new_n7898), .Y(new_n7950_1));
  nand_5 g05602(.A(new_n7950_1), .B(new_n7892), .Y(new_n7951));
  nand_5 g05603(.A(new_n7951), .B(new_n7891), .Y(new_n7952));
  nand_5 g05604(.A(new_n7816), .B(new_n7805), .Y(new_n7953));
  nand_5 g05605(.A(new_n7953), .B(new_n7815), .Y(new_n7954));
  nand_5 g05606(.A(new_n7809), .B(new_n7807), .Y(new_n7955));
  nand_5 g05607(.A(new_n7955), .B(new_n7811_1), .Y(new_n7956));
  not_8  g05608(.A(new_n7956), .Y(new_n7957));
  not_8  g05609(.A(n23697), .Y(new_n7958));
  nand_5 g05610(.A(new_n4942), .B(new_n7958), .Y(new_n7959_1));
  nand_5 g05611(.A(n25475), .B(n23697), .Y(new_n7960));
  nand_5 g05612(.A(new_n7960), .B(new_n7959_1), .Y(new_n7961));
  xor_4  g05613(.A(new_n7961), .B(new_n7957), .Y(new_n7962));
  not_8  g05614(.A(new_n7962), .Y(new_n7963_1));
  nand_5 g05615(.A(new_n7963_1), .B(n25345), .Y(new_n7964));
  nand_5 g05616(.A(new_n7962), .B(new_n6238), .Y(new_n7965));
  nand_5 g05617(.A(new_n7965), .B(new_n7964), .Y(new_n7966));
  xor_4  g05618(.A(new_n7966), .B(new_n7954), .Y(new_n7967));
  not_8  g05619(.A(new_n7967), .Y(new_n7968_1));
  nand_5 g05620(.A(new_n7888), .B(new_n7877), .Y(new_n7969));
  nand_5 g05621(.A(new_n7969), .B(new_n7887), .Y(new_n7970));
  nand_5 g05622(.A(new_n7881), .B(new_n7879), .Y(new_n7971));
  nand_5 g05623(.A(new_n7971), .B(new_n7883), .Y(new_n7972));
  not_8  g05624(.A(new_n7972), .Y(new_n7973));
  not_8  g05625(.A(n21915), .Y(new_n7974));
  nand_5 g05626(.A(new_n7974), .B(new_n6386), .Y(new_n7975));
  nand_5 g05627(.A(n21915), .B(n15182), .Y(new_n7976));
  nand_5 g05628(.A(new_n7976), .B(new_n7975), .Y(new_n7977));
  xor_4  g05629(.A(new_n7977), .B(new_n7973), .Y(new_n7978));
  not_8  g05630(.A(new_n7978), .Y(new_n7979));
  nand_5 g05631(.A(new_n7979), .B(n17351), .Y(new_n7980));
  nand_5 g05632(.A(new_n7978), .B(new_n6388), .Y(new_n7981));
  nand_5 g05633(.A(new_n7981), .B(new_n7980), .Y(new_n7982));
  xor_4  g05634(.A(new_n7982), .B(new_n7970), .Y(new_n7983));
  nand_5 g05635(.A(new_n7983), .B(new_n7968_1), .Y(new_n7984));
  not_8  g05636(.A(new_n7984), .Y(new_n7985));
  or_5   g05637(.A(new_n7983), .B(new_n7968_1), .Y(new_n7986));
  not_8  g05638(.A(new_n7986), .Y(new_n7987));
  nor_5  g05639(.A(new_n7987), .B(new_n7985), .Y(new_n7988));
  xor_4  g05640(.A(new_n7988), .B(new_n7952), .Y(n723));
  not_8  g05641(.A(n8305), .Y(new_n7990));
  not_8  g05642(.A(n8856), .Y(new_n7991));
  nand_5 g05643(.A(new_n7991), .B(new_n7990), .Y(new_n7992_1));
  nand_5 g05644(.A(n8856), .B(n8305), .Y(new_n7993));
  not_8  g05645(.A(n12861), .Y(new_n7994));
  nand_5 g05646(.A(new_n3849), .B(new_n7994), .Y(new_n7995));
  nand_5 g05647(.A(n14130), .B(n12861), .Y(new_n7996));
  not_8  g05648(.A(n13333), .Y(new_n7997));
  not_8  g05649(.A(n16482), .Y(new_n7998));
  nand_5 g05650(.A(new_n7998), .B(new_n7997), .Y(new_n7999_1));
  nand_5 g05651(.A(n16482), .B(n13333), .Y(new_n8000));
  not_8  g05652(.A(n2210), .Y(new_n8001));
  nand_5 g05653(.A(new_n2599), .B(new_n8001), .Y(new_n8002));
  nand_5 g05654(.A(n9942), .B(n2210), .Y(new_n8003));
  nand_5 g05655(.A(new_n5864), .B(new_n5862), .Y(new_n8004));
  nand_5 g05656(.A(new_n8004), .B(new_n5863), .Y(new_n8005));
  nand_5 g05657(.A(new_n8005), .B(new_n8003), .Y(new_n8006_1));
  nand_5 g05658(.A(new_n8006_1), .B(new_n8002), .Y(new_n8007));
  nand_5 g05659(.A(new_n8007), .B(new_n8000), .Y(new_n8008));
  nand_5 g05660(.A(new_n8008), .B(new_n7999_1), .Y(new_n8009));
  nand_5 g05661(.A(new_n8009), .B(new_n7996), .Y(new_n8010));
  nand_5 g05662(.A(new_n8010), .B(new_n7995), .Y(new_n8011));
  nand_5 g05663(.A(new_n8011), .B(new_n7993), .Y(new_n8012));
  nand_5 g05664(.A(new_n8012), .B(new_n7992_1), .Y(new_n8013));
  not_8  g05665(.A(new_n8013), .Y(new_n8014));
  not_8  g05666(.A(n22253), .Y(new_n8015));
  not_8  g05667(.A(n22442), .Y(new_n8016));
  nand_5 g05668(.A(new_n8016), .B(new_n8015), .Y(new_n8017));
  nand_5 g05669(.A(n22442), .B(n22253), .Y(new_n8018));
  not_8  g05670(.A(n468), .Y(new_n8019));
  not_8  g05671(.A(n1255), .Y(new_n8020));
  nand_5 g05672(.A(new_n8020), .B(new_n8019), .Y(new_n8021));
  nand_5 g05673(.A(n1255), .B(n468), .Y(new_n8022));
  not_8  g05674(.A(n5400), .Y(new_n8023));
  not_8  g05675(.A(n9512), .Y(new_n8024));
  nand_5 g05676(.A(new_n8024), .B(new_n8023), .Y(new_n8025));
  nand_5 g05677(.A(n9512), .B(n5400), .Y(new_n8026));
  not_8  g05678(.A(n16608), .Y(new_n8027_1));
  not_8  g05679(.A(n23923), .Y(new_n8028));
  nand_5 g05680(.A(new_n8028), .B(new_n8027_1), .Y(new_n8029));
  nand_5 g05681(.A(n23923), .B(n16608), .Y(new_n8030));
  not_8  g05682(.A(n329), .Y(new_n8031_1));
  nand_5 g05683(.A(new_n5317), .B(new_n8031_1), .Y(new_n8032));
  nand_5 g05684(.A(n21735), .B(n329), .Y(new_n8033));
  not_8  g05685(.A(n2409), .Y(new_n8034));
  not_8  g05686(.A(n8869), .Y(new_n8035));
  nand_5 g05687(.A(new_n8035), .B(new_n5230), .Y(new_n8036));
  nand_5 g05688(.A(n8869), .B(n1738), .Y(new_n8037));
  not_8  g05689(.A(n10372), .Y(new_n8038));
  nand_5 g05690(.A(new_n5234), .B(new_n8038), .Y(new_n8039));
  nand_5 g05691(.A(n12152), .B(n10372), .Y(new_n8040));
  nand_5 g05692(.A(n19107), .B(n7428), .Y(new_n8041));
  nand_5 g05693(.A(new_n8041), .B(new_n8040), .Y(new_n8042_1));
  nand_5 g05694(.A(new_n8042_1), .B(new_n8039), .Y(new_n8043));
  nand_5 g05695(.A(new_n8043), .B(new_n8037), .Y(new_n8044));
  nand_5 g05696(.A(new_n8044), .B(new_n8036), .Y(new_n8045));
  nand_5 g05697(.A(new_n8045), .B(new_n8034), .Y(new_n8046));
  not_8  g05698(.A(new_n8046), .Y(new_n8047));
  nor_5  g05699(.A(new_n8045), .B(new_n8034), .Y(new_n8048));
  nor_5  g05700(.A(new_n8048), .B(n14071), .Y(new_n8049));
  nor_5  g05701(.A(new_n8049), .B(new_n8047), .Y(new_n8050));
  or_5   g05702(.A(new_n8050), .B(n24085), .Y(new_n8051));
  not_8  g05703(.A(n24170), .Y(new_n8052_1));
  nand_5 g05704(.A(new_n8050), .B(n24085), .Y(new_n8053));
  nand_5 g05705(.A(new_n8053), .B(new_n8052_1), .Y(new_n8054));
  nand_5 g05706(.A(new_n8054), .B(new_n8051), .Y(new_n8055));
  nand_5 g05707(.A(new_n8055), .B(new_n8033), .Y(new_n8056));
  nand_5 g05708(.A(new_n8056), .B(new_n8032), .Y(new_n8057));
  nand_5 g05709(.A(new_n8057), .B(new_n8030), .Y(new_n8058));
  nand_5 g05710(.A(new_n8058), .B(new_n8029), .Y(new_n8059));
  nand_5 g05711(.A(new_n8059), .B(new_n8026), .Y(new_n8060));
  nand_5 g05712(.A(new_n8060), .B(new_n8025), .Y(new_n8061));
  nand_5 g05713(.A(new_n8061), .B(new_n8022), .Y(new_n8062));
  nand_5 g05714(.A(new_n8062), .B(new_n8021), .Y(new_n8063));
  nand_5 g05715(.A(new_n8063), .B(new_n8018), .Y(new_n8064));
  nand_5 g05716(.A(new_n8064), .B(new_n8017), .Y(new_n8065));
  nand_5 g05717(.A(new_n8065), .B(new_n8014), .Y(new_n8066));
  nor_5  g05718(.A(new_n8065), .B(new_n8014), .Y(new_n8067_1));
  not_8  g05719(.A(new_n8067_1), .Y(new_n8068));
  nand_5 g05720(.A(new_n8068), .B(new_n8066), .Y(new_n8069));
  nand_5 g05721(.A(new_n7993), .B(new_n7992_1), .Y(new_n8070));
  xor_4  g05722(.A(new_n8070), .B(new_n8011), .Y(new_n8071));
  nand_5 g05723(.A(new_n8018), .B(new_n8017), .Y(new_n8072));
  xnor_4 g05724(.A(new_n8072), .B(new_n8063), .Y(new_n8073));
  or_5   g05725(.A(new_n8073), .B(new_n8071), .Y(new_n8074));
  nand_5 g05726(.A(new_n8073), .B(new_n8071), .Y(new_n8075));
  nand_5 g05727(.A(new_n7996), .B(new_n7995), .Y(new_n8076));
  xor_4  g05728(.A(new_n8076), .B(new_n8009), .Y(new_n8077));
  not_8  g05729(.A(new_n8077), .Y(new_n8078));
  nand_5 g05730(.A(new_n8022), .B(new_n8021), .Y(new_n8079));
  xor_4  g05731(.A(new_n8079), .B(new_n8061), .Y(new_n8080));
  nand_5 g05732(.A(new_n8080), .B(new_n8078), .Y(new_n8081));
  or_5   g05733(.A(new_n8080), .B(new_n8078), .Y(new_n8082));
  nand_5 g05734(.A(new_n8000), .B(new_n7999_1), .Y(new_n8083));
  xor_4  g05735(.A(new_n8083), .B(new_n8007), .Y(new_n8084));
  not_8  g05736(.A(new_n8084), .Y(new_n8085));
  nand_5 g05737(.A(new_n8026), .B(new_n8025), .Y(new_n8086));
  xor_4  g05738(.A(new_n8086), .B(new_n8059), .Y(new_n8087));
  nand_5 g05739(.A(new_n8087), .B(new_n8085), .Y(new_n8088));
  or_5   g05740(.A(new_n8087), .B(new_n8085), .Y(new_n8089));
  nand_5 g05741(.A(new_n8003), .B(new_n8002), .Y(new_n8090));
  xor_4  g05742(.A(new_n8090), .B(new_n8005), .Y(new_n8091));
  nand_5 g05743(.A(new_n8030), .B(new_n8029), .Y(new_n8092));
  xor_4  g05744(.A(new_n8092), .B(new_n8057), .Y(new_n8093));
  not_8  g05745(.A(new_n8093), .Y(new_n8094));
  or_5   g05746(.A(new_n8094), .B(new_n8091), .Y(new_n8095_1));
  nand_5 g05747(.A(new_n8094), .B(new_n8091), .Y(new_n8096));
  nand_5 g05748(.A(new_n8033), .B(new_n8032), .Y(new_n8097));
  xnor_4 g05749(.A(new_n8097), .B(new_n8055), .Y(new_n8098));
  or_5   g05750(.A(new_n8098), .B(new_n5866), .Y(new_n8099));
  nand_5 g05751(.A(new_n8098), .B(new_n5866), .Y(new_n8100));
  and_5  g05752(.A(new_n8053), .B(new_n8051), .Y(new_n8101));
  xor_4  g05753(.A(new_n8101), .B(new_n8052_1), .Y(new_n8102));
  or_5   g05754(.A(new_n8102), .B(new_n5796), .Y(new_n8103_1));
  nand_5 g05755(.A(new_n8102), .B(new_n5796), .Y(new_n8104));
  nor_5  g05756(.A(new_n8048), .B(new_n8047), .Y(new_n8105));
  xor_4  g05757(.A(new_n8105), .B(new_n5226_1), .Y(new_n8106));
  or_5   g05758(.A(new_n8106), .B(new_n5765_1), .Y(new_n8107));
  nand_5 g05759(.A(new_n8106), .B(new_n5765_1), .Y(new_n8108));
  nand_5 g05760(.A(new_n8037), .B(new_n8036), .Y(new_n8109_1));
  xor_4  g05761(.A(new_n8109_1), .B(new_n8043), .Y(new_n8110));
  nand_5 g05762(.A(new_n8110), .B(new_n5757), .Y(new_n8111));
  or_5   g05763(.A(new_n8110), .B(new_n5757), .Y(new_n8112));
  nand_5 g05764(.A(new_n8040), .B(new_n8039), .Y(new_n8113));
  xor_4  g05765(.A(new_n8113), .B(new_n8041), .Y(new_n8114));
  nand_5 g05766(.A(new_n8114), .B(new_n5749), .Y(new_n8115));
  or_5   g05767(.A(new_n8114), .B(new_n5749), .Y(new_n8116));
  xor_4  g05768(.A(n19107), .B(n7428), .Y(new_n8117));
  nor_5  g05769(.A(new_n8117), .B(new_n5745), .Y(new_n8118));
  not_8  g05770(.A(new_n8118), .Y(new_n8119));
  nand_5 g05771(.A(new_n8119), .B(new_n8116), .Y(new_n8120));
  nand_5 g05772(.A(new_n8120), .B(new_n8115), .Y(new_n8121));
  nand_5 g05773(.A(new_n8121), .B(new_n8112), .Y(new_n8122));
  nand_5 g05774(.A(new_n8122), .B(new_n8111), .Y(new_n8123));
  nand_5 g05775(.A(new_n8123), .B(new_n8108), .Y(new_n8124));
  nand_5 g05776(.A(new_n8124), .B(new_n8107), .Y(new_n8125));
  nand_5 g05777(.A(new_n8125), .B(new_n8104), .Y(new_n8126));
  nand_5 g05778(.A(new_n8126), .B(new_n8103_1), .Y(new_n8127_1));
  nand_5 g05779(.A(new_n8127_1), .B(new_n8100), .Y(new_n8128));
  nand_5 g05780(.A(new_n8128), .B(new_n8099), .Y(new_n8129));
  nand_5 g05781(.A(new_n8129), .B(new_n8096), .Y(new_n8130_1));
  nand_5 g05782(.A(new_n8130_1), .B(new_n8095_1), .Y(new_n8131));
  nand_5 g05783(.A(new_n8131), .B(new_n8089), .Y(new_n8132));
  nand_5 g05784(.A(new_n8132), .B(new_n8088), .Y(new_n8133));
  nand_5 g05785(.A(new_n8133), .B(new_n8082), .Y(new_n8134));
  nand_5 g05786(.A(new_n8134), .B(new_n8081), .Y(new_n8135_1));
  nand_5 g05787(.A(new_n8135_1), .B(new_n8075), .Y(new_n8136));
  nand_5 g05788(.A(new_n8136), .B(new_n8074), .Y(new_n8137));
  xor_4  g05789(.A(new_n8137), .B(new_n8069), .Y(new_n8138));
  not_8  g05790(.A(new_n8138), .Y(new_n8139_1));
  not_8  g05791(.A(n26986), .Y(new_n8140));
  nand_5 g05792(.A(new_n8140), .B(n2272), .Y(new_n8141));
  not_8  g05793(.A(n2272), .Y(new_n8142));
  nand_5 g05794(.A(n26986), .B(new_n8142), .Y(new_n8143));
  not_8  g05795(.A(n21287), .Y(new_n8144));
  nand_5 g05796(.A(n25331), .B(new_n8144), .Y(new_n8145));
  not_8  g05797(.A(n25331), .Y(new_n8146));
  nand_5 g05798(.A(new_n8146), .B(n21287), .Y(new_n8147));
  not_8  g05799(.A(n4256), .Y(new_n8148_1));
  nand_5 g05800(.A(n18483), .B(new_n8148_1), .Y(new_n8149_1));
  not_8  g05801(.A(n18483), .Y(new_n8150));
  nand_5 g05802(.A(new_n8150), .B(n4256), .Y(new_n8151));
  nand_5 g05803(.A(new_n2569), .B(n21934), .Y(new_n8152));
  not_8  g05804(.A(n21934), .Y(new_n8153));
  nand_5 g05805(.A(n22332), .B(new_n8153), .Y(new_n8154));
  nand_5 g05806(.A(new_n2474), .B(n18901), .Y(new_n8155));
  not_8  g05807(.A(n18901), .Y(new_n8156));
  nand_5 g05808(.A(n18907), .B(new_n8156), .Y(new_n8157));
  nand_5 g05809(.A(n4376), .B(new_n2411), .Y(new_n8158));
  not_8  g05810(.A(n4376), .Y(new_n8159_1));
  nand_5 g05811(.A(new_n8159_1), .B(n2731), .Y(new_n8160));
  nand_5 g05812(.A(new_n2402), .B(n14570), .Y(new_n8161));
  not_8  g05813(.A(n14570), .Y(new_n8162));
  nand_5 g05814(.A(n19911), .B(new_n8162), .Y(new_n8163));
  nand_5 g05815(.A(n23775), .B(new_n2393), .Y(new_n8164));
  not_8  g05816(.A(n23775), .Y(new_n8165));
  nand_5 g05817(.A(new_n8165), .B(n13708), .Y(new_n8166));
  nand_5 g05818(.A(new_n2384), .B(n8259), .Y(new_n8167));
  not_8  g05819(.A(n8259), .Y(new_n8168));
  nand_5 g05820(.A(n18409), .B(new_n8168), .Y(new_n8169));
  not_8  g05821(.A(n11479), .Y(new_n8170));
  nand_5 g05822(.A(new_n8170), .B(n5704), .Y(new_n8171));
  nand_5 g05823(.A(new_n8171), .B(new_n8169), .Y(new_n8172));
  nand_5 g05824(.A(new_n8172), .B(new_n8167), .Y(new_n8173));
  nand_5 g05825(.A(new_n8173), .B(new_n8166), .Y(new_n8174));
  nand_5 g05826(.A(new_n8174), .B(new_n8164), .Y(new_n8175));
  nand_5 g05827(.A(new_n8175), .B(new_n8163), .Y(new_n8176));
  nand_5 g05828(.A(new_n8176), .B(new_n8161), .Y(new_n8177));
  nand_5 g05829(.A(new_n8177), .B(new_n8160), .Y(new_n8178));
  nand_5 g05830(.A(new_n8178), .B(new_n8158), .Y(new_n8179_1));
  nand_5 g05831(.A(new_n8179_1), .B(new_n8157), .Y(new_n8180));
  nand_5 g05832(.A(new_n8180), .B(new_n8155), .Y(new_n8181));
  nand_5 g05833(.A(new_n8181), .B(new_n8154), .Y(new_n8182));
  nand_5 g05834(.A(new_n8182), .B(new_n8152), .Y(new_n8183));
  nand_5 g05835(.A(new_n8183), .B(new_n8151), .Y(new_n8184));
  nand_5 g05836(.A(new_n8184), .B(new_n8149_1), .Y(new_n8185));
  nand_5 g05837(.A(new_n8185), .B(new_n8147), .Y(new_n8186));
  nand_5 g05838(.A(new_n8186), .B(new_n8145), .Y(new_n8187));
  nand_5 g05839(.A(new_n8187), .B(new_n8143), .Y(new_n8188));
  nand_5 g05840(.A(new_n8188), .B(new_n8141), .Y(new_n8189));
  nand_5 g05841(.A(new_n8189), .B(new_n8139_1), .Y(new_n8190));
  not_8  g05842(.A(new_n8190), .Y(new_n8191));
  nor_5  g05843(.A(new_n8189), .B(new_n8139_1), .Y(new_n8192));
  nor_5  g05844(.A(new_n8192), .B(new_n8191), .Y(new_n8193));
  nand_5 g05845(.A(new_n8143), .B(new_n8141), .Y(new_n8194_1));
  xor_4  g05846(.A(new_n8194_1), .B(new_n8187), .Y(new_n8195));
  nand_5 g05847(.A(new_n8075), .B(new_n8074), .Y(new_n8196));
  xor_4  g05848(.A(new_n8196), .B(new_n8135_1), .Y(new_n8197));
  nand_5 g05849(.A(new_n8197), .B(new_n8195), .Y(new_n8198));
  or_5   g05850(.A(new_n8197), .B(new_n8195), .Y(new_n8199));
  nand_5 g05851(.A(new_n8147), .B(new_n8145), .Y(new_n8200));
  xor_4  g05852(.A(new_n8200), .B(new_n8185), .Y(new_n8201));
  nand_5 g05853(.A(new_n8082), .B(new_n8081), .Y(new_n8202));
  xor_4  g05854(.A(new_n8202), .B(new_n8133), .Y(new_n8203));
  nand_5 g05855(.A(new_n8203), .B(new_n8201), .Y(new_n8204));
  or_5   g05856(.A(new_n8203), .B(new_n8201), .Y(new_n8205));
  nand_5 g05857(.A(new_n8151), .B(new_n8149_1), .Y(new_n8206));
  xor_4  g05858(.A(new_n8206), .B(new_n8183), .Y(new_n8207));
  nand_5 g05859(.A(new_n8089), .B(new_n8088), .Y(new_n8208));
  xor_4  g05860(.A(new_n8208), .B(new_n8131), .Y(new_n8209));
  nand_5 g05861(.A(new_n8209), .B(new_n8207), .Y(new_n8210));
  or_5   g05862(.A(new_n8209), .B(new_n8207), .Y(new_n8211));
  nand_5 g05863(.A(new_n8154), .B(new_n8152), .Y(new_n8212));
  xor_4  g05864(.A(new_n8212), .B(new_n8181), .Y(new_n8213));
  nand_5 g05865(.A(new_n8096), .B(new_n8095_1), .Y(new_n8214));
  xor_4  g05866(.A(new_n8214), .B(new_n8129), .Y(new_n8215_1));
  nand_5 g05867(.A(new_n8215_1), .B(new_n8213), .Y(new_n8216));
  or_5   g05868(.A(new_n8215_1), .B(new_n8213), .Y(new_n8217));
  nand_5 g05869(.A(new_n8157), .B(new_n8155), .Y(new_n8218));
  xor_4  g05870(.A(new_n8218), .B(new_n8179_1), .Y(new_n8219));
  nand_5 g05871(.A(new_n8100), .B(new_n8099), .Y(new_n8220));
  xor_4  g05872(.A(new_n8220), .B(new_n8127_1), .Y(new_n8221));
  nand_5 g05873(.A(new_n8221), .B(new_n8219), .Y(new_n8222));
  or_5   g05874(.A(new_n8221), .B(new_n8219), .Y(new_n8223));
  nand_5 g05875(.A(new_n8160), .B(new_n8158), .Y(new_n8224));
  xor_4  g05876(.A(new_n8224), .B(new_n8177), .Y(new_n8225));
  nand_5 g05877(.A(new_n8104), .B(new_n8103_1), .Y(new_n8226));
  xor_4  g05878(.A(new_n8226), .B(new_n8125), .Y(new_n8227));
  nand_5 g05879(.A(new_n8227), .B(new_n8225), .Y(new_n8228));
  or_5   g05880(.A(new_n8227), .B(new_n8225), .Y(new_n8229));
  nand_5 g05881(.A(new_n8163), .B(new_n8161), .Y(new_n8230));
  xor_4  g05882(.A(new_n8230), .B(new_n8175), .Y(new_n8231));
  nand_5 g05883(.A(new_n8108), .B(new_n8107), .Y(new_n8232));
  xor_4  g05884(.A(new_n8232), .B(new_n8123), .Y(new_n8233));
  nand_5 g05885(.A(new_n8233), .B(new_n8231), .Y(new_n8234));
  or_5   g05886(.A(new_n8233), .B(new_n8231), .Y(new_n8235));
  nand_5 g05887(.A(new_n8166), .B(new_n8164), .Y(new_n8236));
  xor_4  g05888(.A(new_n8236), .B(new_n8173), .Y(new_n8237));
  nand_5 g05889(.A(new_n8112), .B(new_n8111), .Y(new_n8238));
  xor_4  g05890(.A(new_n8238), .B(new_n8121), .Y(new_n8239));
  nand_5 g05891(.A(new_n8239), .B(new_n8237), .Y(new_n8240));
  or_5   g05892(.A(new_n8239), .B(new_n8237), .Y(new_n8241));
  nand_5 g05893(.A(new_n8117), .B(new_n5745), .Y(new_n8242));
  nand_5 g05894(.A(new_n8242), .B(new_n8119), .Y(new_n8243));
  nand_5 g05895(.A(n11479), .B(new_n2377), .Y(new_n8244_1));
  nand_5 g05896(.A(new_n8244_1), .B(new_n8171), .Y(new_n8245));
  nand_5 g05897(.A(new_n8245), .B(new_n8243), .Y(new_n8246));
  not_8  g05898(.A(new_n8171), .Y(new_n8247));
  and_5  g05899(.A(new_n8169), .B(new_n8167), .Y(new_n8248));
  xor_4  g05900(.A(new_n8248), .B(new_n8247), .Y(new_n8249));
  or_5   g05901(.A(new_n8249), .B(new_n8246), .Y(new_n8250));
  nand_5 g05902(.A(new_n8249), .B(new_n8246), .Y(new_n8251));
  nand_5 g05903(.A(new_n8116), .B(new_n8115), .Y(new_n8252));
  xor_4  g05904(.A(new_n8252), .B(new_n8119), .Y(new_n8253));
  not_8  g05905(.A(new_n8253), .Y(new_n8254));
  nand_5 g05906(.A(new_n8254), .B(new_n8251), .Y(new_n8255_1));
  nand_5 g05907(.A(new_n8255_1), .B(new_n8250), .Y(new_n8256_1));
  not_8  g05908(.A(new_n8256_1), .Y(new_n8257));
  nand_5 g05909(.A(new_n8257), .B(new_n8241), .Y(new_n8258));
  nand_5 g05910(.A(new_n8258), .B(new_n8240), .Y(new_n8259_1));
  nand_5 g05911(.A(new_n8259_1), .B(new_n8235), .Y(new_n8260));
  nand_5 g05912(.A(new_n8260), .B(new_n8234), .Y(new_n8261));
  nand_5 g05913(.A(new_n8261), .B(new_n8229), .Y(new_n8262));
  nand_5 g05914(.A(new_n8262), .B(new_n8228), .Y(new_n8263));
  nand_5 g05915(.A(new_n8263), .B(new_n8223), .Y(new_n8264));
  nand_5 g05916(.A(new_n8264), .B(new_n8222), .Y(new_n8265));
  nand_5 g05917(.A(new_n8265), .B(new_n8217), .Y(new_n8266));
  nand_5 g05918(.A(new_n8266), .B(new_n8216), .Y(new_n8267_1));
  nand_5 g05919(.A(new_n8267_1), .B(new_n8211), .Y(new_n8268));
  nand_5 g05920(.A(new_n8268), .B(new_n8210), .Y(new_n8269));
  nand_5 g05921(.A(new_n8269), .B(new_n8205), .Y(new_n8270));
  nand_5 g05922(.A(new_n8270), .B(new_n8204), .Y(new_n8271));
  nand_5 g05923(.A(new_n8271), .B(new_n8199), .Y(new_n8272));
  nand_5 g05924(.A(new_n8272), .B(new_n8198), .Y(new_n8273));
  xor_4  g05925(.A(new_n8273), .B(new_n8193), .Y(n735));
  nand_5 g05926(.A(n21138), .B(n14230), .Y(new_n8275));
  not_8  g05927(.A(n21138), .Y(new_n8276_1));
  nand_5 g05928(.A(new_n8276_1), .B(new_n7513), .Y(new_n8277));
  and_5  g05929(.A(new_n8277), .B(new_n8275), .Y(new_n8278));
  not_8  g05930(.A(new_n8278), .Y(new_n8279));
  nand_5 g05931(.A(new_n7786), .B(n19234), .Y(new_n8280));
  nand_5 g05932(.A(new_n7933), .B(new_n2744), .Y(new_n8281));
  and_5  g05933(.A(new_n8281), .B(new_n8280), .Y(new_n8282));
  nand_5 g05934(.A(new_n8282), .B(n26167), .Y(new_n8283));
  not_8  g05935(.A(n26167), .Y(new_n8284));
  not_8  g05936(.A(new_n8282), .Y(new_n8285_1));
  nand_5 g05937(.A(new_n8285_1), .B(new_n8284), .Y(new_n8286));
  and_5  g05938(.A(new_n8286), .B(new_n8283), .Y(new_n8287));
  or_5   g05939(.A(new_n8287), .B(new_n8279), .Y(new_n8288_1));
  nand_5 g05940(.A(new_n8287), .B(new_n8279), .Y(new_n8289));
  nand_5 g05941(.A(new_n8289), .B(new_n8288_1), .Y(n779));
  not_8  g05942(.A(n17458), .Y(new_n8291));
  nand_5 g05943(.A(new_n8291), .B(n8526), .Y(new_n8292));
  nand_5 g05944(.A(n17458), .B(new_n6846), .Y(new_n8293));
  not_8  g05945(.A(n1222), .Y(new_n8294));
  nand_5 g05946(.A(n2816), .B(new_n8294), .Y(new_n8295));
  nand_5 g05947(.A(new_n6849), .B(n1222), .Y(new_n8296));
  not_8  g05948(.A(n25240), .Y(new_n8297));
  nand_5 g05949(.A(new_n8297), .B(n20359), .Y(new_n8298));
  nand_5 g05950(.A(n25240), .B(new_n6855), .Y(new_n8299));
  not_8  g05951(.A(n10125), .Y(new_n8300));
  nand_5 g05952(.A(new_n8300), .B(n4409), .Y(new_n8301));
  nand_5 g05953(.A(n10125), .B(new_n6861_1), .Y(new_n8302));
  not_8  g05954(.A(n8067), .Y(new_n8303));
  nand_5 g05955(.A(new_n8303), .B(n3570), .Y(new_n8304));
  nand_5 g05956(.A(n8067), .B(new_n6867_1), .Y(new_n8305_1));
  not_8  g05957(.A(n20923), .Y(new_n8306_1));
  nand_5 g05958(.A(new_n8306_1), .B(n13668), .Y(new_n8307));
  nand_5 g05959(.A(n20923), .B(new_n4782), .Y(new_n8308));
  nand_5 g05960(.A(n21276), .B(new_n7606), .Y(new_n8309_1));
  nand_5 g05961(.A(new_n6878), .B(n18157), .Y(new_n8310));
  nand_5 g05962(.A(n26748), .B(new_n7538), .Y(new_n8311));
  nand_5 g05963(.A(new_n6884), .B(n12161), .Y(new_n8312));
  nand_5 g05964(.A(n10057), .B(new_n7519), .Y(new_n8313));
  nand_5 g05965(.A(new_n4654), .B(n5026), .Y(new_n8314));
  nand_5 g05966(.A(new_n4653), .B(n8581), .Y(new_n8315));
  nand_5 g05967(.A(new_n8315), .B(new_n8314), .Y(new_n8316));
  nand_5 g05968(.A(new_n8316), .B(new_n8313), .Y(new_n8317));
  nand_5 g05969(.A(new_n8317), .B(new_n8312), .Y(new_n8318));
  nand_5 g05970(.A(new_n8318), .B(new_n8311), .Y(new_n8319));
  nand_5 g05971(.A(new_n8319), .B(new_n8310), .Y(new_n8320_1));
  nand_5 g05972(.A(new_n8320_1), .B(new_n8309_1), .Y(new_n8321_1));
  nand_5 g05973(.A(new_n8321_1), .B(new_n8308), .Y(new_n8322));
  nand_5 g05974(.A(new_n8322), .B(new_n8307), .Y(new_n8323));
  nand_5 g05975(.A(new_n8323), .B(new_n8305_1), .Y(new_n8324_1));
  nand_5 g05976(.A(new_n8324_1), .B(new_n8304), .Y(new_n8325));
  nand_5 g05977(.A(new_n8325), .B(new_n8302), .Y(new_n8326));
  nand_5 g05978(.A(new_n8326), .B(new_n8301), .Y(new_n8327));
  nand_5 g05979(.A(new_n8327), .B(new_n8299), .Y(new_n8328));
  nand_5 g05980(.A(new_n8328), .B(new_n8298), .Y(new_n8329));
  nand_5 g05981(.A(new_n8329), .B(new_n8296), .Y(new_n8330));
  nand_5 g05982(.A(new_n8330), .B(new_n8295), .Y(new_n8331));
  nand_5 g05983(.A(new_n8331), .B(new_n8293), .Y(new_n8332));
  nand_5 g05984(.A(new_n8332), .B(new_n8292), .Y(new_n8333));
  not_8  g05985(.A(new_n8333), .Y(new_n8334));
  not_8  g05986(.A(n19282), .Y(new_n8335));
  nand_5 g05987(.A(n26986), .B(new_n8335), .Y(new_n8336));
  nand_5 g05988(.A(new_n8140), .B(n19282), .Y(new_n8337));
  nand_5 g05989(.A(n21287), .B(new_n3295), .Y(new_n8338));
  nand_5 g05990(.A(new_n8144), .B(n12657), .Y(new_n8339_1));
  nand_5 g05991(.A(new_n3195), .B(n4256), .Y(new_n8340));
  nand_5 g05992(.A(n17077), .B(new_n8148_1), .Y(new_n8341));
  nand_5 g05993(.A(new_n4283), .B(new_n4280), .Y(new_n8342));
  nand_5 g05994(.A(new_n8342), .B(new_n4282), .Y(new_n8343));
  nand_5 g05995(.A(new_n8343), .B(new_n8341), .Y(new_n8344));
  nand_5 g05996(.A(new_n8344), .B(new_n8340), .Y(new_n8345));
  nand_5 g05997(.A(new_n8345), .B(new_n8339_1), .Y(new_n8346));
  nand_5 g05998(.A(new_n8346), .B(new_n8338), .Y(new_n8347));
  nand_5 g05999(.A(new_n8347), .B(new_n8337), .Y(new_n8348));
  nand_5 g06000(.A(new_n8348), .B(new_n8336), .Y(new_n8349));
  not_8  g06001(.A(new_n8349), .Y(new_n8350));
  nand_5 g06002(.A(new_n8350), .B(new_n8334), .Y(new_n8351));
  nand_5 g06003(.A(new_n8349), .B(new_n8333), .Y(new_n8352));
  nand_5 g06004(.A(new_n8352), .B(new_n8351), .Y(new_n8353));
  not_8  g06005(.A(new_n8353), .Y(new_n8354));
  nand_5 g06006(.A(new_n8293), .B(new_n8292), .Y(new_n8355));
  xor_4  g06007(.A(new_n8355), .B(new_n8331), .Y(new_n8356));
  nand_5 g06008(.A(new_n8337), .B(new_n8336), .Y(new_n8357));
  xor_4  g06009(.A(new_n8357), .B(new_n8347), .Y(new_n8358));
  nand_5 g06010(.A(new_n8358), .B(new_n8356), .Y(new_n8359));
  not_8  g06011(.A(new_n8356), .Y(new_n8360));
  not_8  g06012(.A(new_n8358), .Y(new_n8361));
  nand_5 g06013(.A(new_n8361), .B(new_n8360), .Y(new_n8362));
  nand_5 g06014(.A(new_n8296), .B(new_n8295), .Y(new_n8363_1));
  xor_4  g06015(.A(new_n8363_1), .B(new_n8329), .Y(new_n8364));
  nand_5 g06016(.A(new_n8339_1), .B(new_n8338), .Y(new_n8365));
  xor_4  g06017(.A(new_n8365), .B(new_n8345), .Y(new_n8366));
  nand_5 g06018(.A(new_n8366), .B(new_n8364), .Y(new_n8367));
  or_5   g06019(.A(new_n8366), .B(new_n8364), .Y(new_n8368));
  nand_5 g06020(.A(new_n8299), .B(new_n8298), .Y(new_n8369));
  xor_4  g06021(.A(new_n8369), .B(new_n8327), .Y(new_n8370));
  nand_5 g06022(.A(new_n8341), .B(new_n8340), .Y(new_n8371));
  xor_4  g06023(.A(new_n8371), .B(new_n8343), .Y(new_n8372));
  nand_5 g06024(.A(new_n8372), .B(new_n8370), .Y(new_n8373));
  or_5   g06025(.A(new_n8372), .B(new_n8370), .Y(new_n8374));
  nand_5 g06026(.A(new_n8302), .B(new_n8301), .Y(new_n8375));
  xor_4  g06027(.A(new_n8375), .B(new_n8325), .Y(new_n8376_1));
  not_8  g06028(.A(new_n8376_1), .Y(new_n8377));
  or_5   g06029(.A(new_n8377), .B(new_n4285), .Y(new_n8378));
  nand_5 g06030(.A(new_n8377), .B(new_n4285), .Y(new_n8379));
  nand_5 g06031(.A(new_n8305_1), .B(new_n8304), .Y(new_n8380));
  xor_4  g06032(.A(new_n8380), .B(new_n8323), .Y(new_n8381_1));
  nand_5 g06033(.A(new_n8381_1), .B(new_n4135), .Y(new_n8382));
  not_8  g06034(.A(new_n8381_1), .Y(new_n8383));
  nand_5 g06035(.A(new_n8383), .B(new_n4136), .Y(new_n8384));
  nand_5 g06036(.A(new_n8308), .B(new_n8307), .Y(new_n8385));
  xor_4  g06037(.A(new_n8385), .B(new_n8321_1), .Y(new_n8386));
  nand_5 g06038(.A(new_n8386), .B(new_n4080), .Y(new_n8387));
  not_8  g06039(.A(new_n8386), .Y(new_n8388));
  nand_5 g06040(.A(new_n8388), .B(new_n4081), .Y(new_n8389));
  nand_5 g06041(.A(new_n8310), .B(new_n8309_1), .Y(new_n8390));
  xor_4  g06042(.A(new_n8390), .B(new_n8319), .Y(new_n8391));
  nand_5 g06043(.A(new_n8391), .B(new_n4097), .Y(new_n8392));
  nor_5  g06044(.A(new_n8391), .B(new_n4097), .Y(new_n8393));
  not_8  g06045(.A(new_n8393), .Y(new_n8394));
  nand_5 g06046(.A(new_n8312), .B(new_n8311), .Y(new_n8395));
  xor_4  g06047(.A(new_n8395), .B(new_n8317), .Y(new_n8396));
  nand_5 g06048(.A(new_n8396), .B(new_n4118), .Y(new_n8397));
  not_8  g06049(.A(new_n8396), .Y(new_n8398));
  nand_5 g06050(.A(new_n8398), .B(new_n4119_1), .Y(new_n8399_1));
  and_5  g06051(.A(new_n8314), .B(new_n8313), .Y(new_n8400));
  xor_4  g06052(.A(new_n8400), .B(new_n8315), .Y(new_n8401));
  not_8  g06053(.A(new_n8401), .Y(new_n8402));
  nand_5 g06054(.A(new_n8402), .B(new_n4105), .Y(new_n8403));
  nand_5 g06055(.A(new_n8401), .B(new_n4104), .Y(new_n8404));
  nand_5 g06056(.A(n8920), .B(new_n7526), .Y(new_n8405_1));
  and_5  g06057(.A(new_n8405_1), .B(new_n8315), .Y(new_n8406));
  not_8  g06058(.A(new_n8406), .Y(new_n8407));
  nand_5 g06059(.A(new_n8407), .B(new_n4113), .Y(new_n8408_1));
  nand_5 g06060(.A(new_n8408_1), .B(new_n8404), .Y(new_n8409));
  nand_5 g06061(.A(new_n8409), .B(new_n8403), .Y(new_n8410));
  nand_5 g06062(.A(new_n8410), .B(new_n8399_1), .Y(new_n8411));
  nand_5 g06063(.A(new_n8411), .B(new_n8397), .Y(new_n8412));
  nand_5 g06064(.A(new_n8412), .B(new_n8394), .Y(new_n8413));
  nand_5 g06065(.A(new_n8413), .B(new_n8392), .Y(new_n8414));
  nand_5 g06066(.A(new_n8414), .B(new_n8389), .Y(new_n8415));
  nand_5 g06067(.A(new_n8415), .B(new_n8387), .Y(new_n8416));
  nand_5 g06068(.A(new_n8416), .B(new_n8384), .Y(new_n8417_1));
  nand_5 g06069(.A(new_n8417_1), .B(new_n8382), .Y(new_n8418));
  nand_5 g06070(.A(new_n8418), .B(new_n8379), .Y(new_n8419));
  nand_5 g06071(.A(new_n8419), .B(new_n8378), .Y(new_n8420));
  nand_5 g06072(.A(new_n8420), .B(new_n8374), .Y(new_n8421));
  nand_5 g06073(.A(new_n8421), .B(new_n8373), .Y(new_n8422));
  nand_5 g06074(.A(new_n8422), .B(new_n8368), .Y(new_n8423));
  nand_5 g06075(.A(new_n8423), .B(new_n8367), .Y(new_n8424));
  nand_5 g06076(.A(new_n8424), .B(new_n8362), .Y(new_n8425));
  nand_5 g06077(.A(new_n8425), .B(new_n8359), .Y(new_n8426));
  nor_5  g06078(.A(new_n8426), .B(new_n8354), .Y(new_n8427));
  nand_5 g06079(.A(new_n8426), .B(new_n8354), .Y(new_n8428));
  not_8  g06080(.A(new_n8428), .Y(new_n8429));
  nor_5  g06081(.A(new_n8429), .B(new_n8427), .Y(new_n8430));
  not_8  g06082(.A(n11898), .Y(new_n8431));
  nand_5 g06083(.A(new_n8431), .B(n2979), .Y(new_n8432_1));
  nand_5 g06084(.A(n11898), .B(new_n5369), .Y(new_n8433));
  not_8  g06085(.A(n19941), .Y(new_n8434));
  nand_5 g06086(.A(new_n8434), .B(n647), .Y(new_n8435));
  nand_5 g06087(.A(n19941), .B(new_n5370), .Y(new_n8436));
  not_8  g06088(.A(n1099), .Y(new_n8437));
  nand_5 g06089(.A(n20409), .B(new_n8437), .Y(new_n8438));
  nand_5 g06090(.A(new_n5375), .B(n1099), .Y(new_n8439_1));
  nand_5 g06091(.A(n25749), .B(new_n4298), .Y(new_n8440));
  nand_5 g06092(.A(new_n4293), .B(n2113), .Y(new_n8441));
  not_8  g06093(.A(n21134), .Y(new_n8442));
  nand_5 g06094(.A(new_n8442), .B(n3161), .Y(new_n8443));
  nand_5 g06095(.A(n21134), .B(new_n4219), .Y(new_n8444));
  nand_5 g06096(.A(n9003), .B(new_n4178), .Y(new_n8445));
  nand_5 g06097(.A(new_n5384), .B(n6369), .Y(new_n8446));
  nand_5 g06098(.A(new_n4641), .B(n4957), .Y(new_n8447));
  nand_5 g06099(.A(n25797), .B(new_n4189), .Y(new_n8448));
  nand_5 g06100(.A(new_n4147), .B(n7524), .Y(new_n8449));
  nand_5 g06101(.A(n15967), .B(new_n4195), .Y(new_n8450));
  nand_5 g06102(.A(n15743), .B(new_n4148), .Y(new_n8451));
  nand_5 g06103(.A(new_n4201), .B(n13319), .Y(new_n8452));
  nand_5 g06104(.A(n25435), .B(new_n5469), .Y(new_n8453_1));
  nand_5 g06105(.A(new_n8453_1), .B(new_n8452), .Y(new_n8454));
  nand_5 g06106(.A(new_n8454), .B(new_n8451), .Y(new_n8455));
  nand_5 g06107(.A(new_n8455), .B(new_n8450), .Y(new_n8456));
  nand_5 g06108(.A(new_n8456), .B(new_n8449), .Y(new_n8457));
  nand_5 g06109(.A(new_n8457), .B(new_n8448), .Y(new_n8458));
  nand_5 g06110(.A(new_n8458), .B(new_n8447), .Y(new_n8459));
  nand_5 g06111(.A(new_n8459), .B(new_n8446), .Y(new_n8460));
  nand_5 g06112(.A(new_n8460), .B(new_n8445), .Y(new_n8461));
  nand_5 g06113(.A(new_n8461), .B(new_n8444), .Y(new_n8462));
  nand_5 g06114(.A(new_n8462), .B(new_n8443), .Y(new_n8463));
  nand_5 g06115(.A(new_n8463), .B(new_n8441), .Y(new_n8464));
  nand_5 g06116(.A(new_n8464), .B(new_n8440), .Y(new_n8465));
  nand_5 g06117(.A(new_n8465), .B(new_n8439_1), .Y(new_n8466));
  nand_5 g06118(.A(new_n8466), .B(new_n8438), .Y(new_n8467));
  nand_5 g06119(.A(new_n8467), .B(new_n8436), .Y(new_n8468));
  nand_5 g06120(.A(new_n8468), .B(new_n8435), .Y(new_n8469));
  nand_5 g06121(.A(new_n8469), .B(new_n8433), .Y(new_n8470));
  nand_5 g06122(.A(new_n8470), .B(new_n8432_1), .Y(new_n8471));
  nor_5  g06123(.A(new_n8471), .B(new_n8430), .Y(new_n8472));
  not_8  g06124(.A(new_n8430), .Y(new_n8473));
  not_8  g06125(.A(new_n8471), .Y(new_n8474));
  nor_5  g06126(.A(new_n8474), .B(new_n8473), .Y(new_n8475));
  nor_5  g06127(.A(new_n8475), .B(new_n8472), .Y(new_n8476));
  nand_5 g06128(.A(new_n8359), .B(new_n8362), .Y(new_n8477));
  xor_4  g06129(.A(new_n8477), .B(new_n8424), .Y(new_n8478));
  not_8  g06130(.A(new_n8478), .Y(new_n8479));
  nand_5 g06131(.A(new_n8433), .B(new_n8432_1), .Y(new_n8480_1));
  xor_4  g06132(.A(new_n8480_1), .B(new_n8469), .Y(new_n8481));
  or_5   g06133(.A(new_n8481), .B(new_n8479), .Y(new_n8482));
  nand_5 g06134(.A(new_n8481), .B(new_n8479), .Y(new_n8483));
  nand_5 g06135(.A(new_n8367), .B(new_n8368), .Y(new_n8484));
  xor_4  g06136(.A(new_n8484), .B(new_n8422), .Y(new_n8485));
  not_8  g06137(.A(new_n8485), .Y(new_n8486));
  nand_5 g06138(.A(new_n8436), .B(new_n8435), .Y(new_n8487));
  xor_4  g06139(.A(new_n8487), .B(new_n8467), .Y(new_n8488));
  or_5   g06140(.A(new_n8488), .B(new_n8486), .Y(new_n8489_1));
  nand_5 g06141(.A(new_n8488), .B(new_n8486), .Y(new_n8490));
  nand_5 g06142(.A(new_n8373), .B(new_n8374), .Y(new_n8491));
  xor_4  g06143(.A(new_n8491), .B(new_n8420), .Y(new_n8492));
  not_8  g06144(.A(new_n8492), .Y(new_n8493));
  nand_5 g06145(.A(new_n8439_1), .B(new_n8438), .Y(new_n8494));
  xor_4  g06146(.A(new_n8494), .B(new_n8465), .Y(new_n8495));
  or_5   g06147(.A(new_n8495), .B(new_n8493), .Y(new_n8496));
  nand_5 g06148(.A(new_n8495), .B(new_n8493), .Y(new_n8497));
  nand_5 g06149(.A(new_n8379), .B(new_n8378), .Y(new_n8498));
  xor_4  g06150(.A(new_n8498), .B(new_n8418), .Y(new_n8499));
  not_8  g06151(.A(new_n8499), .Y(new_n8500));
  nand_5 g06152(.A(new_n8441), .B(new_n8440), .Y(new_n8501));
  xor_4  g06153(.A(new_n8501), .B(new_n8463), .Y(new_n8502));
  or_5   g06154(.A(new_n8502), .B(new_n8500), .Y(new_n8503));
  nand_5 g06155(.A(new_n8502), .B(new_n8500), .Y(new_n8504));
  nand_5 g06156(.A(new_n8384), .B(new_n8382), .Y(new_n8505_1));
  xor_4  g06157(.A(new_n8505_1), .B(new_n8416), .Y(new_n8506));
  not_8  g06158(.A(new_n8506), .Y(new_n8507));
  nand_5 g06159(.A(new_n8444), .B(new_n8443), .Y(new_n8508));
  xor_4  g06160(.A(new_n8508), .B(new_n8461), .Y(new_n8509));
  or_5   g06161(.A(new_n8509), .B(new_n8507), .Y(new_n8510_1));
  nand_5 g06162(.A(new_n8509), .B(new_n8507), .Y(new_n8511));
  nand_5 g06163(.A(new_n8389), .B(new_n8387), .Y(new_n8512));
  xor_4  g06164(.A(new_n8512), .B(new_n8414), .Y(new_n8513));
  not_8  g06165(.A(new_n8513), .Y(new_n8514));
  nand_5 g06166(.A(new_n8446), .B(new_n8445), .Y(new_n8515));
  xor_4  g06167(.A(new_n8515), .B(new_n8459), .Y(new_n8516));
  or_5   g06168(.A(new_n8516), .B(new_n8514), .Y(new_n8517));
  nand_5 g06169(.A(new_n8516), .B(new_n8514), .Y(new_n8518));
  nand_5 g06170(.A(new_n8394), .B(new_n8392), .Y(new_n8519_1));
  xor_4  g06171(.A(new_n8519_1), .B(new_n8412), .Y(new_n8520));
  not_8  g06172(.A(new_n8520), .Y(new_n8521));
  nand_5 g06173(.A(new_n8448), .B(new_n8447), .Y(new_n8522));
  xor_4  g06174(.A(new_n8522), .B(new_n8457), .Y(new_n8523));
  or_5   g06175(.A(new_n8523), .B(new_n8521), .Y(new_n8524));
  nand_5 g06176(.A(new_n8523), .B(new_n8521), .Y(new_n8525));
  nand_5 g06177(.A(new_n8399_1), .B(new_n8397), .Y(new_n8526_1));
  xor_4  g06178(.A(new_n8526_1), .B(new_n8410), .Y(new_n8527));
  not_8  g06179(.A(new_n8527), .Y(new_n8528));
  nand_5 g06180(.A(new_n8450), .B(new_n8449), .Y(new_n8529));
  xor_4  g06181(.A(new_n8529), .B(new_n8455), .Y(new_n8530));
  or_5   g06182(.A(new_n8530), .B(new_n8528), .Y(new_n8531));
  nand_5 g06183(.A(new_n8530), .B(new_n8528), .Y(new_n8532));
  not_8  g06184(.A(new_n8408_1), .Y(new_n8533));
  nor_5  g06185(.A(new_n8407), .B(new_n4113), .Y(new_n8534));
  or_5   g06186(.A(new_n8534), .B(new_n8533), .Y(new_n8535_1));
  xor_4  g06187(.A(n25435), .B(new_n5469), .Y(new_n8536));
  nor_5  g06188(.A(new_n8536), .B(new_n8535_1), .Y(new_n8537));
  nand_5 g06189(.A(new_n8452), .B(new_n8451), .Y(new_n8538));
  xnor_4 g06190(.A(new_n8538), .B(new_n8453_1), .Y(new_n8539));
  nand_5 g06191(.A(new_n8539), .B(new_n8537), .Y(new_n8540));
  not_8  g06192(.A(new_n8540), .Y(new_n8541));
  nand_5 g06193(.A(new_n8404), .B(new_n8403), .Y(new_n8542));
  xor_4  g06194(.A(new_n8542), .B(new_n8533), .Y(new_n8543));
  nor_5  g06195(.A(new_n8539), .B(new_n8537), .Y(new_n8544));
  nor_5  g06196(.A(new_n8544), .B(new_n8543), .Y(new_n8545));
  nor_5  g06197(.A(new_n8545), .B(new_n8541), .Y(new_n8546));
  not_8  g06198(.A(new_n8546), .Y(new_n8547));
  nand_5 g06199(.A(new_n8547), .B(new_n8532), .Y(new_n8548));
  nand_5 g06200(.A(new_n8548), .B(new_n8531), .Y(new_n8549));
  nand_5 g06201(.A(new_n8549), .B(new_n8525), .Y(new_n8550_1));
  nand_5 g06202(.A(new_n8550_1), .B(new_n8524), .Y(new_n8551));
  nand_5 g06203(.A(new_n8551), .B(new_n8518), .Y(new_n8552));
  nand_5 g06204(.A(new_n8552), .B(new_n8517), .Y(new_n8553));
  nand_5 g06205(.A(new_n8553), .B(new_n8511), .Y(new_n8554));
  nand_5 g06206(.A(new_n8554), .B(new_n8510_1), .Y(new_n8555));
  nand_5 g06207(.A(new_n8555), .B(new_n8504), .Y(new_n8556));
  nand_5 g06208(.A(new_n8556), .B(new_n8503), .Y(new_n8557));
  nand_5 g06209(.A(new_n8557), .B(new_n8497), .Y(new_n8558));
  nand_5 g06210(.A(new_n8558), .B(new_n8496), .Y(new_n8559));
  nand_5 g06211(.A(new_n8559), .B(new_n8490), .Y(new_n8560));
  nand_5 g06212(.A(new_n8560), .B(new_n8489_1), .Y(new_n8561));
  nand_5 g06213(.A(new_n8561), .B(new_n8483), .Y(new_n8562));
  nand_5 g06214(.A(new_n8562), .B(new_n8482), .Y(new_n8563_1));
  xor_4  g06215(.A(new_n8563_1), .B(new_n8476), .Y(n809));
  not_8  g06216(.A(n1654), .Y(new_n8565));
  nand_5 g06217(.A(new_n8148_1), .B(new_n8565), .Y(new_n8566));
  nand_5 g06218(.A(n4256), .B(n1654), .Y(new_n8567));
  nand_5 g06219(.A(new_n8567), .B(new_n8566), .Y(new_n8568));
  nand_5 g06220(.A(new_n2574), .B(new_n2571), .Y(new_n8569));
  nand_5 g06221(.A(new_n8569), .B(new_n2570_1), .Y(new_n8570));
  not_8  g06222(.A(new_n8570), .Y(new_n8571));
  xor_4  g06223(.A(new_n8571), .B(new_n8568), .Y(new_n8572));
  nand_5 g06224(.A(new_n8572), .B(new_n2577), .Y(new_n8573));
  not_8  g06225(.A(n14440), .Y(new_n8574));
  nand_5 g06226(.A(new_n8144), .B(new_n8574), .Y(new_n8575));
  nand_5 g06227(.A(n21287), .B(n14440), .Y(new_n8576));
  nand_5 g06228(.A(new_n8576), .B(new_n8575), .Y(new_n8577));
  nand_5 g06229(.A(new_n8570), .B(new_n8567), .Y(new_n8578));
  nand_5 g06230(.A(new_n8578), .B(new_n8566), .Y(new_n8579));
  xnor_4 g06231(.A(new_n8579), .B(new_n8577), .Y(new_n8580));
  not_8  g06232(.A(new_n8580), .Y(new_n8581_1));
  nor_5  g06233(.A(new_n8581_1), .B(new_n8573), .Y(new_n8582));
  nand_5 g06234(.A(n26986), .B(n22626), .Y(new_n8583));
  not_8  g06235(.A(n22626), .Y(new_n8584));
  nand_5 g06236(.A(new_n8140), .B(new_n8584), .Y(new_n8585));
  nand_5 g06237(.A(new_n8585), .B(new_n8583), .Y(new_n8586));
  nand_5 g06238(.A(new_n8579), .B(new_n8576), .Y(new_n8587));
  nand_5 g06239(.A(new_n8587), .B(new_n8575), .Y(new_n8588));
  not_8  g06240(.A(new_n8588), .Y(new_n8589));
  xor_4  g06241(.A(new_n8589), .B(new_n8586), .Y(new_n8590));
  nand_5 g06242(.A(new_n8590), .B(new_n8582), .Y(new_n8591));
  nand_5 g06243(.A(new_n8588), .B(new_n8583), .Y(new_n8592));
  nand_5 g06244(.A(new_n8592), .B(new_n8585), .Y(new_n8593));
  not_8  g06245(.A(new_n8593), .Y(new_n8594_1));
  nor_5  g06246(.A(new_n8594_1), .B(new_n8591), .Y(new_n8595));
  xor_4  g06247(.A(new_n8594_1), .B(new_n8591), .Y(new_n8596));
  not_8  g06248(.A(n3425), .Y(new_n8597));
  nand_5 g06249(.A(new_n6233_1), .B(new_n8597), .Y(new_n8598));
  nand_5 g06250(.A(n13494), .B(n3425), .Y(new_n8599));
  nand_5 g06251(.A(new_n6238), .B(new_n3442), .Y(new_n8600));
  nand_5 g06252(.A(n25345), .B(n9967), .Y(new_n8601));
  nand_5 g06253(.A(new_n6062), .B(new_n6242), .Y(new_n8602));
  nand_5 g06254(.A(n20946), .B(n9655), .Y(new_n8603));
  nand_5 g06255(.A(new_n2587), .B(new_n2582_1), .Y(new_n8604));
  nand_5 g06256(.A(new_n8604), .B(new_n2586), .Y(new_n8605));
  nand_5 g06257(.A(new_n8605), .B(new_n8603), .Y(new_n8606));
  nand_5 g06258(.A(new_n8606), .B(new_n8602), .Y(new_n8607));
  nand_5 g06259(.A(new_n8607), .B(new_n8601), .Y(new_n8608_1));
  nand_5 g06260(.A(new_n8608_1), .B(new_n8600), .Y(new_n8609));
  nand_5 g06261(.A(new_n8609), .B(new_n8599), .Y(new_n8610));
  nand_5 g06262(.A(new_n8610), .B(new_n8598), .Y(new_n8611));
  not_8  g06263(.A(new_n8611), .Y(new_n8612));
  or_5   g06264(.A(new_n8612), .B(new_n8596), .Y(new_n8613));
  not_8  g06265(.A(new_n8582), .Y(new_n8614_1));
  not_8  g06266(.A(new_n8590), .Y(new_n8615));
  nand_5 g06267(.A(new_n8615), .B(new_n8614_1), .Y(new_n8616));
  and_5  g06268(.A(new_n8616), .B(new_n8591), .Y(new_n8617));
  nand_5 g06269(.A(new_n8599), .B(new_n8598), .Y(new_n8618));
  xor_4  g06270(.A(new_n8618), .B(new_n8609), .Y(new_n8619));
  nand_5 g06271(.A(new_n8619), .B(new_n8617), .Y(new_n8620_1));
  or_5   g06272(.A(new_n8619), .B(new_n8617), .Y(new_n8621));
  nand_5 g06273(.A(new_n8581_1), .B(new_n8573), .Y(new_n8622));
  and_5  g06274(.A(new_n8622), .B(new_n8614_1), .Y(new_n8623));
  nand_5 g06275(.A(new_n8601), .B(new_n8600), .Y(new_n8624));
  xor_4  g06276(.A(new_n8624), .B(new_n8607), .Y(new_n8625));
  nand_5 g06277(.A(new_n8625), .B(new_n8623), .Y(new_n8626));
  or_5   g06278(.A(new_n8625), .B(new_n8623), .Y(new_n8627));
  not_8  g06279(.A(new_n8572), .Y(new_n8628));
  nand_5 g06280(.A(new_n8628), .B(new_n2578_1), .Y(new_n8629));
  and_5  g06281(.A(new_n8629), .B(new_n8573), .Y(new_n8630));
  nand_5 g06282(.A(new_n8603), .B(new_n8602), .Y(new_n8631));
  xor_4  g06283(.A(new_n8631), .B(new_n8605), .Y(new_n8632));
  nand_5 g06284(.A(new_n8632), .B(new_n8630), .Y(new_n8633));
  or_5   g06285(.A(new_n8632), .B(new_n8630), .Y(new_n8634));
  nand_5 g06286(.A(new_n2592), .B(new_n2567), .Y(new_n8635));
  nand_5 g06287(.A(new_n8635), .B(new_n2591), .Y(new_n8636));
  nand_5 g06288(.A(new_n8636), .B(new_n8634), .Y(new_n8637_1));
  nand_5 g06289(.A(new_n8637_1), .B(new_n8633), .Y(new_n8638_1));
  nand_5 g06290(.A(new_n8638_1), .B(new_n8627), .Y(new_n8639));
  nand_5 g06291(.A(new_n8639), .B(new_n8626), .Y(new_n8640));
  nand_5 g06292(.A(new_n8640), .B(new_n8621), .Y(new_n8641));
  nand_5 g06293(.A(new_n8641), .B(new_n8620_1), .Y(new_n8642));
  nand_5 g06294(.A(new_n8642), .B(new_n8613), .Y(new_n8643));
  nand_5 g06295(.A(new_n8612), .B(new_n8596), .Y(new_n8644));
  nand_5 g06296(.A(new_n8644), .B(new_n8643), .Y(new_n8645));
  nor_5  g06297(.A(new_n8645), .B(new_n8595), .Y(new_n8646));
  nand_5 g06298(.A(new_n8335), .B(n2978), .Y(new_n8647));
  not_8  g06299(.A(n2978), .Y(new_n8648));
  nand_5 g06300(.A(n19282), .B(new_n8648), .Y(new_n8649));
  nand_5 g06301(.A(n23697), .B(new_n3295), .Y(new_n8650));
  nand_5 g06302(.A(new_n7958), .B(n12657), .Y(new_n8651));
  nand_5 g06303(.A(new_n3195), .B(n2289), .Y(new_n8652));
  nand_5 g06304(.A(n17077), .B(new_n7810), .Y(new_n8653));
  nand_5 g06305(.A(new_n3109), .B(n1112), .Y(new_n8654));
  nand_5 g06306(.A(n26510), .B(new_n7757), .Y(new_n8655));
  nand_5 g06307(.A(new_n3073), .B(n20179), .Y(new_n8656_1));
  nand_5 g06308(.A(n23068), .B(new_n7729), .Y(new_n8657));
  nand_5 g06309(.A(new_n3079), .B(n19228), .Y(new_n8658));
  nand_5 g06310(.A(n19514), .B(new_n7732), .Y(new_n8659));
  nand_5 g06311(.A(n15539), .B(new_n3084), .Y(new_n8660));
  nand_5 g06312(.A(new_n7735), .B(n10053), .Y(new_n8661));
  nand_5 g06313(.A(new_n3085), .B(n8052), .Y(new_n8662_1));
  nand_5 g06314(.A(n8399), .B(new_n7738), .Y(new_n8663));
  nand_5 g06315(.A(n10158), .B(new_n3090), .Y(new_n8664));
  nand_5 g06316(.A(new_n7741), .B(n9507), .Y(new_n8665));
  nand_5 g06317(.A(n26979), .B(new_n7784), .Y(new_n8666));
  nand_5 g06318(.A(new_n8666), .B(new_n8665), .Y(new_n8667));
  nand_5 g06319(.A(new_n8667), .B(new_n8664), .Y(new_n8668));
  nand_5 g06320(.A(new_n8668), .B(new_n8663), .Y(new_n8669));
  nand_5 g06321(.A(new_n8669), .B(new_n8662_1), .Y(new_n8670));
  nand_5 g06322(.A(new_n8670), .B(new_n8661), .Y(new_n8671));
  nand_5 g06323(.A(new_n8671), .B(new_n8660), .Y(new_n8672));
  nand_5 g06324(.A(new_n8672), .B(new_n8659), .Y(new_n8673));
  nand_5 g06325(.A(new_n8673), .B(new_n8658), .Y(new_n8674));
  nand_5 g06326(.A(new_n8674), .B(new_n8657), .Y(new_n8675));
  nand_5 g06327(.A(new_n8675), .B(new_n8656_1), .Y(new_n8676));
  nand_5 g06328(.A(new_n8676), .B(new_n8655), .Y(new_n8677));
  nand_5 g06329(.A(new_n8677), .B(new_n8654), .Y(new_n8678_1));
  nand_5 g06330(.A(new_n8678_1), .B(new_n8653), .Y(new_n8679));
  nand_5 g06331(.A(new_n8679), .B(new_n8652), .Y(new_n8680));
  nand_5 g06332(.A(new_n8680), .B(new_n8651), .Y(new_n8681));
  nand_5 g06333(.A(new_n8681), .B(new_n8650), .Y(new_n8682));
  nand_5 g06334(.A(new_n8682), .B(new_n8649), .Y(new_n8683));
  nand_5 g06335(.A(new_n8683), .B(new_n8647), .Y(new_n8684));
  nor_5  g06336(.A(new_n8684), .B(new_n8646), .Y(new_n8685));
  not_8  g06337(.A(new_n8646), .Y(new_n8686));
  not_8  g06338(.A(new_n8684), .Y(new_n8687_1));
  nor_5  g06339(.A(new_n8687_1), .B(new_n8686), .Y(new_n8688));
  nor_5  g06340(.A(new_n8688), .B(new_n8685), .Y(new_n8689));
  nand_5 g06341(.A(new_n8644), .B(new_n8613), .Y(new_n8690));
  xor_4  g06342(.A(new_n8690), .B(new_n8642), .Y(new_n8691));
  nor_5  g06343(.A(new_n8691), .B(new_n8684), .Y(new_n8692));
  not_8  g06344(.A(new_n8691), .Y(new_n8693));
  nor_5  g06345(.A(new_n8693), .B(new_n8687_1), .Y(new_n8694_1));
  nand_5 g06346(.A(new_n8649), .B(new_n8647), .Y(new_n8695));
  xor_4  g06347(.A(new_n8695), .B(new_n8682), .Y(new_n8696));
  nand_5 g06348(.A(new_n8621), .B(new_n8620_1), .Y(new_n8697));
  xor_4  g06349(.A(new_n8697), .B(new_n8640), .Y(new_n8698));
  nand_5 g06350(.A(new_n8698), .B(new_n8696), .Y(new_n8699));
  or_5   g06351(.A(new_n8698), .B(new_n8696), .Y(new_n8700));
  nand_5 g06352(.A(new_n8651), .B(new_n8650), .Y(new_n8701));
  xor_4  g06353(.A(new_n8701), .B(new_n8680), .Y(new_n8702));
  nand_5 g06354(.A(new_n8627), .B(new_n8626), .Y(new_n8703));
  xor_4  g06355(.A(new_n8703), .B(new_n8638_1), .Y(new_n8704));
  nand_5 g06356(.A(new_n8704), .B(new_n8702), .Y(new_n8705));
  or_5   g06357(.A(new_n8704), .B(new_n8702), .Y(new_n8706));
  nand_5 g06358(.A(new_n8653), .B(new_n8652), .Y(new_n8707));
  xor_4  g06359(.A(new_n8707), .B(new_n8678_1), .Y(new_n8708));
  nand_5 g06360(.A(new_n8634), .B(new_n8633), .Y(new_n8709));
  xor_4  g06361(.A(new_n8709), .B(new_n8636), .Y(new_n8710));
  nand_5 g06362(.A(new_n8710), .B(new_n8708), .Y(new_n8711));
  or_5   g06363(.A(new_n8710), .B(new_n8708), .Y(new_n8712));
  nand_5 g06364(.A(new_n8655), .B(new_n8654), .Y(new_n8713));
  xor_4  g06365(.A(new_n8713), .B(new_n8676), .Y(new_n8714));
  nand_5 g06366(.A(new_n8714), .B(new_n2594), .Y(new_n8715));
  or_5   g06367(.A(new_n8714), .B(new_n2594), .Y(new_n8716_1));
  nand_5 g06368(.A(new_n8657), .B(new_n8656_1), .Y(new_n8717));
  xor_4  g06369(.A(new_n8717), .B(new_n8674), .Y(new_n8718));
  nand_5 g06370(.A(new_n8718), .B(new_n2489), .Y(new_n8719));
  or_5   g06371(.A(new_n8718), .B(new_n2489), .Y(new_n8720));
  nand_5 g06372(.A(new_n8659), .B(new_n8658), .Y(new_n8721_1));
  xor_4  g06373(.A(new_n8721_1), .B(new_n8672), .Y(new_n8722));
  nand_5 g06374(.A(new_n8722), .B(new_n2526), .Y(new_n8723));
  or_5   g06375(.A(new_n8722), .B(new_n2526), .Y(new_n8724));
  nand_5 g06376(.A(new_n8661), .B(new_n8660), .Y(new_n8725));
  xor_4  g06377(.A(new_n8725), .B(new_n8670), .Y(new_n8726));
  nand_5 g06378(.A(new_n8726), .B(new_n2532), .Y(new_n8727));
  or_5   g06379(.A(new_n8726), .B(new_n2532), .Y(new_n8728));
  nand_5 g06380(.A(new_n8663), .B(new_n8662_1), .Y(new_n8729));
  xor_4  g06381(.A(new_n8729), .B(new_n8668), .Y(new_n8730));
  nand_5 g06382(.A(new_n8730), .B(new_n2538), .Y(new_n8731));
  or_5   g06383(.A(new_n8730), .B(new_n2538), .Y(new_n8732));
  xor_4  g06384(.A(n26979), .B(new_n7784), .Y(new_n8733));
  nor_5  g06385(.A(new_n8733), .B(new_n2544), .Y(new_n8734));
  and_5  g06386(.A(new_n8665), .B(new_n8664), .Y(new_n8735));
  xor_4  g06387(.A(new_n8735), .B(new_n8666), .Y(new_n8736));
  or_5   g06388(.A(new_n8736), .B(new_n8734), .Y(new_n8737));
  nand_5 g06389(.A(new_n8736), .B(new_n8734), .Y(new_n8738));
  nand_5 g06390(.A(new_n8738), .B(new_n2553_1), .Y(new_n8739));
  nand_5 g06391(.A(new_n8739), .B(new_n8737), .Y(new_n8740));
  nand_5 g06392(.A(new_n8740), .B(new_n8732), .Y(new_n8741));
  nand_5 g06393(.A(new_n8741), .B(new_n8731), .Y(new_n8742));
  nand_5 g06394(.A(new_n8742), .B(new_n8728), .Y(new_n8743));
  nand_5 g06395(.A(new_n8743), .B(new_n8727), .Y(new_n8744_1));
  nand_5 g06396(.A(new_n8744_1), .B(new_n8724), .Y(new_n8745_1));
  nand_5 g06397(.A(new_n8745_1), .B(new_n8723), .Y(new_n8746));
  nand_5 g06398(.A(new_n8746), .B(new_n8720), .Y(new_n8747));
  nand_5 g06399(.A(new_n8747), .B(new_n8719), .Y(new_n8748));
  nand_5 g06400(.A(new_n8748), .B(new_n8716_1), .Y(new_n8749));
  nand_5 g06401(.A(new_n8749), .B(new_n8715), .Y(new_n8750));
  nand_5 g06402(.A(new_n8750), .B(new_n8712), .Y(new_n8751));
  nand_5 g06403(.A(new_n8751), .B(new_n8711), .Y(new_n8752));
  nand_5 g06404(.A(new_n8752), .B(new_n8706), .Y(new_n8753));
  nand_5 g06405(.A(new_n8753), .B(new_n8705), .Y(new_n8754));
  nand_5 g06406(.A(new_n8754), .B(new_n8700), .Y(new_n8755));
  nand_5 g06407(.A(new_n8755), .B(new_n8699), .Y(new_n8756));
  nor_5  g06408(.A(new_n8756), .B(new_n8694_1), .Y(new_n8757));
  nor_5  g06409(.A(new_n8757), .B(new_n8692), .Y(new_n8758));
  xor_4  g06410(.A(new_n8758), .B(new_n8689), .Y(n819));
  nand_5 g06411(.A(new_n8584), .B(n8856), .Y(new_n8760));
  nand_5 g06412(.A(n22626), .B(new_n7991), .Y(new_n8761));
  nand_5 g06413(.A(new_n8574), .B(n14130), .Y(new_n8762));
  nand_5 g06414(.A(n14440), .B(new_n3849), .Y(new_n8763));
  nand_5 g06415(.A(n16482), .B(new_n8565), .Y(new_n8764));
  nand_5 g06416(.A(new_n7998), .B(n1654), .Y(new_n8765));
  nand_5 g06417(.A(new_n2568), .B(n9942), .Y(new_n8766));
  nand_5 g06418(.A(n13783), .B(new_n2599), .Y(new_n8767));
  nand_5 g06419(.A(new_n2475), .B(n25643), .Y(new_n8768));
  nand_5 g06420(.A(n26660), .B(new_n2516), .Y(new_n8769));
  nand_5 g06421(.A(n9557), .B(new_n2412), .Y(new_n8770));
  nand_5 g06422(.A(new_n2490), .B(n3018), .Y(new_n8771));
  nand_5 g06423(.A(new_n2401), .B(n3136), .Y(new_n8772));
  nand_5 g06424(.A(n3480), .B(new_n2494), .Y(new_n8773));
  nand_5 g06425(.A(new_n2394), .B(n6385), .Y(new_n8774));
  nand_5 g06426(.A(n16722), .B(new_n2498), .Y(new_n8775));
  nand_5 g06427(.A(n20138), .B(new_n2383), .Y(new_n8776));
  nand_5 g06428(.A(new_n2502), .B(n11486), .Y(new_n8777));
  nand_5 g06429(.A(n13781), .B(new_n3850_1), .Y(new_n8778));
  nand_5 g06430(.A(new_n8778), .B(new_n8777), .Y(new_n8779));
  nand_5 g06431(.A(new_n8779), .B(new_n8776), .Y(new_n8780));
  nand_5 g06432(.A(new_n8780), .B(new_n8775), .Y(new_n8781));
  nand_5 g06433(.A(new_n8781), .B(new_n8774), .Y(new_n8782_1));
  nand_5 g06434(.A(new_n8782_1), .B(new_n8773), .Y(new_n8783));
  nand_5 g06435(.A(new_n8783), .B(new_n8772), .Y(new_n8784));
  nand_5 g06436(.A(new_n8784), .B(new_n8771), .Y(new_n8785));
  nand_5 g06437(.A(new_n8785), .B(new_n8770), .Y(new_n8786));
  nand_5 g06438(.A(new_n8786), .B(new_n8769), .Y(new_n8787));
  nand_5 g06439(.A(new_n8787), .B(new_n8768), .Y(new_n8788));
  nand_5 g06440(.A(new_n8788), .B(new_n8767), .Y(new_n8789));
  nand_5 g06441(.A(new_n8789), .B(new_n8766), .Y(new_n8790));
  nand_5 g06442(.A(new_n8790), .B(new_n8765), .Y(new_n8791));
  nand_5 g06443(.A(new_n8791), .B(new_n8764), .Y(new_n8792));
  nand_5 g06444(.A(new_n8792), .B(new_n8763), .Y(new_n8793));
  nand_5 g06445(.A(new_n8793), .B(new_n8762), .Y(new_n8794));
  nand_5 g06446(.A(new_n8794), .B(new_n8761), .Y(new_n8795));
  nand_5 g06447(.A(new_n8795), .B(new_n8760), .Y(new_n8796));
  not_8  g06448(.A(new_n8796), .Y(new_n8797));
  not_8  g06449(.A(n25120), .Y(new_n8798));
  nand_5 g06450(.A(new_n8798), .B(n3582), .Y(new_n8799));
  nand_5 g06451(.A(n25120), .B(new_n6795), .Y(new_n8800));
  not_8  g06452(.A(n8363), .Y(new_n8801));
  nand_5 g06453(.A(new_n8801), .B(n2145), .Y(new_n8802));
  nand_5 g06454(.A(n8363), .B(new_n6799), .Y(new_n8803_1));
  not_8  g06455(.A(n14680), .Y(new_n8804));
  nand_5 g06456(.A(new_n8804), .B(n5031), .Y(new_n8805));
  nand_5 g06457(.A(n14680), .B(new_n6803), .Y(new_n8806_1));
  not_8  g06458(.A(n17250), .Y(new_n8807));
  nand_5 g06459(.A(new_n8807), .B(n11044), .Y(new_n8808));
  nand_5 g06460(.A(n17250), .B(new_n6808), .Y(new_n8809_1));
  not_8  g06461(.A(n23160), .Y(new_n8810));
  nand_5 g06462(.A(new_n8810), .B(n2421), .Y(new_n8811));
  nand_5 g06463(.A(n23160), .B(new_n6811), .Y(new_n8812));
  not_8  g06464(.A(n16524), .Y(new_n8813));
  nand_5 g06465(.A(new_n8813), .B(n987), .Y(new_n8814));
  nand_5 g06466(.A(n16524), .B(new_n6814_1), .Y(new_n8815));
  nand_5 g06467(.A(n20478), .B(new_n7605), .Y(new_n8816));
  nand_5 g06468(.A(new_n6817), .B(n11056), .Y(new_n8817));
  nand_5 g06469(.A(n26882), .B(new_n7539), .Y(new_n8818));
  nand_5 g06470(.A(new_n6820), .B(n15271), .Y(new_n8819));
  nand_5 g06471(.A(new_n6544), .B(n22619), .Y(new_n8820));
  nand_5 g06472(.A(n25877), .B(new_n6823), .Y(new_n8821_1));
  nand_5 g06473(.A(n24323), .B(new_n6561), .Y(new_n8822));
  nand_5 g06474(.A(new_n8822), .B(new_n8821_1), .Y(new_n8823));
  nand_5 g06475(.A(new_n8823), .B(new_n8820), .Y(new_n8824_1));
  nand_5 g06476(.A(new_n8824_1), .B(new_n8819), .Y(new_n8825));
  nand_5 g06477(.A(new_n8825), .B(new_n8818), .Y(new_n8826));
  nand_5 g06478(.A(new_n8826), .B(new_n8817), .Y(new_n8827_1));
  nand_5 g06479(.A(new_n8827_1), .B(new_n8816), .Y(new_n8828));
  nand_5 g06480(.A(new_n8828), .B(new_n8815), .Y(new_n8829));
  nand_5 g06481(.A(new_n8829), .B(new_n8814), .Y(new_n8830));
  nand_5 g06482(.A(new_n8830), .B(new_n8812), .Y(new_n8831));
  nand_5 g06483(.A(new_n8831), .B(new_n8811), .Y(new_n8832));
  nand_5 g06484(.A(new_n8832), .B(new_n8809_1), .Y(new_n8833));
  nand_5 g06485(.A(new_n8833), .B(new_n8808), .Y(new_n8834));
  nand_5 g06486(.A(new_n8834), .B(new_n8806_1), .Y(new_n8835));
  nand_5 g06487(.A(new_n8835), .B(new_n8805), .Y(new_n8836));
  nand_5 g06488(.A(new_n8836), .B(new_n8803_1), .Y(new_n8837));
  nand_5 g06489(.A(new_n8837), .B(new_n8802), .Y(new_n8838));
  nand_5 g06490(.A(new_n8838), .B(new_n8800), .Y(new_n8839));
  nand_5 g06491(.A(new_n8839), .B(new_n8799), .Y(new_n8840));
  not_8  g06492(.A(new_n8840), .Y(new_n8841));
  nand_5 g06493(.A(new_n8841), .B(new_n8797), .Y(new_n8842));
  nand_5 g06494(.A(new_n8840), .B(new_n8796), .Y(new_n8843));
  nand_5 g06495(.A(new_n8843), .B(new_n8842), .Y(new_n8844));
  not_8  g06496(.A(new_n8844), .Y(new_n8845));
  nand_5 g06497(.A(new_n8800), .B(new_n8799), .Y(new_n8846));
  xor_4  g06498(.A(new_n8846), .B(new_n8838), .Y(new_n8847));
  nand_5 g06499(.A(new_n8761), .B(new_n8760), .Y(new_n8848));
  xor_4  g06500(.A(new_n8848), .B(new_n8794), .Y(new_n8849_1));
  nand_5 g06501(.A(new_n8849_1), .B(new_n8847), .Y(new_n8850));
  or_5   g06502(.A(new_n8849_1), .B(new_n8847), .Y(new_n8851));
  nand_5 g06503(.A(new_n8803_1), .B(new_n8802), .Y(new_n8852));
  xor_4  g06504(.A(new_n8852), .B(new_n8836), .Y(new_n8853));
  nand_5 g06505(.A(new_n8763), .B(new_n8762), .Y(new_n8854));
  xor_4  g06506(.A(new_n8854), .B(new_n8792), .Y(new_n8855));
  nand_5 g06507(.A(new_n8855), .B(new_n8853), .Y(new_n8856_1));
  not_8  g06508(.A(new_n8853), .Y(new_n8857));
  not_8  g06509(.A(new_n8855), .Y(new_n8858));
  nand_5 g06510(.A(new_n8858), .B(new_n8857), .Y(new_n8859));
  nand_5 g06511(.A(new_n8806_1), .B(new_n8805), .Y(new_n8860));
  xor_4  g06512(.A(new_n8860), .B(new_n8834), .Y(new_n8861_1));
  nand_5 g06513(.A(new_n8765), .B(new_n8764), .Y(new_n8862_1));
  xor_4  g06514(.A(new_n8862_1), .B(new_n8790), .Y(new_n8863));
  nand_5 g06515(.A(new_n8863), .B(new_n8861_1), .Y(new_n8864));
  not_8  g06516(.A(new_n8861_1), .Y(new_n8865));
  not_8  g06517(.A(new_n8863), .Y(new_n8866));
  nand_5 g06518(.A(new_n8866), .B(new_n8865), .Y(new_n8867));
  nand_5 g06519(.A(new_n8809_1), .B(new_n8808), .Y(new_n8868));
  xor_4  g06520(.A(new_n8868), .B(new_n8832), .Y(new_n8869_1));
  nand_5 g06521(.A(new_n8767), .B(new_n8766), .Y(new_n8870));
  xor_4  g06522(.A(new_n8870), .B(new_n8788), .Y(new_n8871));
  nand_5 g06523(.A(new_n8871), .B(new_n8869_1), .Y(new_n8872));
  not_8  g06524(.A(new_n8869_1), .Y(new_n8873));
  not_8  g06525(.A(new_n8871), .Y(new_n8874));
  nand_5 g06526(.A(new_n8874), .B(new_n8873), .Y(new_n8875));
  nand_5 g06527(.A(new_n8812), .B(new_n8811), .Y(new_n8876));
  xor_4  g06528(.A(new_n8876), .B(new_n8830), .Y(new_n8877));
  nand_5 g06529(.A(new_n8769), .B(new_n8768), .Y(new_n8878));
  xor_4  g06530(.A(new_n8878), .B(new_n8786), .Y(new_n8879));
  nand_5 g06531(.A(new_n8879), .B(new_n8877), .Y(new_n8880));
  not_8  g06532(.A(new_n8877), .Y(new_n8881));
  not_8  g06533(.A(new_n8879), .Y(new_n8882));
  nand_5 g06534(.A(new_n8882), .B(new_n8881), .Y(new_n8883));
  nand_5 g06535(.A(new_n8815), .B(new_n8814), .Y(new_n8884_1));
  xor_4  g06536(.A(new_n8884_1), .B(new_n8828), .Y(new_n8885));
  nand_5 g06537(.A(new_n8771), .B(new_n8770), .Y(new_n8886));
  xor_4  g06538(.A(new_n8886), .B(new_n8784), .Y(new_n8887));
  nand_5 g06539(.A(new_n8887), .B(new_n8885), .Y(new_n8888));
  not_8  g06540(.A(new_n8885), .Y(new_n8889));
  not_8  g06541(.A(new_n8887), .Y(new_n8890));
  nand_5 g06542(.A(new_n8890), .B(new_n8889), .Y(new_n8891));
  nand_5 g06543(.A(new_n8817), .B(new_n8816), .Y(new_n8892));
  xor_4  g06544(.A(new_n8892), .B(new_n8826), .Y(new_n8893));
  nand_5 g06545(.A(new_n8773), .B(new_n8772), .Y(new_n8894));
  xor_4  g06546(.A(new_n8894), .B(new_n8782_1), .Y(new_n8895));
  nand_5 g06547(.A(new_n8895), .B(new_n8893), .Y(new_n8896));
  not_8  g06548(.A(new_n8893), .Y(new_n8897));
  not_8  g06549(.A(new_n8895), .Y(new_n8898));
  nand_5 g06550(.A(new_n8898), .B(new_n8897), .Y(new_n8899));
  nand_5 g06551(.A(new_n8819), .B(new_n8818), .Y(new_n8900));
  xor_4  g06552(.A(new_n8900), .B(new_n8824_1), .Y(new_n8901));
  nand_5 g06553(.A(new_n8775), .B(new_n8774), .Y(new_n8902));
  xor_4  g06554(.A(new_n8902), .B(new_n8780), .Y(new_n8903));
  nand_5 g06555(.A(new_n8903), .B(new_n8901), .Y(new_n8904));
  not_8  g06556(.A(new_n8901), .Y(new_n8905));
  not_8  g06557(.A(new_n8903), .Y(new_n8906));
  nand_5 g06558(.A(new_n8906), .B(new_n8905), .Y(new_n8907));
  and_5  g06559(.A(new_n8821_1), .B(new_n8820), .Y(new_n8908));
  xor_4  g06560(.A(new_n8908), .B(new_n8822), .Y(new_n8909_1));
  not_8  g06561(.A(new_n8909_1), .Y(new_n8910));
  and_5  g06562(.A(new_n8777), .B(new_n8776), .Y(new_n8911_1));
  xor_4  g06563(.A(new_n8911_1), .B(new_n8778), .Y(new_n8912));
  not_8  g06564(.A(new_n8912), .Y(new_n8913));
  nand_5 g06565(.A(new_n8913), .B(new_n8910), .Y(new_n8914));
  nand_5 g06566(.A(new_n8912), .B(new_n8909_1), .Y(new_n8915));
  nand_5 g06567(.A(new_n6537), .B(n6775), .Y(new_n8916));
  nand_5 g06568(.A(new_n8916), .B(new_n8822), .Y(new_n8917));
  nand_5 g06569(.A(new_n2378), .B(n9251), .Y(new_n8918));
  nand_5 g06570(.A(new_n8918), .B(new_n8778), .Y(new_n8919));
  nand_5 g06571(.A(new_n8919), .B(new_n8917), .Y(new_n8920_1));
  nand_5 g06572(.A(new_n8920_1), .B(new_n8915), .Y(new_n8921));
  nand_5 g06573(.A(new_n8921), .B(new_n8914), .Y(new_n8922));
  nand_5 g06574(.A(new_n8922), .B(new_n8907), .Y(new_n8923));
  nand_5 g06575(.A(new_n8923), .B(new_n8904), .Y(new_n8924));
  nand_5 g06576(.A(new_n8924), .B(new_n8899), .Y(new_n8925));
  nand_5 g06577(.A(new_n8925), .B(new_n8896), .Y(new_n8926));
  nand_5 g06578(.A(new_n8926), .B(new_n8891), .Y(new_n8927));
  nand_5 g06579(.A(new_n8927), .B(new_n8888), .Y(new_n8928));
  nand_5 g06580(.A(new_n8928), .B(new_n8883), .Y(new_n8929));
  nand_5 g06581(.A(new_n8929), .B(new_n8880), .Y(new_n8930));
  nand_5 g06582(.A(new_n8930), .B(new_n8875), .Y(new_n8931));
  nand_5 g06583(.A(new_n8931), .B(new_n8872), .Y(new_n8932));
  nand_5 g06584(.A(new_n8932), .B(new_n8867), .Y(new_n8933));
  nand_5 g06585(.A(new_n8933), .B(new_n8864), .Y(new_n8934));
  nand_5 g06586(.A(new_n8934), .B(new_n8859), .Y(new_n8935));
  nand_5 g06587(.A(new_n8935), .B(new_n8856_1), .Y(new_n8936));
  nand_5 g06588(.A(new_n8936), .B(new_n8851), .Y(new_n8937));
  nand_5 g06589(.A(new_n8937), .B(new_n8850), .Y(new_n8938));
  nor_5  g06590(.A(new_n8938), .B(new_n8845), .Y(new_n8939));
  nand_5 g06591(.A(new_n8938), .B(new_n8845), .Y(new_n8940));
  not_8  g06592(.A(new_n8940), .Y(new_n8941));
  nor_5  g06593(.A(new_n8941), .B(new_n8939), .Y(new_n8942));
  not_8  g06594(.A(new_n8942), .Y(new_n8943_1));
  nand_5 g06595(.A(new_n5468), .B(new_n5394), .Y(new_n8944));
  or_5   g06596(.A(new_n8944), .B(n19680), .Y(new_n8945));
  nor_5  g06597(.A(new_n8945), .B(n7421), .Y(new_n8946));
  nand_5 g06598(.A(new_n8946), .B(new_n5385), .Y(new_n8947));
  nor_5  g06599(.A(new_n8947), .B(n11630), .Y(new_n8948));
  nand_5 g06600(.A(new_n8948), .B(new_n5378), .Y(new_n8949));
  nor_5  g06601(.A(new_n8949), .B(n18227), .Y(new_n8950));
  nand_5 g06602(.A(new_n8950), .B(new_n5371), .Y(new_n8951));
  nor_5  g06603(.A(new_n8951), .B(n9554), .Y(new_n8952));
  not_8  g06604(.A(new_n8952), .Y(new_n8953));
  nand_5 g06605(.A(new_n8951), .B(n9554), .Y(new_n8954));
  nand_5 g06606(.A(new_n8954), .B(new_n8953), .Y(new_n8955));
  nand_5 g06607(.A(new_n8955), .B(new_n5419), .Y(new_n8956));
  not_8  g06608(.A(new_n8956), .Y(new_n8957));
  xor_4  g06609(.A(new_n8950), .B(n26408), .Y(new_n8958));
  nand_5 g06610(.A(new_n8958), .B(new_n3694), .Y(new_n8959));
  nor_5  g06611(.A(new_n8958), .B(new_n3694), .Y(new_n8960));
  not_8  g06612(.A(new_n8960), .Y(new_n8961));
  xor_4  g06613(.A(new_n8949), .B(new_n5374), .Y(new_n8962));
  nand_5 g06614(.A(new_n8962), .B(new_n3778), .Y(new_n8963));
  nor_5  g06615(.A(new_n8962), .B(new_n3778), .Y(new_n8964_1));
  not_8  g06616(.A(new_n8964_1), .Y(new_n8965));
  xor_4  g06617(.A(new_n8948), .B(n7377), .Y(new_n8966));
  nand_5 g06618(.A(new_n8966), .B(new_n3695), .Y(new_n8967));
  nor_5  g06619(.A(new_n8966), .B(new_n3695), .Y(new_n8968));
  not_8  g06620(.A(new_n8968), .Y(new_n8969));
  xor_4  g06621(.A(new_n8947), .B(new_n5381), .Y(new_n8970));
  nand_5 g06622(.A(new_n8970), .B(new_n3793), .Y(new_n8971_1));
  nor_5  g06623(.A(new_n8970), .B(new_n3793), .Y(new_n8972));
  not_8  g06624(.A(new_n8972), .Y(new_n8973));
  xor_4  g06625(.A(new_n8946), .B(new_n5385), .Y(new_n8974));
  or_5   g06626(.A(new_n8974), .B(n9598), .Y(new_n8975));
  nand_5 g06627(.A(new_n8974), .B(n9598), .Y(new_n8976));
  xor_4  g06628(.A(new_n8945), .B(n7421), .Y(new_n8977));
  or_5   g06629(.A(new_n8977), .B(n22290), .Y(new_n8978));
  nand_5 g06630(.A(new_n8977), .B(n22290), .Y(new_n8979));
  nand_5 g06631(.A(new_n8944), .B(n19680), .Y(new_n8980));
  and_5  g06632(.A(new_n8980), .B(new_n8945), .Y(new_n8981));
  or_5   g06633(.A(new_n8981), .B(n11273), .Y(new_n8982_1));
  nand_5 g06634(.A(new_n8981), .B(n11273), .Y(new_n8983));
  nand_5 g06635(.A(n15508), .B(n2809), .Y(new_n8984));
  and_5  g06636(.A(new_n8984), .B(new_n8944), .Y(new_n8985));
  or_5   g06637(.A(new_n8985), .B(n25565), .Y(new_n8986));
  nand_5 g06638(.A(new_n8985), .B(n25565), .Y(new_n8987));
  nand_5 g06639(.A(n21993), .B(n15508), .Y(new_n8988));
  nand_5 g06640(.A(new_n8988), .B(new_n8987), .Y(new_n8989));
  nand_5 g06641(.A(new_n8989), .B(new_n8986), .Y(new_n8990));
  nand_5 g06642(.A(new_n8990), .B(new_n8983), .Y(new_n8991));
  nand_5 g06643(.A(new_n8991), .B(new_n8982_1), .Y(new_n8992));
  nand_5 g06644(.A(new_n8992), .B(new_n8979), .Y(new_n8993_1));
  nand_5 g06645(.A(new_n8993_1), .B(new_n8978), .Y(new_n8994));
  nand_5 g06646(.A(new_n8994), .B(new_n8976), .Y(new_n8995));
  nand_5 g06647(.A(new_n8995), .B(new_n8975), .Y(new_n8996));
  nand_5 g06648(.A(new_n8996), .B(new_n8973), .Y(new_n8997));
  nand_5 g06649(.A(new_n8997), .B(new_n8971_1), .Y(new_n8998));
  nand_5 g06650(.A(new_n8998), .B(new_n8969), .Y(new_n8999));
  nand_5 g06651(.A(new_n8999), .B(new_n8967), .Y(new_n9000));
  nand_5 g06652(.A(new_n9000), .B(new_n8965), .Y(new_n9001));
  nand_5 g06653(.A(new_n9001), .B(new_n8963), .Y(new_n9002));
  nand_5 g06654(.A(new_n9002), .B(new_n8961), .Y(new_n9003_1));
  nand_5 g06655(.A(new_n9003_1), .B(new_n8959), .Y(new_n9004));
  nor_5  g06656(.A(new_n9004), .B(new_n8957), .Y(new_n9005));
  nor_5  g06657(.A(new_n8955), .B(new_n5419), .Y(new_n9006));
  not_8  g06658(.A(new_n9006), .Y(new_n9007));
  nand_5 g06659(.A(new_n9007), .B(new_n8953), .Y(new_n9008));
  nor_5  g06660(.A(new_n9008), .B(new_n9005), .Y(new_n9009));
  nand_5 g06661(.A(new_n9009), .B(new_n8943_1), .Y(new_n9010));
  not_8  g06662(.A(new_n9009), .Y(new_n9011));
  nand_5 g06663(.A(new_n9011), .B(new_n8942), .Y(new_n9012_1));
  nand_5 g06664(.A(new_n9012_1), .B(new_n9010), .Y(new_n9013));
  nand_5 g06665(.A(new_n8851), .B(new_n8850), .Y(new_n9014));
  xor_4  g06666(.A(new_n9014), .B(new_n8936), .Y(new_n9015));
  not_8  g06667(.A(new_n9015), .Y(new_n9016));
  nand_5 g06668(.A(new_n9007), .B(new_n8956), .Y(new_n9017));
  xor_4  g06669(.A(new_n9017), .B(new_n9004), .Y(new_n9018));
  not_8  g06670(.A(new_n9018), .Y(new_n9019));
  nand_5 g06671(.A(new_n9019), .B(new_n9016), .Y(new_n9020));
  nand_5 g06672(.A(new_n9018), .B(new_n9015), .Y(new_n9021));
  nand_5 g06673(.A(new_n8859), .B(new_n8856_1), .Y(new_n9022));
  xor_4  g06674(.A(new_n9022), .B(new_n8934), .Y(new_n9023));
  nand_5 g06675(.A(new_n8961), .B(new_n8959), .Y(new_n9024));
  xor_4  g06676(.A(new_n9024), .B(new_n9002), .Y(new_n9025));
  or_5   g06677(.A(new_n9025), .B(new_n9023), .Y(new_n9026));
  nand_5 g06678(.A(new_n9025), .B(new_n9023), .Y(new_n9027));
  nand_5 g06679(.A(new_n8867), .B(new_n8864), .Y(new_n9028));
  xor_4  g06680(.A(new_n9028), .B(new_n8932), .Y(new_n9029));
  nand_5 g06681(.A(new_n8965), .B(new_n8963), .Y(new_n9030));
  xor_4  g06682(.A(new_n9030), .B(new_n9000), .Y(new_n9031));
  or_5   g06683(.A(new_n9031), .B(new_n9029), .Y(new_n9032_1));
  nand_5 g06684(.A(new_n9031), .B(new_n9029), .Y(new_n9033));
  nand_5 g06685(.A(new_n8875), .B(new_n8872), .Y(new_n9034));
  xor_4  g06686(.A(new_n9034), .B(new_n8930), .Y(new_n9035));
  not_8  g06687(.A(new_n9035), .Y(new_n9036));
  nand_5 g06688(.A(new_n8969), .B(new_n8967), .Y(new_n9037));
  xor_4  g06689(.A(new_n9037), .B(new_n8998), .Y(new_n9038));
  not_8  g06690(.A(new_n9038), .Y(new_n9039));
  nand_5 g06691(.A(new_n9039), .B(new_n9036), .Y(new_n9040));
  nand_5 g06692(.A(new_n9038), .B(new_n9035), .Y(new_n9041));
  nand_5 g06693(.A(new_n8883), .B(new_n8880), .Y(new_n9042_1));
  xor_4  g06694(.A(new_n9042_1), .B(new_n8928), .Y(new_n9043));
  not_8  g06695(.A(new_n9043), .Y(new_n9044));
  nand_5 g06696(.A(new_n8973), .B(new_n8971_1), .Y(new_n9045));
  xor_4  g06697(.A(new_n9045), .B(new_n8996), .Y(new_n9046_1));
  not_8  g06698(.A(new_n9046_1), .Y(new_n9047_1));
  nand_5 g06699(.A(new_n9047_1), .B(new_n9044), .Y(new_n9048));
  nand_5 g06700(.A(new_n9046_1), .B(new_n9043), .Y(new_n9049));
  nand_5 g06701(.A(new_n8891), .B(new_n8888), .Y(new_n9050));
  xor_4  g06702(.A(new_n9050), .B(new_n8926), .Y(new_n9051));
  not_8  g06703(.A(new_n9051), .Y(new_n9052));
  nand_5 g06704(.A(new_n8976), .B(new_n8975), .Y(new_n9053));
  xor_4  g06705(.A(new_n9053), .B(new_n8994), .Y(new_n9054));
  not_8  g06706(.A(new_n9054), .Y(new_n9055));
  nand_5 g06707(.A(new_n9055), .B(new_n9052), .Y(new_n9056));
  nand_5 g06708(.A(new_n9054), .B(new_n9051), .Y(new_n9057));
  nand_5 g06709(.A(new_n8899), .B(new_n8896), .Y(new_n9058));
  xor_4  g06710(.A(new_n9058), .B(new_n8924), .Y(new_n9059));
  not_8  g06711(.A(new_n9059), .Y(new_n9060));
  nand_5 g06712(.A(new_n8979), .B(new_n8978), .Y(new_n9061));
  xor_4  g06713(.A(new_n9061), .B(new_n8992), .Y(new_n9062));
  not_8  g06714(.A(new_n9062), .Y(new_n9063));
  nand_5 g06715(.A(new_n9063), .B(new_n9060), .Y(new_n9064));
  nand_5 g06716(.A(new_n9062), .B(new_n9059), .Y(new_n9065));
  nand_5 g06717(.A(new_n8907), .B(new_n8904), .Y(new_n9066));
  xor_4  g06718(.A(new_n9066), .B(new_n8922), .Y(new_n9067));
  xor_4  g06719(.A(new_n8919), .B(new_n8917), .Y(new_n9068));
  nand_5 g06720(.A(new_n3697), .B(new_n5468), .Y(new_n9069));
  nand_5 g06721(.A(new_n9069), .B(new_n8988), .Y(new_n9070));
  not_8  g06722(.A(new_n9070), .Y(new_n9071));
  nand_5 g06723(.A(new_n9071), .B(new_n9068), .Y(new_n9072));
  not_8  g06724(.A(new_n9072), .Y(new_n9073));
  and_5  g06725(.A(new_n8987), .B(new_n8986), .Y(new_n9074));
  nand_5 g06726(.A(new_n9074), .B(new_n9073), .Y(new_n9075));
  xor_4  g06727(.A(new_n9074), .B(new_n8988), .Y(new_n9076));
  nand_5 g06728(.A(new_n9076), .B(new_n9072), .Y(new_n9077));
  nand_5 g06729(.A(new_n8915), .B(new_n8914), .Y(new_n9078));
  xor_4  g06730(.A(new_n9078), .B(new_n8920_1), .Y(new_n9079));
  nand_5 g06731(.A(new_n9079), .B(new_n9077), .Y(new_n9080));
  nand_5 g06732(.A(new_n9080), .B(new_n9075), .Y(new_n9081));
  or_5   g06733(.A(new_n9081), .B(new_n9067), .Y(new_n9082));
  nand_5 g06734(.A(new_n9081), .B(new_n9067), .Y(new_n9083));
  nand_5 g06735(.A(new_n8983), .B(new_n8982_1), .Y(new_n9084));
  xor_4  g06736(.A(new_n9084), .B(new_n8990), .Y(new_n9085));
  not_8  g06737(.A(new_n9085), .Y(new_n9086));
  nand_5 g06738(.A(new_n9086), .B(new_n9083), .Y(new_n9087));
  nand_5 g06739(.A(new_n9087), .B(new_n9082), .Y(new_n9088));
  nand_5 g06740(.A(new_n9088), .B(new_n9065), .Y(new_n9089));
  nand_5 g06741(.A(new_n9089), .B(new_n9064), .Y(new_n9090_1));
  nand_5 g06742(.A(new_n9090_1), .B(new_n9057), .Y(new_n9091));
  nand_5 g06743(.A(new_n9091), .B(new_n9056), .Y(new_n9092));
  nand_5 g06744(.A(new_n9092), .B(new_n9049), .Y(new_n9093));
  nand_5 g06745(.A(new_n9093), .B(new_n9048), .Y(new_n9094));
  nand_5 g06746(.A(new_n9094), .B(new_n9041), .Y(new_n9095));
  nand_5 g06747(.A(new_n9095), .B(new_n9040), .Y(new_n9096));
  nand_5 g06748(.A(new_n9096), .B(new_n9033), .Y(new_n9097));
  nand_5 g06749(.A(new_n9097), .B(new_n9032_1), .Y(new_n9098));
  nand_5 g06750(.A(new_n9098), .B(new_n9027), .Y(new_n9099));
  nand_5 g06751(.A(new_n9099), .B(new_n9026), .Y(new_n9100));
  nand_5 g06752(.A(new_n9100), .B(new_n9021), .Y(new_n9101));
  nand_5 g06753(.A(new_n9101), .B(new_n9020), .Y(new_n9102));
  xor_4  g06754(.A(new_n9102), .B(new_n9013), .Y(n829));
  not_8  g06755(.A(n14826), .Y(new_n9104_1));
  nand_5 g06756(.A(new_n4850_1), .B(new_n9104_1), .Y(new_n9105));
  nand_5 g06757(.A(n23272), .B(n14826), .Y(new_n9106));
  not_8  g06758(.A(n23493), .Y(new_n9107));
  nand_5 g06759(.A(new_n9107), .B(new_n4856), .Y(new_n9108));
  nand_5 g06760(.A(n23493), .B(n11481), .Y(new_n9109));
  not_8  g06761(.A(n10275), .Y(new_n9110));
  nand_5 g06762(.A(new_n4862), .B(new_n9110), .Y(new_n9111));
  nand_5 g06763(.A(n16439), .B(n10275), .Y(new_n9112));
  not_8  g06764(.A(n15146), .Y(new_n9113));
  nand_5 g06765(.A(new_n4868), .B(new_n9113), .Y(new_n9114));
  nand_5 g06766(.A(n15241), .B(n15146), .Y(new_n9115));
  not_8  g06767(.A(n11579), .Y(new_n9116));
  nand_5 g06768(.A(new_n9116), .B(new_n4874), .Y(new_n9117));
  nand_5 g06769(.A(n11579), .B(n7678), .Y(new_n9118));
  nand_5 g06770(.A(n3785), .B(n21), .Y(new_n9119));
  not_8  g06771(.A(n21), .Y(new_n9120));
  nand_5 g06772(.A(new_n4880), .B(new_n9120), .Y(new_n9121));
  not_8  g06773(.A(n1682), .Y(new_n9122));
  not_8  g06774(.A(n7963), .Y(new_n9123));
  nand_5 g06775(.A(new_n9123), .B(new_n4892), .Y(new_n9124));
  nand_5 g06776(.A(n7963), .B(n5822), .Y(new_n9125));
  not_8  g06777(.A(n10017), .Y(new_n9126));
  nand_5 g06778(.A(new_n4898), .B(new_n9126), .Y(new_n9127));
  nand_5 g06779(.A(n26443), .B(n10017), .Y(new_n9128));
  nand_5 g06780(.A(new_n9128), .B(new_n2612), .Y(new_n9129_1));
  nand_5 g06781(.A(new_n9129_1), .B(new_n9127), .Y(new_n9130));
  nand_5 g06782(.A(new_n9130), .B(new_n9125), .Y(new_n9131));
  nand_5 g06783(.A(new_n9131), .B(new_n9124), .Y(new_n9132));
  nand_5 g06784(.A(new_n9132), .B(new_n9122), .Y(new_n9133));
  not_8  g06785(.A(new_n9133), .Y(new_n9134));
  nor_5  g06786(.A(new_n9132), .B(new_n9122), .Y(new_n9135));
  nor_5  g06787(.A(new_n9135), .B(n20250), .Y(new_n9136));
  nor_5  g06788(.A(new_n9136), .B(new_n9134), .Y(new_n9137));
  nand_5 g06789(.A(new_n9137), .B(new_n9121), .Y(new_n9138));
  and_5  g06790(.A(new_n9138), .B(new_n9119), .Y(new_n9139));
  nand_5 g06791(.A(new_n9139), .B(new_n9118), .Y(new_n9140));
  nand_5 g06792(.A(new_n9140), .B(new_n9117), .Y(new_n9141));
  nand_5 g06793(.A(new_n9141), .B(new_n9115), .Y(new_n9142));
  nand_5 g06794(.A(new_n9142), .B(new_n9114), .Y(new_n9143));
  nand_5 g06795(.A(new_n9143), .B(new_n9112), .Y(new_n9144));
  nand_5 g06796(.A(new_n9144), .B(new_n9111), .Y(new_n9145));
  nand_5 g06797(.A(new_n9145), .B(new_n9109), .Y(new_n9146_1));
  nand_5 g06798(.A(new_n9146_1), .B(new_n9108), .Y(new_n9147));
  nand_5 g06799(.A(new_n9147), .B(new_n9106), .Y(new_n9148));
  nand_5 g06800(.A(new_n9148), .B(new_n9105), .Y(new_n9149));
  not_8  g06801(.A(new_n9149), .Y(new_n9150));
  not_8  g06802(.A(n22764), .Y(new_n9151));
  nand_5 g06803(.A(new_n9106), .B(new_n9105), .Y(new_n9152));
  xor_4  g06804(.A(new_n9152), .B(new_n9147), .Y(new_n9153));
  nand_5 g06805(.A(new_n9153), .B(new_n9151), .Y(new_n9154));
  not_8  g06806(.A(new_n9153), .Y(new_n9155));
  nand_5 g06807(.A(new_n9155), .B(n22764), .Y(new_n9156));
  not_8  g06808(.A(n26264), .Y(new_n9157));
  nand_5 g06809(.A(new_n9109), .B(new_n9108), .Y(new_n9158));
  xor_4  g06810(.A(new_n9158), .B(new_n9145), .Y(new_n9159));
  nand_5 g06811(.A(new_n9159), .B(new_n9157), .Y(new_n9160));
  not_8  g06812(.A(new_n9159), .Y(new_n9161));
  nand_5 g06813(.A(new_n9161), .B(n26264), .Y(new_n9162));
  not_8  g06814(.A(n7841), .Y(new_n9163));
  nand_5 g06815(.A(new_n9112), .B(new_n9111), .Y(new_n9164_1));
  xor_4  g06816(.A(new_n9164_1), .B(new_n9143), .Y(new_n9165));
  nand_5 g06817(.A(new_n9165), .B(new_n9163), .Y(new_n9166_1));
  not_8  g06818(.A(new_n9165), .Y(new_n9167));
  nand_5 g06819(.A(new_n9167), .B(n7841), .Y(new_n9168));
  not_8  g06820(.A(n16812), .Y(new_n9169));
  nand_5 g06821(.A(new_n9115), .B(new_n9114), .Y(new_n9170));
  xor_4  g06822(.A(new_n9170), .B(new_n9141), .Y(new_n9171));
  nand_5 g06823(.A(new_n9171), .B(new_n9169), .Y(new_n9172_1));
  not_8  g06824(.A(new_n9171), .Y(new_n9173));
  nand_5 g06825(.A(new_n9173), .B(n16812), .Y(new_n9174));
  not_8  g06826(.A(n25068), .Y(new_n9175));
  nand_5 g06827(.A(new_n9118), .B(new_n9117), .Y(new_n9176));
  xor_4  g06828(.A(new_n9176), .B(new_n9139), .Y(new_n9177));
  nand_5 g06829(.A(new_n9177), .B(new_n9175), .Y(new_n9178));
  not_8  g06830(.A(new_n9177), .Y(new_n9179));
  nand_5 g06831(.A(new_n9179), .B(n25068), .Y(new_n9180));
  not_8  g06832(.A(n2331), .Y(new_n9181));
  nand_5 g06833(.A(new_n9121), .B(new_n9119), .Y(new_n9182_1));
  xor_4  g06834(.A(new_n9182_1), .B(new_n9137), .Y(new_n9183));
  not_8  g06835(.A(new_n9183), .Y(new_n9184));
  nand_5 g06836(.A(new_n9184), .B(new_n9181), .Y(new_n9185));
  nand_5 g06837(.A(new_n9183), .B(n2331), .Y(new_n9186));
  not_8  g06838(.A(n22631), .Y(new_n9187));
  nor_5  g06839(.A(new_n9135), .B(new_n9134), .Y(new_n9188));
  xor_4  g06840(.A(new_n9188), .B(new_n4886), .Y(new_n9189));
  not_8  g06841(.A(new_n9189), .Y(new_n9190));
  nand_5 g06842(.A(new_n9190), .B(new_n9187), .Y(new_n9191_1));
  nand_5 g06843(.A(new_n9189), .B(n22631), .Y(new_n9192));
  not_8  g06844(.A(n16743), .Y(new_n9193));
  nand_5 g06845(.A(new_n9125), .B(new_n9124), .Y(new_n9194));
  xor_4  g06846(.A(new_n9194), .B(new_n9130), .Y(new_n9195));
  nand_5 g06847(.A(new_n9195), .B(new_n9193), .Y(new_n9196));
  not_8  g06848(.A(new_n9195), .Y(new_n9197));
  nand_5 g06849(.A(new_n9197), .B(n16743), .Y(new_n9198));
  nand_5 g06850(.A(new_n2616), .B(new_n2611), .Y(new_n9199));
  nand_5 g06851(.A(new_n9199), .B(n15258), .Y(new_n9200));
  or_5   g06852(.A(new_n9199), .B(n15258), .Y(new_n9201));
  nand_5 g06853(.A(new_n9128), .B(new_n9127), .Y(new_n9202));
  not_8  g06854(.A(new_n9202), .Y(new_n9203));
  xor_4  g06855(.A(new_n9203), .B(new_n2612), .Y(new_n9204));
  nand_5 g06856(.A(new_n9204), .B(new_n9201), .Y(new_n9205));
  nand_5 g06857(.A(new_n9205), .B(new_n9200), .Y(new_n9206));
  not_8  g06858(.A(new_n9206), .Y(new_n9207));
  nand_5 g06859(.A(new_n9207), .B(new_n9198), .Y(new_n9208));
  nand_5 g06860(.A(new_n9208), .B(new_n9196), .Y(new_n9209));
  nand_5 g06861(.A(new_n9209), .B(new_n9192), .Y(new_n9210));
  nand_5 g06862(.A(new_n9210), .B(new_n9191_1), .Y(new_n9211));
  nand_5 g06863(.A(new_n9211), .B(new_n9186), .Y(new_n9212));
  nand_5 g06864(.A(new_n9212), .B(new_n9185), .Y(new_n9213));
  nand_5 g06865(.A(new_n9213), .B(new_n9180), .Y(new_n9214));
  nand_5 g06866(.A(new_n9214), .B(new_n9178), .Y(new_n9215));
  nand_5 g06867(.A(new_n9215), .B(new_n9174), .Y(new_n9216));
  nand_5 g06868(.A(new_n9216), .B(new_n9172_1), .Y(new_n9217_1));
  nand_5 g06869(.A(new_n9217_1), .B(new_n9168), .Y(new_n9218));
  nand_5 g06870(.A(new_n9218), .B(new_n9166_1), .Y(new_n9219));
  nand_5 g06871(.A(new_n9219), .B(new_n9162), .Y(new_n9220_1));
  nand_5 g06872(.A(new_n9220_1), .B(new_n9160), .Y(new_n9221));
  nand_5 g06873(.A(new_n9221), .B(new_n9156), .Y(new_n9222));
  nand_5 g06874(.A(new_n9222), .B(new_n9154), .Y(new_n9223));
  nor_5  g06875(.A(new_n9223), .B(new_n9150), .Y(new_n9224));
  not_8  g06876(.A(new_n9224), .Y(new_n9225));
  nand_5 g06877(.A(new_n9223), .B(new_n9150), .Y(new_n9226));
  and_5  g06878(.A(new_n9226), .B(new_n9225), .Y(new_n9227));
  not_8  g06879(.A(new_n9227), .Y(new_n9228));
  not_8  g06880(.A(n18105), .Y(new_n9229));
  nand_5 g06881(.A(new_n9229), .B(n12702), .Y(new_n9230));
  nand_5 g06882(.A(n26797), .B(new_n4928), .Y(new_n9231));
  nand_5 g06883(.A(new_n6168), .B(n24196), .Y(new_n9232));
  not_8  g06884(.A(n16376), .Y(new_n9233));
  nand_5 g06885(.A(n23913), .B(new_n9233), .Y(new_n9234));
  not_8  g06886(.A(n23913), .Y(new_n9235));
  nand_5 g06887(.A(new_n9235), .B(n16376), .Y(new_n9236));
  nand_5 g06888(.A(new_n4929), .B(n22554), .Y(new_n9237));
  nand_5 g06889(.A(n25381), .B(new_n6169), .Y(new_n9238));
  not_8  g06890(.A(n12587), .Y(new_n9239));
  nand_5 g06891(.A(n20429), .B(new_n9239), .Y(new_n9240));
  not_8  g06892(.A(n20429), .Y(new_n9241));
  nand_5 g06893(.A(new_n9241), .B(n12587), .Y(new_n9242));
  nand_5 g06894(.A(n3909), .B(new_n4930), .Y(new_n9243));
  nand_5 g06895(.A(new_n6170), .B(n268), .Y(new_n9244));
  not_8  g06896(.A(n24879), .Y(new_n9245));
  nand_5 g06897(.A(new_n9245), .B(n23974), .Y(new_n9246_1));
  not_8  g06898(.A(n23974), .Y(new_n9247));
  nand_5 g06899(.A(n24879), .B(new_n9247), .Y(new_n9248));
  not_8  g06900(.A(n6785), .Y(new_n9249));
  nand_5 g06901(.A(new_n9249), .B(n2146), .Y(new_n9250));
  not_8  g06902(.A(n2146), .Y(new_n9251_1));
  nand_5 g06903(.A(n6785), .B(new_n9251_1), .Y(new_n9252));
  nand_5 g06904(.A(new_n4931), .B(n22173), .Y(new_n9253));
  nand_5 g06905(.A(n24032), .B(new_n6171_1), .Y(new_n9254));
  nand_5 g06906(.A(new_n9254), .B(new_n2621), .Y(new_n9255));
  nand_5 g06907(.A(new_n9255), .B(new_n9253), .Y(new_n9256));
  nand_5 g06908(.A(new_n9256), .B(new_n9252), .Y(new_n9257));
  nand_5 g06909(.A(new_n9257), .B(new_n9250), .Y(new_n9258));
  nand_5 g06910(.A(new_n9258), .B(new_n9248), .Y(new_n9259_1));
  nand_5 g06911(.A(new_n9259_1), .B(new_n9246_1), .Y(new_n9260));
  nand_5 g06912(.A(new_n9260), .B(new_n9244), .Y(new_n9261_1));
  nand_5 g06913(.A(new_n9261_1), .B(new_n9243), .Y(new_n9262));
  nand_5 g06914(.A(new_n9262), .B(new_n9242), .Y(new_n9263));
  nand_5 g06915(.A(new_n9263), .B(new_n9240), .Y(new_n9264));
  nand_5 g06916(.A(new_n9264), .B(new_n9238), .Y(new_n9265));
  nand_5 g06917(.A(new_n9265), .B(new_n9237), .Y(new_n9266));
  nand_5 g06918(.A(new_n9266), .B(new_n9236), .Y(new_n9267));
  nand_5 g06919(.A(new_n9267), .B(new_n9234), .Y(new_n9268));
  nand_5 g06920(.A(new_n9268), .B(new_n9232), .Y(new_n9269));
  nand_5 g06921(.A(new_n9269), .B(new_n9231), .Y(new_n9270));
  not_8  g06922(.A(n12702), .Y(new_n9271));
  nand_5 g06923(.A(n18105), .B(new_n9271), .Y(new_n9272));
  nand_5 g06924(.A(new_n9272), .B(new_n9270), .Y(new_n9273));
  nand_5 g06925(.A(new_n9273), .B(new_n9230), .Y(new_n9274));
  not_8  g06926(.A(n1536), .Y(new_n9275));
  nand_5 g06927(.A(new_n9272), .B(new_n9230), .Y(new_n9276));
  xor_4  g06928(.A(new_n9276), .B(new_n9270), .Y(new_n9277));
  nand_5 g06929(.A(new_n9277), .B(new_n9275), .Y(new_n9278));
  not_8  g06930(.A(new_n9277), .Y(new_n9279));
  nand_5 g06931(.A(new_n9279), .B(n1536), .Y(new_n9280));
  not_8  g06932(.A(n19454), .Y(new_n9281));
  nand_5 g06933(.A(new_n9232), .B(new_n9231), .Y(new_n9282));
  xor_4  g06934(.A(new_n9282), .B(new_n9268), .Y(new_n9283));
  nand_5 g06935(.A(new_n9283), .B(new_n9281), .Y(new_n9284));
  not_8  g06936(.A(new_n9283), .Y(new_n9285));
  nand_5 g06937(.A(new_n9285), .B(n19454), .Y(new_n9286));
  not_8  g06938(.A(n9445), .Y(new_n9287_1));
  nand_5 g06939(.A(new_n9236), .B(new_n9234), .Y(new_n9288));
  xor_4  g06940(.A(new_n9288), .B(new_n9266), .Y(new_n9289));
  nand_5 g06941(.A(new_n9289), .B(new_n9287_1), .Y(new_n9290));
  not_8  g06942(.A(new_n9289), .Y(new_n9291));
  nand_5 g06943(.A(new_n9291), .B(n9445), .Y(new_n9292));
  not_8  g06944(.A(n1279), .Y(new_n9293));
  nand_5 g06945(.A(new_n9238), .B(new_n9237), .Y(new_n9294));
  xor_4  g06946(.A(new_n9294), .B(new_n9264), .Y(new_n9295));
  nand_5 g06947(.A(new_n9295), .B(new_n9293), .Y(new_n9296));
  not_8  g06948(.A(new_n9295), .Y(new_n9297));
  nand_5 g06949(.A(new_n9297), .B(n1279), .Y(new_n9298));
  not_8  g06950(.A(n8324), .Y(new_n9299));
  nand_5 g06951(.A(new_n9242), .B(new_n9240), .Y(new_n9300));
  xor_4  g06952(.A(new_n9300), .B(new_n9262), .Y(new_n9301));
  nand_5 g06953(.A(new_n9301), .B(new_n9299), .Y(new_n9302));
  not_8  g06954(.A(new_n9301), .Y(new_n9303));
  nand_5 g06955(.A(new_n9303), .B(n8324), .Y(new_n9304));
  not_8  g06956(.A(n12546), .Y(new_n9305));
  nand_5 g06957(.A(new_n9244), .B(new_n9243), .Y(new_n9306));
  xor_4  g06958(.A(new_n9306), .B(new_n9260), .Y(new_n9307));
  nand_5 g06959(.A(new_n9307), .B(new_n9305), .Y(new_n9308_1));
  not_8  g06960(.A(new_n9307), .Y(new_n9309));
  nand_5 g06961(.A(new_n9309), .B(n12546), .Y(new_n9310));
  not_8  g06962(.A(n21078), .Y(new_n9311));
  nand_5 g06963(.A(new_n9248), .B(new_n9246_1), .Y(new_n9312));
  xor_4  g06964(.A(new_n9312), .B(new_n9258), .Y(new_n9313));
  nand_5 g06965(.A(new_n9313), .B(new_n9311), .Y(new_n9314));
  not_8  g06966(.A(new_n9313), .Y(new_n9315));
  nand_5 g06967(.A(new_n9315), .B(n21078), .Y(new_n9316));
  not_8  g06968(.A(n24485), .Y(new_n9317));
  nand_5 g06969(.A(new_n9252), .B(new_n9250), .Y(new_n9318_1));
  xor_4  g06970(.A(new_n9318_1), .B(new_n9256), .Y(new_n9319));
  nand_5 g06971(.A(new_n9319), .B(new_n9317), .Y(new_n9320));
  not_8  g06972(.A(new_n9319), .Y(new_n9321));
  nand_5 g06973(.A(new_n9321), .B(n24485), .Y(new_n9322));
  not_8  g06974(.A(n2420), .Y(new_n9323_1));
  and_5  g06975(.A(new_n9254), .B(new_n9253), .Y(new_n9324));
  xor_4  g06976(.A(new_n9324), .B(new_n2621), .Y(new_n9325));
  not_8  g06977(.A(new_n9325), .Y(new_n9326));
  nand_5 g06978(.A(new_n9326), .B(new_n9323_1), .Y(new_n9327));
  not_8  g06979(.A(new_n2624), .Y(new_n9328));
  nand_5 g06980(.A(new_n9328), .B(n22201), .Y(new_n9329));
  nand_5 g06981(.A(new_n9325), .B(n2420), .Y(new_n9330));
  nand_5 g06982(.A(new_n9330), .B(new_n9329), .Y(new_n9331));
  nand_5 g06983(.A(new_n9331), .B(new_n9327), .Y(new_n9332));
  nand_5 g06984(.A(new_n9332), .B(new_n9322), .Y(new_n9333));
  nand_5 g06985(.A(new_n9333), .B(new_n9320), .Y(new_n9334));
  nand_5 g06986(.A(new_n9334), .B(new_n9316), .Y(new_n9335));
  nand_5 g06987(.A(new_n9335), .B(new_n9314), .Y(new_n9336));
  nand_5 g06988(.A(new_n9336), .B(new_n9310), .Y(new_n9337));
  nand_5 g06989(.A(new_n9337), .B(new_n9308_1), .Y(new_n9338));
  nand_5 g06990(.A(new_n9338), .B(new_n9304), .Y(new_n9339));
  nand_5 g06991(.A(new_n9339), .B(new_n9302), .Y(new_n9340));
  nand_5 g06992(.A(new_n9340), .B(new_n9298), .Y(new_n9341));
  nand_5 g06993(.A(new_n9341), .B(new_n9296), .Y(new_n9342));
  nand_5 g06994(.A(new_n9342), .B(new_n9292), .Y(new_n9343));
  nand_5 g06995(.A(new_n9343), .B(new_n9290), .Y(new_n9344_1));
  nand_5 g06996(.A(new_n9344_1), .B(new_n9286), .Y(new_n9345));
  nand_5 g06997(.A(new_n9345), .B(new_n9284), .Y(new_n9346));
  nand_5 g06998(.A(new_n9346), .B(new_n9280), .Y(new_n9347));
  nand_5 g06999(.A(new_n9347), .B(new_n9278), .Y(new_n9348));
  xnor_4 g07000(.A(new_n9348), .B(new_n9274), .Y(new_n9349));
  nand_5 g07001(.A(new_n9349), .B(new_n9228), .Y(new_n9350));
  nand_5 g07002(.A(new_n9280), .B(new_n9278), .Y(new_n9351));
  xor_4  g07003(.A(new_n9351), .B(new_n9346), .Y(new_n9352));
  nand_5 g07004(.A(new_n9154), .B(new_n9156), .Y(new_n9353));
  xor_4  g07005(.A(new_n9353), .B(new_n9221), .Y(new_n9354));
  nand_5 g07006(.A(new_n9354), .B(new_n9352), .Y(new_n9355));
  or_5   g07007(.A(new_n9354), .B(new_n9352), .Y(new_n9356));
  nand_5 g07008(.A(new_n9286), .B(new_n9284), .Y(new_n9357));
  xor_4  g07009(.A(new_n9357), .B(new_n9344_1), .Y(new_n9358));
  nand_5 g07010(.A(new_n9160), .B(new_n9162), .Y(new_n9359));
  xor_4  g07011(.A(new_n9359), .B(new_n9219), .Y(new_n9360));
  nand_5 g07012(.A(new_n9360), .B(new_n9358), .Y(new_n9361));
  or_5   g07013(.A(new_n9360), .B(new_n9358), .Y(new_n9362));
  nand_5 g07014(.A(new_n9292), .B(new_n9290), .Y(new_n9363));
  xor_4  g07015(.A(new_n9363), .B(new_n9342), .Y(new_n9364_1));
  nand_5 g07016(.A(new_n9166_1), .B(new_n9168), .Y(new_n9365));
  xor_4  g07017(.A(new_n9365), .B(new_n9217_1), .Y(new_n9366));
  nand_5 g07018(.A(new_n9366), .B(new_n9364_1), .Y(new_n9367));
  or_5   g07019(.A(new_n9366), .B(new_n9364_1), .Y(new_n9368));
  nand_5 g07020(.A(new_n9298), .B(new_n9296), .Y(new_n9369));
  xor_4  g07021(.A(new_n9369), .B(new_n9340), .Y(new_n9370));
  nand_5 g07022(.A(new_n9172_1), .B(new_n9174), .Y(new_n9371_1));
  xor_4  g07023(.A(new_n9371_1), .B(new_n9215), .Y(new_n9372_1));
  nand_5 g07024(.A(new_n9372_1), .B(new_n9370), .Y(new_n9373));
  or_5   g07025(.A(new_n9372_1), .B(new_n9370), .Y(new_n9374));
  nand_5 g07026(.A(new_n9304), .B(new_n9302), .Y(new_n9375));
  xor_4  g07027(.A(new_n9375), .B(new_n9338), .Y(new_n9376));
  nand_5 g07028(.A(new_n9178), .B(new_n9180), .Y(new_n9377));
  xor_4  g07029(.A(new_n9377), .B(new_n9213), .Y(new_n9378));
  nand_5 g07030(.A(new_n9378), .B(new_n9376), .Y(new_n9379));
  or_5   g07031(.A(new_n9378), .B(new_n9376), .Y(new_n9380_1));
  nand_5 g07032(.A(new_n9310), .B(new_n9308_1), .Y(new_n9381));
  xor_4  g07033(.A(new_n9381), .B(new_n9336), .Y(new_n9382_1));
  nand_5 g07034(.A(new_n9185), .B(new_n9186), .Y(new_n9383));
  xor_4  g07035(.A(new_n9383), .B(new_n9211), .Y(new_n9384));
  nand_5 g07036(.A(new_n9384), .B(new_n9382_1), .Y(new_n9385));
  or_5   g07037(.A(new_n9384), .B(new_n9382_1), .Y(new_n9386));
  nand_5 g07038(.A(new_n9316), .B(new_n9314), .Y(new_n9387));
  xor_4  g07039(.A(new_n9387), .B(new_n9334), .Y(new_n9388));
  nand_5 g07040(.A(new_n9191_1), .B(new_n9192), .Y(new_n9389));
  xor_4  g07041(.A(new_n9389), .B(new_n9209), .Y(new_n9390));
  nand_5 g07042(.A(new_n9390), .B(new_n9388), .Y(new_n9391));
  or_5   g07043(.A(new_n9390), .B(new_n9388), .Y(new_n9392));
  nand_5 g07044(.A(new_n9322), .B(new_n9320), .Y(new_n9393));
  xor_4  g07045(.A(new_n9393), .B(new_n9332), .Y(new_n9394));
  nand_5 g07046(.A(new_n9198), .B(new_n9196), .Y(new_n9395));
  xor_4  g07047(.A(new_n9395), .B(new_n9207), .Y(new_n9396_1));
  nand_5 g07048(.A(new_n9396_1), .B(new_n9394), .Y(new_n9397));
  or_5   g07049(.A(new_n9396_1), .B(new_n9394), .Y(new_n9398));
  nand_5 g07050(.A(new_n9330), .B(new_n9327), .Y(new_n9399_1));
  xor_4  g07051(.A(new_n9399_1), .B(new_n9329), .Y(new_n9400));
  nand_5 g07052(.A(new_n9200), .B(new_n9201), .Y(new_n9401));
  xor_4  g07053(.A(new_n9401), .B(new_n9204), .Y(new_n9402));
  not_8  g07054(.A(new_n9402), .Y(new_n9403_1));
  nor_5  g07055(.A(new_n9403_1), .B(new_n9400), .Y(new_n9404));
  and_5  g07056(.A(new_n9403_1), .B(new_n9400), .Y(new_n9405));
  nor_5  g07057(.A(new_n9405), .B(new_n2627), .Y(new_n9406));
  nor_5  g07058(.A(new_n9406), .B(new_n9404), .Y(new_n9407));
  nand_5 g07059(.A(new_n9407), .B(new_n9398), .Y(new_n9408));
  nand_5 g07060(.A(new_n9408), .B(new_n9397), .Y(new_n9409));
  nand_5 g07061(.A(new_n9409), .B(new_n9392), .Y(new_n9410));
  nand_5 g07062(.A(new_n9410), .B(new_n9391), .Y(new_n9411));
  nand_5 g07063(.A(new_n9411), .B(new_n9386), .Y(new_n9412));
  nand_5 g07064(.A(new_n9412), .B(new_n9385), .Y(new_n9413));
  nand_5 g07065(.A(new_n9413), .B(new_n9380_1), .Y(new_n9414));
  nand_5 g07066(.A(new_n9414), .B(new_n9379), .Y(new_n9415));
  nand_5 g07067(.A(new_n9415), .B(new_n9374), .Y(new_n9416));
  nand_5 g07068(.A(new_n9416), .B(new_n9373), .Y(new_n9417));
  nand_5 g07069(.A(new_n9417), .B(new_n9368), .Y(new_n9418));
  nand_5 g07070(.A(new_n9418), .B(new_n9367), .Y(new_n9419_1));
  nand_5 g07071(.A(new_n9419_1), .B(new_n9362), .Y(new_n9420));
  nand_5 g07072(.A(new_n9420), .B(new_n9361), .Y(new_n9421));
  nand_5 g07073(.A(new_n9421), .B(new_n9356), .Y(new_n9422));
  nand_5 g07074(.A(new_n9422), .B(new_n9355), .Y(new_n9423_1));
  nand_5 g07075(.A(new_n9423_1), .B(new_n9350), .Y(new_n9424));
  or_5   g07076(.A(new_n9349), .B(new_n9228), .Y(new_n9425));
  nand_5 g07077(.A(new_n9425), .B(new_n9424), .Y(new_n9426));
  nor_5  g07078(.A(new_n9348), .B(new_n9274), .Y(new_n9427));
  xor_4  g07079(.A(new_n9427), .B(new_n9225), .Y(new_n9428));
  xor_4  g07080(.A(new_n9428), .B(new_n9426), .Y(n849));
  nor_5  g07081(.A(new_n2554), .B(new_n2550), .Y(new_n9430_1));
  xor_4  g07082(.A(new_n9430_1), .B(new_n2552), .Y(n858));
  nand_5 g07083(.A(new_n3744), .B(new_n3827), .Y(new_n9432));
  or_5   g07084(.A(new_n9432), .B(n10096), .Y(new_n9433));
  nor_5  g07085(.A(new_n9433), .B(n14790), .Y(new_n9434));
  nand_5 g07086(.A(new_n9434), .B(new_n3732), .Y(new_n9435_1));
  nor_5  g07087(.A(new_n9435_1), .B(n21674), .Y(new_n9436));
  nand_5 g07088(.A(new_n9436), .B(new_n3724), .Y(new_n9437));
  nor_5  g07089(.A(new_n9437), .B(n18444), .Y(new_n9438));
  nand_5 g07090(.A(new_n9438), .B(new_n3716), .Y(new_n9439));
  xor_4  g07091(.A(new_n9439), .B(n3506), .Y(new_n9440));
  xor_4  g07092(.A(new_n9440), .B(n1314), .Y(new_n9441));
  xor_4  g07093(.A(new_n9438), .B(new_n3716), .Y(new_n9442));
  or_5   g07094(.A(new_n9442), .B(n3306), .Y(new_n9443));
  nand_5 g07095(.A(new_n9442), .B(n3306), .Y(new_n9444));
  xor_4  g07096(.A(new_n9437), .B(n18444), .Y(new_n9445_1));
  or_5   g07097(.A(new_n9445_1), .B(n22335), .Y(new_n9446));
  nand_5 g07098(.A(new_n9445_1), .B(n22335), .Y(new_n9447));
  xor_4  g07099(.A(new_n9436), .B(new_n3724), .Y(new_n9448));
  or_5   g07100(.A(new_n9448), .B(n24048), .Y(new_n9449));
  nand_5 g07101(.A(new_n9448), .B(n24048), .Y(new_n9450));
  xor_4  g07102(.A(new_n9435_1), .B(n21674), .Y(new_n9451_1));
  or_5   g07103(.A(new_n9451_1), .B(n1525), .Y(new_n9452));
  nand_5 g07104(.A(new_n9451_1), .B(n1525), .Y(new_n9453));
  xor_4  g07105(.A(new_n9434), .B(new_n3732), .Y(new_n9454));
  or_5   g07106(.A(new_n9454), .B(n16988), .Y(new_n9455));
  nand_5 g07107(.A(new_n9454), .B(n16988), .Y(new_n9456));
  xor_4  g07108(.A(new_n9433), .B(n14790), .Y(new_n9457));
  or_5   g07109(.A(new_n9457), .B(n21779), .Y(new_n9458_1));
  nand_5 g07110(.A(new_n9457), .B(n21779), .Y(new_n9459_1));
  nand_5 g07111(.A(new_n9432), .B(n10096), .Y(new_n9460_1));
  and_5  g07112(.A(new_n9460_1), .B(new_n9433), .Y(new_n9461));
  or_5   g07113(.A(new_n9461), .B(n5376), .Y(new_n9462));
  nand_5 g07114(.A(new_n9461), .B(n5376), .Y(new_n9463));
  nand_5 g07115(.A(n16994), .B(n9246), .Y(new_n9464));
  and_5  g07116(.A(new_n9464), .B(new_n9432), .Y(new_n9465));
  or_5   g07117(.A(new_n9465), .B(n5128), .Y(new_n9466));
  nand_5 g07118(.A(new_n9465), .B(n5128), .Y(new_n9467));
  nand_5 g07119(.A(n23120), .B(n9246), .Y(new_n9468));
  nand_5 g07120(.A(new_n9468), .B(new_n9467), .Y(new_n9469));
  nand_5 g07121(.A(new_n9469), .B(new_n9466), .Y(new_n9470));
  nand_5 g07122(.A(new_n9470), .B(new_n9463), .Y(new_n9471));
  nand_5 g07123(.A(new_n9471), .B(new_n9462), .Y(new_n9472));
  nand_5 g07124(.A(new_n9472), .B(new_n9459_1), .Y(new_n9473));
  nand_5 g07125(.A(new_n9473), .B(new_n9458_1), .Y(new_n9474));
  nand_5 g07126(.A(new_n9474), .B(new_n9456), .Y(new_n9475));
  nand_5 g07127(.A(new_n9475), .B(new_n9455), .Y(new_n9476));
  nand_5 g07128(.A(new_n9476), .B(new_n9453), .Y(new_n9477));
  nand_5 g07129(.A(new_n9477), .B(new_n9452), .Y(new_n9478));
  nand_5 g07130(.A(new_n9478), .B(new_n9450), .Y(new_n9479));
  nand_5 g07131(.A(new_n9479), .B(new_n9449), .Y(new_n9480));
  nand_5 g07132(.A(new_n9480), .B(new_n9447), .Y(new_n9481));
  nand_5 g07133(.A(new_n9481), .B(new_n9446), .Y(new_n9482));
  nand_5 g07134(.A(new_n9482), .B(new_n9444), .Y(new_n9483));
  nand_5 g07135(.A(new_n9483), .B(new_n9443), .Y(new_n9484));
  xor_4  g07136(.A(new_n9484), .B(new_n9441), .Y(new_n9485));
  or_5   g07137(.A(new_n9485), .B(n22442), .Y(new_n9486));
  nand_5 g07138(.A(new_n9485), .B(n22442), .Y(new_n9487));
  nand_5 g07139(.A(new_n9444), .B(new_n9443), .Y(new_n9488));
  xor_4  g07140(.A(new_n9488), .B(new_n9482), .Y(new_n9489));
  nand_5 g07141(.A(new_n9489), .B(new_n8019), .Y(new_n9490));
  or_5   g07142(.A(new_n9489), .B(new_n8019), .Y(new_n9491));
  nand_5 g07143(.A(new_n9447), .B(new_n9446), .Y(new_n9492));
  xor_4  g07144(.A(new_n9492), .B(new_n9480), .Y(new_n9493_1));
  nand_5 g07145(.A(new_n9493_1), .B(new_n8023), .Y(new_n9494));
  or_5   g07146(.A(new_n9493_1), .B(new_n8023), .Y(new_n9495));
  nand_5 g07147(.A(new_n9450), .B(new_n9449), .Y(new_n9496));
  xor_4  g07148(.A(new_n9496), .B(new_n9478), .Y(new_n9497));
  nand_5 g07149(.A(new_n9497), .B(new_n8028), .Y(new_n9498));
  not_8  g07150(.A(new_n9498), .Y(new_n9499));
  nor_5  g07151(.A(new_n9497), .B(new_n8028), .Y(new_n9500));
  nand_5 g07152(.A(new_n9453), .B(new_n9452), .Y(new_n9501));
  xor_4  g07153(.A(new_n9501), .B(new_n9476), .Y(new_n9502));
  nand_5 g07154(.A(new_n9502), .B(new_n8031_1), .Y(new_n9503));
  not_8  g07155(.A(new_n9503), .Y(new_n9504));
  not_8  g07156(.A(new_n9502), .Y(new_n9505));
  nand_5 g07157(.A(new_n9505), .B(n329), .Y(new_n9506));
  not_8  g07158(.A(new_n9506), .Y(new_n9507_1));
  nand_5 g07159(.A(new_n9459_1), .B(new_n9458_1), .Y(new_n9508_1));
  xor_4  g07160(.A(new_n9508_1), .B(new_n9472), .Y(new_n9509));
  nand_5 g07161(.A(new_n9509), .B(new_n8034), .Y(new_n9510));
  or_5   g07162(.A(new_n9509), .B(new_n8034), .Y(new_n9511));
  nand_5 g07163(.A(new_n9463), .B(new_n9462), .Y(new_n9512_1));
  xor_4  g07164(.A(new_n9512_1), .B(new_n9470), .Y(new_n9513));
  nand_5 g07165(.A(new_n9513), .B(new_n8035), .Y(new_n9514));
  nor_5  g07166(.A(new_n9513), .B(new_n8035), .Y(new_n9515));
  not_8  g07167(.A(new_n9515), .Y(new_n9516));
  and_5  g07168(.A(new_n9467), .B(new_n9466), .Y(new_n9517));
  xor_4  g07169(.A(new_n9517), .B(new_n9468), .Y(new_n9518));
  or_5   g07170(.A(new_n9518), .B(n10372), .Y(new_n9519));
  nand_5 g07171(.A(new_n9518), .B(n10372), .Y(new_n9520));
  nand_5 g07172(.A(new_n5144), .B(new_n3827), .Y(new_n9521));
  nand_5 g07173(.A(new_n9521), .B(new_n9468), .Y(new_n9522));
  nand_5 g07174(.A(new_n9522), .B(n7428), .Y(new_n9523));
  nand_5 g07175(.A(new_n9523), .B(new_n9520), .Y(new_n9524));
  nand_5 g07176(.A(new_n9524), .B(new_n9519), .Y(new_n9525));
  nand_5 g07177(.A(new_n9525), .B(new_n9516), .Y(new_n9526));
  nand_5 g07178(.A(new_n9526), .B(new_n9514), .Y(new_n9527));
  nand_5 g07179(.A(new_n9527), .B(new_n9511), .Y(new_n9528));
  nand_5 g07180(.A(new_n9528), .B(new_n9510), .Y(new_n9529));
  nand_5 g07181(.A(new_n9529), .B(new_n8052_1), .Y(new_n9530));
  not_8  g07182(.A(new_n9530), .Y(new_n9531));
  nor_5  g07183(.A(new_n9529), .B(new_n8052_1), .Y(new_n9532));
  nand_5 g07184(.A(new_n9456), .B(new_n9455), .Y(new_n9533));
  xnor_4 g07185(.A(new_n9533), .B(new_n9474), .Y(new_n9534));
  nor_5  g07186(.A(new_n9534), .B(new_n9532), .Y(new_n9535));
  nor_5  g07187(.A(new_n9535), .B(new_n9531), .Y(new_n9536));
  nor_5  g07188(.A(new_n9536), .B(new_n9507_1), .Y(new_n9537));
  nor_5  g07189(.A(new_n9537), .B(new_n9504), .Y(new_n9538));
  nor_5  g07190(.A(new_n9538), .B(new_n9500), .Y(new_n9539));
  nor_5  g07191(.A(new_n9539), .B(new_n9499), .Y(new_n9540));
  not_8  g07192(.A(new_n9540), .Y(new_n9541));
  nand_5 g07193(.A(new_n9541), .B(new_n9495), .Y(new_n9542));
  nand_5 g07194(.A(new_n9542), .B(new_n9494), .Y(new_n9543));
  nand_5 g07195(.A(new_n9543), .B(new_n9491), .Y(new_n9544));
  nand_5 g07196(.A(new_n9544), .B(new_n9490), .Y(new_n9545));
  nand_5 g07197(.A(new_n9545), .B(new_n9487), .Y(new_n9546));
  nand_5 g07198(.A(new_n9546), .B(new_n9486), .Y(new_n9547));
  nor_5  g07199(.A(new_n9440), .B(n1314), .Y(new_n9548));
  nor_5  g07200(.A(new_n9484), .B(new_n9548), .Y(new_n9549));
  or_5   g07201(.A(new_n9439), .B(n3506), .Y(new_n9550));
  nand_5 g07202(.A(new_n9440), .B(n1314), .Y(new_n9551));
  nand_5 g07203(.A(new_n9551), .B(new_n9550), .Y(new_n9552_1));
  nor_5  g07204(.A(new_n9552_1), .B(new_n9549), .Y(new_n9553));
  not_8  g07205(.A(new_n9553), .Y(new_n9554_1));
  xor_4  g07206(.A(new_n9554_1), .B(new_n9547), .Y(new_n9555));
  nor_5  g07207(.A(new_n3904), .B(n25494), .Y(new_n9556_1));
  nor_5  g07208(.A(new_n9556_1), .B(new_n3903), .Y(new_n9557_1));
  nand_5 g07209(.A(new_n3859), .B(new_n7991), .Y(new_n9558_1));
  nand_5 g07210(.A(new_n3904), .B(n25494), .Y(new_n9559));
  nand_5 g07211(.A(new_n9559), .B(new_n9558_1), .Y(new_n9560));
  nor_5  g07212(.A(new_n9560), .B(new_n9557_1), .Y(new_n9561));
  nand_5 g07213(.A(new_n3980), .B(new_n3910), .Y(new_n9562));
  nand_5 g07214(.A(new_n9562), .B(new_n3908), .Y(new_n9563));
  nor_5  g07215(.A(new_n9563), .B(new_n9561), .Y(new_n9564));
  nand_5 g07216(.A(new_n9563), .B(new_n9561), .Y(new_n9565));
  not_8  g07217(.A(new_n9565), .Y(new_n9566));
  nor_5  g07218(.A(new_n9566), .B(new_n9564), .Y(new_n9567));
  or_5   g07219(.A(new_n9567), .B(new_n9555), .Y(new_n9568));
  nand_5 g07220(.A(new_n9567), .B(new_n9555), .Y(new_n9569));
  nand_5 g07221(.A(new_n9569), .B(new_n9568), .Y(new_n9570));
  nand_5 g07222(.A(new_n9487), .B(new_n9486), .Y(new_n9571));
  xor_4  g07223(.A(new_n9571), .B(new_n9545), .Y(new_n9572));
  nand_5 g07224(.A(new_n9572), .B(new_n3981), .Y(new_n9573));
  or_5   g07225(.A(new_n9572), .B(new_n3981), .Y(new_n9574));
  nand_5 g07226(.A(new_n9491), .B(new_n9490), .Y(new_n9575));
  xor_4  g07227(.A(new_n9575), .B(new_n9543), .Y(new_n9576));
  nand_5 g07228(.A(new_n9576), .B(new_n3987), .Y(new_n9577));
  or_5   g07229(.A(new_n9576), .B(new_n3987), .Y(new_n9578));
  nand_5 g07230(.A(new_n9495), .B(new_n9494), .Y(new_n9579));
  xor_4  g07231(.A(new_n9579), .B(new_n9541), .Y(new_n9580));
  nand_5 g07232(.A(new_n9580), .B(new_n3996), .Y(new_n9581));
  or_5   g07233(.A(new_n9580), .B(new_n3996), .Y(new_n9582));
  nor_5  g07234(.A(new_n9500), .B(new_n9499), .Y(new_n9583));
  xor_4  g07235(.A(new_n9583), .B(new_n9538), .Y(new_n9584));
  nand_5 g07236(.A(new_n9584), .B(new_n4001), .Y(new_n9585));
  or_5   g07237(.A(new_n9584), .B(new_n4001), .Y(new_n9586));
  nand_5 g07238(.A(new_n9506), .B(new_n9503), .Y(new_n9587));
  xor_4  g07239(.A(new_n9587), .B(new_n9536), .Y(new_n9588));
  or_5   g07240(.A(new_n9588), .B(new_n4009), .Y(new_n9589));
  nand_5 g07241(.A(new_n9588), .B(new_n4009), .Y(new_n9590));
  nor_5  g07242(.A(new_n9532), .B(new_n9531), .Y(new_n9591));
  xor_4  g07243(.A(new_n9591), .B(new_n9534), .Y(new_n9592));
  nand_5 g07244(.A(new_n9592), .B(new_n4017), .Y(new_n9593));
  or_5   g07245(.A(new_n9592), .B(new_n4017), .Y(new_n9594));
  nand_5 g07246(.A(new_n9511), .B(new_n9510), .Y(new_n9595));
  xor_4  g07247(.A(new_n9595), .B(new_n9527), .Y(new_n9596));
  nand_5 g07248(.A(new_n9596), .B(new_n4024), .Y(new_n9597));
  or_5   g07249(.A(new_n9596), .B(new_n4024), .Y(new_n9598_1));
  nand_5 g07250(.A(new_n9516), .B(new_n9514), .Y(new_n9599));
  xor_4  g07251(.A(new_n9599), .B(new_n9525), .Y(new_n9600));
  nand_5 g07252(.A(new_n9600), .B(new_n4029), .Y(new_n9601));
  nor_5  g07253(.A(new_n9600), .B(new_n4029), .Y(new_n9602));
  not_8  g07254(.A(new_n9602), .Y(new_n9603));
  xor_4  g07255(.A(new_n9522), .B(n7428), .Y(new_n9604));
  nor_5  g07256(.A(new_n9604), .B(new_n4043), .Y(new_n9605));
  not_8  g07257(.A(new_n9605), .Y(new_n9606));
  nor_5  g07258(.A(new_n9606), .B(new_n4037), .Y(new_n9607));
  nand_5 g07259(.A(new_n9606), .B(new_n4038), .Y(new_n9608));
  not_8  g07260(.A(new_n9608), .Y(new_n9609));
  nand_5 g07261(.A(new_n9520), .B(new_n9519), .Y(new_n9610));
  xor_4  g07262(.A(new_n9610), .B(new_n9523), .Y(new_n9611));
  nor_5  g07263(.A(new_n9611), .B(new_n9609), .Y(new_n9612));
  nor_5  g07264(.A(new_n9612), .B(new_n9607), .Y(new_n9613));
  nand_5 g07265(.A(new_n9613), .B(new_n9603), .Y(new_n9614));
  nand_5 g07266(.A(new_n9614), .B(new_n9601), .Y(new_n9615));
  nand_5 g07267(.A(new_n9615), .B(new_n9598_1), .Y(new_n9616_1));
  nand_5 g07268(.A(new_n9616_1), .B(new_n9597), .Y(new_n9617));
  nand_5 g07269(.A(new_n9617), .B(new_n9594), .Y(new_n9618));
  nand_5 g07270(.A(new_n9618), .B(new_n9593), .Y(new_n9619));
  nand_5 g07271(.A(new_n9619), .B(new_n9590), .Y(new_n9620));
  nand_5 g07272(.A(new_n9620), .B(new_n9589), .Y(new_n9621));
  nand_5 g07273(.A(new_n9621), .B(new_n9586), .Y(new_n9622_1));
  nand_5 g07274(.A(new_n9622_1), .B(new_n9585), .Y(new_n9623));
  nand_5 g07275(.A(new_n9623), .B(new_n9582), .Y(new_n9624));
  nand_5 g07276(.A(new_n9624), .B(new_n9581), .Y(new_n9625));
  nand_5 g07277(.A(new_n9625), .B(new_n9578), .Y(new_n9626_1));
  nand_5 g07278(.A(new_n9626_1), .B(new_n9577), .Y(new_n9627));
  nand_5 g07279(.A(new_n9627), .B(new_n9574), .Y(new_n9628));
  nand_5 g07280(.A(new_n9628), .B(new_n9573), .Y(new_n9629));
  xor_4  g07281(.A(new_n9629), .B(new_n9570), .Y(n873));
  nand_5 g07282(.A(n24618), .B(new_n2393), .Y(new_n9631));
  nand_5 g07283(.A(new_n2354), .B(n13708), .Y(new_n9632));
  nand_5 g07284(.A(new_n2384), .B(n3952), .Y(new_n9633_1));
  nand_5 g07285(.A(n18409), .B(new_n2357), .Y(new_n9634));
  nand_5 g07286(.A(new_n2443), .B(n5704), .Y(new_n9635_1));
  nand_5 g07287(.A(new_n9635_1), .B(new_n9634), .Y(new_n9636));
  nand_5 g07288(.A(new_n9636), .B(new_n9633_1), .Y(new_n9637));
  nand_5 g07289(.A(new_n9637), .B(new_n9632), .Y(new_n9638));
  nand_5 g07290(.A(new_n9638), .B(new_n9631), .Y(new_n9639));
  nand_5 g07291(.A(n24278), .B(new_n2402), .Y(new_n9640));
  nand_5 g07292(.A(new_n2350), .B(n19911), .Y(new_n9641));
  nand_5 g07293(.A(new_n9641), .B(new_n9640), .Y(new_n9642));
  xor_4  g07294(.A(new_n9642), .B(new_n9639), .Y(new_n9643));
  nand_5 g07295(.A(new_n9643), .B(new_n5828), .Y(new_n9644));
  or_5   g07296(.A(new_n9643), .B(new_n5828), .Y(new_n9645));
  nand_5 g07297(.A(new_n9632), .B(new_n9631), .Y(new_n9646_1));
  xor_4  g07298(.A(new_n9646_1), .B(new_n9637), .Y(new_n9647));
  nand_5 g07299(.A(new_n9647), .B(new_n5834_1), .Y(new_n9648_1));
  or_5   g07300(.A(new_n9647), .B(new_n5834_1), .Y(new_n9649));
  xor_4  g07301(.A(n12315), .B(new_n2377), .Y(new_n9650));
  nor_5  g07302(.A(new_n9650), .B(new_n5839), .Y(new_n9651));
  nand_5 g07303(.A(new_n9651), .B(new_n5847), .Y(new_n9652));
  or_5   g07304(.A(new_n9651), .B(new_n5847), .Y(new_n9653));
  nand_5 g07305(.A(new_n9634), .B(new_n9633_1), .Y(new_n9654));
  xnor_4 g07306(.A(new_n9654), .B(new_n9635_1), .Y(new_n9655_1));
  nand_5 g07307(.A(new_n9655_1), .B(new_n9653), .Y(new_n9656));
  nand_5 g07308(.A(new_n9656), .B(new_n9652), .Y(new_n9657));
  not_8  g07309(.A(new_n9657), .Y(new_n9658));
  nand_5 g07310(.A(new_n9658), .B(new_n9649), .Y(new_n9659));
  nand_5 g07311(.A(new_n9659), .B(new_n9648_1), .Y(new_n9660));
  nand_5 g07312(.A(new_n9660), .B(new_n9645), .Y(new_n9661));
  nand_5 g07313(.A(new_n9661), .B(new_n9644), .Y(new_n9662));
  not_8  g07314(.A(new_n5804), .Y(new_n9663));
  nand_5 g07315(.A(new_n9641), .B(new_n9639), .Y(new_n9664));
  nand_5 g07316(.A(new_n9664), .B(new_n9640), .Y(new_n9665));
  nand_5 g07317(.A(n4812), .B(new_n2411), .Y(new_n9666));
  nand_5 g07318(.A(new_n2371), .B(n2731), .Y(new_n9667));
  nand_5 g07319(.A(new_n9667), .B(new_n9666), .Y(new_n9668));
  xnor_4 g07320(.A(new_n9668), .B(new_n9665), .Y(new_n9669));
  or_5   g07321(.A(new_n9669), .B(new_n9663), .Y(new_n9670));
  nand_5 g07322(.A(new_n9669), .B(new_n9663), .Y(new_n9671));
  nand_5 g07323(.A(new_n9671), .B(new_n9670), .Y(new_n9672));
  xor_4  g07324(.A(new_n9672), .B(new_n9662), .Y(n879));
  nand_5 g07325(.A(new_n7573), .B(n14684), .Y(new_n9674));
  nand_5 g07326(.A(new_n7572_1), .B(new_n4620), .Y(new_n9675));
  nand_5 g07327(.A(new_n7555), .B(n6631), .Y(new_n9676));
  nand_5 g07328(.A(new_n7554), .B(new_n4621), .Y(new_n9677));
  nand_5 g07329(.A(new_n7560), .B(n24732), .Y(new_n9678));
  not_8  g07330(.A(new_n9678), .Y(new_n9679));
  nand_5 g07331(.A(new_n9679), .B(new_n9677), .Y(new_n9680));
  nand_5 g07332(.A(new_n9680), .B(new_n9676), .Y(new_n9681));
  nand_5 g07333(.A(new_n9681), .B(new_n9675), .Y(new_n9682));
  nand_5 g07334(.A(new_n9682), .B(new_n9674), .Y(new_n9683));
  nand_5 g07335(.A(new_n7625), .B(n17035), .Y(new_n9684));
  nand_5 g07336(.A(new_n7624), .B(new_n4642), .Y(new_n9685));
  nand_5 g07337(.A(new_n9685), .B(new_n9684), .Y(new_n9686));
  xor_4  g07338(.A(new_n9686), .B(new_n9683), .Y(new_n9687));
  not_8  g07339(.A(new_n9687), .Y(new_n9688));
  or_5   g07340(.A(new_n9204), .B(new_n7519), .Y(new_n9689_1));
  nand_5 g07341(.A(new_n9204), .B(new_n7519), .Y(new_n9690));
  nand_5 g07342(.A(new_n2616), .B(n8581), .Y(new_n9691));
  not_8  g07343(.A(new_n9691), .Y(new_n9692));
  nand_5 g07344(.A(new_n9692), .B(new_n9690), .Y(new_n9693));
  nand_5 g07345(.A(new_n9693), .B(new_n9689_1), .Y(new_n9694));
  nand_5 g07346(.A(new_n9195), .B(n12161), .Y(new_n9695_1));
  nand_5 g07347(.A(new_n9197), .B(new_n7538), .Y(new_n9696));
  nand_5 g07348(.A(new_n9696), .B(new_n9695_1), .Y(new_n9697));
  xor_4  g07349(.A(new_n9697), .B(new_n9694), .Y(new_n9698));
  nand_5 g07350(.A(new_n9674), .B(new_n9675), .Y(new_n9699_1));
  xor_4  g07351(.A(new_n9699_1), .B(new_n9681), .Y(new_n9700));
  not_8  g07352(.A(new_n9700), .Y(new_n9701));
  nand_5 g07353(.A(new_n9701), .B(new_n9698), .Y(new_n9702));
  or_5   g07354(.A(new_n9701), .B(new_n9698), .Y(new_n9703));
  nand_5 g07355(.A(new_n9689_1), .B(new_n9690), .Y(new_n9704));
  xor_4  g07356(.A(new_n9704), .B(new_n9692), .Y(new_n9705));
  nand_5 g07357(.A(new_n9676), .B(new_n9677), .Y(new_n9706));
  xor_4  g07358(.A(new_n9706), .B(new_n9679), .Y(new_n9707));
  not_8  g07359(.A(new_n9707), .Y(new_n9708));
  nand_5 g07360(.A(new_n9708), .B(new_n9705), .Y(new_n9709));
  nor_5  g07361(.A(new_n9708), .B(new_n9705), .Y(new_n9710));
  not_8  g07362(.A(new_n9710), .Y(new_n9711));
  nand_5 g07363(.A(new_n7591), .B(new_n4622), .Y(new_n9712));
  and_5  g07364(.A(new_n9712), .B(new_n9678), .Y(new_n9713));
  not_8  g07365(.A(new_n2616), .Y(new_n9714));
  nand_5 g07366(.A(new_n9714), .B(new_n7526), .Y(new_n9715));
  nand_5 g07367(.A(new_n9715), .B(new_n9691), .Y(new_n9716));
  nand_5 g07368(.A(new_n9716), .B(new_n9713), .Y(new_n9717));
  not_8  g07369(.A(new_n9717), .Y(new_n9718));
  nand_5 g07370(.A(new_n9718), .B(new_n9711), .Y(new_n9719));
  nand_5 g07371(.A(new_n9719), .B(new_n9709), .Y(new_n9720));
  nand_5 g07372(.A(new_n9720), .B(new_n9703), .Y(new_n9721));
  nand_5 g07373(.A(new_n9721), .B(new_n9702), .Y(new_n9722));
  nand_5 g07374(.A(new_n9696), .B(new_n9694), .Y(new_n9723));
  nand_5 g07375(.A(new_n9723), .B(new_n9695_1), .Y(new_n9724));
  nand_5 g07376(.A(new_n9190), .B(n18157), .Y(new_n9725));
  nand_5 g07377(.A(new_n9189), .B(new_n7606), .Y(new_n9726_1));
  nand_5 g07378(.A(new_n9726_1), .B(new_n9725), .Y(new_n9727));
  xnor_4 g07379(.A(new_n9727), .B(new_n9724), .Y(new_n9728));
  not_8  g07380(.A(new_n9728), .Y(new_n9729));
  nand_5 g07381(.A(new_n9729), .B(new_n9722), .Y(new_n9730));
  nor_5  g07382(.A(new_n9729), .B(new_n9722), .Y(new_n9731));
  not_8  g07383(.A(new_n9731), .Y(new_n9732));
  nand_5 g07384(.A(new_n9732), .B(new_n9730), .Y(new_n9733));
  xor_4  g07385(.A(new_n9733), .B(new_n9688), .Y(n887));
  nand_5 g07386(.A(new_n6874), .B(n20826), .Y(new_n9735));
  nand_5 g07387(.A(new_n6875), .B(new_n5526), .Y(new_n9736));
  nand_5 g07388(.A(new_n6880), .B(n7305), .Y(new_n9737));
  nand_5 g07389(.A(new_n6881), .B(new_n5532_1), .Y(new_n9738));
  nand_5 g07390(.A(new_n6886), .B(n25872), .Y(new_n9739));
  nand_5 g07391(.A(new_n6887), .B(new_n5538), .Y(new_n9740));
  nand_5 g07392(.A(new_n6891), .B(n20259), .Y(new_n9741));
  nand_5 g07393(.A(new_n6892), .B(new_n5544), .Y(new_n9742));
  nand_5 g07394(.A(new_n6563), .B(n3925), .Y(new_n9743));
  not_8  g07395(.A(new_n9743), .Y(new_n9744));
  nand_5 g07396(.A(new_n9744), .B(new_n9742), .Y(new_n9745));
  nand_5 g07397(.A(new_n9745), .B(new_n9741), .Y(new_n9746));
  nand_5 g07398(.A(new_n9746), .B(new_n9740), .Y(new_n9747));
  nand_5 g07399(.A(new_n9747), .B(new_n9739), .Y(new_n9748));
  nand_5 g07400(.A(new_n9748), .B(new_n9738), .Y(new_n9749));
  nand_5 g07401(.A(new_n9749), .B(new_n9737), .Y(new_n9750));
  nand_5 g07402(.A(new_n9750), .B(new_n9736), .Y(new_n9751));
  nand_5 g07403(.A(new_n9751), .B(new_n9735), .Y(new_n9752));
  nand_5 g07404(.A(new_n6869), .B(n22198), .Y(new_n9753_1));
  nand_5 g07405(.A(new_n6870), .B(new_n5520), .Y(new_n9754));
  nand_5 g07406(.A(new_n9754), .B(new_n9753_1), .Y(new_n9755));
  xor_4  g07407(.A(new_n9755), .B(new_n9752), .Y(new_n9756));
  not_8  g07408(.A(n18537), .Y(new_n9757));
  nand_5 g07409(.A(new_n3127), .B(new_n9757), .Y(new_n9758));
  nand_5 g07410(.A(new_n3126_1), .B(n18537), .Y(new_n9759));
  not_8  g07411(.A(n7057), .Y(new_n9760));
  nand_5 g07412(.A(new_n3135), .B(new_n9760), .Y(new_n9761_1));
  nand_5 g07413(.A(new_n3134), .B(n7057), .Y(new_n9762));
  nand_5 g07414(.A(new_n3144), .B(new_n5709), .Y(new_n9763_1));
  nand_5 g07415(.A(new_n3143), .B(n8381), .Y(new_n9764));
  not_8  g07416(.A(n20235), .Y(new_n9765));
  nand_5 g07417(.A(new_n3161_1), .B(n12495), .Y(new_n9766));
  nand_5 g07418(.A(new_n9766), .B(new_n9765), .Y(new_n9767_1));
  not_8  g07419(.A(new_n9766), .Y(new_n9768));
  nand_5 g07420(.A(new_n9768), .B(n20235), .Y(new_n9769));
  nand_5 g07421(.A(new_n9769), .B(new_n3152), .Y(new_n9770));
  nand_5 g07422(.A(new_n9770), .B(new_n9767_1), .Y(new_n9771_1));
  nand_5 g07423(.A(new_n9771_1), .B(new_n9764), .Y(new_n9772));
  nand_5 g07424(.A(new_n9772), .B(new_n9763_1), .Y(new_n9773));
  nand_5 g07425(.A(new_n9773), .B(new_n9762), .Y(new_n9774));
  nand_5 g07426(.A(new_n9774), .B(new_n9761_1), .Y(new_n9775));
  nand_5 g07427(.A(new_n9775), .B(new_n9759), .Y(new_n9776));
  nand_5 g07428(.A(new_n9776), .B(new_n9758), .Y(new_n9777));
  not_8  g07429(.A(n1163), .Y(new_n9778_1));
  nand_5 g07430(.A(new_n3119), .B(new_n9778_1), .Y(new_n9779));
  nand_5 g07431(.A(new_n3118), .B(n1163), .Y(new_n9780));
  nand_5 g07432(.A(new_n9780), .B(new_n9779), .Y(new_n9781));
  xor_4  g07433(.A(new_n9781), .B(new_n9777), .Y(new_n9782));
  nand_5 g07434(.A(new_n9782), .B(new_n9756), .Y(new_n9783_1));
  or_5   g07435(.A(new_n9782), .B(new_n9756), .Y(new_n9784));
  nand_5 g07436(.A(new_n9735), .B(new_n9736), .Y(new_n9785));
  xor_4  g07437(.A(new_n9785), .B(new_n9750), .Y(new_n9786));
  nand_5 g07438(.A(new_n9758), .B(new_n9759), .Y(new_n9787));
  xor_4  g07439(.A(new_n9787), .B(new_n9775), .Y(new_n9788));
  nand_5 g07440(.A(new_n9788), .B(new_n9786), .Y(new_n9789));
  or_5   g07441(.A(new_n9788), .B(new_n9786), .Y(new_n9790));
  nand_5 g07442(.A(new_n9737), .B(new_n9738), .Y(new_n9791));
  xor_4  g07443(.A(new_n9791), .B(new_n9748), .Y(new_n9792));
  nand_5 g07444(.A(new_n9761_1), .B(new_n9762), .Y(new_n9793));
  xor_4  g07445(.A(new_n9793), .B(new_n9773), .Y(new_n9794));
  nand_5 g07446(.A(new_n9794), .B(new_n9792), .Y(new_n9795));
  or_5   g07447(.A(new_n9794), .B(new_n9792), .Y(new_n9796));
  nand_5 g07448(.A(new_n9739), .B(new_n9740), .Y(new_n9797));
  xor_4  g07449(.A(new_n9797), .B(new_n9746), .Y(new_n9798));
  nand_5 g07450(.A(new_n9763_1), .B(new_n9764), .Y(new_n9799));
  xor_4  g07451(.A(new_n9799), .B(new_n9771_1), .Y(new_n9800));
  nand_5 g07452(.A(new_n9800), .B(new_n9798), .Y(new_n9801));
  or_5   g07453(.A(new_n9800), .B(new_n9798), .Y(new_n9802));
  nand_5 g07454(.A(new_n9741), .B(new_n9742), .Y(new_n9803_1));
  xor_4  g07455(.A(new_n9803_1), .B(new_n9744), .Y(new_n9804));
  not_8  g07456(.A(new_n9804), .Y(new_n9805));
  and_5  g07457(.A(new_n9767_1), .B(new_n9769), .Y(new_n9806));
  xor_4  g07458(.A(new_n9806), .B(new_n3152), .Y(new_n9807));
  or_5   g07459(.A(new_n9807), .B(new_n9805), .Y(new_n9808));
  nand_5 g07460(.A(new_n9807), .B(new_n9805), .Y(new_n9809));
  nand_5 g07461(.A(new_n6565), .B(new_n5549), .Y(new_n9810));
  and_5  g07462(.A(new_n9810), .B(new_n9743), .Y(new_n9811));
  nand_5 g07463(.A(new_n3162), .B(new_n5669), .Y(new_n9812));
  nand_5 g07464(.A(new_n9812), .B(new_n9766), .Y(new_n9813));
  nand_5 g07465(.A(new_n9813), .B(new_n9811), .Y(new_n9814));
  nand_5 g07466(.A(new_n9814), .B(new_n9809), .Y(new_n9815));
  nand_5 g07467(.A(new_n9815), .B(new_n9808), .Y(new_n9816));
  nand_5 g07468(.A(new_n9816), .B(new_n9802), .Y(new_n9817));
  nand_5 g07469(.A(new_n9817), .B(new_n9801), .Y(new_n9818));
  nand_5 g07470(.A(new_n9818), .B(new_n9796), .Y(new_n9819));
  nand_5 g07471(.A(new_n9819), .B(new_n9795), .Y(new_n9820));
  nand_5 g07472(.A(new_n9820), .B(new_n9790), .Y(new_n9821));
  nand_5 g07473(.A(new_n9821), .B(new_n9789), .Y(new_n9822));
  nand_5 g07474(.A(new_n9822), .B(new_n9784), .Y(new_n9823));
  nand_5 g07475(.A(new_n9823), .B(new_n9783_1), .Y(new_n9824));
  not_8  g07476(.A(new_n9824), .Y(new_n9825));
  nand_5 g07477(.A(new_n9754), .B(new_n9752), .Y(new_n9826));
  nand_5 g07478(.A(new_n9826), .B(new_n9753_1), .Y(new_n9827));
  nand_5 g07479(.A(new_n6863_1), .B(n24327), .Y(new_n9828));
  nand_5 g07480(.A(new_n6864), .B(new_n5514), .Y(new_n9829));
  nand_5 g07481(.A(new_n9829), .B(new_n9828), .Y(new_n9830));
  xor_4  g07482(.A(new_n9830), .B(new_n9827), .Y(new_n9831));
  nand_5 g07483(.A(new_n9780), .B(new_n9777), .Y(new_n9832_1));
  nand_5 g07484(.A(new_n9832_1), .B(new_n9779), .Y(new_n9833_1));
  not_8  g07485(.A(n25119), .Y(new_n9834));
  nand_5 g07486(.A(new_n3071), .B(new_n9834), .Y(new_n9835));
  nand_5 g07487(.A(new_n3115), .B(n25119), .Y(new_n9836));
  nand_5 g07488(.A(new_n9836), .B(new_n9835), .Y(new_n9837));
  xor_4  g07489(.A(new_n9837), .B(new_n9833_1), .Y(new_n9838_1));
  or_5   g07490(.A(new_n9838_1), .B(new_n9831), .Y(new_n9839));
  nand_5 g07491(.A(new_n9838_1), .B(new_n9831), .Y(new_n9840));
  nand_5 g07492(.A(new_n9840), .B(new_n9839), .Y(new_n9841));
  xor_4  g07493(.A(new_n9841), .B(new_n9825), .Y(n904));
  nand_5 g07494(.A(new_n7784), .B(new_n7741), .Y(new_n9843));
  nand_5 g07495(.A(n18962), .B(n10158), .Y(new_n9844));
  and_5  g07496(.A(new_n9844), .B(new_n9843), .Y(new_n9845));
  not_8  g07497(.A(new_n9845), .Y(new_n9846));
  nand_5 g07498(.A(new_n9846), .B(new_n3552), .Y(new_n9847));
  nand_5 g07499(.A(new_n9845), .B(n20794), .Y(new_n9848));
  nand_5 g07500(.A(n23333), .B(n18962), .Y(new_n9849));
  nand_5 g07501(.A(new_n9849), .B(new_n9848), .Y(new_n9850));
  nand_5 g07502(.A(new_n9850), .B(new_n9847), .Y(new_n9851));
  not_8  g07503(.A(new_n9851), .Y(new_n9852));
  or_5   g07504(.A(new_n9843), .B(n8052), .Y(new_n9853));
  nand_5 g07505(.A(new_n9843), .B(n8052), .Y(new_n9854));
  and_5  g07506(.A(new_n9854), .B(new_n9853), .Y(new_n9855));
  not_8  g07507(.A(new_n9855), .Y(new_n9856));
  nand_5 g07508(.A(new_n9856), .B(new_n3548), .Y(new_n9857));
  nand_5 g07509(.A(new_n9855), .B(n14603), .Y(new_n9858));
  nand_5 g07510(.A(new_n9858), .B(new_n9857), .Y(new_n9859));
  xor_4  g07511(.A(new_n9859), .B(new_n9852), .Y(new_n9860));
  not_8  g07512(.A(new_n9860), .Y(new_n9861));
  nand_5 g07513(.A(new_n9861), .B(n24786), .Y(new_n9862));
  nand_5 g07514(.A(new_n9860), .B(new_n4596), .Y(new_n9863));
  nand_5 g07515(.A(new_n3654), .B(new_n7784), .Y(new_n9864));
  and_5  g07516(.A(new_n9864), .B(new_n9849), .Y(new_n9865));
  nand_5 g07517(.A(new_n9865), .B(n23065), .Y(new_n9866));
  not_8  g07518(.A(new_n9866), .Y(new_n9867_1));
  nand_5 g07519(.A(new_n9848), .B(new_n9847), .Y(new_n9868));
  not_8  g07520(.A(new_n9868), .Y(new_n9869));
  nand_5 g07521(.A(new_n9869), .B(new_n9867_1), .Y(new_n9870));
  nand_5 g07522(.A(new_n9869), .B(new_n9849), .Y(new_n9871));
  nor_5  g07523(.A(new_n9869), .B(new_n9849), .Y(new_n9872_1));
  nor_5  g07524(.A(new_n9872_1), .B(new_n9867_1), .Y(new_n9873));
  nand_5 g07525(.A(new_n9873), .B(new_n9871), .Y(new_n9874));
  nand_5 g07526(.A(new_n9874), .B(n27120), .Y(new_n9875));
  nand_5 g07527(.A(new_n9875), .B(new_n9870), .Y(new_n9876));
  nand_5 g07528(.A(new_n9876), .B(new_n9863), .Y(new_n9877));
  nand_5 g07529(.A(new_n9877), .B(new_n9862), .Y(new_n9878));
  not_8  g07530(.A(new_n9878), .Y(new_n9879));
  nand_5 g07531(.A(new_n9858), .B(new_n9851), .Y(new_n9880));
  nand_5 g07532(.A(new_n9880), .B(new_n9857), .Y(new_n9881));
  not_8  g07533(.A(new_n9881), .Y(new_n9882));
  nor_5  g07534(.A(new_n9853), .B(n15539), .Y(new_n9883));
  not_8  g07535(.A(new_n9883), .Y(new_n9884));
  nand_5 g07536(.A(new_n9853), .B(n15539), .Y(new_n9885));
  and_5  g07537(.A(new_n9885), .B(new_n9884), .Y(new_n9886));
  not_8  g07538(.A(new_n9886), .Y(new_n9887));
  nand_5 g07539(.A(new_n9887), .B(new_n3639), .Y(new_n9888));
  nand_5 g07540(.A(new_n9886), .B(n18737), .Y(new_n9889));
  nand_5 g07541(.A(new_n9889), .B(new_n9888), .Y(new_n9890_1));
  xor_4  g07542(.A(new_n9890_1), .B(new_n9882), .Y(new_n9891));
  not_8  g07543(.A(new_n9891), .Y(new_n9892));
  nand_5 g07544(.A(new_n9892), .B(n25370), .Y(new_n9893));
  nand_5 g07545(.A(new_n9891), .B(new_n7825), .Y(new_n9894));
  nand_5 g07546(.A(new_n9894), .B(new_n9893), .Y(new_n9895));
  xor_4  g07547(.A(new_n9895), .B(new_n9879), .Y(new_n9896));
  or_5   g07548(.A(new_n9896), .B(new_n7675), .Y(new_n9897));
  not_8  g07549(.A(new_n9897), .Y(new_n9898));
  nand_5 g07550(.A(new_n9896), .B(new_n7675), .Y(new_n9899));
  not_8  g07551(.A(new_n9899), .Y(new_n9900));
  and_5  g07552(.A(new_n9874), .B(new_n9870), .Y(new_n9901));
  xor_4  g07553(.A(new_n9901), .B(new_n4553), .Y(new_n9902));
  nand_5 g07554(.A(new_n9902), .B(new_n7664), .Y(new_n9903));
  or_5   g07555(.A(new_n9902), .B(new_n7664), .Y(new_n9904));
  nor_5  g07556(.A(new_n9865), .B(n23065), .Y(new_n9905));
  nor_5  g07557(.A(new_n9905), .B(new_n9867_1), .Y(new_n9906));
  nand_5 g07558(.A(new_n9906), .B(new_n7656), .Y(new_n9907));
  nand_5 g07559(.A(new_n9907), .B(new_n9904), .Y(new_n9908));
  nand_5 g07560(.A(new_n9908), .B(new_n9903), .Y(new_n9909));
  nand_5 g07561(.A(new_n9909), .B(new_n7651), .Y(new_n9910));
  not_8  g07562(.A(new_n9910), .Y(new_n9911));
  nor_5  g07563(.A(new_n9909), .B(new_n7651), .Y(new_n9912));
  nand_5 g07564(.A(new_n9863), .B(new_n9862), .Y(new_n9913));
  xor_4  g07565(.A(new_n9913), .B(new_n9876), .Y(new_n9914));
  not_8  g07566(.A(new_n9914), .Y(new_n9915));
  nor_5  g07567(.A(new_n9915), .B(new_n9912), .Y(new_n9916));
  nor_5  g07568(.A(new_n9916), .B(new_n9911), .Y(new_n9917_1));
  nor_5  g07569(.A(new_n9917_1), .B(new_n9900), .Y(new_n9918));
  nor_5  g07570(.A(new_n9918), .B(new_n9898), .Y(new_n9919_1));
  not_8  g07571(.A(new_n9919_1), .Y(new_n9920));
  nand_5 g07572(.A(new_n9894), .B(new_n9878), .Y(new_n9921));
  nand_5 g07573(.A(new_n9921), .B(new_n9893), .Y(new_n9922));
  not_8  g07574(.A(new_n9922), .Y(new_n9923));
  nand_5 g07575(.A(new_n9889), .B(new_n9881), .Y(new_n9924));
  nand_5 g07576(.A(new_n9924), .B(new_n9888), .Y(new_n9925));
  not_8  g07577(.A(new_n9925), .Y(new_n9926_1));
  nand_5 g07578(.A(new_n9883), .B(new_n7732), .Y(new_n9927));
  nand_5 g07579(.A(new_n9884), .B(n19228), .Y(new_n9928));
  and_5  g07580(.A(new_n9928), .B(new_n9927), .Y(new_n9929));
  not_8  g07581(.A(new_n9929), .Y(new_n9930));
  nand_5 g07582(.A(new_n9930), .B(new_n3567), .Y(new_n9931));
  nand_5 g07583(.A(new_n9929), .B(n21471), .Y(new_n9932));
  nand_5 g07584(.A(new_n9932), .B(new_n9931), .Y(new_n9933));
  xor_4  g07585(.A(new_n9933), .B(new_n9926_1), .Y(new_n9934_1));
  nand_5 g07586(.A(new_n9934_1), .B(new_n7822), .Y(new_n9935));
  or_5   g07587(.A(new_n9934_1), .B(new_n7822), .Y(new_n9936));
  nand_5 g07588(.A(new_n9936), .B(new_n9935), .Y(new_n9937));
  xor_4  g07589(.A(new_n9937), .B(new_n9923), .Y(new_n9938_1));
  or_5   g07590(.A(new_n9938_1), .B(new_n7716), .Y(new_n9939));
  nand_5 g07591(.A(new_n9938_1), .B(new_n7716), .Y(new_n9940));
  nand_5 g07592(.A(new_n9940), .B(new_n9939), .Y(new_n9941));
  xor_4  g07593(.A(new_n9941), .B(new_n9920), .Y(n948));
  not_8  g07594(.A(n25972), .Y(new_n9943));
  nand_5 g07595(.A(new_n9943), .B(n10250), .Y(new_n9944));
  nand_5 g07596(.A(n25972), .B(new_n7040), .Y(new_n9945));
  nand_5 g07597(.A(new_n9945), .B(new_n9944), .Y(new_n9946_1));
  nand_5 g07598(.A(n21915), .B(new_n6991), .Y(new_n9947));
  nand_5 g07599(.A(new_n7974), .B(n7674), .Y(new_n9948));
  nand_5 g07600(.A(n13775), .B(new_n6997), .Y(new_n9949));
  nand_5 g07601(.A(new_n7882), .B(n6397), .Y(new_n9950));
  nand_5 g07602(.A(new_n7003), .B(n1293), .Y(new_n9951));
  nand_5 g07603(.A(n19196), .B(new_n7838), .Y(new_n9952));
  nand_5 g07604(.A(new_n7118), .B(n19042), .Y(new_n9953));
  nand_5 g07605(.A(n23586), .B(new_n7819), .Y(new_n9954));
  nand_5 g07606(.A(new_n7009), .B(n19472), .Y(new_n9955));
  nand_5 g07607(.A(n21226), .B(new_n7822), .Y(new_n9956));
  nand_5 g07608(.A(n25370), .B(new_n7012), .Y(new_n9957));
  nand_5 g07609(.A(new_n7825), .B(n4426), .Y(new_n9958));
  nand_5 g07610(.A(n24786), .B(new_n4606), .Y(new_n9959));
  nand_5 g07611(.A(new_n4596), .B(n20036), .Y(new_n9960));
  nand_5 g07612(.A(n27120), .B(new_n4561), .Y(new_n9961));
  nand_5 g07613(.A(new_n4553), .B(n11192), .Y(new_n9962));
  nand_5 g07614(.A(new_n4542), .B(n9380), .Y(new_n9963));
  nand_5 g07615(.A(new_n9963), .B(new_n9962), .Y(new_n9964));
  nand_5 g07616(.A(new_n9964), .B(new_n9961), .Y(new_n9965));
  nand_5 g07617(.A(new_n9965), .B(new_n9960), .Y(new_n9966));
  nand_5 g07618(.A(new_n9966), .B(new_n9959), .Y(new_n9967_1));
  nand_5 g07619(.A(new_n9967_1), .B(new_n9958), .Y(new_n9968_1));
  nand_5 g07620(.A(new_n9968_1), .B(new_n9957), .Y(new_n9969));
  nand_5 g07621(.A(new_n9969), .B(new_n9956), .Y(new_n9970));
  nand_5 g07622(.A(new_n9970), .B(new_n9955), .Y(new_n9971));
  nand_5 g07623(.A(new_n9971), .B(new_n9954), .Y(new_n9972));
  nand_5 g07624(.A(new_n9972), .B(new_n9953), .Y(new_n9973));
  nand_5 g07625(.A(new_n9973), .B(new_n9952), .Y(new_n9974));
  nand_5 g07626(.A(new_n9974), .B(new_n9951), .Y(new_n9975));
  nand_5 g07627(.A(new_n9975), .B(new_n9950), .Y(new_n9976));
  nand_5 g07628(.A(new_n9976), .B(new_n9949), .Y(new_n9977));
  nand_5 g07629(.A(new_n9977), .B(new_n9948), .Y(new_n9978));
  nand_5 g07630(.A(new_n9978), .B(new_n9947), .Y(new_n9979));
  xnor_4 g07631(.A(new_n9979), .B(new_n9946_1), .Y(new_n9980));
  not_8  g07632(.A(n15258), .Y(new_n9981));
  nand_5 g07633(.A(new_n9981), .B(new_n2611), .Y(new_n9982));
  or_5   g07634(.A(new_n9982), .B(n16743), .Y(new_n9983));
  nor_5  g07635(.A(new_n9983), .B(n22631), .Y(new_n9984));
  nand_5 g07636(.A(new_n9984), .B(new_n9181), .Y(new_n9985));
  nor_5  g07637(.A(new_n9985), .B(n25068), .Y(new_n9986));
  nand_5 g07638(.A(new_n9986), .B(new_n9169), .Y(new_n9987));
  nor_5  g07639(.A(new_n9987), .B(n7841), .Y(new_n9988));
  nand_5 g07640(.A(new_n9988), .B(new_n9157), .Y(new_n9989));
  not_8  g07641(.A(new_n9989), .Y(new_n9990));
  nor_5  g07642(.A(new_n9988), .B(new_n9157), .Y(new_n9991));
  nor_5  g07643(.A(new_n9991), .B(new_n9990), .Y(new_n9992));
  or_5   g07644(.A(new_n9992), .B(n15077), .Y(new_n9993));
  nand_5 g07645(.A(new_n9992), .B(n15077), .Y(new_n9994));
  xor_4  g07646(.A(new_n9987), .B(n7841), .Y(new_n9995));
  or_5   g07647(.A(new_n9995), .B(n3710), .Y(new_n9996));
  nand_5 g07648(.A(new_n9995), .B(n3710), .Y(new_n9997));
  xor_4  g07649(.A(new_n9986), .B(new_n9169), .Y(new_n9998));
  or_5   g07650(.A(new_n9998), .B(n26318), .Y(new_n9999));
  nand_5 g07651(.A(new_n9998), .B(n26318), .Y(new_n10000));
  xor_4  g07652(.A(new_n9985), .B(n25068), .Y(new_n10001));
  or_5   g07653(.A(new_n10001), .B(n26054), .Y(new_n10002));
  nand_5 g07654(.A(new_n10001), .B(n26054), .Y(new_n10003));
  xor_4  g07655(.A(new_n9984), .B(new_n9181), .Y(new_n10004));
  or_5   g07656(.A(new_n10004), .B(n19081), .Y(new_n10005));
  nand_5 g07657(.A(new_n10004), .B(n19081), .Y(new_n10006));
  xor_4  g07658(.A(new_n9983), .B(n22631), .Y(new_n10007));
  or_5   g07659(.A(new_n10007), .B(n8309), .Y(new_n10008));
  nand_5 g07660(.A(new_n10007), .B(n8309), .Y(new_n10009_1));
  nand_5 g07661(.A(new_n9982), .B(n16743), .Y(new_n10010_1));
  and_5  g07662(.A(new_n10010_1), .B(new_n9983), .Y(new_n10011));
  or_5   g07663(.A(new_n10011), .B(n19144), .Y(new_n10012));
  nand_5 g07664(.A(new_n10011), .B(n19144), .Y(new_n10013));
  nand_5 g07665(.A(n15258), .B(n4588), .Y(new_n10014));
  and_5  g07666(.A(new_n10014), .B(new_n9982), .Y(new_n10015));
  or_5   g07667(.A(new_n10015), .B(n12593), .Y(new_n10016));
  nand_5 g07668(.A(n13714), .B(n4588), .Y(new_n10017_1));
  nand_5 g07669(.A(new_n10015), .B(n12593), .Y(new_n10018_1));
  nand_5 g07670(.A(new_n10018_1), .B(new_n10017_1), .Y(new_n10019_1));
  nand_5 g07671(.A(new_n10019_1), .B(new_n10016), .Y(new_n10020));
  nand_5 g07672(.A(new_n10020), .B(new_n10013), .Y(new_n10021_1));
  nand_5 g07673(.A(new_n10021_1), .B(new_n10012), .Y(new_n10022));
  nand_5 g07674(.A(new_n10022), .B(new_n10009_1), .Y(new_n10023));
  nand_5 g07675(.A(new_n10023), .B(new_n10008), .Y(new_n10024));
  nand_5 g07676(.A(new_n10024), .B(new_n10006), .Y(new_n10025));
  nand_5 g07677(.A(new_n10025), .B(new_n10005), .Y(new_n10026));
  nand_5 g07678(.A(new_n10026), .B(new_n10003), .Y(new_n10027));
  nand_5 g07679(.A(new_n10027), .B(new_n10002), .Y(new_n10028));
  nand_5 g07680(.A(new_n10028), .B(new_n10000), .Y(new_n10029));
  nand_5 g07681(.A(new_n10029), .B(new_n9999), .Y(new_n10030));
  nand_5 g07682(.A(new_n10030), .B(new_n9997), .Y(new_n10031));
  nand_5 g07683(.A(new_n10031), .B(new_n9996), .Y(new_n10032));
  nand_5 g07684(.A(new_n10032), .B(new_n9994), .Y(new_n10033));
  nand_5 g07685(.A(new_n10033), .B(new_n9993), .Y(new_n10034));
  xor_4  g07686(.A(new_n9989), .B(n22764), .Y(new_n10035));
  xor_4  g07687(.A(new_n10035), .B(n12507), .Y(new_n10036));
  xor_4  g07688(.A(new_n10036), .B(new_n10034), .Y(new_n10037));
  nand_5 g07689(.A(n20040), .B(new_n8648), .Y(new_n10038));
  nand_5 g07690(.A(new_n2648), .B(n2978), .Y(new_n10039));
  nand_5 g07691(.A(new_n10039), .B(new_n10038), .Y(new_n10040));
  nand_5 g07692(.A(n23697), .B(new_n2652), .Y(new_n10041));
  nand_5 g07693(.A(new_n7958), .B(n19531), .Y(new_n10042));
  not_8  g07694(.A(n18345), .Y(new_n10043));
  nand_5 g07695(.A(new_n10043), .B(n2289), .Y(new_n10044));
  nand_5 g07696(.A(n18345), .B(new_n7810), .Y(new_n10045));
  nand_5 g07697(.A(new_n2658), .B(n1112), .Y(new_n10046));
  nand_5 g07698(.A(n13190), .B(new_n7757), .Y(new_n10047));
  not_8  g07699(.A(n3460), .Y(new_n10048));
  nand_5 g07700(.A(n20179), .B(new_n10048), .Y(new_n10049));
  nand_5 g07701(.A(new_n7729), .B(n3460), .Y(new_n10050));
  nand_5 g07702(.A(n19228), .B(new_n2663), .Y(new_n10051));
  nand_5 g07703(.A(new_n7732), .B(n5226), .Y(new_n10052));
  not_8  g07704(.A(n17664), .Y(new_n10053_1));
  nand_5 g07705(.A(new_n10053_1), .B(n15539), .Y(new_n10054));
  nand_5 g07706(.A(n17664), .B(new_n7735), .Y(new_n10055_1));
  nand_5 g07707(.A(new_n2669), .B(n8052), .Y(new_n10056));
  nand_5 g07708(.A(n23369), .B(new_n7738), .Y(new_n10057_1));
  nand_5 g07709(.A(n10158), .B(new_n2673), .Y(new_n10058));
  nand_5 g07710(.A(new_n7741), .B(n1136), .Y(new_n10059));
  nand_5 g07711(.A(n19234), .B(new_n7784), .Y(new_n10060));
  nand_5 g07712(.A(new_n10060), .B(new_n10059), .Y(new_n10061));
  nand_5 g07713(.A(new_n10061), .B(new_n10058), .Y(new_n10062));
  nand_5 g07714(.A(new_n10062), .B(new_n10057_1), .Y(new_n10063));
  nand_5 g07715(.A(new_n10063), .B(new_n10056), .Y(new_n10064));
  nand_5 g07716(.A(new_n10064), .B(new_n10055_1), .Y(new_n10065));
  nand_5 g07717(.A(new_n10065), .B(new_n10054), .Y(new_n10066));
  nand_5 g07718(.A(new_n10066), .B(new_n10052), .Y(new_n10067));
  nand_5 g07719(.A(new_n10067), .B(new_n10051), .Y(new_n10068));
  nand_5 g07720(.A(new_n10068), .B(new_n10050), .Y(new_n10069));
  nand_5 g07721(.A(new_n10069), .B(new_n10049), .Y(new_n10070));
  nand_5 g07722(.A(new_n10070), .B(new_n10047), .Y(new_n10071));
  nand_5 g07723(.A(new_n10071), .B(new_n10046), .Y(new_n10072));
  nand_5 g07724(.A(new_n10072), .B(new_n10045), .Y(new_n10073));
  nand_5 g07725(.A(new_n10073), .B(new_n10044), .Y(new_n10074));
  nand_5 g07726(.A(new_n10074), .B(new_n10042), .Y(new_n10075));
  nand_5 g07727(.A(new_n10075), .B(new_n10041), .Y(new_n10076));
  not_8  g07728(.A(new_n10076), .Y(new_n10077));
  xor_4  g07729(.A(new_n10077), .B(new_n10040), .Y(new_n10078));
  not_8  g07730(.A(new_n10078), .Y(new_n10079));
  or_5   g07731(.A(new_n10079), .B(new_n10037), .Y(new_n10080));
  nand_5 g07732(.A(new_n10079), .B(new_n10037), .Y(new_n10081));
  nand_5 g07733(.A(new_n10081), .B(new_n10080), .Y(new_n10082));
  nand_5 g07734(.A(new_n9994), .B(new_n9993), .Y(new_n10083));
  xor_4  g07735(.A(new_n10083), .B(new_n10032), .Y(new_n10084));
  nand_5 g07736(.A(new_n10042), .B(new_n10041), .Y(new_n10085));
  xor_4  g07737(.A(new_n10085), .B(new_n10074), .Y(new_n10086));
  not_8  g07738(.A(new_n10086), .Y(new_n10087));
  nand_5 g07739(.A(new_n10087), .B(new_n10084), .Y(new_n10088));
  or_5   g07740(.A(new_n10087), .B(new_n10084), .Y(new_n10089));
  nand_5 g07741(.A(new_n10045), .B(new_n10044), .Y(new_n10090));
  xor_4  g07742(.A(new_n10090), .B(new_n10072), .Y(new_n10091));
  not_8  g07743(.A(new_n10091), .Y(new_n10092));
  nand_5 g07744(.A(new_n9997), .B(new_n9996), .Y(new_n10093));
  xor_4  g07745(.A(new_n10093), .B(new_n10030), .Y(new_n10094));
  nand_5 g07746(.A(new_n10094), .B(new_n10092), .Y(new_n10095));
  nor_5  g07747(.A(new_n10094), .B(new_n10092), .Y(new_n10096_1));
  not_8  g07748(.A(new_n10096_1), .Y(new_n10097));
  nand_5 g07749(.A(new_n10047), .B(new_n10046), .Y(new_n10098));
  xor_4  g07750(.A(new_n10098), .B(new_n10070), .Y(new_n10099));
  not_8  g07751(.A(new_n10099), .Y(new_n10100));
  nand_5 g07752(.A(new_n10000), .B(new_n9999), .Y(new_n10101_1));
  xor_4  g07753(.A(new_n10101_1), .B(new_n10028), .Y(new_n10102));
  nand_5 g07754(.A(new_n10102), .B(new_n10100), .Y(new_n10103));
  nor_5  g07755(.A(new_n10102), .B(new_n10100), .Y(new_n10104));
  not_8  g07756(.A(new_n10104), .Y(new_n10105));
  nand_5 g07757(.A(new_n10050), .B(new_n10049), .Y(new_n10106));
  xor_4  g07758(.A(new_n10106), .B(new_n10068), .Y(new_n10107));
  not_8  g07759(.A(new_n10107), .Y(new_n10108));
  nand_5 g07760(.A(new_n10003), .B(new_n10002), .Y(new_n10109));
  xor_4  g07761(.A(new_n10109), .B(new_n10026), .Y(new_n10110));
  nand_5 g07762(.A(new_n10110), .B(new_n10108), .Y(new_n10111_1));
  nor_5  g07763(.A(new_n10110), .B(new_n10108), .Y(new_n10112));
  not_8  g07764(.A(new_n10112), .Y(new_n10113));
  nand_5 g07765(.A(new_n10052), .B(new_n10051), .Y(new_n10114));
  xor_4  g07766(.A(new_n10114), .B(new_n10066), .Y(new_n10115));
  not_8  g07767(.A(new_n10115), .Y(new_n10116));
  nand_5 g07768(.A(new_n10006), .B(new_n10005), .Y(new_n10117_1));
  xor_4  g07769(.A(new_n10117_1), .B(new_n10024), .Y(new_n10118));
  nand_5 g07770(.A(new_n10118), .B(new_n10116), .Y(new_n10119));
  nor_5  g07771(.A(new_n10118), .B(new_n10116), .Y(new_n10120));
  nand_5 g07772(.A(new_n10055_1), .B(new_n10054), .Y(new_n10121));
  xor_4  g07773(.A(new_n10121), .B(new_n10064), .Y(new_n10122));
  not_8  g07774(.A(new_n10122), .Y(new_n10123));
  nand_5 g07775(.A(new_n10009_1), .B(new_n10008), .Y(new_n10124));
  xor_4  g07776(.A(new_n10124), .B(new_n10022), .Y(new_n10125_1));
  or_5   g07777(.A(new_n10125_1), .B(new_n10123), .Y(new_n10126));
  nand_5 g07778(.A(new_n10125_1), .B(new_n10123), .Y(new_n10127));
  nand_5 g07779(.A(new_n10057_1), .B(new_n10056), .Y(new_n10128));
  xor_4  g07780(.A(new_n10128), .B(new_n10062), .Y(new_n10129));
  not_8  g07781(.A(new_n10129), .Y(new_n10130));
  nand_5 g07782(.A(new_n10013), .B(new_n10012), .Y(new_n10131));
  xor_4  g07783(.A(new_n10131), .B(new_n10020), .Y(new_n10132));
  nand_5 g07784(.A(new_n10132), .B(new_n10130), .Y(new_n10133));
  or_5   g07785(.A(new_n10132), .B(new_n10130), .Y(new_n10134));
  nand_5 g07786(.A(new_n2744), .B(n18962), .Y(new_n10135));
  and_5  g07787(.A(new_n10135), .B(new_n10060), .Y(new_n10136));
  not_8  g07788(.A(new_n10136), .Y(new_n10137));
  not_8  g07789(.A(n13714), .Y(new_n10138));
  nand_5 g07790(.A(new_n10138), .B(new_n2611), .Y(new_n10139));
  and_5  g07791(.A(new_n10139), .B(new_n10017_1), .Y(new_n10140));
  nand_5 g07792(.A(new_n10140), .B(new_n10137), .Y(new_n10141));
  nand_5 g07793(.A(new_n10059), .B(new_n10058), .Y(new_n10142));
  xnor_4 g07794(.A(new_n10142), .B(new_n10060), .Y(new_n10143));
  not_8  g07795(.A(new_n10143), .Y(new_n10144));
  or_5   g07796(.A(new_n10144), .B(new_n10141), .Y(new_n10145));
  nand_5 g07797(.A(new_n10144), .B(new_n10141), .Y(new_n10146));
  nand_5 g07798(.A(new_n10018_1), .B(new_n10016), .Y(new_n10147));
  xnor_4 g07799(.A(new_n10147), .B(new_n10017_1), .Y(new_n10148));
  not_8  g07800(.A(new_n10148), .Y(new_n10149));
  nand_5 g07801(.A(new_n10149), .B(new_n10146), .Y(new_n10150));
  nand_5 g07802(.A(new_n10150), .B(new_n10145), .Y(new_n10151));
  nand_5 g07803(.A(new_n10151), .B(new_n10134), .Y(new_n10152));
  nand_5 g07804(.A(new_n10152), .B(new_n10133), .Y(new_n10153));
  not_8  g07805(.A(new_n10153), .Y(new_n10154));
  nand_5 g07806(.A(new_n10154), .B(new_n10127), .Y(new_n10155));
  nand_5 g07807(.A(new_n10155), .B(new_n10126), .Y(new_n10156));
  or_5   g07808(.A(new_n10156), .B(new_n10120), .Y(new_n10157));
  nand_5 g07809(.A(new_n10157), .B(new_n10119), .Y(new_n10158_1));
  nand_5 g07810(.A(new_n10158_1), .B(new_n10113), .Y(new_n10159));
  nand_5 g07811(.A(new_n10159), .B(new_n10111_1), .Y(new_n10160));
  nand_5 g07812(.A(new_n10160), .B(new_n10105), .Y(new_n10161));
  nand_5 g07813(.A(new_n10161), .B(new_n10103), .Y(new_n10162));
  nand_5 g07814(.A(new_n10162), .B(new_n10097), .Y(new_n10163));
  nand_5 g07815(.A(new_n10163), .B(new_n10095), .Y(new_n10164));
  nand_5 g07816(.A(new_n10164), .B(new_n10089), .Y(new_n10165_1));
  nand_5 g07817(.A(new_n10165_1), .B(new_n10088), .Y(new_n10166));
  xnor_4 g07818(.A(new_n10166), .B(new_n10082), .Y(new_n10167));
  nand_5 g07819(.A(new_n10167), .B(new_n9980), .Y(new_n10168));
  or_5   g07820(.A(new_n10167), .B(new_n9980), .Y(new_n10169));
  nand_5 g07821(.A(new_n10169), .B(new_n10168), .Y(new_n10170));
  nand_5 g07822(.A(new_n9948), .B(new_n9947), .Y(new_n10171));
  xor_4  g07823(.A(new_n10171), .B(new_n9977), .Y(new_n10172));
  nand_5 g07824(.A(new_n10089), .B(new_n10088), .Y(new_n10173));
  xor_4  g07825(.A(new_n10173), .B(new_n10164), .Y(new_n10174));
  nand_5 g07826(.A(new_n10174), .B(new_n10172), .Y(new_n10175));
  not_8  g07827(.A(new_n10175), .Y(new_n10176));
  nor_5  g07828(.A(new_n10174), .B(new_n10172), .Y(new_n10177));
  nand_5 g07829(.A(new_n9950), .B(new_n9949), .Y(new_n10178));
  xor_4  g07830(.A(new_n10178), .B(new_n9975), .Y(new_n10179));
  nand_5 g07831(.A(new_n10097), .B(new_n10095), .Y(new_n10180));
  xor_4  g07832(.A(new_n10180), .B(new_n10162), .Y(new_n10181));
  nand_5 g07833(.A(new_n10181), .B(new_n10179), .Y(new_n10182));
  not_8  g07834(.A(new_n10182), .Y(new_n10183));
  nor_5  g07835(.A(new_n10181), .B(new_n10179), .Y(new_n10184));
  nand_5 g07836(.A(new_n9952), .B(new_n9951), .Y(new_n10185));
  xor_4  g07837(.A(new_n10185), .B(new_n9973), .Y(new_n10186));
  nand_5 g07838(.A(new_n10105), .B(new_n10103), .Y(new_n10187));
  xor_4  g07839(.A(new_n10187), .B(new_n10160), .Y(new_n10188));
  nand_5 g07840(.A(new_n10188), .B(new_n10186), .Y(new_n10189));
  not_8  g07841(.A(new_n10189), .Y(new_n10190));
  nor_5  g07842(.A(new_n10188), .B(new_n10186), .Y(new_n10191));
  nand_5 g07843(.A(new_n9954), .B(new_n9953), .Y(new_n10192));
  xor_4  g07844(.A(new_n10192), .B(new_n9971), .Y(new_n10193));
  nand_5 g07845(.A(new_n10113), .B(new_n10111_1), .Y(new_n10194));
  xor_4  g07846(.A(new_n10194), .B(new_n10158_1), .Y(new_n10195));
  nand_5 g07847(.A(new_n10195), .B(new_n10193), .Y(new_n10196));
  not_8  g07848(.A(new_n10196), .Y(new_n10197));
  nor_5  g07849(.A(new_n10195), .B(new_n10193), .Y(new_n10198));
  nand_5 g07850(.A(new_n9956), .B(new_n9955), .Y(new_n10199));
  xor_4  g07851(.A(new_n10199), .B(new_n9969), .Y(new_n10200));
  not_8  g07852(.A(new_n10120), .Y(new_n10201_1));
  nand_5 g07853(.A(new_n10201_1), .B(new_n10119), .Y(new_n10202));
  xor_4  g07854(.A(new_n10202), .B(new_n10156), .Y(new_n10203));
  not_8  g07855(.A(new_n10203), .Y(new_n10204));
  nand_5 g07856(.A(new_n10204), .B(new_n10200), .Y(new_n10205));
  not_8  g07857(.A(new_n10205), .Y(new_n10206));
  nor_5  g07858(.A(new_n10204), .B(new_n10200), .Y(new_n10207));
  nand_5 g07859(.A(new_n9958), .B(new_n9957), .Y(new_n10208));
  xor_4  g07860(.A(new_n10208), .B(new_n9967_1), .Y(new_n10209));
  nand_5 g07861(.A(new_n10127), .B(new_n10126), .Y(new_n10210));
  xor_4  g07862(.A(new_n10210), .B(new_n10153), .Y(new_n10211));
  or_5   g07863(.A(new_n10211), .B(new_n10209), .Y(new_n10212));
  nand_5 g07864(.A(new_n10211), .B(new_n10209), .Y(new_n10213));
  nand_5 g07865(.A(new_n9960), .B(new_n9959), .Y(new_n10214));
  xor_4  g07866(.A(new_n10214), .B(new_n9965), .Y(new_n10215));
  nand_5 g07867(.A(new_n10133), .B(new_n10134), .Y(new_n10216));
  xor_4  g07868(.A(new_n10216), .B(new_n10151), .Y(new_n10217));
  or_5   g07869(.A(new_n10217), .B(new_n10215), .Y(new_n10218));
  nand_5 g07870(.A(new_n10217), .B(new_n10215), .Y(new_n10219));
  xor_4  g07871(.A(n23065), .B(new_n4545), .Y(new_n10220));
  not_8  g07872(.A(new_n10220), .Y(new_n10221));
  not_8  g07873(.A(new_n10141), .Y(new_n10222));
  nor_5  g07874(.A(new_n10140), .B(new_n10137), .Y(new_n10223));
  nor_5  g07875(.A(new_n10223), .B(new_n10222), .Y(new_n10224));
  nand_5 g07876(.A(new_n10224), .B(new_n10221), .Y(new_n10225));
  not_8  g07877(.A(new_n10225), .Y(new_n10226));
  nand_5 g07878(.A(new_n9962), .B(new_n9961), .Y(new_n10227));
  xnor_4 g07879(.A(new_n10227), .B(new_n9963), .Y(new_n10228));
  nand_5 g07880(.A(new_n10228), .B(new_n10226), .Y(new_n10229));
  not_8  g07881(.A(new_n10229), .Y(new_n10230));
  nor_5  g07882(.A(new_n10228), .B(new_n10226), .Y(new_n10231));
  nand_5 g07883(.A(new_n10145), .B(new_n10146), .Y(new_n10232));
  xor_4  g07884(.A(new_n10232), .B(new_n10149), .Y(new_n10233));
  nor_5  g07885(.A(new_n10233), .B(new_n10231), .Y(new_n10234));
  nor_5  g07886(.A(new_n10234), .B(new_n10230), .Y(new_n10235));
  not_8  g07887(.A(new_n10235), .Y(new_n10236_1));
  nand_5 g07888(.A(new_n10236_1), .B(new_n10219), .Y(new_n10237));
  nand_5 g07889(.A(new_n10237), .B(new_n10218), .Y(new_n10238));
  nand_5 g07890(.A(new_n10238), .B(new_n10213), .Y(new_n10239_1));
  nand_5 g07891(.A(new_n10239_1), .B(new_n10212), .Y(new_n10240));
  nor_5  g07892(.A(new_n10240), .B(new_n10207), .Y(new_n10241));
  nor_5  g07893(.A(new_n10241), .B(new_n10206), .Y(new_n10242));
  nor_5  g07894(.A(new_n10242), .B(new_n10198), .Y(new_n10243));
  nor_5  g07895(.A(new_n10243), .B(new_n10197), .Y(new_n10244_1));
  nor_5  g07896(.A(new_n10244_1), .B(new_n10191), .Y(new_n10245));
  nor_5  g07897(.A(new_n10245), .B(new_n10190), .Y(new_n10246));
  nor_5  g07898(.A(new_n10246), .B(new_n10184), .Y(new_n10247));
  nor_5  g07899(.A(new_n10247), .B(new_n10183), .Y(new_n10248));
  nor_5  g07900(.A(new_n10248), .B(new_n10177), .Y(new_n10249));
  nor_5  g07901(.A(new_n10249), .B(new_n10176), .Y(new_n10250_1));
  not_8  g07902(.A(new_n10250_1), .Y(new_n10251));
  xor_4  g07903(.A(new_n10251), .B(new_n10170), .Y(n957));
  nand_5 g07904(.A(new_n10137), .B(n20385), .Y(new_n10253));
  not_8  g07905(.A(new_n10253), .Y(new_n10254));
  nor_5  g07906(.A(new_n10137), .B(n20385), .Y(new_n10255));
  or_5   g07907(.A(new_n10255), .B(new_n10254), .Y(new_n10256));
  not_8  g07908(.A(new_n10256), .Y(new_n10257));
  nand_5 g07909(.A(n26167), .B(n24129), .Y(new_n10258));
  not_8  g07910(.A(new_n10258), .Y(new_n10259));
  nor_5  g07911(.A(n26167), .B(n24129), .Y(new_n10260));
  nor_5  g07912(.A(new_n10260), .B(new_n10259), .Y(new_n10261_1));
  not_8  g07913(.A(new_n10261_1), .Y(new_n10262_1));
  nand_5 g07914(.A(new_n10262_1), .B(n21138), .Y(new_n10263));
  nand_5 g07915(.A(new_n10261_1), .B(new_n8276_1), .Y(new_n10264));
  nand_5 g07916(.A(new_n10264), .B(new_n10263), .Y(new_n10265));
  nand_5 g07917(.A(new_n10265), .B(new_n10257), .Y(new_n10266));
  not_8  g07918(.A(new_n10266), .Y(new_n10267));
  nor_5  g07919(.A(new_n10265), .B(new_n10257), .Y(new_n10268));
  nor_5  g07920(.A(new_n10268), .B(new_n10267), .Y(n980));
  xor_4  g07921(.A(new_n8841), .B(new_n4849), .Y(new_n10270));
  nand_5 g07922(.A(new_n8847), .B(new_n4852), .Y(new_n10271));
  not_8  g07923(.A(new_n8847), .Y(new_n10272));
  nand_5 g07924(.A(new_n10272), .B(new_n4854), .Y(new_n10273));
  nand_5 g07925(.A(new_n8853), .B(new_n4858_1), .Y(new_n10274));
  nand_5 g07926(.A(new_n8857), .B(new_n4860), .Y(new_n10275_1));
  nand_5 g07927(.A(new_n8861_1), .B(new_n4864), .Y(new_n10276));
  nand_5 g07928(.A(new_n8865), .B(new_n4866), .Y(new_n10277));
  nand_5 g07929(.A(new_n8869_1), .B(new_n4870), .Y(new_n10278));
  nand_5 g07930(.A(new_n8873), .B(new_n4872), .Y(new_n10279));
  nand_5 g07931(.A(new_n8877), .B(new_n4876), .Y(new_n10280));
  nand_5 g07932(.A(new_n8881), .B(new_n4878), .Y(new_n10281));
  nand_5 g07933(.A(new_n8885), .B(new_n4882), .Y(new_n10282));
  nand_5 g07934(.A(new_n8889), .B(new_n4884), .Y(new_n10283));
  nand_5 g07935(.A(new_n8893), .B(new_n4888), .Y(new_n10284));
  nand_5 g07936(.A(new_n8897), .B(new_n4890), .Y(new_n10285));
  nand_5 g07937(.A(new_n8901), .B(new_n4894), .Y(new_n10286));
  nand_5 g07938(.A(new_n8905), .B(new_n4896), .Y(new_n10287_1));
  nand_5 g07939(.A(new_n8910), .B(new_n4901), .Y(new_n10288));
  nand_5 g07940(.A(new_n8909_1), .B(new_n4900), .Y(new_n10289));
  nand_5 g07941(.A(new_n8917), .B(new_n4906), .Y(new_n10290));
  nand_5 g07942(.A(new_n10290), .B(new_n10289), .Y(new_n10291));
  nand_5 g07943(.A(new_n10291), .B(new_n10288), .Y(new_n10292));
  nand_5 g07944(.A(new_n10292), .B(new_n10287_1), .Y(new_n10293));
  nand_5 g07945(.A(new_n10293), .B(new_n10286), .Y(new_n10294));
  nand_5 g07946(.A(new_n10294), .B(new_n10285), .Y(new_n10295_1));
  nand_5 g07947(.A(new_n10295_1), .B(new_n10284), .Y(new_n10296));
  nand_5 g07948(.A(new_n10296), .B(new_n10283), .Y(new_n10297));
  nand_5 g07949(.A(new_n10297), .B(new_n10282), .Y(new_n10298));
  nand_5 g07950(.A(new_n10298), .B(new_n10281), .Y(new_n10299));
  nand_5 g07951(.A(new_n10299), .B(new_n10280), .Y(new_n10300));
  nand_5 g07952(.A(new_n10300), .B(new_n10279), .Y(new_n10301));
  nand_5 g07953(.A(new_n10301), .B(new_n10278), .Y(new_n10302));
  nand_5 g07954(.A(new_n10302), .B(new_n10277), .Y(new_n10303));
  nand_5 g07955(.A(new_n10303), .B(new_n10276), .Y(new_n10304));
  nand_5 g07956(.A(new_n10304), .B(new_n10275_1), .Y(new_n10305));
  nand_5 g07957(.A(new_n10305), .B(new_n10274), .Y(new_n10306));
  nand_5 g07958(.A(new_n10306), .B(new_n10273), .Y(new_n10307));
  nand_5 g07959(.A(new_n10307), .B(new_n10271), .Y(new_n10308));
  nor_5  g07960(.A(new_n10308), .B(new_n10270), .Y(new_n10309));
  not_8  g07961(.A(new_n10309), .Y(new_n10310));
  nand_5 g07962(.A(new_n10308), .B(new_n10270), .Y(new_n10311));
  and_5  g07963(.A(new_n10311), .B(new_n10310), .Y(new_n10312));
  not_8  g07964(.A(new_n10312), .Y(new_n10313));
  not_8  g07965(.A(n12650), .Y(new_n10314));
  nand_5 g07966(.A(n16544), .B(new_n10314), .Y(new_n10315));
  not_8  g07967(.A(n16544), .Y(new_n10316));
  nand_5 g07968(.A(new_n10316), .B(n12650), .Y(new_n10317));
  not_8  g07969(.A(n10201), .Y(new_n10318));
  nand_5 g07970(.A(new_n10318), .B(n6814), .Y(new_n10319));
  nand_5 g07971(.A(n10201), .B(new_n3286), .Y(new_n10320));
  not_8  g07972(.A(n10593), .Y(new_n10321_1));
  nand_5 g07973(.A(n19701), .B(new_n10321_1), .Y(new_n10322));
  nand_5 g07974(.A(new_n3186), .B(n10593), .Y(new_n10323));
  not_8  g07975(.A(n18290), .Y(new_n10324));
  nand_5 g07976(.A(n23529), .B(new_n10324), .Y(new_n10325));
  nand_5 g07977(.A(new_n3068), .B(n18290), .Y(new_n10326_1));
  not_8  g07978(.A(n11580), .Y(new_n10327_1));
  nand_5 g07979(.A(n24620), .B(new_n10327_1), .Y(new_n10328));
  nand_5 g07980(.A(new_n3035), .B(n11580), .Y(new_n10329));
  not_8  g07981(.A(n15884), .Y(new_n10330_1));
  nand_5 g07982(.A(new_n10330_1), .B(n5211), .Y(new_n10331));
  nand_5 g07983(.A(n15884), .B(new_n3038), .Y(new_n10332));
  not_8  g07984(.A(n6356), .Y(new_n10333));
  nand_5 g07985(.A(n12956), .B(new_n10333), .Y(new_n10334));
  nand_5 g07986(.A(new_n3043), .B(n6356), .Y(new_n10335));
  nand_5 g07987(.A(new_n6205), .B(n18295), .Y(new_n10336));
  nand_5 g07988(.A(n27104), .B(new_n3046), .Y(new_n10337));
  not_8  g07989(.A(n27188), .Y(new_n10338));
  nand_5 g07990(.A(new_n10338), .B(n6502), .Y(new_n10339));
  nand_5 g07991(.A(n27188), .B(new_n3051), .Y(new_n10340_1));
  nand_5 g07992(.A(new_n3159), .B(n6611), .Y(new_n10341));
  nand_5 g07993(.A(new_n10341), .B(new_n10340_1), .Y(new_n10342));
  nand_5 g07994(.A(new_n10342), .B(new_n10339), .Y(new_n10343));
  nand_5 g07995(.A(new_n10343), .B(new_n10337), .Y(new_n10344));
  nand_5 g07996(.A(new_n10344), .B(new_n10336), .Y(new_n10345_1));
  nand_5 g07997(.A(new_n10345_1), .B(new_n10335), .Y(new_n10346));
  nand_5 g07998(.A(new_n10346), .B(new_n10334), .Y(new_n10347));
  nand_5 g07999(.A(new_n10347), .B(new_n10332), .Y(new_n10348));
  nand_5 g08000(.A(new_n10348), .B(new_n10331), .Y(new_n10349));
  nand_5 g08001(.A(new_n10349), .B(new_n10329), .Y(new_n10350));
  nand_5 g08002(.A(new_n10350), .B(new_n10328), .Y(new_n10351));
  nand_5 g08003(.A(new_n10351), .B(new_n10326_1), .Y(new_n10352));
  nand_5 g08004(.A(new_n10352), .B(new_n10325), .Y(new_n10353));
  nand_5 g08005(.A(new_n10353), .B(new_n10323), .Y(new_n10354));
  nand_5 g08006(.A(new_n10354), .B(new_n10322), .Y(new_n10355));
  nand_5 g08007(.A(new_n10355), .B(new_n10320), .Y(new_n10356_1));
  nand_5 g08008(.A(new_n10356_1), .B(new_n10319), .Y(new_n10357));
  nand_5 g08009(.A(new_n10357), .B(new_n10317), .Y(new_n10358));
  nand_5 g08010(.A(new_n10358), .B(new_n10315), .Y(new_n10359));
  nor_5  g08011(.A(new_n10359), .B(new_n10313), .Y(new_n10360));
  not_8  g08012(.A(new_n10359), .Y(new_n10361));
  nor_5  g08013(.A(new_n10361), .B(new_n10312), .Y(new_n10362));
  or_5   g08014(.A(new_n10362), .B(new_n10360), .Y(new_n10363));
  nand_5 g08015(.A(new_n10273), .B(new_n10271), .Y(new_n10364));
  xor_4  g08016(.A(new_n10364), .B(new_n10306), .Y(new_n10365));
  not_8  g08017(.A(new_n10365), .Y(new_n10366));
  nand_5 g08018(.A(new_n10317), .B(new_n10315), .Y(new_n10367));
  xor_4  g08019(.A(new_n10367), .B(new_n10357), .Y(new_n10368));
  nand_5 g08020(.A(new_n10368), .B(new_n10366), .Y(new_n10369));
  or_5   g08021(.A(new_n10368), .B(new_n10366), .Y(new_n10370));
  nand_5 g08022(.A(new_n10275_1), .B(new_n10274), .Y(new_n10371));
  xor_4  g08023(.A(new_n10371), .B(new_n10304), .Y(new_n10372_1));
  not_8  g08024(.A(new_n10372_1), .Y(new_n10373));
  nand_5 g08025(.A(new_n10320), .B(new_n10319), .Y(new_n10374));
  xor_4  g08026(.A(new_n10374), .B(new_n10355), .Y(new_n10375));
  nand_5 g08027(.A(new_n10375), .B(new_n10373), .Y(new_n10376));
  or_5   g08028(.A(new_n10375), .B(new_n10373), .Y(new_n10377));
  nand_5 g08029(.A(new_n10277), .B(new_n10276), .Y(new_n10378));
  xor_4  g08030(.A(new_n10378), .B(new_n10302), .Y(new_n10379));
  not_8  g08031(.A(new_n10379), .Y(new_n10380));
  nand_5 g08032(.A(new_n10323), .B(new_n10322), .Y(new_n10381));
  xor_4  g08033(.A(new_n10381), .B(new_n10353), .Y(new_n10382));
  nand_5 g08034(.A(new_n10382), .B(new_n10380), .Y(new_n10383));
  or_5   g08035(.A(new_n10382), .B(new_n10380), .Y(new_n10384));
  nand_5 g08036(.A(new_n10279), .B(new_n10278), .Y(new_n10385_1));
  xor_4  g08037(.A(new_n10385_1), .B(new_n10300), .Y(new_n10386));
  nand_5 g08038(.A(new_n10326_1), .B(new_n10325), .Y(new_n10387_1));
  xor_4  g08039(.A(new_n10387_1), .B(new_n10351), .Y(new_n10388_1));
  not_8  g08040(.A(new_n10388_1), .Y(new_n10389));
  or_5   g08041(.A(new_n10389), .B(new_n10386), .Y(new_n10390_1));
  nand_5 g08042(.A(new_n10389), .B(new_n10386), .Y(new_n10391));
  nand_5 g08043(.A(new_n10281), .B(new_n10280), .Y(new_n10392));
  xor_4  g08044(.A(new_n10392), .B(new_n10298), .Y(new_n10393));
  not_8  g08045(.A(new_n10393), .Y(new_n10394));
  nand_5 g08046(.A(new_n10329), .B(new_n10328), .Y(new_n10395));
  xor_4  g08047(.A(new_n10395), .B(new_n10349), .Y(new_n10396));
  nand_5 g08048(.A(new_n10396), .B(new_n10394), .Y(new_n10397));
  or_5   g08049(.A(new_n10396), .B(new_n10394), .Y(new_n10398));
  nand_5 g08050(.A(new_n10283), .B(new_n10282), .Y(new_n10399));
  xor_4  g08051(.A(new_n10399), .B(new_n10296), .Y(new_n10400));
  not_8  g08052(.A(new_n10400), .Y(new_n10401));
  nand_5 g08053(.A(new_n10332), .B(new_n10331), .Y(new_n10402));
  xor_4  g08054(.A(new_n10402), .B(new_n10347), .Y(new_n10403));
  nand_5 g08055(.A(new_n10403), .B(new_n10401), .Y(new_n10404_1));
  or_5   g08056(.A(new_n10403), .B(new_n10401), .Y(new_n10405_1));
  nand_5 g08057(.A(new_n10285), .B(new_n10284), .Y(new_n10406));
  xor_4  g08058(.A(new_n10406), .B(new_n10294), .Y(new_n10407));
  not_8  g08059(.A(new_n10407), .Y(new_n10408));
  nand_5 g08060(.A(new_n10335), .B(new_n10334), .Y(new_n10409_1));
  xor_4  g08061(.A(new_n10409_1), .B(new_n10345_1), .Y(new_n10410));
  nand_5 g08062(.A(new_n10410), .B(new_n10408), .Y(new_n10411_1));
  or_5   g08063(.A(new_n10410), .B(new_n10408), .Y(new_n10412));
  nand_5 g08064(.A(new_n10287_1), .B(new_n10286), .Y(new_n10413));
  xor_4  g08065(.A(new_n10413), .B(new_n10292), .Y(new_n10414));
  not_8  g08066(.A(new_n10414), .Y(new_n10415));
  nand_5 g08067(.A(new_n10337), .B(new_n10336), .Y(new_n10416));
  xor_4  g08068(.A(new_n10416), .B(new_n10343), .Y(new_n10417));
  nand_5 g08069(.A(new_n10417), .B(new_n10415), .Y(new_n10418));
  or_5   g08070(.A(new_n10417), .B(new_n10415), .Y(new_n10419));
  not_8  g08071(.A(new_n10290), .Y(new_n10420_1));
  nor_5  g08072(.A(new_n8917), .B(new_n4906), .Y(new_n10421));
  nor_5  g08073(.A(new_n10421), .B(new_n10420_1), .Y(new_n10422));
  not_8  g08074(.A(new_n10422), .Y(new_n10423));
  xor_4  g08075(.A(n15780), .B(new_n6339_1), .Y(new_n10424));
  nor_5  g08076(.A(new_n10424), .B(new_n10423), .Y(new_n10425));
  nand_5 g08077(.A(new_n10340_1), .B(new_n10339), .Y(new_n10426));
  xnor_4 g08078(.A(new_n10426), .B(new_n10341), .Y(new_n10427));
  nand_5 g08079(.A(new_n10427), .B(new_n10425), .Y(new_n10428));
  not_8  g08080(.A(new_n10428), .Y(new_n10429));
  nand_5 g08081(.A(new_n10289), .B(new_n10288), .Y(new_n10430));
  xor_4  g08082(.A(new_n10430), .B(new_n10290), .Y(new_n10431));
  not_8  g08083(.A(new_n10431), .Y(new_n10432_1));
  nor_5  g08084(.A(new_n10427), .B(new_n10425), .Y(new_n10433));
  nor_5  g08085(.A(new_n10433), .B(new_n10432_1), .Y(new_n10434));
  nor_5  g08086(.A(new_n10434), .B(new_n10429), .Y(new_n10435));
  nand_5 g08087(.A(new_n10435), .B(new_n10419), .Y(new_n10436));
  and_5  g08088(.A(new_n10436), .B(new_n10418), .Y(new_n10437));
  not_8  g08089(.A(new_n10437), .Y(new_n10438));
  nand_5 g08090(.A(new_n10438), .B(new_n10412), .Y(new_n10439));
  nand_5 g08091(.A(new_n10439), .B(new_n10411_1), .Y(new_n10440));
  nand_5 g08092(.A(new_n10440), .B(new_n10405_1), .Y(new_n10441));
  nand_5 g08093(.A(new_n10441), .B(new_n10404_1), .Y(new_n10442));
  nand_5 g08094(.A(new_n10442), .B(new_n10398), .Y(new_n10443));
  nand_5 g08095(.A(new_n10443), .B(new_n10397), .Y(new_n10444));
  nand_5 g08096(.A(new_n10444), .B(new_n10391), .Y(new_n10445));
  nand_5 g08097(.A(new_n10445), .B(new_n10390_1), .Y(new_n10446));
  nand_5 g08098(.A(new_n10446), .B(new_n10384), .Y(new_n10447));
  nand_5 g08099(.A(new_n10447), .B(new_n10383), .Y(new_n10448));
  nand_5 g08100(.A(new_n10448), .B(new_n10377), .Y(new_n10449));
  nand_5 g08101(.A(new_n10449), .B(new_n10376), .Y(new_n10450));
  nand_5 g08102(.A(new_n10450), .B(new_n10370), .Y(new_n10451));
  nand_5 g08103(.A(new_n10451), .B(new_n10369), .Y(new_n10452));
  xor_4  g08104(.A(new_n10452), .B(new_n10363), .Y(n982));
  not_8  g08105(.A(n3279), .Y(new_n10454));
  not_8  g08106(.A(n14702), .Y(new_n10455));
  not_8  g08107(.A(n2547), .Y(new_n10456));
  not_8  g08108(.A(n7339), .Y(new_n10457));
  not_8  g08109(.A(n26808), .Y(new_n10458));
  nand_5 g08110(.A(new_n10458), .B(new_n10457), .Y(new_n10459));
  or_5   g08111(.A(new_n10459), .B(n1667), .Y(new_n10460));
  nor_5  g08112(.A(new_n10460), .B(n2680), .Y(new_n10461));
  nand_5 g08113(.A(new_n10461), .B(new_n10456), .Y(new_n10462));
  nor_5  g08114(.A(new_n10462), .B(n2999), .Y(new_n10463));
  nand_5 g08115(.A(new_n10463), .B(new_n10455), .Y(new_n10464));
  nor_5  g08116(.A(new_n10464), .B(n13914), .Y(new_n10465));
  nand_5 g08117(.A(new_n10465), .B(new_n10454), .Y(new_n10466));
  xor_4  g08118(.A(new_n10466), .B(n4306), .Y(new_n10467));
  not_8  g08119(.A(n23166), .Y(new_n10468));
  nand_5 g08120(.A(new_n10468), .B(n18105), .Y(new_n10469));
  nand_5 g08121(.A(n23166), .B(new_n9229), .Y(new_n10470));
  nand_5 g08122(.A(new_n10470), .B(new_n10469), .Y(new_n10471));
  nand_5 g08123(.A(new_n4928), .B(n10577), .Y(new_n10472));
  not_8  g08124(.A(n10577), .Y(new_n10473));
  nand_5 g08125(.A(n24196), .B(new_n10473), .Y(new_n10474));
  nand_5 g08126(.A(new_n9233), .B(n6381), .Y(new_n10475));
  not_8  g08127(.A(n6381), .Y(new_n10476));
  nand_5 g08128(.A(n16376), .B(new_n10476), .Y(new_n10477));
  nand_5 g08129(.A(new_n4929), .B(n14345), .Y(new_n10478));
  not_8  g08130(.A(n14345), .Y(new_n10479));
  nand_5 g08131(.A(n25381), .B(new_n10479), .Y(new_n10480));
  nand_5 g08132(.A(new_n9239), .B(n11356), .Y(new_n10481));
  not_8  g08133(.A(n11356), .Y(new_n10482));
  nand_5 g08134(.A(n12587), .B(new_n10482), .Y(new_n10483));
  nand_5 g08135(.A(n3164), .B(new_n4930), .Y(new_n10484_1));
  not_8  g08136(.A(n3164), .Y(new_n10485));
  nand_5 g08137(.A(new_n10485), .B(n268), .Y(new_n10486));
  nand_5 g08138(.A(new_n9245), .B(n10611), .Y(new_n10487));
  nand_5 g08139(.A(n24879), .B(new_n7620), .Y(new_n10488));
  nand_5 g08140(.A(new_n9249), .B(n2783), .Y(new_n10489_1));
  nand_5 g08141(.A(n6785), .B(new_n7569_1), .Y(new_n10490));
  nand_5 g08142(.A(new_n4931), .B(n15490), .Y(new_n10491));
  nand_5 g08143(.A(n24032), .B(new_n7550), .Y(new_n10492));
  nand_5 g08144(.A(n22843), .B(new_n7558_1), .Y(new_n10493));
  nand_5 g08145(.A(new_n10493), .B(new_n10492), .Y(new_n10494));
  nand_5 g08146(.A(new_n10494), .B(new_n10491), .Y(new_n10495));
  nand_5 g08147(.A(new_n10495), .B(new_n10490), .Y(new_n10496));
  nand_5 g08148(.A(new_n10496), .B(new_n10489_1), .Y(new_n10497));
  nand_5 g08149(.A(new_n10497), .B(new_n10488), .Y(new_n10498));
  nand_5 g08150(.A(new_n10498), .B(new_n10487), .Y(new_n10499));
  nand_5 g08151(.A(new_n10499), .B(new_n10486), .Y(new_n10500));
  nand_5 g08152(.A(new_n10500), .B(new_n10484_1), .Y(new_n10501));
  nand_5 g08153(.A(new_n10501), .B(new_n10483), .Y(new_n10502));
  nand_5 g08154(.A(new_n10502), .B(new_n10481), .Y(new_n10503));
  nand_5 g08155(.A(new_n10503), .B(new_n10480), .Y(new_n10504));
  nand_5 g08156(.A(new_n10504), .B(new_n10478), .Y(new_n10505));
  nand_5 g08157(.A(new_n10505), .B(new_n10477), .Y(new_n10506));
  nand_5 g08158(.A(new_n10506), .B(new_n10475), .Y(new_n10507));
  nand_5 g08159(.A(new_n10507), .B(new_n10474), .Y(new_n10508));
  nand_5 g08160(.A(new_n10508), .B(new_n10472), .Y(new_n10509));
  not_8  g08161(.A(new_n10509), .Y(new_n10510));
  xor_4  g08162(.A(new_n10510), .B(new_n10471), .Y(new_n10511));
  nand_5 g08163(.A(new_n10511), .B(new_n10467), .Y(new_n10512));
  or_5   g08164(.A(new_n10511), .B(new_n10467), .Y(new_n10513));
  nand_5 g08165(.A(new_n10513), .B(new_n10512), .Y(new_n10514_1));
  xor_4  g08166(.A(new_n10465), .B(new_n10454), .Y(new_n10515));
  nand_5 g08167(.A(new_n10474), .B(new_n10472), .Y(new_n10516));
  xor_4  g08168(.A(new_n10516), .B(new_n10507), .Y(new_n10517));
  not_8  g08169(.A(new_n10517), .Y(new_n10518));
  or_5   g08170(.A(new_n10518), .B(new_n10515), .Y(new_n10519));
  nand_5 g08171(.A(new_n10518), .B(new_n10515), .Y(new_n10520));
  xor_4  g08172(.A(new_n10464), .B(n13914), .Y(new_n10521));
  nand_5 g08173(.A(new_n10477), .B(new_n10475), .Y(new_n10522));
  xor_4  g08174(.A(new_n10522), .B(new_n10505), .Y(new_n10523));
  not_8  g08175(.A(new_n10523), .Y(new_n10524));
  or_5   g08176(.A(new_n10524), .B(new_n10521), .Y(new_n10525_1));
  nand_5 g08177(.A(new_n10524), .B(new_n10521), .Y(new_n10526));
  xor_4  g08178(.A(new_n10463), .B(new_n10455), .Y(new_n10527));
  nand_5 g08179(.A(new_n10480), .B(new_n10478), .Y(new_n10528));
  xor_4  g08180(.A(new_n10528), .B(new_n10503), .Y(new_n10529));
  not_8  g08181(.A(new_n10529), .Y(new_n10530));
  or_5   g08182(.A(new_n10530), .B(new_n10527), .Y(new_n10531));
  nand_5 g08183(.A(new_n10530), .B(new_n10527), .Y(new_n10532));
  xor_4  g08184(.A(new_n10462), .B(n2999), .Y(new_n10533));
  nand_5 g08185(.A(new_n10483), .B(new_n10481), .Y(new_n10534));
  xor_4  g08186(.A(new_n10534), .B(new_n10501), .Y(new_n10535));
  not_8  g08187(.A(new_n10535), .Y(new_n10536));
  or_5   g08188(.A(new_n10536), .B(new_n10533), .Y(new_n10537));
  nand_5 g08189(.A(new_n10536), .B(new_n10533), .Y(new_n10538));
  xor_4  g08190(.A(new_n10461), .B(new_n10456), .Y(new_n10539));
  nand_5 g08191(.A(new_n10486), .B(new_n10484_1), .Y(new_n10540_1));
  xor_4  g08192(.A(new_n10540_1), .B(new_n10499), .Y(new_n10541));
  not_8  g08193(.A(new_n10541), .Y(new_n10542));
  or_5   g08194(.A(new_n10542), .B(new_n10539), .Y(new_n10543));
  nand_5 g08195(.A(new_n10542), .B(new_n10539), .Y(new_n10544));
  xor_4  g08196(.A(new_n10460), .B(n2680), .Y(new_n10545));
  nand_5 g08197(.A(new_n10488), .B(new_n10487), .Y(new_n10546));
  xor_4  g08198(.A(new_n10546), .B(new_n10497), .Y(new_n10547));
  not_8  g08199(.A(new_n10547), .Y(new_n10548));
  or_5   g08200(.A(new_n10548), .B(new_n10545), .Y(new_n10549));
  nand_5 g08201(.A(new_n10548), .B(new_n10545), .Y(new_n10550));
  nand_5 g08202(.A(new_n10459), .B(n1667), .Y(new_n10551));
  and_5  g08203(.A(new_n10551), .B(new_n10460), .Y(new_n10552));
  nand_5 g08204(.A(new_n10490), .B(new_n10489_1), .Y(new_n10553));
  xor_4  g08205(.A(new_n10553), .B(new_n10495), .Y(new_n10554));
  not_8  g08206(.A(new_n10554), .Y(new_n10555));
  or_5   g08207(.A(new_n10555), .B(new_n10552), .Y(new_n10556));
  nand_5 g08208(.A(new_n10555), .B(new_n10552), .Y(new_n10557));
  nand_5 g08209(.A(n26808), .B(n7339), .Y(new_n10558));
  and_5  g08210(.A(new_n10558), .B(new_n10459), .Y(new_n10559));
  and_5  g08211(.A(new_n10492), .B(new_n10491), .Y(new_n10560));
  xor_4  g08212(.A(new_n10560), .B(new_n10493), .Y(new_n10561_1));
  or_5   g08213(.A(new_n10561_1), .B(new_n10559), .Y(new_n10562));
  nand_5 g08214(.A(new_n10561_1), .B(new_n10559), .Y(new_n10563));
  nand_5 g08215(.A(new_n2622), .B(n18), .Y(new_n10564_1));
  and_5  g08216(.A(new_n10564_1), .B(new_n10493), .Y(new_n10565));
  not_8  g08217(.A(new_n10565), .Y(new_n10566));
  nand_5 g08218(.A(new_n10566), .B(n26808), .Y(new_n10567));
  nand_5 g08219(.A(new_n10567), .B(new_n10563), .Y(new_n10568));
  nand_5 g08220(.A(new_n10568), .B(new_n10562), .Y(new_n10569));
  nand_5 g08221(.A(new_n10569), .B(new_n10557), .Y(new_n10570));
  nand_5 g08222(.A(new_n10570), .B(new_n10556), .Y(new_n10571));
  nand_5 g08223(.A(new_n10571), .B(new_n10550), .Y(new_n10572));
  nand_5 g08224(.A(new_n10572), .B(new_n10549), .Y(new_n10573));
  nand_5 g08225(.A(new_n10573), .B(new_n10544), .Y(new_n10574));
  nand_5 g08226(.A(new_n10574), .B(new_n10543), .Y(new_n10575));
  nand_5 g08227(.A(new_n10575), .B(new_n10538), .Y(new_n10576));
  nand_5 g08228(.A(new_n10576), .B(new_n10537), .Y(new_n10577_1));
  nand_5 g08229(.A(new_n10577_1), .B(new_n10532), .Y(new_n10578));
  nand_5 g08230(.A(new_n10578), .B(new_n10531), .Y(new_n10579));
  nand_5 g08231(.A(new_n10579), .B(new_n10526), .Y(new_n10580));
  nand_5 g08232(.A(new_n10580), .B(new_n10525_1), .Y(new_n10581));
  nand_5 g08233(.A(new_n10581), .B(new_n10520), .Y(new_n10582));
  nand_5 g08234(.A(new_n10582), .B(new_n10519), .Y(new_n10583));
  not_8  g08235(.A(new_n10583), .Y(new_n10584));
  xor_4  g08236(.A(new_n10584), .B(new_n10514_1), .Y(new_n10585));
  not_8  g08237(.A(new_n10585), .Y(new_n10586));
  or_5   g08238(.A(new_n10586), .B(new_n5052), .Y(new_n10587));
  nand_5 g08239(.A(new_n10586), .B(new_n5052), .Y(new_n10588_1));
  nand_5 g08240(.A(new_n10588_1), .B(new_n10587), .Y(new_n10589));
  nand_5 g08241(.A(new_n10520), .B(new_n10519), .Y(new_n10590));
  xor_4  g08242(.A(new_n10590), .B(new_n10581), .Y(new_n10591));
  nand_5 g08243(.A(new_n10591), .B(new_n5059), .Y(new_n10592));
  nor_5  g08244(.A(new_n10591), .B(new_n5059), .Y(new_n10593_1));
  not_8  g08245(.A(new_n10593_1), .Y(new_n10594));
  nand_5 g08246(.A(new_n10526), .B(new_n10525_1), .Y(new_n10595_1));
  xor_4  g08247(.A(new_n10595_1), .B(new_n10579), .Y(new_n10596));
  nand_5 g08248(.A(new_n10596), .B(new_n5066), .Y(new_n10597));
  nor_5  g08249(.A(new_n10596), .B(new_n5066), .Y(new_n10598));
  not_8  g08250(.A(new_n10598), .Y(new_n10599));
  nand_5 g08251(.A(new_n10532), .B(new_n10531), .Y(new_n10600));
  xor_4  g08252(.A(new_n10600), .B(new_n10577_1), .Y(new_n10601));
  nand_5 g08253(.A(new_n10601), .B(new_n5073), .Y(new_n10602));
  or_5   g08254(.A(new_n10601), .B(new_n5073), .Y(new_n10603));
  nand_5 g08255(.A(new_n10538), .B(new_n10537), .Y(new_n10604));
  xor_4  g08256(.A(new_n10604), .B(new_n10575), .Y(new_n10605));
  nand_5 g08257(.A(new_n10605), .B(new_n5079), .Y(new_n10606));
  nor_5  g08258(.A(new_n10605), .B(new_n5079), .Y(new_n10607));
  not_8  g08259(.A(new_n10607), .Y(new_n10608));
  nand_5 g08260(.A(new_n10544), .B(new_n10543), .Y(new_n10609));
  xor_4  g08261(.A(new_n10609), .B(new_n10573), .Y(new_n10610));
  nand_5 g08262(.A(new_n10610), .B(new_n5085), .Y(new_n10611_1));
  nor_5  g08263(.A(new_n10610), .B(new_n5085), .Y(new_n10612));
  not_8  g08264(.A(new_n10612), .Y(new_n10613));
  nand_5 g08265(.A(new_n10550), .B(new_n10549), .Y(new_n10614_1));
  xor_4  g08266(.A(new_n10614_1), .B(new_n10571), .Y(new_n10615));
  nand_5 g08267(.A(new_n10615), .B(new_n5091), .Y(new_n10616));
  nor_5  g08268(.A(new_n10615), .B(new_n5091), .Y(new_n10617_1));
  not_8  g08269(.A(new_n10617_1), .Y(new_n10618));
  nand_5 g08270(.A(new_n10557), .B(new_n10556), .Y(new_n10619));
  xor_4  g08271(.A(new_n10619), .B(new_n10569), .Y(new_n10620));
  nand_5 g08272(.A(new_n10620), .B(new_n5097), .Y(new_n10621));
  nor_5  g08273(.A(new_n10620), .B(new_n5097), .Y(new_n10622));
  not_8  g08274(.A(new_n10622), .Y(new_n10623));
  nand_5 g08275(.A(new_n10563), .B(new_n10562), .Y(new_n10624));
  xor_4  g08276(.A(new_n10624), .B(new_n10567), .Y(new_n10625));
  nand_5 g08277(.A(new_n10625), .B(new_n5105), .Y(new_n10626));
  not_8  g08278(.A(new_n10625), .Y(new_n10627));
  nand_5 g08279(.A(new_n10627), .B(new_n5104), .Y(new_n10628_1));
  nand_5 g08280(.A(new_n10565), .B(new_n10458), .Y(new_n10629));
  nand_5 g08281(.A(new_n10629), .B(new_n10567), .Y(new_n10630));
  nor_5  g08282(.A(new_n10630), .B(new_n5112), .Y(new_n10631));
  nand_5 g08283(.A(new_n10631), .B(new_n10628_1), .Y(new_n10632));
  nand_5 g08284(.A(new_n10632), .B(new_n10626), .Y(new_n10633));
  nand_5 g08285(.A(new_n10633), .B(new_n10623), .Y(new_n10634));
  nand_5 g08286(.A(new_n10634), .B(new_n10621), .Y(new_n10635));
  nand_5 g08287(.A(new_n10635), .B(new_n10618), .Y(new_n10636));
  nand_5 g08288(.A(new_n10636), .B(new_n10616), .Y(new_n10637));
  nand_5 g08289(.A(new_n10637), .B(new_n10613), .Y(new_n10638));
  nand_5 g08290(.A(new_n10638), .B(new_n10611_1), .Y(new_n10639));
  nand_5 g08291(.A(new_n10639), .B(new_n10608), .Y(new_n10640));
  nand_5 g08292(.A(new_n10640), .B(new_n10606), .Y(new_n10641));
  nand_5 g08293(.A(new_n10641), .B(new_n10603), .Y(new_n10642));
  nand_5 g08294(.A(new_n10642), .B(new_n10602), .Y(new_n10643));
  nand_5 g08295(.A(new_n10643), .B(new_n10599), .Y(new_n10644));
  nand_5 g08296(.A(new_n10644), .B(new_n10597), .Y(new_n10645));
  nand_5 g08297(.A(new_n10645), .B(new_n10594), .Y(new_n10646));
  nand_5 g08298(.A(new_n10646), .B(new_n10592), .Y(new_n10647_1));
  xnor_4 g08299(.A(new_n10647_1), .B(new_n10589), .Y(n984));
  nand_5 g08300(.A(new_n10603), .B(new_n10602), .Y(new_n10649));
  xnor_4 g08301(.A(new_n10649), .B(new_n10641), .Y(n1005));
  nand_5 g08302(.A(new_n3618_1), .B(new_n3619), .Y(new_n10651));
  xnor_4 g08303(.A(new_n10651), .B(new_n3679_1), .Y(n1016));
  nand_5 g08304(.A(new_n4463), .B(new_n4462), .Y(new_n10653_1));
  xnor_4 g08305(.A(new_n10653_1), .B(new_n4481), .Y(n1020));
  nand_5 g08306(.A(new_n10333), .B(new_n3007), .Y(new_n10655));
  nand_5 g08307(.A(n6356), .B(n4665), .Y(new_n10656));
  nand_5 g08308(.A(new_n6205), .B(new_n3010_1), .Y(new_n10657));
  nand_5 g08309(.A(n27104), .B(n19005), .Y(new_n10658));
  nand_5 g08310(.A(new_n10338), .B(new_n3013), .Y(new_n10659));
  nand_5 g08311(.A(n27188), .B(n4326), .Y(new_n10660));
  nand_5 g08312(.A(n6611), .B(n5438), .Y(new_n10661));
  nand_5 g08313(.A(new_n10661), .B(new_n10660), .Y(new_n10662));
  nand_5 g08314(.A(new_n10662), .B(new_n10659), .Y(new_n10663));
  nand_5 g08315(.A(new_n10663), .B(new_n10658), .Y(new_n10664));
  nand_5 g08316(.A(new_n10664), .B(new_n10657), .Y(new_n10665));
  nand_5 g08317(.A(new_n10665), .B(new_n10656), .Y(new_n10666));
  nand_5 g08318(.A(new_n10666), .B(new_n10655), .Y(new_n10667));
  not_8  g08319(.A(new_n10667), .Y(new_n10668));
  nand_5 g08320(.A(new_n10668), .B(n5213), .Y(new_n10669));
  nand_5 g08321(.A(new_n10667), .B(new_n3004), .Y(new_n10670));
  and_5  g08322(.A(new_n10670), .B(new_n10669), .Y(new_n10671));
  xor_4  g08323(.A(new_n10671), .B(new_n10330_1), .Y(new_n10672));
  not_8  g08324(.A(new_n10672), .Y(new_n10673));
  nand_5 g08325(.A(new_n10673), .B(n5211), .Y(new_n10674));
  nand_5 g08326(.A(new_n10672), .B(new_n3038), .Y(new_n10675));
  nand_5 g08327(.A(new_n10656), .B(new_n10655), .Y(new_n10676));
  xor_4  g08328(.A(new_n10676), .B(new_n10665), .Y(new_n10677));
  nand_5 g08329(.A(new_n10677), .B(n12956), .Y(new_n10678));
  not_8  g08330(.A(new_n10677), .Y(new_n10679));
  nand_5 g08331(.A(new_n10679), .B(new_n3043), .Y(new_n10680));
  nand_5 g08332(.A(new_n10658), .B(new_n10657), .Y(new_n10681));
  xor_4  g08333(.A(new_n10681), .B(new_n10663), .Y(new_n10682));
  nand_5 g08334(.A(new_n10682), .B(n18295), .Y(new_n10683));
  not_8  g08335(.A(new_n10682), .Y(new_n10684));
  nand_5 g08336(.A(new_n10684), .B(new_n3046), .Y(new_n10685));
  nand_5 g08337(.A(new_n10660), .B(new_n10659), .Y(new_n10686));
  xor_4  g08338(.A(new_n10686), .B(new_n10661), .Y(new_n10687));
  nand_5 g08339(.A(new_n10687), .B(n6502), .Y(new_n10688));
  not_8  g08340(.A(new_n10687), .Y(new_n10689));
  nand_5 g08341(.A(new_n10689), .B(new_n3051), .Y(new_n10690));
  nand_5 g08342(.A(new_n6339_1), .B(new_n3015), .Y(new_n10691));
  and_5  g08343(.A(new_n10691), .B(new_n10661), .Y(new_n10692_1));
  nand_5 g08344(.A(new_n10692_1), .B(n15780), .Y(new_n10693));
  not_8  g08345(.A(new_n10693), .Y(new_n10694_1));
  nand_5 g08346(.A(new_n10694_1), .B(new_n10690), .Y(new_n10695));
  nand_5 g08347(.A(new_n10695), .B(new_n10688), .Y(new_n10696));
  nand_5 g08348(.A(new_n10696), .B(new_n10685), .Y(new_n10697));
  nand_5 g08349(.A(new_n10697), .B(new_n10683), .Y(new_n10698));
  nand_5 g08350(.A(new_n10698), .B(new_n10680), .Y(new_n10699));
  nand_5 g08351(.A(new_n10699), .B(new_n10678), .Y(new_n10700));
  nand_5 g08352(.A(new_n10700), .B(new_n10675), .Y(new_n10701_1));
  nand_5 g08353(.A(new_n10701_1), .B(new_n10674), .Y(new_n10702));
  nand_5 g08354(.A(new_n10669), .B(new_n10330_1), .Y(new_n10703));
  nand_5 g08355(.A(new_n10703), .B(new_n10670), .Y(new_n10704));
  not_8  g08356(.A(new_n10704), .Y(new_n10705));
  nand_5 g08357(.A(new_n10705), .B(n2035), .Y(new_n10706));
  nand_5 g08358(.A(new_n10704), .B(new_n3000), .Y(new_n10707));
  and_5  g08359(.A(new_n10707), .B(new_n10706), .Y(new_n10708));
  xor_4  g08360(.A(new_n10708), .B(new_n10327_1), .Y(new_n10709));
  not_8  g08361(.A(new_n10709), .Y(new_n10710_1));
  nand_5 g08362(.A(new_n10710_1), .B(n24620), .Y(new_n10711));
  nand_5 g08363(.A(new_n10709), .B(new_n3035), .Y(new_n10712_1));
  nand_5 g08364(.A(new_n10712_1), .B(new_n10711), .Y(new_n10713));
  xor_4  g08365(.A(new_n10713), .B(new_n10702), .Y(new_n10714));
  nand_5 g08366(.A(new_n6878), .B(new_n7605), .Y(new_n10715));
  nand_5 g08367(.A(n21276), .B(n11056), .Y(new_n10716));
  nand_5 g08368(.A(new_n6884), .B(new_n7539), .Y(new_n10717));
  nand_5 g08369(.A(n26748), .B(n15271), .Y(new_n10718));
  nand_5 g08370(.A(new_n6544), .B(new_n4654), .Y(new_n10719));
  nand_5 g08371(.A(n25877), .B(n10057), .Y(new_n10720));
  nand_5 g08372(.A(n24323), .B(n8920), .Y(new_n10721));
  nand_5 g08373(.A(new_n10721), .B(new_n10720), .Y(new_n10722));
  nand_5 g08374(.A(new_n10722), .B(new_n10719), .Y(new_n10723));
  nand_5 g08375(.A(new_n10723), .B(new_n10718), .Y(new_n10724));
  nand_5 g08376(.A(new_n10724), .B(new_n10717), .Y(new_n10725));
  nand_5 g08377(.A(new_n10725), .B(new_n10716), .Y(new_n10726));
  nand_5 g08378(.A(new_n10726), .B(new_n10715), .Y(new_n10727));
  not_8  g08379(.A(new_n10727), .Y(new_n10728));
  nand_5 g08380(.A(n16524), .B(n13668), .Y(new_n10729));
  nand_5 g08381(.A(new_n8813), .B(new_n4782), .Y(new_n10730));
  nand_5 g08382(.A(new_n10730), .B(new_n10729), .Y(new_n10731));
  xor_4  g08383(.A(new_n10731), .B(new_n10728), .Y(new_n10732));
  nand_5 g08384(.A(new_n10732), .B(new_n6814_1), .Y(new_n10733));
  not_8  g08385(.A(new_n10732), .Y(new_n10734));
  nand_5 g08386(.A(new_n10734), .B(n987), .Y(new_n10735));
  nand_5 g08387(.A(new_n10716), .B(new_n10715), .Y(new_n10736));
  xor_4  g08388(.A(new_n10736), .B(new_n10725), .Y(new_n10737));
  not_8  g08389(.A(new_n10737), .Y(new_n10738));
  nand_5 g08390(.A(new_n10738), .B(new_n6817), .Y(new_n10739_1));
  nand_5 g08391(.A(new_n10737), .B(n20478), .Y(new_n10740));
  nand_5 g08392(.A(new_n10718), .B(new_n10717), .Y(new_n10741));
  xor_4  g08393(.A(new_n10741), .B(new_n10723), .Y(new_n10742));
  not_8  g08394(.A(new_n10742), .Y(new_n10743));
  nand_5 g08395(.A(new_n10743), .B(new_n6820), .Y(new_n10744));
  nand_5 g08396(.A(new_n10742), .B(n26882), .Y(new_n10745));
  not_8  g08397(.A(new_n10721), .Y(new_n10746));
  nand_5 g08398(.A(new_n10720), .B(new_n10719), .Y(new_n10747));
  xor_4  g08399(.A(new_n10747), .B(new_n10746), .Y(new_n10748));
  nand_5 g08400(.A(new_n10748), .B(new_n6823), .Y(new_n10749));
  not_8  g08401(.A(new_n10748), .Y(new_n10750));
  nand_5 g08402(.A(new_n10750), .B(n22619), .Y(new_n10751));
  nand_5 g08403(.A(new_n6537), .B(new_n4653), .Y(new_n10752));
  nand_5 g08404(.A(new_n10752), .B(new_n10721), .Y(new_n10753));
  not_8  g08405(.A(new_n10753), .Y(new_n10754));
  nand_5 g08406(.A(new_n10754), .B(n6775), .Y(new_n10755));
  nand_5 g08407(.A(new_n10755), .B(new_n10751), .Y(new_n10756_1));
  nand_5 g08408(.A(new_n10756_1), .B(new_n10749), .Y(new_n10757));
  nand_5 g08409(.A(new_n10757), .B(new_n10745), .Y(new_n10758));
  nand_5 g08410(.A(new_n10758), .B(new_n10744), .Y(new_n10759));
  nand_5 g08411(.A(new_n10759), .B(new_n10740), .Y(new_n10760));
  nand_5 g08412(.A(new_n10760), .B(new_n10739_1), .Y(new_n10761));
  nand_5 g08413(.A(new_n10761), .B(new_n10735), .Y(new_n10762));
  nand_5 g08414(.A(new_n10762), .B(new_n10733), .Y(new_n10763_1));
  nand_5 g08415(.A(new_n10729), .B(new_n10727), .Y(new_n10764));
  nand_5 g08416(.A(new_n10764), .B(new_n10730), .Y(new_n10765));
  not_8  g08417(.A(new_n10765), .Y(new_n10766));
  nand_5 g08418(.A(n23160), .B(n3570), .Y(new_n10767));
  nand_5 g08419(.A(new_n8810), .B(new_n6867_1), .Y(new_n10768));
  nand_5 g08420(.A(new_n10768), .B(new_n10767), .Y(new_n10769));
  xor_4  g08421(.A(new_n10769), .B(new_n10766), .Y(new_n10770));
  nand_5 g08422(.A(new_n10770), .B(new_n6811), .Y(new_n10771));
  not_8  g08423(.A(new_n10770), .Y(new_n10772));
  nand_5 g08424(.A(new_n10772), .B(n2421), .Y(new_n10773));
  nand_5 g08425(.A(new_n10773), .B(new_n10771), .Y(new_n10774));
  xor_4  g08426(.A(new_n10774), .B(new_n10763_1), .Y(new_n10775_1));
  or_5   g08427(.A(new_n10775_1), .B(new_n10714), .Y(new_n10776));
  nand_5 g08428(.A(new_n10775_1), .B(new_n10714), .Y(new_n10777));
  nand_5 g08429(.A(new_n10733), .B(new_n10735), .Y(new_n10778));
  xor_4  g08430(.A(new_n10778), .B(new_n10761), .Y(new_n10779));
  nand_5 g08431(.A(new_n10674), .B(new_n10675), .Y(new_n10780_1));
  xor_4  g08432(.A(new_n10780_1), .B(new_n10700), .Y(new_n10781));
  or_5   g08433(.A(new_n10781), .B(new_n10779), .Y(new_n10782));
  nand_5 g08434(.A(new_n10781), .B(new_n10779), .Y(new_n10783));
  nand_5 g08435(.A(new_n10678), .B(new_n10680), .Y(new_n10784));
  xor_4  g08436(.A(new_n10784), .B(new_n10698), .Y(new_n10785));
  nand_5 g08437(.A(new_n10739_1), .B(new_n10740), .Y(new_n10786));
  xor_4  g08438(.A(new_n10786), .B(new_n10759), .Y(new_n10787));
  or_5   g08439(.A(new_n10787), .B(new_n10785), .Y(new_n10788));
  nand_5 g08440(.A(new_n10787), .B(new_n10785), .Y(new_n10789));
  nand_5 g08441(.A(new_n10683), .B(new_n10685), .Y(new_n10790));
  xor_4  g08442(.A(new_n10790), .B(new_n10696), .Y(new_n10791));
  nand_5 g08443(.A(new_n10744), .B(new_n10745), .Y(new_n10792_1));
  xor_4  g08444(.A(new_n10792_1), .B(new_n10757), .Y(new_n10793));
  or_5   g08445(.A(new_n10793), .B(new_n10791), .Y(new_n10794));
  nand_5 g08446(.A(new_n10793), .B(new_n10791), .Y(new_n10795));
  nand_5 g08447(.A(new_n10749), .B(new_n10751), .Y(new_n10796));
  xor_4  g08448(.A(new_n10796), .B(new_n10755), .Y(new_n10797));
  nand_5 g08449(.A(new_n10688), .B(new_n10690), .Y(new_n10798));
  xor_4  g08450(.A(new_n10798), .B(new_n10694_1), .Y(new_n10799));
  or_5   g08451(.A(new_n10799), .B(new_n10797), .Y(new_n10800));
  nand_5 g08452(.A(new_n10799), .B(new_n10797), .Y(new_n10801));
  nand_5 g08453(.A(new_n10753), .B(new_n6561), .Y(new_n10802));
  and_5  g08454(.A(new_n10802), .B(new_n10755), .Y(new_n10803));
  not_8  g08455(.A(new_n10692_1), .Y(new_n10804));
  nand_5 g08456(.A(new_n10804), .B(new_n3159), .Y(new_n10805));
  nand_5 g08457(.A(new_n10805), .B(new_n10693), .Y(new_n10806));
  nand_5 g08458(.A(new_n10806), .B(new_n10803), .Y(new_n10807));
  nand_5 g08459(.A(new_n10807), .B(new_n10801), .Y(new_n10808));
  nand_5 g08460(.A(new_n10808), .B(new_n10800), .Y(new_n10809));
  nand_5 g08461(.A(new_n10809), .B(new_n10795), .Y(new_n10810));
  nand_5 g08462(.A(new_n10810), .B(new_n10794), .Y(new_n10811));
  nand_5 g08463(.A(new_n10811), .B(new_n10789), .Y(new_n10812));
  nand_5 g08464(.A(new_n10812), .B(new_n10788), .Y(new_n10813));
  nand_5 g08465(.A(new_n10813), .B(new_n10783), .Y(new_n10814));
  nand_5 g08466(.A(new_n10814), .B(new_n10782), .Y(new_n10815));
  nand_5 g08467(.A(new_n10815), .B(new_n10777), .Y(new_n10816));
  nand_5 g08468(.A(new_n10816), .B(new_n10776), .Y(new_n10817_1));
  nand_5 g08469(.A(new_n10712_1), .B(new_n10702), .Y(new_n10818));
  nand_5 g08470(.A(new_n10818), .B(new_n10711), .Y(new_n10819));
  not_8  g08471(.A(new_n10819), .Y(new_n10820));
  nand_5 g08472(.A(new_n10706), .B(new_n10327_1), .Y(new_n10821));
  nand_5 g08473(.A(new_n10821), .B(new_n10707), .Y(new_n10822));
  nand_5 g08474(.A(new_n10324), .B(new_n2997), .Y(new_n10823));
  nand_5 g08475(.A(n18290), .B(n12875), .Y(new_n10824));
  nand_5 g08476(.A(new_n10824), .B(new_n10823), .Y(new_n10825));
  xor_4  g08477(.A(new_n10825), .B(new_n10822), .Y(new_n10826));
  nand_5 g08478(.A(new_n10826), .B(n23529), .Y(new_n10827));
  not_8  g08479(.A(new_n10826), .Y(new_n10828));
  nand_5 g08480(.A(new_n10828), .B(new_n3068), .Y(new_n10829));
  nand_5 g08481(.A(new_n10829), .B(new_n10827), .Y(new_n10830));
  xor_4  g08482(.A(new_n10830), .B(new_n10820), .Y(new_n10831));
  nand_5 g08483(.A(new_n10773), .B(new_n10763_1), .Y(new_n10832));
  nand_5 g08484(.A(new_n10832), .B(new_n10771), .Y(new_n10833));
  nand_5 g08485(.A(new_n10767), .B(new_n10765), .Y(new_n10834_1));
  nand_5 g08486(.A(new_n10834_1), .B(new_n10768), .Y(new_n10835));
  not_8  g08487(.A(new_n10835), .Y(new_n10836));
  nand_5 g08488(.A(new_n8807), .B(new_n6861_1), .Y(new_n10837));
  nand_5 g08489(.A(n17250), .B(n4409), .Y(new_n10838));
  nand_5 g08490(.A(new_n10838), .B(new_n10837), .Y(new_n10839));
  xor_4  g08491(.A(new_n10839), .B(new_n10836), .Y(new_n10840));
  nand_5 g08492(.A(new_n10840), .B(new_n6808), .Y(new_n10841));
  not_8  g08493(.A(new_n10840), .Y(new_n10842));
  nand_5 g08494(.A(new_n10842), .B(n11044), .Y(new_n10843));
  nand_5 g08495(.A(new_n10843), .B(new_n10841), .Y(new_n10844));
  xor_4  g08496(.A(new_n10844), .B(new_n10833), .Y(new_n10845));
  not_8  g08497(.A(new_n10845), .Y(new_n10846));
  nand_5 g08498(.A(new_n10846), .B(new_n10831), .Y(new_n10847));
  not_8  g08499(.A(new_n10831), .Y(new_n10848));
  nand_5 g08500(.A(new_n10845), .B(new_n10848), .Y(new_n10849));
  nand_5 g08501(.A(new_n10849), .B(new_n10847), .Y(new_n10850));
  xnor_4 g08502(.A(new_n10850), .B(new_n10817_1), .Y(n1044));
  nand_5 g08503(.A(n6775), .B(n3925), .Y(new_n10852));
  nand_5 g08504(.A(new_n6823), .B(new_n6561), .Y(new_n10853));
  nand_5 g08505(.A(n22619), .B(n6775), .Y(new_n10854));
  and_5  g08506(.A(new_n10854), .B(new_n10853), .Y(new_n10855));
  nand_5 g08507(.A(new_n10855), .B(n20259), .Y(new_n10856));
  or_5   g08508(.A(new_n10855), .B(n20259), .Y(new_n10857));
  nand_5 g08509(.A(new_n10857), .B(new_n10856), .Y(new_n10858));
  xor_4  g08510(.A(new_n10858), .B(new_n10852), .Y(new_n10859));
  nand_5 g08511(.A(new_n10859), .B(new_n6534), .Y(new_n10860));
  nand_5 g08512(.A(new_n10858), .B(new_n6533), .Y(new_n10861));
  nand_5 g08513(.A(new_n6561), .B(new_n5549), .Y(new_n10862));
  and_5  g08514(.A(new_n10862), .B(new_n10852), .Y(new_n10863));
  nand_5 g08515(.A(new_n10863), .B(new_n6536), .Y(new_n10864));
  not_8  g08516(.A(new_n10864), .Y(new_n10865));
  nand_5 g08517(.A(new_n10865), .B(new_n10861), .Y(new_n10866));
  nand_5 g08518(.A(new_n10866), .B(new_n10860), .Y(new_n10867));
  nand_5 g08519(.A(new_n6531), .B(new_n6525), .Y(new_n10868));
  nand_5 g08520(.A(new_n10868), .B(new_n6530), .Y(new_n10869));
  not_8  g08521(.A(new_n10869), .Y(new_n10870));
  or_5   g08522(.A(new_n6526), .B(n16396), .Y(new_n10871));
  nand_5 g08523(.A(new_n6526), .B(n16396), .Y(new_n10872));
  and_5  g08524(.A(new_n10872), .B(new_n10871), .Y(new_n10873));
  not_8  g08525(.A(new_n10873), .Y(new_n10874_1));
  nand_5 g08526(.A(new_n10874_1), .B(new_n2394), .Y(new_n10875));
  nand_5 g08527(.A(new_n10873), .B(n16722), .Y(new_n10876));
  nand_5 g08528(.A(new_n10876), .B(new_n10875), .Y(new_n10877));
  xor_4  g08529(.A(new_n10877), .B(new_n10870), .Y(new_n10878));
  not_8  g08530(.A(new_n10878), .Y(new_n10879));
  nand_5 g08531(.A(new_n10856), .B(new_n10852), .Y(new_n10880));
  nand_5 g08532(.A(new_n10880), .B(new_n10857), .Y(new_n10881));
  not_8  g08533(.A(new_n10881), .Y(new_n10882));
  not_8  g08534(.A(new_n10853), .Y(new_n10883));
  nand_5 g08535(.A(new_n10883), .B(new_n6820), .Y(new_n10884));
  nand_5 g08536(.A(new_n10853), .B(n26882), .Y(new_n10885));
  nand_5 g08537(.A(new_n10885), .B(new_n10884), .Y(new_n10886));
  nand_5 g08538(.A(new_n10886), .B(new_n5538), .Y(new_n10887));
  nor_5  g08539(.A(new_n10886), .B(new_n5538), .Y(new_n10888));
  not_8  g08540(.A(new_n10888), .Y(new_n10889));
  nand_5 g08541(.A(new_n10889), .B(new_n10887), .Y(new_n10890));
  xor_4  g08542(.A(new_n10890), .B(new_n10882), .Y(new_n10891));
  not_8  g08543(.A(new_n10891), .Y(new_n10892));
  nand_5 g08544(.A(new_n10892), .B(new_n10879), .Y(new_n10893));
  nand_5 g08545(.A(new_n10891), .B(new_n10878), .Y(new_n10894));
  nand_5 g08546(.A(new_n10894), .B(new_n10893), .Y(new_n10895));
  xor_4  g08547(.A(new_n10895), .B(new_n10867), .Y(new_n10896));
  nand_5 g08548(.A(n20235), .B(new_n3051), .Y(new_n10897));
  nand_5 g08549(.A(new_n9765), .B(n6502), .Y(new_n10898));
  nand_5 g08550(.A(n15780), .B(new_n5669), .Y(new_n10899));
  nand_5 g08551(.A(new_n10899), .B(new_n10898), .Y(new_n10900));
  nand_5 g08552(.A(new_n10900), .B(new_n10897), .Y(new_n10901));
  nand_5 g08553(.A(new_n3046), .B(n8381), .Y(new_n10902));
  nand_5 g08554(.A(n18295), .B(new_n5709), .Y(new_n10903));
  nand_5 g08555(.A(new_n10903), .B(new_n10902), .Y(new_n10904));
  xor_4  g08556(.A(new_n10904), .B(new_n10901), .Y(new_n10905));
  or_5   g08557(.A(new_n10905), .B(new_n10896), .Y(new_n10906));
  nand_5 g08558(.A(new_n10905), .B(new_n10896), .Y(new_n10907));
  not_8  g08559(.A(new_n10863), .Y(new_n10908));
  nand_5 g08560(.A(new_n10908), .B(new_n6553), .Y(new_n10909));
  and_5  g08561(.A(new_n10909), .B(new_n10864), .Y(new_n10910));
  not_8  g08562(.A(new_n10910), .Y(new_n10911));
  xor_4  g08563(.A(n15780), .B(new_n5669), .Y(new_n10912));
  nor_5  g08564(.A(new_n10912), .B(new_n10911), .Y(new_n10913));
  and_5  g08565(.A(new_n10898), .B(new_n10897), .Y(new_n10914));
  xor_4  g08566(.A(new_n10914), .B(new_n10899), .Y(new_n10915));
  nand_5 g08567(.A(new_n10915), .B(new_n10913), .Y(new_n10916));
  not_8  g08568(.A(new_n10859), .Y(new_n10917));
  nand_5 g08569(.A(new_n10917), .B(new_n6533), .Y(new_n10918));
  nand_5 g08570(.A(new_n10918), .B(new_n10860), .Y(new_n10919));
  xor_4  g08571(.A(new_n10919), .B(new_n10864), .Y(new_n10920));
  or_5   g08572(.A(new_n10915), .B(new_n10913), .Y(new_n10921));
  nand_5 g08573(.A(new_n10921), .B(new_n10920), .Y(new_n10922));
  nand_5 g08574(.A(new_n10922), .B(new_n10916), .Y(new_n10923));
  nand_5 g08575(.A(new_n10923), .B(new_n10907), .Y(new_n10924_1));
  nand_5 g08576(.A(new_n10924_1), .B(new_n10906), .Y(new_n10925));
  nand_5 g08577(.A(new_n10894), .B(new_n10867), .Y(new_n10926));
  nand_5 g08578(.A(new_n10926), .B(new_n10893), .Y(new_n10927));
  not_8  g08579(.A(new_n10927), .Y(new_n10928));
  nand_5 g08580(.A(new_n10889), .B(new_n10881), .Y(new_n10929));
  nand_5 g08581(.A(new_n10929), .B(new_n10887), .Y(new_n10930));
  not_8  g08582(.A(new_n10884), .Y(new_n10931));
  nand_5 g08583(.A(new_n10931), .B(new_n6817), .Y(new_n10932));
  nand_5 g08584(.A(new_n10884), .B(n20478), .Y(new_n10933));
  and_5  g08585(.A(new_n10933), .B(new_n10932), .Y(new_n10934));
  or_5   g08586(.A(new_n10934), .B(n7305), .Y(new_n10935));
  nand_5 g08587(.A(new_n10934), .B(n7305), .Y(new_n10936));
  nand_5 g08588(.A(new_n10936), .B(new_n10935), .Y(new_n10937));
  xor_4  g08589(.A(new_n10937), .B(new_n10930), .Y(new_n10938));
  not_8  g08590(.A(new_n10938), .Y(new_n10939));
  nand_5 g08591(.A(new_n10876), .B(new_n10869), .Y(new_n10940));
  nand_5 g08592(.A(new_n10940), .B(new_n10875), .Y(new_n10941));
  not_8  g08593(.A(new_n10941), .Y(new_n10942));
  nor_5  g08594(.A(new_n10871), .B(n25074), .Y(new_n10943_1));
  not_8  g08595(.A(new_n10943_1), .Y(new_n10944));
  nand_5 g08596(.A(new_n10871), .B(n25074), .Y(new_n10945));
  and_5  g08597(.A(new_n10945), .B(new_n10944), .Y(new_n10946));
  not_8  g08598(.A(new_n10946), .Y(new_n10947));
  nand_5 g08599(.A(new_n10947), .B(new_n2401), .Y(new_n10948));
  nand_5 g08600(.A(new_n10946), .B(n3480), .Y(new_n10949));
  nand_5 g08601(.A(new_n10949), .B(new_n10948), .Y(new_n10950));
  xor_4  g08602(.A(new_n10950), .B(new_n10942), .Y(new_n10951));
  nand_5 g08603(.A(new_n10951), .B(new_n10939), .Y(new_n10952));
  not_8  g08604(.A(new_n10951), .Y(new_n10953));
  nand_5 g08605(.A(new_n10953), .B(new_n10938), .Y(new_n10954));
  nand_5 g08606(.A(new_n10954), .B(new_n10952), .Y(new_n10955));
  xor_4  g08607(.A(new_n10955), .B(new_n10928), .Y(new_n10956));
  nand_5 g08608(.A(new_n10903), .B(new_n10901), .Y(new_n10957));
  nand_5 g08609(.A(new_n10957), .B(new_n10902), .Y(new_n10958));
  nand_5 g08610(.A(new_n3043), .B(n7057), .Y(new_n10959));
  nand_5 g08611(.A(n12956), .B(new_n9760), .Y(new_n10960));
  nand_5 g08612(.A(new_n10960), .B(new_n10959), .Y(new_n10961_1));
  xnor_4 g08613(.A(new_n10961_1), .B(new_n10958), .Y(new_n10962));
  nand_5 g08614(.A(new_n10962), .B(new_n10956), .Y(new_n10963));
  or_5   g08615(.A(new_n10962), .B(new_n10956), .Y(new_n10964));
  nand_5 g08616(.A(new_n10964), .B(new_n10963), .Y(new_n10965));
  xnor_4 g08617(.A(new_n10965), .B(new_n10925), .Y(n1060));
  nand_5 g08618(.A(new_n3624), .B(new_n3625), .Y(new_n10967));
  xnor_4 g08619(.A(new_n10967), .B(new_n3677), .Y(n1069));
  not_8  g08620(.A(n21749), .Y(new_n10969));
  not_8  g08621(.A(n26744), .Y(new_n10970));
  nand_5 g08622(.A(new_n10970), .B(new_n10969), .Y(new_n10971));
  nand_5 g08623(.A(n26744), .B(n21749), .Y(new_n10972));
  not_8  g08624(.A(n7769), .Y(new_n10973));
  not_8  g08625(.A(n26625), .Y(new_n10974));
  nand_5 g08626(.A(new_n10974), .B(new_n10973), .Y(new_n10975));
  nand_5 g08627(.A(n26625), .B(n7769), .Y(new_n10976));
  nand_5 g08628(.A(new_n10976), .B(new_n8275), .Y(new_n10977));
  nand_5 g08629(.A(new_n10977), .B(new_n10975), .Y(new_n10978));
  nand_5 g08630(.A(new_n10978), .B(new_n10972), .Y(new_n10979));
  nand_5 g08631(.A(new_n10979), .B(new_n10971), .Y(new_n10980));
  nand_5 g08632(.A(n11566), .B(n1558), .Y(new_n10981));
  not_8  g08633(.A(n1558), .Y(new_n10982));
  not_8  g08634(.A(n11566), .Y(new_n10983));
  nand_5 g08635(.A(new_n10983), .B(new_n10982), .Y(new_n10984));
  nand_5 g08636(.A(new_n10984), .B(new_n10981), .Y(new_n10985));
  xnor_4 g08637(.A(new_n10985), .B(new_n10980), .Y(new_n10986));
  not_8  g08638(.A(new_n10986), .Y(new_n10987));
  nand_5 g08639(.A(new_n7792), .B(new_n2673), .Y(new_n10988));
  nand_5 g08640(.A(new_n7791), .B(n1136), .Y(new_n10989));
  nand_5 g08641(.A(new_n10989), .B(new_n8280), .Y(new_n10990));
  nand_5 g08642(.A(new_n10990), .B(new_n10988), .Y(new_n10991));
  nand_5 g08643(.A(new_n7782), .B(new_n2669), .Y(new_n10992));
  nand_5 g08644(.A(new_n7780_1), .B(n23369), .Y(new_n10993));
  nand_5 g08645(.A(new_n10993), .B(new_n10992), .Y(new_n10994));
  xor_4  g08646(.A(new_n10994), .B(new_n10991), .Y(new_n10995));
  not_8  g08647(.A(new_n10995), .Y(new_n10996));
  not_8  g08648(.A(n17095), .Y(new_n10997));
  not_8  g08649(.A(n22591), .Y(new_n10998));
  nand_5 g08650(.A(new_n8284), .B(new_n10998), .Y(new_n10999));
  not_8  g08651(.A(new_n10999), .Y(new_n11000));
  nand_5 g08652(.A(new_n11000), .B(new_n10997), .Y(new_n11001));
  not_8  g08653(.A(new_n11001), .Y(new_n11002));
  nor_5  g08654(.A(new_n11000), .B(new_n10997), .Y(new_n11003));
  or_5   g08655(.A(new_n11003), .B(new_n11002), .Y(new_n11004));
  or_5   g08656(.A(new_n11004), .B(new_n10996), .Y(new_n11005_1));
  nand_5 g08657(.A(new_n11004), .B(new_n10996), .Y(new_n11006));
  not_8  g08658(.A(new_n8283), .Y(new_n11007));
  nand_5 g08659(.A(new_n11007), .B(new_n10998), .Y(new_n11008));
  not_8  g08660(.A(new_n11008), .Y(new_n11009));
  nand_5 g08661(.A(new_n10988), .B(new_n10989), .Y(new_n11010));
  xor_4  g08662(.A(new_n11010), .B(new_n8280), .Y(new_n11011_1));
  not_8  g08663(.A(new_n11011_1), .Y(new_n11012));
  nor_5  g08664(.A(new_n8284), .B(new_n10998), .Y(new_n11013));
  nor_5  g08665(.A(new_n11013), .B(new_n11000), .Y(new_n11014));
  nor_5  g08666(.A(new_n11014), .B(new_n11007), .Y(new_n11015));
  nor_5  g08667(.A(new_n11015), .B(new_n11012), .Y(new_n11016));
  nor_5  g08668(.A(new_n11016), .B(new_n11009), .Y(new_n11017));
  not_8  g08669(.A(new_n11017), .Y(new_n11018));
  nand_5 g08670(.A(new_n11018), .B(new_n11006), .Y(new_n11019));
  nand_5 g08671(.A(new_n11019), .B(new_n11005_1), .Y(new_n11020));
  nand_5 g08672(.A(new_n10993), .B(new_n10991), .Y(new_n11021));
  nand_5 g08673(.A(new_n11021), .B(new_n10992), .Y(new_n11022));
  nand_5 g08674(.A(new_n7777), .B(new_n10053_1), .Y(new_n11023_1));
  nand_5 g08675(.A(new_n7775), .B(n17664), .Y(new_n11024));
  nand_5 g08676(.A(new_n11024), .B(new_n11023_1), .Y(new_n11025_1));
  xor_4  g08677(.A(new_n11025_1), .B(new_n11022), .Y(new_n11026));
  not_8  g08678(.A(new_n11026), .Y(new_n11027));
  not_8  g08679(.A(n15378), .Y(new_n11028));
  nand_5 g08680(.A(new_n11002), .B(new_n11028), .Y(new_n11029));
  nand_5 g08681(.A(new_n11001), .B(n15378), .Y(new_n11030));
  nand_5 g08682(.A(new_n11030), .B(new_n11029), .Y(new_n11031));
  or_5   g08683(.A(new_n11031), .B(new_n11027), .Y(new_n11032));
  nand_5 g08684(.A(new_n11031), .B(new_n11027), .Y(new_n11033));
  nand_5 g08685(.A(new_n11033), .B(new_n11032), .Y(new_n11034));
  xor_4  g08686(.A(new_n11034), .B(new_n11020), .Y(new_n11035));
  nand_5 g08687(.A(new_n11035), .B(new_n10987), .Y(new_n11036));
  or_5   g08688(.A(new_n11035), .B(new_n10987), .Y(new_n11037));
  nand_5 g08689(.A(new_n10972), .B(new_n10971), .Y(new_n11038));
  xor_4  g08690(.A(new_n11038), .B(new_n10978), .Y(new_n11039));
  not_8  g08691(.A(new_n11039), .Y(new_n11040));
  nand_5 g08692(.A(new_n11006), .B(new_n11005_1), .Y(new_n11041));
  xor_4  g08693(.A(new_n11041), .B(new_n11017), .Y(new_n11042));
  or_5   g08694(.A(new_n11042), .B(new_n11040), .Y(new_n11043));
  nand_5 g08695(.A(new_n11042), .B(new_n11040), .Y(new_n11044_1));
  nor_5  g08696(.A(new_n11015), .B(new_n11009), .Y(new_n11045));
  xor_4  g08697(.A(new_n11045), .B(new_n11012), .Y(new_n11046));
  nand_5 g08698(.A(new_n10976), .B(new_n10975), .Y(new_n11047));
  xor_4  g08699(.A(new_n11047), .B(new_n8275), .Y(new_n11048));
  nand_5 g08700(.A(new_n11048), .B(new_n11046), .Y(new_n11049));
  not_8  g08701(.A(new_n11049), .Y(new_n11050));
  or_5   g08702(.A(new_n11048), .B(new_n11046), .Y(new_n11051));
  not_8  g08703(.A(new_n11051), .Y(new_n11052));
  nor_5  g08704(.A(new_n11052), .B(new_n8288_1), .Y(new_n11053));
  nor_5  g08705(.A(new_n11053), .B(new_n11050), .Y(new_n11054));
  not_8  g08706(.A(new_n11054), .Y(new_n11055));
  nand_5 g08707(.A(new_n11055), .B(new_n11044_1), .Y(new_n11056_1));
  nand_5 g08708(.A(new_n11056_1), .B(new_n11043), .Y(new_n11057));
  nand_5 g08709(.A(new_n11057), .B(new_n11037), .Y(new_n11058));
  nand_5 g08710(.A(new_n11058), .B(new_n11036), .Y(new_n11059));
  nand_5 g08711(.A(new_n10981), .B(new_n10980), .Y(new_n11060));
  nand_5 g08712(.A(new_n11060), .B(new_n10984), .Y(new_n11061));
  not_8  g08713(.A(n3959), .Y(new_n11062));
  not_8  g08714(.A(n9832), .Y(new_n11063_1));
  nand_5 g08715(.A(new_n11063_1), .B(new_n11062), .Y(new_n11064));
  nand_5 g08716(.A(n9832), .B(n3959), .Y(new_n11065));
  nand_5 g08717(.A(new_n11065), .B(new_n11064), .Y(new_n11066));
  xnor_4 g08718(.A(new_n11066), .B(new_n11061), .Y(new_n11067));
  not_8  g08719(.A(new_n11067), .Y(new_n11068));
  nand_5 g08720(.A(new_n11033), .B(new_n11020), .Y(new_n11069));
  nand_5 g08721(.A(new_n11069), .B(new_n11032), .Y(new_n11070));
  nand_5 g08722(.A(new_n11024), .B(new_n11022), .Y(new_n11071));
  nand_5 g08723(.A(new_n11071), .B(new_n11023_1), .Y(new_n11072));
  not_8  g08724(.A(new_n11072), .Y(new_n11073));
  nand_5 g08725(.A(new_n7772), .B(new_n2663), .Y(new_n11074));
  nand_5 g08726(.A(new_n7770), .B(n5226), .Y(new_n11075));
  nand_5 g08727(.A(new_n11075), .B(new_n11074), .Y(new_n11076));
  xor_4  g08728(.A(new_n11076), .B(new_n11073), .Y(new_n11077));
  not_8  g08729(.A(new_n11077), .Y(new_n11078_1));
  or_5   g08730(.A(new_n11029), .B(n19575), .Y(new_n11079));
  nand_5 g08731(.A(new_n11029), .B(n19575), .Y(new_n11080_1));
  and_5  g08732(.A(new_n11080_1), .B(new_n11079), .Y(new_n11081));
  nand_5 g08733(.A(new_n11081), .B(new_n11078_1), .Y(new_n11082));
  or_5   g08734(.A(new_n11081), .B(new_n11078_1), .Y(new_n11083));
  nand_5 g08735(.A(new_n11083), .B(new_n11082), .Y(new_n11084));
  xor_4  g08736(.A(new_n11084), .B(new_n11070), .Y(new_n11085));
  nand_5 g08737(.A(new_n11085), .B(new_n11068), .Y(new_n11086));
  or_5   g08738(.A(new_n11085), .B(new_n11068), .Y(new_n11087));
  nand_5 g08739(.A(new_n11087), .B(new_n11086), .Y(new_n11088));
  xor_4  g08740(.A(new_n11088), .B(new_n11059), .Y(n1111));
  nand_5 g08741(.A(new_n2716), .B(new_n4952_1), .Y(new_n11090));
  nand_5 g08742(.A(new_n2713), .B(n12446), .Y(new_n11091));
  or_5   g08743(.A(new_n2719), .B(n11011), .Y(new_n11092));
  nand_5 g08744(.A(new_n2719), .B(n11011), .Y(new_n11093));
  nand_5 g08745(.A(new_n2726), .B(new_n6249), .Y(new_n11094_1));
  nand_5 g08746(.A(new_n2723), .B(n16029), .Y(new_n11095));
  or_5   g08747(.A(new_n2729), .B(n16476), .Y(new_n11096));
  nand_5 g08748(.A(new_n2729), .B(n16476), .Y(new_n11097));
  nand_5 g08749(.A(new_n2736), .B(new_n6255), .Y(new_n11098));
  nand_5 g08750(.A(new_n2733), .B(n11615), .Y(new_n11099));
  nand_5 g08751(.A(new_n2742), .B(new_n6258), .Y(new_n11100));
  nand_5 g08752(.A(new_n2739), .B(n22433), .Y(new_n11101_1));
  nand_5 g08753(.A(new_n2746), .B(n14090), .Y(new_n11102));
  nand_5 g08754(.A(new_n11102), .B(new_n11101_1), .Y(new_n11103_1));
  nand_5 g08755(.A(new_n11103_1), .B(new_n11100), .Y(new_n11104));
  nand_5 g08756(.A(new_n11104), .B(new_n11099), .Y(new_n11105));
  nand_5 g08757(.A(new_n11105), .B(new_n11098), .Y(new_n11106));
  nand_5 g08758(.A(new_n11106), .B(new_n11097), .Y(new_n11107));
  nand_5 g08759(.A(new_n11107), .B(new_n11096), .Y(new_n11108));
  nand_5 g08760(.A(new_n11108), .B(new_n11095), .Y(new_n11109));
  nand_5 g08761(.A(new_n11109), .B(new_n11094_1), .Y(new_n11110));
  nand_5 g08762(.A(new_n11110), .B(new_n11093), .Y(new_n11111));
  nand_5 g08763(.A(new_n11111), .B(new_n11092), .Y(new_n11112));
  nand_5 g08764(.A(new_n11112), .B(new_n11091), .Y(new_n11113));
  nand_5 g08765(.A(new_n11113), .B(new_n11090), .Y(new_n11114));
  nand_5 g08766(.A(new_n2710), .B(new_n6240), .Y(new_n11115));
  nand_5 g08767(.A(new_n2707), .B(n23849), .Y(new_n11116));
  nand_5 g08768(.A(new_n11116), .B(new_n11115), .Y(new_n11117));
  xor_4  g08769(.A(new_n11117), .B(new_n11114), .Y(new_n11118));
  not_8  g08770(.A(new_n2858_1), .Y(new_n11119));
  nand_5 g08771(.A(new_n10943_1), .B(new_n3078), .Y(new_n11120_1));
  nor_5  g08772(.A(new_n11120_1), .B(n20929), .Y(new_n11121_1));
  nand_5 g08773(.A(new_n11121_1), .B(new_n3108), .Y(new_n11122));
  not_8  g08774(.A(new_n11122), .Y(new_n11123));
  nor_5  g08775(.A(new_n11121_1), .B(new_n3108), .Y(new_n11124));
  nor_5  g08776(.A(new_n11124), .B(new_n11123), .Y(new_n11125));
  not_8  g08777(.A(new_n11125), .Y(new_n11126));
  nand_5 g08778(.A(new_n11126), .B(new_n11119), .Y(new_n11127_1));
  nand_5 g08779(.A(new_n11125), .B(new_n2858_1), .Y(new_n11128));
  not_8  g08780(.A(new_n2864), .Y(new_n11129));
  xor_4  g08781(.A(new_n11120_1), .B(n20929), .Y(new_n11130));
  not_8  g08782(.A(new_n11130), .Y(new_n11131));
  nand_5 g08783(.A(new_n11131), .B(new_n11129), .Y(new_n11132_1));
  nand_5 g08784(.A(new_n11130), .B(new_n2864), .Y(new_n11133));
  not_8  g08785(.A(new_n2869), .Y(new_n11134_1));
  nand_5 g08786(.A(new_n10944), .B(n8006), .Y(new_n11135));
  and_5  g08787(.A(new_n11135), .B(new_n11120_1), .Y(new_n11136));
  not_8  g08788(.A(new_n11136), .Y(new_n11137));
  nand_5 g08789(.A(new_n11137), .B(new_n11134_1), .Y(new_n11138_1));
  nand_5 g08790(.A(new_n11136), .B(new_n2869), .Y(new_n11139));
  nand_5 g08791(.A(new_n10947), .B(new_n2875), .Y(new_n11140));
  nand_5 g08792(.A(new_n10946), .B(new_n2874), .Y(new_n11141));
  nand_5 g08793(.A(new_n10874_1), .B(new_n2883), .Y(new_n11142));
  nand_5 g08794(.A(new_n10873), .B(new_n2884), .Y(new_n11143));
  nand_5 g08795(.A(new_n6529), .B(new_n2889), .Y(new_n11144));
  nand_5 g08796(.A(new_n6528), .B(new_n2890), .Y(new_n11145));
  nand_5 g08797(.A(new_n2893), .B(new_n3163), .Y(new_n11146));
  not_8  g08798(.A(new_n11146), .Y(new_n11147));
  nand_5 g08799(.A(new_n11147), .B(new_n11145), .Y(new_n11148));
  nand_5 g08800(.A(new_n11148), .B(new_n11144), .Y(new_n11149));
  nand_5 g08801(.A(new_n11149), .B(new_n11143), .Y(new_n11150));
  nand_5 g08802(.A(new_n11150), .B(new_n11142), .Y(new_n11151));
  nand_5 g08803(.A(new_n11151), .B(new_n11141), .Y(new_n11152));
  nand_5 g08804(.A(new_n11152), .B(new_n11140), .Y(new_n11153));
  nand_5 g08805(.A(new_n11153), .B(new_n11139), .Y(new_n11154));
  nand_5 g08806(.A(new_n11154), .B(new_n11138_1), .Y(new_n11155));
  nand_5 g08807(.A(new_n11155), .B(new_n11133), .Y(new_n11156));
  nand_5 g08808(.A(new_n11156), .B(new_n11132_1), .Y(new_n11157));
  nand_5 g08809(.A(new_n11157), .B(new_n11128), .Y(new_n11158));
  nand_5 g08810(.A(new_n11158), .B(new_n11127_1), .Y(new_n11159));
  not_8  g08811(.A(new_n2853_1), .Y(new_n11160));
  nand_5 g08812(.A(new_n11123), .B(new_n3194), .Y(new_n11161));
  nand_5 g08813(.A(new_n11122), .B(n11841), .Y(new_n11162));
  and_5  g08814(.A(new_n11162), .B(new_n11161), .Y(new_n11163));
  not_8  g08815(.A(new_n11163), .Y(new_n11164));
  nand_5 g08816(.A(new_n11164), .B(new_n11160), .Y(new_n11165));
  nand_5 g08817(.A(new_n11163), .B(new_n2853_1), .Y(new_n11166));
  nand_5 g08818(.A(new_n11166), .B(new_n11165), .Y(new_n11167));
  xor_4  g08819(.A(new_n11167), .B(new_n11159), .Y(new_n11168));
  or_5   g08820(.A(new_n11168), .B(new_n11118), .Y(new_n11169));
  nand_5 g08821(.A(new_n11168), .B(new_n11118), .Y(new_n11170));
  nand_5 g08822(.A(new_n11090), .B(new_n11091), .Y(new_n11171));
  xor_4  g08823(.A(new_n11171), .B(new_n11112), .Y(new_n11172));
  nand_5 g08824(.A(new_n11127_1), .B(new_n11128), .Y(new_n11173));
  xor_4  g08825(.A(new_n11173), .B(new_n11157), .Y(new_n11174));
  or_5   g08826(.A(new_n11174), .B(new_n11172), .Y(new_n11175));
  nand_5 g08827(.A(new_n11174), .B(new_n11172), .Y(new_n11176));
  nand_5 g08828(.A(new_n11092), .B(new_n11093), .Y(new_n11177));
  xor_4  g08829(.A(new_n11177), .B(new_n11110), .Y(new_n11178));
  nand_5 g08830(.A(new_n11132_1), .B(new_n11133), .Y(new_n11179));
  xor_4  g08831(.A(new_n11179), .B(new_n11155), .Y(new_n11180));
  or_5   g08832(.A(new_n11180), .B(new_n11178), .Y(new_n11181));
  nand_5 g08833(.A(new_n11180), .B(new_n11178), .Y(new_n11182_1));
  nand_5 g08834(.A(new_n11094_1), .B(new_n11095), .Y(new_n11183));
  xor_4  g08835(.A(new_n11183), .B(new_n11108), .Y(new_n11184_1));
  nand_5 g08836(.A(new_n11138_1), .B(new_n11139), .Y(new_n11185));
  xor_4  g08837(.A(new_n11185), .B(new_n11153), .Y(new_n11186));
  or_5   g08838(.A(new_n11186), .B(new_n11184_1), .Y(new_n11187));
  nand_5 g08839(.A(new_n11186), .B(new_n11184_1), .Y(new_n11188));
  nand_5 g08840(.A(new_n11140), .B(new_n11141), .Y(new_n11189));
  xor_4  g08841(.A(new_n11189), .B(new_n11151), .Y(new_n11190));
  nand_5 g08842(.A(new_n11096), .B(new_n11097), .Y(new_n11191));
  xor_4  g08843(.A(new_n11191), .B(new_n11106), .Y(new_n11192_1));
  or_5   g08844(.A(new_n11192_1), .B(new_n11190), .Y(new_n11193));
  nand_5 g08845(.A(new_n11192_1), .B(new_n11190), .Y(new_n11194));
  nand_5 g08846(.A(new_n11098), .B(new_n11099), .Y(new_n11195));
  xor_4  g08847(.A(new_n11195), .B(new_n11104), .Y(new_n11196));
  nand_5 g08848(.A(new_n11142), .B(new_n11143), .Y(new_n11197));
  xor_4  g08849(.A(new_n11197), .B(new_n11149), .Y(new_n11198));
  or_5   g08850(.A(new_n11198), .B(new_n11196), .Y(new_n11199));
  nand_5 g08851(.A(new_n11198), .B(new_n11196), .Y(new_n11200));
  nand_5 g08852(.A(new_n11144), .B(new_n11145), .Y(new_n11201_1));
  xor_4  g08853(.A(new_n11201_1), .B(new_n11147), .Y(new_n11202));
  nand_5 g08854(.A(new_n11100), .B(new_n11101_1), .Y(new_n11203));
  xor_4  g08855(.A(new_n11203), .B(new_n11102), .Y(new_n11204));
  or_5   g08856(.A(new_n11204), .B(new_n11202), .Y(new_n11205));
  nand_5 g08857(.A(new_n11204), .B(new_n11202), .Y(new_n11206));
  nand_5 g08858(.A(new_n2974), .B(new_n2631), .Y(new_n11207));
  and_5  g08859(.A(new_n11207), .B(new_n11102), .Y(new_n11208));
  xor_4  g08860(.A(new_n2893), .B(n2088), .Y(new_n11209));
  nand_5 g08861(.A(new_n11209), .B(new_n11208), .Y(new_n11210));
  nand_5 g08862(.A(new_n11210), .B(new_n11206), .Y(new_n11211));
  nand_5 g08863(.A(new_n11211), .B(new_n11205), .Y(new_n11212));
  nand_5 g08864(.A(new_n11212), .B(new_n11200), .Y(new_n11213));
  nand_5 g08865(.A(new_n11213), .B(new_n11199), .Y(new_n11214));
  nand_5 g08866(.A(new_n11214), .B(new_n11194), .Y(new_n11215));
  nand_5 g08867(.A(new_n11215), .B(new_n11193), .Y(new_n11216));
  nand_5 g08868(.A(new_n11216), .B(new_n11188), .Y(new_n11217));
  nand_5 g08869(.A(new_n11217), .B(new_n11187), .Y(new_n11218));
  nand_5 g08870(.A(new_n11218), .B(new_n11182_1), .Y(new_n11219));
  nand_5 g08871(.A(new_n11219), .B(new_n11181), .Y(new_n11220_1));
  nand_5 g08872(.A(new_n11220_1), .B(new_n11176), .Y(new_n11221));
  nand_5 g08873(.A(new_n11221), .B(new_n11175), .Y(new_n11222));
  nand_5 g08874(.A(new_n11222), .B(new_n11170), .Y(new_n11223_1));
  nand_5 g08875(.A(new_n11223_1), .B(new_n11169), .Y(new_n11224));
  nand_5 g08876(.A(new_n11116), .B(new_n11114), .Y(new_n11225));
  nand_5 g08877(.A(new_n11225), .B(new_n11115), .Y(new_n11226));
  nand_5 g08878(.A(new_n2704), .B(new_n4942), .Y(new_n11227));
  nand_5 g08879(.A(new_n2701), .B(n25475), .Y(new_n11228));
  nand_5 g08880(.A(new_n11228), .B(new_n11227), .Y(new_n11229));
  xor_4  g08881(.A(new_n11229), .B(new_n11226), .Y(new_n11230));
  nand_5 g08882(.A(new_n11166), .B(new_n11159), .Y(new_n11231));
  nand_5 g08883(.A(new_n11231), .B(new_n11165), .Y(new_n11232));
  not_8  g08884(.A(new_n11232), .Y(new_n11233));
  not_8  g08885(.A(new_n2848), .Y(new_n11234_1));
  or_5   g08886(.A(new_n11161), .B(n27089), .Y(new_n11235));
  nand_5 g08887(.A(new_n11161), .B(n27089), .Y(new_n11236));
  and_5  g08888(.A(new_n11236), .B(new_n11235), .Y(new_n11237));
  not_8  g08889(.A(new_n11237), .Y(new_n11238));
  nand_5 g08890(.A(new_n11238), .B(new_n11234_1), .Y(new_n11239));
  nand_5 g08891(.A(new_n11237), .B(new_n2848), .Y(new_n11240));
  nand_5 g08892(.A(new_n11240), .B(new_n11239), .Y(new_n11241));
  xor_4  g08893(.A(new_n11241), .B(new_n11233), .Y(new_n11242));
  not_8  g08894(.A(new_n11242), .Y(new_n11243));
  nand_5 g08895(.A(new_n11243), .B(new_n11230), .Y(new_n11244));
  not_8  g08896(.A(new_n11230), .Y(new_n11245_1));
  nand_5 g08897(.A(new_n11242), .B(new_n11245_1), .Y(new_n11246));
  nand_5 g08898(.A(new_n11246), .B(new_n11244), .Y(new_n11247));
  xor_4  g08899(.A(new_n11247), .B(new_n11224), .Y(n1119));
  nand_5 g08900(.A(new_n9065), .B(new_n9064), .Y(new_n11249));
  xor_4  g08901(.A(new_n11249), .B(new_n9088), .Y(n1120));
  not_8  g08902(.A(new_n8919), .Y(new_n11251));
  nand_5 g08903(.A(n9246), .B(n3925), .Y(new_n11252));
  nand_5 g08904(.A(new_n3827), .B(new_n5549), .Y(new_n11253));
  nand_5 g08905(.A(new_n11253), .B(new_n11252), .Y(new_n11254));
  xor_4  g08906(.A(new_n11254), .B(new_n11251), .Y(new_n11255));
  not_8  g08907(.A(n7428), .Y(new_n11256));
  nand_5 g08908(.A(n12495), .B(new_n11256), .Y(new_n11257));
  nand_5 g08909(.A(new_n5669), .B(n7428), .Y(new_n11258));
  nand_5 g08910(.A(new_n11258), .B(new_n11257), .Y(new_n11259));
  nand_5 g08911(.A(new_n11259), .B(new_n11255), .Y(new_n11260));
  not_8  g08912(.A(new_n11260), .Y(new_n11261_1));
  nor_5  g08913(.A(new_n11259), .B(new_n11255), .Y(new_n11262));
  nor_5  g08914(.A(new_n11262), .B(new_n11261_1), .Y(n1196));
  nand_5 g08915(.A(n6794), .B(new_n2506), .Y(new_n11264));
  nand_5 g08916(.A(new_n2442), .B(n2387), .Y(new_n11265));
  nand_5 g08917(.A(new_n11265), .B(new_n11264), .Y(new_n11266_1));
  nand_5 g08918(.A(new_n11266_1), .B(new_n9068), .Y(new_n11267));
  not_8  g08919(.A(new_n11264), .Y(new_n11268));
  nand_5 g08920(.A(new_n2358), .B(n19494), .Y(new_n11269));
  nand_5 g08921(.A(n20077), .B(new_n2504), .Y(new_n11270));
  and_5  g08922(.A(new_n11270), .B(new_n11269), .Y(new_n11271));
  xor_4  g08923(.A(new_n11271), .B(new_n11268), .Y(new_n11272));
  or_5   g08924(.A(new_n11272), .B(new_n11267), .Y(new_n11273_1));
  nand_5 g08925(.A(new_n11272), .B(new_n11267), .Y(new_n11274));
  nand_5 g08926(.A(new_n11274), .B(new_n9079), .Y(new_n11275_1));
  nand_5 g08927(.A(new_n11275_1), .B(new_n11273_1), .Y(new_n11276));
  nand_5 g08928(.A(new_n11270), .B(new_n11264), .Y(new_n11277));
  nand_5 g08929(.A(new_n11277), .B(new_n11269), .Y(new_n11278));
  nand_5 g08930(.A(n16223), .B(new_n2353), .Y(new_n11279));
  nand_5 g08931(.A(new_n2500), .B(n15636), .Y(new_n11280));
  nand_5 g08932(.A(new_n11280), .B(new_n11279), .Y(new_n11281));
  xnor_4 g08933(.A(new_n11281), .B(new_n11278), .Y(new_n11282));
  nand_5 g08934(.A(new_n11282), .B(new_n9067), .Y(new_n11283));
  not_8  g08935(.A(new_n11283), .Y(new_n11284));
  nor_5  g08936(.A(new_n11282), .B(new_n9067), .Y(new_n11285));
  nor_5  g08937(.A(new_n11285), .B(new_n11284), .Y(new_n11286));
  xor_4  g08938(.A(new_n11286), .B(new_n11276), .Y(n1237));
  not_8  g08939(.A(new_n6516), .Y(new_n11288));
  nand_5 g08940(.A(new_n11288), .B(new_n6433), .Y(new_n11289));
  xnor_4 g08941(.A(new_n11289), .B(new_n6514_1), .Y(n1239));
  nand_5 g08942(.A(new_n9151), .B(new_n9275), .Y(new_n11291));
  nand_5 g08943(.A(n22764), .B(n1536), .Y(new_n11292));
  nand_5 g08944(.A(new_n11292), .B(new_n11291), .Y(new_n11293));
  nand_5 g08945(.A(new_n9157), .B(new_n9281), .Y(new_n11294));
  not_8  g08946(.A(new_n11294), .Y(new_n11295));
  nand_5 g08947(.A(n26264), .B(n19454), .Y(new_n11296));
  not_8  g08948(.A(new_n11296), .Y(new_n11297));
  nand_5 g08949(.A(new_n9287_1), .B(new_n9163), .Y(new_n11298));
  not_8  g08950(.A(new_n11298), .Y(new_n11299));
  nand_5 g08951(.A(n9445), .B(n7841), .Y(new_n11300));
  not_8  g08952(.A(new_n11300), .Y(new_n11301));
  nand_5 g08953(.A(new_n9169), .B(new_n9293), .Y(new_n11302_1));
  not_8  g08954(.A(new_n11302_1), .Y(new_n11303));
  nand_5 g08955(.A(n16812), .B(n1279), .Y(new_n11304));
  not_8  g08956(.A(new_n11304), .Y(new_n11305));
  nand_5 g08957(.A(new_n9317), .B(new_n9193), .Y(new_n11306));
  nand_5 g08958(.A(n24485), .B(n16743), .Y(new_n11307));
  nand_5 g08959(.A(new_n9981), .B(new_n9323_1), .Y(new_n11308));
  nand_5 g08960(.A(n15258), .B(n2420), .Y(new_n11309));
  nand_5 g08961(.A(n22201), .B(n4588), .Y(new_n11310));
  nand_5 g08962(.A(new_n11310), .B(new_n11309), .Y(new_n11311));
  nand_5 g08963(.A(new_n11311), .B(new_n11308), .Y(new_n11312));
  nand_5 g08964(.A(new_n11312), .B(new_n11307), .Y(new_n11313_1));
  nand_5 g08965(.A(new_n11313_1), .B(new_n11306), .Y(new_n11314));
  nand_5 g08966(.A(new_n11314), .B(new_n9311), .Y(new_n11315));
  not_8  g08967(.A(new_n11315), .Y(new_n11316));
  nor_5  g08968(.A(new_n11314), .B(new_n9311), .Y(new_n11317));
  nor_5  g08969(.A(new_n11317), .B(n22631), .Y(new_n11318));
  nor_5  g08970(.A(new_n11318), .B(new_n11316), .Y(new_n11319));
  or_5   g08971(.A(new_n11319), .B(n2331), .Y(new_n11320));
  nand_5 g08972(.A(new_n11319), .B(n2331), .Y(new_n11321));
  nand_5 g08973(.A(new_n11321), .B(new_n9305), .Y(new_n11322));
  nand_5 g08974(.A(new_n11322), .B(new_n11320), .Y(new_n11323));
  nand_5 g08975(.A(new_n11323), .B(new_n9299), .Y(new_n11324));
  not_8  g08976(.A(new_n11324), .Y(new_n11325_1));
  nor_5  g08977(.A(new_n11323), .B(new_n9299), .Y(new_n11326_1));
  nor_5  g08978(.A(new_n11326_1), .B(n25068), .Y(new_n11327));
  nor_5  g08979(.A(new_n11327), .B(new_n11325_1), .Y(new_n11328));
  nor_5  g08980(.A(new_n11328), .B(new_n11305), .Y(new_n11329));
  nor_5  g08981(.A(new_n11329), .B(new_n11303), .Y(new_n11330_1));
  nor_5  g08982(.A(new_n11330_1), .B(new_n11301), .Y(new_n11331));
  nor_5  g08983(.A(new_n11331), .B(new_n11299), .Y(new_n11332));
  nor_5  g08984(.A(new_n11332), .B(new_n11297), .Y(new_n11333));
  nor_5  g08985(.A(new_n11333), .B(new_n11295), .Y(new_n11334));
  not_8  g08986(.A(new_n11334), .Y(new_n11335));
  xor_4  g08987(.A(new_n11335), .B(new_n11293), .Y(new_n11336));
  nand_5 g08988(.A(new_n11336), .B(n2416), .Y(new_n11337));
  not_8  g08989(.A(new_n11337), .Y(new_n11338));
  nor_5  g08990(.A(new_n11336), .B(n2416), .Y(new_n11339));
  not_8  g08991(.A(n21905), .Y(new_n11340));
  nand_5 g08992(.A(new_n11296), .B(new_n11294), .Y(new_n11341));
  xor_4  g08993(.A(new_n11341), .B(new_n11332), .Y(new_n11342));
  or_5   g08994(.A(new_n11342), .B(new_n11340), .Y(new_n11343));
  nand_5 g08995(.A(new_n11342), .B(new_n11340), .Y(new_n11344));
  not_8  g08996(.A(n22918), .Y(new_n11345));
  nand_5 g08997(.A(new_n11300), .B(new_n11298), .Y(new_n11346));
  xor_4  g08998(.A(new_n11346), .B(new_n11330_1), .Y(new_n11347_1));
  or_5   g08999(.A(new_n11347_1), .B(new_n11345), .Y(new_n11348_1));
  nand_5 g09000(.A(new_n11347_1), .B(new_n11345), .Y(new_n11349));
  not_8  g09001(.A(n25923), .Y(new_n11350));
  nand_5 g09002(.A(new_n11304), .B(new_n11302_1), .Y(new_n11351));
  xor_4  g09003(.A(new_n11351), .B(new_n11328), .Y(new_n11352_1));
  or_5   g09004(.A(new_n11352_1), .B(new_n11350), .Y(new_n11353));
  nand_5 g09005(.A(new_n11352_1), .B(new_n11350), .Y(new_n11354));
  not_8  g09006(.A(n6790), .Y(new_n11355));
  nor_5  g09007(.A(new_n11326_1), .B(new_n11325_1), .Y(new_n11356_1));
  xor_4  g09008(.A(new_n11356_1), .B(new_n9175), .Y(new_n11357));
  or_5   g09009(.A(new_n11357), .B(new_n11355), .Y(new_n11358));
  nand_5 g09010(.A(new_n11357), .B(new_n11355), .Y(new_n11359));
  not_8  g09011(.A(n22879), .Y(new_n11360));
  and_5  g09012(.A(new_n11321), .B(new_n11320), .Y(new_n11361));
  xor_4  g09013(.A(new_n11361), .B(new_n9305), .Y(new_n11362));
  or_5   g09014(.A(new_n11362), .B(new_n11360), .Y(new_n11363));
  nand_5 g09015(.A(new_n11362), .B(new_n11360), .Y(new_n11364));
  not_8  g09016(.A(n2117), .Y(new_n11365));
  nor_5  g09017(.A(new_n11317), .B(new_n11316), .Y(new_n11366));
  xor_4  g09018(.A(new_n11366), .B(new_n9187), .Y(new_n11367));
  or_5   g09019(.A(new_n11367), .B(new_n11365), .Y(new_n11368));
  nand_5 g09020(.A(new_n11367), .B(new_n11365), .Y(new_n11369));
  nand_5 g09021(.A(new_n11307), .B(new_n11306), .Y(new_n11370));
  xor_4  g09022(.A(new_n11370), .B(new_n11312), .Y(new_n11371));
  nand_5 g09023(.A(new_n11371), .B(n5882), .Y(new_n11372));
  or_5   g09024(.A(new_n11371), .B(n5882), .Y(new_n11373));
  nand_5 g09025(.A(new_n11309), .B(new_n11308), .Y(new_n11374));
  xor_4  g09026(.A(new_n11374), .B(new_n11310), .Y(new_n11375_1));
  nand_5 g09027(.A(new_n11375_1), .B(n11775), .Y(new_n11376));
  or_5   g09028(.A(new_n11375_1), .B(n11775), .Y(new_n11377));
  not_8  g09029(.A(n27134), .Y(new_n11378));
  nand_5 g09030(.A(new_n2619_1), .B(new_n2611), .Y(new_n11379_1));
  nand_5 g09031(.A(new_n11379_1), .B(new_n11310), .Y(new_n11380));
  nor_5  g09032(.A(new_n11380), .B(new_n11378), .Y(new_n11381));
  nand_5 g09033(.A(new_n11381), .B(new_n11377), .Y(new_n11382));
  nand_5 g09034(.A(new_n11382), .B(new_n11376), .Y(new_n11383));
  nand_5 g09035(.A(new_n11383), .B(new_n11373), .Y(new_n11384));
  nand_5 g09036(.A(new_n11384), .B(new_n11372), .Y(new_n11385));
  nand_5 g09037(.A(new_n11385), .B(new_n11369), .Y(new_n11386_1));
  nand_5 g09038(.A(new_n11386_1), .B(new_n11368), .Y(new_n11387));
  nand_5 g09039(.A(new_n11387), .B(new_n11364), .Y(new_n11388));
  nand_5 g09040(.A(new_n11388), .B(new_n11363), .Y(new_n11389));
  nand_5 g09041(.A(new_n11389), .B(new_n11359), .Y(new_n11390));
  nand_5 g09042(.A(new_n11390), .B(new_n11358), .Y(new_n11391_1));
  nand_5 g09043(.A(new_n11391_1), .B(new_n11354), .Y(new_n11392));
  nand_5 g09044(.A(new_n11392), .B(new_n11353), .Y(new_n11393));
  nand_5 g09045(.A(new_n11393), .B(new_n11349), .Y(new_n11394));
  nand_5 g09046(.A(new_n11394), .B(new_n11348_1), .Y(new_n11395));
  nand_5 g09047(.A(new_n11395), .B(new_n11344), .Y(new_n11396));
  nand_5 g09048(.A(new_n11396), .B(new_n11343), .Y(new_n11397));
  not_8  g09049(.A(new_n11397), .Y(new_n11398_1));
  nor_5  g09050(.A(new_n11398_1), .B(new_n11339), .Y(new_n11399));
  nor_5  g09051(.A(new_n11399), .B(new_n11338), .Y(new_n11400));
  nand_5 g09052(.A(new_n11335), .B(new_n11292), .Y(new_n11401));
  nand_5 g09053(.A(new_n11401), .B(new_n11291), .Y(new_n11402));
  or_5   g09054(.A(new_n11402), .B(new_n11400), .Y(new_n11403_1));
  not_8  g09055(.A(n13549), .Y(new_n11404));
  nand_5 g09056(.A(new_n9104_1), .B(new_n11404), .Y(new_n11405));
  nand_5 g09057(.A(n14826), .B(n13549), .Y(new_n11406));
  nand_5 g09058(.A(new_n11406), .B(new_n11405), .Y(new_n11407));
  not_8  g09059(.A(new_n11407), .Y(new_n11408));
  not_8  g09060(.A(n5532), .Y(new_n11409));
  nand_5 g09061(.A(new_n9113), .B(new_n11409), .Y(new_n11410));
  nand_5 g09062(.A(n15146), .B(n5532), .Y(new_n11411));
  not_8  g09063(.A(n3962), .Y(new_n11412));
  nand_5 g09064(.A(new_n9116), .B(new_n11412), .Y(new_n11413));
  nand_5 g09065(.A(n11579), .B(n3962), .Y(new_n11414));
  not_8  g09066(.A(n23513), .Y(new_n11415));
  nand_5 g09067(.A(new_n11415), .B(new_n9120), .Y(new_n11416));
  nand_5 g09068(.A(n23513), .B(n21), .Y(new_n11417));
  not_8  g09069(.A(n6427), .Y(new_n11418));
  nand_5 g09070(.A(new_n11418), .B(new_n9122), .Y(new_n11419_1));
  nand_5 g09071(.A(n6427), .B(n1682), .Y(new_n11420));
  not_8  g09072(.A(n6590), .Y(new_n11421));
  nand_5 g09073(.A(new_n9123), .B(new_n11421), .Y(new_n11422));
  nand_5 g09074(.A(n7963), .B(n6590), .Y(new_n11423));
  not_8  g09075(.A(n20349), .Y(new_n11424_1));
  nand_5 g09076(.A(new_n11424_1), .B(new_n9126), .Y(new_n11425));
  nand_5 g09077(.A(n20349), .B(n10017), .Y(new_n11426));
  nand_5 g09078(.A(n15936), .B(n3618), .Y(new_n11427));
  nand_5 g09079(.A(new_n11427), .B(new_n11426), .Y(new_n11428));
  nand_5 g09080(.A(new_n11428), .B(new_n11425), .Y(new_n11429));
  nand_5 g09081(.A(new_n11429), .B(new_n11423), .Y(new_n11430));
  nand_5 g09082(.A(new_n11430), .B(new_n11422), .Y(new_n11431));
  nand_5 g09083(.A(new_n11431), .B(new_n11420), .Y(new_n11432));
  nand_5 g09084(.A(new_n11432), .B(new_n11419_1), .Y(new_n11433));
  nand_5 g09085(.A(new_n11433), .B(new_n11417), .Y(new_n11434));
  nand_5 g09086(.A(new_n11434), .B(new_n11416), .Y(new_n11435));
  nand_5 g09087(.A(new_n11435), .B(new_n11414), .Y(new_n11436));
  nand_5 g09088(.A(new_n11436), .B(new_n11413), .Y(new_n11437));
  nand_5 g09089(.A(new_n11437), .B(new_n11411), .Y(new_n11438));
  nand_5 g09090(.A(new_n11438), .B(new_n11410), .Y(new_n11439_1));
  nand_5 g09091(.A(n22359), .B(n10275), .Y(new_n11440));
  nand_5 g09092(.A(new_n11440), .B(new_n11439_1), .Y(new_n11441));
  not_8  g09093(.A(n22359), .Y(new_n11442));
  nand_5 g09094(.A(new_n11442), .B(new_n9110), .Y(new_n11443));
  nand_5 g09095(.A(new_n11443), .B(new_n11441), .Y(new_n11444));
  nand_5 g09096(.A(n23493), .B(n8405), .Y(new_n11445));
  nand_5 g09097(.A(new_n11445), .B(new_n11444), .Y(new_n11446));
  not_8  g09098(.A(n8405), .Y(new_n11447));
  nand_5 g09099(.A(new_n9107), .B(new_n11447), .Y(new_n11448));
  nand_5 g09100(.A(new_n11448), .B(new_n11446), .Y(new_n11449));
  xor_4  g09101(.A(new_n11449), .B(new_n11408), .Y(new_n11450));
  or_5   g09102(.A(new_n11450), .B(new_n9229), .Y(new_n11451));
  nand_5 g09103(.A(new_n11450), .B(new_n9229), .Y(new_n11452));
  nand_5 g09104(.A(n23493), .B(new_n11447), .Y(new_n11453));
  nand_5 g09105(.A(new_n9107), .B(n8405), .Y(new_n11454));
  nand_5 g09106(.A(new_n11454), .B(new_n11453), .Y(new_n11455_1));
  xor_4  g09107(.A(new_n11455_1), .B(new_n11444), .Y(new_n11456));
  or_5   g09108(.A(new_n11456), .B(new_n4928), .Y(new_n11457));
  nand_5 g09109(.A(new_n11456), .B(new_n4928), .Y(new_n11458));
  nand_5 g09110(.A(new_n11442), .B(n10275), .Y(new_n11459));
  nand_5 g09111(.A(n22359), .B(new_n9110), .Y(new_n11460));
  nand_5 g09112(.A(new_n11460), .B(new_n11459), .Y(new_n11461));
  xor_4  g09113(.A(new_n11461), .B(new_n11439_1), .Y(new_n11462_1));
  or_5   g09114(.A(new_n11462_1), .B(new_n9233), .Y(new_n11463));
  nand_5 g09115(.A(new_n11462_1), .B(new_n9233), .Y(new_n11464));
  nand_5 g09116(.A(new_n11411), .B(new_n11410), .Y(new_n11465));
  not_8  g09117(.A(new_n11465), .Y(new_n11466));
  xor_4  g09118(.A(new_n11466), .B(new_n11437), .Y(new_n11467));
  or_5   g09119(.A(new_n11467), .B(new_n4929), .Y(new_n11468));
  nand_5 g09120(.A(new_n11467), .B(new_n4929), .Y(new_n11469));
  nand_5 g09121(.A(new_n11414), .B(new_n11413), .Y(new_n11470_1));
  not_8  g09122(.A(new_n11470_1), .Y(new_n11471));
  xor_4  g09123(.A(new_n11471), .B(new_n11435), .Y(new_n11472_1));
  or_5   g09124(.A(new_n11472_1), .B(new_n9239), .Y(new_n11473_1));
  nand_5 g09125(.A(new_n11472_1), .B(new_n9239), .Y(new_n11474));
  nand_5 g09126(.A(new_n11417), .B(new_n11416), .Y(new_n11475));
  not_8  g09127(.A(new_n11475), .Y(new_n11476));
  xor_4  g09128(.A(new_n11476), .B(new_n11433), .Y(new_n11477));
  or_5   g09129(.A(new_n11477), .B(new_n4930), .Y(new_n11478));
  nand_5 g09130(.A(new_n11477), .B(new_n4930), .Y(new_n11479_1));
  nand_5 g09131(.A(new_n11420), .B(new_n11419_1), .Y(new_n11480));
  not_8  g09132(.A(new_n11480), .Y(new_n11481_1));
  xor_4  g09133(.A(new_n11481_1), .B(new_n11431), .Y(new_n11482));
  or_5   g09134(.A(new_n11482), .B(new_n9245), .Y(new_n11483));
  nand_5 g09135(.A(new_n11482), .B(new_n9245), .Y(new_n11484));
  nand_5 g09136(.A(new_n11423), .B(new_n11422), .Y(new_n11485));
  not_8  g09137(.A(new_n11485), .Y(new_n11486_1));
  xor_4  g09138(.A(new_n11486_1), .B(new_n11429), .Y(new_n11487));
  or_5   g09139(.A(new_n11487), .B(new_n9249), .Y(new_n11488));
  nand_5 g09140(.A(new_n11487), .B(new_n9249), .Y(new_n11489));
  nand_5 g09141(.A(new_n11426), .B(new_n11425), .Y(new_n11490));
  xor_4  g09142(.A(new_n11490), .B(new_n11427), .Y(new_n11491));
  nand_5 g09143(.A(new_n11491), .B(n24032), .Y(new_n11492));
  nor_5  g09144(.A(new_n11491), .B(n24032), .Y(new_n11493));
  nand_5 g09145(.A(n15936), .B(new_n2614), .Y(new_n11494));
  not_8  g09146(.A(new_n11494), .Y(new_n11495));
  nor_5  g09147(.A(n15936), .B(new_n2614), .Y(new_n11496_1));
  nor_5  g09148(.A(new_n11496_1), .B(new_n11495), .Y(new_n11497));
  not_8  g09149(.A(new_n11497), .Y(new_n11498));
  nand_5 g09150(.A(new_n11498), .B(n22843), .Y(new_n11499));
  or_5   g09151(.A(new_n11499), .B(new_n11493), .Y(new_n11500));
  nand_5 g09152(.A(new_n11500), .B(new_n11492), .Y(new_n11501));
  nand_5 g09153(.A(new_n11501), .B(new_n11489), .Y(new_n11502));
  nand_5 g09154(.A(new_n11502), .B(new_n11488), .Y(new_n11503_1));
  nand_5 g09155(.A(new_n11503_1), .B(new_n11484), .Y(new_n11504));
  nand_5 g09156(.A(new_n11504), .B(new_n11483), .Y(new_n11505));
  nand_5 g09157(.A(new_n11505), .B(new_n11479_1), .Y(new_n11506_1));
  nand_5 g09158(.A(new_n11506_1), .B(new_n11478), .Y(new_n11507));
  nand_5 g09159(.A(new_n11507), .B(new_n11474), .Y(new_n11508));
  nand_5 g09160(.A(new_n11508), .B(new_n11473_1), .Y(new_n11509));
  nand_5 g09161(.A(new_n11509), .B(new_n11469), .Y(new_n11510));
  nand_5 g09162(.A(new_n11510), .B(new_n11468), .Y(new_n11511));
  nand_5 g09163(.A(new_n11511), .B(new_n11464), .Y(new_n11512));
  nand_5 g09164(.A(new_n11512), .B(new_n11463), .Y(new_n11513));
  nand_5 g09165(.A(new_n11513), .B(new_n11458), .Y(new_n11514));
  nand_5 g09166(.A(new_n11514), .B(new_n11457), .Y(new_n11515_1));
  nand_5 g09167(.A(new_n11515_1), .B(new_n11452), .Y(new_n11516));
  nand_5 g09168(.A(new_n11516), .B(new_n11451), .Y(new_n11517));
  nand_5 g09169(.A(new_n11449), .B(new_n11406), .Y(new_n11518));
  nand_5 g09170(.A(new_n11518), .B(new_n11405), .Y(new_n11519));
  not_8  g09171(.A(new_n11519), .Y(new_n11520));
  nand_5 g09172(.A(new_n11520), .B(new_n11517), .Y(new_n11521));
  not_8  g09173(.A(new_n11521), .Y(new_n11522));
  nand_5 g09174(.A(new_n11522), .B(new_n11403_1), .Y(new_n11523));
  or_5   g09175(.A(new_n11522), .B(new_n11403_1), .Y(new_n11524));
  nand_5 g09176(.A(new_n11524), .B(new_n11523), .Y(new_n11525));
  xor_4  g09177(.A(new_n11402), .B(new_n11400), .Y(new_n11526));
  nor_5  g09178(.A(new_n11520), .B(new_n11517), .Y(new_n11527));
  nor_5  g09179(.A(new_n11527), .B(new_n11522), .Y(new_n11528));
  not_8  g09180(.A(new_n11528), .Y(new_n11529));
  and_5  g09181(.A(new_n11529), .B(new_n11526), .Y(new_n11530));
  nor_5  g09182(.A(new_n11529), .B(new_n11526), .Y(new_n11531));
  nor_5  g09183(.A(new_n11339), .B(new_n11338), .Y(new_n11532));
  xor_4  g09184(.A(new_n11532), .B(new_n11397), .Y(new_n11533));
  nand_5 g09185(.A(new_n11452), .B(new_n11451), .Y(new_n11534));
  xor_4  g09186(.A(new_n11534), .B(new_n11515_1), .Y(new_n11535));
  and_5  g09187(.A(new_n11535), .B(new_n11533), .Y(new_n11536));
  nor_5  g09188(.A(new_n11535), .B(new_n11533), .Y(new_n11537));
  nand_5 g09189(.A(new_n11344), .B(new_n11343), .Y(new_n11538_1));
  xor_4  g09190(.A(new_n11538_1), .B(new_n11395), .Y(new_n11539));
  nand_5 g09191(.A(new_n11458), .B(new_n11457), .Y(new_n11540));
  xor_4  g09192(.A(new_n11540), .B(new_n11513), .Y(new_n11541));
  not_8  g09193(.A(new_n11541), .Y(new_n11542));
  nand_5 g09194(.A(new_n11542), .B(new_n11539), .Y(new_n11543));
  or_5   g09195(.A(new_n11542), .B(new_n11539), .Y(new_n11544));
  nand_5 g09196(.A(new_n11349), .B(new_n11348_1), .Y(new_n11545));
  xor_4  g09197(.A(new_n11545), .B(new_n11393), .Y(new_n11546));
  nand_5 g09198(.A(new_n11464), .B(new_n11463), .Y(new_n11547));
  xor_4  g09199(.A(new_n11547), .B(new_n11511), .Y(new_n11548_1));
  not_8  g09200(.A(new_n11548_1), .Y(new_n11549));
  nand_5 g09201(.A(new_n11549), .B(new_n11546), .Y(new_n11550));
  nor_5  g09202(.A(new_n11549), .B(new_n11546), .Y(new_n11551));
  not_8  g09203(.A(new_n11551), .Y(new_n11552));
  nand_5 g09204(.A(new_n11354), .B(new_n11353), .Y(new_n11553));
  xor_4  g09205(.A(new_n11553), .B(new_n11391_1), .Y(new_n11554));
  nand_5 g09206(.A(new_n11469), .B(new_n11468), .Y(new_n11555));
  xor_4  g09207(.A(new_n11555), .B(new_n11509), .Y(new_n11556));
  not_8  g09208(.A(new_n11556), .Y(new_n11557));
  nand_5 g09209(.A(new_n11557), .B(new_n11554), .Y(new_n11558));
  nor_5  g09210(.A(new_n11557), .B(new_n11554), .Y(new_n11559));
  not_8  g09211(.A(new_n11559), .Y(new_n11560));
  nand_5 g09212(.A(new_n11359), .B(new_n11358), .Y(new_n11561));
  xor_4  g09213(.A(new_n11561), .B(new_n11389), .Y(new_n11562));
  nand_5 g09214(.A(new_n11474), .B(new_n11473_1), .Y(new_n11563));
  xor_4  g09215(.A(new_n11563), .B(new_n11507), .Y(new_n11564_1));
  not_8  g09216(.A(new_n11564_1), .Y(new_n11565));
  nand_5 g09217(.A(new_n11565), .B(new_n11562), .Y(new_n11566_1));
  or_5   g09218(.A(new_n11565), .B(new_n11562), .Y(new_n11567));
  nand_5 g09219(.A(new_n11364), .B(new_n11363), .Y(new_n11568));
  xor_4  g09220(.A(new_n11568), .B(new_n11387), .Y(new_n11569));
  nand_5 g09221(.A(new_n11479_1), .B(new_n11478), .Y(new_n11570));
  xor_4  g09222(.A(new_n11570), .B(new_n11505), .Y(new_n11571));
  not_8  g09223(.A(new_n11571), .Y(new_n11572));
  nand_5 g09224(.A(new_n11572), .B(new_n11569), .Y(new_n11573));
  or_5   g09225(.A(new_n11572), .B(new_n11569), .Y(new_n11574));
  nand_5 g09226(.A(new_n11369), .B(new_n11368), .Y(new_n11575));
  xor_4  g09227(.A(new_n11575), .B(new_n11385), .Y(new_n11576));
  nand_5 g09228(.A(new_n11484), .B(new_n11483), .Y(new_n11577));
  xor_4  g09229(.A(new_n11577), .B(new_n11503_1), .Y(new_n11578));
  not_8  g09230(.A(new_n11578), .Y(new_n11579_1));
  nand_5 g09231(.A(new_n11579_1), .B(new_n11576), .Y(new_n11580_1));
  or_5   g09232(.A(new_n11579_1), .B(new_n11576), .Y(new_n11581));
  nand_5 g09233(.A(new_n11373), .B(new_n11372), .Y(new_n11582));
  xor_4  g09234(.A(new_n11582), .B(new_n11383), .Y(new_n11583));
  nand_5 g09235(.A(new_n11489), .B(new_n11488), .Y(new_n11584));
  xor_4  g09236(.A(new_n11584), .B(new_n11501), .Y(new_n11585));
  not_8  g09237(.A(new_n11585), .Y(new_n11586));
  nand_5 g09238(.A(new_n11586), .B(new_n11583), .Y(new_n11587));
  or_5   g09239(.A(new_n11586), .B(new_n11583), .Y(new_n11588));
  nand_5 g09240(.A(new_n11377), .B(new_n11376), .Y(new_n11589));
  xor_4  g09241(.A(new_n11589), .B(new_n11381), .Y(new_n11590));
  not_8  g09242(.A(new_n11493), .Y(new_n11591_1));
  nand_5 g09243(.A(new_n11591_1), .B(new_n11492), .Y(new_n11592));
  xor_4  g09244(.A(new_n11592), .B(new_n11499), .Y(new_n11593));
  nand_5 g09245(.A(new_n11593), .B(new_n11590), .Y(new_n11594));
  nor_5  g09246(.A(new_n11593), .B(new_n11590), .Y(new_n11595));
  not_8  g09247(.A(new_n11595), .Y(new_n11596));
  xor_4  g09248(.A(new_n11380), .B(new_n11378), .Y(new_n11597));
  nand_5 g09249(.A(new_n11497), .B(new_n2622), .Y(new_n11598));
  and_5  g09250(.A(new_n11598), .B(new_n11499), .Y(new_n11599));
  not_8  g09251(.A(new_n11599), .Y(new_n11600));
  nor_5  g09252(.A(new_n11600), .B(new_n11597), .Y(new_n11601));
  nand_5 g09253(.A(new_n11601), .B(new_n11596), .Y(new_n11602));
  nand_5 g09254(.A(new_n11602), .B(new_n11594), .Y(new_n11603));
  nand_5 g09255(.A(new_n11603), .B(new_n11588), .Y(new_n11604));
  nand_5 g09256(.A(new_n11604), .B(new_n11587), .Y(new_n11605));
  nand_5 g09257(.A(new_n11605), .B(new_n11581), .Y(new_n11606));
  nand_5 g09258(.A(new_n11606), .B(new_n11580_1), .Y(new_n11607_1));
  nand_5 g09259(.A(new_n11607_1), .B(new_n11574), .Y(new_n11608));
  nand_5 g09260(.A(new_n11608), .B(new_n11573), .Y(new_n11609));
  nand_5 g09261(.A(new_n11609), .B(new_n11567), .Y(new_n11610));
  nand_5 g09262(.A(new_n11610), .B(new_n11566_1), .Y(new_n11611));
  nand_5 g09263(.A(new_n11611), .B(new_n11560), .Y(new_n11612));
  nand_5 g09264(.A(new_n11612), .B(new_n11558), .Y(new_n11613));
  nand_5 g09265(.A(new_n11613), .B(new_n11552), .Y(new_n11614));
  nand_5 g09266(.A(new_n11614), .B(new_n11550), .Y(new_n11615_1));
  nand_5 g09267(.A(new_n11615_1), .B(new_n11544), .Y(new_n11616));
  nand_5 g09268(.A(new_n11616), .B(new_n11543), .Y(new_n11617));
  nor_5  g09269(.A(new_n11617), .B(new_n11537), .Y(new_n11618));
  nor_5  g09270(.A(new_n11618), .B(new_n11536), .Y(new_n11619));
  nor_5  g09271(.A(new_n11619), .B(new_n11531), .Y(new_n11620));
  nor_5  g09272(.A(new_n11620), .B(new_n11530), .Y(new_n11621));
  xor_4  g09273(.A(new_n11621), .B(new_n11525), .Y(n1302));
  not_8  g09274(.A(n11220), .Y(new_n11623));
  nand_5 g09275(.A(new_n10314), .B(new_n11623), .Y(new_n11624));
  nand_5 g09276(.A(new_n3276), .B(new_n10318), .Y(new_n11625));
  nand_5 g09277(.A(new_n10321_1), .B(new_n3030_1), .Y(new_n11626));
  nand_5 g09278(.A(new_n10824), .B(new_n10822), .Y(new_n11627));
  nand_5 g09279(.A(new_n11627), .B(new_n10823), .Y(new_n11628));
  nand_5 g09280(.A(n10593), .B(n1662), .Y(new_n11629));
  nand_5 g09281(.A(new_n11629), .B(new_n11628), .Y(new_n11630_1));
  nand_5 g09282(.A(new_n11630_1), .B(new_n11626), .Y(new_n11631));
  nand_5 g09283(.A(n22379), .B(n10201), .Y(new_n11632));
  nand_5 g09284(.A(new_n11632), .B(new_n11631), .Y(new_n11633));
  nand_5 g09285(.A(new_n11633), .B(new_n11625), .Y(new_n11634));
  nand_5 g09286(.A(n12650), .B(n11220), .Y(new_n11635));
  nand_5 g09287(.A(new_n11635), .B(new_n11634), .Y(new_n11636));
  nand_5 g09288(.A(new_n11636), .B(new_n11624), .Y(new_n11637));
  not_8  g09289(.A(new_n11637), .Y(new_n11638));
  nand_5 g09290(.A(new_n2839), .B(new_n2780), .Y(new_n11639));
  nand_5 g09291(.A(new_n11639), .B(new_n2783_1), .Y(new_n11640));
  nand_5 g09292(.A(new_n11640), .B(new_n11638), .Y(new_n11641));
  not_8  g09293(.A(new_n11640), .Y(new_n11642));
  nand_5 g09294(.A(new_n11642), .B(new_n11637), .Y(new_n11643));
  nand_5 g09295(.A(new_n11643), .B(new_n11641), .Y(new_n11644));
  nand_5 g09296(.A(new_n11635), .B(new_n11624), .Y(new_n11645));
  xor_4  g09297(.A(new_n11645), .B(new_n11634), .Y(new_n11646));
  not_8  g09298(.A(new_n11646), .Y(new_n11647_1));
  nand_5 g09299(.A(new_n11647_1), .B(new_n2840), .Y(new_n11648));
  nand_5 g09300(.A(new_n11646), .B(new_n2841), .Y(new_n11649));
  nand_5 g09301(.A(new_n11632), .B(new_n11625), .Y(new_n11650));
  xor_4  g09302(.A(new_n11650), .B(new_n11631), .Y(new_n11651));
  not_8  g09303(.A(new_n11651), .Y(new_n11652));
  nand_5 g09304(.A(new_n11652), .B(new_n11234_1), .Y(new_n11653));
  nand_5 g09305(.A(new_n11651), .B(new_n2848), .Y(new_n11654));
  nand_5 g09306(.A(new_n11629), .B(new_n11626), .Y(new_n11655));
  xor_4  g09307(.A(new_n11655), .B(new_n11628), .Y(new_n11656));
  not_8  g09308(.A(new_n11656), .Y(new_n11657));
  nand_5 g09309(.A(new_n11657), .B(new_n11160), .Y(new_n11658));
  nand_5 g09310(.A(new_n11656), .B(new_n2853_1), .Y(new_n11659));
  nand_5 g09311(.A(new_n10828), .B(new_n11119), .Y(new_n11660));
  nand_5 g09312(.A(new_n10826), .B(new_n2858_1), .Y(new_n11661));
  nand_5 g09313(.A(new_n10709), .B(new_n11129), .Y(new_n11662));
  nand_5 g09314(.A(new_n10710_1), .B(new_n2864), .Y(new_n11663));
  nand_5 g09315(.A(new_n10672), .B(new_n11134_1), .Y(new_n11664));
  nand_5 g09316(.A(new_n10673), .B(new_n2869), .Y(new_n11665));
  nand_5 g09317(.A(new_n10679), .B(new_n2875), .Y(new_n11666));
  nand_5 g09318(.A(new_n10677), .B(new_n2874), .Y(new_n11667_1));
  nand_5 g09319(.A(new_n10684), .B(new_n2883), .Y(new_n11668));
  nand_5 g09320(.A(new_n10682), .B(new_n2884), .Y(new_n11669));
  nand_5 g09321(.A(new_n10689), .B(new_n2889), .Y(new_n11670));
  nand_5 g09322(.A(new_n10687), .B(new_n2890), .Y(new_n11671));
  nand_5 g09323(.A(new_n10804), .B(new_n2893), .Y(new_n11672));
  not_8  g09324(.A(new_n11672), .Y(new_n11673));
  nand_5 g09325(.A(new_n11673), .B(new_n11671), .Y(new_n11674_1));
  nand_5 g09326(.A(new_n11674_1), .B(new_n11670), .Y(new_n11675));
  nand_5 g09327(.A(new_n11675), .B(new_n11669), .Y(new_n11676));
  nand_5 g09328(.A(new_n11676), .B(new_n11668), .Y(new_n11677));
  nand_5 g09329(.A(new_n11677), .B(new_n11667_1), .Y(new_n11678));
  nand_5 g09330(.A(new_n11678), .B(new_n11666), .Y(new_n11679));
  nand_5 g09331(.A(new_n11679), .B(new_n11665), .Y(new_n11680));
  nand_5 g09332(.A(new_n11680), .B(new_n11664), .Y(new_n11681));
  nand_5 g09333(.A(new_n11681), .B(new_n11663), .Y(new_n11682_1));
  nand_5 g09334(.A(new_n11682_1), .B(new_n11662), .Y(new_n11683));
  nand_5 g09335(.A(new_n11683), .B(new_n11661), .Y(new_n11684));
  nand_5 g09336(.A(new_n11684), .B(new_n11660), .Y(new_n11685));
  nand_5 g09337(.A(new_n11685), .B(new_n11659), .Y(new_n11686));
  nand_5 g09338(.A(new_n11686), .B(new_n11658), .Y(new_n11687));
  nand_5 g09339(.A(new_n11687), .B(new_n11654), .Y(new_n11688));
  nand_5 g09340(.A(new_n11688), .B(new_n11653), .Y(new_n11689));
  nand_5 g09341(.A(new_n11689), .B(new_n11649), .Y(new_n11690));
  nand_5 g09342(.A(new_n11690), .B(new_n11648), .Y(new_n11691));
  xor_4  g09343(.A(new_n11691), .B(new_n11644), .Y(new_n11692));
  not_8  g09344(.A(new_n11692), .Y(new_n11693));
  not_8  g09345(.A(n13951), .Y(new_n11694));
  nand_5 g09346(.A(new_n11694), .B(n12507), .Y(new_n11695));
  not_8  g09347(.A(n12507), .Y(new_n11696));
  nand_5 g09348(.A(n13951), .B(new_n11696), .Y(new_n11697));
  nand_5 g09349(.A(new_n2766), .B(n15077), .Y(new_n11698));
  not_8  g09350(.A(n15077), .Y(new_n11699));
  nand_5 g09351(.A(n22793), .B(new_n11699), .Y(new_n11700));
  not_8  g09352(.A(n8439), .Y(new_n11701));
  nand_5 g09353(.A(new_n11701), .B(n3710), .Y(new_n11702));
  not_8  g09354(.A(n3710), .Y(new_n11703));
  nand_5 g09355(.A(n8439), .B(new_n11703), .Y(new_n11704));
  nand_5 g09356(.A(n26318), .B(new_n2767), .Y(new_n11705));
  not_8  g09357(.A(n26318), .Y(new_n11706));
  nand_5 g09358(.A(new_n11706), .B(n25523), .Y(new_n11707));
  not_8  g09359(.A(n5579), .Y(new_n11708));
  nand_5 g09360(.A(n26054), .B(new_n11708), .Y(new_n11709));
  not_8  g09361(.A(n26054), .Y(new_n11710_1));
  nand_5 g09362(.A(new_n11710_1), .B(n5579), .Y(new_n11711));
  nand_5 g09363(.A(new_n2768), .B(n19081), .Y(new_n11712_1));
  not_8  g09364(.A(n19081), .Y(new_n11713));
  nand_5 g09365(.A(n23430), .B(new_n11713), .Y(new_n11714));
  nand_5 g09366(.A(new_n2876), .B(n8309), .Y(new_n11715));
  not_8  g09367(.A(n8309), .Y(new_n11716));
  nand_5 g09368(.A(n10411), .B(new_n11716), .Y(new_n11717));
  not_8  g09369(.A(n16971), .Y(new_n11718));
  nand_5 g09370(.A(n19144), .B(new_n11718), .Y(new_n11719));
  not_8  g09371(.A(n19144), .Y(new_n11720));
  nand_5 g09372(.A(new_n11720), .B(n16971), .Y(new_n11721));
  nand_5 g09373(.A(n12593), .B(new_n2769), .Y(new_n11722));
  not_8  g09374(.A(n12593), .Y(new_n11723));
  nand_5 g09375(.A(new_n11723), .B(n11503), .Y(new_n11724_1));
  nand_5 g09376(.A(n18151), .B(new_n10138), .Y(new_n11725));
  nand_5 g09377(.A(new_n11725), .B(new_n11724_1), .Y(new_n11726));
  nand_5 g09378(.A(new_n11726), .B(new_n11722), .Y(new_n11727));
  nand_5 g09379(.A(new_n11727), .B(new_n11721), .Y(new_n11728));
  nand_5 g09380(.A(new_n11728), .B(new_n11719), .Y(new_n11729));
  nand_5 g09381(.A(new_n11729), .B(new_n11717), .Y(new_n11730));
  nand_5 g09382(.A(new_n11730), .B(new_n11715), .Y(new_n11731));
  nand_5 g09383(.A(new_n11731), .B(new_n11714), .Y(new_n11732));
  nand_5 g09384(.A(new_n11732), .B(new_n11712_1), .Y(new_n11733));
  nand_5 g09385(.A(new_n11733), .B(new_n11711), .Y(new_n11734));
  nand_5 g09386(.A(new_n11734), .B(new_n11709), .Y(new_n11735));
  nand_5 g09387(.A(new_n11735), .B(new_n11707), .Y(new_n11736_1));
  nand_5 g09388(.A(new_n11736_1), .B(new_n11705), .Y(new_n11737));
  nand_5 g09389(.A(new_n11737), .B(new_n11704), .Y(new_n11738));
  nand_5 g09390(.A(new_n11738), .B(new_n11702), .Y(new_n11739));
  nand_5 g09391(.A(new_n11739), .B(new_n11700), .Y(new_n11740));
  nand_5 g09392(.A(new_n11740), .B(new_n11698), .Y(new_n11741_1));
  nand_5 g09393(.A(new_n11741_1), .B(new_n11697), .Y(new_n11742));
  nand_5 g09394(.A(new_n11742), .B(new_n11695), .Y(new_n11743));
  nor_5  g09395(.A(new_n11743), .B(new_n11693), .Y(new_n11744));
  not_8  g09396(.A(new_n11743), .Y(new_n11745));
  nor_5  g09397(.A(new_n11745), .B(new_n11692), .Y(new_n11746));
  or_5   g09398(.A(new_n11746), .B(new_n11744), .Y(new_n11747));
  nand_5 g09399(.A(new_n11697), .B(new_n11695), .Y(new_n11748));
  xor_4  g09400(.A(new_n11748), .B(new_n11741_1), .Y(new_n11749_1));
  nand_5 g09401(.A(new_n11648), .B(new_n11649), .Y(new_n11750));
  xor_4  g09402(.A(new_n11750), .B(new_n11689), .Y(new_n11751));
  not_8  g09403(.A(new_n11751), .Y(new_n11752));
  nand_5 g09404(.A(new_n11752), .B(new_n11749_1), .Y(new_n11753));
  or_5   g09405(.A(new_n11752), .B(new_n11749_1), .Y(new_n11754));
  nand_5 g09406(.A(new_n11700), .B(new_n11698), .Y(new_n11755));
  xor_4  g09407(.A(new_n11755), .B(new_n11739), .Y(new_n11756));
  nand_5 g09408(.A(new_n11653), .B(new_n11654), .Y(new_n11757));
  xor_4  g09409(.A(new_n11757), .B(new_n11687), .Y(new_n11758));
  not_8  g09410(.A(new_n11758), .Y(new_n11759));
  nand_5 g09411(.A(new_n11759), .B(new_n11756), .Y(new_n11760));
  or_5   g09412(.A(new_n11759), .B(new_n11756), .Y(new_n11761));
  nand_5 g09413(.A(new_n11704), .B(new_n11702), .Y(new_n11762));
  xor_4  g09414(.A(new_n11762), .B(new_n11737), .Y(new_n11763));
  nand_5 g09415(.A(new_n11658), .B(new_n11659), .Y(new_n11764));
  xor_4  g09416(.A(new_n11764), .B(new_n11685), .Y(new_n11765));
  not_8  g09417(.A(new_n11765), .Y(new_n11766));
  nand_5 g09418(.A(new_n11766), .B(new_n11763), .Y(new_n11767));
  or_5   g09419(.A(new_n11766), .B(new_n11763), .Y(new_n11768));
  nand_5 g09420(.A(new_n11707), .B(new_n11705), .Y(new_n11769));
  xor_4  g09421(.A(new_n11769), .B(new_n11735), .Y(new_n11770_1));
  nand_5 g09422(.A(new_n11660), .B(new_n11661), .Y(new_n11771_1));
  xor_4  g09423(.A(new_n11771_1), .B(new_n11683), .Y(new_n11772));
  not_8  g09424(.A(new_n11772), .Y(new_n11773));
  nand_5 g09425(.A(new_n11773), .B(new_n11770_1), .Y(new_n11774));
  or_5   g09426(.A(new_n11773), .B(new_n11770_1), .Y(new_n11775_1));
  nand_5 g09427(.A(new_n11711), .B(new_n11709), .Y(new_n11776));
  xor_4  g09428(.A(new_n11776), .B(new_n11733), .Y(new_n11777));
  nand_5 g09429(.A(new_n11662), .B(new_n11663), .Y(new_n11778));
  xor_4  g09430(.A(new_n11778), .B(new_n11681), .Y(new_n11779));
  not_8  g09431(.A(new_n11779), .Y(new_n11780));
  nand_5 g09432(.A(new_n11780), .B(new_n11777), .Y(new_n11781));
  or_5   g09433(.A(new_n11780), .B(new_n11777), .Y(new_n11782));
  nand_5 g09434(.A(new_n11714), .B(new_n11712_1), .Y(new_n11783));
  xor_4  g09435(.A(new_n11783), .B(new_n11731), .Y(new_n11784));
  nand_5 g09436(.A(new_n11664), .B(new_n11665), .Y(new_n11785));
  xor_4  g09437(.A(new_n11785), .B(new_n11679), .Y(new_n11786));
  not_8  g09438(.A(new_n11786), .Y(new_n11787));
  nand_5 g09439(.A(new_n11787), .B(new_n11784), .Y(new_n11788));
  or_5   g09440(.A(new_n11787), .B(new_n11784), .Y(new_n11789));
  nand_5 g09441(.A(new_n11717), .B(new_n11715), .Y(new_n11790));
  xor_4  g09442(.A(new_n11790), .B(new_n11729), .Y(new_n11791));
  nand_5 g09443(.A(new_n11666), .B(new_n11667_1), .Y(new_n11792));
  xor_4  g09444(.A(new_n11792), .B(new_n11677), .Y(new_n11793));
  not_8  g09445(.A(new_n11793), .Y(new_n11794));
  nand_5 g09446(.A(new_n11794), .B(new_n11791), .Y(new_n11795));
  nor_5  g09447(.A(new_n11794), .B(new_n11791), .Y(new_n11796));
  not_8  g09448(.A(new_n11796), .Y(new_n11797));
  nand_5 g09449(.A(new_n11721), .B(new_n11719), .Y(new_n11798));
  xor_4  g09450(.A(new_n11798), .B(new_n11727), .Y(new_n11799));
  nand_5 g09451(.A(new_n11668), .B(new_n11669), .Y(new_n11800));
  xor_4  g09452(.A(new_n11800), .B(new_n11675), .Y(new_n11801));
  not_8  g09453(.A(new_n11801), .Y(new_n11802));
  or_5   g09454(.A(new_n11802), .B(new_n11799), .Y(new_n11803));
  nand_5 g09455(.A(new_n11802), .B(new_n11799), .Y(new_n11804));
  xor_4  g09456(.A(new_n10692_1), .B(new_n2893), .Y(new_n11805));
  nand_5 g09457(.A(new_n2770), .B(n13714), .Y(new_n11806));
  nand_5 g09458(.A(new_n11806), .B(new_n11725), .Y(new_n11807));
  nand_5 g09459(.A(new_n11807), .B(new_n11805), .Y(new_n11808));
  not_8  g09460(.A(new_n11725), .Y(new_n11809));
  and_5  g09461(.A(new_n11724_1), .B(new_n11722), .Y(new_n11810));
  xor_4  g09462(.A(new_n11810), .B(new_n11809), .Y(new_n11811));
  or_5   g09463(.A(new_n11811), .B(new_n11808), .Y(new_n11812));
  nand_5 g09464(.A(new_n11811), .B(new_n11808), .Y(new_n11813));
  nand_5 g09465(.A(new_n11670), .B(new_n11671), .Y(new_n11814));
  xor_4  g09466(.A(new_n11814), .B(new_n11673), .Y(new_n11815));
  nand_5 g09467(.A(new_n11815), .B(new_n11813), .Y(new_n11816));
  nand_5 g09468(.A(new_n11816), .B(new_n11812), .Y(new_n11817));
  nand_5 g09469(.A(new_n11817), .B(new_n11804), .Y(new_n11818_1));
  nand_5 g09470(.A(new_n11818_1), .B(new_n11803), .Y(new_n11819));
  not_8  g09471(.A(new_n11819), .Y(new_n11820));
  nand_5 g09472(.A(new_n11820), .B(new_n11797), .Y(new_n11821));
  nand_5 g09473(.A(new_n11821), .B(new_n11795), .Y(new_n11822));
  nand_5 g09474(.A(new_n11822), .B(new_n11789), .Y(new_n11823));
  nand_5 g09475(.A(new_n11823), .B(new_n11788), .Y(new_n11824));
  nand_5 g09476(.A(new_n11824), .B(new_n11782), .Y(new_n11825));
  nand_5 g09477(.A(new_n11825), .B(new_n11781), .Y(new_n11826));
  nand_5 g09478(.A(new_n11826), .B(new_n11775_1), .Y(new_n11827));
  nand_5 g09479(.A(new_n11827), .B(new_n11774), .Y(new_n11828));
  nand_5 g09480(.A(new_n11828), .B(new_n11768), .Y(new_n11829));
  nand_5 g09481(.A(new_n11829), .B(new_n11767), .Y(new_n11830));
  nand_5 g09482(.A(new_n11830), .B(new_n11761), .Y(new_n11831));
  nand_5 g09483(.A(new_n11831), .B(new_n11760), .Y(new_n11832));
  nand_5 g09484(.A(new_n11832), .B(new_n11754), .Y(new_n11833));
  nand_5 g09485(.A(new_n11833), .B(new_n11753), .Y(new_n11834));
  xor_4  g09486(.A(new_n11834), .B(new_n11747), .Y(n1332));
  nand_5 g09487(.A(new_n6593), .B(new_n4376_1), .Y(new_n11836));
  nor_5  g09488(.A(new_n11836), .B(n10405), .Y(new_n11837_1));
  nand_5 g09489(.A(new_n11837_1), .B(new_n4438), .Y(new_n11838));
  nor_5  g09490(.A(new_n11838), .B(n20151), .Y(new_n11839));
  nand_5 g09491(.A(new_n11839), .B(new_n6394), .Y(new_n11840));
  nor_5  g09492(.A(new_n11840), .B(n27037), .Y(new_n11841_1));
  nand_5 g09493(.A(new_n11841_1), .B(new_n6386), .Y(new_n11842_1));
  xor_4  g09494(.A(new_n11842_1), .B(n8614), .Y(new_n11843_1));
  not_8  g09495(.A(new_n11843_1), .Y(new_n11844));
  or_5   g09496(.A(new_n6585), .B(n5330), .Y(new_n11845));
  nor_5  g09497(.A(new_n11845), .B(n5451), .Y(new_n11846));
  nand_5 g09498(.A(new_n11846), .B(new_n4359), .Y(new_n11847));
  nor_5  g09499(.A(new_n11847), .B(n13677), .Y(new_n11848));
  nand_5 g09500(.A(new_n11848), .B(new_n7179), .Y(new_n11849));
  nor_5  g09501(.A(new_n11849), .B(n7692), .Y(new_n11850));
  nand_5 g09502(.A(new_n11850), .B(new_n7171), .Y(new_n11851));
  nand_5 g09503(.A(new_n11851), .B(n15766), .Y(new_n11852));
  nor_5  g09504(.A(new_n11851), .B(n15766), .Y(new_n11853));
  not_8  g09505(.A(new_n11853), .Y(new_n11854));
  and_5  g09506(.A(new_n11854), .B(new_n11852), .Y(new_n11855));
  nand_5 g09507(.A(new_n11855), .B(n23895), .Y(new_n11856));
  not_8  g09508(.A(new_n11855), .Y(new_n11857));
  nand_5 g09509(.A(new_n11857), .B(new_n6384), .Y(new_n11858));
  nand_5 g09510(.A(new_n11858), .B(new_n11856), .Y(new_n11859));
  xor_4  g09511(.A(new_n11850), .B(new_n7171), .Y(new_n11860));
  not_8  g09512(.A(new_n11860), .Y(new_n11861));
  nand_5 g09513(.A(new_n11861), .B(new_n6388), .Y(new_n11862));
  nand_5 g09514(.A(new_n11860), .B(n17351), .Y(new_n11863));
  xor_4  g09515(.A(new_n11849), .B(n7692), .Y(new_n11864));
  not_8  g09516(.A(new_n11864), .Y(new_n11865));
  nand_5 g09517(.A(new_n11865), .B(new_n6392), .Y(new_n11866));
  nand_5 g09518(.A(new_n11864), .B(n11736), .Y(new_n11867));
  xor_4  g09519(.A(new_n11848), .B(new_n7179), .Y(new_n11868));
  not_8  g09520(.A(new_n11868), .Y(new_n11869));
  nand_5 g09521(.A(new_n11869), .B(new_n6396), .Y(new_n11870));
  nand_5 g09522(.A(new_n11868), .B(n23200), .Y(new_n11871));
  xor_4  g09523(.A(new_n11847), .B(n13677), .Y(new_n11872));
  not_8  g09524(.A(new_n11872), .Y(new_n11873));
  nand_5 g09525(.A(new_n11873), .B(new_n6399), .Y(new_n11874));
  nand_5 g09526(.A(new_n11872), .B(n17959), .Y(new_n11875));
  xor_4  g09527(.A(new_n11846), .B(new_n4359), .Y(new_n11876));
  not_8  g09528(.A(new_n11876), .Y(new_n11877));
  nand_5 g09529(.A(new_n11877), .B(new_n6402), .Y(new_n11878));
  nand_5 g09530(.A(new_n11876), .B(n7566), .Y(new_n11879));
  xor_4  g09531(.A(new_n11845), .B(n5451), .Y(new_n11880));
  not_8  g09532(.A(new_n11880), .Y(new_n11881));
  nand_5 g09533(.A(new_n11881), .B(new_n6405), .Y(new_n11882));
  nand_5 g09534(.A(new_n11880), .B(n7731), .Y(new_n11883));
  nand_5 g09535(.A(new_n6585), .B(n5330), .Y(new_n11884));
  and_5  g09536(.A(new_n11884), .B(new_n11845), .Y(new_n11885));
  not_8  g09537(.A(new_n11885), .Y(new_n11886));
  nand_5 g09538(.A(new_n11886), .B(new_n6408), .Y(new_n11887));
  nand_5 g09539(.A(new_n11885), .B(n12341), .Y(new_n11888));
  nand_5 g09540(.A(new_n6590_1), .B(new_n6577), .Y(new_n11889));
  nand_5 g09541(.A(new_n11889), .B(new_n6589), .Y(new_n11890));
  nand_5 g09542(.A(new_n11890), .B(new_n11888), .Y(new_n11891));
  nand_5 g09543(.A(new_n11891), .B(new_n11887), .Y(new_n11892));
  nand_5 g09544(.A(new_n11892), .B(new_n11883), .Y(new_n11893));
  nand_5 g09545(.A(new_n11893), .B(new_n11882), .Y(new_n11894));
  nand_5 g09546(.A(new_n11894), .B(new_n11879), .Y(new_n11895));
  nand_5 g09547(.A(new_n11895), .B(new_n11878), .Y(new_n11896));
  nand_5 g09548(.A(new_n11896), .B(new_n11875), .Y(new_n11897));
  nand_5 g09549(.A(new_n11897), .B(new_n11874), .Y(new_n11898_1));
  nand_5 g09550(.A(new_n11898_1), .B(new_n11871), .Y(new_n11899));
  nand_5 g09551(.A(new_n11899), .B(new_n11870), .Y(new_n11900));
  nand_5 g09552(.A(new_n11900), .B(new_n11867), .Y(new_n11901));
  nand_5 g09553(.A(new_n11901), .B(new_n11866), .Y(new_n11902));
  nand_5 g09554(.A(new_n11902), .B(new_n11863), .Y(new_n11903));
  nand_5 g09555(.A(new_n11903), .B(new_n11862), .Y(new_n11904));
  not_8  g09556(.A(new_n11904), .Y(new_n11905_1));
  xor_4  g09557(.A(new_n11905_1), .B(new_n11859), .Y(new_n11906));
  nand_5 g09558(.A(new_n11906), .B(new_n11844), .Y(new_n11907));
  xor_4  g09559(.A(new_n11841_1), .B(new_n6386), .Y(new_n11908));
  nand_5 g09560(.A(new_n11863), .B(new_n11862), .Y(new_n11909));
  xor_4  g09561(.A(new_n11909), .B(new_n11902), .Y(new_n11910));
  nand_5 g09562(.A(new_n11910), .B(new_n11908), .Y(new_n11911));
  or_5   g09563(.A(new_n11910), .B(new_n11908), .Y(new_n11912));
  xor_4  g09564(.A(new_n11840), .B(n27037), .Y(new_n11913));
  nand_5 g09565(.A(new_n11867), .B(new_n11866), .Y(new_n11914));
  xor_4  g09566(.A(new_n11914), .B(new_n11900), .Y(new_n11915));
  nand_5 g09567(.A(new_n11915), .B(new_n11913), .Y(new_n11916));
  or_5   g09568(.A(new_n11915), .B(new_n11913), .Y(new_n11917));
  xor_4  g09569(.A(new_n11839), .B(new_n6394), .Y(new_n11918));
  nand_5 g09570(.A(new_n11871), .B(new_n11870), .Y(new_n11919));
  xor_4  g09571(.A(new_n11919), .B(new_n11898_1), .Y(new_n11920));
  nand_5 g09572(.A(new_n11920), .B(new_n11918), .Y(new_n11921));
  or_5   g09573(.A(new_n11920), .B(new_n11918), .Y(new_n11922));
  xor_4  g09574(.A(new_n11838), .B(n20151), .Y(new_n11923));
  nand_5 g09575(.A(new_n11875), .B(new_n11874), .Y(new_n11924));
  xor_4  g09576(.A(new_n11924), .B(new_n11896), .Y(new_n11925));
  nand_5 g09577(.A(new_n11925), .B(new_n11923), .Y(new_n11926_1));
  nor_5  g09578(.A(new_n11925), .B(new_n11923), .Y(new_n11927));
  not_8  g09579(.A(new_n11927), .Y(new_n11928));
  xor_4  g09580(.A(new_n11837_1), .B(new_n4438), .Y(new_n11929));
  nand_5 g09581(.A(new_n11879), .B(new_n11878), .Y(new_n11930));
  xor_4  g09582(.A(new_n11930), .B(new_n11894), .Y(new_n11931));
  nand_5 g09583(.A(new_n11931), .B(new_n11929), .Y(new_n11932));
  nor_5  g09584(.A(new_n11931), .B(new_n11929), .Y(new_n11933));
  not_8  g09585(.A(new_n11933), .Y(new_n11934));
  xor_4  g09586(.A(new_n11836), .B(new_n4396), .Y(new_n11935));
  nand_5 g09587(.A(new_n11883), .B(new_n11882), .Y(new_n11936));
  xor_4  g09588(.A(new_n11936), .B(new_n11892), .Y(new_n11937));
  not_8  g09589(.A(new_n11937), .Y(new_n11938));
  or_5   g09590(.A(new_n11938), .B(new_n11935), .Y(new_n11939));
  nand_5 g09591(.A(new_n11938), .B(new_n11935), .Y(new_n11940));
  xor_4  g09592(.A(new_n6593), .B(n11302), .Y(new_n11941));
  nand_5 g09593(.A(new_n11888), .B(new_n11887), .Y(new_n11942));
  xor_4  g09594(.A(new_n11942), .B(new_n11890), .Y(new_n11943));
  not_8  g09595(.A(new_n11943), .Y(new_n11944));
  or_5   g09596(.A(new_n11944), .B(new_n11941), .Y(new_n11945));
  nand_5 g09597(.A(new_n11944), .B(new_n11941), .Y(new_n11946));
  nor_5  g09598(.A(new_n6598), .B(new_n6592), .Y(new_n11947));
  nor_5  g09599(.A(new_n11947), .B(new_n6596_1), .Y(new_n11948));
  nand_5 g09600(.A(new_n11948), .B(new_n11946), .Y(new_n11949));
  nand_5 g09601(.A(new_n11949), .B(new_n11945), .Y(new_n11950));
  nand_5 g09602(.A(new_n11950), .B(new_n11940), .Y(new_n11951));
  nand_5 g09603(.A(new_n11951), .B(new_n11939), .Y(new_n11952));
  nand_5 g09604(.A(new_n11952), .B(new_n11934), .Y(new_n11953));
  nand_5 g09605(.A(new_n11953), .B(new_n11932), .Y(new_n11954));
  nand_5 g09606(.A(new_n11954), .B(new_n11928), .Y(new_n11955));
  nand_5 g09607(.A(new_n11955), .B(new_n11926_1), .Y(new_n11956));
  nand_5 g09608(.A(new_n11956), .B(new_n11922), .Y(new_n11957));
  nand_5 g09609(.A(new_n11957), .B(new_n11921), .Y(new_n11958));
  nand_5 g09610(.A(new_n11958), .B(new_n11917), .Y(new_n11959));
  nand_5 g09611(.A(new_n11959), .B(new_n11916), .Y(new_n11960));
  nand_5 g09612(.A(new_n11960), .B(new_n11912), .Y(new_n11961));
  nand_5 g09613(.A(new_n11961), .B(new_n11911), .Y(new_n11962));
  nand_5 g09614(.A(new_n11962), .B(new_n11907), .Y(new_n11963));
  nor_5  g09615(.A(new_n11842_1), .B(n8614), .Y(new_n11964));
  not_8  g09616(.A(new_n11906), .Y(new_n11965_1));
  nand_5 g09617(.A(new_n11965_1), .B(new_n11843_1), .Y(new_n11966));
  not_8  g09618(.A(new_n11966), .Y(new_n11967));
  nor_5  g09619(.A(new_n11967), .B(new_n11964), .Y(new_n11968));
  nand_5 g09620(.A(new_n11968), .B(new_n11963), .Y(new_n11969));
  nand_5 g09621(.A(new_n11905_1), .B(new_n11858), .Y(new_n11970));
  not_8  g09622(.A(new_n11970), .Y(new_n11971));
  nand_5 g09623(.A(new_n11856), .B(new_n11854), .Y(new_n11972));
  nor_5  g09624(.A(new_n11972), .B(new_n11971), .Y(new_n11973));
  nor_5  g09625(.A(new_n11973), .B(new_n11969), .Y(new_n11974));
  not_8  g09626(.A(new_n11974), .Y(new_n11975));
  not_8  g09627(.A(new_n6379_1), .Y(new_n11976));
  nand_5 g09628(.A(new_n6279), .B(n14692), .Y(new_n11977));
  not_8  g09629(.A(n14692), .Y(new_n11978));
  nand_5 g09630(.A(new_n6280), .B(new_n11978), .Y(new_n11979));
  not_8  g09631(.A(n4100), .Y(new_n11980_1));
  nand_5 g09632(.A(new_n6284), .B(new_n11980_1), .Y(new_n11981));
  nand_5 g09633(.A(new_n6285), .B(n4100), .Y(new_n11982));
  not_8  g09634(.A(n21957), .Y(new_n11983));
  nand_5 g09635(.A(new_n6291), .B(new_n11983), .Y(new_n11984));
  nand_5 g09636(.A(new_n6292), .B(n21957), .Y(new_n11985));
  not_8  g09637(.A(n15761), .Y(new_n11986));
  nand_5 g09638(.A(new_n6299), .B(new_n11986), .Y(new_n11987));
  nand_5 g09639(.A(new_n6300), .B(n15761), .Y(new_n11988));
  not_8  g09640(.A(n11201), .Y(new_n11989));
  nand_5 g09641(.A(new_n6307), .B(new_n11989), .Y(new_n11990));
  nand_5 g09642(.A(new_n6308_1), .B(n11201), .Y(new_n11991));
  not_8  g09643(.A(n18690), .Y(new_n11992));
  nand_5 g09644(.A(new_n6315), .B(new_n11992), .Y(new_n11993));
  nand_5 g09645(.A(new_n6316), .B(n18690), .Y(new_n11994));
  not_8  g09646(.A(n12153), .Y(new_n11995));
  nand_5 g09647(.A(new_n6323_1), .B(new_n11995), .Y(new_n11996));
  nand_5 g09648(.A(new_n6324), .B(n12153), .Y(new_n11997));
  not_8  g09649(.A(n13044), .Y(new_n11998));
  nand_5 g09650(.A(new_n6330_1), .B(new_n11998), .Y(new_n11999));
  nand_5 g09651(.A(new_n6331), .B(n13044), .Y(new_n12000_1));
  nand_5 g09652(.A(new_n6604), .B(new_n6601), .Y(new_n12001));
  nand_5 g09653(.A(new_n12001), .B(new_n6603), .Y(new_n12002));
  nand_5 g09654(.A(new_n12002), .B(new_n12000_1), .Y(new_n12003_1));
  nand_5 g09655(.A(new_n12003_1), .B(new_n11999), .Y(new_n12004));
  nand_5 g09656(.A(new_n12004), .B(new_n11997), .Y(new_n12005));
  nand_5 g09657(.A(new_n12005), .B(new_n11996), .Y(new_n12006));
  nand_5 g09658(.A(new_n12006), .B(new_n11994), .Y(new_n12007));
  nand_5 g09659(.A(new_n12007), .B(new_n11993), .Y(new_n12008));
  nand_5 g09660(.A(new_n12008), .B(new_n11991), .Y(new_n12009));
  nand_5 g09661(.A(new_n12009), .B(new_n11990), .Y(new_n12010));
  nand_5 g09662(.A(new_n12010), .B(new_n11988), .Y(new_n12011_1));
  nand_5 g09663(.A(new_n12011_1), .B(new_n11987), .Y(new_n12012));
  nand_5 g09664(.A(new_n12012), .B(new_n11985), .Y(new_n12013));
  nand_5 g09665(.A(new_n12013), .B(new_n11984), .Y(new_n12014));
  nand_5 g09666(.A(new_n12014), .B(new_n11982), .Y(new_n12015));
  nand_5 g09667(.A(new_n12015), .B(new_n11981), .Y(new_n12016));
  not_8  g09668(.A(new_n12016), .Y(new_n12017));
  nand_5 g09669(.A(new_n12017), .B(new_n11979), .Y(new_n12018));
  nand_5 g09670(.A(new_n12018), .B(new_n11977), .Y(new_n12019));
  nand_5 g09671(.A(new_n12019), .B(new_n11976), .Y(new_n12020));
  nand_5 g09672(.A(new_n12020), .B(new_n11975), .Y(new_n12021));
  not_8  g09673(.A(new_n12020), .Y(new_n12022));
  nand_5 g09674(.A(new_n12022), .B(new_n11974), .Y(new_n12023));
  nand_5 g09675(.A(new_n12023), .B(new_n12021), .Y(new_n12024));
  xor_4  g09676(.A(new_n11973), .B(new_n11969), .Y(new_n12025));
  nor_5  g09677(.A(new_n12019), .B(new_n11976), .Y(new_n12026));
  nor_5  g09678(.A(new_n12026), .B(new_n12022), .Y(new_n12027));
  not_8  g09679(.A(new_n12027), .Y(new_n12028));
  nand_5 g09680(.A(new_n12028), .B(new_n12025), .Y(new_n12029));
  nor_5  g09681(.A(new_n12028), .B(new_n12025), .Y(new_n12030));
  not_8  g09682(.A(new_n12030), .Y(new_n12031));
  nand_5 g09683(.A(new_n11977), .B(new_n11979), .Y(new_n12032));
  xor_4  g09684(.A(new_n12032), .B(new_n12016), .Y(new_n12033));
  and_5  g09685(.A(new_n11966), .B(new_n11907), .Y(new_n12034));
  xor_4  g09686(.A(new_n12034), .B(new_n11962), .Y(new_n12035));
  or_5   g09687(.A(new_n12035), .B(new_n12033), .Y(new_n12036));
  nand_5 g09688(.A(new_n12035), .B(new_n12033), .Y(new_n12037));
  nand_5 g09689(.A(new_n11982), .B(new_n11981), .Y(new_n12038));
  xor_4  g09690(.A(new_n12038), .B(new_n12014), .Y(new_n12039));
  not_8  g09691(.A(new_n12039), .Y(new_n12040));
  nand_5 g09692(.A(new_n11912), .B(new_n11911), .Y(new_n12041));
  xor_4  g09693(.A(new_n12041), .B(new_n11960), .Y(new_n12042));
  nand_5 g09694(.A(new_n12042), .B(new_n12040), .Y(new_n12043));
  or_5   g09695(.A(new_n12042), .B(new_n12040), .Y(new_n12044));
  nand_5 g09696(.A(new_n11985), .B(new_n11984), .Y(new_n12045));
  xor_4  g09697(.A(new_n12045), .B(new_n12012), .Y(new_n12046));
  not_8  g09698(.A(new_n12046), .Y(new_n12047));
  nand_5 g09699(.A(new_n11917), .B(new_n11916), .Y(new_n12048));
  xor_4  g09700(.A(new_n12048), .B(new_n11958), .Y(new_n12049));
  nand_5 g09701(.A(new_n12049), .B(new_n12047), .Y(new_n12050));
  or_5   g09702(.A(new_n12049), .B(new_n12047), .Y(new_n12051));
  nand_5 g09703(.A(new_n11988), .B(new_n11987), .Y(new_n12052));
  xor_4  g09704(.A(new_n12052), .B(new_n12010), .Y(new_n12053));
  not_8  g09705(.A(new_n12053), .Y(new_n12054));
  nand_5 g09706(.A(new_n11922), .B(new_n11921), .Y(new_n12055));
  xor_4  g09707(.A(new_n12055), .B(new_n11956), .Y(new_n12056));
  or_5   g09708(.A(new_n12056), .B(new_n12054), .Y(new_n12057));
  nand_5 g09709(.A(new_n12056), .B(new_n12054), .Y(new_n12058));
  nand_5 g09710(.A(new_n11991), .B(new_n11990), .Y(new_n12059));
  xor_4  g09711(.A(new_n12059), .B(new_n12008), .Y(new_n12060));
  nand_5 g09712(.A(new_n11928), .B(new_n11926_1), .Y(new_n12061));
  xor_4  g09713(.A(new_n12061), .B(new_n11954), .Y(new_n12062));
  not_8  g09714(.A(new_n12062), .Y(new_n12063));
  nand_5 g09715(.A(new_n12063), .B(new_n12060), .Y(new_n12064));
  nor_5  g09716(.A(new_n12063), .B(new_n12060), .Y(new_n12065));
  not_8  g09717(.A(new_n12065), .Y(new_n12066));
  nand_5 g09718(.A(new_n11994), .B(new_n11993), .Y(new_n12067));
  xor_4  g09719(.A(new_n12067), .B(new_n12006), .Y(new_n12068));
  not_8  g09720(.A(new_n12068), .Y(new_n12069));
  nand_5 g09721(.A(new_n11934), .B(new_n11932), .Y(new_n12070));
  xor_4  g09722(.A(new_n12070), .B(new_n11952), .Y(new_n12071));
  or_5   g09723(.A(new_n12071), .B(new_n12069), .Y(new_n12072_1));
  nand_5 g09724(.A(new_n12071), .B(new_n12069), .Y(new_n12073));
  nand_5 g09725(.A(new_n11997), .B(new_n11996), .Y(new_n12074));
  xor_4  g09726(.A(new_n12074), .B(new_n12004), .Y(new_n12075));
  not_8  g09727(.A(new_n12075), .Y(new_n12076));
  nand_5 g09728(.A(new_n11940), .B(new_n11939), .Y(new_n12077));
  xor_4  g09729(.A(new_n12077), .B(new_n11950), .Y(new_n12078));
  or_5   g09730(.A(new_n12078), .B(new_n12076), .Y(new_n12079));
  nand_5 g09731(.A(new_n12078), .B(new_n12076), .Y(new_n12080));
  nand_5 g09732(.A(new_n11946), .B(new_n11945), .Y(new_n12081));
  xor_4  g09733(.A(new_n12081), .B(new_n11948), .Y(new_n12082));
  nand_5 g09734(.A(new_n12000_1), .B(new_n11999), .Y(new_n12083));
  xor_4  g09735(.A(new_n12083), .B(new_n12002), .Y(new_n12084));
  not_8  g09736(.A(new_n12084), .Y(new_n12085));
  nand_5 g09737(.A(new_n12085), .B(new_n12082), .Y(new_n12086));
  or_5   g09738(.A(new_n12085), .B(new_n12082), .Y(new_n12087));
  nand_5 g09739(.A(new_n6608), .B(new_n6584), .Y(new_n12088));
  nand_5 g09740(.A(new_n12088), .B(new_n6607), .Y(new_n12089));
  nand_5 g09741(.A(new_n12089), .B(new_n12087), .Y(new_n12090));
  and_5  g09742(.A(new_n12090), .B(new_n12086), .Y(new_n12091));
  nand_5 g09743(.A(new_n12091), .B(new_n12080), .Y(new_n12092));
  nand_5 g09744(.A(new_n12092), .B(new_n12079), .Y(new_n12093));
  nand_5 g09745(.A(new_n12093), .B(new_n12073), .Y(new_n12094));
  nand_5 g09746(.A(new_n12094), .B(new_n12072_1), .Y(new_n12095));
  nand_5 g09747(.A(new_n12095), .B(new_n12066), .Y(new_n12096));
  nand_5 g09748(.A(new_n12096), .B(new_n12064), .Y(new_n12097));
  nand_5 g09749(.A(new_n12097), .B(new_n12058), .Y(new_n12098));
  and_5  g09750(.A(new_n12098), .B(new_n12057), .Y(new_n12099));
  nand_5 g09751(.A(new_n12099), .B(new_n12051), .Y(new_n12100));
  nand_5 g09752(.A(new_n12100), .B(new_n12050), .Y(new_n12101));
  nand_5 g09753(.A(new_n12101), .B(new_n12044), .Y(new_n12102));
  nand_5 g09754(.A(new_n12102), .B(new_n12043), .Y(new_n12103));
  nand_5 g09755(.A(new_n12103), .B(new_n12037), .Y(new_n12104));
  nand_5 g09756(.A(new_n12104), .B(new_n12036), .Y(new_n12105));
  nand_5 g09757(.A(new_n12105), .B(new_n12031), .Y(new_n12106));
  nand_5 g09758(.A(new_n12106), .B(new_n12029), .Y(new_n12107));
  xor_4  g09759(.A(new_n12107), .B(new_n12024), .Y(n1357));
  nand_5 g09760(.A(new_n9177), .B(n8067), .Y(new_n12109));
  nand_5 g09761(.A(new_n9179), .B(new_n8303), .Y(new_n12110));
  nand_5 g09762(.A(new_n9184), .B(n20923), .Y(new_n12111));
  nand_5 g09763(.A(new_n9183), .B(new_n8306_1), .Y(new_n12112));
  nand_5 g09764(.A(new_n9726_1), .B(new_n9724), .Y(new_n12113_1));
  nand_5 g09765(.A(new_n12113_1), .B(new_n9725), .Y(new_n12114));
  nand_5 g09766(.A(new_n12114), .B(new_n12112), .Y(new_n12115));
  nand_5 g09767(.A(new_n12115), .B(new_n12111), .Y(new_n12116));
  nand_5 g09768(.A(new_n12116), .B(new_n12110), .Y(new_n12117));
  nand_5 g09769(.A(new_n12117), .B(new_n12109), .Y(new_n12118));
  nand_5 g09770(.A(new_n9171), .B(n10125), .Y(new_n12119));
  nand_5 g09771(.A(new_n9173), .B(new_n8300), .Y(new_n12120));
  nand_5 g09772(.A(new_n12120), .B(new_n12119), .Y(new_n12121_1));
  xor_4  g09773(.A(new_n12121_1), .B(new_n12118), .Y(new_n12122));
  nand_5 g09774(.A(new_n4178), .B(new_n10485), .Y(new_n12123));
  nand_5 g09775(.A(n6369), .B(n3164), .Y(new_n12124));
  nand_5 g09776(.A(new_n7622), .B(new_n7618), .Y(new_n12125));
  nand_5 g09777(.A(new_n12125), .B(new_n7621), .Y(new_n12126));
  nand_5 g09778(.A(new_n12126), .B(new_n12124), .Y(new_n12127));
  nand_5 g09779(.A(new_n12127), .B(new_n12123), .Y(new_n12128));
  not_8  g09780(.A(new_n12128), .Y(new_n12129));
  nand_5 g09781(.A(n21134), .B(n11356), .Y(new_n12130));
  nand_5 g09782(.A(new_n8442), .B(new_n10482), .Y(new_n12131_1));
  nand_5 g09783(.A(new_n12131_1), .B(new_n12130), .Y(new_n12132));
  xor_4  g09784(.A(new_n12132), .B(new_n12129), .Y(new_n12133));
  not_8  g09785(.A(new_n12133), .Y(new_n12134));
  nand_5 g09786(.A(new_n12134), .B(n26452), .Y(new_n12135));
  not_8  g09787(.A(n26452), .Y(new_n12136));
  nand_5 g09788(.A(new_n12133), .B(new_n12136), .Y(new_n12137));
  nand_5 g09789(.A(new_n12124), .B(new_n12123), .Y(new_n12138));
  xor_4  g09790(.A(new_n12138), .B(new_n12126), .Y(new_n12139));
  nand_5 g09791(.A(new_n12139), .B(n19905), .Y(new_n12140));
  not_8  g09792(.A(new_n12139), .Y(new_n12141));
  nand_5 g09793(.A(new_n12141), .B(new_n4768), .Y(new_n12142));
  nand_5 g09794(.A(new_n9685), .B(new_n9683), .Y(new_n12143));
  nand_5 g09795(.A(new_n12143), .B(new_n9684), .Y(new_n12144));
  nand_5 g09796(.A(new_n12144), .B(new_n12142), .Y(new_n12145));
  nand_5 g09797(.A(new_n12145), .B(new_n12140), .Y(new_n12146_1));
  nand_5 g09798(.A(new_n12146_1), .B(new_n12137), .Y(new_n12147));
  nand_5 g09799(.A(new_n12147), .B(new_n12135), .Y(new_n12148));
  nand_5 g09800(.A(new_n12130), .B(new_n12128), .Y(new_n12149));
  nand_5 g09801(.A(new_n12149), .B(new_n12131_1), .Y(new_n12150));
  not_8  g09802(.A(new_n12150), .Y(new_n12151));
  nand_5 g09803(.A(n14345), .B(n2113), .Y(new_n12152_1));
  nand_5 g09804(.A(new_n10479), .B(new_n4298), .Y(new_n12153_1));
  nand_5 g09805(.A(new_n12153_1), .B(new_n12152_1), .Y(new_n12154));
  xor_4  g09806(.A(new_n12154), .B(new_n12151), .Y(new_n12155));
  not_8  g09807(.A(new_n12155), .Y(new_n12156));
  nand_5 g09808(.A(new_n12156), .B(n15546), .Y(new_n12157_1));
  not_8  g09809(.A(n15546), .Y(new_n12158_1));
  nand_5 g09810(.A(new_n12155), .B(new_n12158_1), .Y(new_n12159));
  nand_5 g09811(.A(new_n12159), .B(new_n12157_1), .Y(new_n12160));
  xor_4  g09812(.A(new_n12160), .B(new_n12148), .Y(new_n12161_1));
  not_8  g09813(.A(new_n12161_1), .Y(new_n12162));
  nand_5 g09814(.A(new_n12162), .B(new_n12122), .Y(new_n12163));
  nor_5  g09815(.A(new_n12162), .B(new_n12122), .Y(new_n12164));
  not_8  g09816(.A(new_n12164), .Y(new_n12165));
  nand_5 g09817(.A(new_n12109), .B(new_n12110), .Y(new_n12166));
  xor_4  g09818(.A(new_n12166), .B(new_n12116), .Y(new_n12167));
  nand_5 g09819(.A(new_n12135), .B(new_n12137), .Y(new_n12168));
  xor_4  g09820(.A(new_n12168), .B(new_n12146_1), .Y(new_n12169));
  not_8  g09821(.A(new_n12169), .Y(new_n12170));
  nand_5 g09822(.A(new_n12170), .B(new_n12167), .Y(new_n12171));
  nor_5  g09823(.A(new_n12170), .B(new_n12167), .Y(new_n12172));
  not_8  g09824(.A(new_n12172), .Y(new_n12173));
  nand_5 g09825(.A(new_n12111), .B(new_n12112), .Y(new_n12174));
  xor_4  g09826(.A(new_n12174), .B(new_n12114), .Y(new_n12175));
  nand_5 g09827(.A(new_n12140), .B(new_n12142), .Y(new_n12176));
  xor_4  g09828(.A(new_n12176), .B(new_n12144), .Y(new_n12177));
  not_8  g09829(.A(new_n12177), .Y(new_n12178));
  nand_5 g09830(.A(new_n12178), .B(new_n12175), .Y(new_n12179_1));
  nor_5  g09831(.A(new_n12178), .B(new_n12175), .Y(new_n12180));
  not_8  g09832(.A(new_n12180), .Y(new_n12181));
  nand_5 g09833(.A(new_n9732), .B(new_n9688), .Y(new_n12182));
  nand_5 g09834(.A(new_n12182), .B(new_n9730), .Y(new_n12183));
  nand_5 g09835(.A(new_n12183), .B(new_n12181), .Y(new_n12184));
  nand_5 g09836(.A(new_n12184), .B(new_n12179_1), .Y(new_n12185));
  nand_5 g09837(.A(new_n12185), .B(new_n12173), .Y(new_n12186));
  nand_5 g09838(.A(new_n12186), .B(new_n12171), .Y(new_n12187));
  nand_5 g09839(.A(new_n12187), .B(new_n12165), .Y(new_n12188));
  nand_5 g09840(.A(new_n12188), .B(new_n12163), .Y(new_n12189));
  nand_5 g09841(.A(new_n12120), .B(new_n12118), .Y(new_n12190));
  nand_5 g09842(.A(new_n12190), .B(new_n12119), .Y(new_n12191));
  nand_5 g09843(.A(new_n9165), .B(n25240), .Y(new_n12192_1));
  nand_5 g09844(.A(new_n9167), .B(new_n8297), .Y(new_n12193));
  nand_5 g09845(.A(new_n12193), .B(new_n12192_1), .Y(new_n12194));
  xnor_4 g09846(.A(new_n12194), .B(new_n12191), .Y(new_n12195));
  nand_5 g09847(.A(new_n12159), .B(new_n12148), .Y(new_n12196));
  nand_5 g09848(.A(new_n12196), .B(new_n12157_1), .Y(new_n12197));
  nand_5 g09849(.A(new_n12152_1), .B(new_n12150), .Y(new_n12198));
  nand_5 g09850(.A(new_n12198), .B(new_n12153_1), .Y(new_n12199));
  not_8  g09851(.A(new_n12199), .Y(new_n12200));
  nand_5 g09852(.A(new_n10476), .B(new_n8437), .Y(new_n12201));
  nand_5 g09853(.A(n6381), .B(n1099), .Y(new_n12202));
  nand_5 g09854(.A(new_n12202), .B(new_n12201), .Y(new_n12203));
  xor_4  g09855(.A(new_n12203), .B(new_n12200), .Y(new_n12204));
  not_8  g09856(.A(new_n12204), .Y(new_n12205));
  nand_5 g09857(.A(new_n12205), .B(n5077), .Y(new_n12206));
  not_8  g09858(.A(n5077), .Y(new_n12207));
  nand_5 g09859(.A(new_n12204), .B(new_n12207), .Y(new_n12208));
  nand_5 g09860(.A(new_n12208), .B(new_n12206), .Y(new_n12209_1));
  xor_4  g09861(.A(new_n12209_1), .B(new_n12197), .Y(new_n12210));
  or_5   g09862(.A(new_n12210), .B(new_n12195), .Y(new_n12211));
  nand_5 g09863(.A(new_n12210), .B(new_n12195), .Y(new_n12212));
  nand_5 g09864(.A(new_n12212), .B(new_n12211), .Y(new_n12213));
  xor_4  g09865(.A(new_n12213), .B(new_n12189), .Y(n1371));
  nand_5 g09866(.A(new_n10949), .B(new_n10941), .Y(new_n12215));
  nand_5 g09867(.A(new_n12215), .B(new_n10948), .Y(new_n12216));
  nand_5 g09868(.A(new_n11137), .B(new_n2412), .Y(new_n12217));
  nand_5 g09869(.A(new_n11136), .B(n3018), .Y(new_n12218));
  nand_5 g09870(.A(new_n12218), .B(new_n12217), .Y(new_n12219));
  xor_4  g09871(.A(new_n12219), .B(new_n12216), .Y(new_n12220));
  not_8  g09872(.A(new_n12220), .Y(new_n12221));
  nand_5 g09873(.A(new_n4886), .B(n11056), .Y(new_n12222));
  nand_5 g09874(.A(n20250), .B(new_n7605), .Y(new_n12223_1));
  nand_5 g09875(.A(n15271), .B(new_n4892), .Y(new_n12224));
  nand_5 g09876(.A(new_n7539), .B(n5822), .Y(new_n12225_1));
  nand_5 g09877(.A(new_n6545), .B(new_n6538), .Y(new_n12226));
  nand_5 g09878(.A(new_n12226), .B(new_n6543), .Y(new_n12227));
  nand_5 g09879(.A(new_n12227), .B(new_n12225_1), .Y(new_n12228_1));
  nand_5 g09880(.A(new_n12228_1), .B(new_n12224), .Y(new_n12229));
  nand_5 g09881(.A(new_n12229), .B(new_n12223_1), .Y(new_n12230));
  nand_5 g09882(.A(new_n12230), .B(new_n12222), .Y(new_n12231));
  nand_5 g09883(.A(n16524), .B(new_n4880), .Y(new_n12232));
  nand_5 g09884(.A(new_n8813), .B(n3785), .Y(new_n12233));
  nand_5 g09885(.A(new_n12233), .B(new_n12232), .Y(new_n12234));
  xor_4  g09886(.A(new_n12234), .B(new_n12231), .Y(new_n12235_1));
  nand_5 g09887(.A(new_n12235_1), .B(new_n12221), .Y(new_n12236));
  not_8  g09888(.A(new_n12235_1), .Y(new_n12237));
  nand_5 g09889(.A(new_n12237), .B(new_n12220), .Y(new_n12238));
  nand_5 g09890(.A(new_n12223_1), .B(new_n12222), .Y(new_n12239));
  xor_4  g09891(.A(new_n12239), .B(new_n12229), .Y(new_n12240));
  nand_5 g09892(.A(new_n12240), .B(new_n10951), .Y(new_n12241));
  not_8  g09893(.A(new_n12240), .Y(new_n12242));
  nand_5 g09894(.A(new_n12242), .B(new_n10953), .Y(new_n12243));
  nand_5 g09895(.A(new_n12225_1), .B(new_n12224), .Y(new_n12244));
  xor_4  g09896(.A(new_n12244), .B(new_n12227), .Y(new_n12245));
  nand_5 g09897(.A(new_n12245), .B(new_n10878), .Y(new_n12246));
  not_8  g09898(.A(new_n12245), .Y(new_n12247));
  nand_5 g09899(.A(new_n12247), .B(new_n10879), .Y(new_n12248));
  nand_5 g09900(.A(new_n6550), .B(new_n6533), .Y(new_n12249));
  nand_5 g09901(.A(new_n12249), .B(new_n6549), .Y(new_n12250));
  nand_5 g09902(.A(new_n12250), .B(new_n12248), .Y(new_n12251));
  nand_5 g09903(.A(new_n12251), .B(new_n12246), .Y(new_n12252));
  nand_5 g09904(.A(new_n12252), .B(new_n12243), .Y(new_n12253));
  nand_5 g09905(.A(new_n12253), .B(new_n12241), .Y(new_n12254));
  nand_5 g09906(.A(new_n12254), .B(new_n12238), .Y(new_n12255));
  nand_5 g09907(.A(new_n12255), .B(new_n12236), .Y(new_n12256));
  nand_5 g09908(.A(new_n12218), .B(new_n12216), .Y(new_n12257));
  nand_5 g09909(.A(new_n12257), .B(new_n12217), .Y(new_n12258));
  nand_5 g09910(.A(new_n11131), .B(new_n2475), .Y(new_n12259));
  nand_5 g09911(.A(new_n11130), .B(n26660), .Y(new_n12260));
  nand_5 g09912(.A(new_n12260), .B(new_n12259), .Y(new_n12261));
  xor_4  g09913(.A(new_n12261), .B(new_n12258), .Y(new_n12262));
  not_8  g09914(.A(new_n12262), .Y(new_n12263));
  nand_5 g09915(.A(new_n12233), .B(new_n12231), .Y(new_n12264));
  nand_5 g09916(.A(new_n12264), .B(new_n12232), .Y(new_n12265));
  nand_5 g09917(.A(n23160), .B(new_n4874), .Y(new_n12266));
  nand_5 g09918(.A(new_n8810), .B(n7678), .Y(new_n12267));
  nand_5 g09919(.A(new_n12267), .B(new_n12266), .Y(new_n12268));
  xor_4  g09920(.A(new_n12268), .B(new_n12265), .Y(new_n12269));
  nand_5 g09921(.A(new_n12269), .B(new_n12263), .Y(new_n12270));
  not_8  g09922(.A(new_n12269), .Y(new_n12271));
  nand_5 g09923(.A(new_n12271), .B(new_n12262), .Y(new_n12272));
  nand_5 g09924(.A(new_n12272), .B(new_n12270), .Y(new_n12273));
  xor_4  g09925(.A(new_n12273), .B(new_n12256), .Y(new_n12274));
  not_8  g09926(.A(new_n12274), .Y(new_n12275));
  nand_5 g09927(.A(new_n12275), .B(new_n6307), .Y(new_n12276));
  nand_5 g09928(.A(new_n12274), .B(new_n6308_1), .Y(new_n12277));
  nand_5 g09929(.A(new_n12236), .B(new_n12238), .Y(new_n12278));
  xor_4  g09930(.A(new_n12278), .B(new_n12254), .Y(new_n12279));
  not_8  g09931(.A(new_n12279), .Y(new_n12280));
  nand_5 g09932(.A(new_n12280), .B(new_n6315), .Y(new_n12281));
  nand_5 g09933(.A(new_n12279), .B(new_n6316), .Y(new_n12282));
  nand_5 g09934(.A(new_n12241), .B(new_n12243), .Y(new_n12283));
  xor_4  g09935(.A(new_n12283), .B(new_n12252), .Y(new_n12284));
  not_8  g09936(.A(new_n12284), .Y(new_n12285));
  nand_5 g09937(.A(new_n12285), .B(new_n6323_1), .Y(new_n12286));
  nand_5 g09938(.A(new_n12284), .B(new_n6324), .Y(new_n12287));
  nand_5 g09939(.A(new_n12246), .B(new_n12248), .Y(new_n12288));
  xor_4  g09940(.A(new_n12288), .B(new_n12250), .Y(new_n12289));
  not_8  g09941(.A(new_n12289), .Y(new_n12290));
  nand_5 g09942(.A(new_n12290), .B(new_n6330_1), .Y(new_n12291));
  nand_5 g09943(.A(new_n12289), .B(new_n6331), .Y(new_n12292));
  nand_5 g09944(.A(new_n6557), .B(new_n6552), .Y(new_n12293));
  nand_5 g09945(.A(new_n12293), .B(new_n6556_1), .Y(new_n12294));
  nand_5 g09946(.A(new_n12294), .B(new_n12292), .Y(new_n12295));
  nand_5 g09947(.A(new_n12295), .B(new_n12291), .Y(new_n12296));
  nand_5 g09948(.A(new_n12296), .B(new_n12287), .Y(new_n12297));
  nand_5 g09949(.A(new_n12297), .B(new_n12286), .Y(new_n12298));
  nand_5 g09950(.A(new_n12298), .B(new_n12282), .Y(new_n12299));
  nand_5 g09951(.A(new_n12299), .B(new_n12281), .Y(new_n12300));
  nand_5 g09952(.A(new_n12300), .B(new_n12277), .Y(new_n12301));
  nand_5 g09953(.A(new_n12301), .B(new_n12276), .Y(new_n12302_1));
  nand_5 g09954(.A(new_n12272), .B(new_n12256), .Y(new_n12303));
  nand_5 g09955(.A(new_n12303), .B(new_n12270), .Y(new_n12304_1));
  not_8  g09956(.A(new_n12304_1), .Y(new_n12305));
  nand_5 g09957(.A(new_n12260), .B(new_n12258), .Y(new_n12306));
  nand_5 g09958(.A(new_n12306), .B(new_n12259), .Y(new_n12307));
  not_8  g09959(.A(new_n12307), .Y(new_n12308));
  nand_5 g09960(.A(new_n11126), .B(new_n2568), .Y(new_n12309));
  nand_5 g09961(.A(new_n11125), .B(n13783), .Y(new_n12310));
  nand_5 g09962(.A(new_n12310), .B(new_n12309), .Y(new_n12311));
  xor_4  g09963(.A(new_n12311), .B(new_n12308), .Y(new_n12312));
  nand_5 g09964(.A(new_n12267), .B(new_n12265), .Y(new_n12313));
  nand_5 g09965(.A(new_n12313), .B(new_n12266), .Y(new_n12314));
  not_8  g09966(.A(new_n12314), .Y(new_n12315_1));
  nand_5 g09967(.A(n17250), .B(new_n4868), .Y(new_n12316));
  nand_5 g09968(.A(new_n8807), .B(n15241), .Y(new_n12317));
  nand_5 g09969(.A(new_n12317), .B(new_n12316), .Y(new_n12318));
  xor_4  g09970(.A(new_n12318), .B(new_n12315_1), .Y(new_n12319));
  not_8  g09971(.A(new_n12319), .Y(new_n12320));
  nand_5 g09972(.A(new_n12320), .B(new_n12312), .Y(new_n12321));
  not_8  g09973(.A(new_n12312), .Y(new_n12322));
  nand_5 g09974(.A(new_n12319), .B(new_n12322), .Y(new_n12323));
  nand_5 g09975(.A(new_n12323), .B(new_n12321), .Y(new_n12324_1));
  xor_4  g09976(.A(new_n12324_1), .B(new_n12305), .Y(new_n12325_1));
  nand_5 g09977(.A(new_n12325_1), .B(new_n6299), .Y(new_n12326));
  not_8  g09978(.A(new_n12325_1), .Y(new_n12327));
  nand_5 g09979(.A(new_n12327), .B(new_n6300), .Y(new_n12328));
  nand_5 g09980(.A(new_n12328), .B(new_n12326), .Y(new_n12329_1));
  xor_4  g09981(.A(new_n12329_1), .B(new_n12302_1), .Y(n1385));
  nand_5 g09982(.A(n26808), .B(n24732), .Y(new_n12331));
  nand_5 g09983(.A(new_n10458), .B(new_n4622), .Y(new_n12332));
  nand_5 g09984(.A(new_n12332), .B(new_n12331), .Y(new_n12333));
  not_8  g09985(.A(new_n12331), .Y(new_n12334));
  nand_5 g09986(.A(n7339), .B(n6631), .Y(new_n12335));
  nand_5 g09987(.A(new_n10457), .B(new_n4621), .Y(new_n12336));
  nand_5 g09988(.A(new_n12336), .B(new_n12335), .Y(new_n12337));
  xor_4  g09989(.A(new_n12337), .B(new_n12334), .Y(new_n12338));
  nand_5 g09990(.A(new_n12338), .B(new_n12333), .Y(new_n12339));
  nand_5 g09991(.A(new_n12335), .B(new_n12331), .Y(new_n12340));
  nand_5 g09992(.A(new_n12340), .B(new_n12336), .Y(new_n12341_1));
  not_8  g09993(.A(new_n12341_1), .Y(new_n12342));
  not_8  g09994(.A(n1667), .Y(new_n12343));
  nand_5 g09995(.A(new_n4620), .B(new_n12343), .Y(new_n12344));
  nand_5 g09996(.A(n14684), .B(n1667), .Y(new_n12345));
  nand_5 g09997(.A(new_n12345), .B(new_n12344), .Y(new_n12346_1));
  xor_4  g09998(.A(new_n12346_1), .B(new_n12342), .Y(new_n12347));
  not_8  g09999(.A(new_n12347), .Y(new_n12348));
  nor_5  g10000(.A(new_n12348), .B(new_n12339), .Y(new_n12349_1));
  nand_5 g10001(.A(new_n12345), .B(new_n12341_1), .Y(new_n12350));
  nand_5 g10002(.A(new_n12350), .B(new_n12344), .Y(new_n12351));
  not_8  g10003(.A(new_n12351), .Y(new_n12352));
  nand_5 g10004(.A(new_n12352), .B(n2680), .Y(new_n12353));
  not_8  g10005(.A(n2680), .Y(new_n12354));
  nand_5 g10006(.A(new_n12351), .B(new_n12354), .Y(new_n12355));
  and_5  g10007(.A(new_n12355), .B(new_n12353), .Y(new_n12356));
  xor_4  g10008(.A(new_n12356), .B(new_n4642), .Y(new_n12357));
  nand_5 g10009(.A(new_n12357), .B(new_n12349_1), .Y(new_n12358));
  nand_5 g10010(.A(new_n12353), .B(new_n4642), .Y(new_n12359));
  nand_5 g10011(.A(new_n12359), .B(new_n12355), .Y(new_n12360));
  nand_5 g10012(.A(new_n4768), .B(new_n10456), .Y(new_n12361));
  nand_5 g10013(.A(n19905), .B(n2547), .Y(new_n12362));
  nand_5 g10014(.A(new_n12362), .B(new_n12361), .Y(new_n12363));
  xor_4  g10015(.A(new_n12363), .B(new_n12360), .Y(new_n12364_1));
  nor_5  g10016(.A(new_n12364_1), .B(new_n12358), .Y(new_n12365));
  not_8  g10017(.A(n2999), .Y(new_n12366));
  nand_5 g10018(.A(new_n12136), .B(new_n12366), .Y(new_n12367));
  nand_5 g10019(.A(n26452), .B(n2999), .Y(new_n12368));
  nand_5 g10020(.A(new_n12368), .B(new_n12367), .Y(new_n12369));
  nand_5 g10021(.A(new_n12362), .B(new_n12360), .Y(new_n12370));
  nand_5 g10022(.A(new_n12370), .B(new_n12361), .Y(new_n12371));
  xor_4  g10023(.A(new_n12371), .B(new_n12369), .Y(new_n12372));
  not_8  g10024(.A(new_n12372), .Y(new_n12373));
  nand_5 g10025(.A(new_n12373), .B(new_n12365), .Y(new_n12374));
  nand_5 g10026(.A(new_n12158_1), .B(new_n10455), .Y(new_n12375));
  nand_5 g10027(.A(n15546), .B(n14702), .Y(new_n12376));
  nand_5 g10028(.A(new_n12376), .B(new_n12375), .Y(new_n12377));
  nand_5 g10029(.A(new_n12371), .B(new_n12368), .Y(new_n12378));
  nand_5 g10030(.A(new_n12378), .B(new_n12367), .Y(new_n12379));
  xor_4  g10031(.A(new_n12379), .B(new_n12377), .Y(new_n12380_1));
  nor_5  g10032(.A(new_n12380_1), .B(new_n12374), .Y(new_n12381));
  not_8  g10033(.A(n13914), .Y(new_n12382));
  nand_5 g10034(.A(new_n12382), .B(new_n12207), .Y(new_n12383_1));
  nand_5 g10035(.A(n13914), .B(n5077), .Y(new_n12384_1));
  nand_5 g10036(.A(new_n12384_1), .B(new_n12383_1), .Y(new_n12385));
  nand_5 g10037(.A(new_n12379), .B(new_n12376), .Y(new_n12386));
  nand_5 g10038(.A(new_n12386), .B(new_n12375), .Y(new_n12387));
  xor_4  g10039(.A(new_n12387), .B(new_n12385), .Y(new_n12388));
  not_8  g10040(.A(new_n12388), .Y(new_n12389));
  nand_5 g10041(.A(new_n12389), .B(new_n12381), .Y(new_n12390));
  not_8  g10042(.A(new_n12390), .Y(new_n12391));
  not_8  g10043(.A(n18035), .Y(new_n12392));
  nand_5 g10044(.A(new_n12392), .B(new_n10454), .Y(new_n12393));
  nand_5 g10045(.A(n18035), .B(n3279), .Y(new_n12394));
  nand_5 g10046(.A(new_n12394), .B(new_n12393), .Y(new_n12395));
  nand_5 g10047(.A(new_n12387), .B(new_n12384_1), .Y(new_n12396));
  nand_5 g10048(.A(new_n12396), .B(new_n12383_1), .Y(new_n12397_1));
  xor_4  g10049(.A(new_n12397_1), .B(new_n12395), .Y(new_n12398_1));
  not_8  g10050(.A(new_n12398_1), .Y(new_n12399));
  nand_5 g10051(.A(new_n12399), .B(new_n12391), .Y(new_n12400));
  nand_5 g10052(.A(n8827), .B(n4306), .Y(new_n12401));
  not_8  g10053(.A(n4306), .Y(new_n12402));
  not_8  g10054(.A(n8827), .Y(new_n12403));
  nand_5 g10055(.A(new_n12403), .B(new_n12402), .Y(new_n12404));
  nand_5 g10056(.A(new_n12404), .B(new_n12401), .Y(new_n12405));
  nand_5 g10057(.A(new_n12397_1), .B(new_n12394), .Y(new_n12406));
  nand_5 g10058(.A(new_n12406), .B(new_n12393), .Y(new_n12407));
  xor_4  g10059(.A(new_n12407), .B(new_n12405), .Y(new_n12408_1));
  or_5   g10060(.A(new_n12408_1), .B(new_n12400), .Y(new_n12409));
  nand_5 g10061(.A(new_n12408_1), .B(new_n12400), .Y(new_n12410));
  and_5  g10062(.A(new_n12410), .B(new_n12409), .Y(new_n12411));
  nand_5 g10063(.A(new_n12411), .B(new_n9153), .Y(new_n12412));
  or_5   g10064(.A(new_n12411), .B(new_n9153), .Y(new_n12413));
  nand_5 g10065(.A(new_n12413), .B(new_n12412), .Y(new_n12414));
  nand_5 g10066(.A(new_n12398_1), .B(new_n12390), .Y(new_n12415));
  and_5  g10067(.A(new_n12415), .B(new_n12400), .Y(new_n12416));
  nand_5 g10068(.A(new_n12416), .B(new_n9159), .Y(new_n12417));
  or_5   g10069(.A(new_n12416), .B(new_n9159), .Y(new_n12418));
  not_8  g10070(.A(new_n12381), .Y(new_n12419));
  nand_5 g10071(.A(new_n12388), .B(new_n12419), .Y(new_n12420));
  and_5  g10072(.A(new_n12420), .B(new_n12390), .Y(new_n12421));
  nand_5 g10073(.A(new_n12421), .B(new_n9165), .Y(new_n12422));
  or_5   g10074(.A(new_n12421), .B(new_n9165), .Y(new_n12423));
  nand_5 g10075(.A(new_n12380_1), .B(new_n12374), .Y(new_n12424));
  and_5  g10076(.A(new_n12424), .B(new_n12419), .Y(new_n12425));
  nand_5 g10077(.A(new_n12425), .B(new_n9171), .Y(new_n12426));
  or_5   g10078(.A(new_n12425), .B(new_n9171), .Y(new_n12427));
  not_8  g10079(.A(new_n12365), .Y(new_n12428));
  nand_5 g10080(.A(new_n12372), .B(new_n12428), .Y(new_n12429));
  and_5  g10081(.A(new_n12429), .B(new_n12374), .Y(new_n12430));
  nand_5 g10082(.A(new_n12430), .B(new_n9177), .Y(new_n12431));
  or_5   g10083(.A(new_n12430), .B(new_n9177), .Y(new_n12432));
  nand_5 g10084(.A(new_n12364_1), .B(new_n12358), .Y(new_n12433));
  and_5  g10085(.A(new_n12433), .B(new_n12428), .Y(new_n12434));
  nand_5 g10086(.A(new_n12434), .B(new_n9184), .Y(new_n12435));
  or_5   g10087(.A(new_n12434), .B(new_n9184), .Y(new_n12436));
  not_8  g10088(.A(new_n12357), .Y(new_n12437));
  xor_4  g10089(.A(new_n12437), .B(new_n12349_1), .Y(new_n12438));
  or_5   g10090(.A(new_n12438), .B(new_n9189), .Y(new_n12439));
  nand_5 g10091(.A(new_n12438), .B(new_n9189), .Y(new_n12440));
  xor_4  g10092(.A(new_n12347), .B(new_n12339), .Y(new_n12441));
  or_5   g10093(.A(new_n12441), .B(new_n9197), .Y(new_n12442));
  nand_5 g10094(.A(new_n12441), .B(new_n9197), .Y(new_n12443));
  not_8  g10095(.A(new_n12333), .Y(new_n12444));
  nand_5 g10096(.A(new_n12444), .B(new_n2616), .Y(new_n12445));
  or_5   g10097(.A(new_n12445), .B(new_n9202), .Y(new_n12446_1));
  nand_5 g10098(.A(new_n12445), .B(new_n9204), .Y(new_n12447));
  xor_4  g10099(.A(new_n12338), .B(new_n12444), .Y(new_n12448));
  not_8  g10100(.A(new_n12448), .Y(new_n12449_1));
  nand_5 g10101(.A(new_n12449_1), .B(new_n12447), .Y(new_n12450));
  nand_5 g10102(.A(new_n12450), .B(new_n12446_1), .Y(new_n12451));
  nand_5 g10103(.A(new_n12451), .B(new_n12443), .Y(new_n12452));
  nand_5 g10104(.A(new_n12452), .B(new_n12442), .Y(new_n12453));
  nand_5 g10105(.A(new_n12453), .B(new_n12440), .Y(new_n12454));
  nand_5 g10106(.A(new_n12454), .B(new_n12439), .Y(new_n12455));
  nand_5 g10107(.A(new_n12455), .B(new_n12436), .Y(new_n12456));
  nand_5 g10108(.A(new_n12456), .B(new_n12435), .Y(new_n12457));
  nand_5 g10109(.A(new_n12457), .B(new_n12432), .Y(new_n12458));
  nand_5 g10110(.A(new_n12458), .B(new_n12431), .Y(new_n12459));
  nand_5 g10111(.A(new_n12459), .B(new_n12427), .Y(new_n12460));
  nand_5 g10112(.A(new_n12460), .B(new_n12426), .Y(new_n12461_1));
  nand_5 g10113(.A(new_n12461_1), .B(new_n12423), .Y(new_n12462_1));
  nand_5 g10114(.A(new_n12462_1), .B(new_n12422), .Y(new_n12463));
  nand_5 g10115(.A(new_n12463), .B(new_n12418), .Y(new_n12464));
  nand_5 g10116(.A(new_n12464), .B(new_n12417), .Y(new_n12465));
  xor_4  g10117(.A(new_n12465), .B(new_n12414), .Y(new_n12466));
  nand_5 g10118(.A(new_n12466), .B(new_n10511), .Y(new_n12467_1));
  or_5   g10119(.A(new_n12466), .B(new_n10511), .Y(new_n12468));
  nand_5 g10120(.A(new_n12468), .B(new_n12467_1), .Y(new_n12469_1));
  nand_5 g10121(.A(new_n12418), .B(new_n12417), .Y(new_n12470));
  xor_4  g10122(.A(new_n12470), .B(new_n12463), .Y(new_n12471));
  nand_5 g10123(.A(new_n12471), .B(new_n10518), .Y(new_n12472));
  or_5   g10124(.A(new_n12471), .B(new_n10518), .Y(new_n12473));
  nand_5 g10125(.A(new_n12423), .B(new_n12422), .Y(new_n12474));
  xor_4  g10126(.A(new_n12474), .B(new_n12461_1), .Y(new_n12475));
  nand_5 g10127(.A(new_n12475), .B(new_n10524), .Y(new_n12476));
  or_5   g10128(.A(new_n12475), .B(new_n10524), .Y(new_n12477));
  nand_5 g10129(.A(new_n12427), .B(new_n12426), .Y(new_n12478));
  xor_4  g10130(.A(new_n12478), .B(new_n12459), .Y(new_n12479));
  nand_5 g10131(.A(new_n12479), .B(new_n10530), .Y(new_n12480));
  or_5   g10132(.A(new_n12479), .B(new_n10530), .Y(new_n12481));
  nand_5 g10133(.A(new_n12432), .B(new_n12431), .Y(new_n12482));
  xor_4  g10134(.A(new_n12482), .B(new_n12457), .Y(new_n12483));
  nand_5 g10135(.A(new_n12483), .B(new_n10536), .Y(new_n12484));
  or_5   g10136(.A(new_n12483), .B(new_n10536), .Y(new_n12485));
  nand_5 g10137(.A(new_n12436), .B(new_n12435), .Y(new_n12486));
  xor_4  g10138(.A(new_n12486), .B(new_n12455), .Y(new_n12487));
  nand_5 g10139(.A(new_n12487), .B(new_n10542), .Y(new_n12488));
  or_5   g10140(.A(new_n12487), .B(new_n10542), .Y(new_n12489));
  nand_5 g10141(.A(new_n12440), .B(new_n12439), .Y(new_n12490));
  xor_4  g10142(.A(new_n12490), .B(new_n12453), .Y(new_n12491));
  nand_5 g10143(.A(new_n12491), .B(new_n10548), .Y(new_n12492));
  or_5   g10144(.A(new_n12491), .B(new_n10548), .Y(new_n12493));
  nand_5 g10145(.A(new_n12443), .B(new_n12442), .Y(new_n12494));
  xor_4  g10146(.A(new_n12494), .B(new_n12451), .Y(new_n12495_1));
  nand_5 g10147(.A(new_n12495_1), .B(new_n10555), .Y(new_n12496));
  nor_5  g10148(.A(new_n12495_1), .B(new_n10555), .Y(new_n12497));
  not_8  g10149(.A(new_n12497), .Y(new_n12498));
  not_8  g10150(.A(new_n10561_1), .Y(new_n12499));
  nand_5 g10151(.A(new_n12333), .B(new_n9714), .Y(new_n12500));
  and_5  g10152(.A(new_n12500), .B(new_n12445), .Y(new_n12501));
  or_5   g10153(.A(new_n12501), .B(new_n10565), .Y(new_n12502));
  or_5   g10154(.A(new_n12502), .B(new_n12499), .Y(new_n12503));
  nand_5 g10155(.A(new_n12502), .B(new_n12499), .Y(new_n12504));
  nand_5 g10156(.A(new_n12447), .B(new_n12446_1), .Y(new_n12505));
  xor_4  g10157(.A(new_n12505), .B(new_n12448), .Y(new_n12506));
  not_8  g10158(.A(new_n12506), .Y(new_n12507_1));
  nand_5 g10159(.A(new_n12507_1), .B(new_n12504), .Y(new_n12508));
  nand_5 g10160(.A(new_n12508), .B(new_n12503), .Y(new_n12509));
  nand_5 g10161(.A(new_n12509), .B(new_n12498), .Y(new_n12510));
  nand_5 g10162(.A(new_n12510), .B(new_n12496), .Y(new_n12511));
  nand_5 g10163(.A(new_n12511), .B(new_n12493), .Y(new_n12512));
  nand_5 g10164(.A(new_n12512), .B(new_n12492), .Y(new_n12513));
  nand_5 g10165(.A(new_n12513), .B(new_n12489), .Y(new_n12514));
  nand_5 g10166(.A(new_n12514), .B(new_n12488), .Y(new_n12515_1));
  nand_5 g10167(.A(new_n12515_1), .B(new_n12485), .Y(new_n12516_1));
  nand_5 g10168(.A(new_n12516_1), .B(new_n12484), .Y(new_n12517));
  nand_5 g10169(.A(new_n12517), .B(new_n12481), .Y(new_n12518));
  nand_5 g10170(.A(new_n12518), .B(new_n12480), .Y(new_n12519));
  nand_5 g10171(.A(new_n12519), .B(new_n12477), .Y(new_n12520));
  nand_5 g10172(.A(new_n12520), .B(new_n12476), .Y(new_n12521));
  nand_5 g10173(.A(new_n12521), .B(new_n12473), .Y(new_n12522));
  nand_5 g10174(.A(new_n12522), .B(new_n12472), .Y(new_n12523));
  xor_4  g10175(.A(new_n12523), .B(new_n12469_1), .Y(n1498));
  nand_5 g10176(.A(n20658), .B(n9090), .Y(new_n12525));
  not_8  g10177(.A(n9090), .Y(new_n12526));
  nand_5 g10178(.A(new_n5469), .B(new_n12526), .Y(new_n12527));
  and_5  g10179(.A(new_n12527), .B(new_n12525), .Y(new_n12528));
  nand_5 g10180(.A(new_n12528), .B(new_n6767), .Y(new_n12529));
  not_8  g10181(.A(new_n12529), .Y(new_n12530));
  nor_5  g10182(.A(new_n12528), .B(new_n6767), .Y(new_n12531));
  nor_5  g10183(.A(new_n12531), .B(new_n12530), .Y(new_n12532));
  nand_5 g10184(.A(new_n12532), .B(new_n5633), .Y(new_n12533));
  not_8  g10185(.A(new_n12533), .Y(new_n12534));
  nor_5  g10186(.A(new_n12532), .B(new_n5633), .Y(new_n12535));
  nor_5  g10187(.A(new_n12535), .B(new_n12534), .Y(n1501));
  nand_5 g10188(.A(new_n11065), .B(new_n11061), .Y(new_n12537));
  nand_5 g10189(.A(new_n12537), .B(new_n11064), .Y(new_n12538));
  not_8  g10190(.A(n21222), .Y(new_n12539));
  not_8  g10191(.A(n26565), .Y(new_n12540_1));
  nand_5 g10192(.A(new_n12540_1), .B(new_n12539), .Y(new_n12541));
  nand_5 g10193(.A(n26565), .B(n21222), .Y(new_n12542));
  nand_5 g10194(.A(new_n12542), .B(new_n12541), .Y(new_n12543));
  xor_4  g10195(.A(new_n12543), .B(new_n12538), .Y(new_n12544));
  not_8  g10196(.A(n25094), .Y(new_n12545_1));
  not_8  g10197(.A(n11473), .Y(new_n12546_1));
  not_8  g10198(.A(n15506), .Y(new_n12547));
  nand_5 g10199(.A(new_n12547), .B(new_n12546_1), .Y(new_n12548));
  or_5   g10200(.A(new_n12548), .B(n5131), .Y(new_n12549));
  nor_5  g10201(.A(new_n12549), .B(n21538), .Y(new_n12550));
  nand_5 g10202(.A(new_n12550), .B(new_n12545_1), .Y(new_n12551));
  not_8  g10203(.A(new_n12551), .Y(new_n12552_1));
  nor_5  g10204(.A(new_n12550), .B(new_n12545_1), .Y(new_n12553));
  nor_5  g10205(.A(new_n12553), .B(new_n12552_1), .Y(new_n12554));
  nand_5 g10206(.A(new_n12554), .B(new_n11184_1), .Y(new_n12555));
  not_8  g10207(.A(new_n11184_1), .Y(new_n12556));
  not_8  g10208(.A(new_n12554), .Y(new_n12557));
  nand_5 g10209(.A(new_n12557), .B(new_n12556), .Y(new_n12558));
  not_8  g10210(.A(n21538), .Y(new_n12559));
  xor_4  g10211(.A(new_n12549), .B(new_n12559), .Y(new_n12560));
  not_8  g10212(.A(new_n12560), .Y(new_n12561));
  nand_5 g10213(.A(new_n12561), .B(new_n11192_1), .Y(new_n12562_1));
  or_5   g10214(.A(new_n12561), .B(new_n11192_1), .Y(new_n12563));
  nand_5 g10215(.A(new_n12548), .B(n5131), .Y(new_n12564));
  and_5  g10216(.A(new_n12564), .B(new_n12549), .Y(new_n12565));
  nand_5 g10217(.A(new_n12565), .B(new_n11196), .Y(new_n12566_1));
  not_8  g10218(.A(new_n11196), .Y(new_n12567));
  not_8  g10219(.A(new_n12565), .Y(new_n12568));
  nand_5 g10220(.A(new_n12568), .B(new_n12567), .Y(new_n12569_1));
  nand_5 g10221(.A(new_n11208), .B(n15506), .Y(new_n12570));
  or_5   g10222(.A(new_n12570), .B(n11473), .Y(new_n12571));
  nand_5 g10223(.A(n15506), .B(n11473), .Y(new_n12572));
  and_5  g10224(.A(new_n12572), .B(new_n12548), .Y(new_n12573));
  not_8  g10225(.A(new_n12573), .Y(new_n12574));
  nand_5 g10226(.A(new_n12574), .B(new_n12570), .Y(new_n12575));
  nand_5 g10227(.A(new_n12575), .B(new_n11204), .Y(new_n12576));
  nand_5 g10228(.A(new_n12576), .B(new_n12571), .Y(new_n12577));
  nand_5 g10229(.A(new_n12577), .B(new_n12569_1), .Y(new_n12578));
  nand_5 g10230(.A(new_n12578), .B(new_n12566_1), .Y(new_n12579));
  nand_5 g10231(.A(new_n12579), .B(new_n12563), .Y(new_n12580));
  nand_5 g10232(.A(new_n12580), .B(new_n12562_1), .Y(new_n12581));
  nand_5 g10233(.A(new_n12581), .B(new_n12558), .Y(new_n12582));
  nand_5 g10234(.A(new_n12582), .B(new_n12555), .Y(new_n12583));
  not_8  g10235(.A(n1611), .Y(new_n12584));
  nand_5 g10236(.A(new_n12552_1), .B(new_n12584), .Y(new_n12585));
  nand_5 g10237(.A(new_n12551), .B(n1611), .Y(new_n12586));
  and_5  g10238(.A(new_n12586), .B(new_n12585), .Y(new_n12587_1));
  nand_5 g10239(.A(new_n12587_1), .B(new_n11178), .Y(new_n12588));
  not_8  g10240(.A(new_n11178), .Y(new_n12589));
  not_8  g10241(.A(new_n12587_1), .Y(new_n12590));
  nand_5 g10242(.A(new_n12590), .B(new_n12589), .Y(new_n12591));
  nand_5 g10243(.A(new_n12591), .B(new_n12588), .Y(new_n12592));
  xor_4  g10244(.A(new_n12592), .B(new_n12583), .Y(new_n12593_1));
  or_5   g10245(.A(new_n12593_1), .B(new_n12544), .Y(new_n12594));
  nand_5 g10246(.A(new_n12593_1), .B(new_n12544), .Y(new_n12595));
  nand_5 g10247(.A(new_n12555), .B(new_n12558), .Y(new_n12596));
  xor_4  g10248(.A(new_n12596), .B(new_n12581), .Y(new_n12597));
  or_5   g10249(.A(new_n12597), .B(new_n11068), .Y(new_n12598));
  nand_5 g10250(.A(new_n12597), .B(new_n11068), .Y(new_n12599));
  nand_5 g10251(.A(new_n12562_1), .B(new_n12563), .Y(new_n12600));
  xor_4  g10252(.A(new_n12600), .B(new_n12579), .Y(new_n12601));
  or_5   g10253(.A(new_n12601), .B(new_n10987), .Y(new_n12602));
  nand_5 g10254(.A(new_n12601), .B(new_n10987), .Y(new_n12603));
  nand_5 g10255(.A(new_n12566_1), .B(new_n12569_1), .Y(new_n12604));
  xor_4  g10256(.A(new_n12604), .B(new_n12577), .Y(new_n12605));
  nand_5 g10257(.A(new_n12605), .B(new_n11039), .Y(new_n12606));
  or_5   g10258(.A(new_n12605), .B(new_n11039), .Y(new_n12607_1));
  not_8  g10259(.A(new_n11048), .Y(new_n12608));
  not_8  g10260(.A(new_n11208), .Y(new_n12609));
  nand_5 g10261(.A(new_n12609), .B(new_n12547), .Y(new_n12610));
  and_5  g10262(.A(new_n12610), .B(new_n12570), .Y(new_n12611));
  not_8  g10263(.A(new_n12611), .Y(new_n12612));
  nand_5 g10264(.A(new_n12612), .B(new_n8278), .Y(new_n12613));
  or_5   g10265(.A(new_n12613), .B(new_n12608), .Y(new_n12614));
  nand_5 g10266(.A(new_n12613), .B(new_n12608), .Y(new_n12615));
  nand_5 g10267(.A(new_n12575), .B(new_n12571), .Y(new_n12616));
  xor_4  g10268(.A(new_n12616), .B(new_n11204), .Y(new_n12617));
  nand_5 g10269(.A(new_n12617), .B(new_n12615), .Y(new_n12618));
  nand_5 g10270(.A(new_n12618), .B(new_n12614), .Y(new_n12619));
  nand_5 g10271(.A(new_n12619), .B(new_n12607_1), .Y(new_n12620_1));
  and_5  g10272(.A(new_n12620_1), .B(new_n12606), .Y(new_n12621_1));
  nand_5 g10273(.A(new_n12621_1), .B(new_n12603), .Y(new_n12622));
  nand_5 g10274(.A(new_n12622), .B(new_n12602), .Y(new_n12623));
  nand_5 g10275(.A(new_n12623), .B(new_n12599), .Y(new_n12624));
  nand_5 g10276(.A(new_n12624), .B(new_n12598), .Y(new_n12625));
  nand_5 g10277(.A(new_n12625), .B(new_n12595), .Y(new_n12626_1));
  nand_5 g10278(.A(new_n12626_1), .B(new_n12594), .Y(new_n12627));
  nand_5 g10279(.A(new_n12542), .B(new_n12538), .Y(new_n12628));
  nand_5 g10280(.A(new_n12628), .B(new_n12541), .Y(new_n12629));
  not_8  g10281(.A(new_n12629), .Y(new_n12630));
  not_8  g10282(.A(n3366), .Y(new_n12631));
  not_8  g10283(.A(n20470), .Y(new_n12632));
  nand_5 g10284(.A(new_n12632), .B(new_n12631), .Y(new_n12633));
  nand_5 g10285(.A(n20470), .B(n3366), .Y(new_n12634));
  nand_5 g10286(.A(new_n12634), .B(new_n12633), .Y(new_n12635));
  xor_4  g10287(.A(new_n12635), .B(new_n12630), .Y(new_n12636));
  nand_5 g10288(.A(new_n12591), .B(new_n12583), .Y(new_n12637));
  nand_5 g10289(.A(new_n12637), .B(new_n12588), .Y(new_n12638));
  or_5   g10290(.A(new_n12585), .B(n752), .Y(new_n12639));
  nand_5 g10291(.A(new_n12585), .B(n752), .Y(new_n12640));
  and_5  g10292(.A(new_n12640), .B(new_n12639), .Y(new_n12641));
  nand_5 g10293(.A(new_n12641), .B(new_n11172), .Y(new_n12642));
  not_8  g10294(.A(new_n11172), .Y(new_n12643));
  not_8  g10295(.A(new_n12641), .Y(new_n12644));
  nand_5 g10296(.A(new_n12644), .B(new_n12643), .Y(new_n12645));
  nand_5 g10297(.A(new_n12645), .B(new_n12642), .Y(new_n12646));
  xnor_4 g10298(.A(new_n12646), .B(new_n12638), .Y(new_n12647));
  nand_5 g10299(.A(new_n12647), .B(new_n12636), .Y(new_n12648));
  not_8  g10300(.A(new_n12648), .Y(new_n12649));
  nor_5  g10301(.A(new_n12647), .B(new_n12636), .Y(new_n12650_1));
  nor_5  g10302(.A(new_n12650_1), .B(new_n12649), .Y(new_n12651));
  xor_4  g10303(.A(new_n12651), .B(new_n12627), .Y(n1518));
  nand_5 g10304(.A(new_n10076), .B(new_n10038), .Y(new_n12653));
  nand_5 g10305(.A(new_n12653), .B(new_n10039), .Y(new_n12654_1));
  nand_5 g10306(.A(n17458), .B(new_n9104_1), .Y(new_n12655));
  nand_5 g10307(.A(new_n8291), .B(n14826), .Y(new_n12656));
  nand_5 g10308(.A(new_n9107), .B(n1222), .Y(new_n12657_1));
  nand_5 g10309(.A(n23493), .B(new_n8294), .Y(new_n12658));
  nand_5 g10310(.A(n25240), .B(new_n9110), .Y(new_n12659));
  nand_5 g10311(.A(new_n8297), .B(n10275), .Y(new_n12660));
  nand_5 g10312(.A(new_n9113), .B(n10125), .Y(new_n12661));
  nand_5 g10313(.A(n15146), .B(new_n8300), .Y(new_n12662));
  nand_5 g10314(.A(new_n9116), .B(n8067), .Y(new_n12663));
  nand_5 g10315(.A(n11579), .B(new_n8303), .Y(new_n12664));
  nand_5 g10316(.A(n20923), .B(new_n9120), .Y(new_n12665_1));
  nand_5 g10317(.A(new_n8306_1), .B(n21), .Y(new_n12666));
  nand_5 g10318(.A(n18157), .B(new_n9122), .Y(new_n12667));
  nand_5 g10319(.A(new_n7606), .B(n1682), .Y(new_n12668));
  nand_5 g10320(.A(n12161), .B(new_n9123), .Y(new_n12669));
  nand_5 g10321(.A(new_n7538), .B(n7963), .Y(new_n12670_1));
  nand_5 g10322(.A(new_n9126), .B(n5026), .Y(new_n12671));
  nand_5 g10323(.A(n10017), .B(new_n7519), .Y(new_n12672));
  nand_5 g10324(.A(new_n7526), .B(n3618), .Y(new_n12673));
  nand_5 g10325(.A(new_n12673), .B(new_n12672), .Y(new_n12674));
  nand_5 g10326(.A(new_n12674), .B(new_n12671), .Y(new_n12675));
  nand_5 g10327(.A(new_n12675), .B(new_n12670_1), .Y(new_n12676));
  nand_5 g10328(.A(new_n12676), .B(new_n12669), .Y(new_n12677));
  nand_5 g10329(.A(new_n12677), .B(new_n12668), .Y(new_n12678));
  nand_5 g10330(.A(new_n12678), .B(new_n12667), .Y(new_n12679));
  nand_5 g10331(.A(new_n12679), .B(new_n12666), .Y(new_n12680));
  nand_5 g10332(.A(new_n12680), .B(new_n12665_1), .Y(new_n12681));
  nand_5 g10333(.A(new_n12681), .B(new_n12664), .Y(new_n12682));
  nand_5 g10334(.A(new_n12682), .B(new_n12663), .Y(new_n12683));
  nand_5 g10335(.A(new_n12683), .B(new_n12662), .Y(new_n12684));
  nand_5 g10336(.A(new_n12684), .B(new_n12661), .Y(new_n12685));
  nand_5 g10337(.A(new_n12685), .B(new_n12660), .Y(new_n12686));
  nand_5 g10338(.A(new_n12686), .B(new_n12659), .Y(new_n12687));
  nand_5 g10339(.A(new_n12687), .B(new_n12658), .Y(new_n12688));
  nand_5 g10340(.A(new_n12688), .B(new_n12657_1), .Y(new_n12689));
  nand_5 g10341(.A(new_n12689), .B(new_n12656), .Y(new_n12690));
  nand_5 g10342(.A(new_n12690), .B(new_n12655), .Y(new_n12691));
  nor_5  g10343(.A(new_n4793), .B(n12821), .Y(new_n12692));
  nand_5 g10344(.A(new_n12692), .B(new_n2798), .Y(new_n12693));
  nor_5  g10345(.A(new_n12693), .B(n7330), .Y(new_n12694));
  nand_5 g10346(.A(new_n12694), .B(new_n2785), .Y(new_n12695));
  nand_5 g10347(.A(new_n12695), .B(n2944), .Y(new_n12696));
  nor_5  g10348(.A(new_n12695), .B(n2944), .Y(new_n12697));
  not_8  g10349(.A(new_n12697), .Y(new_n12698));
  and_5  g10350(.A(new_n12698), .B(new_n12696), .Y(new_n12699));
  not_8  g10351(.A(new_n12699), .Y(new_n12700));
  nand_5 g10352(.A(new_n12700), .B(new_n8335), .Y(new_n12701));
  not_8  g10353(.A(new_n12701), .Y(new_n12702_1));
  xor_4  g10354(.A(new_n12694), .B(new_n2785), .Y(new_n12703));
  not_8  g10355(.A(new_n12703), .Y(new_n12704));
  nand_5 g10356(.A(new_n12704), .B(new_n3295), .Y(new_n12705));
  nand_5 g10357(.A(new_n12703), .B(n12657), .Y(new_n12706));
  xor_4  g10358(.A(new_n12693), .B(n7330), .Y(new_n12707_1));
  not_8  g10359(.A(new_n12707_1), .Y(new_n12708));
  nand_5 g10360(.A(new_n12708), .B(new_n3195), .Y(new_n12709));
  nand_5 g10361(.A(new_n12707_1), .B(n17077), .Y(new_n12710));
  xor_4  g10362(.A(new_n12692), .B(new_n2798), .Y(new_n12711));
  not_8  g10363(.A(new_n12711), .Y(new_n12712));
  nand_5 g10364(.A(new_n12712), .B(new_n3109), .Y(new_n12713));
  nand_5 g10365(.A(new_n12711), .B(n26510), .Y(new_n12714));
  xor_4  g10366(.A(new_n4793), .B(n12821), .Y(new_n12715));
  not_8  g10367(.A(new_n12715), .Y(new_n12716));
  nand_5 g10368(.A(new_n12716), .B(new_n3073), .Y(new_n12717));
  nand_5 g10369(.A(new_n12715), .B(n23068), .Y(new_n12718));
  nand_5 g10370(.A(new_n4798), .B(new_n4791), .Y(new_n12719));
  nand_5 g10371(.A(new_n12719), .B(new_n4797), .Y(new_n12720));
  nand_5 g10372(.A(new_n12720), .B(new_n12718), .Y(new_n12721));
  nand_5 g10373(.A(new_n12721), .B(new_n12717), .Y(new_n12722));
  nand_5 g10374(.A(new_n12722), .B(new_n12714), .Y(new_n12723));
  nand_5 g10375(.A(new_n12723), .B(new_n12713), .Y(new_n12724));
  nand_5 g10376(.A(new_n12724), .B(new_n12710), .Y(new_n12725_1));
  nand_5 g10377(.A(new_n12725_1), .B(new_n12709), .Y(new_n12726));
  nand_5 g10378(.A(new_n12726), .B(new_n12706), .Y(new_n12727_1));
  nand_5 g10379(.A(new_n12727_1), .B(new_n12705), .Y(new_n12728));
  nor_5  g10380(.A(new_n12728), .B(new_n12702_1), .Y(new_n12729));
  nand_5 g10381(.A(new_n12699), .B(n19282), .Y(new_n12730));
  nand_5 g10382(.A(new_n12730), .B(new_n12698), .Y(new_n12731));
  nor_5  g10383(.A(new_n12731), .B(new_n12729), .Y(new_n12732));
  not_8  g10384(.A(new_n12732), .Y(new_n12733));
  nand_5 g10385(.A(new_n12733), .B(new_n12691), .Y(new_n12734));
  not_8  g10386(.A(new_n12734), .Y(new_n12735));
  not_8  g10387(.A(new_n12691), .Y(new_n12736));
  nand_5 g10388(.A(new_n12732), .B(new_n12736), .Y(new_n12737));
  nand_5 g10389(.A(new_n12737), .B(new_n12734), .Y(new_n12738));
  nand_5 g10390(.A(new_n12656), .B(new_n12655), .Y(new_n12739));
  xor_4  g10391(.A(new_n12739), .B(new_n12689), .Y(new_n12740_1));
  nand_5 g10392(.A(new_n12730), .B(new_n12701), .Y(new_n12741));
  xor_4  g10393(.A(new_n12741), .B(new_n12728), .Y(new_n12742_1));
  not_8  g10394(.A(new_n12742_1), .Y(new_n12743));
  nand_5 g10395(.A(new_n12743), .B(new_n12740_1), .Y(new_n12744));
  not_8  g10396(.A(new_n12740_1), .Y(new_n12745));
  nand_5 g10397(.A(new_n12742_1), .B(new_n12745), .Y(new_n12746_1));
  nand_5 g10398(.A(new_n12658), .B(new_n12657_1), .Y(new_n12747));
  xor_4  g10399(.A(new_n12747), .B(new_n12687), .Y(new_n12748));
  nand_5 g10400(.A(new_n12706), .B(new_n12705), .Y(new_n12749));
  xor_4  g10401(.A(new_n12749), .B(new_n12726), .Y(new_n12750));
  not_8  g10402(.A(new_n12750), .Y(new_n12751));
  nand_5 g10403(.A(new_n12751), .B(new_n12748), .Y(new_n12752));
  or_5   g10404(.A(new_n12751), .B(new_n12748), .Y(new_n12753));
  nand_5 g10405(.A(new_n12660), .B(new_n12659), .Y(new_n12754));
  xor_4  g10406(.A(new_n12754), .B(new_n12685), .Y(new_n12755));
  nand_5 g10407(.A(new_n12710), .B(new_n12709), .Y(new_n12756_1));
  xor_4  g10408(.A(new_n12756_1), .B(new_n12724), .Y(new_n12757));
  not_8  g10409(.A(new_n12757), .Y(new_n12758));
  nand_5 g10410(.A(new_n12758), .B(new_n12755), .Y(new_n12759));
  or_5   g10411(.A(new_n12758), .B(new_n12755), .Y(new_n12760));
  nand_5 g10412(.A(new_n12662), .B(new_n12661), .Y(new_n12761));
  xor_4  g10413(.A(new_n12761), .B(new_n12683), .Y(new_n12762));
  nand_5 g10414(.A(new_n12714), .B(new_n12713), .Y(new_n12763));
  xor_4  g10415(.A(new_n12763), .B(new_n12722), .Y(new_n12764));
  not_8  g10416(.A(new_n12764), .Y(new_n12765));
  nand_5 g10417(.A(new_n12765), .B(new_n12762), .Y(new_n12766));
  or_5   g10418(.A(new_n12765), .B(new_n12762), .Y(new_n12767));
  nand_5 g10419(.A(new_n12664), .B(new_n12663), .Y(new_n12768));
  xor_4  g10420(.A(new_n12768), .B(new_n12681), .Y(new_n12769));
  nand_5 g10421(.A(new_n12718), .B(new_n12717), .Y(new_n12770));
  xor_4  g10422(.A(new_n12770), .B(new_n12720), .Y(new_n12771));
  not_8  g10423(.A(new_n12771), .Y(new_n12772));
  nand_5 g10424(.A(new_n12772), .B(new_n12769), .Y(new_n12773));
  or_5   g10425(.A(new_n12772), .B(new_n12769), .Y(new_n12774));
  nand_5 g10426(.A(new_n12666), .B(new_n12665_1), .Y(new_n12775));
  xor_4  g10427(.A(new_n12775), .B(new_n12679), .Y(new_n12776));
  nand_5 g10428(.A(new_n12776), .B(new_n4800), .Y(new_n12777));
  not_8  g10429(.A(new_n12776), .Y(new_n12778));
  nand_5 g10430(.A(new_n12778), .B(new_n4802), .Y(new_n12779));
  nand_5 g10431(.A(new_n12668), .B(new_n12667), .Y(new_n12780));
  xor_4  g10432(.A(new_n12780), .B(new_n12677), .Y(new_n12781));
  nand_5 g10433(.A(new_n12781), .B(new_n4729), .Y(new_n12782));
  or_5   g10434(.A(new_n12781), .B(new_n4729), .Y(new_n12783_1));
  nand_5 g10435(.A(new_n12670_1), .B(new_n12669), .Y(new_n12784));
  xor_4  g10436(.A(new_n12784), .B(new_n12675), .Y(new_n12785));
  nand_5 g10437(.A(new_n12785), .B(new_n4687), .Y(new_n12786));
  not_8  g10438(.A(new_n12785), .Y(new_n12787));
  nand_5 g10439(.A(new_n12787), .B(new_n4688), .Y(new_n12788));
  nand_5 g10440(.A(new_n12672), .B(new_n12671), .Y(new_n12789));
  xnor_4 g10441(.A(new_n12789), .B(new_n12673), .Y(new_n12790));
  not_8  g10442(.A(new_n12790), .Y(new_n12791));
  nand_5 g10443(.A(n8581), .B(new_n2614), .Y(new_n12792));
  and_5  g10444(.A(new_n12792), .B(new_n12673), .Y(new_n12793));
  not_8  g10445(.A(new_n12793), .Y(new_n12794));
  nand_5 g10446(.A(new_n12794), .B(new_n4701), .Y(new_n12795));
  nand_5 g10447(.A(new_n12795), .B(new_n12791), .Y(new_n12796));
  or_5   g10448(.A(new_n12795), .B(new_n12791), .Y(new_n12797));
  nand_5 g10449(.A(new_n12797), .B(new_n4694), .Y(new_n12798));
  nand_5 g10450(.A(new_n12798), .B(new_n12796), .Y(new_n12799));
  nand_5 g10451(.A(new_n12799), .B(new_n12788), .Y(new_n12800));
  nand_5 g10452(.A(new_n12800), .B(new_n12786), .Y(new_n12801_1));
  nand_5 g10453(.A(new_n12801_1), .B(new_n12783_1), .Y(new_n12802));
  nand_5 g10454(.A(new_n12802), .B(new_n12782), .Y(new_n12803));
  nand_5 g10455(.A(new_n12803), .B(new_n12779), .Y(new_n12804));
  nand_5 g10456(.A(new_n12804), .B(new_n12777), .Y(new_n12805));
  nand_5 g10457(.A(new_n12805), .B(new_n12774), .Y(new_n12806));
  nand_5 g10458(.A(new_n12806), .B(new_n12773), .Y(new_n12807));
  nand_5 g10459(.A(new_n12807), .B(new_n12767), .Y(new_n12808));
  nand_5 g10460(.A(new_n12808), .B(new_n12766), .Y(new_n12809));
  nand_5 g10461(.A(new_n12809), .B(new_n12760), .Y(new_n12810));
  nand_5 g10462(.A(new_n12810), .B(new_n12759), .Y(new_n12811_1));
  nand_5 g10463(.A(new_n12811_1), .B(new_n12753), .Y(new_n12812_1));
  nand_5 g10464(.A(new_n12812_1), .B(new_n12752), .Y(new_n12813));
  nand_5 g10465(.A(new_n12813), .B(new_n12746_1), .Y(new_n12814));
  nand_5 g10466(.A(new_n12814), .B(new_n12744), .Y(new_n12815));
  nor_5  g10467(.A(new_n12815), .B(new_n12738), .Y(new_n12816_1));
  nor_5  g10468(.A(new_n12816_1), .B(new_n12735), .Y(new_n12817));
  xor_4  g10469(.A(new_n12817), .B(new_n12654_1), .Y(new_n12818));
  xor_4  g10470(.A(new_n12815), .B(new_n12738), .Y(new_n12819));
  not_8  g10471(.A(new_n12819), .Y(new_n12820));
  nand_5 g10472(.A(new_n12820), .B(new_n12654_1), .Y(new_n12821_1));
  not_8  g10473(.A(new_n12654_1), .Y(new_n12822));
  nand_5 g10474(.A(new_n12819), .B(new_n12822), .Y(new_n12823));
  nand_5 g10475(.A(new_n12744), .B(new_n12746_1), .Y(new_n12824));
  xor_4  g10476(.A(new_n12824), .B(new_n12813), .Y(new_n12825));
  not_8  g10477(.A(new_n12825), .Y(new_n12826));
  nand_5 g10478(.A(new_n12826), .B(new_n10079), .Y(new_n12827));
  nand_5 g10479(.A(new_n12825), .B(new_n10078), .Y(new_n12828));
  nand_5 g10480(.A(new_n12752), .B(new_n12753), .Y(new_n12829));
  xor_4  g10481(.A(new_n12829), .B(new_n12811_1), .Y(new_n12830));
  not_8  g10482(.A(new_n12830), .Y(new_n12831));
  nand_5 g10483(.A(new_n12831), .B(new_n10086), .Y(new_n12832));
  nand_5 g10484(.A(new_n12830), .B(new_n10087), .Y(new_n12833));
  nand_5 g10485(.A(new_n12759), .B(new_n12760), .Y(new_n12834));
  xor_4  g10486(.A(new_n12834), .B(new_n12809), .Y(new_n12835));
  not_8  g10487(.A(new_n12835), .Y(new_n12836));
  nand_5 g10488(.A(new_n12836), .B(new_n10091), .Y(new_n12837));
  nand_5 g10489(.A(new_n12835), .B(new_n10092), .Y(new_n12838));
  nand_5 g10490(.A(new_n12766), .B(new_n12767), .Y(new_n12839));
  xor_4  g10491(.A(new_n12839), .B(new_n12807), .Y(new_n12840));
  not_8  g10492(.A(new_n12840), .Y(new_n12841));
  nand_5 g10493(.A(new_n12841), .B(new_n10099), .Y(new_n12842));
  nand_5 g10494(.A(new_n12840), .B(new_n10100), .Y(new_n12843_1));
  nand_5 g10495(.A(new_n12773), .B(new_n12774), .Y(new_n12844));
  xor_4  g10496(.A(new_n12844), .B(new_n12805), .Y(new_n12845));
  not_8  g10497(.A(new_n12845), .Y(new_n12846));
  nand_5 g10498(.A(new_n12846), .B(new_n10107), .Y(new_n12847));
  nand_5 g10499(.A(new_n12845), .B(new_n10108), .Y(new_n12848));
  nand_5 g10500(.A(new_n12777), .B(new_n12779), .Y(new_n12849));
  xor_4  g10501(.A(new_n12849), .B(new_n12803), .Y(new_n12850));
  not_8  g10502(.A(new_n12850), .Y(new_n12851));
  nand_5 g10503(.A(new_n12851), .B(new_n10115), .Y(new_n12852));
  nand_5 g10504(.A(new_n12850), .B(new_n10116), .Y(new_n12853));
  nand_5 g10505(.A(new_n12782), .B(new_n12783_1), .Y(new_n12854));
  xor_4  g10506(.A(new_n12854), .B(new_n12801_1), .Y(new_n12855));
  not_8  g10507(.A(new_n12855), .Y(new_n12856));
  nand_5 g10508(.A(new_n12856), .B(new_n10122), .Y(new_n12857));
  nand_5 g10509(.A(new_n12855), .B(new_n10123), .Y(new_n12858));
  nand_5 g10510(.A(new_n12786), .B(new_n12788), .Y(new_n12859));
  xor_4  g10511(.A(new_n12859), .B(new_n12799), .Y(new_n12860));
  not_8  g10512(.A(new_n12860), .Y(new_n12861_1));
  nand_5 g10513(.A(new_n12861_1), .B(new_n10129), .Y(new_n12862));
  nand_5 g10514(.A(new_n12860), .B(new_n10130), .Y(new_n12863));
  not_8  g10515(.A(new_n12795), .Y(new_n12864_1));
  nor_5  g10516(.A(new_n12794), .B(new_n4701), .Y(new_n12865_1));
  nor_5  g10517(.A(new_n12865_1), .B(new_n12864_1), .Y(new_n12866));
  nand_5 g10518(.A(new_n12866), .B(new_n10137), .Y(new_n12867));
  nand_5 g10519(.A(new_n12867), .B(new_n10144), .Y(new_n12868));
  or_5   g10520(.A(new_n12867), .B(new_n10144), .Y(new_n12869));
  nand_5 g10521(.A(new_n12796), .B(new_n12797), .Y(new_n12870_1));
  xor_4  g10522(.A(new_n12870_1), .B(new_n4695), .Y(new_n12871_1));
  nand_5 g10523(.A(new_n12871_1), .B(new_n12869), .Y(new_n12872));
  nand_5 g10524(.A(new_n12872), .B(new_n12868), .Y(new_n12873_1));
  nand_5 g10525(.A(new_n12873_1), .B(new_n12863), .Y(new_n12874));
  nand_5 g10526(.A(new_n12874), .B(new_n12862), .Y(new_n12875_1));
  nand_5 g10527(.A(new_n12875_1), .B(new_n12858), .Y(new_n12876));
  nand_5 g10528(.A(new_n12876), .B(new_n12857), .Y(new_n12877));
  nand_5 g10529(.A(new_n12877), .B(new_n12853), .Y(new_n12878));
  nand_5 g10530(.A(new_n12878), .B(new_n12852), .Y(new_n12879));
  nand_5 g10531(.A(new_n12879), .B(new_n12848), .Y(new_n12880));
  nand_5 g10532(.A(new_n12880), .B(new_n12847), .Y(new_n12881));
  nand_5 g10533(.A(new_n12881), .B(new_n12843_1), .Y(new_n12882));
  nand_5 g10534(.A(new_n12882), .B(new_n12842), .Y(new_n12883));
  nand_5 g10535(.A(new_n12883), .B(new_n12838), .Y(new_n12884));
  nand_5 g10536(.A(new_n12884), .B(new_n12837), .Y(new_n12885));
  nand_5 g10537(.A(new_n12885), .B(new_n12833), .Y(new_n12886));
  nand_5 g10538(.A(new_n12886), .B(new_n12832), .Y(new_n12887));
  nand_5 g10539(.A(new_n12887), .B(new_n12828), .Y(new_n12888));
  nand_5 g10540(.A(new_n12888), .B(new_n12827), .Y(new_n12889));
  nand_5 g10541(.A(new_n12889), .B(new_n12823), .Y(new_n12890));
  nand_5 g10542(.A(new_n12890), .B(new_n12821_1), .Y(new_n12891));
  xor_4  g10543(.A(new_n12891), .B(new_n12818), .Y(n1527));
  not_8  g10544(.A(new_n9029), .Y(new_n12893));
  nand_5 g10545(.A(new_n2585), .B(n10739), .Y(new_n12894));
  nand_5 g10546(.A(n13490), .B(new_n2601), .Y(new_n12895));
  nand_5 g10547(.A(new_n2467), .B(n21753), .Y(new_n12896));
  nand_5 g10548(.A(n22660), .B(new_n2518), .Y(new_n12897));
  nand_5 g10549(.A(n21832), .B(new_n2370), .Y(new_n12898));
  nand_5 g10550(.A(new_n2492), .B(n1777), .Y(new_n12899));
  nand_5 g10551(.A(n26913), .B(new_n2349), .Y(new_n12900_1));
  nand_5 g10552(.A(new_n2496), .B(n8745), .Y(new_n12901));
  nand_5 g10553(.A(new_n11280), .B(new_n11278), .Y(new_n12902));
  nand_5 g10554(.A(new_n12902), .B(new_n11279), .Y(new_n12903));
  nand_5 g10555(.A(new_n12903), .B(new_n12901), .Y(new_n12904_1));
  nand_5 g10556(.A(new_n12904_1), .B(new_n12900_1), .Y(new_n12905));
  nand_5 g10557(.A(new_n12905), .B(new_n12899), .Y(new_n12906));
  nand_5 g10558(.A(new_n12906), .B(new_n12898), .Y(new_n12907));
  nand_5 g10559(.A(new_n12907), .B(new_n12897), .Y(new_n12908));
  nand_5 g10560(.A(new_n12908), .B(new_n12896), .Y(new_n12909));
  nand_5 g10561(.A(new_n12909), .B(new_n12895), .Y(new_n12910));
  nand_5 g10562(.A(new_n12910), .B(new_n12894), .Y(new_n12911));
  nand_5 g10563(.A(n13074), .B(new_n6242), .Y(new_n12912));
  nand_5 g10564(.A(new_n3321), .B(n9655), .Y(new_n12913));
  nand_5 g10565(.A(new_n12913), .B(new_n12912), .Y(new_n12914));
  xor_4  g10566(.A(new_n12914), .B(new_n12911), .Y(new_n12915));
  or_5   g10567(.A(new_n12915), .B(new_n12893), .Y(new_n12916));
  nand_5 g10568(.A(new_n12915), .B(new_n12893), .Y(new_n12917_1));
  nand_5 g10569(.A(new_n12895), .B(new_n12894), .Y(new_n12918));
  xor_4  g10570(.A(new_n12918), .B(new_n12909), .Y(new_n12919));
  or_5   g10571(.A(new_n12919), .B(new_n9036), .Y(new_n12920));
  nand_5 g10572(.A(new_n12919), .B(new_n9036), .Y(new_n12921));
  nand_5 g10573(.A(new_n12897), .B(new_n12896), .Y(new_n12922));
  xor_4  g10574(.A(new_n12922), .B(new_n12907), .Y(new_n12923));
  or_5   g10575(.A(new_n12923), .B(new_n9044), .Y(new_n12924));
  nand_5 g10576(.A(new_n12923), .B(new_n9044), .Y(new_n12925));
  nand_5 g10577(.A(new_n12899), .B(new_n12898), .Y(new_n12926));
  xor_4  g10578(.A(new_n12926), .B(new_n12905), .Y(new_n12927));
  or_5   g10579(.A(new_n12927), .B(new_n9052), .Y(new_n12928));
  nand_5 g10580(.A(new_n12927), .B(new_n9052), .Y(new_n12929));
  nand_5 g10581(.A(new_n12901), .B(new_n12900_1), .Y(new_n12930));
  xor_4  g10582(.A(new_n12930), .B(new_n12903), .Y(new_n12931));
  or_5   g10583(.A(new_n12931), .B(new_n9060), .Y(new_n12932));
  nand_5 g10584(.A(new_n12931), .B(new_n9060), .Y(new_n12933));
  not_8  g10585(.A(new_n11276), .Y(new_n12934));
  nor_5  g10586(.A(new_n11285), .B(new_n12934), .Y(new_n12935));
  nor_5  g10587(.A(new_n12935), .B(new_n11284), .Y(new_n12936));
  not_8  g10588(.A(new_n12936), .Y(new_n12937));
  nand_5 g10589(.A(new_n12937), .B(new_n12933), .Y(new_n12938));
  nand_5 g10590(.A(new_n12938), .B(new_n12932), .Y(new_n12939));
  nand_5 g10591(.A(new_n12939), .B(new_n12929), .Y(new_n12940));
  nand_5 g10592(.A(new_n12940), .B(new_n12928), .Y(new_n12941_1));
  nand_5 g10593(.A(new_n12941_1), .B(new_n12925), .Y(new_n12942_1));
  nand_5 g10594(.A(new_n12942_1), .B(new_n12924), .Y(new_n12943));
  nand_5 g10595(.A(new_n12943), .B(new_n12921), .Y(new_n12944));
  nand_5 g10596(.A(new_n12944), .B(new_n12920), .Y(new_n12945));
  nand_5 g10597(.A(new_n12945), .B(new_n12917_1), .Y(new_n12946));
  nand_5 g10598(.A(new_n12946), .B(new_n12916), .Y(new_n12947));
  nand_5 g10599(.A(new_n12913), .B(new_n12911), .Y(new_n12948));
  nand_5 g10600(.A(new_n12948), .B(new_n12912), .Y(new_n12949));
  nand_5 g10601(.A(new_n6238), .B(n23463), .Y(new_n12950));
  nand_5 g10602(.A(n25345), .B(new_n3318), .Y(new_n12951));
  nand_5 g10603(.A(new_n12951), .B(new_n12950), .Y(new_n12952));
  xnor_4 g10604(.A(new_n12952), .B(new_n12949), .Y(new_n12953));
  nand_5 g10605(.A(new_n12953), .B(new_n9023), .Y(new_n12954));
  or_5   g10606(.A(new_n12953), .B(new_n9023), .Y(new_n12955));
  nand_5 g10607(.A(new_n12955), .B(new_n12954), .Y(new_n12956_1));
  xnor_4 g10608(.A(new_n12956_1), .B(new_n12947), .Y(n1580));
  not_8  g10609(.A(new_n8535_1), .Y(new_n12958));
  xor_4  g10610(.A(n18962), .B(new_n2443), .Y(new_n12959));
  not_8  g10611(.A(new_n12959), .Y(new_n12960));
  nand_5 g10612(.A(new_n12960), .B(new_n12958), .Y(new_n12961));
  not_8  g10613(.A(new_n12961), .Y(new_n12962));
  nand_5 g10614(.A(n18962), .B(new_n2443), .Y(new_n12963));
  nand_5 g10615(.A(new_n7741), .B(n3952), .Y(new_n12964));
  nand_5 g10616(.A(n10158), .B(new_n2357), .Y(new_n12965));
  nand_5 g10617(.A(new_n12965), .B(new_n12964), .Y(new_n12966));
  xnor_4 g10618(.A(new_n12966), .B(new_n12963), .Y(new_n12967));
  nand_5 g10619(.A(new_n12967), .B(new_n12962), .Y(new_n12968));
  nor_5  g10620(.A(new_n12967), .B(new_n12962), .Y(new_n12969));
  not_8  g10621(.A(new_n12969), .Y(new_n12970));
  nand_5 g10622(.A(new_n12970), .B(new_n12968), .Y(new_n12971));
  xor_4  g10623(.A(new_n12971), .B(new_n8543), .Y(n1586));
  not_8  g10624(.A(n10117), .Y(new_n12973));
  nand_5 g10625(.A(new_n12973), .B(n3306), .Y(new_n12974));
  or_5   g10626(.A(new_n12973), .B(n3306), .Y(new_n12975));
  not_8  g10627(.A(n13460), .Y(new_n12976));
  nand_5 g10628(.A(n22335), .B(new_n12976), .Y(new_n12977));
  nor_5  g10629(.A(n22335), .B(new_n12976), .Y(new_n12978_1));
  not_8  g10630(.A(new_n12978_1), .Y(new_n12979));
  not_8  g10631(.A(n6104), .Y(new_n12980_1));
  nand_5 g10632(.A(n24048), .B(new_n12980_1), .Y(new_n12981));
  nor_5  g10633(.A(n24048), .B(new_n12980_1), .Y(new_n12982));
  not_8  g10634(.A(new_n12982), .Y(new_n12983));
  nand_5 g10635(.A(new_n5295), .B(new_n5291), .Y(new_n12984));
  nand_5 g10636(.A(new_n12984), .B(new_n5294), .Y(new_n12985_1));
  nand_5 g10637(.A(new_n12985_1), .B(new_n12983), .Y(new_n12986));
  nand_5 g10638(.A(new_n12986), .B(new_n12981), .Y(new_n12987_1));
  nand_5 g10639(.A(new_n12987_1), .B(new_n12979), .Y(new_n12988));
  nand_5 g10640(.A(new_n12988), .B(new_n12977), .Y(new_n12989));
  nand_5 g10641(.A(new_n12989), .B(new_n12975), .Y(new_n12990));
  nand_5 g10642(.A(new_n12990), .B(new_n12974), .Y(new_n12991));
  not_8  g10643(.A(new_n12991), .Y(new_n12992_1));
  not_8  g10644(.A(n25494), .Y(new_n12993));
  nand_5 g10645(.A(new_n12993), .B(n1314), .Y(new_n12994));
  or_5   g10646(.A(new_n12993), .B(n1314), .Y(new_n12995));
  nand_5 g10647(.A(new_n12995), .B(new_n12994), .Y(new_n12996));
  xor_4  g10648(.A(new_n12996), .B(new_n12992_1), .Y(new_n12997));
  not_8  g10649(.A(n23717), .Y(new_n12998));
  or_5   g10650(.A(n25296), .B(new_n12998), .Y(new_n12999));
  nand_5 g10651(.A(n25296), .B(new_n12998), .Y(new_n13000));
  nand_5 g10652(.A(new_n13000), .B(new_n12999), .Y(new_n13001));
  not_8  g10653(.A(n7788), .Y(new_n13002));
  or_5   g10654(.A(n20013), .B(new_n13002), .Y(new_n13003));
  nand_5 g10655(.A(n20013), .B(new_n13002), .Y(new_n13004));
  not_8  g10656(.A(n1320), .Y(new_n13005_1));
  nand_5 g10657(.A(n5443), .B(new_n13005_1), .Y(new_n13006));
  nor_5  g10658(.A(n5443), .B(new_n13005_1), .Y(new_n13007));
  not_8  g10659(.A(new_n13007), .Y(new_n13008));
  nand_5 g10660(.A(new_n7471), .B(new_n7467), .Y(new_n13009));
  nand_5 g10661(.A(new_n13009), .B(new_n7470), .Y(new_n13010));
  nand_5 g10662(.A(new_n13010), .B(new_n13008), .Y(new_n13011));
  nand_5 g10663(.A(new_n13011), .B(new_n13006), .Y(new_n13012));
  nand_5 g10664(.A(new_n13012), .B(new_n13004), .Y(new_n13013));
  nand_5 g10665(.A(new_n13013), .B(new_n13003), .Y(new_n13014));
  not_8  g10666(.A(new_n13014), .Y(new_n13015));
  xor_4  g10667(.A(new_n13015), .B(new_n13001), .Y(new_n13016));
  nand_5 g10668(.A(new_n13016), .B(new_n12997), .Y(new_n13017));
  not_8  g10669(.A(new_n12997), .Y(new_n13018));
  not_8  g10670(.A(new_n13016), .Y(new_n13019));
  nand_5 g10671(.A(new_n13019), .B(new_n13018), .Y(new_n13020));
  nand_5 g10672(.A(new_n13020), .B(new_n13017), .Y(new_n13021));
  nand_5 g10673(.A(new_n12975), .B(new_n12974), .Y(new_n13022));
  xor_4  g10674(.A(new_n13022), .B(new_n12989), .Y(new_n13023));
  nand_5 g10675(.A(new_n13004), .B(new_n13003), .Y(new_n13024));
  xor_4  g10676(.A(new_n13024), .B(new_n13012), .Y(new_n13025));
  nand_5 g10677(.A(new_n13025), .B(new_n13023), .Y(new_n13026_1));
  not_8  g10678(.A(new_n13023), .Y(new_n13027));
  not_8  g10679(.A(new_n13025), .Y(new_n13028));
  nand_5 g10680(.A(new_n13028), .B(new_n13027), .Y(new_n13029));
  nand_5 g10681(.A(new_n12979), .B(new_n12977), .Y(new_n13030));
  xor_4  g10682(.A(new_n13030), .B(new_n12987_1), .Y(new_n13031));
  nand_5 g10683(.A(new_n13008), .B(new_n13006), .Y(new_n13032));
  xor_4  g10684(.A(new_n13032), .B(new_n13010), .Y(new_n13033));
  nand_5 g10685(.A(new_n13033), .B(new_n13031), .Y(new_n13034));
  or_5   g10686(.A(new_n13033), .B(new_n13031), .Y(new_n13035));
  nand_5 g10687(.A(new_n12983), .B(new_n12981), .Y(new_n13036));
  xor_4  g10688(.A(new_n13036), .B(new_n12985_1), .Y(new_n13037));
  nand_5 g10689(.A(new_n13037), .B(new_n7474), .Y(new_n13038));
  not_8  g10690(.A(new_n13037), .Y(new_n13039));
  nand_5 g10691(.A(new_n13039), .B(new_n7473), .Y(new_n13040));
  nand_5 g10692(.A(new_n5310), .B(new_n5289), .Y(new_n13041));
  nand_5 g10693(.A(new_n13041), .B(new_n5309), .Y(new_n13042));
  nand_5 g10694(.A(new_n13042), .B(new_n13040), .Y(new_n13043_1));
  nand_5 g10695(.A(new_n13043_1), .B(new_n13038), .Y(new_n13044_1));
  nand_5 g10696(.A(new_n13044_1), .B(new_n13035), .Y(new_n13045));
  nand_5 g10697(.A(new_n13045), .B(new_n13034), .Y(new_n13046));
  nand_5 g10698(.A(new_n13046), .B(new_n13029), .Y(new_n13047));
  nand_5 g10699(.A(new_n13047), .B(new_n13026_1), .Y(new_n13048_1));
  xor_4  g10700(.A(new_n13048_1), .B(new_n13021), .Y(new_n13049));
  not_8  g10701(.A(n1483), .Y(new_n13050));
  nand_5 g10702(.A(n19539), .B(new_n13050), .Y(new_n13051));
  nor_5  g10703(.A(n19539), .B(new_n13050), .Y(new_n13052));
  not_8  g10704(.A(new_n13052), .Y(new_n13053));
  nand_5 g10705(.A(new_n13053), .B(new_n13051), .Y(new_n13054_1));
  not_8  g10706(.A(n8194), .Y(new_n13055));
  or_5   g10707(.A(n24093), .B(new_n13055), .Y(new_n13056));
  nand_5 g10708(.A(n24093), .B(new_n13055), .Y(new_n13057));
  not_8  g10709(.A(n23035), .Y(new_n13058));
  nand_5 g10710(.A(n23657), .B(new_n13058), .Y(new_n13059));
  nor_5  g10711(.A(n23657), .B(new_n13058), .Y(new_n13060));
  not_8  g10712(.A(new_n13060), .Y(new_n13061));
  nand_5 g10713(.A(new_n7484), .B(new_n7479), .Y(new_n13062));
  nand_5 g10714(.A(new_n13062), .B(new_n7482), .Y(new_n13063));
  nand_5 g10715(.A(new_n13063), .B(new_n13061), .Y(new_n13064));
  nand_5 g10716(.A(new_n13064), .B(new_n13059), .Y(new_n13065));
  nand_5 g10717(.A(new_n13065), .B(new_n13057), .Y(new_n13066));
  nand_5 g10718(.A(new_n13066), .B(new_n13056), .Y(new_n13067));
  not_8  g10719(.A(new_n13067), .Y(new_n13068));
  xor_4  g10720(.A(new_n13068), .B(new_n13054_1), .Y(new_n13069));
  nand_5 g10721(.A(new_n13069), .B(new_n13049), .Y(new_n13070));
  or_5   g10722(.A(new_n13069), .B(new_n13049), .Y(new_n13071));
  nand_5 g10723(.A(new_n13071), .B(new_n13070), .Y(new_n13072));
  nand_5 g10724(.A(new_n13057), .B(new_n13056), .Y(new_n13073));
  xor_4  g10725(.A(new_n13073), .B(new_n13065), .Y(new_n13074_1));
  not_8  g10726(.A(new_n13074_1), .Y(new_n13075));
  nand_5 g10727(.A(new_n13026_1), .B(new_n13029), .Y(new_n13076));
  xor_4  g10728(.A(new_n13076), .B(new_n13046), .Y(new_n13077));
  nand_5 g10729(.A(new_n13077), .B(new_n13075), .Y(new_n13078));
  not_8  g10730(.A(new_n13077), .Y(new_n13079));
  nand_5 g10731(.A(new_n13079), .B(new_n13074_1), .Y(new_n13080));
  nand_5 g10732(.A(new_n13061), .B(new_n13059), .Y(new_n13081));
  xor_4  g10733(.A(new_n13081), .B(new_n13063), .Y(new_n13082_1));
  not_8  g10734(.A(new_n13082_1), .Y(new_n13083));
  nand_5 g10735(.A(new_n13034), .B(new_n13035), .Y(new_n13084));
  xor_4  g10736(.A(new_n13084), .B(new_n13044_1), .Y(new_n13085));
  nand_5 g10737(.A(new_n13085), .B(new_n13083), .Y(new_n13086));
  not_8  g10738(.A(new_n13085), .Y(new_n13087));
  nand_5 g10739(.A(new_n13087), .B(new_n13082_1), .Y(new_n13088));
  nand_5 g10740(.A(new_n13038), .B(new_n13040), .Y(new_n13089));
  xor_4  g10741(.A(new_n13089), .B(new_n13042), .Y(new_n13090));
  nand_5 g10742(.A(new_n13090), .B(new_n7486), .Y(new_n13091));
  not_8  g10743(.A(new_n13090), .Y(new_n13092));
  nand_5 g10744(.A(new_n13092), .B(new_n7487), .Y(new_n13093));
  nand_5 g10745(.A(new_n7413), .B(new_n5312), .Y(new_n13094));
  or_5   g10746(.A(new_n7413), .B(new_n5312), .Y(new_n13095));
  nand_5 g10747(.A(new_n7328), .B(new_n5222), .Y(new_n13096_1));
  nand_5 g10748(.A(new_n7327), .B(new_n5223), .Y(new_n13097));
  nand_5 g10749(.A(new_n7375), .B(new_n5253), .Y(new_n13098));
  nand_5 g10750(.A(new_n7374), .B(new_n5254), .Y(new_n13099));
  nand_5 g10751(.A(new_n7381), .B(new_n5260), .Y(new_n13100));
  or_5   g10752(.A(new_n7381), .B(new_n5260), .Y(new_n13101));
  nand_5 g10753(.A(new_n7390_1), .B(new_n5266), .Y(new_n13102));
  or_5   g10754(.A(new_n13102), .B(new_n7387), .Y(new_n13103));
  nand_5 g10755(.A(new_n13102), .B(new_n7387), .Y(new_n13104));
  nand_5 g10756(.A(new_n13104), .B(new_n5276), .Y(new_n13105));
  nand_5 g10757(.A(new_n13105), .B(new_n13103), .Y(new_n13106));
  nand_5 g10758(.A(new_n13106), .B(new_n13101), .Y(new_n13107));
  nand_5 g10759(.A(new_n13107), .B(new_n13100), .Y(new_n13108));
  nand_5 g10760(.A(new_n13108), .B(new_n13099), .Y(new_n13109));
  nand_5 g10761(.A(new_n13109), .B(new_n13098), .Y(new_n13110_1));
  nand_5 g10762(.A(new_n13110_1), .B(new_n13097), .Y(new_n13111));
  nand_5 g10763(.A(new_n13111), .B(new_n13096_1), .Y(new_n13112));
  nand_5 g10764(.A(new_n13112), .B(new_n13095), .Y(new_n13113));
  nand_5 g10765(.A(new_n13113), .B(new_n13094), .Y(new_n13114));
  nand_5 g10766(.A(new_n13114), .B(new_n13093), .Y(new_n13115));
  nand_5 g10767(.A(new_n13115), .B(new_n13091), .Y(new_n13116_1));
  nand_5 g10768(.A(new_n13116_1), .B(new_n13088), .Y(new_n13117));
  nand_5 g10769(.A(new_n13117), .B(new_n13086), .Y(new_n13118));
  nand_5 g10770(.A(new_n13118), .B(new_n13080), .Y(new_n13119));
  nand_5 g10771(.A(new_n13119), .B(new_n13078), .Y(new_n13120));
  not_8  g10772(.A(new_n13120), .Y(new_n13121));
  xor_4  g10773(.A(new_n13121), .B(new_n13072), .Y(n1590));
  nand_5 g10774(.A(new_n8728), .B(new_n8727), .Y(new_n13123));
  xor_4  g10775(.A(new_n13123), .B(new_n8742), .Y(n1602));
  nand_5 g10776(.A(new_n2922), .B(new_n2921), .Y(new_n13125));
  xnor_4 g10777(.A(new_n13125), .B(new_n2992), .Y(n1634));
  nand_5 g10778(.A(new_n13078), .B(new_n13080), .Y(new_n13127));
  xnor_4 g10779(.A(new_n13127), .B(new_n13118), .Y(n1636));
  nand_5 g10780(.A(new_n7960), .B(new_n7956), .Y(new_n13129));
  nand_5 g10781(.A(new_n13129), .B(new_n7959_1), .Y(new_n13130));
  nand_5 g10782(.A(new_n13130), .B(new_n8648), .Y(new_n13131));
  not_8  g10783(.A(new_n13131), .Y(new_n13132));
  nor_5  g10784(.A(new_n13130), .B(new_n8648), .Y(new_n13133));
  nor_5  g10785(.A(new_n13133), .B(n18880), .Y(new_n13134));
  nor_5  g10786(.A(new_n13134), .B(new_n13132), .Y(new_n13135));
  not_8  g10787(.A(new_n13135), .Y(new_n13136));
  nor_5  g10788(.A(new_n13133), .B(new_n13132), .Y(new_n13137_1));
  xor_4  g10789(.A(new_n13137_1), .B(new_n4966_1), .Y(new_n13138));
  nand_5 g10790(.A(new_n13138), .B(new_n2648), .Y(new_n13139));
  not_8  g10791(.A(new_n13138), .Y(new_n13140));
  nand_5 g10792(.A(new_n13140), .B(n20040), .Y(new_n13141_1));
  nand_5 g10793(.A(new_n7962), .B(new_n2652), .Y(new_n13142));
  nand_5 g10794(.A(new_n7963_1), .B(n19531), .Y(new_n13143));
  nand_5 g10795(.A(new_n7813), .B(new_n10043), .Y(new_n13144_1));
  nand_5 g10796(.A(new_n7814), .B(n18345), .Y(new_n13145));
  nand_5 g10797(.A(new_n7760), .B(new_n2658), .Y(new_n13146));
  nand_5 g10798(.A(new_n7761), .B(n13190), .Y(new_n13147));
  nand_5 g10799(.A(new_n7767), .B(new_n10048), .Y(new_n13148));
  nand_5 g10800(.A(new_n7765), .B(n3460), .Y(new_n13149));
  nand_5 g10801(.A(new_n11075), .B(new_n11072), .Y(new_n13150));
  nand_5 g10802(.A(new_n13150), .B(new_n11074), .Y(new_n13151));
  nand_5 g10803(.A(new_n13151), .B(new_n13149), .Y(new_n13152));
  nand_5 g10804(.A(new_n13152), .B(new_n13148), .Y(new_n13153));
  nand_5 g10805(.A(new_n13153), .B(new_n13147), .Y(new_n13154));
  nand_5 g10806(.A(new_n13154), .B(new_n13146), .Y(new_n13155));
  nand_5 g10807(.A(new_n13155), .B(new_n13145), .Y(new_n13156));
  nand_5 g10808(.A(new_n13156), .B(new_n13144_1), .Y(new_n13157));
  nand_5 g10809(.A(new_n13157), .B(new_n13143), .Y(new_n13158));
  nand_5 g10810(.A(new_n13158), .B(new_n13142), .Y(new_n13159));
  nand_5 g10811(.A(new_n13159), .B(new_n13141_1), .Y(new_n13160));
  nand_5 g10812(.A(new_n13160), .B(new_n13139), .Y(new_n13161));
  nor_5  g10813(.A(new_n13161), .B(new_n13136), .Y(new_n13162));
  not_8  g10814(.A(new_n13162), .Y(new_n13163));
  nand_5 g10815(.A(new_n13161), .B(new_n13136), .Y(new_n13164));
  and_5  g10816(.A(new_n13164), .B(new_n13163), .Y(new_n13165));
  not_8  g10817(.A(n17037), .Y(new_n13166));
  not_8  g10818(.A(n26191), .Y(new_n13167));
  nor_5  g10819(.A(new_n11079), .B(n26512), .Y(new_n13168_1));
  nand_5 g10820(.A(new_n13168_1), .B(new_n13167), .Y(new_n13169));
  nor_5  g10821(.A(new_n13169), .B(n5386), .Y(new_n13170));
  nand_5 g10822(.A(new_n13170), .B(new_n13166), .Y(new_n13171));
  nor_5  g10823(.A(new_n13171), .B(n7569), .Y(new_n13172));
  xor_4  g10824(.A(new_n13172), .B(new_n13165), .Y(new_n13173));
  nand_5 g10825(.A(new_n13139), .B(new_n13141_1), .Y(new_n13174));
  xor_4  g10826(.A(new_n13174), .B(new_n13159), .Y(new_n13175));
  not_8  g10827(.A(new_n13175), .Y(new_n13176));
  not_8  g10828(.A(new_n13172), .Y(new_n13177));
  nand_5 g10829(.A(new_n13171), .B(n7569), .Y(new_n13178));
  nand_5 g10830(.A(new_n13178), .B(new_n13177), .Y(new_n13179));
  or_5   g10831(.A(new_n13179), .B(new_n13176), .Y(new_n13180));
  nand_5 g10832(.A(new_n13179), .B(new_n13176), .Y(new_n13181));
  nand_5 g10833(.A(new_n13142), .B(new_n13143), .Y(new_n13182));
  xor_4  g10834(.A(new_n13182), .B(new_n13157), .Y(new_n13183));
  not_8  g10835(.A(new_n13183), .Y(new_n13184));
  xor_4  g10836(.A(new_n13170), .B(n17037), .Y(new_n13185));
  or_5   g10837(.A(new_n13185), .B(new_n13184), .Y(new_n13186));
  nand_5 g10838(.A(new_n13185), .B(new_n13184), .Y(new_n13187));
  nand_5 g10839(.A(new_n13144_1), .B(new_n13145), .Y(new_n13188));
  xor_4  g10840(.A(new_n13188), .B(new_n13155), .Y(new_n13189));
  not_8  g10841(.A(new_n13189), .Y(new_n13190_1));
  not_8  g10842(.A(n5386), .Y(new_n13191));
  xor_4  g10843(.A(new_n13169), .B(new_n13191), .Y(new_n13192));
  or_5   g10844(.A(new_n13192), .B(new_n13190_1), .Y(new_n13193));
  nand_5 g10845(.A(new_n13192), .B(new_n13190_1), .Y(new_n13194));
  nand_5 g10846(.A(new_n13146), .B(new_n13147), .Y(new_n13195));
  xor_4  g10847(.A(new_n13195), .B(new_n13153), .Y(new_n13196));
  not_8  g10848(.A(new_n13196), .Y(new_n13197));
  xor_4  g10849(.A(new_n13168_1), .B(n26191), .Y(new_n13198_1));
  or_5   g10850(.A(new_n13198_1), .B(new_n13197), .Y(new_n13199_1));
  nand_5 g10851(.A(new_n13198_1), .B(new_n13197), .Y(new_n13200));
  nand_5 g10852(.A(new_n13148), .B(new_n13149), .Y(new_n13201));
  xor_4  g10853(.A(new_n13201), .B(new_n13151), .Y(new_n13202));
  xor_4  g10854(.A(new_n11079), .B(n26512), .Y(new_n13203));
  nand_5 g10855(.A(new_n13203), .B(new_n13202), .Y(new_n13204_1));
  or_5   g10856(.A(new_n13203), .B(new_n13202), .Y(new_n13205));
  nand_5 g10857(.A(new_n11083), .B(new_n11070), .Y(new_n13206));
  nand_5 g10858(.A(new_n13206), .B(new_n11082), .Y(new_n13207));
  nand_5 g10859(.A(new_n13207), .B(new_n13205), .Y(new_n13208));
  nand_5 g10860(.A(new_n13208), .B(new_n13204_1), .Y(new_n13209_1));
  nand_5 g10861(.A(new_n13209_1), .B(new_n13200), .Y(new_n13210));
  nand_5 g10862(.A(new_n13210), .B(new_n13199_1), .Y(new_n13211));
  nand_5 g10863(.A(new_n13211), .B(new_n13194), .Y(new_n13212));
  nand_5 g10864(.A(new_n13212), .B(new_n13193), .Y(new_n13213));
  nand_5 g10865(.A(new_n13213), .B(new_n13187), .Y(new_n13214));
  nand_5 g10866(.A(new_n13214), .B(new_n13186), .Y(new_n13215));
  nand_5 g10867(.A(new_n13215), .B(new_n13181), .Y(new_n13216));
  nand_5 g10868(.A(new_n13216), .B(new_n13180), .Y(new_n13217));
  xor_4  g10869(.A(new_n13217), .B(new_n13173), .Y(new_n13218));
  not_8  g10870(.A(n4514), .Y(new_n13219));
  not_8  g10871(.A(n10514), .Y(new_n13220));
  nand_5 g10872(.A(new_n13220), .B(new_n13219), .Y(new_n13221));
  nand_5 g10873(.A(n10514), .B(n4514), .Y(new_n13222));
  not_8  g10874(.A(n3984), .Y(new_n13223));
  not_8  g10875(.A(n18649), .Y(new_n13224));
  nand_5 g10876(.A(new_n13224), .B(new_n13223), .Y(new_n13225));
  nand_5 g10877(.A(n18649), .B(n3984), .Y(new_n13226));
  not_8  g10878(.A(n6218), .Y(new_n13227));
  not_8  g10879(.A(n19652), .Y(new_n13228));
  nand_5 g10880(.A(new_n13228), .B(new_n13227), .Y(new_n13229));
  nand_5 g10881(.A(n19652), .B(n6218), .Y(new_n13230));
  nand_5 g10882(.A(new_n12634), .B(new_n12629), .Y(new_n13231));
  nand_5 g10883(.A(new_n13231), .B(new_n12633), .Y(new_n13232));
  nand_5 g10884(.A(new_n13232), .B(new_n13230), .Y(new_n13233));
  nand_5 g10885(.A(new_n13233), .B(new_n13229), .Y(new_n13234));
  nand_5 g10886(.A(new_n13234), .B(new_n13226), .Y(new_n13235));
  nand_5 g10887(.A(new_n13235), .B(new_n13225), .Y(new_n13236));
  nand_5 g10888(.A(new_n13236), .B(new_n13222), .Y(new_n13237));
  nand_5 g10889(.A(new_n13237), .B(new_n13221), .Y(new_n13238));
  not_8  g10890(.A(new_n13238), .Y(new_n13239));
  or_5   g10891(.A(new_n13239), .B(new_n13218), .Y(new_n13240));
  nand_5 g10892(.A(new_n13239), .B(new_n13218), .Y(new_n13241));
  nand_5 g10893(.A(new_n13241), .B(new_n13240), .Y(new_n13242));
  nand_5 g10894(.A(new_n13222), .B(new_n13221), .Y(new_n13243));
  xor_4  g10895(.A(new_n13243), .B(new_n13236), .Y(new_n13244));
  nand_5 g10896(.A(new_n13181), .B(new_n13180), .Y(new_n13245));
  xor_4  g10897(.A(new_n13245), .B(new_n13215), .Y(new_n13246));
  nand_5 g10898(.A(new_n13246), .B(new_n13244), .Y(new_n13247));
  or_5   g10899(.A(new_n13246), .B(new_n13244), .Y(new_n13248));
  nand_5 g10900(.A(new_n13226), .B(new_n13225), .Y(new_n13249));
  xor_4  g10901(.A(new_n13249), .B(new_n13234), .Y(new_n13250));
  nand_5 g10902(.A(new_n13187), .B(new_n13186), .Y(new_n13251));
  xor_4  g10903(.A(new_n13251), .B(new_n13213), .Y(new_n13252));
  nand_5 g10904(.A(new_n13252), .B(new_n13250), .Y(new_n13253));
  or_5   g10905(.A(new_n13252), .B(new_n13250), .Y(new_n13254));
  nand_5 g10906(.A(new_n13230), .B(new_n13229), .Y(new_n13255));
  xor_4  g10907(.A(new_n13255), .B(new_n13232), .Y(new_n13256));
  nand_5 g10908(.A(new_n13194), .B(new_n13193), .Y(new_n13257));
  xor_4  g10909(.A(new_n13257), .B(new_n13211), .Y(new_n13258));
  nand_5 g10910(.A(new_n13258), .B(new_n13256), .Y(new_n13259));
  or_5   g10911(.A(new_n13258), .B(new_n13256), .Y(new_n13260));
  nand_5 g10912(.A(new_n13200), .B(new_n13199_1), .Y(new_n13261));
  xor_4  g10913(.A(new_n13261), .B(new_n13209_1), .Y(new_n13262));
  not_8  g10914(.A(new_n13262), .Y(new_n13263_1));
  or_5   g10915(.A(new_n13263_1), .B(new_n12636), .Y(new_n13264));
  nand_5 g10916(.A(new_n13263_1), .B(new_n12636), .Y(new_n13265));
  nand_5 g10917(.A(new_n13205), .B(new_n13204_1), .Y(new_n13266));
  xor_4  g10918(.A(new_n13266), .B(new_n13207), .Y(new_n13267));
  nand_5 g10919(.A(new_n13267), .B(new_n12544), .Y(new_n13268));
  nor_5  g10920(.A(new_n13267), .B(new_n12544), .Y(new_n13269));
  not_8  g10921(.A(new_n13269), .Y(new_n13270_1));
  nand_5 g10922(.A(new_n11087), .B(new_n11059), .Y(new_n13271));
  nand_5 g10923(.A(new_n13271), .B(new_n11086), .Y(new_n13272));
  nand_5 g10924(.A(new_n13272), .B(new_n13270_1), .Y(new_n13273_1));
  nand_5 g10925(.A(new_n13273_1), .B(new_n13268), .Y(new_n13274));
  nand_5 g10926(.A(new_n13274), .B(new_n13265), .Y(new_n13275));
  nand_5 g10927(.A(new_n13275), .B(new_n13264), .Y(new_n13276));
  nand_5 g10928(.A(new_n13276), .B(new_n13260), .Y(new_n13277));
  nand_5 g10929(.A(new_n13277), .B(new_n13259), .Y(new_n13278));
  nand_5 g10930(.A(new_n13278), .B(new_n13254), .Y(new_n13279));
  nand_5 g10931(.A(new_n13279), .B(new_n13253), .Y(new_n13280));
  nand_5 g10932(.A(new_n13280), .B(new_n13248), .Y(new_n13281));
  nand_5 g10933(.A(new_n13281), .B(new_n13247), .Y(new_n13282));
  xor_4  g10934(.A(new_n13282), .B(new_n13242), .Y(n1684));
  not_8  g10935(.A(n23912), .Y(new_n13284));
  nand_5 g10936(.A(new_n7059), .B(n3984), .Y(new_n13285_1));
  nand_5 g10937(.A(new_n7057_1), .B(new_n13223), .Y(new_n13286));
  nand_5 g10938(.A(new_n13286), .B(new_n13285_1), .Y(new_n13287));
  nand_5 g10939(.A(new_n7062), .B(new_n13228), .Y(new_n13288));
  nand_5 g10940(.A(new_n7064), .B(n19652), .Y(new_n13289));
  nand_5 g10941(.A(new_n7068), .B(new_n12631), .Y(new_n13290));
  nand_5 g10942(.A(new_n7067), .B(n3366), .Y(new_n13291));
  nand_5 g10943(.A(new_n4517), .B(new_n12540_1), .Y(new_n13292));
  nand_5 g10944(.A(new_n4516), .B(n26565), .Y(new_n13293));
  nand_5 g10945(.A(new_n4443), .B(new_n11062), .Y(new_n13294));
  nand_5 g10946(.A(new_n4442), .B(n3959), .Y(new_n13295));
  nand_5 g10947(.A(new_n4401_1), .B(new_n10983), .Y(new_n13296));
  nand_5 g10948(.A(new_n4400), .B(n11566), .Y(new_n13297));
  nand_5 g10949(.A(new_n4383), .B(new_n10970), .Y(new_n13298));
  nand_5 g10950(.A(new_n4382), .B(n26744), .Y(new_n13299));
  nand_5 g10951(.A(new_n4389), .B(new_n10974), .Y(new_n13300));
  nand_5 g10952(.A(new_n4388), .B(n26625), .Y(new_n13301));
  nand_5 g10953(.A(n19922), .B(n14230), .Y(new_n13302));
  nand_5 g10954(.A(new_n13302), .B(new_n13301), .Y(new_n13303));
  nand_5 g10955(.A(new_n13303), .B(new_n13300), .Y(new_n13304));
  nand_5 g10956(.A(new_n13304), .B(new_n13299), .Y(new_n13305));
  nand_5 g10957(.A(new_n13305), .B(new_n13298), .Y(new_n13306));
  nand_5 g10958(.A(new_n13306), .B(new_n13297), .Y(new_n13307));
  nand_5 g10959(.A(new_n13307), .B(new_n13296), .Y(new_n13308));
  nand_5 g10960(.A(new_n13308), .B(new_n13295), .Y(new_n13309));
  nand_5 g10961(.A(new_n13309), .B(new_n13294), .Y(new_n13310));
  nand_5 g10962(.A(new_n13310), .B(new_n13293), .Y(new_n13311));
  nand_5 g10963(.A(new_n13311), .B(new_n13292), .Y(new_n13312));
  nand_5 g10964(.A(new_n13312), .B(new_n13291), .Y(new_n13313));
  nand_5 g10965(.A(new_n13313), .B(new_n13290), .Y(new_n13314));
  nand_5 g10966(.A(new_n13314), .B(new_n13289), .Y(new_n13315));
  nand_5 g10967(.A(new_n13315), .B(new_n13288), .Y(new_n13316));
  xnor_4 g10968(.A(new_n13316), .B(new_n13287), .Y(new_n13317));
  or_5   g10969(.A(new_n13317), .B(n13026), .Y(new_n13318));
  nand_5 g10970(.A(new_n13317), .B(n13026), .Y(new_n13319_1));
  nand_5 g10971(.A(new_n13289), .B(new_n13288), .Y(new_n13320));
  xor_4  g10972(.A(new_n13320), .B(new_n13314), .Y(new_n13321));
  not_8  g10973(.A(new_n13321), .Y(new_n13322));
  or_5   g10974(.A(new_n13322), .B(n2175), .Y(new_n13323));
  nand_5 g10975(.A(new_n13322), .B(n2175), .Y(new_n13324));
  nand_5 g10976(.A(new_n13291), .B(new_n13290), .Y(new_n13325));
  xor_4  g10977(.A(new_n13325), .B(new_n13312), .Y(new_n13326));
  not_8  g10978(.A(new_n13326), .Y(new_n13327));
  or_5   g10979(.A(new_n13327), .B(n752), .Y(new_n13328));
  nand_5 g10980(.A(new_n13327), .B(n752), .Y(new_n13329));
  nand_5 g10981(.A(new_n13293), .B(new_n13292), .Y(new_n13330));
  xor_4  g10982(.A(new_n13330), .B(new_n13310), .Y(new_n13331));
  nand_5 g10983(.A(new_n13331), .B(new_n12584), .Y(new_n13332));
  or_5   g10984(.A(new_n13331), .B(new_n12584), .Y(new_n13333_1));
  nand_5 g10985(.A(new_n13295), .B(new_n13294), .Y(new_n13334));
  xor_4  g10986(.A(new_n13334), .B(new_n13308), .Y(new_n13335));
  nand_5 g10987(.A(new_n13335), .B(new_n12545_1), .Y(new_n13336));
  or_5   g10988(.A(new_n13335), .B(new_n12545_1), .Y(new_n13337));
  nand_5 g10989(.A(new_n13297), .B(new_n13296), .Y(new_n13338_1));
  xor_4  g10990(.A(new_n13338_1), .B(new_n13306), .Y(new_n13339));
  nand_5 g10991(.A(new_n13339), .B(new_n12559), .Y(new_n13340));
  or_5   g10992(.A(new_n13339), .B(new_n12559), .Y(new_n13341));
  not_8  g10993(.A(n5131), .Y(new_n13342));
  nand_5 g10994(.A(new_n13299), .B(new_n13298), .Y(new_n13343));
  xor_4  g10995(.A(new_n13343), .B(new_n13304), .Y(new_n13344));
  nand_5 g10996(.A(new_n13344), .B(new_n13342), .Y(new_n13345));
  nor_5  g10997(.A(new_n13344), .B(new_n13342), .Y(new_n13346));
  not_8  g10998(.A(new_n13346), .Y(new_n13347));
  nand_5 g10999(.A(new_n13301), .B(new_n13300), .Y(new_n13348));
  xnor_4 g11000(.A(new_n13348), .B(new_n13302), .Y(new_n13349));
  nand_5 g11001(.A(new_n13349), .B(n11473), .Y(new_n13350));
  nand_5 g11002(.A(new_n4378), .B(new_n7513), .Y(new_n13351));
  and_5  g11003(.A(new_n13351), .B(new_n13302), .Y(new_n13352));
  or_5   g11004(.A(new_n13352), .B(new_n12547), .Y(new_n13353));
  nand_5 g11005(.A(new_n13353), .B(new_n13350), .Y(new_n13354));
  nor_5  g11006(.A(new_n13349), .B(n11473), .Y(new_n13355));
  not_8  g11007(.A(new_n13355), .Y(new_n13356));
  nand_5 g11008(.A(new_n13356), .B(new_n13354), .Y(new_n13357));
  nand_5 g11009(.A(new_n13357), .B(new_n13347), .Y(new_n13358));
  nand_5 g11010(.A(new_n13358), .B(new_n13345), .Y(new_n13359));
  nand_5 g11011(.A(new_n13359), .B(new_n13341), .Y(new_n13360));
  nand_5 g11012(.A(new_n13360), .B(new_n13340), .Y(new_n13361));
  nand_5 g11013(.A(new_n13361), .B(new_n13337), .Y(new_n13362));
  nand_5 g11014(.A(new_n13362), .B(new_n13336), .Y(new_n13363));
  nand_5 g11015(.A(new_n13363), .B(new_n13333_1), .Y(new_n13364));
  nand_5 g11016(.A(new_n13364), .B(new_n13332), .Y(new_n13365));
  nand_5 g11017(.A(new_n13365), .B(new_n13329), .Y(new_n13366));
  nand_5 g11018(.A(new_n13366), .B(new_n13328), .Y(new_n13367_1));
  nand_5 g11019(.A(new_n13367_1), .B(new_n13324), .Y(new_n13368));
  nand_5 g11020(.A(new_n13368), .B(new_n13323), .Y(new_n13369));
  nand_5 g11021(.A(new_n13369), .B(new_n13319_1), .Y(new_n13370));
  nand_5 g11022(.A(new_n13370), .B(new_n13318), .Y(new_n13371));
  nand_5 g11023(.A(new_n13371), .B(new_n13284), .Y(new_n13372));
  not_8  g11024(.A(new_n13372), .Y(new_n13373));
  nor_5  g11025(.A(new_n13371), .B(new_n13284), .Y(new_n13374));
  nand_5 g11026(.A(new_n7053), .B(n4514), .Y(new_n13375));
  nand_5 g11027(.A(new_n7054), .B(new_n13219), .Y(new_n13376));
  nand_5 g11028(.A(new_n13376), .B(new_n13375), .Y(new_n13377));
  nand_5 g11029(.A(new_n13316), .B(new_n13285_1), .Y(new_n13378));
  nand_5 g11030(.A(new_n13378), .B(new_n13286), .Y(new_n13379));
  not_8  g11031(.A(new_n13379), .Y(new_n13380));
  xor_4  g11032(.A(new_n13380), .B(new_n13377), .Y(new_n13381));
  nor_5  g11033(.A(new_n13381), .B(new_n13374), .Y(new_n13382));
  nor_5  g11034(.A(new_n13382), .B(new_n13373), .Y(new_n13383));
  nand_5 g11035(.A(new_n13380), .B(new_n13376), .Y(new_n13384));
  not_8  g11036(.A(new_n13384), .Y(new_n13385));
  nand_5 g11037(.A(new_n13375), .B(new_n7052), .Y(new_n13386));
  nor_5  g11038(.A(new_n13386), .B(new_n13385), .Y(new_n13387));
  nor_5  g11039(.A(new_n13387), .B(new_n13383), .Y(new_n13388));
  or_5   g11040(.A(new_n4984), .B(n15766), .Y(new_n13389));
  nand_5 g11041(.A(new_n4984), .B(n15766), .Y(new_n13390));
  or_5   g11042(.A(new_n4989), .B(n25629), .Y(new_n13391));
  nand_5 g11043(.A(new_n4989), .B(n25629), .Y(new_n13392));
  or_5   g11044(.A(new_n4994), .B(n7692), .Y(new_n13393));
  nand_5 g11045(.A(new_n4994), .B(n7692), .Y(new_n13394));
  or_5   g11046(.A(new_n4999), .B(n23039), .Y(new_n13395));
  nand_5 g11047(.A(new_n4999), .B(n23039), .Y(new_n13396));
  nand_5 g11048(.A(new_n4504), .B(new_n4488), .Y(new_n13397));
  nand_5 g11049(.A(new_n13397), .B(new_n4502), .Y(new_n13398));
  nand_5 g11050(.A(new_n13398), .B(new_n13396), .Y(new_n13399));
  nand_5 g11051(.A(new_n13399), .B(new_n13395), .Y(new_n13400));
  nand_5 g11052(.A(new_n13400), .B(new_n13394), .Y(new_n13401));
  nand_5 g11053(.A(new_n13401), .B(new_n13393), .Y(new_n13402));
  nand_5 g11054(.A(new_n13402), .B(new_n13392), .Y(new_n13403));
  nand_5 g11055(.A(new_n13403), .B(new_n13391), .Y(new_n13404));
  nand_5 g11056(.A(new_n13404), .B(new_n13390), .Y(new_n13405));
  nand_5 g11057(.A(new_n13405), .B(new_n13389), .Y(new_n13406));
  nor_5  g11058(.A(new_n13406), .B(new_n4979), .Y(new_n13407_1));
  nand_5 g11059(.A(new_n13407_1), .B(new_n13388), .Y(new_n13408));
  or_5   g11060(.A(new_n13407_1), .B(new_n13388), .Y(new_n13409_1));
  nand_5 g11061(.A(new_n13409_1), .B(new_n13408), .Y(new_n13410));
  not_8  g11062(.A(new_n13407_1), .Y(new_n13411));
  nand_5 g11063(.A(new_n13406), .B(new_n4979), .Y(new_n13412));
  and_5  g11064(.A(new_n13412), .B(new_n13411), .Y(new_n13413));
  xor_4  g11065(.A(new_n13387), .B(new_n13383), .Y(new_n13414));
  or_5   g11066(.A(new_n13414), .B(new_n13413), .Y(new_n13415));
  nand_5 g11067(.A(new_n13414), .B(new_n13413), .Y(new_n13416));
  nor_5  g11068(.A(new_n13374), .B(new_n13373), .Y(new_n13417));
  xor_4  g11069(.A(new_n13417), .B(new_n13381), .Y(new_n13418));
  nand_5 g11070(.A(new_n13389), .B(new_n13390), .Y(new_n13419_1));
  xor_4  g11071(.A(new_n13419_1), .B(new_n13404), .Y(new_n13420));
  not_8  g11072(.A(new_n13420), .Y(new_n13421));
  nand_5 g11073(.A(new_n13421), .B(new_n13418), .Y(new_n13422));
  not_8  g11074(.A(new_n13422), .Y(new_n13423));
  nor_5  g11075(.A(new_n13421), .B(new_n13418), .Y(new_n13424_1));
  nand_5 g11076(.A(new_n13319_1), .B(new_n13318), .Y(new_n13425));
  xor_4  g11077(.A(new_n13425), .B(new_n13369), .Y(new_n13426));
  nand_5 g11078(.A(new_n13391), .B(new_n13392), .Y(new_n13427));
  xor_4  g11079(.A(new_n13427), .B(new_n13402), .Y(new_n13428));
  not_8  g11080(.A(new_n13428), .Y(new_n13429));
  nand_5 g11081(.A(new_n13429), .B(new_n13426), .Y(new_n13430));
  or_5   g11082(.A(new_n13429), .B(new_n13426), .Y(new_n13431));
  nand_5 g11083(.A(new_n13324), .B(new_n13323), .Y(new_n13432));
  xor_4  g11084(.A(new_n13432), .B(new_n13367_1), .Y(new_n13433));
  nand_5 g11085(.A(new_n13393), .B(new_n13394), .Y(new_n13434));
  xor_4  g11086(.A(new_n13434), .B(new_n13400), .Y(new_n13435));
  not_8  g11087(.A(new_n13435), .Y(new_n13436));
  nand_5 g11088(.A(new_n13436), .B(new_n13433), .Y(new_n13437));
  or_5   g11089(.A(new_n13436), .B(new_n13433), .Y(new_n13438));
  nand_5 g11090(.A(new_n13395), .B(new_n13396), .Y(new_n13439));
  xor_4  g11091(.A(new_n13439), .B(new_n13398), .Y(new_n13440));
  not_8  g11092(.A(new_n13440), .Y(new_n13441));
  nand_5 g11093(.A(new_n13329), .B(new_n13328), .Y(new_n13442));
  xor_4  g11094(.A(new_n13442), .B(new_n13365), .Y(new_n13443));
  nand_5 g11095(.A(new_n13443), .B(new_n13441), .Y(new_n13444));
  or_5   g11096(.A(new_n13443), .B(new_n13441), .Y(new_n13445));
  nand_5 g11097(.A(new_n13333_1), .B(new_n13332), .Y(new_n13446));
  xor_4  g11098(.A(new_n13446), .B(new_n13363), .Y(new_n13447));
  nand_5 g11099(.A(new_n13447), .B(new_n4507), .Y(new_n13448));
  or_5   g11100(.A(new_n13447), .B(new_n4507), .Y(new_n13449));
  nand_5 g11101(.A(new_n13337), .B(new_n13336), .Y(new_n13450));
  xor_4  g11102(.A(new_n13450), .B(new_n13361), .Y(new_n13451));
  nand_5 g11103(.A(new_n13451), .B(new_n4375), .Y(new_n13452));
  or_5   g11104(.A(new_n13451), .B(new_n4375), .Y(new_n13453_1));
  nand_5 g11105(.A(new_n13341), .B(new_n13340), .Y(new_n13454));
  xor_4  g11106(.A(new_n13454), .B(new_n13359), .Y(new_n13455));
  nand_5 g11107(.A(new_n13455), .B(new_n4459), .Y(new_n13456_1));
  or_5   g11108(.A(new_n13455), .B(new_n4459), .Y(new_n13457_1));
  nand_5 g11109(.A(new_n13347), .B(new_n13345), .Y(new_n13458));
  xor_4  g11110(.A(new_n13458), .B(new_n13357), .Y(new_n13459));
  nand_5 g11111(.A(new_n13459), .B(new_n4466), .Y(new_n13460_1));
  nor_5  g11112(.A(new_n13459), .B(new_n4466), .Y(new_n13461));
  not_8  g11113(.A(new_n13461), .Y(new_n13462));
  not_8  g11114(.A(new_n4472), .Y(new_n13463));
  nand_5 g11115(.A(new_n13356), .B(new_n13350), .Y(new_n13464));
  xor_4  g11116(.A(new_n13464), .B(new_n13353), .Y(new_n13465));
  nand_5 g11117(.A(new_n13465), .B(new_n13463), .Y(new_n13466));
  nor_5  g11118(.A(new_n13465), .B(new_n13463), .Y(new_n13467));
  not_8  g11119(.A(new_n13467), .Y(new_n13468));
  nand_5 g11120(.A(new_n13352), .B(new_n12547), .Y(new_n13469));
  nand_5 g11121(.A(new_n13469), .B(new_n13353), .Y(new_n13470));
  nand_5 g11122(.A(new_n13470), .B(new_n2635), .Y(new_n13471));
  nand_5 g11123(.A(new_n13471), .B(new_n13468), .Y(new_n13472));
  nand_5 g11124(.A(new_n13472), .B(new_n13466), .Y(new_n13473));
  nand_5 g11125(.A(new_n13473), .B(new_n13462), .Y(new_n13474));
  nand_5 g11126(.A(new_n13474), .B(new_n13460_1), .Y(new_n13475));
  nand_5 g11127(.A(new_n13475), .B(new_n13457_1), .Y(new_n13476));
  nand_5 g11128(.A(new_n13476), .B(new_n13456_1), .Y(new_n13477_1));
  nand_5 g11129(.A(new_n13477_1), .B(new_n13453_1), .Y(new_n13478));
  nand_5 g11130(.A(new_n13478), .B(new_n13452), .Y(new_n13479));
  nand_5 g11131(.A(new_n13479), .B(new_n13449), .Y(new_n13480));
  nand_5 g11132(.A(new_n13480), .B(new_n13448), .Y(new_n13481));
  nand_5 g11133(.A(new_n13481), .B(new_n13445), .Y(new_n13482));
  nand_5 g11134(.A(new_n13482), .B(new_n13444), .Y(new_n13483));
  nand_5 g11135(.A(new_n13483), .B(new_n13438), .Y(new_n13484_1));
  nand_5 g11136(.A(new_n13484_1), .B(new_n13437), .Y(new_n13485));
  nand_5 g11137(.A(new_n13485), .B(new_n13431), .Y(new_n13486_1));
  nand_5 g11138(.A(new_n13486_1), .B(new_n13430), .Y(new_n13487_1));
  not_8  g11139(.A(new_n13487_1), .Y(new_n13488));
  nor_5  g11140(.A(new_n13488), .B(new_n13424_1), .Y(new_n13489));
  nor_5  g11141(.A(new_n13489), .B(new_n13423), .Y(new_n13490_1));
  not_8  g11142(.A(new_n13490_1), .Y(new_n13491));
  nand_5 g11143(.A(new_n13491), .B(new_n13416), .Y(new_n13492));
  nand_5 g11144(.A(new_n13492), .B(new_n13415), .Y(new_n13493));
  not_8  g11145(.A(new_n13493), .Y(new_n13494_1));
  xor_4  g11146(.A(new_n13494_1), .B(new_n13410), .Y(n1701));
  nand_5 g11147(.A(new_n4238), .B(new_n4237), .Y(new_n13496));
  xnor_4 g11148(.A(new_n13496), .B(new_n4274), .Y(n1703));
  nand_5 g11149(.A(new_n5064_1), .B(new_n5062_1), .Y(new_n13498));
  xnor_4 g11150(.A(new_n13498), .B(new_n5127), .Y(n1721));
  nor_5  g11151(.A(new_n10452), .B(new_n10362), .Y(new_n13500_1));
  nor_5  g11152(.A(new_n13500_1), .B(new_n10360), .Y(new_n13501_1));
  nand_5 g11153(.A(new_n8840), .B(new_n4849), .Y(new_n13502));
  nand_5 g11154(.A(new_n10310), .B(new_n13502), .Y(new_n13503));
  nor_5  g11155(.A(new_n13503), .B(new_n10361), .Y(new_n13504));
  nor_5  g11156(.A(new_n13504), .B(new_n13501_1), .Y(new_n13505));
  not_8  g11157(.A(new_n13503), .Y(new_n13506_1));
  nor_5  g11158(.A(new_n13506_1), .B(new_n10359), .Y(new_n13507));
  nor_5  g11159(.A(new_n13507), .B(new_n13500_1), .Y(new_n13508));
  nor_5  g11160(.A(new_n13508), .B(new_n13505), .Y(n1760));
  nand_5 g11161(.A(new_n4470), .B(new_n4469), .Y(new_n13510));
  xnor_4 g11162(.A(new_n13510), .B(new_n4479), .Y(n1791));
  xor_4  g11163(.A(new_n3658), .B(new_n3656), .Y(n1808));
  nand_5 g11164(.A(new_n6233_1), .B(n4319), .Y(new_n13513));
  nand_5 g11165(.A(n13494), .B(new_n3313), .Y(new_n13514));
  nand_5 g11166(.A(new_n12951), .B(new_n12949), .Y(new_n13515));
  nand_5 g11167(.A(new_n13515), .B(new_n12950), .Y(new_n13516));
  nand_5 g11168(.A(new_n13516), .B(new_n13514), .Y(new_n13517));
  nand_5 g11169(.A(new_n13517), .B(new_n13513), .Y(new_n13518));
  nor_5  g11170(.A(new_n13518), .B(new_n8942), .Y(new_n13519));
  and_5  g11171(.A(new_n13518), .B(new_n8942), .Y(new_n13520));
  nand_5 g11172(.A(new_n13514), .B(new_n13513), .Y(new_n13521));
  xor_4  g11173(.A(new_n13521), .B(new_n13516), .Y(new_n13522));
  or_5   g11174(.A(new_n13522), .B(new_n9016), .Y(new_n13523));
  nand_5 g11175(.A(new_n13522), .B(new_n9016), .Y(new_n13524));
  nand_5 g11176(.A(new_n12955), .B(new_n12947), .Y(new_n13525));
  nand_5 g11177(.A(new_n13525), .B(new_n12954), .Y(new_n13526));
  nand_5 g11178(.A(new_n13526), .B(new_n13524), .Y(new_n13527));
  and_5  g11179(.A(new_n13527), .B(new_n13523), .Y(new_n13528));
  nor_5  g11180(.A(new_n13528), .B(new_n13520), .Y(new_n13529));
  nor_5  g11181(.A(new_n13529), .B(new_n13519), .Y(new_n13530));
  nand_5 g11182(.A(new_n8940), .B(new_n8842), .Y(new_n13531));
  and_5  g11183(.A(new_n13531), .B(new_n13518), .Y(new_n13532));
  nor_5  g11184(.A(new_n13532), .B(new_n13530), .Y(new_n13533));
  nor_5  g11185(.A(new_n13531), .B(new_n13518), .Y(new_n13534));
  nor_5  g11186(.A(new_n13534), .B(new_n13529), .Y(new_n13535));
  nor_5  g11187(.A(new_n13535), .B(new_n13533), .Y(n1821));
  not_8  g11188(.A(new_n7935), .Y(new_n13537));
  xor_4  g11189(.A(new_n7937_1), .B(new_n13537), .Y(n1832));
  nand_5 g11190(.A(new_n4139), .B(new_n6807), .Y(new_n13539));
  nor_5  g11191(.A(new_n13539), .B(n11926), .Y(new_n13540));
  nand_5 g11192(.A(new_n13540), .B(new_n6800), .Y(new_n13541));
  nor_5  g11193(.A(new_n13541), .B(n21784), .Y(new_n13542));
  not_8  g11194(.A(new_n13542), .Y(new_n13543));
  nand_5 g11195(.A(new_n13541), .B(n21784), .Y(new_n13544));
  and_5  g11196(.A(new_n13544), .B(new_n13543), .Y(new_n13545));
  nand_5 g11197(.A(new_n13545), .B(new_n8361), .Y(new_n13546));
  or_5   g11198(.A(new_n13545), .B(new_n8361), .Y(new_n13547));
  nand_5 g11199(.A(new_n13547), .B(new_n13546), .Y(new_n13548_1));
  xor_4  g11200(.A(new_n13540), .B(n5521), .Y(new_n13549_1));
  nand_5 g11201(.A(new_n13549_1), .B(new_n8366), .Y(new_n13550));
  not_8  g11202(.A(new_n13550), .Y(new_n13551_1));
  nor_5  g11203(.A(new_n13549_1), .B(new_n8366), .Y(new_n13552));
  xor_4  g11204(.A(new_n13539), .B(new_n6804), .Y(new_n13553));
  nand_5 g11205(.A(new_n13553), .B(new_n8372), .Y(new_n13554));
  not_8  g11206(.A(new_n13554), .Y(new_n13555));
  nor_5  g11207(.A(new_n13553), .B(new_n8372), .Y(new_n13556));
  nand_5 g11208(.A(new_n4287), .B(new_n4278), .Y(new_n13557));
  and_5  g11209(.A(new_n13557), .B(new_n4288), .Y(new_n13558));
  nor_5  g11210(.A(new_n13558), .B(new_n13556), .Y(new_n13559));
  nor_5  g11211(.A(new_n13559), .B(new_n13555), .Y(new_n13560));
  nor_5  g11212(.A(new_n13560), .B(new_n13552), .Y(new_n13561));
  nor_5  g11213(.A(new_n13561), .B(new_n13551_1), .Y(new_n13562));
  not_8  g11214(.A(new_n13562), .Y(new_n13563));
  xor_4  g11215(.A(new_n13563), .B(new_n13548_1), .Y(new_n13564));
  not_8  g11216(.A(n2160), .Y(new_n13565));
  nand_5 g11217(.A(n9934), .B(n2272), .Y(new_n13566));
  nand_5 g11218(.A(new_n5326), .B(new_n8142), .Y(new_n13567));
  nand_5 g11219(.A(new_n13567), .B(new_n13566), .Y(new_n13568));
  nand_5 g11220(.A(new_n8146), .B(new_n5363), .Y(new_n13569));
  nand_5 g11221(.A(n25331), .B(n18496), .Y(new_n13570));
  nand_5 g11222(.A(new_n5588), .B(new_n8150), .Y(new_n13571));
  nand_5 g11223(.A(n26224), .B(n18483), .Y(new_n13572));
  nand_5 g11224(.A(new_n8153), .B(new_n4297), .Y(new_n13573));
  nand_5 g11225(.A(n21934), .B(n19327), .Y(new_n13574));
  nand_5 g11226(.A(new_n4222), .B(new_n8156), .Y(new_n13575));
  nand_5 g11227(.A(n22597), .B(n18901), .Y(new_n13576));
  nand_5 g11228(.A(new_n4177), .B(new_n8159_1), .Y(new_n13577));
  nand_5 g11229(.A(n26107), .B(n4376), .Y(new_n13578));
  nand_5 g11230(.A(new_n8162), .B(new_n4146_1), .Y(new_n13579));
  nand_5 g11231(.A(n14570), .B(n342), .Y(new_n13580));
  nand_5 g11232(.A(new_n4160), .B(new_n8165), .Y(new_n13581));
  nand_5 g11233(.A(n26553), .B(n23775), .Y(new_n13582));
  nand_5 g11234(.A(new_n8168), .B(new_n5331), .Y(new_n13583));
  nand_5 g11235(.A(n8259), .B(n4964), .Y(new_n13584));
  nand_5 g11236(.A(n11479), .B(n7876), .Y(new_n13585));
  nand_5 g11237(.A(new_n13585), .B(new_n13584), .Y(new_n13586));
  nand_5 g11238(.A(new_n13586), .B(new_n13583), .Y(new_n13587));
  nand_5 g11239(.A(new_n13587), .B(new_n13582), .Y(new_n13588));
  nand_5 g11240(.A(new_n13588), .B(new_n13581), .Y(new_n13589));
  nand_5 g11241(.A(new_n13589), .B(new_n13580), .Y(new_n13590));
  nand_5 g11242(.A(new_n13590), .B(new_n13579), .Y(new_n13591));
  nand_5 g11243(.A(new_n13591), .B(new_n13578), .Y(new_n13592));
  nand_5 g11244(.A(new_n13592), .B(new_n13577), .Y(new_n13593));
  nand_5 g11245(.A(new_n13593), .B(new_n13576), .Y(new_n13594));
  nand_5 g11246(.A(new_n13594), .B(new_n13575), .Y(new_n13595));
  nand_5 g11247(.A(new_n13595), .B(new_n13574), .Y(new_n13596));
  nand_5 g11248(.A(new_n13596), .B(new_n13573), .Y(new_n13597));
  nand_5 g11249(.A(new_n13597), .B(new_n13572), .Y(new_n13598));
  nand_5 g11250(.A(new_n13598), .B(new_n13571), .Y(new_n13599));
  nand_5 g11251(.A(new_n13599), .B(new_n13570), .Y(new_n13600));
  nand_5 g11252(.A(new_n13600), .B(new_n13569), .Y(new_n13601));
  not_8  g11253(.A(new_n13601), .Y(new_n13602_1));
  xor_4  g11254(.A(new_n13602_1), .B(new_n13568), .Y(new_n13603));
  not_8  g11255(.A(new_n13603), .Y(new_n13604));
  nand_5 g11256(.A(new_n13604), .B(new_n13565), .Y(new_n13605));
  nand_5 g11257(.A(new_n13603), .B(n2160), .Y(new_n13606));
  nand_5 g11258(.A(new_n13606), .B(new_n13605), .Y(new_n13607));
  nand_5 g11259(.A(new_n13570), .B(new_n13569), .Y(new_n13608));
  xor_4  g11260(.A(new_n13608), .B(new_n13599), .Y(new_n13609));
  nand_5 g11261(.A(new_n13609), .B(new_n3287), .Y(new_n13610));
  not_8  g11262(.A(new_n13610), .Y(new_n13611));
  nor_5  g11263(.A(new_n13609), .B(new_n3287), .Y(new_n13612));
  nand_5 g11264(.A(new_n13572), .B(new_n13571), .Y(new_n13613));
  xor_4  g11265(.A(new_n13613), .B(new_n13597), .Y(new_n13614));
  nand_5 g11266(.A(new_n13614), .B(new_n3185), .Y(new_n13615));
  or_5   g11267(.A(new_n13614), .B(new_n3185), .Y(new_n13616));
  nand_5 g11268(.A(new_n13574), .B(new_n13573), .Y(new_n13617));
  xor_4  g11269(.A(new_n13617), .B(new_n13595), .Y(new_n13618));
  nand_5 g11270(.A(new_n13618), .B(new_n3067_1), .Y(new_n13619));
  or_5   g11271(.A(new_n13618), .B(new_n3067_1), .Y(new_n13620));
  nand_5 g11272(.A(new_n13576), .B(new_n13575), .Y(new_n13621));
  xor_4  g11273(.A(new_n13621), .B(new_n13593), .Y(new_n13622));
  nand_5 g11274(.A(new_n13622), .B(new_n3034), .Y(new_n13623));
  nor_5  g11275(.A(new_n13622), .B(new_n3034), .Y(new_n13624));
  not_8  g11276(.A(new_n13624), .Y(new_n13625));
  nand_5 g11277(.A(new_n13578), .B(new_n13577), .Y(new_n13626_1));
  xor_4  g11278(.A(new_n13626_1), .B(new_n13591), .Y(new_n13627));
  nand_5 g11279(.A(new_n13627), .B(new_n3039), .Y(new_n13628));
  nor_5  g11280(.A(new_n13627), .B(new_n3039), .Y(new_n13629));
  not_8  g11281(.A(new_n13629), .Y(new_n13630));
  nand_5 g11282(.A(new_n13580), .B(new_n13579), .Y(new_n13631));
  xor_4  g11283(.A(new_n13631), .B(new_n13589), .Y(new_n13632));
  nand_5 g11284(.A(new_n13632), .B(new_n3042), .Y(new_n13633));
  nor_5  g11285(.A(new_n13632), .B(new_n3042), .Y(new_n13634));
  not_8  g11286(.A(new_n13634), .Y(new_n13635));
  nand_5 g11287(.A(new_n13582), .B(new_n13581), .Y(new_n13636));
  xor_4  g11288(.A(new_n13636), .B(new_n13587), .Y(new_n13637));
  nand_5 g11289(.A(new_n13637), .B(new_n3047), .Y(new_n13638));
  nor_5  g11290(.A(new_n13637), .B(new_n3047), .Y(new_n13639));
  nand_5 g11291(.A(new_n8170), .B(new_n4207), .Y(new_n13640));
  and_5  g11292(.A(new_n13640), .B(new_n13585), .Y(new_n13641));
  or_5   g11293(.A(new_n13641), .B(new_n3158), .Y(new_n13642));
  nor_5  g11294(.A(new_n13642), .B(new_n3050), .Y(new_n13643));
  not_8  g11295(.A(new_n13643), .Y(new_n13644));
  nand_5 g11296(.A(new_n13642), .B(new_n3050), .Y(new_n13645));
  nand_5 g11297(.A(new_n13584), .B(new_n13583), .Y(new_n13646));
  xor_4  g11298(.A(new_n13646), .B(new_n13585), .Y(new_n13647));
  not_8  g11299(.A(new_n13647), .Y(new_n13648));
  nand_5 g11300(.A(new_n13648), .B(new_n13645), .Y(new_n13649));
  nand_5 g11301(.A(new_n13649), .B(new_n13644), .Y(new_n13650));
  or_5   g11302(.A(new_n13650), .B(new_n13639), .Y(new_n13651));
  nand_5 g11303(.A(new_n13651), .B(new_n13638), .Y(new_n13652));
  nand_5 g11304(.A(new_n13652), .B(new_n13635), .Y(new_n13653));
  nand_5 g11305(.A(new_n13653), .B(new_n13633), .Y(new_n13654));
  nand_5 g11306(.A(new_n13654), .B(new_n13630), .Y(new_n13655));
  nand_5 g11307(.A(new_n13655), .B(new_n13628), .Y(new_n13656));
  nand_5 g11308(.A(new_n13656), .B(new_n13625), .Y(new_n13657));
  nand_5 g11309(.A(new_n13657), .B(new_n13623), .Y(new_n13658));
  nand_5 g11310(.A(new_n13658), .B(new_n13620), .Y(new_n13659));
  nand_5 g11311(.A(new_n13659), .B(new_n13619), .Y(new_n13660));
  nand_5 g11312(.A(new_n13660), .B(new_n13616), .Y(new_n13661));
  nand_5 g11313(.A(new_n13661), .B(new_n13615), .Y(new_n13662));
  not_8  g11314(.A(new_n13662), .Y(new_n13663));
  nor_5  g11315(.A(new_n13663), .B(new_n13612), .Y(new_n13664));
  nor_5  g11316(.A(new_n13664), .B(new_n13611), .Y(new_n13665));
  xor_4  g11317(.A(new_n13665), .B(new_n13607), .Y(new_n13666));
  nand_5 g11318(.A(new_n13666), .B(new_n13564), .Y(new_n13667));
  or_5   g11319(.A(new_n13666), .B(new_n13564), .Y(new_n13668_1));
  nand_5 g11320(.A(new_n13668_1), .B(new_n13667), .Y(new_n13669));
  nor_5  g11321(.A(new_n13552), .B(new_n13551_1), .Y(new_n13670));
  xor_4  g11322(.A(new_n13670), .B(new_n13560), .Y(new_n13671));
  nor_5  g11323(.A(new_n13612), .B(new_n13611), .Y(new_n13672));
  xor_4  g11324(.A(new_n13672), .B(new_n13662), .Y(new_n13673));
  nand_5 g11325(.A(new_n13673), .B(new_n13671), .Y(new_n13674));
  nor_5  g11326(.A(new_n13673), .B(new_n13671), .Y(new_n13675));
  not_8  g11327(.A(new_n13675), .Y(new_n13676));
  nor_5  g11328(.A(new_n13556), .B(new_n13555), .Y(new_n13677_1));
  xor_4  g11329(.A(new_n13677_1), .B(new_n13558), .Y(new_n13678));
  not_8  g11330(.A(new_n13678), .Y(new_n13679));
  nand_5 g11331(.A(new_n13616), .B(new_n13615), .Y(new_n13680));
  xor_4  g11332(.A(new_n13680), .B(new_n13660), .Y(new_n13681));
  or_5   g11333(.A(new_n13681), .B(new_n13679), .Y(new_n13682));
  nand_5 g11334(.A(new_n13681), .B(new_n13679), .Y(new_n13683_1));
  nand_5 g11335(.A(new_n13620), .B(new_n13619), .Y(new_n13684));
  xor_4  g11336(.A(new_n13684), .B(new_n13658), .Y(new_n13685));
  not_8  g11337(.A(new_n13685), .Y(new_n13686));
  nand_5 g11338(.A(new_n13686), .B(new_n4290), .Y(new_n13687));
  not_8  g11339(.A(new_n13687), .Y(new_n13688));
  nor_5  g11340(.A(new_n13686), .B(new_n4290), .Y(new_n13689));
  nand_5 g11341(.A(new_n13625), .B(new_n13623), .Y(new_n13690));
  xor_4  g11342(.A(new_n13690), .B(new_n13656), .Y(new_n13691));
  not_8  g11343(.A(new_n13691), .Y(new_n13692));
  nand_5 g11344(.A(new_n13692), .B(new_n4145), .Y(new_n13693));
  nor_5  g11345(.A(new_n13692), .B(new_n4145), .Y(new_n13694));
  not_8  g11346(.A(new_n13694), .Y(new_n13695));
  not_8  g11347(.A(new_n4240), .Y(new_n13696));
  nand_5 g11348(.A(new_n13630), .B(new_n13628), .Y(new_n13697));
  xor_4  g11349(.A(new_n13697), .B(new_n13654), .Y(new_n13698));
  or_5   g11350(.A(new_n13698), .B(new_n13696), .Y(new_n13699));
  nand_5 g11351(.A(new_n13698), .B(new_n13696), .Y(new_n13700));
  nand_5 g11352(.A(new_n13635), .B(new_n13633), .Y(new_n13701));
  xor_4  g11353(.A(new_n13701), .B(new_n13652), .Y(new_n13702));
  not_8  g11354(.A(new_n13702), .Y(new_n13703));
  nand_5 g11355(.A(new_n13703), .B(new_n4246), .Y(new_n13704));
  nor_5  g11356(.A(new_n13703), .B(new_n4246), .Y(new_n13705));
  not_8  g11357(.A(new_n13639), .Y(new_n13706));
  nand_5 g11358(.A(new_n13706), .B(new_n13638), .Y(new_n13707));
  xor_4  g11359(.A(new_n13707), .B(new_n13650), .Y(new_n13708_1));
  nand_5 g11360(.A(new_n13708_1), .B(new_n4252), .Y(new_n13709));
  not_8  g11361(.A(new_n13709), .Y(new_n13710_1));
  nor_5  g11362(.A(new_n13708_1), .B(new_n4252), .Y(new_n13711));
  not_8  g11363(.A(new_n4264), .Y(new_n13712));
  xor_4  g11364(.A(new_n13641), .B(new_n3158), .Y(new_n13713));
  nor_5  g11365(.A(new_n13713), .B(new_n13712), .Y(new_n13714_1));
  nand_5 g11366(.A(new_n13644), .B(new_n13645), .Y(new_n13715));
  xor_4  g11367(.A(new_n13715), .B(new_n13648), .Y(new_n13716));
  nand_5 g11368(.A(new_n13716), .B(new_n13714_1), .Y(new_n13717));
  or_5   g11369(.A(new_n13716), .B(new_n13714_1), .Y(new_n13718));
  nand_5 g11370(.A(new_n13718), .B(new_n4258), .Y(new_n13719_1));
  nand_5 g11371(.A(new_n13719_1), .B(new_n13717), .Y(new_n13720));
  not_8  g11372(.A(new_n13720), .Y(new_n13721));
  nor_5  g11373(.A(new_n13721), .B(new_n13711), .Y(new_n13722_1));
  nor_5  g11374(.A(new_n13722_1), .B(new_n13710_1), .Y(new_n13723));
  or_5   g11375(.A(new_n13723), .B(new_n13705), .Y(new_n13724));
  nand_5 g11376(.A(new_n13724), .B(new_n13704), .Y(new_n13725));
  nand_5 g11377(.A(new_n13725), .B(new_n13700), .Y(new_n13726));
  nand_5 g11378(.A(new_n13726), .B(new_n13699), .Y(new_n13727));
  nand_5 g11379(.A(new_n13727), .B(new_n13695), .Y(new_n13728));
  nand_5 g11380(.A(new_n13728), .B(new_n13693), .Y(new_n13729));
  not_8  g11381(.A(new_n13729), .Y(new_n13730));
  nor_5  g11382(.A(new_n13730), .B(new_n13689), .Y(new_n13731));
  nor_5  g11383(.A(new_n13731), .B(new_n13688), .Y(new_n13732));
  not_8  g11384(.A(new_n13732), .Y(new_n13733));
  nand_5 g11385(.A(new_n13733), .B(new_n13683_1), .Y(new_n13734));
  nand_5 g11386(.A(new_n13734), .B(new_n13682), .Y(new_n13735));
  nand_5 g11387(.A(new_n13735), .B(new_n13676), .Y(new_n13736));
  nand_5 g11388(.A(new_n13736), .B(new_n13674), .Y(new_n13737));
  not_8  g11389(.A(new_n13737), .Y(new_n13738));
  xor_4  g11390(.A(new_n13738), .B(new_n13669), .Y(n1859));
  nor_5  g11391(.A(new_n5826), .B(new_n5825), .Y(new_n13740));
  xor_4  g11392(.A(new_n13740), .B(new_n5856), .Y(n1860));
  nand_5 g11393(.A(new_n7976), .B(new_n7972), .Y(new_n13742));
  nand_5 g11394(.A(new_n13742), .B(new_n7975), .Y(new_n13743));
  nand_5 g11395(.A(new_n13743), .B(new_n6382), .Y(new_n13744));
  not_8  g11396(.A(new_n13744), .Y(new_n13745));
  nor_5  g11397(.A(new_n13743), .B(new_n6382), .Y(new_n13746));
  nor_5  g11398(.A(new_n13746), .B(n25972), .Y(new_n13747));
  nor_5  g11399(.A(new_n13747), .B(new_n13745), .Y(new_n13748));
  nor_5  g11400(.A(new_n13746), .B(new_n13745), .Y(new_n13749));
  xor_4  g11401(.A(new_n13749), .B(new_n9943), .Y(new_n13750));
  not_8  g11402(.A(new_n13750), .Y(new_n13751));
  nand_5 g11403(.A(new_n13751), .B(n10250), .Y(new_n13752));
  nand_5 g11404(.A(new_n13750), .B(new_n7040), .Y(new_n13753));
  nand_5 g11405(.A(new_n7979), .B(n7674), .Y(new_n13754_1));
  nand_5 g11406(.A(new_n7978), .B(new_n6991), .Y(new_n13755));
  nand_5 g11407(.A(new_n7886), .B(n6397), .Y(new_n13756));
  nand_5 g11408(.A(new_n7885), .B(new_n6997), .Y(new_n13757));
  nand_5 g11409(.A(new_n7842), .B(n19196), .Y(new_n13758));
  nand_5 g11410(.A(new_n7841_1), .B(new_n7003), .Y(new_n13759));
  nand_5 g11411(.A(new_n7846), .B(n23586), .Y(new_n13760));
  nand_5 g11412(.A(new_n7848), .B(new_n7118), .Y(new_n13761));
  nand_5 g11413(.A(new_n7851), .B(n21226), .Y(new_n13762));
  nand_5 g11414(.A(new_n7853), .B(new_n7009), .Y(new_n13763));
  nand_5 g11415(.A(new_n7856), .B(n4426), .Y(new_n13764_1));
  nand_5 g11416(.A(new_n7858), .B(new_n7012), .Y(new_n13765));
  nand_5 g11417(.A(new_n4612), .B(n20036), .Y(new_n13766));
  nand_5 g11418(.A(new_n4600), .B(new_n4606), .Y(new_n13767));
  nand_5 g11419(.A(new_n4566), .B(n11192), .Y(new_n13768));
  nand_5 g11420(.A(new_n4557), .B(new_n4561), .Y(new_n13769));
  nand_5 g11421(.A(new_n4544), .B(n9380), .Y(new_n13770));
  not_8  g11422(.A(new_n13770), .Y(new_n13771));
  nand_5 g11423(.A(new_n13771), .B(new_n13769), .Y(new_n13772));
  nand_5 g11424(.A(new_n13772), .B(new_n13768), .Y(new_n13773));
  nand_5 g11425(.A(new_n13773), .B(new_n13767), .Y(new_n13774));
  nand_5 g11426(.A(new_n13774), .B(new_n13766), .Y(new_n13775_1));
  nand_5 g11427(.A(new_n13775_1), .B(new_n13765), .Y(new_n13776));
  nand_5 g11428(.A(new_n13776), .B(new_n13764_1), .Y(new_n13777));
  nand_5 g11429(.A(new_n13777), .B(new_n13763), .Y(new_n13778));
  nand_5 g11430(.A(new_n13778), .B(new_n13762), .Y(new_n13779));
  nand_5 g11431(.A(new_n13779), .B(new_n13761), .Y(new_n13780));
  nand_5 g11432(.A(new_n13780), .B(new_n13760), .Y(new_n13781_1));
  nand_5 g11433(.A(new_n13781_1), .B(new_n13759), .Y(new_n13782));
  nand_5 g11434(.A(new_n13782), .B(new_n13758), .Y(new_n13783_1));
  nand_5 g11435(.A(new_n13783_1), .B(new_n13757), .Y(new_n13784));
  nand_5 g11436(.A(new_n13784), .B(new_n13756), .Y(new_n13785));
  nand_5 g11437(.A(new_n13785), .B(new_n13755), .Y(new_n13786));
  nand_5 g11438(.A(new_n13786), .B(new_n13754_1), .Y(new_n13787));
  nand_5 g11439(.A(new_n13787), .B(new_n13753), .Y(new_n13788));
  nand_5 g11440(.A(new_n13788), .B(new_n13752), .Y(new_n13789));
  nand_5 g11441(.A(new_n13789), .B(new_n13748), .Y(new_n13790));
  nand_5 g11442(.A(new_n13790), .B(new_n13162), .Y(new_n13791));
  or_5   g11443(.A(new_n13790), .B(new_n13162), .Y(new_n13792));
  not_8  g11444(.A(new_n13165), .Y(new_n13793));
  xor_4  g11445(.A(new_n13789), .B(new_n13748), .Y(new_n13794));
  or_5   g11446(.A(new_n13794), .B(new_n13793), .Y(new_n13795));
  nand_5 g11447(.A(new_n13794), .B(new_n13793), .Y(new_n13796));
  nand_5 g11448(.A(new_n13752), .B(new_n13753), .Y(new_n13797));
  xor_4  g11449(.A(new_n13797), .B(new_n13787), .Y(new_n13798_1));
  nand_5 g11450(.A(new_n13798_1), .B(new_n13175), .Y(new_n13799));
  or_5   g11451(.A(new_n13798_1), .B(new_n13175), .Y(new_n13800));
  nand_5 g11452(.A(new_n13754_1), .B(new_n13755), .Y(new_n13801));
  xor_4  g11453(.A(new_n13801), .B(new_n13785), .Y(new_n13802));
  nand_5 g11454(.A(new_n13802), .B(new_n13183), .Y(new_n13803));
  or_5   g11455(.A(new_n13802), .B(new_n13183), .Y(new_n13804));
  nand_5 g11456(.A(new_n13756), .B(new_n13757), .Y(new_n13805));
  xor_4  g11457(.A(new_n13805), .B(new_n13783_1), .Y(new_n13806));
  nand_5 g11458(.A(new_n13806), .B(new_n13189), .Y(new_n13807));
  or_5   g11459(.A(new_n13806), .B(new_n13189), .Y(new_n13808));
  nand_5 g11460(.A(new_n13758), .B(new_n13759), .Y(new_n13809));
  xor_4  g11461(.A(new_n13809), .B(new_n13781_1), .Y(new_n13810));
  nand_5 g11462(.A(new_n13810), .B(new_n13196), .Y(new_n13811));
  or_5   g11463(.A(new_n13810), .B(new_n13196), .Y(new_n13812));
  nand_5 g11464(.A(new_n13760), .B(new_n13761), .Y(new_n13813));
  xor_4  g11465(.A(new_n13813), .B(new_n13779), .Y(new_n13814));
  nand_5 g11466(.A(new_n13814), .B(new_n13202), .Y(new_n13815));
  or_5   g11467(.A(new_n13814), .B(new_n13202), .Y(new_n13816));
  nand_5 g11468(.A(new_n13762), .B(new_n13763), .Y(new_n13817));
  xor_4  g11469(.A(new_n13817), .B(new_n13777), .Y(new_n13818));
  nand_5 g11470(.A(new_n13818), .B(new_n11078_1), .Y(new_n13819));
  or_5   g11471(.A(new_n13818), .B(new_n11078_1), .Y(new_n13820));
  nand_5 g11472(.A(new_n13764_1), .B(new_n13765), .Y(new_n13821));
  xor_4  g11473(.A(new_n13821), .B(new_n13775_1), .Y(new_n13822));
  nand_5 g11474(.A(new_n13822), .B(new_n11026), .Y(new_n13823));
  or_5   g11475(.A(new_n13822), .B(new_n11026), .Y(new_n13824));
  nand_5 g11476(.A(new_n13766), .B(new_n13767), .Y(new_n13825));
  xor_4  g11477(.A(new_n13825), .B(new_n13773), .Y(new_n13826));
  nand_5 g11478(.A(new_n13826), .B(new_n10995), .Y(new_n13827));
  or_5   g11479(.A(new_n13826), .B(new_n10995), .Y(new_n13828));
  nand_5 g11480(.A(new_n13768), .B(new_n13769), .Y(new_n13829));
  xor_4  g11481(.A(new_n13829), .B(new_n13771), .Y(new_n13830));
  nand_5 g11482(.A(new_n13830), .B(new_n11011_1), .Y(new_n13831));
  or_5   g11483(.A(new_n13830), .B(new_n11011_1), .Y(new_n13832));
  nor_5  g11484(.A(new_n4544), .B(n9380), .Y(new_n13833));
  nor_5  g11485(.A(new_n13833), .B(new_n13771), .Y(new_n13834));
  nor_5  g11486(.A(new_n13834), .B(new_n8285_1), .Y(new_n13835_1));
  nand_5 g11487(.A(new_n13835_1), .B(new_n13832), .Y(new_n13836));
  nand_5 g11488(.A(new_n13836), .B(new_n13831), .Y(new_n13837));
  nand_5 g11489(.A(new_n13837), .B(new_n13828), .Y(new_n13838));
  nand_5 g11490(.A(new_n13838), .B(new_n13827), .Y(new_n13839));
  nand_5 g11491(.A(new_n13839), .B(new_n13824), .Y(new_n13840));
  nand_5 g11492(.A(new_n13840), .B(new_n13823), .Y(new_n13841));
  nand_5 g11493(.A(new_n13841), .B(new_n13820), .Y(new_n13842));
  nand_5 g11494(.A(new_n13842), .B(new_n13819), .Y(new_n13843));
  nand_5 g11495(.A(new_n13843), .B(new_n13816), .Y(new_n13844));
  nand_5 g11496(.A(new_n13844), .B(new_n13815), .Y(new_n13845));
  nand_5 g11497(.A(new_n13845), .B(new_n13812), .Y(new_n13846));
  nand_5 g11498(.A(new_n13846), .B(new_n13811), .Y(new_n13847));
  nand_5 g11499(.A(new_n13847), .B(new_n13808), .Y(new_n13848));
  nand_5 g11500(.A(new_n13848), .B(new_n13807), .Y(new_n13849));
  nand_5 g11501(.A(new_n13849), .B(new_n13804), .Y(new_n13850_1));
  nand_5 g11502(.A(new_n13850_1), .B(new_n13803), .Y(new_n13851_1));
  nand_5 g11503(.A(new_n13851_1), .B(new_n13800), .Y(new_n13852));
  nand_5 g11504(.A(new_n13852), .B(new_n13799), .Y(new_n13853));
  nand_5 g11505(.A(new_n13853), .B(new_n13796), .Y(new_n13854));
  nand_5 g11506(.A(new_n13854), .B(new_n13795), .Y(new_n13855));
  nand_5 g11507(.A(new_n13855), .B(new_n13792), .Y(new_n13856));
  nand_5 g11508(.A(new_n13856), .B(new_n13791), .Y(n1861));
  nand_5 g11509(.A(new_n10138), .B(new_n11723), .Y(new_n13858));
  not_8  g11510(.A(new_n13858), .Y(new_n13859));
  nand_5 g11511(.A(new_n13859), .B(new_n11720), .Y(new_n13860));
  nor_5  g11512(.A(new_n13860), .B(n8309), .Y(new_n13861));
  nand_5 g11513(.A(new_n13861), .B(new_n11713), .Y(new_n13862));
  not_8  g11514(.A(new_n13862), .Y(new_n13863));
  nor_5  g11515(.A(new_n13861), .B(new_n11713), .Y(new_n13864));
  nor_5  g11516(.A(new_n13864), .B(new_n13863), .Y(new_n13865));
  nand_5 g11517(.A(new_n13865), .B(new_n6045), .Y(new_n13866));
  or_5   g11518(.A(new_n13865), .B(new_n6045), .Y(new_n13867));
  xor_4  g11519(.A(new_n13860), .B(new_n11716), .Y(new_n13868));
  or_5   g11520(.A(new_n13868), .B(new_n6012_1), .Y(new_n13869));
  nand_5 g11521(.A(new_n13868), .B(new_n6012_1), .Y(new_n13870));
  nand_5 g11522(.A(new_n13858), .B(n19144), .Y(new_n13871));
  nand_5 g11523(.A(new_n13871), .B(new_n13860), .Y(new_n13872));
  or_5   g11524(.A(new_n13872), .B(new_n6019), .Y(new_n13873));
  nand_5 g11525(.A(new_n13872), .B(new_n6019), .Y(new_n13874));
  nand_5 g11526(.A(new_n6030), .B(n13714), .Y(new_n13875));
  nand_5 g11527(.A(n13714), .B(n12593), .Y(new_n13876));
  nand_5 g11528(.A(new_n13876), .B(new_n13858), .Y(new_n13877));
  nand_5 g11529(.A(new_n13877), .B(new_n13875), .Y(new_n13878));
  not_8  g11530(.A(new_n13878), .Y(new_n13879));
  nor_5  g11531(.A(new_n13875), .B(n12593), .Y(new_n13880));
  nor_5  g11532(.A(new_n13880), .B(new_n6023), .Y(new_n13881));
  nor_5  g11533(.A(new_n13881), .B(new_n13879), .Y(new_n13882));
  nand_5 g11534(.A(new_n13882), .B(new_n13874), .Y(new_n13883));
  nand_5 g11535(.A(new_n13883), .B(new_n13873), .Y(new_n13884));
  nand_5 g11536(.A(new_n13884), .B(new_n13870), .Y(new_n13885));
  nand_5 g11537(.A(new_n13885), .B(new_n13869), .Y(new_n13886));
  nand_5 g11538(.A(new_n13886), .B(new_n13867), .Y(new_n13887));
  nand_5 g11539(.A(new_n13887), .B(new_n13866), .Y(new_n13888));
  nand_5 g11540(.A(new_n13863), .B(new_n11710_1), .Y(new_n13889));
  not_8  g11541(.A(new_n13889), .Y(new_n13890));
  nor_5  g11542(.A(new_n13863), .B(new_n11710_1), .Y(new_n13891));
  nor_5  g11543(.A(new_n13891), .B(new_n13890), .Y(new_n13892));
  nand_5 g11544(.A(new_n13892), .B(new_n5997), .Y(new_n13893));
  or_5   g11545(.A(new_n13892), .B(new_n5997), .Y(new_n13894));
  nand_5 g11546(.A(new_n13894), .B(new_n13893), .Y(new_n13895));
  xor_4  g11547(.A(new_n13895), .B(new_n13888), .Y(new_n13896));
  nand_5 g11548(.A(new_n9930), .B(new_n8386), .Y(new_n13897));
  nand_5 g11549(.A(new_n9929), .B(new_n8388), .Y(new_n13898));
  nand_5 g11550(.A(new_n9887), .B(new_n8391), .Y(new_n13899));
  not_8  g11551(.A(new_n8391), .Y(new_n13900));
  nand_5 g11552(.A(new_n9886), .B(new_n13900), .Y(new_n13901));
  nand_5 g11553(.A(new_n9856), .B(new_n8396), .Y(new_n13902));
  nand_5 g11554(.A(new_n9855), .B(new_n8398), .Y(new_n13903));
  nand_5 g11555(.A(new_n9846), .B(new_n8402), .Y(new_n13904));
  nand_5 g11556(.A(new_n9845), .B(new_n8401), .Y(new_n13905));
  nand_5 g11557(.A(new_n8407), .B(n18962), .Y(new_n13906));
  nand_5 g11558(.A(new_n13906), .B(new_n13905), .Y(new_n13907));
  nand_5 g11559(.A(new_n13907), .B(new_n13904), .Y(new_n13908));
  nand_5 g11560(.A(new_n13908), .B(new_n13903), .Y(new_n13909));
  nand_5 g11561(.A(new_n13909), .B(new_n13902), .Y(new_n13910));
  nand_5 g11562(.A(new_n13910), .B(new_n13901), .Y(new_n13911));
  nand_5 g11563(.A(new_n13911), .B(new_n13899), .Y(new_n13912_1));
  nand_5 g11564(.A(new_n13912_1), .B(new_n13898), .Y(new_n13913));
  nand_5 g11565(.A(new_n13913), .B(new_n13897), .Y(new_n13914_1));
  nor_5  g11566(.A(new_n9927), .B(n20179), .Y(new_n13915));
  not_8  g11567(.A(new_n13915), .Y(new_n13916));
  nand_5 g11568(.A(new_n9927), .B(n20179), .Y(new_n13917));
  and_5  g11569(.A(new_n13917), .B(new_n13916), .Y(new_n13918));
  not_8  g11570(.A(new_n13918), .Y(new_n13919));
  nand_5 g11571(.A(new_n13919), .B(new_n8381_1), .Y(new_n13920));
  nand_5 g11572(.A(new_n13918), .B(new_n8383), .Y(new_n13921));
  nand_5 g11573(.A(new_n13921), .B(new_n13920), .Y(new_n13922_1));
  xnor_4 g11574(.A(new_n13922_1), .B(new_n13914_1), .Y(new_n13923_1));
  nand_5 g11575(.A(new_n13923_1), .B(new_n13896), .Y(new_n13924));
  not_8  g11576(.A(new_n13924), .Y(new_n13925));
  nor_5  g11577(.A(new_n13923_1), .B(new_n13896), .Y(new_n13926));
  nand_5 g11578(.A(new_n13867), .B(new_n13866), .Y(new_n13927));
  xor_4  g11579(.A(new_n13927), .B(new_n13886), .Y(new_n13928));
  not_8  g11580(.A(new_n13928), .Y(new_n13929));
  nand_5 g11581(.A(new_n13898), .B(new_n13897), .Y(new_n13930));
  xor_4  g11582(.A(new_n13930), .B(new_n13912_1), .Y(new_n13931));
  or_5   g11583(.A(new_n13931), .B(new_n13929), .Y(new_n13932));
  nand_5 g11584(.A(new_n13931), .B(new_n13929), .Y(new_n13933));
  nand_5 g11585(.A(new_n13870), .B(new_n13869), .Y(new_n13934));
  xor_4  g11586(.A(new_n13934), .B(new_n13884), .Y(new_n13935));
  not_8  g11587(.A(new_n13935), .Y(new_n13936));
  nand_5 g11588(.A(new_n13901), .B(new_n13899), .Y(new_n13937));
  xor_4  g11589(.A(new_n13937), .B(new_n13910), .Y(new_n13938));
  or_5   g11590(.A(new_n13938), .B(new_n13936), .Y(new_n13939));
  not_8  g11591(.A(new_n13939), .Y(new_n13940));
  nand_5 g11592(.A(new_n13938), .B(new_n13936), .Y(new_n13941));
  not_8  g11593(.A(new_n13941), .Y(new_n13942));
  nand_5 g11594(.A(new_n13874), .B(new_n13873), .Y(new_n13943));
  xor_4  g11595(.A(new_n13943), .B(new_n13882), .Y(new_n13944));
  not_8  g11596(.A(new_n13944), .Y(new_n13945));
  nand_5 g11597(.A(new_n13903), .B(new_n13902), .Y(new_n13946));
  xor_4  g11598(.A(new_n13946), .B(new_n13908), .Y(new_n13947));
  nand_5 g11599(.A(new_n13947), .B(new_n13945), .Y(new_n13948));
  nor_5  g11600(.A(new_n13947), .B(new_n13945), .Y(new_n13949));
  nor_5  g11601(.A(new_n13880), .B(new_n13879), .Y(new_n13950));
  xor_4  g11602(.A(new_n13950), .B(new_n6023), .Y(new_n13951_1));
  nand_5 g11603(.A(new_n13905), .B(new_n13904), .Y(new_n13952));
  xor_4  g11604(.A(new_n13952), .B(new_n13906), .Y(new_n13953));
  nand_5 g11605(.A(new_n13953), .B(new_n13951_1), .Y(new_n13954));
  not_8  g11606(.A(new_n13954), .Y(new_n13955));
  nor_5  g11607(.A(new_n13953), .B(new_n13951_1), .Y(new_n13956));
  xor_4  g11608(.A(new_n6030), .B(n13714), .Y(new_n13957));
  xor_4  g11609(.A(new_n8406), .B(new_n7784), .Y(new_n13958));
  nand_5 g11610(.A(new_n13958), .B(new_n13957), .Y(new_n13959));
  nor_5  g11611(.A(new_n13959), .B(new_n13956), .Y(new_n13960));
  nor_5  g11612(.A(new_n13960), .B(new_n13955), .Y(new_n13961));
  or_5   g11613(.A(new_n13961), .B(new_n13949), .Y(new_n13962));
  nand_5 g11614(.A(new_n13962), .B(new_n13948), .Y(new_n13963));
  nor_5  g11615(.A(new_n13963), .B(new_n13942), .Y(new_n13964));
  nor_5  g11616(.A(new_n13964), .B(new_n13940), .Y(new_n13965));
  not_8  g11617(.A(new_n13965), .Y(new_n13966));
  nand_5 g11618(.A(new_n13966), .B(new_n13933), .Y(new_n13967));
  nand_5 g11619(.A(new_n13967), .B(new_n13932), .Y(new_n13968));
  not_8  g11620(.A(new_n13968), .Y(new_n13969));
  nor_5  g11621(.A(new_n13969), .B(new_n13926), .Y(new_n13970));
  nor_5  g11622(.A(new_n13970), .B(new_n13925), .Y(new_n13971));
  not_8  g11623(.A(new_n13971), .Y(new_n13972));
  nand_5 g11624(.A(new_n13894), .B(new_n13888), .Y(new_n13973));
  nand_5 g11625(.A(new_n13973), .B(new_n13893), .Y(new_n13974));
  xor_4  g11626(.A(new_n13889), .B(n26318), .Y(new_n13975));
  nand_5 g11627(.A(new_n13975), .B(new_n5990), .Y(new_n13976));
  or_5   g11628(.A(new_n13975), .B(new_n5990), .Y(new_n13977));
  nand_5 g11629(.A(new_n13977), .B(new_n13976), .Y(new_n13978));
  xor_4  g11630(.A(new_n13978), .B(new_n13974), .Y(new_n13979));
  not_8  g11631(.A(new_n13979), .Y(new_n13980));
  nand_5 g11632(.A(new_n13921), .B(new_n13914_1), .Y(new_n13981));
  nand_5 g11633(.A(new_n13981), .B(new_n13920), .Y(new_n13982));
  nand_5 g11634(.A(new_n13915), .B(new_n7757), .Y(new_n13983));
  nand_5 g11635(.A(new_n13916), .B(n1112), .Y(new_n13984));
  and_5  g11636(.A(new_n13984), .B(new_n13983), .Y(new_n13985));
  not_8  g11637(.A(new_n13985), .Y(new_n13986));
  nand_5 g11638(.A(new_n13986), .B(new_n8376_1), .Y(new_n13987));
  nand_5 g11639(.A(new_n13985), .B(new_n8377), .Y(new_n13988));
  nand_5 g11640(.A(new_n13988), .B(new_n13987), .Y(new_n13989));
  xor_4  g11641(.A(new_n13989), .B(new_n13982), .Y(new_n13990));
  or_5   g11642(.A(new_n13990), .B(new_n13980), .Y(new_n13991));
  nand_5 g11643(.A(new_n13990), .B(new_n13980), .Y(new_n13992));
  nand_5 g11644(.A(new_n13992), .B(new_n13991), .Y(new_n13993));
  xor_4  g11645(.A(new_n13993), .B(new_n13972), .Y(n1891));
  nand_5 g11646(.A(new_n4377), .B(n6729), .Y(new_n13995));
  nand_5 g11647(.A(n10792), .B(new_n4422), .Y(new_n13996));
  nand_5 g11648(.A(new_n2636), .B(n19922), .Y(new_n13997));
  nand_5 g11649(.A(new_n13997), .B(new_n13996), .Y(new_n13998));
  nand_5 g11650(.A(new_n13998), .B(new_n13995), .Y(new_n13999));
  or_5   g11651(.A(n9323), .B(new_n4408), .Y(new_n14000));
  nand_5 g11652(.A(n9323), .B(new_n4408), .Y(new_n14001));
  nand_5 g11653(.A(new_n14001), .B(new_n14000), .Y(new_n14002));
  xor_4  g11654(.A(new_n14002), .B(new_n13999), .Y(new_n14003));
  or_5   g11655(.A(new_n14003), .B(new_n7446), .Y(new_n14004_1));
  nand_5 g11656(.A(new_n14003), .B(new_n7446), .Y(new_n14005));
  xor_4  g11657(.A(n21687), .B(new_n4378), .Y(new_n14006));
  nor_5  g11658(.A(new_n14006), .B(new_n7449), .Y(new_n14007));
  nand_5 g11659(.A(new_n13996), .B(new_n13995), .Y(new_n14008));
  xnor_4 g11660(.A(new_n14008), .B(new_n13997), .Y(new_n14009));
  nand_5 g11661(.A(new_n14009), .B(new_n14007), .Y(new_n14010));
  not_8  g11662(.A(new_n14010), .Y(new_n14011));
  nor_5  g11663(.A(new_n14009), .B(new_n14007), .Y(new_n14012));
  nor_5  g11664(.A(new_n14012), .B(new_n7455), .Y(new_n14013));
  nor_5  g11665(.A(new_n14013), .B(new_n14011), .Y(new_n14014));
  not_8  g11666(.A(new_n14014), .Y(new_n14015));
  nand_5 g11667(.A(new_n14015), .B(new_n14005), .Y(new_n14016));
  nand_5 g11668(.A(new_n14016), .B(new_n14004_1), .Y(new_n14017));
  nand_5 g11669(.A(new_n14001), .B(new_n13999), .Y(new_n14018));
  nand_5 g11670(.A(new_n14018), .B(new_n14000), .Y(new_n14019));
  or_5   g11671(.A(new_n4407), .B(n1949), .Y(new_n14020));
  nand_5 g11672(.A(new_n4407), .B(n1949), .Y(new_n14021));
  nand_5 g11673(.A(new_n14021), .B(new_n14020), .Y(new_n14022));
  xnor_4 g11674(.A(new_n14022), .B(new_n14019), .Y(new_n14023));
  nand_5 g11675(.A(new_n14023), .B(new_n7442), .Y(new_n14024));
  not_8  g11676(.A(new_n14024), .Y(new_n14025));
  nor_5  g11677(.A(new_n14023), .B(new_n7442), .Y(new_n14026));
  nor_5  g11678(.A(new_n14026), .B(new_n14025), .Y(new_n14027));
  xor_4  g11679(.A(new_n14027), .B(new_n14017), .Y(n1925));
  nand_5 g11680(.A(new_n8720), .B(new_n8719), .Y(new_n14029));
  xor_4  g11681(.A(new_n14029), .B(new_n8746), .Y(n1942));
  nand_5 g11682(.A(new_n7215), .B(new_n7214), .Y(new_n14031));
  xor_4  g11683(.A(new_n14031), .B(new_n7295), .Y(n1972));
  nor_5  g11684(.A(new_n10035), .B(n12507), .Y(new_n14033));
  nor_5  g11685(.A(new_n14033), .B(new_n10034), .Y(new_n14034));
  nand_5 g11686(.A(new_n9990), .B(new_n9151), .Y(new_n14035));
  nand_5 g11687(.A(new_n10035), .B(n12507), .Y(new_n14036_1));
  nand_5 g11688(.A(new_n14036_1), .B(new_n14035), .Y(new_n14037));
  nor_5  g11689(.A(new_n14037), .B(new_n14034), .Y(new_n14038));
  nor_5  g11690(.A(new_n14038), .B(new_n12654_1), .Y(new_n14039));
  nand_5 g11691(.A(new_n10166), .B(new_n10081), .Y(new_n14040));
  nand_5 g11692(.A(new_n14040), .B(new_n10080), .Y(new_n14041));
  nand_5 g11693(.A(new_n14041), .B(new_n14039), .Y(new_n14042));
  nand_5 g11694(.A(new_n14038), .B(new_n12654_1), .Y(new_n14043));
  or_5   g11695(.A(new_n14043), .B(new_n14041), .Y(new_n14044));
  nand_5 g11696(.A(new_n14044), .B(new_n14042), .Y(new_n14045));
  nor_5  g11697(.A(new_n14045), .B(new_n12736), .Y(new_n14046));
  xor_4  g11698(.A(new_n14045), .B(new_n12691), .Y(new_n14047));
  xor_4  g11699(.A(new_n14038), .B(new_n12654_1), .Y(new_n14048));
  xor_4  g11700(.A(new_n14048), .B(new_n14041), .Y(new_n14049));
  nand_5 g11701(.A(new_n14049), .B(new_n12691), .Y(new_n14050));
  not_8  g11702(.A(new_n14049), .Y(new_n14051));
  nand_5 g11703(.A(new_n14051), .B(new_n12736), .Y(new_n14052));
  or_5   g11704(.A(new_n12745), .B(new_n10167), .Y(new_n14053));
  nand_5 g11705(.A(new_n12745), .B(new_n10167), .Y(new_n14054));
  nand_5 g11706(.A(new_n12748), .B(new_n10174), .Y(new_n14055));
  or_5   g11707(.A(new_n12748), .B(new_n10174), .Y(new_n14056));
  or_5   g11708(.A(new_n12755), .B(new_n10181), .Y(new_n14057));
  nand_5 g11709(.A(new_n12755), .B(new_n10181), .Y(new_n14058));
  or_5   g11710(.A(new_n12762), .B(new_n10188), .Y(new_n14059_1));
  nand_5 g11711(.A(new_n12762), .B(new_n10188), .Y(new_n14060));
  or_5   g11712(.A(new_n12769), .B(new_n10195), .Y(new_n14061));
  nand_5 g11713(.A(new_n12769), .B(new_n10195), .Y(new_n14062));
  nand_5 g11714(.A(new_n12778), .B(new_n10203), .Y(new_n14063));
  nand_5 g11715(.A(new_n12776), .B(new_n10204), .Y(new_n14064));
  or_5   g11716(.A(new_n12781), .B(new_n10211), .Y(new_n14065));
  nand_5 g11717(.A(new_n12781), .B(new_n10211), .Y(new_n14066));
  or_5   g11718(.A(new_n12785), .B(new_n10217), .Y(new_n14067));
  nand_5 g11719(.A(new_n12785), .B(new_n10217), .Y(new_n14068));
  nand_5 g11720(.A(new_n12794), .B(new_n10224), .Y(new_n14069));
  or_5   g11721(.A(new_n14069), .B(new_n12791), .Y(new_n14070));
  not_8  g11722(.A(new_n10233), .Y(new_n14071_1));
  nand_5 g11723(.A(new_n14069), .B(new_n12791), .Y(new_n14072));
  nand_5 g11724(.A(new_n14072), .B(new_n14071_1), .Y(new_n14073));
  nand_5 g11725(.A(new_n14073), .B(new_n14070), .Y(new_n14074));
  nand_5 g11726(.A(new_n14074), .B(new_n14068), .Y(new_n14075));
  nand_5 g11727(.A(new_n14075), .B(new_n14067), .Y(new_n14076));
  nand_5 g11728(.A(new_n14076), .B(new_n14066), .Y(new_n14077));
  nand_5 g11729(.A(new_n14077), .B(new_n14065), .Y(new_n14078));
  nand_5 g11730(.A(new_n14078), .B(new_n14064), .Y(new_n14079));
  nand_5 g11731(.A(new_n14079), .B(new_n14063), .Y(new_n14080));
  nand_5 g11732(.A(new_n14080), .B(new_n14062), .Y(new_n14081_1));
  nand_5 g11733(.A(new_n14081_1), .B(new_n14061), .Y(new_n14082));
  nand_5 g11734(.A(new_n14082), .B(new_n14060), .Y(new_n14083));
  nand_5 g11735(.A(new_n14083), .B(new_n14059_1), .Y(new_n14084));
  nand_5 g11736(.A(new_n14084), .B(new_n14058), .Y(new_n14085));
  and_5  g11737(.A(new_n14085), .B(new_n14057), .Y(new_n14086));
  nand_5 g11738(.A(new_n14086), .B(new_n14056), .Y(new_n14087));
  nand_5 g11739(.A(new_n14087), .B(new_n14055), .Y(new_n14088));
  nand_5 g11740(.A(new_n14088), .B(new_n14054), .Y(new_n14089));
  nand_5 g11741(.A(new_n14089), .B(new_n14053), .Y(new_n14090_1));
  nand_5 g11742(.A(new_n14090_1), .B(new_n14052), .Y(new_n14091));
  nand_5 g11743(.A(new_n14091), .B(new_n14050), .Y(new_n14092));
  nor_5  g11744(.A(new_n14092), .B(new_n14047), .Y(new_n14093));
  nor_5  g11745(.A(new_n14093), .B(new_n14046), .Y(n1981));
  nand_5 g11746(.A(new_n14054), .B(new_n14053), .Y(new_n14095_1));
  xor_4  g11747(.A(new_n14095_1), .B(new_n14088), .Y(n2004));
  or_5   g11748(.A(new_n7054), .B(n10018), .Y(new_n14097));
  nand_5 g11749(.A(new_n7054), .B(n10018), .Y(new_n14098));
  not_8  g11750(.A(n2184), .Y(new_n14099));
  nand_5 g11751(.A(new_n7059), .B(new_n14099), .Y(new_n14100));
  nand_5 g11752(.A(new_n7057_1), .B(n2184), .Y(new_n14101));
  not_8  g11753(.A(n3541), .Y(new_n14102));
  nand_5 g11754(.A(new_n7064), .B(new_n14102), .Y(new_n14103));
  nand_5 g11755(.A(new_n7062), .B(n3541), .Y(new_n14104));
  nand_5 g11756(.A(new_n7067), .B(new_n7492), .Y(new_n14105));
  nand_5 g11757(.A(new_n7068), .B(n16818), .Y(new_n14106));
  or_5   g11758(.A(new_n4517), .B(n1269), .Y(new_n14107_1));
  nand_5 g11759(.A(new_n4517), .B(n1269), .Y(new_n14108));
  nand_5 g11760(.A(new_n4442), .B(new_n7361), .Y(new_n14109));
  nand_5 g11761(.A(new_n4443), .B(n14576), .Y(new_n14110));
  or_5   g11762(.A(new_n4401_1), .B(n2985), .Y(new_n14111));
  nand_5 g11763(.A(new_n4401_1), .B(n2985), .Y(new_n14112));
  or_5   g11764(.A(new_n4383), .B(n5605), .Y(new_n14113));
  nand_5 g11765(.A(new_n4383), .B(n5605), .Y(new_n14114));
  nand_5 g11766(.A(new_n4388), .B(new_n7331), .Y(new_n14115));
  nand_5 g11767(.A(new_n4389), .B(n15652), .Y(new_n14116));
  nand_5 g11768(.A(new_n4378), .B(n4939), .Y(new_n14117));
  nand_5 g11769(.A(new_n14117), .B(new_n14116), .Y(new_n14118));
  nand_5 g11770(.A(new_n14118), .B(new_n14115), .Y(new_n14119));
  nand_5 g11771(.A(new_n14119), .B(new_n14114), .Y(new_n14120));
  nand_5 g11772(.A(new_n14120), .B(new_n14113), .Y(new_n14121_1));
  nand_5 g11773(.A(new_n14121_1), .B(new_n14112), .Y(new_n14122));
  nand_5 g11774(.A(new_n14122), .B(new_n14111), .Y(new_n14123));
  nand_5 g11775(.A(new_n14123), .B(new_n14110), .Y(new_n14124));
  nand_5 g11776(.A(new_n14124), .B(new_n14109), .Y(new_n14125));
  nand_5 g11777(.A(new_n14125), .B(new_n14108), .Y(new_n14126_1));
  nand_5 g11778(.A(new_n14126_1), .B(new_n14107_1), .Y(new_n14127));
  nand_5 g11779(.A(new_n14127), .B(new_n14106), .Y(new_n14128));
  nand_5 g11780(.A(new_n14128), .B(new_n14105), .Y(new_n14129));
  nand_5 g11781(.A(new_n14129), .B(new_n14104), .Y(new_n14130_1));
  nand_5 g11782(.A(new_n14130_1), .B(new_n14103), .Y(new_n14131));
  nand_5 g11783(.A(new_n14131), .B(new_n14101), .Y(new_n14132));
  nand_5 g11784(.A(new_n14132), .B(new_n14100), .Y(new_n14133));
  nand_5 g11785(.A(new_n14133), .B(new_n14098), .Y(new_n14134));
  xor_4  g11786(.A(new_n14134), .B(new_n7051), .Y(new_n14135));
  nand_5 g11787(.A(new_n14135), .B(new_n14097), .Y(new_n14136_1));
  nand_5 g11788(.A(new_n14136_1), .B(new_n7044), .Y(new_n14137));
  or_5   g11789(.A(new_n14136_1), .B(new_n7044), .Y(new_n14138));
  and_5  g11790(.A(new_n14138), .B(new_n14137), .Y(new_n14139));
  nand_5 g11791(.A(new_n14098), .B(new_n14097), .Y(new_n14140));
  xor_4  g11792(.A(new_n14140), .B(new_n14133), .Y(new_n14141));
  or_5   g11793(.A(new_n14141), .B(new_n7087), .Y(new_n14142));
  nand_5 g11794(.A(new_n14141), .B(new_n7087), .Y(new_n14143));
  nand_5 g11795(.A(new_n14100), .B(new_n14101), .Y(new_n14144));
  xor_4  g11796(.A(new_n14144), .B(new_n14131), .Y(new_n14145));
  or_5   g11797(.A(new_n14145), .B(new_n7095), .Y(new_n14146));
  nand_5 g11798(.A(new_n14145), .B(new_n7095), .Y(new_n14147_1));
  nand_5 g11799(.A(new_n14103), .B(new_n14104), .Y(new_n14148_1));
  xor_4  g11800(.A(new_n14148_1), .B(new_n14129), .Y(new_n14149));
  or_5   g11801(.A(new_n14149), .B(new_n7103), .Y(new_n14150));
  nand_5 g11802(.A(new_n14149), .B(new_n7103), .Y(new_n14151));
  nand_5 g11803(.A(new_n14105), .B(new_n14106), .Y(new_n14152));
  xor_4  g11804(.A(new_n14152), .B(new_n14127), .Y(new_n14153));
  or_5   g11805(.A(new_n14153), .B(new_n7111), .Y(new_n14154));
  nand_5 g11806(.A(new_n14153), .B(new_n7111), .Y(new_n14155));
  nand_5 g11807(.A(new_n14107_1), .B(new_n14108), .Y(new_n14156));
  xor_4  g11808(.A(new_n14156), .B(new_n14125), .Y(new_n14157));
  or_5   g11809(.A(new_n14157), .B(new_n7120), .Y(new_n14158));
  nand_5 g11810(.A(new_n14157), .B(new_n7120), .Y(new_n14159));
  nand_5 g11811(.A(new_n14109), .B(new_n14110), .Y(new_n14160));
  xor_4  g11812(.A(new_n14160), .B(new_n14123), .Y(new_n14161));
  or_5   g11813(.A(new_n14161), .B(new_n7125), .Y(new_n14162));
  nand_5 g11814(.A(new_n14161), .B(new_n7125), .Y(new_n14163));
  nand_5 g11815(.A(new_n14111), .B(new_n14112), .Y(new_n14164));
  xor_4  g11816(.A(new_n14164), .B(new_n14121_1), .Y(new_n14165));
  or_5   g11817(.A(new_n14165), .B(new_n7128), .Y(new_n14166));
  nand_5 g11818(.A(new_n14165), .B(new_n7128), .Y(new_n14167));
  not_8  g11819(.A(new_n7132), .Y(new_n14168));
  nand_5 g11820(.A(new_n14113), .B(new_n14114), .Y(new_n14169));
  xor_4  g11821(.A(new_n14169), .B(new_n14119), .Y(new_n14170));
  or_5   g11822(.A(new_n14170), .B(new_n14168), .Y(new_n14171));
  nand_5 g11823(.A(new_n14170), .B(new_n14168), .Y(new_n14172));
  xor_4  g11824(.A(n19922), .B(new_n7330_1), .Y(new_n14173));
  not_8  g11825(.A(new_n14173), .Y(new_n14174_1));
  nand_5 g11826(.A(new_n14174_1), .B(new_n7142), .Y(new_n14175));
  not_8  g11827(.A(new_n14175), .Y(new_n14176));
  nand_5 g11828(.A(new_n14176), .B(new_n7136), .Y(new_n14177));
  nand_5 g11829(.A(new_n14175), .B(new_n7137), .Y(new_n14178));
  nand_5 g11830(.A(new_n14115), .B(new_n14116), .Y(new_n14179));
  xnor_4 g11831(.A(new_n14179), .B(new_n14117), .Y(new_n14180));
  nand_5 g11832(.A(new_n14180), .B(new_n14178), .Y(new_n14181));
  nand_5 g11833(.A(new_n14181), .B(new_n14177), .Y(new_n14182));
  nand_5 g11834(.A(new_n14182), .B(new_n14172), .Y(new_n14183));
  nand_5 g11835(.A(new_n14183), .B(new_n14171), .Y(new_n14184));
  nand_5 g11836(.A(new_n14184), .B(new_n14167), .Y(new_n14185));
  nand_5 g11837(.A(new_n14185), .B(new_n14166), .Y(new_n14186));
  nand_5 g11838(.A(new_n14186), .B(new_n14163), .Y(new_n14187));
  nand_5 g11839(.A(new_n14187), .B(new_n14162), .Y(new_n14188));
  nand_5 g11840(.A(new_n14188), .B(new_n14159), .Y(new_n14189));
  nand_5 g11841(.A(new_n14189), .B(new_n14158), .Y(new_n14190_1));
  nand_5 g11842(.A(new_n14190_1), .B(new_n14155), .Y(new_n14191));
  nand_5 g11843(.A(new_n14191), .B(new_n14154), .Y(new_n14192));
  nand_5 g11844(.A(new_n14192), .B(new_n14151), .Y(new_n14193));
  nand_5 g11845(.A(new_n14193), .B(new_n14150), .Y(new_n14194));
  nand_5 g11846(.A(new_n14194), .B(new_n14147_1), .Y(new_n14195));
  nand_5 g11847(.A(new_n14195), .B(new_n14146), .Y(new_n14196));
  nand_5 g11848(.A(new_n14196), .B(new_n14143), .Y(new_n14197));
  nand_5 g11849(.A(new_n14197), .B(new_n14142), .Y(new_n14198));
  xor_4  g11850(.A(new_n14198), .B(new_n14139), .Y(new_n14199));
  nand_5 g11851(.A(new_n7166), .B(n5140), .Y(new_n14200));
  not_8  g11852(.A(n5140), .Y(new_n14201));
  nand_5 g11853(.A(n6105), .B(new_n14201), .Y(new_n14202));
  nand_5 g11854(.A(n6204), .B(new_n7170), .Y(new_n14203));
  not_8  g11855(.A(n6204), .Y(new_n14204));
  nand_5 g11856(.A(new_n14204), .B(n3795), .Y(new_n14205));
  nand_5 g11857(.A(new_n7175), .B(n3349), .Y(new_n14206));
  not_8  g11858(.A(n3349), .Y(new_n14207));
  nand_5 g11859(.A(n25464), .B(new_n14207), .Y(new_n14208));
  nand_5 g11860(.A(new_n7178), .B(n1742), .Y(new_n14209));
  nand_5 g11861(.A(n4590), .B(new_n7491), .Y(new_n14210));
  nand_5 g11862(.A(new_n7182), .B(n4858), .Y(new_n14211_1));
  nand_5 g11863(.A(n26752), .B(new_n7416), .Y(new_n14212));
  nand_5 g11864(.A(n8244), .B(new_n7185), .Y(new_n14213));
  nand_5 g11865(.A(new_n7360), .B(n6513), .Y(new_n14214));
  nand_5 g11866(.A(n9493), .B(new_n7188), .Y(new_n14215));
  nand_5 g11867(.A(new_n7329), .B(n3918), .Y(new_n14216));
  nand_5 g11868(.A(n15167), .B(new_n4586), .Y(new_n14217));
  nand_5 g11869(.A(new_n7341), .B(n919), .Y(new_n14218));
  nand_5 g11870(.A(new_n4535), .B(n21095), .Y(new_n14219));
  nand_5 g11871(.A(n25316), .B(new_n7347), .Y(new_n14220));
  or_5   g11872(.A(new_n4573), .B(n8656), .Y(new_n14221));
  nand_5 g11873(.A(new_n14221), .B(new_n14220), .Y(new_n14222_1));
  nand_5 g11874(.A(new_n14222_1), .B(new_n14219), .Y(new_n14223));
  nand_5 g11875(.A(new_n14223), .B(new_n14218), .Y(new_n14224));
  nand_5 g11876(.A(new_n14224), .B(new_n14217), .Y(new_n14225));
  nand_5 g11877(.A(new_n14225), .B(new_n14216), .Y(new_n14226));
  nand_5 g11878(.A(new_n14226), .B(new_n14215), .Y(new_n14227));
  nand_5 g11879(.A(new_n14227), .B(new_n14214), .Y(new_n14228));
  nand_5 g11880(.A(new_n14228), .B(new_n14213), .Y(new_n14229));
  nand_5 g11881(.A(new_n14229), .B(new_n14212), .Y(new_n14230_1));
  nand_5 g11882(.A(new_n14230_1), .B(new_n14211_1), .Y(new_n14231));
  nand_5 g11883(.A(new_n14231), .B(new_n14210), .Y(new_n14232));
  nand_5 g11884(.A(new_n14232), .B(new_n14209), .Y(new_n14233));
  nand_5 g11885(.A(new_n14233), .B(new_n14208), .Y(new_n14234));
  nand_5 g11886(.A(new_n14234), .B(new_n14206), .Y(new_n14235));
  nand_5 g11887(.A(new_n14235), .B(new_n14205), .Y(new_n14236));
  nand_5 g11888(.A(new_n14236), .B(new_n14203), .Y(new_n14237));
  nand_5 g11889(.A(new_n14237), .B(new_n14202), .Y(new_n14238));
  nand_5 g11890(.A(new_n14238), .B(new_n14200), .Y(new_n14239));
  not_8  g11891(.A(new_n14239), .Y(new_n14240));
  nand_5 g11892(.A(new_n14240), .B(new_n14199), .Y(new_n14241));
  or_5   g11893(.A(new_n14240), .B(new_n14199), .Y(new_n14242));
  nand_5 g11894(.A(new_n14202), .B(new_n14200), .Y(new_n14243));
  xor_4  g11895(.A(new_n14243), .B(new_n14237), .Y(new_n14244));
  nand_5 g11896(.A(new_n14143), .B(new_n14142), .Y(new_n14245));
  xor_4  g11897(.A(new_n14245), .B(new_n14196), .Y(new_n14246));
  nand_5 g11898(.A(new_n14246), .B(new_n14244), .Y(new_n14247));
  or_5   g11899(.A(new_n14246), .B(new_n14244), .Y(new_n14248));
  nand_5 g11900(.A(new_n14205), .B(new_n14203), .Y(new_n14249));
  xor_4  g11901(.A(new_n14249), .B(new_n14235), .Y(new_n14250));
  not_8  g11902(.A(new_n14250), .Y(new_n14251));
  nand_5 g11903(.A(new_n14147_1), .B(new_n14146), .Y(new_n14252));
  xnor_4 g11904(.A(new_n14252), .B(new_n14194), .Y(new_n14253));
  or_5   g11905(.A(new_n14253), .B(new_n14251), .Y(new_n14254));
  nand_5 g11906(.A(new_n14253), .B(new_n14251), .Y(new_n14255));
  nand_5 g11907(.A(new_n14208), .B(new_n14206), .Y(new_n14256));
  xor_4  g11908(.A(new_n14256), .B(new_n14233), .Y(new_n14257));
  not_8  g11909(.A(new_n14257), .Y(new_n14258));
  nand_5 g11910(.A(new_n14151), .B(new_n14150), .Y(new_n14259));
  xnor_4 g11911(.A(new_n14259), .B(new_n14192), .Y(new_n14260));
  or_5   g11912(.A(new_n14260), .B(new_n14258), .Y(new_n14261));
  nand_5 g11913(.A(new_n14260), .B(new_n14258), .Y(new_n14262));
  nand_5 g11914(.A(new_n14210), .B(new_n14209), .Y(new_n14263));
  xor_4  g11915(.A(new_n14263), .B(new_n14231), .Y(new_n14264));
  not_8  g11916(.A(new_n14264), .Y(new_n14265));
  nand_5 g11917(.A(new_n14155), .B(new_n14154), .Y(new_n14266));
  xnor_4 g11918(.A(new_n14266), .B(new_n14190_1), .Y(new_n14267_1));
  or_5   g11919(.A(new_n14267_1), .B(new_n14265), .Y(new_n14268));
  nand_5 g11920(.A(new_n14267_1), .B(new_n14265), .Y(new_n14269));
  nand_5 g11921(.A(new_n14212), .B(new_n14211_1), .Y(new_n14270));
  xor_4  g11922(.A(new_n14270), .B(new_n14229), .Y(new_n14271_1));
  not_8  g11923(.A(new_n14271_1), .Y(new_n14272));
  nand_5 g11924(.A(new_n14159), .B(new_n14158), .Y(new_n14273));
  xnor_4 g11925(.A(new_n14273), .B(new_n14188), .Y(new_n14274));
  or_5   g11926(.A(new_n14274), .B(new_n14272), .Y(new_n14275_1));
  nand_5 g11927(.A(new_n14274), .B(new_n14272), .Y(new_n14276));
  nand_5 g11928(.A(new_n14214), .B(new_n14213), .Y(new_n14277_1));
  xor_4  g11929(.A(new_n14277_1), .B(new_n14227), .Y(new_n14278));
  nand_5 g11930(.A(new_n14163), .B(new_n14162), .Y(new_n14279));
  xor_4  g11931(.A(new_n14279), .B(new_n14186), .Y(new_n14280));
  nand_5 g11932(.A(new_n14280), .B(new_n14278), .Y(new_n14281));
  or_5   g11933(.A(new_n14280), .B(new_n14278), .Y(new_n14282));
  nand_5 g11934(.A(new_n14216), .B(new_n14215), .Y(new_n14283));
  xor_4  g11935(.A(new_n14283), .B(new_n14225), .Y(new_n14284));
  nand_5 g11936(.A(new_n14167), .B(new_n14166), .Y(new_n14285));
  xor_4  g11937(.A(new_n14285), .B(new_n14184), .Y(new_n14286));
  nand_5 g11938(.A(new_n14286), .B(new_n14284), .Y(new_n14287));
  nor_5  g11939(.A(new_n14286), .B(new_n14284), .Y(new_n14288));
  not_8  g11940(.A(new_n14288), .Y(new_n14289));
  nand_5 g11941(.A(new_n14218), .B(new_n14217), .Y(new_n14290));
  xor_4  g11942(.A(new_n14290), .B(new_n14223), .Y(new_n14291));
  nand_5 g11943(.A(new_n14172), .B(new_n14171), .Y(new_n14292));
  xor_4  g11944(.A(new_n14292), .B(new_n14182), .Y(new_n14293));
  nand_5 g11945(.A(new_n14293), .B(new_n14291), .Y(new_n14294_1));
  not_8  g11946(.A(new_n14294_1), .Y(new_n14295));
  nor_5  g11947(.A(new_n14293), .B(new_n14291), .Y(new_n14296));
  nand_5 g11948(.A(new_n4573), .B(n8656), .Y(new_n14297));
  and_5  g11949(.A(new_n14297), .B(new_n14221), .Y(new_n14298));
  nand_5 g11950(.A(new_n14173), .B(new_n7275), .Y(new_n14299));
  nand_5 g11951(.A(new_n14299), .B(new_n14175), .Y(new_n14300));
  nor_5  g11952(.A(new_n14300), .B(new_n14298), .Y(new_n14301));
  and_5  g11953(.A(new_n14220), .B(new_n14219), .Y(new_n14302));
  xor_4  g11954(.A(new_n14302), .B(new_n14221), .Y(new_n14303));
  or_5   g11955(.A(new_n14303), .B(new_n14301), .Y(new_n14304));
  nand_5 g11956(.A(new_n14303), .B(new_n14301), .Y(new_n14305));
  nand_5 g11957(.A(new_n14178), .B(new_n14177), .Y(new_n14306));
  xor_4  g11958(.A(new_n14306), .B(new_n14180), .Y(new_n14307));
  nand_5 g11959(.A(new_n14307), .B(new_n14305), .Y(new_n14308));
  nand_5 g11960(.A(new_n14308), .B(new_n14304), .Y(new_n14309));
  not_8  g11961(.A(new_n14309), .Y(new_n14310_1));
  nor_5  g11962(.A(new_n14310_1), .B(new_n14296), .Y(new_n14311));
  nor_5  g11963(.A(new_n14311), .B(new_n14295), .Y(new_n14312));
  not_8  g11964(.A(new_n14312), .Y(new_n14313));
  nand_5 g11965(.A(new_n14313), .B(new_n14289), .Y(new_n14314));
  nand_5 g11966(.A(new_n14314), .B(new_n14287), .Y(new_n14315));
  nand_5 g11967(.A(new_n14315), .B(new_n14282), .Y(new_n14316));
  nand_5 g11968(.A(new_n14316), .B(new_n14281), .Y(new_n14317));
  nand_5 g11969(.A(new_n14317), .B(new_n14276), .Y(new_n14318));
  nand_5 g11970(.A(new_n14318), .B(new_n14275_1), .Y(new_n14319));
  nand_5 g11971(.A(new_n14319), .B(new_n14269), .Y(new_n14320));
  nand_5 g11972(.A(new_n14320), .B(new_n14268), .Y(new_n14321));
  nand_5 g11973(.A(new_n14321), .B(new_n14262), .Y(new_n14322));
  nand_5 g11974(.A(new_n14322), .B(new_n14261), .Y(new_n14323_1));
  nand_5 g11975(.A(new_n14323_1), .B(new_n14255), .Y(new_n14324));
  nand_5 g11976(.A(new_n14324), .B(new_n14254), .Y(new_n14325));
  nand_5 g11977(.A(new_n14325), .B(new_n14248), .Y(new_n14326_1));
  and_5  g11978(.A(new_n14326_1), .B(new_n14247), .Y(new_n14327));
  nand_5 g11979(.A(new_n14327), .B(new_n14242), .Y(new_n14328));
  nand_5 g11980(.A(new_n14328), .B(new_n14241), .Y(new_n14329));
  nand_5 g11981(.A(new_n14198), .B(new_n14138), .Y(new_n14330));
  nor_5  g11982(.A(new_n14134), .B(new_n7052), .Y(new_n14331));
  not_8  g11983(.A(new_n14137), .Y(new_n14332));
  nor_5  g11984(.A(new_n14332), .B(new_n14331), .Y(new_n14333));
  nand_5 g11985(.A(new_n14333), .B(new_n14330), .Y(new_n14334));
  nor_5  g11986(.A(new_n14334), .B(new_n14329), .Y(n2007));
  nand_5 g11987(.A(new_n10219), .B(new_n10218), .Y(new_n14336));
  xor_4  g11988(.A(new_n14336), .B(new_n10235), .Y(n2061));
  nand_5 g11989(.A(new_n13031), .B(new_n8209), .Y(new_n14338));
  or_5   g11990(.A(new_n13031), .B(new_n8209), .Y(new_n14339));
  nand_5 g11991(.A(new_n13037), .B(new_n8215_1), .Y(new_n14340));
  or_5   g11992(.A(new_n13037), .B(new_n8215_1), .Y(new_n14341));
  nand_5 g11993(.A(new_n8221), .B(new_n5298), .Y(new_n14342_1));
  or_5   g11994(.A(new_n8221), .B(new_n5298), .Y(new_n14343));
  nand_5 g11995(.A(new_n8227), .B(new_n5208), .Y(new_n14344));
  or_5   g11996(.A(new_n8227), .B(new_n5208), .Y(new_n14345_1));
  nand_5 g11997(.A(new_n8233), .B(new_n5154), .Y(new_n14346));
  or_5   g11998(.A(new_n8233), .B(new_n5154), .Y(new_n14347));
  nand_5 g11999(.A(new_n8239), .B(new_n5177), .Y(new_n14348));
  or_5   g12000(.A(new_n8239), .B(new_n5177), .Y(new_n14349));
  nand_5 g12001(.A(new_n8243), .B(new_n5192), .Y(new_n14350));
  nand_5 g12002(.A(new_n14350), .B(new_n5184_1), .Y(new_n14351));
  or_5   g12003(.A(new_n14350), .B(new_n5184_1), .Y(new_n14352));
  nand_5 g12004(.A(new_n14352), .B(new_n8253), .Y(new_n14353_1));
  nand_5 g12005(.A(new_n14353_1), .B(new_n14351), .Y(new_n14354));
  nand_5 g12006(.A(new_n14354), .B(new_n14349), .Y(new_n14355));
  nand_5 g12007(.A(new_n14355), .B(new_n14348), .Y(new_n14356));
  nand_5 g12008(.A(new_n14356), .B(new_n14347), .Y(new_n14357));
  nand_5 g12009(.A(new_n14357), .B(new_n14346), .Y(new_n14358));
  nand_5 g12010(.A(new_n14358), .B(new_n14345_1), .Y(new_n14359));
  nand_5 g12011(.A(new_n14359), .B(new_n14344), .Y(new_n14360));
  nand_5 g12012(.A(new_n14360), .B(new_n14343), .Y(new_n14361));
  nand_5 g12013(.A(new_n14361), .B(new_n14342_1), .Y(new_n14362));
  nand_5 g12014(.A(new_n14362), .B(new_n14341), .Y(new_n14363));
  nand_5 g12015(.A(new_n14363), .B(new_n14340), .Y(new_n14364_1));
  nand_5 g12016(.A(new_n14364_1), .B(new_n14339), .Y(new_n14365));
  nand_5 g12017(.A(new_n14365), .B(new_n14338), .Y(new_n14366));
  or_5   g12018(.A(new_n13023), .B(new_n8203), .Y(new_n14367));
  nand_5 g12019(.A(new_n13023), .B(new_n8203), .Y(new_n14368));
  nand_5 g12020(.A(new_n14368), .B(new_n14367), .Y(new_n14369));
  xor_4  g12021(.A(new_n14369), .B(new_n14366), .Y(n2092));
  nand_5 g12022(.A(new_n2384), .B(new_n2377), .Y(new_n14371));
  or_5   g12023(.A(new_n14371), .B(n13708), .Y(new_n14372));
  nor_5  g12024(.A(new_n14372), .B(n19911), .Y(new_n14373));
  nand_5 g12025(.A(new_n14373), .B(new_n2411), .Y(new_n14374));
  nor_5  g12026(.A(new_n14374), .B(n18907), .Y(new_n14375_1));
  nand_5 g12027(.A(new_n14375_1), .B(new_n2569), .Y(new_n14376));
  nor_5  g12028(.A(new_n14376), .B(n4256), .Y(new_n14377));
  nand_5 g12029(.A(new_n14377), .B(new_n8144), .Y(new_n14378));
  xor_4  g12030(.A(new_n14378), .B(n26986), .Y(new_n14379));
  nor_5  g12031(.A(new_n14379), .B(n8305), .Y(new_n14380));
  xor_4  g12032(.A(new_n14377), .B(n21287), .Y(new_n14381));
  nand_5 g12033(.A(new_n14381), .B(new_n7994), .Y(new_n14382));
  or_5   g12034(.A(new_n14381), .B(new_n7994), .Y(new_n14383));
  xor_4  g12035(.A(new_n14376), .B(n4256), .Y(new_n14384));
  or_5   g12036(.A(new_n14384), .B(n13333), .Y(new_n14385));
  xor_4  g12037(.A(new_n14375_1), .B(new_n2569), .Y(new_n14386));
  or_5   g12038(.A(new_n14386), .B(n2210), .Y(new_n14387));
  xor_4  g12039(.A(new_n14374), .B(n18907), .Y(new_n14388));
  or_5   g12040(.A(new_n14388), .B(n20604), .Y(new_n14389));
  xor_4  g12041(.A(new_n14373), .B(new_n2411), .Y(new_n14390));
  or_5   g12042(.A(new_n14390), .B(n16158), .Y(new_n14391));
  xor_4  g12043(.A(new_n14372), .B(n19911), .Y(new_n14392));
  or_5   g12044(.A(new_n14392), .B(n5752), .Y(new_n14393));
  nand_5 g12045(.A(new_n14371), .B(n13708), .Y(new_n14394));
  and_5  g12046(.A(new_n14394), .B(new_n14372), .Y(new_n14395));
  or_5   g12047(.A(new_n14395), .B(n18171), .Y(new_n14396));
  nand_5 g12048(.A(n18409), .B(n5704), .Y(new_n14397));
  and_5  g12049(.A(new_n14397), .B(new_n14371), .Y(new_n14398));
  or_5   g12050(.A(new_n14398), .B(n25073), .Y(new_n14399));
  nand_5 g12051(.A(n22309), .B(n5704), .Y(new_n14400));
  nand_5 g12052(.A(new_n14398), .B(n25073), .Y(new_n14401));
  nand_5 g12053(.A(new_n14401), .B(new_n14400), .Y(new_n14402));
  nand_5 g12054(.A(new_n14402), .B(new_n14399), .Y(new_n14403));
  nand_5 g12055(.A(new_n14395), .B(n18171), .Y(new_n14404));
  nand_5 g12056(.A(new_n14404), .B(new_n14403), .Y(new_n14405));
  nand_5 g12057(.A(new_n14405), .B(new_n14396), .Y(new_n14406));
  nand_5 g12058(.A(new_n14392), .B(n5752), .Y(new_n14407));
  nand_5 g12059(.A(new_n14407), .B(new_n14406), .Y(new_n14408));
  nand_5 g12060(.A(new_n14408), .B(new_n14393), .Y(new_n14409));
  nand_5 g12061(.A(new_n14390), .B(n16158), .Y(new_n14410));
  nand_5 g12062(.A(new_n14410), .B(new_n14409), .Y(new_n14411));
  nand_5 g12063(.A(new_n14411), .B(new_n14391), .Y(new_n14412_1));
  nand_5 g12064(.A(new_n14388), .B(n20604), .Y(new_n14413));
  nand_5 g12065(.A(new_n14413), .B(new_n14412_1), .Y(new_n14414_1));
  nand_5 g12066(.A(new_n14414_1), .B(new_n14389), .Y(new_n14415));
  nand_5 g12067(.A(new_n14386), .B(n2210), .Y(new_n14416));
  nand_5 g12068(.A(new_n14416), .B(new_n14415), .Y(new_n14417));
  nand_5 g12069(.A(new_n14417), .B(new_n14387), .Y(new_n14418));
  nand_5 g12070(.A(new_n14384), .B(n13333), .Y(new_n14419));
  nand_5 g12071(.A(new_n14419), .B(new_n14418), .Y(new_n14420));
  nand_5 g12072(.A(new_n14420), .B(new_n14385), .Y(new_n14421));
  nand_5 g12073(.A(new_n14421), .B(new_n14383), .Y(new_n14422));
  nand_5 g12074(.A(new_n14422), .B(new_n14382), .Y(new_n14423));
  nor_5  g12075(.A(new_n14423), .B(new_n14380), .Y(new_n14424));
  or_5   g12076(.A(new_n14378), .B(n26986), .Y(new_n14425));
  nand_5 g12077(.A(new_n14379), .B(n8305), .Y(new_n14426));
  nand_5 g12078(.A(new_n14426), .B(new_n14425), .Y(new_n14427));
  nor_5  g12079(.A(new_n14427), .B(new_n14424), .Y(new_n14428));
  xor_4  g12080(.A(new_n14379), .B(n8305), .Y(new_n14429));
  xor_4  g12081(.A(new_n14429), .B(new_n14423), .Y(new_n14430));
  nor_5  g12082(.A(n7876), .B(n4964), .Y(new_n14431));
  nand_5 g12083(.A(new_n14431), .B(new_n4160), .Y(new_n14432));
  nor_5  g12084(.A(new_n14432), .B(n342), .Y(new_n14433));
  nand_5 g12085(.A(new_n14433), .B(new_n4177), .Y(new_n14434));
  nor_5  g12086(.A(new_n14434), .B(n22597), .Y(new_n14435));
  nand_5 g12087(.A(new_n14435), .B(new_n4297), .Y(new_n14436));
  nor_5  g12088(.A(new_n14436), .B(n26224), .Y(new_n14437));
  nand_5 g12089(.A(new_n14437), .B(new_n5363), .Y(new_n14438));
  xor_4  g12090(.A(new_n14438), .B(n9934), .Y(new_n14439));
  not_8  g12091(.A(new_n14439), .Y(new_n14440_1));
  nand_5 g12092(.A(new_n14440_1), .B(new_n14430), .Y(new_n14441));
  nand_5 g12093(.A(new_n14383), .B(new_n14382), .Y(new_n14442));
  xor_4  g12094(.A(new_n14442), .B(new_n14421), .Y(new_n14443));
  xor_4  g12095(.A(new_n14437), .B(new_n5363), .Y(new_n14444));
  nand_5 g12096(.A(new_n14444), .B(new_n14443), .Y(new_n14445));
  or_5   g12097(.A(new_n14444), .B(new_n14443), .Y(new_n14446));
  nand_5 g12098(.A(new_n14419), .B(new_n14385), .Y(new_n14447));
  xor_4  g12099(.A(new_n14447), .B(new_n14418), .Y(new_n14448));
  xor_4  g12100(.A(new_n14436), .B(n26224), .Y(new_n14449));
  nand_5 g12101(.A(new_n14449), .B(new_n14448), .Y(new_n14450));
  or_5   g12102(.A(new_n14449), .B(new_n14448), .Y(new_n14451));
  nand_5 g12103(.A(new_n14416), .B(new_n14387), .Y(new_n14452));
  xor_4  g12104(.A(new_n14452), .B(new_n14415), .Y(new_n14453));
  xor_4  g12105(.A(new_n14435), .B(new_n4297), .Y(new_n14454));
  nand_5 g12106(.A(new_n14454), .B(new_n14453), .Y(new_n14455));
  or_5   g12107(.A(new_n14454), .B(new_n14453), .Y(new_n14456));
  nand_5 g12108(.A(new_n14413), .B(new_n14389), .Y(new_n14457_1));
  xor_4  g12109(.A(new_n14457_1), .B(new_n14412_1), .Y(new_n14458));
  xor_4  g12110(.A(new_n14434), .B(n22597), .Y(new_n14459));
  nand_5 g12111(.A(new_n14459), .B(new_n14458), .Y(new_n14460));
  or_5   g12112(.A(new_n14459), .B(new_n14458), .Y(new_n14461));
  nand_5 g12113(.A(new_n14410), .B(new_n14391), .Y(new_n14462));
  xor_4  g12114(.A(new_n14462), .B(new_n14409), .Y(new_n14463));
  xor_4  g12115(.A(new_n14433), .B(new_n4177), .Y(new_n14464_1));
  nand_5 g12116(.A(new_n14464_1), .B(new_n14463), .Y(new_n14465));
  or_5   g12117(.A(new_n14464_1), .B(new_n14463), .Y(new_n14466));
  nand_5 g12118(.A(new_n14407), .B(new_n14393), .Y(new_n14467));
  xor_4  g12119(.A(new_n14467), .B(new_n14406), .Y(new_n14468));
  xor_4  g12120(.A(new_n14432), .B(n342), .Y(new_n14469));
  nand_5 g12121(.A(new_n14469), .B(new_n14468), .Y(new_n14470));
  or_5   g12122(.A(new_n14469), .B(new_n14468), .Y(new_n14471_1));
  nand_5 g12123(.A(new_n14404), .B(new_n14396), .Y(new_n14472));
  xor_4  g12124(.A(new_n14472), .B(new_n14403), .Y(new_n14473));
  xor_4  g12125(.A(new_n14431), .B(new_n4160), .Y(new_n14474));
  nand_5 g12126(.A(new_n14474), .B(new_n14473), .Y(new_n14475_1));
  nor_5  g12127(.A(new_n14474), .B(new_n14473), .Y(new_n14476));
  not_8  g12128(.A(new_n14476), .Y(new_n14477));
  nand_5 g12129(.A(new_n14401), .B(new_n14399), .Y(new_n14478));
  xor_4  g12130(.A(new_n14478), .B(new_n14400), .Y(new_n14479));
  nor_5  g12131(.A(new_n4207), .B(new_n5331), .Y(new_n14480));
  nor_5  g12132(.A(new_n14480), .B(new_n14431), .Y(new_n14481));
  nand_5 g12133(.A(new_n14481), .B(new_n14479), .Y(new_n14482));
  nor_5  g12134(.A(new_n14481), .B(new_n14479), .Y(new_n14483));
  not_8  g12135(.A(new_n14483), .Y(new_n14484));
  nand_5 g12136(.A(new_n5743), .B(new_n2377), .Y(new_n14485));
  and_5  g12137(.A(new_n14485), .B(new_n14400), .Y(new_n14486));
  nand_5 g12138(.A(new_n14486), .B(n7876), .Y(new_n14487));
  not_8  g12139(.A(new_n14487), .Y(new_n14488));
  nand_5 g12140(.A(new_n14488), .B(new_n14484), .Y(new_n14489));
  nand_5 g12141(.A(new_n14489), .B(new_n14482), .Y(new_n14490));
  nand_5 g12142(.A(new_n14490), .B(new_n14477), .Y(new_n14491));
  nand_5 g12143(.A(new_n14491), .B(new_n14475_1), .Y(new_n14492));
  nand_5 g12144(.A(new_n14492), .B(new_n14471_1), .Y(new_n14493));
  nand_5 g12145(.A(new_n14493), .B(new_n14470), .Y(new_n14494));
  nand_5 g12146(.A(new_n14494), .B(new_n14466), .Y(new_n14495));
  nand_5 g12147(.A(new_n14495), .B(new_n14465), .Y(new_n14496));
  nand_5 g12148(.A(new_n14496), .B(new_n14461), .Y(new_n14497));
  nand_5 g12149(.A(new_n14497), .B(new_n14460), .Y(new_n14498));
  nand_5 g12150(.A(new_n14498), .B(new_n14456), .Y(new_n14499));
  nand_5 g12151(.A(new_n14499), .B(new_n14455), .Y(new_n14500));
  nand_5 g12152(.A(new_n14500), .B(new_n14451), .Y(new_n14501));
  nand_5 g12153(.A(new_n14501), .B(new_n14450), .Y(new_n14502));
  nand_5 g12154(.A(new_n14502), .B(new_n14446), .Y(new_n14503));
  nand_5 g12155(.A(new_n14503), .B(new_n14445), .Y(new_n14504));
  nand_5 g12156(.A(new_n14504), .B(new_n14441), .Y(new_n14505));
  nor_5  g12157(.A(new_n14438), .B(n9934), .Y(new_n14506));
  not_8  g12158(.A(new_n14430), .Y(new_n14507));
  nand_5 g12159(.A(new_n14439), .B(new_n14507), .Y(new_n14508));
  not_8  g12160(.A(new_n14508), .Y(new_n14509));
  nor_5  g12161(.A(new_n14509), .B(new_n14506), .Y(new_n14510_1));
  nand_5 g12162(.A(new_n14510_1), .B(new_n14505), .Y(new_n14511));
  nor_5  g12163(.A(new_n14511), .B(new_n14428), .Y(new_n14512));
  nand_5 g12164(.A(n22253), .B(n10650), .Y(new_n14513));
  not_8  g12165(.A(n10650), .Y(new_n14514));
  nand_5 g12166(.A(new_n8015), .B(new_n14514), .Y(new_n14515));
  nand_5 g12167(.A(new_n14515), .B(new_n14513), .Y(new_n14516));
  not_8  g12168(.A(n12900), .Y(new_n14517));
  nand_5 g12169(.A(new_n14517), .B(new_n8020), .Y(new_n14518));
  nand_5 g12170(.A(n12900), .B(n1255), .Y(new_n14519));
  not_8  g12171(.A(n20411), .Y(new_n14520));
  nand_5 g12172(.A(new_n14520), .B(new_n8024), .Y(new_n14521));
  nand_5 g12173(.A(n20411), .B(n9512), .Y(new_n14522));
  not_8  g12174(.A(n17069), .Y(new_n14523));
  nand_5 g12175(.A(new_n14523), .B(new_n8027_1), .Y(new_n14524));
  nand_5 g12176(.A(n17069), .B(n16608), .Y(new_n14525));
  not_8  g12177(.A(n15918), .Y(new_n14526));
  nand_5 g12178(.A(new_n5317), .B(new_n14526), .Y(new_n14527));
  nand_5 g12179(.A(n21735), .B(n15918), .Y(new_n14528));
  not_8  g12180(.A(n17784), .Y(new_n14529));
  nand_5 g12181(.A(new_n5246), .B(new_n14529), .Y(new_n14530));
  nand_5 g12182(.A(n24085), .B(n17784), .Y(new_n14531));
  not_8  g12183(.A(n14323), .Y(new_n14532));
  nand_5 g12184(.A(new_n14532), .B(new_n5226_1), .Y(new_n14533));
  nand_5 g12185(.A(n14323), .B(n14071), .Y(new_n14534));
  not_8  g12186(.A(n2886), .Y(new_n14535));
  nand_5 g12187(.A(new_n14535), .B(new_n5230), .Y(new_n14536));
  nand_5 g12188(.A(n2886), .B(n1738), .Y(new_n14537));
  not_8  g12189(.A(n1040), .Y(new_n14538));
  nand_5 g12190(.A(new_n5234), .B(new_n14538), .Y(new_n14539));
  nand_5 g12191(.A(n12152), .B(n1040), .Y(new_n14540));
  nand_5 g12192(.A(n19107), .B(n9090), .Y(new_n14541_1));
  nand_5 g12193(.A(new_n14541_1), .B(new_n14540), .Y(new_n14542));
  nand_5 g12194(.A(new_n14542), .B(new_n14539), .Y(new_n14543));
  nand_5 g12195(.A(new_n14543), .B(new_n14537), .Y(new_n14544));
  nand_5 g12196(.A(new_n14544), .B(new_n14536), .Y(new_n14545));
  nand_5 g12197(.A(new_n14545), .B(new_n14534), .Y(new_n14546_1));
  nand_5 g12198(.A(new_n14546_1), .B(new_n14533), .Y(new_n14547_1));
  nand_5 g12199(.A(new_n14547_1), .B(new_n14531), .Y(new_n14548));
  nand_5 g12200(.A(new_n14548), .B(new_n14530), .Y(new_n14549));
  nand_5 g12201(.A(new_n14549), .B(new_n14528), .Y(new_n14550));
  nand_5 g12202(.A(new_n14550), .B(new_n14527), .Y(new_n14551));
  nand_5 g12203(.A(new_n14551), .B(new_n14525), .Y(new_n14552));
  nand_5 g12204(.A(new_n14552), .B(new_n14524), .Y(new_n14553));
  nand_5 g12205(.A(new_n14553), .B(new_n14522), .Y(new_n14554));
  nand_5 g12206(.A(new_n14554), .B(new_n14521), .Y(new_n14555));
  nand_5 g12207(.A(new_n14555), .B(new_n14519), .Y(new_n14556));
  nand_5 g12208(.A(new_n14556), .B(new_n14518), .Y(new_n14557));
  not_8  g12209(.A(new_n14557), .Y(new_n14558));
  xor_4  g12210(.A(new_n14558), .B(new_n14516), .Y(new_n14559));
  or_5   g12211(.A(new_n14559), .B(n2272), .Y(new_n14560));
  nand_5 g12212(.A(new_n14559), .B(n2272), .Y(new_n14561));
  nand_5 g12213(.A(new_n14519), .B(new_n14518), .Y(new_n14562));
  xor_4  g12214(.A(new_n14562), .B(new_n14555), .Y(new_n14563));
  nand_5 g12215(.A(new_n14563), .B(new_n8146), .Y(new_n14564));
  or_5   g12216(.A(new_n14563), .B(new_n8146), .Y(new_n14565));
  nand_5 g12217(.A(new_n14522), .B(new_n14521), .Y(new_n14566));
  xor_4  g12218(.A(new_n14566), .B(new_n14553), .Y(new_n14567));
  nand_5 g12219(.A(new_n14567), .B(new_n8150), .Y(new_n14568));
  or_5   g12220(.A(new_n14567), .B(new_n8150), .Y(new_n14569));
  nand_5 g12221(.A(new_n14525), .B(new_n14524), .Y(new_n14570_1));
  xor_4  g12222(.A(new_n14570_1), .B(new_n14551), .Y(new_n14571));
  nand_5 g12223(.A(new_n14571), .B(new_n8153), .Y(new_n14572));
  or_5   g12224(.A(new_n14571), .B(new_n8153), .Y(new_n14573));
  nand_5 g12225(.A(new_n14528), .B(new_n14527), .Y(new_n14574));
  xor_4  g12226(.A(new_n14574), .B(new_n14549), .Y(new_n14575_1));
  nand_5 g12227(.A(new_n14575_1), .B(new_n8156), .Y(new_n14576_1));
  nor_5  g12228(.A(new_n14575_1), .B(new_n8156), .Y(new_n14577));
  not_8  g12229(.A(new_n14577), .Y(new_n14578));
  nand_5 g12230(.A(new_n14531), .B(new_n14530), .Y(new_n14579));
  xor_4  g12231(.A(new_n14579), .B(new_n14547_1), .Y(new_n14580));
  nand_5 g12232(.A(new_n14580), .B(new_n8159_1), .Y(new_n14581));
  nor_5  g12233(.A(new_n14580), .B(new_n8159_1), .Y(new_n14582));
  not_8  g12234(.A(new_n14582), .Y(new_n14583));
  nand_5 g12235(.A(new_n14534), .B(new_n14533), .Y(new_n14584));
  xor_4  g12236(.A(new_n14584), .B(new_n14545), .Y(new_n14585));
  nand_5 g12237(.A(new_n14585), .B(new_n8162), .Y(new_n14586));
  nor_5  g12238(.A(new_n14585), .B(new_n8162), .Y(new_n14587));
  not_8  g12239(.A(new_n14587), .Y(new_n14588));
  nand_5 g12240(.A(new_n14537), .B(new_n14536), .Y(new_n14589));
  xor_4  g12241(.A(new_n14589), .B(new_n14543), .Y(new_n14590));
  nand_5 g12242(.A(new_n14590), .B(new_n8165), .Y(new_n14591));
  nor_5  g12243(.A(new_n14590), .B(new_n8165), .Y(new_n14592));
  nand_5 g12244(.A(new_n5236), .B(new_n12526), .Y(new_n14593_1));
  and_5  g12245(.A(new_n14593_1), .B(new_n14541_1), .Y(new_n14594));
  or_5   g12246(.A(new_n14594), .B(new_n8170), .Y(new_n14595));
  nor_5  g12247(.A(new_n14595), .B(new_n8168), .Y(new_n14596));
  not_8  g12248(.A(new_n14596), .Y(new_n14597));
  nand_5 g12249(.A(new_n14595), .B(new_n8168), .Y(new_n14598));
  nand_5 g12250(.A(new_n14540), .B(new_n14539), .Y(new_n14599));
  xor_4  g12251(.A(new_n14599), .B(new_n14541_1), .Y(new_n14600));
  not_8  g12252(.A(new_n14600), .Y(new_n14601));
  nand_5 g12253(.A(new_n14601), .B(new_n14598), .Y(new_n14602));
  nand_5 g12254(.A(new_n14602), .B(new_n14597), .Y(new_n14603_1));
  or_5   g12255(.A(new_n14603_1), .B(new_n14592), .Y(new_n14604));
  nand_5 g12256(.A(new_n14604), .B(new_n14591), .Y(new_n14605));
  nand_5 g12257(.A(new_n14605), .B(new_n14588), .Y(new_n14606));
  nand_5 g12258(.A(new_n14606), .B(new_n14586), .Y(new_n14607));
  nand_5 g12259(.A(new_n14607), .B(new_n14583), .Y(new_n14608));
  nand_5 g12260(.A(new_n14608), .B(new_n14581), .Y(new_n14609));
  nand_5 g12261(.A(new_n14609), .B(new_n14578), .Y(new_n14610));
  nand_5 g12262(.A(new_n14610), .B(new_n14576_1), .Y(new_n14611));
  nand_5 g12263(.A(new_n14611), .B(new_n14573), .Y(new_n14612));
  nand_5 g12264(.A(new_n14612), .B(new_n14572), .Y(new_n14613));
  nand_5 g12265(.A(new_n14613), .B(new_n14569), .Y(new_n14614));
  nand_5 g12266(.A(new_n14614), .B(new_n14568), .Y(new_n14615));
  nand_5 g12267(.A(new_n14615), .B(new_n14565), .Y(new_n14616));
  nand_5 g12268(.A(new_n14616), .B(new_n14564), .Y(new_n14617));
  nand_5 g12269(.A(new_n14617), .B(new_n14561), .Y(new_n14618));
  nand_5 g12270(.A(new_n14618), .B(new_n14560), .Y(new_n14619));
  nand_5 g12271(.A(new_n14557), .B(new_n14513), .Y(new_n14620));
  nand_5 g12272(.A(new_n14620), .B(new_n14515), .Y(new_n14621));
  not_8  g12273(.A(new_n14621), .Y(new_n14622));
  nor_5  g12274(.A(new_n14622), .B(new_n14619), .Y(new_n14623));
  xor_4  g12275(.A(new_n14511), .B(new_n14428), .Y(new_n14624));
  xor_4  g12276(.A(new_n14622), .B(new_n14619), .Y(new_n14625));
  nor_5  g12277(.A(new_n14625), .B(new_n14624), .Y(new_n14626));
  nand_5 g12278(.A(new_n14561), .B(new_n14560), .Y(new_n14627));
  xor_4  g12279(.A(new_n14627), .B(new_n14617), .Y(new_n14628));
  and_5  g12280(.A(new_n14508), .B(new_n14441), .Y(new_n14629));
  xor_4  g12281(.A(new_n14629), .B(new_n14504), .Y(new_n14630));
  not_8  g12282(.A(new_n14630), .Y(new_n14631));
  nand_5 g12283(.A(new_n14631), .B(new_n14628), .Y(new_n14632));
  not_8  g12284(.A(new_n14632), .Y(new_n14633_1));
  nor_5  g12285(.A(new_n14631), .B(new_n14628), .Y(new_n14634));
  nand_5 g12286(.A(new_n14446), .B(new_n14445), .Y(new_n14635));
  xor_4  g12287(.A(new_n14635), .B(new_n14502), .Y(new_n14636_1));
  nand_5 g12288(.A(new_n14565), .B(new_n14564), .Y(new_n14637));
  xor_4  g12289(.A(new_n14637), .B(new_n14615), .Y(new_n14638));
  nand_5 g12290(.A(new_n14638), .B(new_n14636_1), .Y(new_n14639));
  not_8  g12291(.A(new_n14639), .Y(new_n14640));
  nor_5  g12292(.A(new_n14638), .B(new_n14636_1), .Y(new_n14641));
  nand_5 g12293(.A(new_n14451), .B(new_n14450), .Y(new_n14642));
  xor_4  g12294(.A(new_n14642), .B(new_n14500), .Y(new_n14643));
  nand_5 g12295(.A(new_n14569), .B(new_n14568), .Y(new_n14644));
  xor_4  g12296(.A(new_n14644), .B(new_n14613), .Y(new_n14645));
  nand_5 g12297(.A(new_n14645), .B(new_n14643), .Y(new_n14646));
  not_8  g12298(.A(new_n14646), .Y(new_n14647));
  nor_5  g12299(.A(new_n14645), .B(new_n14643), .Y(new_n14648));
  nand_5 g12300(.A(new_n14456), .B(new_n14455), .Y(new_n14649));
  xor_4  g12301(.A(new_n14649), .B(new_n14498), .Y(new_n14650));
  nand_5 g12302(.A(new_n14573), .B(new_n14572), .Y(new_n14651));
  xor_4  g12303(.A(new_n14651), .B(new_n14611), .Y(new_n14652));
  nand_5 g12304(.A(new_n14652), .B(new_n14650), .Y(new_n14653));
  not_8  g12305(.A(new_n14653), .Y(new_n14654));
  nor_5  g12306(.A(new_n14652), .B(new_n14650), .Y(new_n14655));
  nand_5 g12307(.A(new_n14461), .B(new_n14460), .Y(new_n14656));
  xor_4  g12308(.A(new_n14656), .B(new_n14496), .Y(new_n14657));
  nand_5 g12309(.A(new_n14578), .B(new_n14576_1), .Y(new_n14658));
  xor_4  g12310(.A(new_n14658), .B(new_n14609), .Y(new_n14659));
  nand_5 g12311(.A(new_n14659), .B(new_n14657), .Y(new_n14660));
  not_8  g12312(.A(new_n14660), .Y(new_n14661));
  nor_5  g12313(.A(new_n14659), .B(new_n14657), .Y(new_n14662));
  nand_5 g12314(.A(new_n14466), .B(new_n14465), .Y(new_n14663));
  xor_4  g12315(.A(new_n14663), .B(new_n14494), .Y(new_n14664));
  nand_5 g12316(.A(new_n14583), .B(new_n14581), .Y(new_n14665));
  xor_4  g12317(.A(new_n14665), .B(new_n14607), .Y(new_n14666));
  nand_5 g12318(.A(new_n14666), .B(new_n14664), .Y(new_n14667));
  or_5   g12319(.A(new_n14666), .B(new_n14664), .Y(new_n14668));
  nand_5 g12320(.A(new_n14471_1), .B(new_n14470), .Y(new_n14669));
  xor_4  g12321(.A(new_n14669), .B(new_n14492), .Y(new_n14670));
  nand_5 g12322(.A(new_n14588), .B(new_n14586), .Y(new_n14671));
  xor_4  g12323(.A(new_n14671), .B(new_n14605), .Y(new_n14672));
  nand_5 g12324(.A(new_n14672), .B(new_n14670), .Y(new_n14673));
  or_5   g12325(.A(new_n14672), .B(new_n14670), .Y(new_n14674));
  not_8  g12326(.A(new_n14592), .Y(new_n14675));
  nand_5 g12327(.A(new_n14675), .B(new_n14591), .Y(new_n14676));
  xor_4  g12328(.A(new_n14676), .B(new_n14603_1), .Y(new_n14677));
  nand_5 g12329(.A(new_n14477), .B(new_n14475_1), .Y(new_n14678));
  xor_4  g12330(.A(new_n14678), .B(new_n14490), .Y(new_n14679));
  not_8  g12331(.A(new_n14679), .Y(new_n14680_1));
  or_5   g12332(.A(new_n14680_1), .B(new_n14677), .Y(new_n14681));
  nand_5 g12333(.A(new_n14680_1), .B(new_n14677), .Y(new_n14682));
  nand_5 g12334(.A(new_n14597), .B(new_n14598), .Y(new_n14683));
  xor_4  g12335(.A(new_n14683), .B(new_n14601), .Y(new_n14684_1));
  nand_5 g12336(.A(new_n14484), .B(new_n14482), .Y(new_n14685));
  xor_4  g12337(.A(new_n14685), .B(new_n14488), .Y(new_n14686));
  not_8  g12338(.A(new_n14686), .Y(new_n14687));
  or_5   g12339(.A(new_n14687), .B(new_n14684_1), .Y(new_n14688));
  nand_5 g12340(.A(new_n14687), .B(new_n14684_1), .Y(new_n14689));
  xor_4  g12341(.A(new_n14594), .B(new_n8170), .Y(new_n14690));
  not_8  g12342(.A(new_n14690), .Y(new_n14691));
  nor_5  g12343(.A(new_n14486), .B(n7876), .Y(new_n14692_1));
  nor_5  g12344(.A(new_n14692_1), .B(new_n14488), .Y(new_n14693));
  nand_5 g12345(.A(new_n14693), .B(new_n14691), .Y(new_n14694));
  nand_5 g12346(.A(new_n14694), .B(new_n14689), .Y(new_n14695));
  nand_5 g12347(.A(new_n14695), .B(new_n14688), .Y(new_n14696));
  nand_5 g12348(.A(new_n14696), .B(new_n14682), .Y(new_n14697));
  nand_5 g12349(.A(new_n14697), .B(new_n14681), .Y(new_n14698));
  nand_5 g12350(.A(new_n14698), .B(new_n14674), .Y(new_n14699));
  nand_5 g12351(.A(new_n14699), .B(new_n14673), .Y(new_n14700));
  nand_5 g12352(.A(new_n14700), .B(new_n14668), .Y(new_n14701_1));
  nand_5 g12353(.A(new_n14701_1), .B(new_n14667), .Y(new_n14702_1));
  not_8  g12354(.A(new_n14702_1), .Y(new_n14703));
  nor_5  g12355(.A(new_n14703), .B(new_n14662), .Y(new_n14704_1));
  nor_5  g12356(.A(new_n14704_1), .B(new_n14661), .Y(new_n14705));
  nor_5  g12357(.A(new_n14705), .B(new_n14655), .Y(new_n14706));
  nor_5  g12358(.A(new_n14706), .B(new_n14654), .Y(new_n14707));
  nor_5  g12359(.A(new_n14707), .B(new_n14648), .Y(new_n14708));
  nor_5  g12360(.A(new_n14708), .B(new_n14647), .Y(new_n14709));
  nor_5  g12361(.A(new_n14709), .B(new_n14641), .Y(new_n14710));
  nor_5  g12362(.A(new_n14710), .B(new_n14640), .Y(new_n14711));
  nor_5  g12363(.A(new_n14711), .B(new_n14634), .Y(new_n14712));
  nor_5  g12364(.A(new_n14712), .B(new_n14633_1), .Y(new_n14713));
  nor_5  g12365(.A(new_n14713), .B(new_n14626), .Y(new_n14714));
  or_5   g12366(.A(new_n14714), .B(new_n14623), .Y(new_n14715));
  nand_5 g12367(.A(new_n14714), .B(new_n14623), .Y(new_n14716));
  nand_5 g12368(.A(new_n14716), .B(new_n14715), .Y(new_n14717));
  nand_5 g12369(.A(new_n14625), .B(new_n14624), .Y(new_n14718));
  nand_5 g12370(.A(new_n14718), .B(new_n14717), .Y(new_n14719));
  xnor_4 g12371(.A(new_n14719), .B(new_n14512), .Y(n2095));
  nand_5 g12372(.A(new_n13094), .B(new_n13095), .Y(new_n14721));
  xnor_4 g12373(.A(new_n14721), .B(new_n13112), .Y(n2105));
  nand_5 g12374(.A(new_n12202), .B(new_n12199), .Y(new_n14723));
  nand_5 g12375(.A(new_n14723), .B(new_n12201), .Y(new_n14724));
  not_8  g12376(.A(new_n14724), .Y(new_n14725));
  nand_5 g12377(.A(new_n8434), .B(new_n10473), .Y(new_n14726));
  nand_5 g12378(.A(n19941), .B(n10577), .Y(new_n14727));
  nand_5 g12379(.A(new_n14727), .B(new_n14726), .Y(new_n14728));
  xor_4  g12380(.A(new_n14728), .B(new_n14725), .Y(new_n14729));
  not_8  g12381(.A(new_n14729), .Y(new_n14730));
  nand_5 g12382(.A(new_n14730), .B(n18035), .Y(new_n14731));
  nand_5 g12383(.A(new_n14729), .B(new_n12392), .Y(new_n14732));
  nand_5 g12384(.A(new_n12208), .B(new_n12197), .Y(new_n14733));
  nand_5 g12385(.A(new_n14733), .B(new_n12206), .Y(new_n14734_1));
  nand_5 g12386(.A(new_n14734_1), .B(new_n14732), .Y(new_n14735));
  nand_5 g12387(.A(new_n14735), .B(new_n14731), .Y(new_n14736));
  nand_5 g12388(.A(new_n14727), .B(new_n14724), .Y(new_n14737));
  nand_5 g12389(.A(new_n14737), .B(new_n14726), .Y(new_n14738));
  not_8  g12390(.A(new_n14738), .Y(new_n14739));
  nand_5 g12391(.A(new_n10468), .B(new_n8431), .Y(new_n14740));
  nand_5 g12392(.A(n23166), .B(n11898), .Y(new_n14741));
  nand_5 g12393(.A(new_n14741), .B(new_n14740), .Y(new_n14742));
  xor_4  g12394(.A(new_n14742), .B(new_n14739), .Y(new_n14743));
  not_8  g12395(.A(new_n14743), .Y(new_n14744));
  nand_5 g12396(.A(new_n14744), .B(n8827), .Y(new_n14745));
  nand_5 g12397(.A(new_n14743), .B(new_n12403), .Y(new_n14746_1));
  nand_5 g12398(.A(new_n14746_1), .B(new_n14745), .Y(new_n14747));
  xor_4  g12399(.A(new_n14747), .B(new_n14736), .Y(new_n14748));
  nand_5 g12400(.A(new_n14748), .B(new_n6911), .Y(new_n14749));
  not_8  g12401(.A(new_n6911), .Y(new_n14750));
  not_8  g12402(.A(new_n14748), .Y(new_n14751));
  nand_5 g12403(.A(new_n14751), .B(new_n14750), .Y(new_n14752));
  nand_5 g12404(.A(new_n14752), .B(new_n14749), .Y(new_n14753));
  not_8  g12405(.A(new_n6916), .Y(new_n14754));
  nand_5 g12406(.A(new_n14731), .B(new_n14732), .Y(new_n14755));
  xor_4  g12407(.A(new_n14755), .B(new_n14734_1), .Y(new_n14756));
  not_8  g12408(.A(new_n14756), .Y(new_n14757));
  nand_5 g12409(.A(new_n14757), .B(new_n14754), .Y(new_n14758));
  nand_5 g12410(.A(new_n14756), .B(new_n6916), .Y(new_n14759));
  or_5   g12411(.A(new_n12210), .B(new_n6923), .Y(new_n14760));
  nand_5 g12412(.A(new_n12210), .B(new_n6923), .Y(new_n14761));
  not_8  g12413(.A(new_n6930), .Y(new_n14762));
  nand_5 g12414(.A(new_n12162), .B(new_n14762), .Y(new_n14763_1));
  nand_5 g12415(.A(new_n12161_1), .B(new_n6930), .Y(new_n14764));
  not_8  g12416(.A(new_n6937), .Y(new_n14765));
  nand_5 g12417(.A(new_n12170), .B(new_n14765), .Y(new_n14766));
  nand_5 g12418(.A(new_n12169), .B(new_n6937), .Y(new_n14767));
  not_8  g12419(.A(new_n6943), .Y(new_n14768));
  nand_5 g12420(.A(new_n12178), .B(new_n14768), .Y(new_n14769));
  nand_5 g12421(.A(new_n12177), .B(new_n6943), .Y(new_n14770));
  not_8  g12422(.A(new_n6950), .Y(new_n14771));
  nand_5 g12423(.A(new_n9688), .B(new_n14771), .Y(new_n14772_1));
  nand_5 g12424(.A(new_n9687), .B(new_n6950), .Y(new_n14773));
  not_8  g12425(.A(new_n6956), .Y(new_n14774));
  nand_5 g12426(.A(new_n9701), .B(new_n14774), .Y(new_n14775));
  nand_5 g12427(.A(new_n9700), .B(new_n6956), .Y(new_n14776));
  nand_5 g12428(.A(new_n9708), .B(new_n6963), .Y(new_n14777));
  nand_5 g12429(.A(new_n9706), .B(new_n6962), .Y(new_n14778));
  not_8  g12430(.A(new_n9713), .Y(new_n14779));
  nor_5  g12431(.A(new_n14779), .B(new_n6567_1), .Y(new_n14780));
  nand_5 g12432(.A(new_n14780), .B(new_n14778), .Y(new_n14781));
  nand_5 g12433(.A(new_n14781), .B(new_n14777), .Y(new_n14782));
  nand_5 g12434(.A(new_n14782), .B(new_n14776), .Y(new_n14783));
  nand_5 g12435(.A(new_n14783), .B(new_n14775), .Y(new_n14784));
  nand_5 g12436(.A(new_n14784), .B(new_n14773), .Y(new_n14785));
  nand_5 g12437(.A(new_n14785), .B(new_n14772_1), .Y(new_n14786));
  nand_5 g12438(.A(new_n14786), .B(new_n14770), .Y(new_n14787));
  nand_5 g12439(.A(new_n14787), .B(new_n14769), .Y(new_n14788));
  nand_5 g12440(.A(new_n14788), .B(new_n14767), .Y(new_n14789));
  nand_5 g12441(.A(new_n14789), .B(new_n14766), .Y(new_n14790_1));
  nand_5 g12442(.A(new_n14790_1), .B(new_n14764), .Y(new_n14791));
  nand_5 g12443(.A(new_n14791), .B(new_n14763_1), .Y(new_n14792));
  nand_5 g12444(.A(new_n14792), .B(new_n14761), .Y(new_n14793));
  nand_5 g12445(.A(new_n14793), .B(new_n14760), .Y(new_n14794));
  nand_5 g12446(.A(new_n14794), .B(new_n14759), .Y(new_n14795));
  nand_5 g12447(.A(new_n14795), .B(new_n14758), .Y(new_n14796));
  xor_4  g12448(.A(new_n14796), .B(new_n14753), .Y(n2122));
  nand_5 g12449(.A(new_n2950), .B(new_n2949), .Y(new_n14798));
  xnor_4 g12450(.A(new_n14798), .B(new_n2984), .Y(n2147));
  nand_5 g12451(.A(new_n12051), .B(new_n12050), .Y(new_n14800));
  xor_4  g12452(.A(new_n14800), .B(new_n12099), .Y(n2209));
  xor_4  g12453(.A(new_n6554), .B(new_n6338), .Y(n2214));
  nand_5 g12454(.A(new_n12855), .B(new_n4736), .Y(new_n14803));
  nand_5 g12455(.A(new_n12856), .B(new_n4651), .Y(new_n14804));
  nand_5 g12456(.A(new_n12861_1), .B(new_n4742), .Y(new_n14805));
  nand_5 g12457(.A(new_n12860), .B(new_n4741), .Y(new_n14806));
  nand_5 g12458(.A(new_n12871_1), .B(new_n4746), .Y(new_n14807));
  or_5   g12459(.A(new_n12871_1), .B(new_n4746), .Y(new_n14808));
  nand_5 g12460(.A(new_n12866), .B(new_n4757), .Y(new_n14809));
  nand_5 g12461(.A(new_n14809), .B(new_n14808), .Y(new_n14810));
  nand_5 g12462(.A(new_n14810), .B(new_n14807), .Y(new_n14811));
  nand_5 g12463(.A(new_n14811), .B(new_n14806), .Y(new_n14812));
  nand_5 g12464(.A(new_n14812), .B(new_n14805), .Y(new_n14813));
  not_8  g12465(.A(new_n14813), .Y(new_n14814));
  nand_5 g12466(.A(new_n14814), .B(new_n14804), .Y(new_n14815));
  nand_5 g12467(.A(new_n14815), .B(new_n14803), .Y(new_n14816));
  nand_5 g12468(.A(new_n12850), .B(new_n4808), .Y(new_n14817));
  nand_5 g12469(.A(new_n12851), .B(new_n4777_1), .Y(new_n14818));
  nand_5 g12470(.A(new_n14818), .B(new_n14817), .Y(new_n14819_1));
  xnor_4 g12471(.A(new_n14819_1), .B(new_n14816), .Y(n2238));
  nand_5 g12472(.A(new_n12853), .B(new_n12852), .Y(new_n14821));
  xor_4  g12473(.A(new_n14821), .B(new_n12877), .Y(n2327));
  nand_5 g12474(.A(new_n6463), .B(new_n6462), .Y(new_n14823));
  xnor_4 g12475(.A(new_n14823), .B(new_n6503), .Y(n2343));
  nand_5 g12476(.A(new_n7630_1), .B(new_n7598_1), .Y(new_n14825));
  nand_5 g12477(.A(new_n14825), .B(new_n7633), .Y(new_n14826_1));
  nand_5 g12478(.A(new_n7612), .B(new_n7600), .Y(new_n14827_1));
  nand_5 g12479(.A(new_n14827_1), .B(new_n7611), .Y(new_n14828));
  not_8  g12480(.A(new_n14828), .Y(new_n14829));
  nand_5 g12481(.A(new_n7608), .B(new_n7603), .Y(new_n14830));
  nand_5 g12482(.A(new_n14830), .B(new_n7607_1), .Y(new_n14831));
  not_8  g12483(.A(new_n14831), .Y(new_n14832));
  nand_5 g12484(.A(new_n8306_1), .B(new_n8813), .Y(new_n14833));
  nand_5 g12485(.A(n20923), .B(n16524), .Y(new_n14834));
  nand_5 g12486(.A(new_n14834), .B(new_n14833), .Y(new_n14835));
  xor_4  g12487(.A(new_n14835), .B(new_n14832), .Y(new_n14836));
  or_5   g12488(.A(new_n14836), .B(new_n4880), .Y(new_n14837));
  nand_5 g12489(.A(new_n14836), .B(new_n4880), .Y(new_n14838));
  nand_5 g12490(.A(new_n14838), .B(new_n14837), .Y(new_n14839_1));
  xor_4  g12491(.A(new_n14839_1), .B(new_n14829), .Y(new_n14840));
  nand_5 g12492(.A(new_n7627), .B(new_n7616_1), .Y(new_n14841));
  nand_5 g12493(.A(new_n14841), .B(new_n7626), .Y(new_n14842));
  nand_5 g12494(.A(new_n12139), .B(n13453), .Y(new_n14843));
  nand_5 g12495(.A(new_n12141), .B(new_n5385), .Y(new_n14844));
  nand_5 g12496(.A(new_n14844), .B(new_n14843), .Y(new_n14845));
  xor_4  g12497(.A(new_n14845), .B(new_n14842), .Y(new_n14846));
  nand_5 g12498(.A(new_n14846), .B(new_n14840), .Y(new_n14847));
  not_8  g12499(.A(new_n14840), .Y(new_n14848));
  not_8  g12500(.A(new_n14846), .Y(new_n14849_1));
  nand_5 g12501(.A(new_n14849_1), .B(new_n14848), .Y(new_n14850));
  nand_5 g12502(.A(new_n14850), .B(new_n14847), .Y(new_n14851));
  xor_4  g12503(.A(new_n14851), .B(new_n14826_1), .Y(n2361));
  xor_4  g12504(.A(new_n4045), .B(new_n4043), .Y(n2363));
  nand_5 g12505(.A(new_n5083), .B(new_n5082_1), .Y(new_n14854));
  xnor_4 g12506(.A(new_n14854), .B(new_n5121), .Y(n2374));
  nand_5 g12507(.A(new_n6639), .B(new_n6631_1), .Y(new_n14856));
  nand_5 g12508(.A(new_n14856), .B(new_n6638), .Y(new_n14857));
  nand_5 g12509(.A(new_n6635), .B(new_n6633), .Y(new_n14858));
  nand_5 g12510(.A(new_n14858), .B(new_n6634_1), .Y(new_n14859));
  nand_5 g12511(.A(new_n14859), .B(new_n4098), .Y(new_n14860));
  not_8  g12512(.A(new_n14860), .Y(new_n14861));
  nor_5  g12513(.A(new_n14859), .B(new_n4098), .Y(new_n14862));
  nor_5  g12514(.A(new_n14862), .B(new_n14861), .Y(new_n14863));
  xor_4  g12515(.A(new_n14863), .B(new_n5532_1), .Y(new_n14864));
  or_5   g12516(.A(new_n14864), .B(new_n5453), .Y(new_n14865));
  nand_5 g12517(.A(new_n14864), .B(new_n5453), .Y(new_n14866));
  nand_5 g12518(.A(new_n14866), .B(new_n14865), .Y(new_n14867));
  xor_4  g12519(.A(new_n14867), .B(new_n14857), .Y(new_n14868));
  or_5   g12520(.A(new_n14868), .B(new_n4192), .Y(new_n14869));
  nand_5 g12521(.A(new_n14868), .B(new_n4192), .Y(new_n14870));
  nand_5 g12522(.A(new_n6643), .B(new_n6629), .Y(new_n14871));
  nand_5 g12523(.A(new_n14871), .B(new_n6642), .Y(new_n14872));
  nand_5 g12524(.A(new_n14872), .B(new_n14870), .Y(new_n14873));
  nand_5 g12525(.A(new_n14873), .B(new_n14869), .Y(new_n14874));
  nor_5  g12526(.A(new_n14862), .B(n7305), .Y(new_n14875));
  nor_5  g12527(.A(new_n14875), .B(new_n14861), .Y(new_n14876));
  not_8  g12528(.A(new_n14876), .Y(new_n14877));
  nand_5 g12529(.A(new_n14877), .B(new_n4082), .Y(new_n14878));
  nand_5 g12530(.A(new_n14876), .B(n626), .Y(new_n14879));
  and_5  g12531(.A(new_n14879), .B(new_n14878), .Y(new_n14880));
  xor_4  g12532(.A(new_n14880), .B(new_n5526), .Y(new_n14881));
  nand_5 g12533(.A(new_n14866), .B(new_n14857), .Y(new_n14882));
  nand_5 g12534(.A(new_n14882), .B(new_n14865), .Y(new_n14883));
  not_8  g12535(.A(new_n14883), .Y(new_n14884));
  or_5   g12536(.A(new_n14884), .B(new_n14881), .Y(new_n14885));
  nand_5 g12537(.A(new_n14884), .B(new_n14881), .Y(new_n14886));
  nand_5 g12538(.A(new_n14886), .B(new_n14885), .Y(new_n14887));
  xor_4  g12539(.A(new_n14887), .B(new_n5447), .Y(new_n14888));
  nand_5 g12540(.A(new_n14888), .B(new_n4186_1), .Y(new_n14889));
  or_5   g12541(.A(new_n14888), .B(new_n4186_1), .Y(new_n14890));
  nand_5 g12542(.A(new_n14890), .B(new_n14889), .Y(new_n14891_1));
  xnor_4 g12543(.A(new_n14891_1), .B(new_n14874), .Y(n2388));
  nand_5 g12544(.A(n11220), .B(n3425), .Y(new_n14893));
  nand_5 g12545(.A(new_n11623), .B(new_n8597), .Y(new_n14894));
  nand_5 g12546(.A(new_n14894), .B(new_n14893), .Y(new_n14895));
  nand_5 g12547(.A(new_n6139), .B(new_n6136), .Y(new_n14896));
  nand_5 g12548(.A(new_n14896), .B(new_n6138), .Y(new_n14897));
  xor_4  g12549(.A(new_n14897), .B(new_n14895), .Y(new_n14898));
  nand_5 g12550(.A(n7335), .B(n2160), .Y(new_n14899_1));
  nand_5 g12551(.A(new_n3314), .B(new_n13565), .Y(new_n14900));
  nand_5 g12552(.A(new_n14900), .B(new_n14899_1), .Y(new_n14901));
  nand_5 g12553(.A(new_n6147), .B(new_n6144), .Y(new_n14902));
  nand_5 g12554(.A(new_n14902), .B(new_n6146), .Y(new_n14903));
  not_8  g12555(.A(new_n14903), .Y(new_n14904));
  xor_4  g12556(.A(new_n14904), .B(new_n14901), .Y(new_n14905));
  or_5   g12557(.A(new_n14905), .B(new_n14898), .Y(new_n14906));
  nand_5 g12558(.A(new_n14905), .B(new_n14898), .Y(new_n14907));
  nand_5 g12559(.A(new_n14907), .B(new_n14906), .Y(new_n14908));
  nand_5 g12560(.A(new_n6151), .B(new_n6134), .Y(new_n14909));
  nand_5 g12561(.A(new_n14909), .B(new_n6150), .Y(new_n14910));
  xor_4  g12562(.A(new_n14910), .B(new_n14908), .Y(new_n14911));
  not_8  g12563(.A(new_n14911), .Y(new_n14912));
  xor_4  g12564(.A(new_n6157), .B(n7593), .Y(new_n14913));
  nand_5 g12565(.A(new_n14913), .B(n5025), .Y(new_n14914));
  nor_5  g12566(.A(new_n14913), .B(n5025), .Y(new_n14915));
  not_8  g12567(.A(new_n14915), .Y(new_n14916));
  nand_5 g12568(.A(new_n14916), .B(new_n14914), .Y(new_n14917));
  nand_5 g12569(.A(new_n6161), .B(new_n6156), .Y(new_n14918));
  nand_5 g12570(.A(new_n14918), .B(new_n6160_1), .Y(new_n14919));
  xor_4  g12571(.A(new_n14919), .B(new_n14917), .Y(new_n14920));
  nand_5 g12572(.A(new_n14920), .B(new_n14912), .Y(new_n14921));
  not_8  g12573(.A(new_n14921), .Y(new_n14922));
  nor_5  g12574(.A(new_n14920), .B(new_n14912), .Y(new_n14923));
  nor_5  g12575(.A(new_n14923), .B(new_n14922), .Y(new_n14924));
  nand_5 g12576(.A(new_n6164), .B(new_n6132), .Y(new_n14925));
  and_5  g12577(.A(new_n14925), .B(new_n6165), .Y(new_n14926));
  xor_4  g12578(.A(new_n14926), .B(new_n14924), .Y(n2440));
  nand_5 g12579(.A(new_n13260), .B(new_n13259), .Y(new_n14928));
  xor_4  g12580(.A(new_n14928), .B(new_n13276), .Y(n2444));
  nand_5 g12581(.A(new_n5702), .B(new_n3508), .Y(new_n14930));
  not_8  g12582(.A(new_n14930), .Y(new_n14931_1));
  nor_5  g12583(.A(new_n5702), .B(new_n3508), .Y(new_n14932));
  nor_5  g12584(.A(new_n14932), .B(new_n14931_1), .Y(n2513));
  not_8  g12585(.A(new_n12525), .Y(new_n14934));
  not_8  g12586(.A(new_n6770), .Y(new_n14935));
  nand_5 g12587(.A(new_n14935), .B(new_n14538), .Y(new_n14936));
  nand_5 g12588(.A(new_n6770), .B(n1040), .Y(new_n14937));
  and_5  g12589(.A(new_n14937), .B(new_n14936), .Y(new_n14938));
  xor_4  g12590(.A(new_n14938), .B(new_n14934), .Y(new_n14939));
  not_8  g12591(.A(new_n14939), .Y(new_n14940));
  nand_5 g12592(.A(new_n14940), .B(new_n6685), .Y(new_n14941));
  nand_5 g12593(.A(new_n14939), .B(n24374), .Y(new_n14942));
  nand_5 g12594(.A(new_n12528), .B(n14575), .Y(new_n14943));
  nand_5 g12595(.A(new_n14943), .B(new_n14942), .Y(new_n14944_1));
  nand_5 g12596(.A(new_n14944_1), .B(new_n14941), .Y(new_n14945));
  nand_5 g12597(.A(new_n14937), .B(new_n12525), .Y(new_n14946));
  nand_5 g12598(.A(new_n14946), .B(new_n14936), .Y(new_n14947));
  nand_5 g12599(.A(new_n6758), .B(new_n14535), .Y(new_n14948));
  nand_5 g12600(.A(new_n6757), .B(n2886), .Y(new_n14949));
  nand_5 g12601(.A(new_n14949), .B(new_n14948), .Y(new_n14950));
  xor_4  g12602(.A(new_n14950), .B(new_n14947), .Y(new_n14951));
  or_5   g12603(.A(new_n14951), .B(n7949), .Y(new_n14952));
  nand_5 g12604(.A(new_n14951), .B(n7949), .Y(new_n14953));
  nand_5 g12605(.A(new_n14953), .B(new_n14952), .Y(new_n14954_1));
  xor_4  g12606(.A(new_n14954_1), .B(new_n14945), .Y(new_n14955));
  or_5   g12607(.A(new_n14955), .B(new_n14680_1), .Y(new_n14956));
  nand_5 g12608(.A(new_n14955), .B(new_n14680_1), .Y(new_n14957));
  nand_5 g12609(.A(new_n14941), .B(new_n14942), .Y(new_n14958));
  xor_4  g12610(.A(new_n14958), .B(new_n14943), .Y(new_n14959));
  or_5   g12611(.A(new_n14959), .B(new_n14687), .Y(new_n14960));
  nand_5 g12612(.A(new_n14959), .B(new_n14687), .Y(new_n14961));
  xor_4  g12613(.A(new_n12528), .B(n14575), .Y(new_n14962));
  nand_5 g12614(.A(new_n14962), .B(new_n14693), .Y(new_n14963));
  nand_5 g12615(.A(new_n14963), .B(new_n14961), .Y(new_n14964));
  nand_5 g12616(.A(new_n14964), .B(new_n14960), .Y(new_n14965));
  nand_5 g12617(.A(new_n14965), .B(new_n14957), .Y(new_n14966));
  nand_5 g12618(.A(new_n14966), .B(new_n14956), .Y(new_n14967));
  not_8  g12619(.A(new_n14967), .Y(new_n14968));
  nand_5 g12620(.A(new_n14953), .B(new_n14945), .Y(new_n14969));
  nand_5 g12621(.A(new_n14969), .B(new_n14952), .Y(new_n14970));
  nand_5 g12622(.A(new_n14949), .B(new_n14947), .Y(new_n14971));
  nand_5 g12623(.A(new_n14971), .B(new_n14948), .Y(new_n14972));
  not_8  g12624(.A(new_n14972), .Y(new_n14973));
  nand_5 g12625(.A(new_n6750), .B(new_n14532), .Y(new_n14974));
  nand_5 g12626(.A(new_n6749), .B(n14323), .Y(new_n14975));
  nand_5 g12627(.A(new_n14975), .B(new_n14974), .Y(new_n14976));
  xor_4  g12628(.A(new_n14976), .B(new_n14973), .Y(new_n14977_1));
  nand_5 g12629(.A(new_n14977_1), .B(new_n6681), .Y(new_n14978));
  not_8  g12630(.A(new_n14977_1), .Y(new_n14979));
  nand_5 g12631(.A(new_n14979), .B(n12562), .Y(new_n14980));
  nand_5 g12632(.A(new_n14980), .B(new_n14978), .Y(new_n14981));
  xor_4  g12633(.A(new_n14981), .B(new_n14970), .Y(new_n14982));
  not_8  g12634(.A(new_n14982), .Y(new_n14983));
  nand_5 g12635(.A(new_n14983), .B(new_n14670), .Y(new_n14984));
  not_8  g12636(.A(new_n14984), .Y(new_n14985));
  nor_5  g12637(.A(new_n14983), .B(new_n14670), .Y(new_n14986));
  nor_5  g12638(.A(new_n14986), .B(new_n14985), .Y(new_n14987));
  xor_4  g12639(.A(new_n14987), .B(new_n14968), .Y(n2515));
  nand_5 g12640(.A(new_n12481), .B(new_n12480), .Y(new_n14989_1));
  xor_4  g12641(.A(new_n14989_1), .B(new_n12517), .Y(n2533));
  nor_5  g12642(.A(new_n8091), .B(new_n5867), .Y(new_n14991));
  nand_5 g12643(.A(new_n14991), .B(new_n8085), .Y(new_n14992));
  or_5   g12644(.A(new_n14992), .B(new_n8077), .Y(new_n14993));
  nor_5  g12645(.A(new_n14993), .B(new_n8071), .Y(new_n14994));
  nand_5 g12646(.A(new_n14994), .B(new_n8013), .Y(new_n14995));
  not_8  g12647(.A(new_n14995), .Y(new_n14996));
  nor_5  g12648(.A(new_n14994), .B(new_n8013), .Y(new_n14997));
  or_5   g12649(.A(new_n14997), .B(new_n14996), .Y(new_n14998));
  nand_5 g12650(.A(new_n14998), .B(new_n3361), .Y(new_n14999));
  xor_4  g12651(.A(new_n14993), .B(new_n8071), .Y(new_n15000));
  nand_5 g12652(.A(new_n15000), .B(new_n3363), .Y(new_n15001));
  or_5   g12653(.A(new_n15000), .B(new_n3363), .Y(new_n15002_1));
  nand_5 g12654(.A(new_n14992), .B(new_n8077), .Y(new_n15003));
  and_5  g12655(.A(new_n15003), .B(new_n14993), .Y(new_n15004_1));
  nand_5 g12656(.A(new_n15004_1), .B(new_n3369), .Y(new_n15005));
  or_5   g12657(.A(new_n15004_1), .B(new_n3369), .Y(new_n15006));
  not_8  g12658(.A(new_n14991), .Y(new_n15007));
  nand_5 g12659(.A(new_n15007), .B(new_n8084), .Y(new_n15008));
  and_5  g12660(.A(new_n15008), .B(new_n14992), .Y(new_n15009));
  nand_5 g12661(.A(new_n15009), .B(new_n3375), .Y(new_n15010));
  or_5   g12662(.A(new_n15009), .B(new_n3375), .Y(new_n15011_1));
  nand_5 g12663(.A(new_n8091), .B(new_n5867), .Y(new_n15012));
  and_5  g12664(.A(new_n15012), .B(new_n15007), .Y(new_n15013));
  nand_5 g12665(.A(new_n15013), .B(new_n3381), .Y(new_n15014));
  or_5   g12666(.A(new_n15013), .B(new_n3381), .Y(new_n15015));
  nand_5 g12667(.A(new_n5871), .B(new_n5860), .Y(new_n15016));
  nand_5 g12668(.A(new_n15016), .B(new_n5870), .Y(new_n15017));
  nand_5 g12669(.A(new_n15017), .B(new_n15015), .Y(new_n15018));
  nand_5 g12670(.A(new_n15018), .B(new_n15014), .Y(new_n15019_1));
  nand_5 g12671(.A(new_n15019_1), .B(new_n15011_1), .Y(new_n15020));
  nand_5 g12672(.A(new_n15020), .B(new_n15010), .Y(new_n15021));
  nand_5 g12673(.A(new_n15021), .B(new_n15006), .Y(new_n15022));
  nand_5 g12674(.A(new_n15022), .B(new_n15005), .Y(new_n15023));
  nand_5 g12675(.A(new_n15023), .B(new_n15002_1), .Y(new_n15024));
  nand_5 g12676(.A(new_n15024), .B(new_n15001), .Y(new_n15025));
  nand_5 g12677(.A(new_n15025), .B(new_n14999), .Y(new_n15026));
  not_8  g12678(.A(new_n15026), .Y(new_n15027));
  or_5   g12679(.A(new_n14998), .B(new_n3361), .Y(new_n15028));
  nand_5 g12680(.A(new_n15028), .B(new_n14995), .Y(new_n15029));
  nor_5  g12681(.A(new_n15029), .B(new_n15027), .Y(new_n15030));
  nand_5 g12682(.A(new_n8140), .B(n3425), .Y(new_n15031_1));
  nand_5 g12683(.A(n26986), .B(new_n8597), .Y(new_n15032));
  nand_5 g12684(.A(new_n8144), .B(n9967), .Y(new_n15033_1));
  nand_5 g12685(.A(n21287), .B(new_n3442), .Y(new_n15034));
  nand_5 g12686(.A(n20946), .B(new_n8148_1), .Y(new_n15035));
  nand_5 g12687(.A(new_n6062), .B(n4256), .Y(new_n15036));
  nand_5 g12688(.A(new_n2569), .B(n7751), .Y(new_n15037));
  nand_5 g12689(.A(n22332), .B(new_n2584), .Y(new_n15038));
  nand_5 g12690(.A(n26823), .B(new_n2474), .Y(new_n15039));
  nand_5 g12691(.A(new_n2468), .B(n18907), .Y(new_n15040));
  nand_5 g12692(.A(new_n9667), .B(new_n9665), .Y(new_n15041));
  nand_5 g12693(.A(new_n15041), .B(new_n9666), .Y(new_n15042));
  nand_5 g12694(.A(new_n15042), .B(new_n15040), .Y(new_n15043));
  nand_5 g12695(.A(new_n15043), .B(new_n15039), .Y(new_n15044));
  nand_5 g12696(.A(new_n15044), .B(new_n15038), .Y(new_n15045));
  nand_5 g12697(.A(new_n15045), .B(new_n15037), .Y(new_n15046));
  nand_5 g12698(.A(new_n15046), .B(new_n15036), .Y(new_n15047));
  nand_5 g12699(.A(new_n15047), .B(new_n15035), .Y(new_n15048));
  nand_5 g12700(.A(new_n15048), .B(new_n15034), .Y(new_n15049));
  nand_5 g12701(.A(new_n15049), .B(new_n15033_1), .Y(new_n15050));
  nand_5 g12702(.A(new_n15050), .B(new_n15032), .Y(new_n15051));
  nand_5 g12703(.A(new_n15051), .B(new_n15031_1), .Y(new_n15052_1));
  nor_5  g12704(.A(new_n15052_1), .B(new_n15030), .Y(new_n15053_1));
  not_8  g12705(.A(new_n15030), .Y(new_n15054));
  not_8  g12706(.A(new_n15052_1), .Y(new_n15055));
  nor_5  g12707(.A(new_n15055), .B(new_n15054), .Y(new_n15056));
  nor_5  g12708(.A(new_n15056), .B(new_n15053_1), .Y(new_n15057));
  nand_5 g12709(.A(new_n15028), .B(new_n14999), .Y(new_n15058));
  xor_4  g12710(.A(new_n15058), .B(new_n15025), .Y(new_n15059));
  nor_5  g12711(.A(new_n15059), .B(new_n15052_1), .Y(new_n15060));
  not_8  g12712(.A(new_n15059), .Y(new_n15061));
  nor_5  g12713(.A(new_n15061), .B(new_n15055), .Y(new_n15062));
  nand_5 g12714(.A(new_n15032), .B(new_n15031_1), .Y(new_n15063));
  xor_4  g12715(.A(new_n15063), .B(new_n15050), .Y(new_n15064));
  nand_5 g12716(.A(new_n15002_1), .B(new_n15001), .Y(new_n15065));
  xor_4  g12717(.A(new_n15065), .B(new_n15023), .Y(new_n15066));
  nand_5 g12718(.A(new_n15066), .B(new_n15064), .Y(new_n15067));
  or_5   g12719(.A(new_n15066), .B(new_n15064), .Y(new_n15068));
  nand_5 g12720(.A(new_n15034), .B(new_n15033_1), .Y(new_n15069));
  xor_4  g12721(.A(new_n15069), .B(new_n15048), .Y(new_n15070));
  nand_5 g12722(.A(new_n15006), .B(new_n15005), .Y(new_n15071));
  xor_4  g12723(.A(new_n15071), .B(new_n15021), .Y(new_n15072));
  nand_5 g12724(.A(new_n15072), .B(new_n15070), .Y(new_n15073));
  or_5   g12725(.A(new_n15072), .B(new_n15070), .Y(new_n15074));
  nand_5 g12726(.A(new_n15036), .B(new_n15035), .Y(new_n15075));
  xor_4  g12727(.A(new_n15075), .B(new_n15046), .Y(new_n15076));
  nand_5 g12728(.A(new_n15011_1), .B(new_n15010), .Y(new_n15077_1));
  xor_4  g12729(.A(new_n15077_1), .B(new_n15019_1), .Y(new_n15078));
  nand_5 g12730(.A(new_n15078), .B(new_n15076), .Y(new_n15079));
  or_5   g12731(.A(new_n15078), .B(new_n15076), .Y(new_n15080));
  nand_5 g12732(.A(new_n15038), .B(new_n15037), .Y(new_n15081));
  xor_4  g12733(.A(new_n15081), .B(new_n15044), .Y(new_n15082_1));
  nand_5 g12734(.A(new_n15015), .B(new_n15014), .Y(new_n15083));
  xor_4  g12735(.A(new_n15083), .B(new_n15017), .Y(new_n15084));
  nand_5 g12736(.A(new_n15084), .B(new_n15082_1), .Y(new_n15085));
  or_5   g12737(.A(new_n15084), .B(new_n15082_1), .Y(new_n15086));
  nand_5 g12738(.A(new_n15040), .B(new_n15039), .Y(new_n15087));
  xor_4  g12739(.A(new_n15087), .B(new_n15042), .Y(new_n15088));
  nand_5 g12740(.A(new_n15088), .B(new_n5873), .Y(new_n15089));
  or_5   g12741(.A(new_n15088), .B(new_n5873), .Y(new_n15090));
  nand_5 g12742(.A(new_n9671), .B(new_n9662), .Y(new_n15091));
  nand_5 g12743(.A(new_n15091), .B(new_n9670), .Y(new_n15092));
  nand_5 g12744(.A(new_n15092), .B(new_n15090), .Y(new_n15093));
  nand_5 g12745(.A(new_n15093), .B(new_n15089), .Y(new_n15094_1));
  nand_5 g12746(.A(new_n15094_1), .B(new_n15086), .Y(new_n15095));
  nand_5 g12747(.A(new_n15095), .B(new_n15085), .Y(new_n15096));
  nand_5 g12748(.A(new_n15096), .B(new_n15080), .Y(new_n15097));
  nand_5 g12749(.A(new_n15097), .B(new_n15079), .Y(new_n15098));
  nand_5 g12750(.A(new_n15098), .B(new_n15074), .Y(new_n15099));
  nand_5 g12751(.A(new_n15099), .B(new_n15073), .Y(new_n15100));
  nand_5 g12752(.A(new_n15100), .B(new_n15068), .Y(new_n15101));
  nand_5 g12753(.A(new_n15101), .B(new_n15067), .Y(new_n15102));
  nor_5  g12754(.A(new_n15102), .B(new_n15062), .Y(new_n15103));
  nor_5  g12755(.A(new_n15103), .B(new_n15060), .Y(new_n15104));
  xor_4  g12756(.A(new_n15104), .B(new_n15057), .Y(n2535));
  nand_5 g12757(.A(new_n5544), .B(new_n5549), .Y(new_n15106));
  nand_5 g12758(.A(n20259), .B(n3925), .Y(new_n15107));
  and_5  g12759(.A(new_n15107), .B(new_n15106), .Y(new_n15108));
  nand_5 g12760(.A(new_n15108), .B(n16994), .Y(new_n15109));
  nand_5 g12761(.A(new_n15109), .B(new_n11252), .Y(new_n15110));
  or_5   g12762(.A(new_n15108), .B(n16994), .Y(new_n15111));
  nand_5 g12763(.A(new_n15111), .B(new_n15110), .Y(new_n15112));
  xor_4  g12764(.A(new_n15106), .B(n25872), .Y(new_n15113));
  nand_5 g12765(.A(new_n15113), .B(n10096), .Y(new_n15114));
  nand_5 g12766(.A(new_n15114), .B(new_n15112), .Y(new_n15115));
  nor_5  g12767(.A(new_n15113), .B(n10096), .Y(new_n15116));
  not_8  g12768(.A(new_n15116), .Y(new_n15117));
  nand_5 g12769(.A(new_n15117), .B(new_n15115), .Y(new_n15118_1));
  or_5   g12770(.A(new_n15106), .B(n25872), .Y(new_n15119));
  xor_4  g12771(.A(new_n15119), .B(n7305), .Y(new_n15120));
  nand_5 g12772(.A(new_n15120), .B(n14790), .Y(new_n15121));
  or_5   g12773(.A(new_n15120), .B(n14790), .Y(new_n15122));
  nand_5 g12774(.A(new_n15122), .B(new_n15121), .Y(new_n15123));
  xor_4  g12775(.A(new_n15123), .B(new_n15118_1), .Y(new_n15124));
  or_5   g12776(.A(new_n15124), .B(new_n8898), .Y(new_n15125));
  nand_5 g12777(.A(new_n15124), .B(new_n8898), .Y(new_n15126));
  nand_5 g12778(.A(new_n15117), .B(new_n15114), .Y(new_n15127));
  xor_4  g12779(.A(new_n15127), .B(new_n15112), .Y(new_n15128_1));
  or_5   g12780(.A(new_n15128_1), .B(new_n8906), .Y(new_n15129));
  nand_5 g12781(.A(new_n15128_1), .B(new_n8906), .Y(new_n15130));
  not_8  g12782(.A(new_n11252), .Y(new_n15131));
  and_5  g12783(.A(new_n15111), .B(new_n15109), .Y(new_n15132));
  xor_4  g12784(.A(new_n15132), .B(new_n15131), .Y(new_n15133));
  or_5   g12785(.A(new_n15133), .B(new_n8912), .Y(new_n15134));
  nor_5  g12786(.A(new_n11254), .B(new_n11251), .Y(new_n15135));
  not_8  g12787(.A(new_n15135), .Y(new_n15136));
  nand_5 g12788(.A(new_n15133), .B(new_n8912), .Y(new_n15137));
  nand_5 g12789(.A(new_n15137), .B(new_n15136), .Y(new_n15138));
  nand_5 g12790(.A(new_n15138), .B(new_n15134), .Y(new_n15139_1));
  nand_5 g12791(.A(new_n15139_1), .B(new_n15130), .Y(new_n15140));
  nand_5 g12792(.A(new_n15140), .B(new_n15129), .Y(new_n15141));
  nand_5 g12793(.A(new_n15141), .B(new_n15126), .Y(new_n15142));
  nand_5 g12794(.A(new_n15142), .B(new_n15125), .Y(new_n15143));
  nand_5 g12795(.A(new_n15121), .B(new_n15118_1), .Y(new_n15144));
  nand_5 g12796(.A(new_n15144), .B(new_n15122), .Y(new_n15145_1));
  nor_5  g12797(.A(new_n15119), .B(n7305), .Y(new_n15146_1));
  xor_4  g12798(.A(new_n15146_1), .B(new_n5526), .Y(new_n15147));
  nand_5 g12799(.A(new_n15147), .B(n17251), .Y(new_n15148));
  or_5   g12800(.A(new_n15147), .B(n17251), .Y(new_n15149));
  nand_5 g12801(.A(new_n15149), .B(new_n15148), .Y(new_n15150));
  xor_4  g12802(.A(new_n15150), .B(new_n15145_1), .Y(new_n15151));
  or_5   g12803(.A(new_n15151), .B(new_n8890), .Y(new_n15152));
  nand_5 g12804(.A(new_n15151), .B(new_n8890), .Y(new_n15153));
  nand_5 g12805(.A(new_n15153), .B(new_n15152), .Y(new_n15154));
  xor_4  g12806(.A(new_n15154), .B(new_n15143), .Y(new_n15155));
  not_8  g12807(.A(new_n15155), .Y(new_n15156));
  nand_5 g12808(.A(new_n9760), .B(n2409), .Y(new_n15157));
  nand_5 g12809(.A(n7057), .B(new_n8034), .Y(new_n15158));
  nand_5 g12810(.A(n8869), .B(new_n5709), .Y(new_n15159));
  nand_5 g12811(.A(new_n8035), .B(n8381), .Y(new_n15160));
  nand_5 g12812(.A(new_n9765), .B(n10372), .Y(new_n15161));
  nand_5 g12813(.A(n20235), .B(new_n8038), .Y(new_n15162));
  nand_5 g12814(.A(new_n15162), .B(new_n11257), .Y(new_n15163));
  nand_5 g12815(.A(new_n15163), .B(new_n15161), .Y(new_n15164));
  nand_5 g12816(.A(new_n15164), .B(new_n15160), .Y(new_n15165_1));
  nand_5 g12817(.A(new_n15165_1), .B(new_n15159), .Y(new_n15166));
  nand_5 g12818(.A(new_n15166), .B(new_n15158), .Y(new_n15167_1));
  nand_5 g12819(.A(new_n15167_1), .B(new_n15157), .Y(new_n15168));
  nand_5 g12820(.A(n24170), .B(new_n9757), .Y(new_n15169));
  nand_5 g12821(.A(new_n8052_1), .B(n18537), .Y(new_n15170));
  nand_5 g12822(.A(new_n15170), .B(new_n15169), .Y(new_n15171));
  xor_4  g12823(.A(new_n15171), .B(new_n15168), .Y(new_n15172));
  or_5   g12824(.A(new_n15172), .B(new_n15156), .Y(new_n15173));
  nand_5 g12825(.A(new_n15172), .B(new_n15156), .Y(new_n15174));
  nand_5 g12826(.A(new_n15126), .B(new_n15125), .Y(new_n15175));
  xor_4  g12827(.A(new_n15175), .B(new_n15141), .Y(new_n15176_1));
  not_8  g12828(.A(new_n15176_1), .Y(new_n15177));
  nand_5 g12829(.A(new_n15158), .B(new_n15157), .Y(new_n15178));
  xor_4  g12830(.A(new_n15178), .B(new_n15166), .Y(new_n15179));
  or_5   g12831(.A(new_n15179), .B(new_n15177), .Y(new_n15180_1));
  nand_5 g12832(.A(new_n15179), .B(new_n15177), .Y(new_n15181));
  nand_5 g12833(.A(new_n15130), .B(new_n15129), .Y(new_n15182_1));
  xor_4  g12834(.A(new_n15182_1), .B(new_n15139_1), .Y(new_n15183));
  not_8  g12835(.A(new_n15183), .Y(new_n15184));
  nand_5 g12836(.A(new_n15160), .B(new_n15159), .Y(new_n15185));
  xor_4  g12837(.A(new_n15185), .B(new_n15164), .Y(new_n15186));
  or_5   g12838(.A(new_n15186), .B(new_n15184), .Y(new_n15187));
  nand_5 g12839(.A(new_n15186), .B(new_n15184), .Y(new_n15188));
  not_8  g12840(.A(new_n11257), .Y(new_n15189));
  and_5  g12841(.A(new_n15162), .B(new_n15161), .Y(new_n15190));
  xor_4  g12842(.A(new_n15190), .B(new_n15189), .Y(new_n15191));
  or_5   g12843(.A(new_n15191), .B(new_n11260), .Y(new_n15192));
  nand_5 g12844(.A(new_n15137), .B(new_n15134), .Y(new_n15193));
  xor_4  g12845(.A(new_n15193), .B(new_n15135), .Y(new_n15194));
  not_8  g12846(.A(new_n15194), .Y(new_n15195));
  nand_5 g12847(.A(new_n15191), .B(new_n11260), .Y(new_n15196));
  nand_5 g12848(.A(new_n15196), .B(new_n15195), .Y(new_n15197));
  nand_5 g12849(.A(new_n15197), .B(new_n15192), .Y(new_n15198));
  nand_5 g12850(.A(new_n15198), .B(new_n15188), .Y(new_n15199));
  nand_5 g12851(.A(new_n15199), .B(new_n15187), .Y(new_n15200));
  nand_5 g12852(.A(new_n15200), .B(new_n15181), .Y(new_n15201));
  nand_5 g12853(.A(new_n15201), .B(new_n15180_1), .Y(new_n15202));
  nand_5 g12854(.A(new_n15202), .B(new_n15174), .Y(new_n15203));
  nand_5 g12855(.A(new_n15203), .B(new_n15173), .Y(new_n15204));
  nand_5 g12856(.A(new_n15153), .B(new_n15143), .Y(new_n15205_1));
  nand_5 g12857(.A(new_n15205_1), .B(new_n15152), .Y(new_n15206));
  nand_5 g12858(.A(new_n15148), .B(new_n15145_1), .Y(new_n15207));
  nand_5 g12859(.A(new_n15207), .B(new_n15149), .Y(new_n15208));
  nand_5 g12860(.A(new_n15146_1), .B(new_n5526), .Y(new_n15209));
  xor_4  g12861(.A(new_n15209), .B(n22198), .Y(new_n15210));
  or_5   g12862(.A(new_n15210), .B(n21674), .Y(new_n15211));
  nand_5 g12863(.A(new_n15210), .B(n21674), .Y(new_n15212));
  nand_5 g12864(.A(new_n15212), .B(new_n15211), .Y(new_n15213));
  xor_4  g12865(.A(new_n15213), .B(new_n15208), .Y(new_n15214));
  or_5   g12866(.A(new_n15214), .B(new_n8882), .Y(new_n15215));
  nand_5 g12867(.A(new_n15214), .B(new_n8882), .Y(new_n15216));
  nand_5 g12868(.A(new_n15216), .B(new_n15215), .Y(new_n15217));
  xor_4  g12869(.A(new_n15217), .B(new_n15206), .Y(new_n15218));
  nand_5 g12870(.A(new_n15170), .B(new_n15168), .Y(new_n15219));
  nand_5 g12871(.A(new_n15219), .B(new_n15169), .Y(new_n15220));
  not_8  g12872(.A(new_n15220), .Y(new_n15221));
  nand_5 g12873(.A(new_n9778_1), .B(n329), .Y(new_n15222));
  nand_5 g12874(.A(n1163), .B(new_n8031_1), .Y(new_n15223));
  nand_5 g12875(.A(new_n15223), .B(new_n15222), .Y(new_n15224));
  xor_4  g12876(.A(new_n15224), .B(new_n15221), .Y(new_n15225));
  nand_5 g12877(.A(new_n15225), .B(new_n15218), .Y(new_n15226));
  not_8  g12878(.A(new_n15218), .Y(new_n15227));
  not_8  g12879(.A(new_n15225), .Y(new_n15228));
  nand_5 g12880(.A(new_n15228), .B(new_n15227), .Y(new_n15229));
  nand_5 g12881(.A(new_n15229), .B(new_n15226), .Y(new_n15230_1));
  xnor_4 g12882(.A(new_n15230_1), .B(new_n15204), .Y(n2537));
  nand_5 g12883(.A(new_n4724), .B(new_n3139), .Y(new_n15232));
  nand_5 g12884(.A(new_n4723), .B(new_n3138), .Y(new_n15233));
  nand_5 g12885(.A(new_n4683), .B(new_n3146), .Y(new_n15234));
  nand_5 g12886(.A(new_n4682), .B(new_n3148), .Y(new_n15235));
  nand_5 g12887(.A(new_n4673), .B(new_n3154), .Y(new_n15236));
  nand_5 g12888(.A(new_n4672), .B(new_n3156), .Y(new_n15237));
  nand_5 g12889(.A(new_n3166), .B(new_n3248), .Y(new_n15238));
  not_8  g12890(.A(new_n15238), .Y(new_n15239));
  nand_5 g12891(.A(new_n15239), .B(new_n15237), .Y(new_n15240));
  nand_5 g12892(.A(new_n15240), .B(new_n15236), .Y(new_n15241_1));
  nand_5 g12893(.A(new_n15241_1), .B(new_n15235), .Y(new_n15242));
  nand_5 g12894(.A(new_n15242), .B(new_n15234), .Y(new_n15243));
  nand_5 g12895(.A(new_n15243), .B(new_n15233), .Y(new_n15244));
  nand_5 g12896(.A(new_n15244), .B(new_n15232), .Y(new_n15245));
  nand_5 g12897(.A(new_n4796), .B(new_n3130), .Y(new_n15246));
  nand_5 g12898(.A(new_n4795), .B(new_n3129), .Y(new_n15247));
  nand_5 g12899(.A(new_n15247), .B(new_n15246), .Y(new_n15248));
  xor_4  g12900(.A(new_n15248), .B(new_n15245), .Y(new_n15249));
  nand_5 g12901(.A(new_n15249), .B(new_n11078_1), .Y(new_n15250));
  or_5   g12902(.A(new_n15249), .B(new_n11078_1), .Y(new_n15251));
  nand_5 g12903(.A(new_n15232), .B(new_n15233), .Y(new_n15252));
  xor_4  g12904(.A(new_n15252), .B(new_n15243), .Y(new_n15253));
  or_5   g12905(.A(new_n15253), .B(new_n11026), .Y(new_n15254));
  nand_5 g12906(.A(new_n15253), .B(new_n11026), .Y(new_n15255_1));
  nand_5 g12907(.A(new_n15234), .B(new_n15235), .Y(new_n15256));
  xor_4  g12908(.A(new_n15256), .B(new_n15241_1), .Y(new_n15257));
  or_5   g12909(.A(new_n15257), .B(new_n10995), .Y(new_n15258_1));
  nand_5 g12910(.A(new_n15257), .B(new_n10995), .Y(new_n15259));
  nand_5 g12911(.A(new_n15236), .B(new_n15237), .Y(new_n15260));
  xor_4  g12912(.A(new_n15260), .B(new_n15239), .Y(new_n15261));
  or_5   g12913(.A(new_n15261), .B(new_n11011_1), .Y(new_n15262));
  nand_5 g12914(.A(new_n15261), .B(new_n11011_1), .Y(new_n15263));
  nand_5 g12915(.A(new_n3244_1), .B(n1152), .Y(new_n15264));
  nand_5 g12916(.A(new_n15264), .B(new_n15238), .Y(new_n15265));
  nand_5 g12917(.A(new_n15265), .B(new_n8282), .Y(new_n15266));
  nand_5 g12918(.A(new_n15266), .B(new_n15263), .Y(new_n15267));
  nand_5 g12919(.A(new_n15267), .B(new_n15262), .Y(new_n15268));
  nand_5 g12920(.A(new_n15268), .B(new_n15259), .Y(new_n15269));
  nand_5 g12921(.A(new_n15269), .B(new_n15258_1), .Y(new_n15270));
  nand_5 g12922(.A(new_n15270), .B(new_n15255_1), .Y(new_n15271_1));
  and_5  g12923(.A(new_n15271_1), .B(new_n15254), .Y(new_n15272));
  nand_5 g12924(.A(new_n15272), .B(new_n15251), .Y(new_n15273));
  nand_5 g12925(.A(new_n15273), .B(new_n15250), .Y(new_n15274));
  not_8  g12926(.A(new_n13202), .Y(new_n15275_1));
  nand_5 g12927(.A(new_n15247), .B(new_n15245), .Y(new_n15276));
  nand_5 g12928(.A(new_n15276), .B(new_n15246), .Y(new_n15277));
  nand_5 g12929(.A(new_n12716), .B(new_n3122), .Y(new_n15278));
  nand_5 g12930(.A(new_n12715), .B(new_n3121), .Y(new_n15279));
  nand_5 g12931(.A(new_n15279), .B(new_n15278), .Y(new_n15280));
  xnor_4 g12932(.A(new_n15280), .B(new_n15277), .Y(new_n15281));
  or_5   g12933(.A(new_n15281), .B(new_n15275_1), .Y(new_n15282));
  nand_5 g12934(.A(new_n15281), .B(new_n15275_1), .Y(new_n15283));
  nand_5 g12935(.A(new_n15283), .B(new_n15282), .Y(new_n15284));
  xnor_4 g12936(.A(new_n15284), .B(new_n15274), .Y(n2553));
  nand_5 g12937(.A(new_n13700), .B(new_n13699), .Y(new_n15286));
  xnor_4 g12938(.A(new_n15286), .B(new_n13725), .Y(n2555));
  nand_5 g12939(.A(new_n12444), .B(n12892), .Y(new_n15288));
  or_5   g12940(.A(new_n12444), .B(n12892), .Y(new_n15289_1));
  and_5  g12941(.A(new_n15289_1), .B(new_n15288), .Y(new_n15290));
  nand_5 g12942(.A(new_n15290), .B(new_n11600), .Y(new_n15291));
  not_8  g12943(.A(new_n15291), .Y(new_n15292));
  not_8  g12944(.A(n12209), .Y(new_n15293));
  or_5   g12945(.A(new_n12338), .B(new_n15293), .Y(new_n15294));
  nand_5 g12946(.A(new_n12338), .B(new_n15293), .Y(new_n15295));
  nand_5 g12947(.A(new_n15295), .B(new_n15294), .Y(new_n15296));
  xor_4  g12948(.A(new_n15296), .B(new_n15288), .Y(new_n15297));
  not_8  g12949(.A(new_n15297), .Y(new_n15298));
  or_5   g12950(.A(new_n15298), .B(new_n11593), .Y(new_n15299));
  nand_5 g12951(.A(new_n15298), .B(new_n11593), .Y(new_n15300_1));
  nand_5 g12952(.A(new_n15300_1), .B(new_n15299), .Y(new_n15301));
  xor_4  g12953(.A(new_n15301), .B(new_n15292), .Y(n2560));
  nand_5 g12954(.A(new_n3909_1), .B(new_n14514), .Y(new_n15303));
  nand_5 g12955(.A(n26180), .B(n10650), .Y(new_n15304));
  nand_5 g12956(.A(new_n3915), .B(new_n14517), .Y(new_n15305));
  nand_5 g12957(.A(n24004), .B(n12900), .Y(new_n15306));
  nand_5 g12958(.A(new_n14520), .B(new_n3921), .Y(new_n15307_1));
  nand_5 g12959(.A(n20411), .B(n12871), .Y(new_n15308));
  nand_5 g12960(.A(new_n3927), .B(new_n14523), .Y(new_n15309));
  nand_5 g12961(.A(n23304), .B(n17069), .Y(new_n15310));
  nand_5 g12962(.A(new_n3957), .B(new_n14538), .Y(new_n15311));
  nand_5 g12963(.A(n8721), .B(n1040), .Y(new_n15312));
  nand_5 g12964(.A(n18578), .B(n9090), .Y(new_n15313));
  nand_5 g12965(.A(new_n15313), .B(new_n15312), .Y(new_n15314));
  nand_5 g12966(.A(new_n15314), .B(new_n15311), .Y(new_n15315));
  nand_5 g12967(.A(new_n15315), .B(new_n14535), .Y(new_n15316));
  not_8  g12968(.A(new_n15316), .Y(new_n15317));
  nor_5  g12969(.A(new_n15315), .B(new_n14535), .Y(new_n15318));
  nor_5  g12970(.A(new_n15318), .B(n14633), .Y(new_n15319));
  nor_5  g12971(.A(new_n15319), .B(new_n15317), .Y(new_n15320));
  or_5   g12972(.A(new_n15320), .B(n4722), .Y(new_n15321));
  nand_5 g12973(.A(new_n15320), .B(n4722), .Y(new_n15322));
  nand_5 g12974(.A(new_n15322), .B(new_n14532), .Y(new_n15323));
  nand_5 g12975(.A(new_n15323), .B(new_n15321), .Y(new_n15324));
  nand_5 g12976(.A(new_n15324), .B(new_n3939), .Y(new_n15325));
  not_8  g12977(.A(new_n15325), .Y(new_n15326));
  nor_5  g12978(.A(new_n15324), .B(new_n3939), .Y(new_n15327_1));
  nor_5  g12979(.A(new_n15327_1), .B(n17784), .Y(new_n15328));
  nor_5  g12980(.A(new_n15328), .B(new_n15326), .Y(new_n15329));
  or_5   g12981(.A(new_n15329), .B(n15918), .Y(new_n15330));
  nand_5 g12982(.A(new_n15329), .B(n15918), .Y(new_n15331));
  nand_5 g12983(.A(new_n15331), .B(new_n3933), .Y(new_n15332_1));
  nand_5 g12984(.A(new_n15332_1), .B(new_n15330), .Y(new_n15333));
  nand_5 g12985(.A(new_n15333), .B(new_n15310), .Y(new_n15334));
  nand_5 g12986(.A(new_n15334), .B(new_n15309), .Y(new_n15335));
  nand_5 g12987(.A(new_n15335), .B(new_n15308), .Y(new_n15336));
  nand_5 g12988(.A(new_n15336), .B(new_n15307_1), .Y(new_n15337));
  nand_5 g12989(.A(new_n15337), .B(new_n15306), .Y(new_n15338));
  nand_5 g12990(.A(new_n15338), .B(new_n15305), .Y(new_n15339));
  nand_5 g12991(.A(new_n15339), .B(new_n15304), .Y(new_n15340));
  nand_5 g12992(.A(new_n15340), .B(new_n15303), .Y(new_n15341));
  nand_5 g12993(.A(new_n6707_1), .B(new_n6662), .Y(new_n15342));
  nand_5 g12994(.A(new_n15342), .B(new_n6664), .Y(new_n15343));
  not_8  g12995(.A(new_n15343), .Y(new_n15344));
  or_5   g12996(.A(new_n15344), .B(new_n15341), .Y(new_n15345_1));
  nand_5 g12997(.A(new_n15344), .B(new_n15341), .Y(new_n15346));
  nand_5 g12998(.A(new_n15304), .B(new_n15303), .Y(new_n15347));
  xor_4  g12999(.A(new_n15347), .B(new_n15339), .Y(new_n15348));
  nand_5 g13000(.A(new_n15348), .B(new_n6709), .Y(new_n15349));
  not_8  g13001(.A(new_n15349), .Y(new_n15350));
  not_8  g13002(.A(new_n15348), .Y(new_n15351));
  nand_5 g13003(.A(new_n15351), .B(new_n6708), .Y(new_n15352));
  not_8  g13004(.A(new_n15352), .Y(new_n15353_1));
  nand_5 g13005(.A(new_n15306), .B(new_n15305), .Y(new_n15354));
  xnor_4 g13006(.A(new_n15354), .B(new_n15337), .Y(new_n15355));
  nand_5 g13007(.A(new_n15355), .B(new_n6717), .Y(new_n15356));
  or_5   g13008(.A(new_n15355), .B(new_n6717), .Y(new_n15357));
  nand_5 g13009(.A(new_n15308), .B(new_n15307_1), .Y(new_n15358));
  xor_4  g13010(.A(new_n15358), .B(new_n15335), .Y(new_n15359));
  or_5   g13011(.A(new_n15359), .B(new_n6726), .Y(new_n15360));
  nand_5 g13012(.A(new_n15359), .B(new_n6726), .Y(new_n15361));
  nand_5 g13013(.A(new_n15310), .B(new_n15309), .Y(new_n15362));
  xnor_4 g13014(.A(new_n15362), .B(new_n15333), .Y(new_n15363));
  nand_5 g13015(.A(new_n15363), .B(new_n6731), .Y(new_n15364));
  or_5   g13016(.A(new_n15363), .B(new_n6731), .Y(new_n15365));
  and_5  g13017(.A(new_n15331), .B(new_n15330), .Y(new_n15366_1));
  xor_4  g13018(.A(new_n15366_1), .B(new_n3933), .Y(new_n15367));
  nand_5 g13019(.A(new_n15367), .B(new_n6738), .Y(new_n15368));
  or_5   g13020(.A(new_n15367), .B(new_n6738), .Y(new_n15369));
  nor_5  g13021(.A(new_n15327_1), .B(new_n15326), .Y(new_n15370));
  xor_4  g13022(.A(new_n15370), .B(n17784), .Y(new_n15371));
  or_5   g13023(.A(new_n15371), .B(new_n6745), .Y(new_n15372));
  nand_5 g13024(.A(new_n15371), .B(new_n6745), .Y(new_n15373));
  and_5  g13025(.A(new_n15322), .B(new_n15321), .Y(new_n15374));
  xor_4  g13026(.A(new_n15374), .B(new_n14532), .Y(new_n15375));
  nand_5 g13027(.A(new_n15375), .B(new_n6753), .Y(new_n15376));
  or_5   g13028(.A(new_n15375), .B(new_n6753), .Y(new_n15377));
  nor_5  g13029(.A(new_n15318), .B(new_n15317), .Y(new_n15378_1));
  xor_4  g13030(.A(new_n15378_1), .B(new_n3951), .Y(new_n15379));
  nand_5 g13031(.A(new_n15379), .B(new_n6760), .Y(new_n15380));
  or_5   g13032(.A(new_n15379), .B(new_n6760), .Y(new_n15381));
  not_8  g13033(.A(new_n15313), .Y(new_n15382_1));
  nor_5  g13034(.A(n18578), .B(n9090), .Y(new_n15383));
  or_5   g13035(.A(new_n15383), .B(new_n15382_1), .Y(new_n15384));
  nand_5 g13036(.A(new_n15384), .B(new_n6767), .Y(new_n15385));
  nand_5 g13037(.A(new_n15385), .B(new_n6774), .Y(new_n15386));
  nand_5 g13038(.A(new_n15312), .B(new_n15311), .Y(new_n15387));
  xor_4  g13039(.A(new_n15387), .B(new_n15382_1), .Y(new_n15388));
  nand_5 g13040(.A(new_n15388), .B(new_n15386), .Y(new_n15389));
  or_5   g13041(.A(new_n15385), .B(new_n6772), .Y(new_n15390));
  nand_5 g13042(.A(new_n15390), .B(new_n15389), .Y(new_n15391));
  nand_5 g13043(.A(new_n15391), .B(new_n15381), .Y(new_n15392));
  nand_5 g13044(.A(new_n15392), .B(new_n15380), .Y(new_n15393));
  nand_5 g13045(.A(new_n15393), .B(new_n15377), .Y(new_n15394));
  nand_5 g13046(.A(new_n15394), .B(new_n15376), .Y(new_n15395));
  nand_5 g13047(.A(new_n15395), .B(new_n15373), .Y(new_n15396));
  nand_5 g13048(.A(new_n15396), .B(new_n15372), .Y(new_n15397));
  nand_5 g13049(.A(new_n15397), .B(new_n15369), .Y(new_n15398));
  nand_5 g13050(.A(new_n15398), .B(new_n15368), .Y(new_n15399));
  nand_5 g13051(.A(new_n15399), .B(new_n15365), .Y(new_n15400));
  nand_5 g13052(.A(new_n15400), .B(new_n15364), .Y(new_n15401));
  nand_5 g13053(.A(new_n15401), .B(new_n15361), .Y(new_n15402));
  nand_5 g13054(.A(new_n15402), .B(new_n15360), .Y(new_n15403));
  nand_5 g13055(.A(new_n15403), .B(new_n15357), .Y(new_n15404));
  nand_5 g13056(.A(new_n15404), .B(new_n15356), .Y(new_n15405));
  nor_5  g13057(.A(new_n15405), .B(new_n15353_1), .Y(new_n15406));
  nor_5  g13058(.A(new_n15406), .B(new_n15350), .Y(new_n15407_1));
  not_8  g13059(.A(new_n15407_1), .Y(new_n15408));
  nand_5 g13060(.A(new_n15408), .B(new_n15346), .Y(new_n15409));
  nand_5 g13061(.A(new_n15409), .B(new_n15345_1), .Y(new_n15410));
  nand_5 g13062(.A(new_n15346), .B(new_n15345_1), .Y(new_n15411));
  xor_4  g13063(.A(new_n15411), .B(new_n15407_1), .Y(new_n15412));
  nand_5 g13064(.A(new_n3765), .B(new_n3714), .Y(new_n15413));
  nand_5 g13065(.A(new_n15413), .B(new_n3712), .Y(new_n15414));
  or_5   g13066(.A(new_n15414), .B(new_n15412), .Y(new_n15415));
  nand_5 g13067(.A(new_n15414), .B(new_n15412), .Y(new_n15416));
  nand_5 g13068(.A(new_n15352), .B(new_n15349), .Y(new_n15417));
  xor_4  g13069(.A(new_n15417), .B(new_n15405), .Y(new_n15418));
  or_5   g13070(.A(new_n15418), .B(new_n3770), .Y(new_n15419));
  not_8  g13071(.A(new_n15419), .Y(new_n15420));
  nand_5 g13072(.A(new_n15418), .B(new_n3770), .Y(new_n15421));
  not_8  g13073(.A(new_n15421), .Y(new_n15422));
  nand_5 g13074(.A(new_n15356), .B(new_n15357), .Y(new_n15423));
  xor_4  g13075(.A(new_n15423), .B(new_n15403), .Y(new_n15424_1));
  nand_5 g13076(.A(new_n15424_1), .B(new_n3775), .Y(new_n15425));
  or_5   g13077(.A(new_n15424_1), .B(new_n3775), .Y(new_n15426));
  nand_5 g13078(.A(new_n15361), .B(new_n15360), .Y(new_n15427));
  xor_4  g13079(.A(new_n15427), .B(new_n15401), .Y(new_n15428_1));
  nand_5 g13080(.A(new_n15428_1), .B(new_n3781_1), .Y(new_n15429));
  or_5   g13081(.A(new_n15428_1), .B(new_n3781_1), .Y(new_n15430));
  nand_5 g13082(.A(new_n15365), .B(new_n15364), .Y(new_n15431));
  xnor_4 g13083(.A(new_n15431), .B(new_n15399), .Y(new_n15432));
  or_5   g13084(.A(new_n15432), .B(new_n3791), .Y(new_n15433));
  nand_5 g13085(.A(new_n15432), .B(new_n3791), .Y(new_n15434));
  nand_5 g13086(.A(new_n15369), .B(new_n15368), .Y(new_n15435_1));
  xor_4  g13087(.A(new_n15435_1), .B(new_n15397), .Y(new_n15436));
  nand_5 g13088(.A(new_n15436), .B(new_n3796), .Y(new_n15437));
  or_5   g13089(.A(new_n15436), .B(new_n3796), .Y(new_n15438_1));
  nand_5 g13090(.A(new_n15373), .B(new_n15372), .Y(new_n15439));
  xor_4  g13091(.A(new_n15439), .B(new_n15395), .Y(new_n15440));
  nand_5 g13092(.A(new_n15440), .B(new_n3802), .Y(new_n15441));
  or_5   g13093(.A(new_n15440), .B(new_n3802), .Y(new_n15442));
  nand_5 g13094(.A(new_n15377), .B(new_n15376), .Y(new_n15443));
  xor_4  g13095(.A(new_n15443), .B(new_n15393), .Y(new_n15444));
  nand_5 g13096(.A(new_n15444), .B(new_n3808), .Y(new_n15445));
  or_5   g13097(.A(new_n15444), .B(new_n3808), .Y(new_n15446));
  nand_5 g13098(.A(new_n15381), .B(new_n15380), .Y(new_n15447));
  xor_4  g13099(.A(new_n15447), .B(new_n15391), .Y(new_n15448));
  nand_5 g13100(.A(new_n15448), .B(new_n3815), .Y(new_n15449));
  or_5   g13101(.A(new_n15448), .B(new_n3815), .Y(new_n15450));
  nand_5 g13102(.A(new_n15390), .B(new_n15386), .Y(new_n15451));
  xor_4  g13103(.A(new_n15451), .B(new_n15388), .Y(new_n15452));
  nand_5 g13104(.A(new_n15452), .B(new_n3824), .Y(new_n15453));
  or_5   g13105(.A(new_n15452), .B(new_n3824), .Y(new_n15454));
  xor_4  g13106(.A(new_n15384), .B(new_n6767), .Y(new_n15455));
  nand_5 g13107(.A(new_n15455), .B(new_n3830), .Y(new_n15456));
  nand_5 g13108(.A(new_n15456), .B(new_n15454), .Y(new_n15457));
  nand_5 g13109(.A(new_n15457), .B(new_n15453), .Y(new_n15458));
  nand_5 g13110(.A(new_n15458), .B(new_n15450), .Y(new_n15459));
  nand_5 g13111(.A(new_n15459), .B(new_n15449), .Y(new_n15460));
  nand_5 g13112(.A(new_n15460), .B(new_n15446), .Y(new_n15461));
  nand_5 g13113(.A(new_n15461), .B(new_n15445), .Y(new_n15462));
  nand_5 g13114(.A(new_n15462), .B(new_n15442), .Y(new_n15463));
  nand_5 g13115(.A(new_n15463), .B(new_n15441), .Y(new_n15464));
  nand_5 g13116(.A(new_n15464), .B(new_n15438_1), .Y(new_n15465_1));
  nand_5 g13117(.A(new_n15465_1), .B(new_n15437), .Y(new_n15466));
  nand_5 g13118(.A(new_n15466), .B(new_n15434), .Y(new_n15467_1));
  nand_5 g13119(.A(new_n15467_1), .B(new_n15433), .Y(new_n15468));
  nand_5 g13120(.A(new_n15468), .B(new_n15430), .Y(new_n15469));
  nand_5 g13121(.A(new_n15469), .B(new_n15429), .Y(new_n15470_1));
  nand_5 g13122(.A(new_n15470_1), .B(new_n15426), .Y(new_n15471));
  nand_5 g13123(.A(new_n15471), .B(new_n15425), .Y(new_n15472));
  nor_5  g13124(.A(new_n15472), .B(new_n15422), .Y(new_n15473));
  nor_5  g13125(.A(new_n15473), .B(new_n15420), .Y(new_n15474));
  not_8  g13126(.A(new_n15474), .Y(new_n15475));
  nand_5 g13127(.A(new_n15475), .B(new_n15416), .Y(new_n15476));
  nand_5 g13128(.A(new_n15476), .B(new_n15415), .Y(new_n15477_1));
  not_8  g13129(.A(new_n15477_1), .Y(new_n15478));
  xor_4  g13130(.A(new_n15478), .B(new_n15410), .Y(n2561));
  nand_5 g13131(.A(new_n9652), .B(new_n9653), .Y(new_n15480));
  xnor_4 g13132(.A(new_n15480), .B(new_n9655_1), .Y(n2573));
  nand_5 g13133(.A(n18151), .B(new_n3248), .Y(new_n15482));
  nand_5 g13134(.A(new_n2770), .B(n1152), .Y(new_n15483));
  and_5  g13135(.A(new_n15483), .B(new_n15482), .Y(new_n15484));
  not_8  g13136(.A(new_n15484), .Y(new_n15485));
  nand_5 g13137(.A(new_n15485), .B(new_n11498), .Y(new_n15486));
  nand_5 g13138(.A(n14148), .B(new_n2769), .Y(new_n15487));
  nand_5 g13139(.A(new_n2809_1), .B(n11503), .Y(new_n15488));
  nand_5 g13140(.A(new_n15488), .B(new_n15487), .Y(new_n15489));
  xor_4  g13141(.A(new_n15489), .B(new_n15482), .Y(new_n15490_1));
  or_5   g13142(.A(new_n15490_1), .B(new_n15486), .Y(new_n15491));
  nand_5 g13143(.A(new_n15490_1), .B(new_n15486), .Y(new_n15492));
  xor_4  g13144(.A(new_n11494), .B(new_n11490), .Y(new_n15493));
  nand_5 g13145(.A(new_n15493), .B(new_n15492), .Y(new_n15494));
  nand_5 g13146(.A(new_n15494), .B(new_n15491), .Y(new_n15495));
  nand_5 g13147(.A(n20349), .B(new_n9126), .Y(new_n15496_1));
  nand_5 g13148(.A(new_n15496_1), .B(new_n11494), .Y(new_n15497));
  nand_5 g13149(.A(new_n11424_1), .B(n10017), .Y(new_n15498));
  nand_5 g13150(.A(new_n15498), .B(new_n15497), .Y(new_n15499));
  xor_4  g13151(.A(new_n15499), .B(new_n11485), .Y(new_n15500));
  nand_5 g13152(.A(new_n15488), .B(new_n15482), .Y(new_n15501_1));
  nand_5 g13153(.A(new_n15501_1), .B(new_n15487), .Y(new_n15502));
  nand_5 g13154(.A(new_n11718), .B(n7149), .Y(new_n15503));
  nand_5 g13155(.A(n16971), .B(new_n2805), .Y(new_n15504));
  nand_5 g13156(.A(new_n15504), .B(new_n15503), .Y(new_n15505));
  xor_4  g13157(.A(new_n15505), .B(new_n15502), .Y(new_n15506_1));
  not_8  g13158(.A(new_n15506_1), .Y(new_n15507));
  nand_5 g13159(.A(new_n15507), .B(new_n15500), .Y(new_n15508_1));
  not_8  g13160(.A(new_n15500), .Y(new_n15509));
  nand_5 g13161(.A(new_n15506_1), .B(new_n15509), .Y(new_n15510));
  nand_5 g13162(.A(new_n15510), .B(new_n15508_1), .Y(new_n15511));
  xor_4  g13163(.A(new_n15511), .B(new_n15495), .Y(new_n15512));
  nand_5 g13164(.A(new_n15293), .B(n6631), .Y(new_n15513));
  nand_5 g13165(.A(n12209), .B(new_n4621), .Y(new_n15514));
  nand_5 g13166(.A(new_n4622), .B(n12892), .Y(new_n15515));
  nand_5 g13167(.A(new_n15515), .B(new_n15514), .Y(new_n15516));
  nand_5 g13168(.A(new_n15516), .B(new_n15513), .Y(new_n15517));
  not_8  g13169(.A(n22588), .Y(new_n15518));
  nand_5 g13170(.A(new_n15518), .B(n14684), .Y(new_n15519));
  nand_5 g13171(.A(n22588), .B(new_n4620), .Y(new_n15520));
  nand_5 g13172(.A(new_n15520), .B(new_n15519), .Y(new_n15521));
  xor_4  g13173(.A(new_n15521), .B(new_n15517), .Y(new_n15522));
  nand_5 g13174(.A(new_n15522), .B(new_n15512), .Y(new_n15523));
  not_8  g13175(.A(new_n15512), .Y(new_n15524));
  not_8  g13176(.A(new_n15522), .Y(new_n15525));
  nand_5 g13177(.A(new_n15525), .B(new_n15524), .Y(new_n15526));
  nand_5 g13178(.A(new_n15484), .B(new_n11497), .Y(new_n15527));
  nand_5 g13179(.A(new_n15527), .B(new_n15486), .Y(new_n15528));
  not_8  g13180(.A(new_n15528), .Y(new_n15529));
  not_8  g13181(.A(new_n15515), .Y(new_n15530));
  nor_5  g13182(.A(new_n4622), .B(n12892), .Y(new_n15531));
  or_5   g13183(.A(new_n15531), .B(new_n15530), .Y(new_n15532));
  nand_5 g13184(.A(new_n15532), .B(new_n15529), .Y(new_n15533));
  nand_5 g13185(.A(new_n15514), .B(new_n15513), .Y(new_n15534));
  xor_4  g13186(.A(new_n15534), .B(new_n15515), .Y(new_n15535));
  nand_5 g13187(.A(new_n15535), .B(new_n15533), .Y(new_n15536));
  or_5   g13188(.A(new_n15535), .B(new_n15533), .Y(new_n15537));
  nand_5 g13189(.A(new_n15491), .B(new_n15492), .Y(new_n15538));
  xor_4  g13190(.A(new_n15538), .B(new_n15493), .Y(new_n15539_1));
  nand_5 g13191(.A(new_n15539_1), .B(new_n15537), .Y(new_n15540));
  nand_5 g13192(.A(new_n15540), .B(new_n15536), .Y(new_n15541));
  nand_5 g13193(.A(new_n15541), .B(new_n15526), .Y(new_n15542));
  nand_5 g13194(.A(new_n15542), .B(new_n15523), .Y(new_n15543));
  nand_5 g13195(.A(new_n15510), .B(new_n15495), .Y(new_n15544));
  nand_5 g13196(.A(new_n15544), .B(new_n15508_1), .Y(new_n15545));
  nand_5 g13197(.A(new_n9123), .B(n6590), .Y(new_n15546_1));
  nand_5 g13198(.A(new_n15546_1), .B(new_n15499), .Y(new_n15547));
  nand_5 g13199(.A(n7963), .B(new_n11421), .Y(new_n15548));
  nand_5 g13200(.A(new_n15548), .B(new_n15547), .Y(new_n15549));
  xor_4  g13201(.A(new_n15549), .B(new_n11480), .Y(new_n15550));
  nand_5 g13202(.A(new_n15504), .B(new_n15502), .Y(new_n15551));
  nand_5 g13203(.A(new_n15551), .B(new_n15503), .Y(new_n15552));
  not_8  g13204(.A(new_n15552), .Y(new_n15553));
  nand_5 g13205(.A(n18558), .B(new_n2876), .Y(new_n15554));
  nand_5 g13206(.A(new_n2872), .B(n10411), .Y(new_n15555_1));
  nand_5 g13207(.A(new_n15555_1), .B(new_n15554), .Y(new_n15556));
  xor_4  g13208(.A(new_n15556), .B(new_n15553), .Y(new_n15557));
  nand_5 g13209(.A(new_n15557), .B(new_n15550), .Y(new_n15558_1));
  not_8  g13210(.A(new_n15550), .Y(new_n15559_1));
  not_8  g13211(.A(new_n15557), .Y(new_n15560));
  nand_5 g13212(.A(new_n15560), .B(new_n15559_1), .Y(new_n15561));
  nand_5 g13213(.A(new_n15561), .B(new_n15558_1), .Y(new_n15562));
  xor_4  g13214(.A(new_n15562), .B(new_n15545), .Y(new_n15563));
  nand_5 g13215(.A(new_n15520), .B(new_n15517), .Y(new_n15564));
  nand_5 g13216(.A(new_n15564), .B(new_n15519), .Y(new_n15565));
  not_8  g13217(.A(new_n15565), .Y(new_n15566));
  not_8  g13218(.A(n19515), .Y(new_n15567));
  nand_5 g13219(.A(new_n15567), .B(n17035), .Y(new_n15568));
  nand_5 g13220(.A(n19515), .B(new_n4642), .Y(new_n15569));
  nand_5 g13221(.A(new_n15569), .B(new_n15568), .Y(new_n15570_1));
  xor_4  g13222(.A(new_n15570_1), .B(new_n15566), .Y(new_n15571));
  not_8  g13223(.A(new_n15571), .Y(new_n15572));
  nand_5 g13224(.A(new_n15572), .B(new_n15563), .Y(new_n15573_1));
  not_8  g13225(.A(new_n15563), .Y(new_n15574));
  nand_5 g13226(.A(new_n15571), .B(new_n15574), .Y(new_n15575));
  nand_5 g13227(.A(new_n15575), .B(new_n15573_1), .Y(new_n15576));
  xor_4  g13228(.A(new_n15576), .B(new_n15543), .Y(n2578));
  nor_5  g13229(.A(new_n13531), .B(new_n9009), .Y(new_n15578));
  xor_4  g13230(.A(new_n13531), .B(new_n9011), .Y(new_n15579));
  nand_5 g13231(.A(new_n9102), .B(new_n9010), .Y(new_n15580));
  nand_5 g13232(.A(new_n15580), .B(new_n9012_1), .Y(new_n15581));
  nor_5  g13233(.A(new_n15581), .B(new_n15579), .Y(new_n15582));
  nor_5  g13234(.A(new_n15582), .B(new_n15578), .Y(n2582));
  nand_5 g13235(.A(new_n4743), .B(new_n4744), .Y(new_n15584));
  xor_4  g13236(.A(new_n15584), .B(new_n4760), .Y(n2602));
  nand_5 g13237(.A(new_n9313), .B(new_n4886), .Y(new_n15586));
  nand_5 g13238(.A(new_n9315), .B(n20250), .Y(new_n15587));
  nand_5 g13239(.A(new_n9319), .B(new_n4892), .Y(new_n15588_1));
  nand_5 g13240(.A(new_n9321), .B(n5822), .Y(new_n15589));
  nand_5 g13241(.A(new_n9326), .B(new_n4898), .Y(new_n15590_1));
  nand_5 g13242(.A(new_n9325), .B(n26443), .Y(new_n15591));
  nand_5 g13243(.A(new_n9328), .B(n1681), .Y(new_n15592));
  nand_5 g13244(.A(new_n15592), .B(new_n15591), .Y(new_n15593));
  nand_5 g13245(.A(new_n15593), .B(new_n15590_1), .Y(new_n15594));
  nand_5 g13246(.A(new_n15594), .B(new_n15589), .Y(new_n15595));
  nand_5 g13247(.A(new_n15595), .B(new_n15588_1), .Y(new_n15596));
  nand_5 g13248(.A(new_n15596), .B(new_n15587), .Y(new_n15597));
  nand_5 g13249(.A(new_n15597), .B(new_n15586), .Y(new_n15598_1));
  nand_5 g13250(.A(new_n9307), .B(new_n4880), .Y(new_n15599));
  nand_5 g13251(.A(new_n9309), .B(n3785), .Y(new_n15600));
  nand_5 g13252(.A(new_n15600), .B(new_n15599), .Y(new_n15601));
  xnor_4 g13253(.A(new_n15601), .B(new_n15598_1), .Y(new_n15602_1));
  nand_5 g13254(.A(new_n2619_1), .B(new_n9323_1), .Y(new_n15603));
  or_5   g13255(.A(new_n15603), .B(n24485), .Y(new_n15604));
  nor_5  g13256(.A(new_n15604), .B(n21078), .Y(new_n15605));
  not_8  g13257(.A(new_n15605), .Y(new_n15606));
  nand_5 g13258(.A(new_n15604), .B(n21078), .Y(new_n15607));
  nand_5 g13259(.A(new_n15607), .B(new_n15606), .Y(new_n15608));
  nand_5 g13260(.A(new_n15608), .B(new_n4336), .Y(new_n15609));
  or_5   g13261(.A(new_n15608), .B(new_n4336), .Y(new_n15610));
  nand_5 g13262(.A(new_n15603), .B(n24485), .Y(new_n15611));
  and_5  g13263(.A(new_n15611), .B(new_n15604), .Y(new_n15612));
  or_5   g13264(.A(new_n15612), .B(new_n4342), .Y(new_n15613));
  nand_5 g13265(.A(new_n15612), .B(new_n4342), .Y(new_n15614_1));
  nand_5 g13266(.A(n22201), .B(n2420), .Y(new_n15615));
  and_5  g13267(.A(new_n15615), .B(new_n15603), .Y(new_n15616));
  or_5   g13268(.A(new_n15616), .B(new_n4351), .Y(new_n15617));
  nand_5 g13269(.A(new_n15616), .B(new_n4351), .Y(new_n15618));
  nand_5 g13270(.A(new_n2634), .B(n22201), .Y(new_n15619));
  nand_5 g13271(.A(new_n15619), .B(new_n15618), .Y(new_n15620));
  nand_5 g13272(.A(new_n15620), .B(new_n15617), .Y(new_n15621));
  nand_5 g13273(.A(new_n15621), .B(new_n15614_1), .Y(new_n15622));
  nand_5 g13274(.A(new_n15622), .B(new_n15613), .Y(new_n15623));
  nand_5 g13275(.A(new_n15623), .B(new_n15610), .Y(new_n15624));
  nand_5 g13276(.A(new_n15624), .B(new_n15609), .Y(new_n15625));
  xor_4  g13277(.A(new_n15605), .B(new_n9305), .Y(new_n15626));
  or_5   g13278(.A(new_n15626), .B(new_n4371), .Y(new_n15627));
  nand_5 g13279(.A(new_n15626), .B(new_n4371), .Y(new_n15628));
  nand_5 g13280(.A(new_n15628), .B(new_n15627), .Y(new_n15629));
  xor_4  g13281(.A(new_n15629), .B(new_n15625), .Y(new_n15630));
  not_8  g13282(.A(new_n15630), .Y(new_n15631));
  or_5   g13283(.A(new_n15631), .B(new_n15602_1), .Y(new_n15632));
  nand_5 g13284(.A(new_n15631), .B(new_n15602_1), .Y(new_n15633));
  nand_5 g13285(.A(new_n15587), .B(new_n15586), .Y(new_n15634));
  xor_4  g13286(.A(new_n15634), .B(new_n15596), .Y(new_n15635));
  nand_5 g13287(.A(new_n15610), .B(new_n15609), .Y(new_n15636_1));
  xor_4  g13288(.A(new_n15636_1), .B(new_n15623), .Y(new_n15637));
  nand_5 g13289(.A(new_n15637), .B(new_n15635), .Y(new_n15638));
  or_5   g13290(.A(new_n15637), .B(new_n15635), .Y(new_n15639));
  nand_5 g13291(.A(new_n15589), .B(new_n15588_1), .Y(new_n15640));
  xor_4  g13292(.A(new_n15640), .B(new_n15594), .Y(new_n15641));
  nand_5 g13293(.A(new_n15614_1), .B(new_n15613), .Y(new_n15642));
  xor_4  g13294(.A(new_n15642), .B(new_n15621), .Y(new_n15643));
  nand_5 g13295(.A(new_n15643), .B(new_n15641), .Y(new_n15644));
  or_5   g13296(.A(new_n15643), .B(new_n15641), .Y(new_n15645));
  nand_5 g13297(.A(new_n15591), .B(new_n15590_1), .Y(new_n15646));
  xor_4  g13298(.A(new_n15646), .B(new_n15592), .Y(new_n15647));
  nand_5 g13299(.A(new_n15618), .B(new_n15617), .Y(new_n15648));
  xor_4  g13300(.A(new_n15648), .B(new_n15619), .Y(new_n15649));
  nand_5 g13301(.A(new_n15649), .B(new_n15647), .Y(new_n15650));
  or_5   g13302(.A(new_n15649), .B(new_n15647), .Y(new_n15651));
  xor_4  g13303(.A(new_n2624), .B(new_n2613), .Y(new_n15652_1));
  not_8  g13304(.A(new_n15652_1), .Y(new_n15653));
  nand_5 g13305(.A(new_n5108), .B(new_n2619_1), .Y(new_n15654));
  nand_5 g13306(.A(new_n15654), .B(new_n15619), .Y(new_n15655));
  nor_5  g13307(.A(new_n15655), .B(new_n15653), .Y(new_n15656));
  nand_5 g13308(.A(new_n15656), .B(new_n15651), .Y(new_n15657));
  nand_5 g13309(.A(new_n15657), .B(new_n15650), .Y(new_n15658));
  nand_5 g13310(.A(new_n15658), .B(new_n15645), .Y(new_n15659));
  nand_5 g13311(.A(new_n15659), .B(new_n15644), .Y(new_n15660));
  nand_5 g13312(.A(new_n15660), .B(new_n15639), .Y(new_n15661));
  nand_5 g13313(.A(new_n15661), .B(new_n15638), .Y(new_n15662_1));
  nand_5 g13314(.A(new_n15662_1), .B(new_n15633), .Y(new_n15663));
  nand_5 g13315(.A(new_n15663), .B(new_n15632), .Y(new_n15664));
  nand_5 g13316(.A(new_n15628), .B(new_n15625), .Y(new_n15665));
  nand_5 g13317(.A(new_n15665), .B(new_n15627), .Y(new_n15666));
  nand_5 g13318(.A(new_n15605), .B(new_n9305), .Y(new_n15667));
  xor_4  g13319(.A(new_n15667), .B(n8324), .Y(new_n15668));
  or_5   g13320(.A(new_n15668), .B(new_n4503), .Y(new_n15669));
  nand_5 g13321(.A(new_n15668), .B(new_n4503), .Y(new_n15670));
  nand_5 g13322(.A(new_n15670), .B(new_n15669), .Y(new_n15671));
  xor_4  g13323(.A(new_n15671), .B(new_n15666), .Y(new_n15672));
  not_8  g13324(.A(new_n15672), .Y(new_n15673));
  nand_5 g13325(.A(new_n15600), .B(new_n15598_1), .Y(new_n15674));
  nand_5 g13326(.A(new_n15674), .B(new_n15599), .Y(new_n15675));
  nand_5 g13327(.A(new_n9301), .B(new_n4874), .Y(new_n15676));
  nand_5 g13328(.A(new_n9303), .B(n7678), .Y(new_n15677));
  nand_5 g13329(.A(new_n15677), .B(new_n15676), .Y(new_n15678));
  xnor_4 g13330(.A(new_n15678), .B(new_n15675), .Y(new_n15679));
  or_5   g13331(.A(new_n15679), .B(new_n15673), .Y(new_n15680));
  nand_5 g13332(.A(new_n15679), .B(new_n15673), .Y(new_n15681));
  nand_5 g13333(.A(new_n15681), .B(new_n15680), .Y(new_n15682));
  xnor_4 g13334(.A(new_n15682), .B(new_n15664), .Y(n2619));
  nand_5 g13335(.A(new_n6711), .B(new_n14514), .Y(new_n15684));
  not_8  g13336(.A(new_n15684), .Y(new_n15685));
  nand_5 g13337(.A(new_n6715), .B(new_n14517), .Y(new_n15686));
  nand_5 g13338(.A(new_n6714), .B(n12900), .Y(new_n15687));
  nand_5 g13339(.A(new_n6722), .B(new_n14520), .Y(new_n15688));
  nand_5 g13340(.A(new_n6721), .B(n20411), .Y(new_n15689));
  nand_5 g13341(.A(new_n6729_1), .B(new_n14523), .Y(new_n15690));
  nand_5 g13342(.A(new_n6728), .B(n17069), .Y(new_n15691));
  nand_5 g13343(.A(new_n6736_1), .B(new_n14526), .Y(new_n15692));
  nand_5 g13344(.A(new_n6735), .B(n15918), .Y(new_n15693));
  nand_5 g13345(.A(new_n6743), .B(new_n14529), .Y(new_n15694));
  nand_5 g13346(.A(new_n6742), .B(n17784), .Y(new_n15695));
  nand_5 g13347(.A(new_n14975), .B(new_n14972), .Y(new_n15696));
  nand_5 g13348(.A(new_n15696), .B(new_n14974), .Y(new_n15697));
  nand_5 g13349(.A(new_n15697), .B(new_n15695), .Y(new_n15698));
  nand_5 g13350(.A(new_n15698), .B(new_n15694), .Y(new_n15699));
  nand_5 g13351(.A(new_n15699), .B(new_n15693), .Y(new_n15700));
  nand_5 g13352(.A(new_n15700), .B(new_n15692), .Y(new_n15701));
  nand_5 g13353(.A(new_n15701), .B(new_n15691), .Y(new_n15702));
  nand_5 g13354(.A(new_n15702), .B(new_n15690), .Y(new_n15703));
  nand_5 g13355(.A(new_n15703), .B(new_n15689), .Y(new_n15704));
  nand_5 g13356(.A(new_n15704), .B(new_n15688), .Y(new_n15705));
  nand_5 g13357(.A(new_n15705), .B(new_n15687), .Y(new_n15706));
  nand_5 g13358(.A(new_n15706), .B(new_n15686), .Y(new_n15707));
  nor_5  g13359(.A(new_n15707), .B(new_n15685), .Y(new_n15708));
  nand_5 g13360(.A(new_n6661), .B(n10650), .Y(new_n15709));
  nand_5 g13361(.A(new_n15709), .B(new_n6660), .Y(new_n15710));
  nor_5  g13362(.A(new_n15710), .B(new_n15708), .Y(new_n15711));
  not_8  g13363(.A(new_n15711), .Y(new_n15712));
  nand_5 g13364(.A(new_n15709), .B(new_n15684), .Y(new_n15713));
  xor_4  g13365(.A(new_n15713), .B(new_n15707), .Y(new_n15714));
  not_8  g13366(.A(new_n15714), .Y(new_n15715));
  nand_5 g13367(.A(new_n15715), .B(new_n6663), .Y(new_n15716_1));
  nand_5 g13368(.A(new_n15714), .B(n6456), .Y(new_n15717));
  nand_5 g13369(.A(new_n15687), .B(new_n15686), .Y(new_n15718));
  xor_4  g13370(.A(new_n15718), .B(new_n15705), .Y(new_n15719));
  not_8  g13371(.A(new_n15719), .Y(new_n15720));
  nand_5 g13372(.A(new_n15720), .B(new_n6666), .Y(new_n15721));
  nand_5 g13373(.A(new_n15719), .B(n4085), .Y(new_n15722));
  nand_5 g13374(.A(new_n15689), .B(new_n15688), .Y(new_n15723));
  xor_4  g13375(.A(new_n15723), .B(new_n15703), .Y(new_n15724));
  not_8  g13376(.A(new_n15724), .Y(new_n15725));
  nand_5 g13377(.A(new_n15725), .B(new_n6669_1), .Y(new_n15726));
  nand_5 g13378(.A(new_n15724), .B(n26725), .Y(new_n15727));
  nand_5 g13379(.A(new_n15691), .B(new_n15690), .Y(new_n15728));
  xor_4  g13380(.A(new_n15728), .B(new_n15701), .Y(new_n15729));
  not_8  g13381(.A(new_n15729), .Y(new_n15730));
  nand_5 g13382(.A(new_n15730), .B(new_n6672), .Y(new_n15731));
  nand_5 g13383(.A(new_n15729), .B(n11980), .Y(new_n15732));
  nand_5 g13384(.A(new_n15693), .B(new_n15692), .Y(new_n15733));
  xor_4  g13385(.A(new_n15733), .B(new_n15699), .Y(new_n15734));
  not_8  g13386(.A(new_n15734), .Y(new_n15735));
  nand_5 g13387(.A(new_n15735), .B(new_n6675), .Y(new_n15736));
  nand_5 g13388(.A(new_n15734), .B(n3253), .Y(new_n15737));
  nand_5 g13389(.A(new_n15695), .B(new_n15694), .Y(new_n15738));
  xor_4  g13390(.A(new_n15738), .B(new_n15697), .Y(new_n15739));
  not_8  g13391(.A(new_n15739), .Y(new_n15740));
  nand_5 g13392(.A(new_n15740), .B(new_n6679), .Y(new_n15741));
  nand_5 g13393(.A(new_n15739), .B(n7759), .Y(new_n15742));
  nand_5 g13394(.A(new_n14980), .B(new_n14970), .Y(new_n15743_1));
  nand_5 g13395(.A(new_n15743_1), .B(new_n14978), .Y(new_n15744));
  nand_5 g13396(.A(new_n15744), .B(new_n15742), .Y(new_n15745));
  nand_5 g13397(.A(new_n15745), .B(new_n15741), .Y(new_n15746));
  nand_5 g13398(.A(new_n15746), .B(new_n15737), .Y(new_n15747));
  nand_5 g13399(.A(new_n15747), .B(new_n15736), .Y(new_n15748));
  nand_5 g13400(.A(new_n15748), .B(new_n15732), .Y(new_n15749_1));
  nand_5 g13401(.A(new_n15749_1), .B(new_n15731), .Y(new_n15750));
  nand_5 g13402(.A(new_n15750), .B(new_n15727), .Y(new_n15751));
  nand_5 g13403(.A(new_n15751), .B(new_n15726), .Y(new_n15752));
  nand_5 g13404(.A(new_n15752), .B(new_n15722), .Y(new_n15753));
  nand_5 g13405(.A(new_n15753), .B(new_n15721), .Y(new_n15754));
  nand_5 g13406(.A(new_n15754), .B(new_n15717), .Y(new_n15755));
  nand_5 g13407(.A(new_n15755), .B(new_n15716_1), .Y(new_n15756));
  nor_5  g13408(.A(new_n15756), .B(new_n15712), .Y(new_n15757));
  nor_5  g13409(.A(new_n15757), .B(new_n14512), .Y(new_n15758));
  and_5  g13410(.A(new_n15757), .B(new_n14512), .Y(new_n15759));
  xor_4  g13411(.A(new_n15756), .B(new_n15712), .Y(new_n15760));
  not_8  g13412(.A(new_n15760), .Y(new_n15761_1));
  nand_5 g13413(.A(new_n15761_1), .B(new_n14624), .Y(new_n15762_1));
  not_8  g13414(.A(new_n15762_1), .Y(new_n15763));
  nor_5  g13415(.A(new_n15761_1), .B(new_n14624), .Y(new_n15764));
  nand_5 g13416(.A(new_n15716_1), .B(new_n15717), .Y(new_n15765));
  xor_4  g13417(.A(new_n15765), .B(new_n15754), .Y(new_n15766_1));
  or_5   g13418(.A(new_n15766_1), .B(new_n14630), .Y(new_n15767));
  nand_5 g13419(.A(new_n15766_1), .B(new_n14630), .Y(new_n15768));
  not_8  g13420(.A(new_n14636_1), .Y(new_n15769));
  nand_5 g13421(.A(new_n15721), .B(new_n15722), .Y(new_n15770));
  xor_4  g13422(.A(new_n15770), .B(new_n15752), .Y(new_n15771));
  or_5   g13423(.A(new_n15771), .B(new_n15769), .Y(new_n15772));
  nand_5 g13424(.A(new_n15771), .B(new_n15769), .Y(new_n15773));
  not_8  g13425(.A(new_n14643), .Y(new_n15774));
  nand_5 g13426(.A(new_n15726), .B(new_n15727), .Y(new_n15775));
  xor_4  g13427(.A(new_n15775), .B(new_n15750), .Y(new_n15776));
  or_5   g13428(.A(new_n15776), .B(new_n15774), .Y(new_n15777));
  nand_5 g13429(.A(new_n15776), .B(new_n15774), .Y(new_n15778));
  not_8  g13430(.A(new_n14650), .Y(new_n15779));
  nand_5 g13431(.A(new_n15731), .B(new_n15732), .Y(new_n15780_1));
  xor_4  g13432(.A(new_n15780_1), .B(new_n15748), .Y(new_n15781));
  or_5   g13433(.A(new_n15781), .B(new_n15779), .Y(new_n15782));
  nand_5 g13434(.A(new_n15781), .B(new_n15779), .Y(new_n15783));
  not_8  g13435(.A(new_n14657), .Y(new_n15784));
  nand_5 g13436(.A(new_n15736), .B(new_n15737), .Y(new_n15785));
  xor_4  g13437(.A(new_n15785), .B(new_n15746), .Y(new_n15786));
  or_5   g13438(.A(new_n15786), .B(new_n15784), .Y(new_n15787));
  nand_5 g13439(.A(new_n15786), .B(new_n15784), .Y(new_n15788));
  not_8  g13440(.A(new_n14664), .Y(new_n15789));
  nand_5 g13441(.A(new_n15741), .B(new_n15742), .Y(new_n15790));
  xor_4  g13442(.A(new_n15790), .B(new_n15744), .Y(new_n15791));
  or_5   g13443(.A(new_n15791), .B(new_n15789), .Y(new_n15792));
  nand_5 g13444(.A(new_n15791), .B(new_n15789), .Y(new_n15793_1));
  nor_5  g13445(.A(new_n14986), .B(new_n14968), .Y(new_n15794));
  nor_5  g13446(.A(new_n15794), .B(new_n14985), .Y(new_n15795));
  not_8  g13447(.A(new_n15795), .Y(new_n15796));
  nand_5 g13448(.A(new_n15796), .B(new_n15793_1), .Y(new_n15797));
  nand_5 g13449(.A(new_n15797), .B(new_n15792), .Y(new_n15798));
  nand_5 g13450(.A(new_n15798), .B(new_n15788), .Y(new_n15799));
  nand_5 g13451(.A(new_n15799), .B(new_n15787), .Y(new_n15800));
  nand_5 g13452(.A(new_n15800), .B(new_n15783), .Y(new_n15801));
  nand_5 g13453(.A(new_n15801), .B(new_n15782), .Y(new_n15802));
  nand_5 g13454(.A(new_n15802), .B(new_n15778), .Y(new_n15803));
  nand_5 g13455(.A(new_n15803), .B(new_n15777), .Y(new_n15804));
  nand_5 g13456(.A(new_n15804), .B(new_n15773), .Y(new_n15805));
  nand_5 g13457(.A(new_n15805), .B(new_n15772), .Y(new_n15806));
  nand_5 g13458(.A(new_n15806), .B(new_n15768), .Y(new_n15807));
  nand_5 g13459(.A(new_n15807), .B(new_n15767), .Y(new_n15808));
  not_8  g13460(.A(new_n15808), .Y(new_n15809));
  nor_5  g13461(.A(new_n15809), .B(new_n15764), .Y(new_n15810));
  nor_5  g13462(.A(new_n15810), .B(new_n15763), .Y(new_n15811));
  nor_5  g13463(.A(new_n15811), .B(new_n15759), .Y(new_n15812_1));
  nor_5  g13464(.A(new_n15812_1), .B(new_n15758), .Y(n2661));
  nand_5 g13465(.A(new_n12863), .B(new_n12862), .Y(new_n15814));
  xor_4  g13466(.A(new_n15814), .B(new_n12873_1), .Y(n2693));
  nand_5 g13467(.A(new_n15490_1), .B(new_n8402), .Y(new_n15816_1));
  nor_5  g13468(.A(new_n15490_1), .B(new_n8402), .Y(new_n15817));
  not_8  g13469(.A(new_n15817), .Y(new_n15818));
  nand_5 g13470(.A(new_n15485), .B(new_n8407), .Y(new_n15819));
  nand_5 g13471(.A(new_n15819), .B(new_n15818), .Y(new_n15820));
  nand_5 g13472(.A(new_n15820), .B(new_n15816_1), .Y(new_n15821));
  not_8  g13473(.A(new_n15821), .Y(new_n15822));
  nand_5 g13474(.A(new_n15506_1), .B(new_n8396), .Y(new_n15823));
  nand_5 g13475(.A(new_n15507), .B(new_n8398), .Y(new_n15824));
  nand_5 g13476(.A(new_n15824), .B(new_n15823), .Y(new_n15825));
  xor_4  g13477(.A(new_n15825), .B(new_n15822), .Y(new_n15826));
  nand_5 g13478(.A(new_n11723), .B(n4326), .Y(new_n15827));
  nand_5 g13479(.A(n12593), .B(new_n3013), .Y(new_n15828));
  nand_5 g13480(.A(n13714), .B(new_n3015), .Y(new_n15829));
  nand_5 g13481(.A(new_n15829), .B(new_n15828), .Y(new_n15830));
  nand_5 g13482(.A(new_n15830), .B(new_n15827), .Y(new_n15831_1));
  nand_5 g13483(.A(new_n11720), .B(n19005), .Y(new_n15832));
  nand_5 g13484(.A(n19144), .B(new_n3010_1), .Y(new_n15833));
  nand_5 g13485(.A(new_n15833), .B(new_n15832), .Y(new_n15834));
  xor_4  g13486(.A(new_n15834), .B(new_n15831_1), .Y(new_n15835));
  or_5   g13487(.A(new_n15835), .B(new_n15826), .Y(new_n15836));
  nand_5 g13488(.A(new_n15835), .B(new_n15826), .Y(new_n15837));
  nand_5 g13489(.A(new_n15484), .B(new_n8406), .Y(new_n15838));
  nand_5 g13490(.A(new_n15838), .B(new_n15819), .Y(new_n15839));
  xor_4  g13491(.A(n13714), .B(new_n3015), .Y(new_n15840));
  nor_5  g13492(.A(new_n15840), .B(new_n15839), .Y(new_n15841));
  nand_5 g13493(.A(new_n15828), .B(new_n15827), .Y(new_n15842));
  xnor_4 g13494(.A(new_n15842), .B(new_n15829), .Y(new_n15843));
  nand_5 g13495(.A(new_n15843), .B(new_n15841), .Y(new_n15844));
  not_8  g13496(.A(new_n15844), .Y(new_n15845));
  nand_5 g13497(.A(new_n15818), .B(new_n15816_1), .Y(new_n15846_1));
  xnor_4 g13498(.A(new_n15846_1), .B(new_n15819), .Y(new_n15847));
  nor_5  g13499(.A(new_n15843), .B(new_n15841), .Y(new_n15848));
  nor_5  g13500(.A(new_n15848), .B(new_n15847), .Y(new_n15849));
  nor_5  g13501(.A(new_n15849), .B(new_n15845), .Y(new_n15850));
  not_8  g13502(.A(new_n15850), .Y(new_n15851));
  nand_5 g13503(.A(new_n15851), .B(new_n15837), .Y(new_n15852));
  nand_5 g13504(.A(new_n15852), .B(new_n15836), .Y(new_n15853));
  nand_5 g13505(.A(new_n15824), .B(new_n15821), .Y(new_n15854));
  nand_5 g13506(.A(new_n15854), .B(new_n15823), .Y(new_n15855));
  not_8  g13507(.A(new_n15855), .Y(new_n15856));
  nand_5 g13508(.A(new_n15560), .B(new_n8391), .Y(new_n15857));
  nand_5 g13509(.A(new_n15557), .B(new_n13900), .Y(new_n15858));
  nand_5 g13510(.A(new_n15858), .B(new_n15857), .Y(new_n15859_1));
  xor_4  g13511(.A(new_n15859_1), .B(new_n15856), .Y(new_n15860));
  not_8  g13512(.A(new_n15860), .Y(new_n15861));
  nand_5 g13513(.A(new_n15833), .B(new_n15831_1), .Y(new_n15862));
  nand_5 g13514(.A(new_n15862), .B(new_n15832), .Y(new_n15863));
  nand_5 g13515(.A(new_n11716), .B(n4665), .Y(new_n15864));
  nand_5 g13516(.A(n8309), .B(new_n3007), .Y(new_n15865));
  nand_5 g13517(.A(new_n15865), .B(new_n15864), .Y(new_n15866));
  xnor_4 g13518(.A(new_n15866), .B(new_n15863), .Y(new_n15867));
  nand_5 g13519(.A(new_n15867), .B(new_n15861), .Y(new_n15868));
  not_8  g13520(.A(new_n15868), .Y(new_n15869_1));
  nor_5  g13521(.A(new_n15867), .B(new_n15861), .Y(new_n15870));
  nor_5  g13522(.A(new_n15870), .B(new_n15869_1), .Y(new_n15871));
  xor_4  g13523(.A(new_n15871), .B(new_n15853), .Y(n2703));
  nand_5 g13524(.A(new_n14773), .B(new_n14772_1), .Y(new_n15873));
  xor_4  g13525(.A(new_n15873), .B(new_n14784), .Y(n2706));
  nor_5  g13526(.A(new_n7493), .B(n3541), .Y(new_n15875));
  nand_5 g13527(.A(new_n15875), .B(new_n14099), .Y(new_n15876));
  nor_5  g13528(.A(new_n15876), .B(n10018), .Y(new_n15877));
  not_8  g13529(.A(new_n15877), .Y(new_n15878));
  nand_5 g13530(.A(new_n15876), .B(n10018), .Y(new_n15879));
  and_5  g13531(.A(new_n15879), .B(new_n15878), .Y(new_n15880));
  not_8  g13532(.A(new_n15880), .Y(new_n15881));
  nand_5 g13533(.A(new_n15881), .B(new_n14201), .Y(new_n15882));
  not_8  g13534(.A(new_n15882), .Y(new_n15883));
  xor_4  g13535(.A(new_n15875), .B(n2184), .Y(new_n15884_1));
  nand_5 g13536(.A(new_n15884_1), .B(new_n14204), .Y(new_n15885_1));
  not_8  g13537(.A(new_n15884_1), .Y(new_n15886));
  nand_5 g13538(.A(new_n15886), .B(n6204), .Y(new_n15887));
  xor_4  g13539(.A(new_n7493), .B(new_n14102), .Y(new_n15888));
  nand_5 g13540(.A(new_n15888), .B(new_n14207), .Y(new_n15889_1));
  not_8  g13541(.A(new_n15888), .Y(new_n15890));
  nand_5 g13542(.A(new_n15890), .B(n3349), .Y(new_n15891));
  nand_5 g13543(.A(new_n7498), .B(new_n7489), .Y(new_n15892));
  nand_5 g13544(.A(new_n15892), .B(new_n7497), .Y(new_n15893));
  nand_5 g13545(.A(new_n15893), .B(new_n15891), .Y(new_n15894));
  nand_5 g13546(.A(new_n15894), .B(new_n15889_1), .Y(new_n15895));
  nand_5 g13547(.A(new_n15895), .B(new_n15887), .Y(new_n15896));
  nand_5 g13548(.A(new_n15896), .B(new_n15885_1), .Y(new_n15897));
  nor_5  g13549(.A(new_n15897), .B(new_n15883), .Y(new_n15898));
  nand_5 g13550(.A(new_n15880), .B(n5140), .Y(new_n15899));
  nand_5 g13551(.A(new_n15899), .B(new_n15878), .Y(new_n15900));
  nor_5  g13552(.A(new_n15900), .B(new_n15898), .Y(new_n15901));
  nand_5 g13553(.A(new_n13067), .B(new_n13051), .Y(new_n15902));
  nand_5 g13554(.A(new_n15902), .B(new_n13053), .Y(new_n15903));
  not_8  g13555(.A(new_n15903), .Y(new_n15904));
  nand_5 g13556(.A(new_n15904), .B(new_n15901), .Y(new_n15905));
  nand_5 g13557(.A(new_n15899), .B(new_n15882), .Y(new_n15906));
  xor_4  g13558(.A(new_n15906), .B(new_n15897), .Y(new_n15907));
  nand_5 g13559(.A(new_n15907), .B(new_n13069), .Y(new_n15908));
  or_5   g13560(.A(new_n15907), .B(new_n13069), .Y(new_n15909));
  nand_5 g13561(.A(new_n15887), .B(new_n15885_1), .Y(new_n15910));
  xor_4  g13562(.A(new_n15910), .B(new_n15895), .Y(new_n15911));
  nand_5 g13563(.A(new_n15911), .B(new_n13075), .Y(new_n15912));
  or_5   g13564(.A(new_n15911), .B(new_n13075), .Y(new_n15913));
  nand_5 g13565(.A(new_n15891), .B(new_n15889_1), .Y(new_n15914));
  xor_4  g13566(.A(new_n15914), .B(new_n15893), .Y(new_n15915));
  nand_5 g13567(.A(new_n15915), .B(new_n13083), .Y(new_n15916));
  nor_5  g13568(.A(new_n15915), .B(new_n13083), .Y(new_n15917_1));
  not_8  g13569(.A(new_n15917_1), .Y(new_n15918_1));
  nand_5 g13570(.A(new_n7502), .B(new_n7476), .Y(new_n15919));
  nand_5 g13571(.A(new_n15919), .B(new_n7501), .Y(new_n15920));
  nand_5 g13572(.A(new_n15920), .B(new_n15918_1), .Y(new_n15921));
  nand_5 g13573(.A(new_n15921), .B(new_n15916), .Y(new_n15922_1));
  nand_5 g13574(.A(new_n15922_1), .B(new_n15913), .Y(new_n15923));
  nand_5 g13575(.A(new_n15923), .B(new_n15912), .Y(new_n15924));
  nand_5 g13576(.A(new_n15924), .B(new_n15909), .Y(new_n15925));
  nand_5 g13577(.A(new_n15925), .B(new_n15908), .Y(new_n15926));
  or_5   g13578(.A(new_n15904), .B(new_n15901), .Y(new_n15927));
  nand_5 g13579(.A(new_n15927), .B(new_n15926), .Y(new_n15928));
  nand_5 g13580(.A(new_n15928), .B(new_n15905), .Y(new_n15929));
  xor_4  g13581(.A(new_n15929), .B(new_n15901), .Y(new_n15930));
  not_8  g13582(.A(n1831), .Y(new_n15931));
  or_5   g13583(.A(n3320), .B(new_n15931), .Y(new_n15932));
  nand_5 g13584(.A(n3320), .B(new_n15931), .Y(new_n15933));
  nand_5 g13585(.A(n13137), .B(new_n7045), .Y(new_n15934));
  nand_5 g13586(.A(new_n6992), .B(n1288), .Y(new_n15935));
  nand_5 g13587(.A(n18452), .B(new_n7061), .Y(new_n15936_1));
  nand_5 g13588(.A(new_n6998_1), .B(n1752), .Y(new_n15937));
  nand_5 g13589(.A(n21317), .B(new_n7046), .Y(new_n15938));
  nand_5 g13590(.A(new_n7004), .B(n13110), .Y(new_n15939));
  or_5   g13591(.A(n25694), .B(new_n4522), .Y(new_n15940));
  nand_5 g13592(.A(n25694), .B(new_n4522), .Y(new_n15941));
  nand_5 g13593(.A(n19789), .B(new_n4439), .Y(new_n15942));
  nand_5 g13594(.A(new_n4523), .B(n15424), .Y(new_n15943));
  nand_5 g13595(.A(new_n14021), .B(new_n14019), .Y(new_n15944));
  nand_5 g13596(.A(new_n15944), .B(new_n14020), .Y(new_n15945));
  nand_5 g13597(.A(new_n15945), .B(new_n15943), .Y(new_n15946));
  nand_5 g13598(.A(new_n15946), .B(new_n15942), .Y(new_n15947_1));
  nand_5 g13599(.A(new_n15947_1), .B(new_n15941), .Y(new_n15948));
  nand_5 g13600(.A(new_n15948), .B(new_n15940), .Y(new_n15949));
  nand_5 g13601(.A(new_n15949), .B(new_n15939), .Y(new_n15950));
  nand_5 g13602(.A(new_n15950), .B(new_n15938), .Y(new_n15951));
  nand_5 g13603(.A(new_n15951), .B(new_n15937), .Y(new_n15952));
  nand_5 g13604(.A(new_n15952), .B(new_n15936_1), .Y(new_n15953));
  nand_5 g13605(.A(new_n15953), .B(new_n15935), .Y(new_n15954));
  nand_5 g13606(.A(new_n15954), .B(new_n15934), .Y(new_n15955));
  nand_5 g13607(.A(new_n15955), .B(new_n15933), .Y(new_n15956_1));
  nand_5 g13608(.A(new_n15956_1), .B(new_n15932), .Y(new_n15957));
  nor_5  g13609(.A(new_n15957), .B(new_n15930), .Y(new_n15958_1));
  and_5  g13610(.A(new_n15957), .B(new_n15930), .Y(new_n15959));
  nor_5  g13611(.A(new_n15959), .B(new_n15958_1), .Y(new_n15960));
  xor_4  g13612(.A(new_n15926), .B(new_n15901), .Y(new_n15961));
  xor_4  g13613(.A(new_n15961), .B(new_n15904), .Y(new_n15962));
  not_8  g13614(.A(new_n15962), .Y(new_n15963));
  nand_5 g13615(.A(new_n15963), .B(new_n15957), .Y(new_n15964));
  or_5   g13616(.A(new_n15963), .B(new_n15957), .Y(new_n15965));
  nand_5 g13617(.A(new_n15933), .B(new_n15932), .Y(new_n15966));
  xor_4  g13618(.A(new_n15966), .B(new_n15955), .Y(new_n15967_1));
  nand_5 g13619(.A(new_n15909), .B(new_n15908), .Y(new_n15968));
  xor_4  g13620(.A(new_n15968), .B(new_n15924), .Y(new_n15969));
  nand_5 g13621(.A(new_n15969), .B(new_n15967_1), .Y(new_n15970));
  not_8  g13622(.A(new_n15970), .Y(new_n15971));
  nor_5  g13623(.A(new_n15969), .B(new_n15967_1), .Y(new_n15972));
  nand_5 g13624(.A(new_n15935), .B(new_n15934), .Y(new_n15973));
  xor_4  g13625(.A(new_n15973), .B(new_n15953), .Y(new_n15974));
  nand_5 g13626(.A(new_n15913), .B(new_n15912), .Y(new_n15975));
  xor_4  g13627(.A(new_n15975), .B(new_n15922_1), .Y(new_n15976));
  nand_5 g13628(.A(new_n15976), .B(new_n15974), .Y(new_n15977));
  not_8  g13629(.A(new_n15977), .Y(new_n15978));
  nor_5  g13630(.A(new_n15976), .B(new_n15974), .Y(new_n15979_1));
  nand_5 g13631(.A(new_n15918_1), .B(new_n15916), .Y(new_n15980));
  xor_4  g13632(.A(new_n15980), .B(new_n15920), .Y(new_n15981));
  nand_5 g13633(.A(new_n15937), .B(new_n15936_1), .Y(new_n15982));
  xor_4  g13634(.A(new_n15982), .B(new_n15951), .Y(new_n15983));
  or_5   g13635(.A(new_n15983), .B(new_n15981), .Y(new_n15984));
  nand_5 g13636(.A(new_n15983), .B(new_n15981), .Y(new_n15985));
  nand_5 g13637(.A(new_n15939), .B(new_n15938), .Y(new_n15986_1));
  xor_4  g13638(.A(new_n15986_1), .B(new_n15949), .Y(new_n15987));
  or_5   g13639(.A(new_n15987), .B(new_n7505), .Y(new_n15988));
  nand_5 g13640(.A(new_n15987), .B(new_n7505), .Y(new_n15989));
  nand_5 g13641(.A(new_n15941), .B(new_n15940), .Y(new_n15990));
  xor_4  g13642(.A(new_n15990), .B(new_n15947_1), .Y(new_n15991));
  or_5   g13643(.A(new_n15991), .B(new_n7430), .Y(new_n15992));
  nand_5 g13644(.A(new_n15991), .B(new_n7430), .Y(new_n15993));
  nand_5 g13645(.A(new_n15943), .B(new_n15942), .Y(new_n15994));
  xor_4  g13646(.A(new_n15994), .B(new_n15945), .Y(new_n15995));
  or_5   g13647(.A(new_n15995), .B(new_n7435), .Y(new_n15996));
  nand_5 g13648(.A(new_n15995), .B(new_n7435), .Y(new_n15997));
  not_8  g13649(.A(new_n14017), .Y(new_n15998));
  nor_5  g13650(.A(new_n14026), .B(new_n15998), .Y(new_n15999));
  nor_5  g13651(.A(new_n15999), .B(new_n14025), .Y(new_n16000));
  not_8  g13652(.A(new_n16000), .Y(new_n16001));
  nand_5 g13653(.A(new_n16001), .B(new_n15997), .Y(new_n16002));
  nand_5 g13654(.A(new_n16002), .B(new_n15996), .Y(new_n16003));
  nand_5 g13655(.A(new_n16003), .B(new_n15993), .Y(new_n16004));
  nand_5 g13656(.A(new_n16004), .B(new_n15992), .Y(new_n16005));
  nand_5 g13657(.A(new_n16005), .B(new_n15989), .Y(new_n16006));
  nand_5 g13658(.A(new_n16006), .B(new_n15988), .Y(new_n16007));
  nand_5 g13659(.A(new_n16007), .B(new_n15985), .Y(new_n16008));
  nand_5 g13660(.A(new_n16008), .B(new_n15984), .Y(new_n16009));
  nor_5  g13661(.A(new_n16009), .B(new_n15979_1), .Y(new_n16010));
  nor_5  g13662(.A(new_n16010), .B(new_n15978), .Y(new_n16011));
  nor_5  g13663(.A(new_n16011), .B(new_n15972), .Y(new_n16012));
  nor_5  g13664(.A(new_n16012), .B(new_n15971), .Y(new_n16013_1));
  not_8  g13665(.A(new_n16013_1), .Y(new_n16014));
  nand_5 g13666(.A(new_n16014), .B(new_n15965), .Y(new_n16015));
  nand_5 g13667(.A(new_n16015), .B(new_n15964), .Y(new_n16016));
  xor_4  g13668(.A(new_n16016), .B(new_n15960), .Y(n2711));
  nand_5 g13669(.A(n15490), .B(new_n10457), .Y(new_n16018));
  nand_5 g13670(.A(new_n7550), .B(n7339), .Y(new_n16019));
  nand_5 g13671(.A(n26808), .B(new_n7558_1), .Y(new_n16020));
  nand_5 g13672(.A(new_n16020), .B(new_n16019), .Y(new_n16021));
  nand_5 g13673(.A(new_n16021), .B(new_n16018), .Y(new_n16022));
  nand_5 g13674(.A(n2783), .B(new_n12343), .Y(new_n16023));
  nand_5 g13675(.A(new_n7569_1), .B(n1667), .Y(new_n16024));
  nand_5 g13676(.A(new_n16024), .B(new_n16023), .Y(new_n16025));
  xor_4  g13677(.A(new_n16025), .B(new_n16022), .Y(new_n16026));
  nand_5 g13678(.A(new_n16026), .B(new_n10415), .Y(new_n16027));
  or_5   g13679(.A(new_n16026), .B(new_n10415), .Y(new_n16028));
  xor_4  g13680(.A(n26808), .B(new_n7558_1), .Y(new_n16029_1));
  nor_5  g13681(.A(new_n16029_1), .B(new_n10423), .Y(new_n16030));
  nand_5 g13682(.A(new_n16019), .B(new_n16018), .Y(new_n16031));
  xnor_4 g13683(.A(new_n16031), .B(new_n16020), .Y(new_n16032));
  and_5  g13684(.A(new_n16032), .B(new_n16030), .Y(new_n16033));
  nor_5  g13685(.A(new_n16032), .B(new_n16030), .Y(new_n16034));
  nor_5  g13686(.A(new_n16034), .B(new_n10432_1), .Y(new_n16035));
  nor_5  g13687(.A(new_n16035), .B(new_n16033), .Y(new_n16036));
  nand_5 g13688(.A(new_n16036), .B(new_n16028), .Y(new_n16037));
  nand_5 g13689(.A(new_n16037), .B(new_n16027), .Y(new_n16038));
  nand_5 g13690(.A(new_n16024), .B(new_n16022), .Y(new_n16039));
  nand_5 g13691(.A(new_n16039), .B(new_n16023), .Y(new_n16040));
  nand_5 g13692(.A(n10611), .B(new_n12354), .Y(new_n16041));
  nand_5 g13693(.A(new_n7620), .B(n2680), .Y(new_n16042));
  nand_5 g13694(.A(new_n16042), .B(new_n16041), .Y(new_n16043));
  xnor_4 g13695(.A(new_n16043), .B(new_n16040), .Y(new_n16044));
  nand_5 g13696(.A(new_n16044), .B(new_n10407), .Y(new_n16045));
  or_5   g13697(.A(new_n16044), .B(new_n10407), .Y(new_n16046));
  nand_5 g13698(.A(new_n16046), .B(new_n16045), .Y(new_n16047));
  xor_4  g13699(.A(new_n16047), .B(new_n16038), .Y(n2761));
  nand_5 g13700(.A(new_n8798), .B(new_n6846), .Y(new_n16049));
  nand_5 g13701(.A(new_n8801), .B(new_n6849), .Y(new_n16050));
  nand_5 g13702(.A(new_n6855), .B(new_n8804), .Y(new_n16051));
  nand_5 g13703(.A(new_n10838), .B(new_n10835), .Y(new_n16052));
  nand_5 g13704(.A(new_n16052), .B(new_n10837), .Y(new_n16053));
  nand_5 g13705(.A(n20359), .B(n14680), .Y(new_n16054));
  nand_5 g13706(.A(new_n16054), .B(new_n16053), .Y(new_n16055));
  nand_5 g13707(.A(new_n16055), .B(new_n16051), .Y(new_n16056));
  nand_5 g13708(.A(n8363), .B(n2816), .Y(new_n16057));
  nand_5 g13709(.A(new_n16057), .B(new_n16056), .Y(new_n16058));
  nand_5 g13710(.A(new_n16058), .B(new_n16050), .Y(new_n16059));
  nand_5 g13711(.A(n25120), .B(n8526), .Y(new_n16060_1));
  nand_5 g13712(.A(new_n16060_1), .B(new_n16059), .Y(new_n16061));
  nand_5 g13713(.A(new_n16061), .B(new_n16049), .Y(new_n16062_1));
  nand_5 g13714(.A(new_n16060_1), .B(new_n16049), .Y(new_n16063));
  xor_4  g13715(.A(new_n16063), .B(new_n16059), .Y(new_n16064));
  not_8  g13716(.A(new_n16064), .Y(new_n16065));
  nand_5 g13717(.A(new_n16065), .B(new_n8291), .Y(new_n16066));
  nand_5 g13718(.A(new_n16064), .B(n17458), .Y(new_n16067));
  nand_5 g13719(.A(new_n16057), .B(new_n16050), .Y(new_n16068_1));
  xor_4  g13720(.A(new_n16068_1), .B(new_n16056), .Y(new_n16069));
  not_8  g13721(.A(new_n16069), .Y(new_n16070));
  nand_5 g13722(.A(new_n16070), .B(new_n8294), .Y(new_n16071));
  nand_5 g13723(.A(new_n16069), .B(n1222), .Y(new_n16072));
  nand_5 g13724(.A(new_n16054), .B(new_n16051), .Y(new_n16073));
  xor_4  g13725(.A(new_n16073), .B(new_n16053), .Y(new_n16074));
  not_8  g13726(.A(new_n16074), .Y(new_n16075));
  nand_5 g13727(.A(new_n16075), .B(new_n8297), .Y(new_n16076));
  nand_5 g13728(.A(new_n16074), .B(n25240), .Y(new_n16077));
  nand_5 g13729(.A(new_n10840), .B(new_n8300), .Y(new_n16078));
  nand_5 g13730(.A(new_n10842), .B(n10125), .Y(new_n16079));
  nand_5 g13731(.A(new_n10770), .B(new_n8303), .Y(new_n16080_1));
  nand_5 g13732(.A(new_n10772), .B(n8067), .Y(new_n16081));
  nand_5 g13733(.A(new_n10732), .B(new_n8306_1), .Y(new_n16082));
  nand_5 g13734(.A(new_n10734), .B(n20923), .Y(new_n16083));
  nand_5 g13735(.A(new_n10738), .B(new_n7606), .Y(new_n16084));
  nand_5 g13736(.A(new_n10737), .B(n18157), .Y(new_n16085));
  nand_5 g13737(.A(new_n10743), .B(new_n7538), .Y(new_n16086));
  nand_5 g13738(.A(new_n10742), .B(n12161), .Y(new_n16087));
  nand_5 g13739(.A(new_n10748), .B(new_n7519), .Y(new_n16088));
  nand_5 g13740(.A(new_n10750), .B(n5026), .Y(new_n16089));
  nand_5 g13741(.A(new_n10754), .B(n8581), .Y(new_n16090));
  nand_5 g13742(.A(new_n16090), .B(new_n16089), .Y(new_n16091));
  nand_5 g13743(.A(new_n16091), .B(new_n16088), .Y(new_n16092));
  nand_5 g13744(.A(new_n16092), .B(new_n16087), .Y(new_n16093));
  nand_5 g13745(.A(new_n16093), .B(new_n16086), .Y(new_n16094));
  nand_5 g13746(.A(new_n16094), .B(new_n16085), .Y(new_n16095));
  nand_5 g13747(.A(new_n16095), .B(new_n16084), .Y(new_n16096));
  nand_5 g13748(.A(new_n16096), .B(new_n16083), .Y(new_n16097));
  nand_5 g13749(.A(new_n16097), .B(new_n16082), .Y(new_n16098_1));
  nand_5 g13750(.A(new_n16098_1), .B(new_n16081), .Y(new_n16099));
  nand_5 g13751(.A(new_n16099), .B(new_n16080_1), .Y(new_n16100));
  nand_5 g13752(.A(new_n16100), .B(new_n16079), .Y(new_n16101));
  nand_5 g13753(.A(new_n16101), .B(new_n16078), .Y(new_n16102));
  nand_5 g13754(.A(new_n16102), .B(new_n16077), .Y(new_n16103));
  nand_5 g13755(.A(new_n16103), .B(new_n16076), .Y(new_n16104));
  nand_5 g13756(.A(new_n16104), .B(new_n16072), .Y(new_n16105));
  nand_5 g13757(.A(new_n16105), .B(new_n16071), .Y(new_n16106));
  nand_5 g13758(.A(new_n16106), .B(new_n16067), .Y(new_n16107));
  nand_5 g13759(.A(new_n16107), .B(new_n16066), .Y(new_n16108));
  nor_5  g13760(.A(new_n16108), .B(new_n16062_1), .Y(new_n16109));
  nor_5  g13761(.A(new_n4299), .B(n1099), .Y(new_n16110_1));
  nand_5 g13762(.A(new_n16110_1), .B(new_n8434), .Y(new_n16111));
  nor_5  g13763(.A(new_n16111), .B(n11898), .Y(new_n16112));
  nand_5 g13764(.A(new_n16112), .B(new_n5493), .Y(new_n16113));
  not_8  g13765(.A(new_n16112), .Y(new_n16114));
  nand_5 g13766(.A(new_n16111), .B(n11898), .Y(new_n16115));
  and_5  g13767(.A(new_n16115), .B(new_n16114), .Y(new_n16116));
  not_8  g13768(.A(new_n16116), .Y(new_n16117));
  nand_5 g13769(.A(new_n16117), .B(new_n5424), .Y(new_n16118));
  nand_5 g13770(.A(new_n16116), .B(new_n5422), .Y(new_n16119));
  xor_4  g13771(.A(new_n16110_1), .B(new_n8434), .Y(new_n16120));
  not_8  g13772(.A(new_n16120), .Y(new_n16121));
  nand_5 g13773(.A(new_n16121), .B(new_n5427), .Y(new_n16122));
  nand_5 g13774(.A(new_n16120), .B(new_n5428), .Y(new_n16123));
  xor_4  g13775(.A(new_n4299), .B(n1099), .Y(new_n16124));
  not_8  g13776(.A(new_n16124), .Y(new_n16125));
  nand_5 g13777(.A(new_n16125), .B(new_n5432), .Y(new_n16126));
  nand_5 g13778(.A(new_n16124), .B(new_n5433), .Y(new_n16127));
  nand_5 g13779(.A(new_n5437), .B(new_n4302), .Y(new_n16128));
  nand_5 g13780(.A(new_n5438_1), .B(new_n4301), .Y(new_n16129));
  nand_5 g13781(.A(new_n5442), .B(new_n4227), .Y(new_n16130));
  nand_5 g13782(.A(new_n5443_1), .B(new_n4226), .Y(new_n16131));
  nand_5 g13783(.A(new_n5447), .B(new_n4182), .Y(new_n16132));
  nand_5 g13784(.A(new_n5448), .B(new_n4181), .Y(new_n16133));
  nand_5 g13785(.A(new_n5453), .B(new_n4157), .Y(new_n16134));
  not_8  g13786(.A(new_n16134), .Y(new_n16135));
  nand_5 g13787(.A(new_n5454), .B(new_n4156), .Y(new_n16136));
  not_8  g13788(.A(new_n16136), .Y(new_n16137));
  nand_5 g13789(.A(new_n5459), .B(new_n4163), .Y(new_n16138));
  not_8  g13790(.A(new_n16138), .Y(new_n16139));
  nand_5 g13791(.A(new_n5460), .B(new_n4162), .Y(new_n16140));
  not_8  g13792(.A(new_n16140), .Y(new_n16141));
  nand_5 g13793(.A(new_n5471), .B(new_n4149), .Y(new_n16142_1));
  nand_5 g13794(.A(new_n16142_1), .B(new_n4167), .Y(new_n16143));
  nand_5 g13795(.A(new_n5471), .B(new_n4151_1), .Y(new_n16144));
  nand_5 g13796(.A(new_n16144), .B(new_n5465), .Y(new_n16145));
  nand_5 g13797(.A(new_n16145), .B(new_n16143), .Y(new_n16146));
  nor_5  g13798(.A(new_n16146), .B(new_n16141), .Y(new_n16147));
  nor_5  g13799(.A(new_n16147), .B(new_n16139), .Y(new_n16148));
  nor_5  g13800(.A(new_n16148), .B(new_n16137), .Y(new_n16149));
  nor_5  g13801(.A(new_n16149), .B(new_n16135), .Y(new_n16150));
  not_8  g13802(.A(new_n16150), .Y(new_n16151));
  nand_5 g13803(.A(new_n16151), .B(new_n16133), .Y(new_n16152));
  nand_5 g13804(.A(new_n16152), .B(new_n16132), .Y(new_n16153));
  nand_5 g13805(.A(new_n16153), .B(new_n16131), .Y(new_n16154));
  nand_5 g13806(.A(new_n16154), .B(new_n16130), .Y(new_n16155));
  nand_5 g13807(.A(new_n16155), .B(new_n16129), .Y(new_n16156));
  nand_5 g13808(.A(new_n16156), .B(new_n16128), .Y(new_n16157));
  nand_5 g13809(.A(new_n16157), .B(new_n16127), .Y(new_n16158_1));
  nand_5 g13810(.A(new_n16158_1), .B(new_n16126), .Y(new_n16159));
  nand_5 g13811(.A(new_n16159), .B(new_n16123), .Y(new_n16160));
  nand_5 g13812(.A(new_n16160), .B(new_n16122), .Y(new_n16161));
  nand_5 g13813(.A(new_n16161), .B(new_n16119), .Y(new_n16162));
  nand_5 g13814(.A(new_n16162), .B(new_n16118), .Y(new_n16163));
  nor_5  g13815(.A(new_n16163), .B(new_n16113), .Y(new_n16164));
  nand_5 g13816(.A(new_n16163), .B(new_n5418), .Y(new_n16165));
  nor_5  g13817(.A(new_n16165), .B(new_n16112), .Y(new_n16166));
  nor_5  g13818(.A(new_n16166), .B(new_n16164), .Y(new_n16167_1));
  nor_5  g13819(.A(new_n16167_1), .B(new_n16109), .Y(new_n16168));
  not_8  g13820(.A(new_n16109), .Y(new_n16169));
  nand_5 g13821(.A(new_n16108), .B(new_n16062_1), .Y(new_n16170));
  and_5  g13822(.A(new_n16170), .B(new_n16169), .Y(new_n16171));
  not_8  g13823(.A(new_n16171), .Y(new_n16172));
  nand_5 g13824(.A(new_n16114), .B(new_n5418), .Y(new_n16173));
  nand_5 g13825(.A(new_n16173), .B(new_n16113), .Y(new_n16174));
  xor_4  g13826(.A(new_n16174), .B(new_n16163), .Y(new_n16175));
  nand_5 g13827(.A(new_n16175), .B(new_n16172), .Y(new_n16176));
  or_5   g13828(.A(new_n16175), .B(new_n16172), .Y(new_n16177));
  nand_5 g13829(.A(new_n16066), .B(new_n16067), .Y(new_n16178));
  xor_4  g13830(.A(new_n16178), .B(new_n16106), .Y(new_n16179));
  nand_5 g13831(.A(new_n16119), .B(new_n16118), .Y(new_n16180));
  xor_4  g13832(.A(new_n16180), .B(new_n16161), .Y(new_n16181));
  or_5   g13833(.A(new_n16181), .B(new_n16179), .Y(new_n16182));
  nand_5 g13834(.A(new_n16181), .B(new_n16179), .Y(new_n16183));
  nand_5 g13835(.A(new_n16071), .B(new_n16072), .Y(new_n16184));
  xor_4  g13836(.A(new_n16184), .B(new_n16104), .Y(new_n16185_1));
  nand_5 g13837(.A(new_n16123), .B(new_n16122), .Y(new_n16186));
  xor_4  g13838(.A(new_n16186), .B(new_n16159), .Y(new_n16187));
  or_5   g13839(.A(new_n16187), .B(new_n16185_1), .Y(new_n16188));
  nand_5 g13840(.A(new_n16187), .B(new_n16185_1), .Y(new_n16189));
  nand_5 g13841(.A(new_n16076), .B(new_n16077), .Y(new_n16190));
  xor_4  g13842(.A(new_n16190), .B(new_n16102), .Y(new_n16191));
  nand_5 g13843(.A(new_n16127), .B(new_n16126), .Y(new_n16192));
  xor_4  g13844(.A(new_n16192), .B(new_n16157), .Y(new_n16193));
  or_5   g13845(.A(new_n16193), .B(new_n16191), .Y(new_n16194));
  nand_5 g13846(.A(new_n16193), .B(new_n16191), .Y(new_n16195));
  nand_5 g13847(.A(new_n16078), .B(new_n16079), .Y(new_n16196_1));
  xor_4  g13848(.A(new_n16196_1), .B(new_n16100), .Y(new_n16197));
  nand_5 g13849(.A(new_n16129), .B(new_n16128), .Y(new_n16198));
  xor_4  g13850(.A(new_n16198), .B(new_n16155), .Y(new_n16199));
  or_5   g13851(.A(new_n16199), .B(new_n16197), .Y(new_n16200));
  nand_5 g13852(.A(new_n16199), .B(new_n16197), .Y(new_n16201));
  nand_5 g13853(.A(new_n16080_1), .B(new_n16081), .Y(new_n16202));
  xor_4  g13854(.A(new_n16202), .B(new_n16098_1), .Y(new_n16203));
  nand_5 g13855(.A(new_n16131), .B(new_n16130), .Y(new_n16204));
  xor_4  g13856(.A(new_n16204), .B(new_n16153), .Y(new_n16205));
  or_5   g13857(.A(new_n16205), .B(new_n16203), .Y(new_n16206_1));
  nand_5 g13858(.A(new_n16205), .B(new_n16203), .Y(new_n16207));
  nand_5 g13859(.A(new_n16082), .B(new_n16083), .Y(new_n16208));
  xor_4  g13860(.A(new_n16208), .B(new_n16096), .Y(new_n16209));
  nand_5 g13861(.A(new_n16133), .B(new_n16132), .Y(new_n16210));
  xor_4  g13862(.A(new_n16210), .B(new_n16151), .Y(new_n16211));
  or_5   g13863(.A(new_n16211), .B(new_n16209), .Y(new_n16212));
  nand_5 g13864(.A(new_n16211), .B(new_n16209), .Y(new_n16213));
  nand_5 g13865(.A(new_n16084), .B(new_n16085), .Y(new_n16214));
  xor_4  g13866(.A(new_n16214), .B(new_n16094), .Y(new_n16215_1));
  not_8  g13867(.A(new_n16215_1), .Y(new_n16216));
  nand_5 g13868(.A(new_n16136), .B(new_n16134), .Y(new_n16217_1));
  xor_4  g13869(.A(new_n16217_1), .B(new_n16148), .Y(new_n16218_1));
  nand_5 g13870(.A(new_n16218_1), .B(new_n16216), .Y(new_n16219_1));
  or_5   g13871(.A(new_n16218_1), .B(new_n16216), .Y(new_n16220));
  nand_5 g13872(.A(new_n16086), .B(new_n16087), .Y(new_n16221));
  xor_4  g13873(.A(new_n16221), .B(new_n16092), .Y(new_n16222));
  not_8  g13874(.A(new_n16222), .Y(new_n16223_1));
  nand_5 g13875(.A(new_n16140), .B(new_n16138), .Y(new_n16224));
  xor_4  g13876(.A(new_n16224), .B(new_n16146), .Y(new_n16225));
  nand_5 g13877(.A(new_n16225), .B(new_n16223_1), .Y(new_n16226));
  or_5   g13878(.A(new_n16225), .B(new_n16223_1), .Y(new_n16227));
  nand_5 g13879(.A(new_n16088), .B(new_n16089), .Y(new_n16228));
  xor_4  g13880(.A(new_n16228), .B(new_n16090), .Y(new_n16229));
  not_8  g13881(.A(new_n16229), .Y(new_n16230_1));
  nand_5 g13882(.A(new_n16144), .B(new_n16143), .Y(new_n16231));
  xor_4  g13883(.A(new_n16231), .B(new_n5465), .Y(new_n16232));
  nand_5 g13884(.A(new_n16232), .B(new_n16230_1), .Y(new_n16233));
  or_5   g13885(.A(new_n16232), .B(new_n16230_1), .Y(new_n16234));
  nand_5 g13886(.A(new_n10753), .B(new_n7526), .Y(new_n16235));
  and_5  g13887(.A(new_n16235), .B(new_n16090), .Y(new_n16236));
  not_8  g13888(.A(new_n16236), .Y(new_n16237));
  xor_4  g13889(.A(new_n5471), .B(new_n4149), .Y(new_n16238));
  or_5   g13890(.A(new_n16238), .B(new_n16237), .Y(new_n16239));
  nand_5 g13891(.A(new_n16239), .B(new_n16234), .Y(new_n16240));
  nand_5 g13892(.A(new_n16240), .B(new_n16233), .Y(new_n16241));
  nand_5 g13893(.A(new_n16241), .B(new_n16227), .Y(new_n16242));
  nand_5 g13894(.A(new_n16242), .B(new_n16226), .Y(new_n16243_1));
  nand_5 g13895(.A(new_n16243_1), .B(new_n16220), .Y(new_n16244));
  nand_5 g13896(.A(new_n16244), .B(new_n16219_1), .Y(new_n16245));
  nand_5 g13897(.A(new_n16245), .B(new_n16213), .Y(new_n16246));
  nand_5 g13898(.A(new_n16246), .B(new_n16212), .Y(new_n16247_1));
  nand_5 g13899(.A(new_n16247_1), .B(new_n16207), .Y(new_n16248));
  nand_5 g13900(.A(new_n16248), .B(new_n16206_1), .Y(new_n16249));
  nand_5 g13901(.A(new_n16249), .B(new_n16201), .Y(new_n16250));
  nand_5 g13902(.A(new_n16250), .B(new_n16200), .Y(new_n16251));
  nand_5 g13903(.A(new_n16251), .B(new_n16195), .Y(new_n16252));
  nand_5 g13904(.A(new_n16252), .B(new_n16194), .Y(new_n16253));
  nand_5 g13905(.A(new_n16253), .B(new_n16189), .Y(new_n16254));
  nand_5 g13906(.A(new_n16254), .B(new_n16188), .Y(new_n16255));
  nand_5 g13907(.A(new_n16255), .B(new_n16183), .Y(new_n16256));
  nand_5 g13908(.A(new_n16256), .B(new_n16182), .Y(new_n16257));
  nand_5 g13909(.A(new_n16257), .B(new_n16177), .Y(new_n16258));
  nand_5 g13910(.A(new_n16258), .B(new_n16176), .Y(new_n16259));
  nor_5  g13911(.A(new_n16259), .B(new_n16168), .Y(new_n16260));
  not_8  g13912(.A(new_n16164), .Y(new_n16261));
  nand_5 g13913(.A(new_n16167_1), .B(new_n16109), .Y(new_n16262));
  nand_5 g13914(.A(new_n16262), .B(new_n16261), .Y(new_n16263));
  nor_5  g13915(.A(new_n16263), .B(new_n16260), .Y(n2774));
  nand_5 g13916(.A(new_n3786), .B(new_n3726), .Y(new_n16265));
  nand_5 g13917(.A(new_n3790), .B(n442), .Y(new_n16266));
  nand_5 g13918(.A(new_n3794_1), .B(new_n3730), .Y(new_n16267));
  or_5   g13919(.A(new_n3794_1), .B(new_n3730), .Y(new_n16268));
  nand_5 g13920(.A(new_n3800), .B(new_n3734), .Y(new_n16269));
  nand_5 g13921(.A(new_n3799), .B(n4913), .Y(new_n16270));
  nand_5 g13922(.A(new_n3806), .B(new_n3738), .Y(new_n16271));
  nand_5 g13923(.A(new_n3805), .B(n604), .Y(new_n16272));
  nand_5 g13924(.A(new_n3813), .B(new_n3742), .Y(new_n16273));
  nand_5 g13925(.A(new_n3812), .B(n16824), .Y(new_n16274));
  nand_5 g13926(.A(new_n3821), .B(new_n3746), .Y(new_n16275_1));
  nand_5 g13927(.A(new_n3820), .B(n16521), .Y(new_n16276));
  nand_5 g13928(.A(n21993), .B(n7139), .Y(new_n16277));
  nand_5 g13929(.A(new_n16277), .B(new_n16276), .Y(new_n16278));
  nand_5 g13930(.A(new_n16278), .B(new_n16275_1), .Y(new_n16279_1));
  nand_5 g13931(.A(new_n16279_1), .B(new_n16274), .Y(new_n16280));
  nand_5 g13932(.A(new_n16280), .B(new_n16273), .Y(new_n16281));
  nand_5 g13933(.A(new_n16281), .B(new_n16272), .Y(new_n16282));
  nand_5 g13934(.A(new_n16282), .B(new_n16271), .Y(new_n16283));
  nand_5 g13935(.A(new_n16283), .B(new_n16270), .Y(new_n16284));
  nand_5 g13936(.A(new_n16284), .B(new_n16269), .Y(new_n16285));
  nand_5 g13937(.A(new_n16285), .B(new_n16268), .Y(new_n16286));
  nand_5 g13938(.A(new_n16286), .B(new_n16267), .Y(new_n16287));
  nand_5 g13939(.A(new_n16287), .B(new_n16266), .Y(new_n16288));
  nand_5 g13940(.A(new_n16288), .B(new_n16265), .Y(new_n16289));
  nand_5 g13941(.A(new_n3779), .B(new_n3722), .Y(new_n16290));
  nand_5 g13942(.A(new_n3783), .B(n13719), .Y(new_n16291));
  nand_5 g13943(.A(new_n16291), .B(new_n16290), .Y(new_n16292));
  xor_4  g13944(.A(new_n16292), .B(new_n16289), .Y(new_n16293));
  or_5   g13945(.A(new_n10932), .B(n987), .Y(new_n16294));
  nor_5  g13946(.A(new_n16294), .B(n2421), .Y(new_n16295));
  not_8  g13947(.A(new_n16295), .Y(new_n16296));
  nand_5 g13948(.A(new_n16294), .B(n2421), .Y(new_n16297));
  and_5  g13949(.A(new_n16297), .B(new_n16296), .Y(new_n16298));
  or_5   g13950(.A(new_n16298), .B(n22198), .Y(new_n16299));
  nand_5 g13951(.A(new_n16298), .B(n22198), .Y(new_n16300));
  nand_5 g13952(.A(new_n10932), .B(n987), .Y(new_n16301));
  and_5  g13953(.A(new_n16301), .B(new_n16294), .Y(new_n16302));
  or_5   g13954(.A(new_n16302), .B(n20826), .Y(new_n16303));
  nand_5 g13955(.A(new_n16302), .B(n20826), .Y(new_n16304));
  nand_5 g13956(.A(new_n10936), .B(new_n10930), .Y(new_n16305));
  nand_5 g13957(.A(new_n16305), .B(new_n10935), .Y(new_n16306));
  nand_5 g13958(.A(new_n16306), .B(new_n16304), .Y(new_n16307));
  nand_5 g13959(.A(new_n16307), .B(new_n16303), .Y(new_n16308));
  nand_5 g13960(.A(new_n16308), .B(new_n16300), .Y(new_n16309));
  nand_5 g13961(.A(new_n16309), .B(new_n16299), .Y(new_n16310));
  nand_5 g13962(.A(new_n16295), .B(new_n6808), .Y(new_n16311));
  nand_5 g13963(.A(new_n16296), .B(n11044), .Y(new_n16312));
  and_5  g13964(.A(new_n16312), .B(new_n16311), .Y(new_n16313));
  or_5   g13965(.A(new_n16313), .B(n24327), .Y(new_n16314));
  nand_5 g13966(.A(new_n16313), .B(n24327), .Y(new_n16315));
  nand_5 g13967(.A(new_n16315), .B(new_n16314), .Y(new_n16316));
  xor_4  g13968(.A(new_n16316), .B(new_n16310), .Y(new_n16317));
  nand_5 g13969(.A(new_n16317), .B(new_n3925_1), .Y(new_n16318));
  not_8  g13970(.A(new_n16317), .Y(new_n16319));
  nand_5 g13971(.A(new_n16319), .B(new_n3928), .Y(new_n16320));
  nand_5 g13972(.A(new_n16300), .B(new_n16299), .Y(new_n16321));
  xor_4  g13973(.A(new_n16321), .B(new_n16308), .Y(new_n16322_1));
  nand_5 g13974(.A(new_n16322_1), .B(new_n3931), .Y(new_n16323));
  not_8  g13975(.A(new_n16322_1), .Y(new_n16324));
  nand_5 g13976(.A(new_n16324), .B(new_n3934_1), .Y(new_n16325));
  nand_5 g13977(.A(new_n16304), .B(new_n16303), .Y(new_n16326));
  xor_4  g13978(.A(new_n16326), .B(new_n16306), .Y(new_n16327_1));
  nand_5 g13979(.A(new_n16327_1), .B(new_n3937), .Y(new_n16328));
  not_8  g13980(.A(new_n16327_1), .Y(new_n16329));
  nand_5 g13981(.A(new_n16329), .B(new_n3940), .Y(new_n16330));
  nand_5 g13982(.A(new_n10938), .B(new_n3943), .Y(new_n16331));
  nand_5 g13983(.A(new_n10939), .B(new_n3946), .Y(new_n16332));
  nand_5 g13984(.A(new_n10892), .B(new_n3949), .Y(new_n16333));
  nand_5 g13985(.A(new_n10891), .B(new_n3952_1), .Y(new_n16334));
  nand_5 g13986(.A(new_n10859), .B(new_n3955), .Y(new_n16335));
  nand_5 g13987(.A(new_n10917), .B(new_n3954), .Y(new_n16336));
  nand_5 g13988(.A(new_n10863), .B(new_n3962_1), .Y(new_n16337));
  not_8  g13989(.A(new_n16337), .Y(new_n16338));
  nand_5 g13990(.A(new_n16338), .B(new_n16336), .Y(new_n16339));
  nand_5 g13991(.A(new_n16339), .B(new_n16335), .Y(new_n16340));
  nand_5 g13992(.A(new_n16340), .B(new_n16334), .Y(new_n16341));
  nand_5 g13993(.A(new_n16341), .B(new_n16333), .Y(new_n16342));
  nand_5 g13994(.A(new_n16342), .B(new_n16332), .Y(new_n16343));
  nand_5 g13995(.A(new_n16343), .B(new_n16331), .Y(new_n16344));
  nand_5 g13996(.A(new_n16344), .B(new_n16330), .Y(new_n16345));
  nand_5 g13997(.A(new_n16345), .B(new_n16328), .Y(new_n16346));
  nand_5 g13998(.A(new_n16346), .B(new_n16325), .Y(new_n16347));
  nand_5 g13999(.A(new_n16347), .B(new_n16323), .Y(new_n16348));
  nand_5 g14000(.A(new_n16348), .B(new_n16320), .Y(new_n16349));
  nand_5 g14001(.A(new_n16349), .B(new_n16318), .Y(new_n16350_1));
  nand_5 g14002(.A(new_n16315), .B(new_n16310), .Y(new_n16351));
  nand_5 g14003(.A(new_n16351), .B(new_n16314), .Y(new_n16352));
  nor_5  g14004(.A(new_n16311), .B(n5031), .Y(new_n16353));
  not_8  g14005(.A(new_n16353), .Y(new_n16354));
  nand_5 g14006(.A(new_n16311), .B(n5031), .Y(new_n16355));
  and_5  g14007(.A(new_n16355), .B(new_n16354), .Y(new_n16356));
  or_5   g14008(.A(new_n16356), .B(n2659), .Y(new_n16357));
  nand_5 g14009(.A(new_n16356), .B(n2659), .Y(new_n16358));
  nand_5 g14010(.A(new_n16358), .B(new_n16357), .Y(new_n16359));
  xor_4  g14011(.A(new_n16359), .B(new_n16352), .Y(new_n16360));
  nand_5 g14012(.A(new_n16360), .B(new_n3919), .Y(new_n16361));
  not_8  g14013(.A(new_n16360), .Y(new_n16362));
  nand_5 g14014(.A(new_n16362), .B(new_n3922), .Y(new_n16363));
  nand_5 g14015(.A(new_n16363), .B(new_n16361), .Y(new_n16364));
  xor_4  g14016(.A(new_n16364), .B(new_n16350_1), .Y(new_n16365));
  not_8  g14017(.A(new_n16365), .Y(new_n16366));
  or_5   g14018(.A(new_n16366), .B(new_n16293), .Y(new_n16367_1));
  not_8  g14019(.A(new_n16367_1), .Y(new_n16368));
  nand_5 g14020(.A(new_n16366), .B(new_n16293), .Y(new_n16369));
  not_8  g14021(.A(new_n16369), .Y(new_n16370));
  nand_5 g14022(.A(new_n16266), .B(new_n16265), .Y(new_n16371));
  xor_4  g14023(.A(new_n16371), .B(new_n16287), .Y(new_n16372));
  nand_5 g14024(.A(new_n16320), .B(new_n16318), .Y(new_n16373));
  xor_4  g14025(.A(new_n16373), .B(new_n16348), .Y(new_n16374));
  not_8  g14026(.A(new_n16374), .Y(new_n16375));
  or_5   g14027(.A(new_n16375), .B(new_n16372), .Y(new_n16376_1));
  not_8  g14028(.A(new_n16376_1), .Y(new_n16377));
  nand_5 g14029(.A(new_n16375), .B(new_n16372), .Y(new_n16378));
  not_8  g14030(.A(new_n16378), .Y(new_n16379_1));
  nand_5 g14031(.A(new_n16268), .B(new_n16267), .Y(new_n16380));
  xor_4  g14032(.A(new_n16380), .B(new_n16285), .Y(new_n16381));
  nand_5 g14033(.A(new_n16325), .B(new_n16323), .Y(new_n16382));
  xor_4  g14034(.A(new_n16382), .B(new_n16346), .Y(new_n16383));
  not_8  g14035(.A(new_n16383), .Y(new_n16384));
  nand_5 g14036(.A(new_n16384), .B(new_n16381), .Y(new_n16385));
  or_5   g14037(.A(new_n16384), .B(new_n16381), .Y(new_n16386));
  nand_5 g14038(.A(new_n16270), .B(new_n16269), .Y(new_n16387));
  xor_4  g14039(.A(new_n16387), .B(new_n16283), .Y(new_n16388));
  nand_5 g14040(.A(new_n16330), .B(new_n16328), .Y(new_n16389));
  xor_4  g14041(.A(new_n16389), .B(new_n16344), .Y(new_n16390));
  not_8  g14042(.A(new_n16390), .Y(new_n16391));
  nand_5 g14043(.A(new_n16391), .B(new_n16388), .Y(new_n16392));
  nor_5  g14044(.A(new_n16391), .B(new_n16388), .Y(new_n16393));
  not_8  g14045(.A(new_n16393), .Y(new_n16394));
  nand_5 g14046(.A(new_n16272), .B(new_n16271), .Y(new_n16395));
  xor_4  g14047(.A(new_n16395), .B(new_n16281), .Y(new_n16396_1));
  nand_5 g14048(.A(new_n16332), .B(new_n16331), .Y(new_n16397));
  xor_4  g14049(.A(new_n16397), .B(new_n16342), .Y(new_n16398_1));
  not_8  g14050(.A(new_n16398_1), .Y(new_n16399));
  nand_5 g14051(.A(new_n16399), .B(new_n16396_1), .Y(new_n16400));
  nor_5  g14052(.A(new_n16399), .B(new_n16396_1), .Y(new_n16401));
  not_8  g14053(.A(new_n16401), .Y(new_n16402));
  nand_5 g14054(.A(new_n16334), .B(new_n16333), .Y(new_n16403));
  xor_4  g14055(.A(new_n16403), .B(new_n16340), .Y(new_n16404));
  not_8  g14056(.A(new_n16404), .Y(new_n16405));
  nand_5 g14057(.A(new_n16274), .B(new_n16273), .Y(new_n16406_1));
  xor_4  g14058(.A(new_n16406_1), .B(new_n16279_1), .Y(new_n16407_1));
  nand_5 g14059(.A(new_n16407_1), .B(new_n16405), .Y(new_n16408));
  or_5   g14060(.A(new_n16407_1), .B(new_n16405), .Y(new_n16409));
  nor_5  g14061(.A(new_n10863), .B(new_n3962_1), .Y(new_n16410));
  nor_5  g14062(.A(new_n16410), .B(new_n16338), .Y(new_n16411));
  not_8  g14063(.A(new_n16411), .Y(new_n16412));
  nand_5 g14064(.A(new_n3697), .B(new_n3748), .Y(new_n16413));
  nand_5 g14065(.A(new_n16413), .B(new_n16277), .Y(new_n16414));
  nor_5  g14066(.A(new_n16414), .B(new_n16412), .Y(new_n16415));
  nand_5 g14067(.A(new_n16276), .B(new_n16275_1), .Y(new_n16416));
  nand_5 g14068(.A(new_n10917), .B(new_n3958), .Y(new_n16417));
  nand_5 g14069(.A(new_n16417), .B(new_n16335), .Y(new_n16418));
  xor_4  g14070(.A(new_n16418), .B(new_n16337), .Y(new_n16419_1));
  not_8  g14071(.A(new_n16419_1), .Y(new_n16420));
  nand_5 g14072(.A(new_n16420), .B(new_n16416), .Y(new_n16421));
  nand_5 g14073(.A(new_n16421), .B(new_n16415), .Y(new_n16422));
  xor_4  g14074(.A(new_n16416), .B(new_n16277), .Y(new_n16423));
  nand_5 g14075(.A(new_n16423), .B(new_n16419_1), .Y(new_n16424_1));
  nand_5 g14076(.A(new_n16424_1), .B(new_n16422), .Y(new_n16425));
  nand_5 g14077(.A(new_n16425), .B(new_n16409), .Y(new_n16426));
  nand_5 g14078(.A(new_n16426), .B(new_n16408), .Y(new_n16427));
  nand_5 g14079(.A(new_n16427), .B(new_n16402), .Y(new_n16428_1));
  nand_5 g14080(.A(new_n16428_1), .B(new_n16400), .Y(new_n16429));
  nand_5 g14081(.A(new_n16429), .B(new_n16394), .Y(new_n16430));
  nand_5 g14082(.A(new_n16430), .B(new_n16392), .Y(new_n16431));
  nand_5 g14083(.A(new_n16431), .B(new_n16386), .Y(new_n16432));
  nand_5 g14084(.A(new_n16432), .B(new_n16385), .Y(new_n16433_1));
  nor_5  g14085(.A(new_n16433_1), .B(new_n16379_1), .Y(new_n16434));
  nor_5  g14086(.A(new_n16434), .B(new_n16377), .Y(new_n16435));
  nor_5  g14087(.A(new_n16435), .B(new_n16370), .Y(new_n16436));
  nor_5  g14088(.A(new_n16436), .B(new_n16368), .Y(new_n16437));
  nand_5 g14089(.A(new_n16363), .B(new_n16350_1), .Y(new_n16438));
  nand_5 g14090(.A(new_n16438), .B(new_n16361), .Y(new_n16439_1));
  nand_5 g14091(.A(new_n16358), .B(new_n16352), .Y(new_n16440_1));
  nand_5 g14092(.A(new_n16440_1), .B(new_n16357), .Y(new_n16441));
  nand_5 g14093(.A(new_n16353), .B(new_n6799), .Y(new_n16442));
  nand_5 g14094(.A(new_n16354), .B(n2145), .Y(new_n16443));
  and_5  g14095(.A(new_n16443), .B(new_n16442), .Y(new_n16444));
  or_5   g14096(.A(new_n16444), .B(n2858), .Y(new_n16445_1));
  nand_5 g14097(.A(new_n16444), .B(n2858), .Y(new_n16446));
  nand_5 g14098(.A(new_n16446), .B(new_n16445_1), .Y(new_n16447));
  xor_4  g14099(.A(new_n16447), .B(new_n16441), .Y(new_n16448));
  nand_5 g14100(.A(new_n16448), .B(new_n3913), .Y(new_n16449));
  not_8  g14101(.A(new_n16448), .Y(new_n16450));
  nand_5 g14102(.A(new_n16450), .B(new_n3916), .Y(new_n16451));
  nand_5 g14103(.A(new_n16451), .B(new_n16449), .Y(new_n16452));
  xor_4  g14104(.A(new_n16452), .B(new_n16439_1), .Y(new_n16453));
  not_8  g14105(.A(new_n16453), .Y(new_n16454));
  nand_5 g14106(.A(new_n16291), .B(new_n16289), .Y(new_n16455));
  nand_5 g14107(.A(new_n16455), .B(new_n16290), .Y(new_n16456));
  nand_5 g14108(.A(new_n3773), .B(new_n3718), .Y(new_n16457));
  or_5   g14109(.A(new_n3773), .B(new_n3718), .Y(new_n16458));
  nand_5 g14110(.A(new_n16458), .B(new_n16457), .Y(new_n16459));
  xor_4  g14111(.A(new_n16459), .B(new_n16456), .Y(new_n16460_1));
  or_5   g14112(.A(new_n16460_1), .B(new_n16454), .Y(new_n16461));
  not_8  g14113(.A(new_n16461), .Y(new_n16462));
  nand_5 g14114(.A(new_n16460_1), .B(new_n16454), .Y(new_n16463));
  not_8  g14115(.A(new_n16463), .Y(new_n16464));
  nor_5  g14116(.A(new_n16464), .B(new_n16462), .Y(new_n16465));
  xor_4  g14117(.A(new_n16465), .B(new_n16437), .Y(n2779));
  not_8  g14118(.A(n25586), .Y(new_n16467));
  nand_5 g14119(.A(new_n11857), .B(new_n16467), .Y(new_n16468));
  nand_5 g14120(.A(new_n11855), .B(n25586), .Y(new_n16469));
  nand_5 g14121(.A(new_n16469), .B(new_n16468), .Y(new_n16470));
  not_8  g14122(.A(n25751), .Y(new_n16471));
  nand_5 g14123(.A(new_n11861), .B(new_n16471), .Y(new_n16472));
  nand_5 g14124(.A(new_n11860), .B(n25751), .Y(new_n16473));
  not_8  g14125(.A(n26053), .Y(new_n16474));
  nand_5 g14126(.A(new_n11865), .B(new_n16474), .Y(new_n16475));
  nand_5 g14127(.A(new_n11864), .B(n26053), .Y(new_n16476_1));
  not_8  g14128(.A(n7917), .Y(new_n16477));
  nand_5 g14129(.A(new_n11869), .B(new_n16477), .Y(new_n16478));
  nand_5 g14130(.A(new_n11868), .B(n7917), .Y(new_n16479));
  not_8  g14131(.A(n17302), .Y(new_n16480));
  nand_5 g14132(.A(new_n11873), .B(new_n16480), .Y(new_n16481_1));
  nand_5 g14133(.A(new_n11872), .B(n17302), .Y(new_n16482_1));
  not_8  g14134(.A(n2013), .Y(new_n16483));
  nand_5 g14135(.A(new_n11877), .B(new_n16483), .Y(new_n16484));
  nand_5 g14136(.A(new_n11876), .B(n2013), .Y(new_n16485));
  not_8  g14137(.A(n23755), .Y(new_n16486));
  nand_5 g14138(.A(new_n11881), .B(new_n16486), .Y(new_n16487));
  nand_5 g14139(.A(new_n11880), .B(n23755), .Y(new_n16488));
  not_8  g14140(.A(n19163), .Y(new_n16489));
  nand_5 g14141(.A(new_n11886), .B(new_n16489), .Y(new_n16490));
  nand_5 g14142(.A(new_n11885), .B(n19163), .Y(new_n16491));
  not_8  g14143(.A(n22358), .Y(new_n16492));
  nand_5 g14144(.A(new_n6588), .B(new_n16492), .Y(new_n16493_1));
  nand_5 g14145(.A(n25926), .B(n9646), .Y(new_n16494));
  nand_5 g14146(.A(new_n6587_1), .B(n22358), .Y(new_n16495));
  nand_5 g14147(.A(new_n16495), .B(new_n16494), .Y(new_n16496));
  nand_5 g14148(.A(new_n16496), .B(new_n16493_1), .Y(new_n16497));
  nand_5 g14149(.A(new_n16497), .B(new_n16491), .Y(new_n16498));
  nand_5 g14150(.A(new_n16498), .B(new_n16490), .Y(new_n16499));
  nand_5 g14151(.A(new_n16499), .B(new_n16488), .Y(new_n16500));
  nand_5 g14152(.A(new_n16500), .B(new_n16487), .Y(new_n16501));
  nand_5 g14153(.A(new_n16501), .B(new_n16485), .Y(new_n16502_1));
  nand_5 g14154(.A(new_n16502_1), .B(new_n16484), .Y(new_n16503));
  nand_5 g14155(.A(new_n16503), .B(new_n16482_1), .Y(new_n16504));
  nand_5 g14156(.A(new_n16504), .B(new_n16481_1), .Y(new_n16505));
  nand_5 g14157(.A(new_n16505), .B(new_n16479), .Y(new_n16506_1));
  nand_5 g14158(.A(new_n16506_1), .B(new_n16478), .Y(new_n16507_1));
  nand_5 g14159(.A(new_n16507_1), .B(new_n16476_1), .Y(new_n16508));
  nand_5 g14160(.A(new_n16508), .B(new_n16475), .Y(new_n16509));
  nand_5 g14161(.A(new_n16509), .B(new_n16473), .Y(new_n16510));
  nand_5 g14162(.A(new_n16510), .B(new_n16472), .Y(new_n16511));
  xor_4  g14163(.A(new_n16511), .B(new_n16470), .Y(new_n16512));
  not_8  g14164(.A(new_n16512), .Y(new_n16513));
  nand_5 g14165(.A(new_n16513), .B(n4514), .Y(new_n16514));
  nand_5 g14166(.A(new_n16512), .B(new_n13219), .Y(new_n16515));
  nand_5 g14167(.A(new_n16515), .B(new_n16514), .Y(new_n16516_1));
  nand_5 g14168(.A(new_n16473), .B(new_n16472), .Y(new_n16517_1));
  xor_4  g14169(.A(new_n16517_1), .B(new_n16509), .Y(new_n16518));
  nand_5 g14170(.A(new_n16518), .B(new_n13223), .Y(new_n16519));
  or_5   g14171(.A(new_n16518), .B(new_n13223), .Y(new_n16520));
  nand_5 g14172(.A(new_n16476_1), .B(new_n16475), .Y(new_n16521_1));
  xor_4  g14173(.A(new_n16521_1), .B(new_n16507_1), .Y(new_n16522));
  nand_5 g14174(.A(new_n16522), .B(new_n13228), .Y(new_n16523));
  or_5   g14175(.A(new_n16522), .B(new_n13228), .Y(new_n16524_1));
  nand_5 g14176(.A(new_n16479), .B(new_n16478), .Y(new_n16525));
  xor_4  g14177(.A(new_n16525), .B(new_n16505), .Y(new_n16526));
  nand_5 g14178(.A(new_n16526), .B(new_n12631), .Y(new_n16527_1));
  or_5   g14179(.A(new_n16526), .B(new_n12631), .Y(new_n16528));
  nand_5 g14180(.A(new_n16482_1), .B(new_n16481_1), .Y(new_n16529));
  xor_4  g14181(.A(new_n16529), .B(new_n16503), .Y(new_n16530));
  nand_5 g14182(.A(new_n16530), .B(new_n12540_1), .Y(new_n16531));
  or_5   g14183(.A(new_n16530), .B(new_n12540_1), .Y(new_n16532));
  nand_5 g14184(.A(new_n16485), .B(new_n16484), .Y(new_n16533));
  xor_4  g14185(.A(new_n16533), .B(new_n16501), .Y(new_n16534));
  nand_5 g14186(.A(new_n16534), .B(new_n11062), .Y(new_n16535));
  or_5   g14187(.A(new_n16534), .B(new_n11062), .Y(new_n16536));
  nand_5 g14188(.A(new_n16488), .B(new_n16487), .Y(new_n16537));
  xor_4  g14189(.A(new_n16537), .B(new_n16499), .Y(new_n16538));
  nand_5 g14190(.A(new_n16538), .B(new_n10983), .Y(new_n16539));
  nor_5  g14191(.A(new_n16538), .B(new_n10983), .Y(new_n16540));
  not_8  g14192(.A(new_n16540), .Y(new_n16541));
  nand_5 g14193(.A(new_n16491), .B(new_n16490), .Y(new_n16542));
  xor_4  g14194(.A(new_n16542), .B(new_n16497), .Y(new_n16543));
  nand_5 g14195(.A(new_n16543), .B(new_n10970), .Y(new_n16544_1));
  nor_5  g14196(.A(new_n16543), .B(new_n10970), .Y(new_n16545));
  not_8  g14197(.A(new_n16545), .Y(new_n16546));
  and_5  g14198(.A(new_n16495), .B(new_n16493_1), .Y(new_n16547));
  xor_4  g14199(.A(new_n16547), .B(new_n16494), .Y(new_n16548));
  nand_5 g14200(.A(new_n16548), .B(n26625), .Y(new_n16549));
  nand_5 g14201(.A(new_n16549), .B(new_n7512), .Y(new_n16550));
  or_5   g14202(.A(new_n16548), .B(n26625), .Y(new_n16551));
  nand_5 g14203(.A(new_n16551), .B(new_n16550), .Y(new_n16552));
  nand_5 g14204(.A(new_n16552), .B(new_n16546), .Y(new_n16553));
  nand_5 g14205(.A(new_n16553), .B(new_n16544_1), .Y(new_n16554_1));
  nand_5 g14206(.A(new_n16554_1), .B(new_n16541), .Y(new_n16555));
  nand_5 g14207(.A(new_n16555), .B(new_n16539), .Y(new_n16556));
  nand_5 g14208(.A(new_n16556), .B(new_n16536), .Y(new_n16557));
  nand_5 g14209(.A(new_n16557), .B(new_n16535), .Y(new_n16558));
  nand_5 g14210(.A(new_n16558), .B(new_n16532), .Y(new_n16559));
  nand_5 g14211(.A(new_n16559), .B(new_n16531), .Y(new_n16560));
  nand_5 g14212(.A(new_n16560), .B(new_n16528), .Y(new_n16561));
  nand_5 g14213(.A(new_n16561), .B(new_n16527_1), .Y(new_n16562));
  nand_5 g14214(.A(new_n16562), .B(new_n16524_1), .Y(new_n16563));
  nand_5 g14215(.A(new_n16563), .B(new_n16523), .Y(new_n16564));
  nand_5 g14216(.A(new_n16564), .B(new_n16520), .Y(new_n16565));
  nand_5 g14217(.A(new_n16565), .B(new_n16519), .Y(new_n16566));
  xnor_4 g14218(.A(new_n16566), .B(new_n16516_1), .Y(new_n16567));
  or_5   g14219(.A(new_n16567), .B(new_n12033), .Y(new_n16568));
  nand_5 g14220(.A(new_n16567), .B(new_n12033), .Y(new_n16569));
  nand_5 g14221(.A(new_n16520), .B(new_n16519), .Y(new_n16570));
  xor_4  g14222(.A(new_n16570), .B(new_n16564), .Y(new_n16571));
  nand_5 g14223(.A(new_n16571), .B(new_n12040), .Y(new_n16572));
  or_5   g14224(.A(new_n16571), .B(new_n12040), .Y(new_n16573));
  nand_5 g14225(.A(new_n16524_1), .B(new_n16523), .Y(new_n16574));
  xor_4  g14226(.A(new_n16574), .B(new_n16562), .Y(new_n16575));
  nand_5 g14227(.A(new_n16575), .B(new_n12047), .Y(new_n16576));
  or_5   g14228(.A(new_n16575), .B(new_n12047), .Y(new_n16577));
  nand_5 g14229(.A(new_n16528), .B(new_n16527_1), .Y(new_n16578));
  xnor_4 g14230(.A(new_n16578), .B(new_n16560), .Y(new_n16579));
  or_5   g14231(.A(new_n16579), .B(new_n12053), .Y(new_n16580));
  nand_5 g14232(.A(new_n16579), .B(new_n12053), .Y(new_n16581));
  nand_5 g14233(.A(new_n16532), .B(new_n16531), .Y(new_n16582));
  xnor_4 g14234(.A(new_n16582), .B(new_n16558), .Y(new_n16583_1));
  or_5   g14235(.A(new_n16583_1), .B(new_n12060), .Y(new_n16584_1));
  nand_5 g14236(.A(new_n16583_1), .B(new_n12060), .Y(new_n16585));
  nand_5 g14237(.A(new_n16536), .B(new_n16535), .Y(new_n16586));
  xor_4  g14238(.A(new_n16586), .B(new_n16556), .Y(new_n16587));
  or_5   g14239(.A(new_n16587), .B(new_n12069), .Y(new_n16588));
  nand_5 g14240(.A(new_n16587), .B(new_n12069), .Y(new_n16589_1));
  nand_5 g14241(.A(new_n16541), .B(new_n16539), .Y(new_n16590));
  xor_4  g14242(.A(new_n16590), .B(new_n16554_1), .Y(new_n16591));
  or_5   g14243(.A(new_n16591), .B(new_n12076), .Y(new_n16592));
  nand_5 g14244(.A(new_n16591), .B(new_n12076), .Y(new_n16593));
  nand_5 g14245(.A(new_n16546), .B(new_n16544_1), .Y(new_n16594));
  xor_4  g14246(.A(new_n16594), .B(new_n16552), .Y(new_n16595));
  or_5   g14247(.A(new_n16595), .B(new_n12085), .Y(new_n16596_1));
  nand_5 g14248(.A(new_n16595), .B(new_n12085), .Y(new_n16597));
  nand_5 g14249(.A(new_n7515), .B(new_n6576_1), .Y(new_n16598));
  nor_5  g14250(.A(new_n16598), .B(new_n6605), .Y(new_n16599));
  not_8  g14251(.A(new_n16599), .Y(new_n16600));
  not_8  g14252(.A(new_n6606), .Y(new_n16601));
  nand_5 g14253(.A(new_n16598), .B(new_n16601), .Y(new_n16602));
  nand_5 g14254(.A(new_n16551), .B(new_n16549), .Y(new_n16603));
  xnor_4 g14255(.A(new_n16603), .B(new_n7512), .Y(new_n16604));
  nand_5 g14256(.A(new_n16604), .B(new_n16602), .Y(new_n16605));
  nand_5 g14257(.A(new_n16605), .B(new_n16600), .Y(new_n16606));
  nand_5 g14258(.A(new_n16606), .B(new_n16597), .Y(new_n16607));
  nand_5 g14259(.A(new_n16607), .B(new_n16596_1), .Y(new_n16608_1));
  nand_5 g14260(.A(new_n16608_1), .B(new_n16593), .Y(new_n16609));
  nand_5 g14261(.A(new_n16609), .B(new_n16592), .Y(new_n16610));
  nand_5 g14262(.A(new_n16610), .B(new_n16589_1), .Y(new_n16611));
  nand_5 g14263(.A(new_n16611), .B(new_n16588), .Y(new_n16612));
  not_8  g14264(.A(new_n16612), .Y(new_n16613));
  nand_5 g14265(.A(new_n16613), .B(new_n16585), .Y(new_n16614));
  nand_5 g14266(.A(new_n16614), .B(new_n16584_1), .Y(new_n16615));
  nand_5 g14267(.A(new_n16615), .B(new_n16581), .Y(new_n16616));
  nand_5 g14268(.A(new_n16616), .B(new_n16580), .Y(new_n16617_1));
  nand_5 g14269(.A(new_n16617_1), .B(new_n16577), .Y(new_n16618));
  nand_5 g14270(.A(new_n16618), .B(new_n16576), .Y(new_n16619));
  nand_5 g14271(.A(new_n16619), .B(new_n16573), .Y(new_n16620));
  nand_5 g14272(.A(new_n16620), .B(new_n16572), .Y(new_n16621));
  nand_5 g14273(.A(new_n16621), .B(new_n16569), .Y(new_n16622));
  nand_5 g14274(.A(new_n16622), .B(new_n16568), .Y(new_n16623));
  nand_5 g14275(.A(new_n16623), .B(new_n12028), .Y(new_n16624));
  not_8  g14276(.A(new_n16624), .Y(new_n16625));
  nor_5  g14277(.A(new_n16623), .B(new_n12028), .Y(new_n16626));
  nor_5  g14278(.A(new_n16626), .B(new_n16625), .Y(new_n16627));
  not_8  g14279(.A(new_n16468), .Y(new_n16628));
  nor_5  g14280(.A(new_n16511), .B(new_n16628), .Y(new_n16629));
  nand_5 g14281(.A(new_n16469), .B(new_n11854), .Y(new_n16630_1));
  nor_5  g14282(.A(new_n16630_1), .B(new_n16629), .Y(new_n16631));
  nand_5 g14283(.A(new_n16566), .B(new_n16514), .Y(new_n16632));
  nand_5 g14284(.A(new_n16632), .B(new_n16515), .Y(new_n16633));
  xor_4  g14285(.A(new_n16633), .B(new_n16631), .Y(new_n16634));
  not_8  g14286(.A(new_n16634), .Y(new_n16635));
  xor_4  g14287(.A(new_n16635), .B(new_n16627), .Y(n2826));
  nand_5 g14288(.A(new_n2693_1), .B(new_n2646_1), .Y(new_n16637));
  nand_5 g14289(.A(new_n16637), .B(new_n2649), .Y(new_n16638));
  not_8  g14290(.A(new_n16638), .Y(new_n16639));
  nand_5 g14291(.A(new_n2764), .B(new_n2698), .Y(new_n16640_1));
  nand_5 g14292(.A(new_n16640_1), .B(new_n2697), .Y(new_n16641));
  nand_5 g14293(.A(new_n16641), .B(new_n16639), .Y(new_n16642));
  not_8  g14294(.A(new_n16642), .Y(new_n16643));
  nand_5 g14295(.A(new_n7092), .B(n5140), .Y(new_n16644));
  nand_5 g14296(.A(new_n7087), .B(new_n14201), .Y(new_n16645));
  nand_5 g14297(.A(new_n7100), .B(n6204), .Y(new_n16646));
  nand_5 g14298(.A(new_n7095), .B(new_n14204), .Y(new_n16647));
  nand_5 g14299(.A(new_n7108), .B(n3349), .Y(new_n16648));
  nand_5 g14300(.A(new_n7103), .B(new_n14207), .Y(new_n16649));
  nand_5 g14301(.A(new_n7116), .B(n1742), .Y(new_n16650));
  nand_5 g14302(.A(new_n7111), .B(new_n7491), .Y(new_n16651));
  not_8  g14303(.A(new_n7120), .Y(new_n16652));
  nand_5 g14304(.A(new_n16652), .B(n4858), .Y(new_n16653));
  nand_5 g14305(.A(new_n7120), .B(new_n7416), .Y(new_n16654));
  nand_5 g14306(.A(new_n7124), .B(n8244), .Y(new_n16655));
  nand_5 g14307(.A(new_n7125), .B(new_n7360), .Y(new_n16656_1));
  nand_5 g14308(.A(new_n7127), .B(n9493), .Y(new_n16657));
  nand_5 g14309(.A(new_n7128), .B(new_n7329), .Y(new_n16658));
  nand_5 g14310(.A(new_n7132), .B(n15167), .Y(new_n16659));
  nand_5 g14311(.A(new_n14168), .B(new_n7341), .Y(new_n16660));
  nand_5 g14312(.A(new_n7138), .B(n21095), .Y(new_n16661));
  nand_5 g14313(.A(new_n7137), .B(new_n7347), .Y(new_n16662));
  nand_5 g14314(.A(new_n7142), .B(n8656), .Y(new_n16663));
  not_8  g14315(.A(new_n16663), .Y(new_n16664));
  nand_5 g14316(.A(new_n16664), .B(new_n16662), .Y(new_n16665));
  nand_5 g14317(.A(new_n16665), .B(new_n16661), .Y(new_n16666));
  nand_5 g14318(.A(new_n16666), .B(new_n16660), .Y(new_n16667));
  nand_5 g14319(.A(new_n16667), .B(new_n16659), .Y(new_n16668));
  nand_5 g14320(.A(new_n16668), .B(new_n16658), .Y(new_n16669));
  nand_5 g14321(.A(new_n16669), .B(new_n16657), .Y(new_n16670));
  nand_5 g14322(.A(new_n16670), .B(new_n16656_1), .Y(new_n16671));
  nand_5 g14323(.A(new_n16671), .B(new_n16655), .Y(new_n16672));
  nand_5 g14324(.A(new_n16672), .B(new_n16654), .Y(new_n16673));
  nand_5 g14325(.A(new_n16673), .B(new_n16653), .Y(new_n16674_1));
  nand_5 g14326(.A(new_n16674_1), .B(new_n16651), .Y(new_n16675));
  nand_5 g14327(.A(new_n16675), .B(new_n16650), .Y(new_n16676));
  nand_5 g14328(.A(new_n16676), .B(new_n16649), .Y(new_n16677));
  nand_5 g14329(.A(new_n16677), .B(new_n16648), .Y(new_n16678));
  nand_5 g14330(.A(new_n16678), .B(new_n16647), .Y(new_n16679));
  nand_5 g14331(.A(new_n16679), .B(new_n16646), .Y(new_n16680));
  nand_5 g14332(.A(new_n16680), .B(new_n16645), .Y(new_n16681));
  nand_5 g14333(.A(new_n16681), .B(new_n16644), .Y(new_n16682_1));
  nand_5 g14334(.A(new_n16682_1), .B(new_n7044), .Y(new_n16683));
  nand_5 g14335(.A(new_n16683), .B(new_n16643), .Y(new_n16684_1));
  or_5   g14336(.A(new_n16683), .B(new_n16643), .Y(new_n16685));
  nand_5 g14337(.A(new_n16685), .B(new_n16684_1), .Y(new_n16686));
  or_5   g14338(.A(new_n16641), .B(new_n16639), .Y(new_n16687));
  and_5  g14339(.A(new_n16687), .B(new_n16642), .Y(new_n16688_1));
  not_8  g14340(.A(new_n16688_1), .Y(new_n16689));
  xor_4  g14341(.A(new_n16682_1), .B(new_n7044), .Y(new_n16690));
  nand_5 g14342(.A(new_n16690), .B(new_n16689), .Y(new_n16691));
  not_8  g14343(.A(new_n16691), .Y(new_n16692));
  nor_5  g14344(.A(new_n16690), .B(new_n16689), .Y(new_n16693));
  not_8  g14345(.A(new_n2765), .Y(new_n16694));
  nand_5 g14346(.A(new_n16644), .B(new_n16645), .Y(new_n16695));
  xor_4  g14347(.A(new_n16695), .B(new_n16680), .Y(new_n16696));
  or_5   g14348(.A(new_n16696), .B(new_n16694), .Y(new_n16697));
  nand_5 g14349(.A(new_n16696), .B(new_n16694), .Y(new_n16698));
  nand_5 g14350(.A(new_n16646), .B(new_n16647), .Y(new_n16699));
  xor_4  g14351(.A(new_n16699), .B(new_n16678), .Y(new_n16700));
  or_5   g14352(.A(new_n16700), .B(new_n2918), .Y(new_n16701));
  nand_5 g14353(.A(new_n16700), .B(new_n2918), .Y(new_n16702));
  nand_5 g14354(.A(new_n16648), .B(new_n16649), .Y(new_n16703));
  xor_4  g14355(.A(new_n16703), .B(new_n16676), .Y(new_n16704));
  not_8  g14356(.A(new_n16704), .Y(new_n16705));
  nand_5 g14357(.A(new_n16705), .B(new_n2924), .Y(new_n16706));
  not_8  g14358(.A(new_n16706), .Y(new_n16707));
  nand_5 g14359(.A(new_n16704), .B(new_n2925), .Y(new_n16708));
  not_8  g14360(.A(new_n16708), .Y(new_n16709));
  nand_5 g14361(.A(new_n16650), .B(new_n16651), .Y(new_n16710));
  xor_4  g14362(.A(new_n16710), .B(new_n16674_1), .Y(new_n16711));
  nand_5 g14363(.A(new_n16711), .B(new_n2932), .Y(new_n16712));
  or_5   g14364(.A(new_n16711), .B(new_n2932), .Y(new_n16713));
  nand_5 g14365(.A(new_n16653), .B(new_n16654), .Y(new_n16714));
  xor_4  g14366(.A(new_n16714), .B(new_n16672), .Y(new_n16715));
  nand_5 g14367(.A(new_n16715), .B(new_n2939), .Y(new_n16716));
  nor_5  g14368(.A(new_n16715), .B(new_n2939), .Y(new_n16717));
  not_8  g14369(.A(new_n16717), .Y(new_n16718));
  nand_5 g14370(.A(new_n16655), .B(new_n16656_1), .Y(new_n16719));
  xor_4  g14371(.A(new_n16719), .B(new_n16670), .Y(new_n16720));
  nand_5 g14372(.A(new_n16720), .B(new_n2946), .Y(new_n16721));
  not_8  g14373(.A(new_n16721), .Y(new_n16722_1));
  nor_5  g14374(.A(new_n16720), .B(new_n2946), .Y(new_n16723));
  nand_5 g14375(.A(new_n16657), .B(new_n16658), .Y(new_n16724));
  xor_4  g14376(.A(new_n16724), .B(new_n16668), .Y(new_n16725));
  nand_5 g14377(.A(new_n16725), .B(new_n2953), .Y(new_n16726));
  not_8  g14378(.A(new_n16726), .Y(new_n16727));
  nor_5  g14379(.A(new_n16725), .B(new_n2953), .Y(new_n16728));
  nand_5 g14380(.A(new_n16659), .B(new_n16660), .Y(new_n16729));
  xor_4  g14381(.A(new_n16729), .B(new_n16666), .Y(new_n16730));
  nand_5 g14382(.A(new_n16730), .B(new_n2960), .Y(new_n16731));
  not_8  g14383(.A(new_n16731), .Y(new_n16732));
  nor_5  g14384(.A(new_n16730), .B(new_n2960), .Y(new_n16733_1));
  nand_5 g14385(.A(new_n16661), .B(new_n16662), .Y(new_n16734));
  xor_4  g14386(.A(new_n16734), .B(new_n16664), .Y(new_n16735));
  nand_5 g14387(.A(new_n16735), .B(new_n2969), .Y(new_n16736));
  not_8  g14388(.A(new_n16735), .Y(new_n16737));
  nand_5 g14389(.A(new_n16737), .B(new_n2967), .Y(new_n16738));
  or_5   g14390(.A(new_n7142), .B(n8656), .Y(new_n16739));
  nand_5 g14391(.A(new_n16739), .B(new_n16663), .Y(new_n16740));
  nand_5 g14392(.A(new_n16740), .B(new_n2976), .Y(new_n16741));
  not_8  g14393(.A(new_n16741), .Y(new_n16742));
  nand_5 g14394(.A(new_n16742), .B(new_n16738), .Y(new_n16743_1));
  nand_5 g14395(.A(new_n16743_1), .B(new_n16736), .Y(new_n16744));
  not_8  g14396(.A(new_n16744), .Y(new_n16745));
  nor_5  g14397(.A(new_n16745), .B(new_n16733_1), .Y(new_n16746));
  nor_5  g14398(.A(new_n16746), .B(new_n16732), .Y(new_n16747));
  nor_5  g14399(.A(new_n16747), .B(new_n16728), .Y(new_n16748));
  nor_5  g14400(.A(new_n16748), .B(new_n16727), .Y(new_n16749));
  nor_5  g14401(.A(new_n16749), .B(new_n16723), .Y(new_n16750));
  nor_5  g14402(.A(new_n16750), .B(new_n16722_1), .Y(new_n16751));
  not_8  g14403(.A(new_n16751), .Y(new_n16752));
  nand_5 g14404(.A(new_n16752), .B(new_n16718), .Y(new_n16753));
  nand_5 g14405(.A(new_n16753), .B(new_n16716), .Y(new_n16754));
  nand_5 g14406(.A(new_n16754), .B(new_n16713), .Y(new_n16755));
  nand_5 g14407(.A(new_n16755), .B(new_n16712), .Y(new_n16756));
  nor_5  g14408(.A(new_n16756), .B(new_n16709), .Y(new_n16757));
  nor_5  g14409(.A(new_n16757), .B(new_n16707), .Y(new_n16758));
  not_8  g14410(.A(new_n16758), .Y(new_n16759));
  nand_5 g14411(.A(new_n16759), .B(new_n16702), .Y(new_n16760));
  nand_5 g14412(.A(new_n16760), .B(new_n16701), .Y(new_n16761));
  nand_5 g14413(.A(new_n16761), .B(new_n16698), .Y(new_n16762));
  nand_5 g14414(.A(new_n16762), .B(new_n16697), .Y(new_n16763));
  not_8  g14415(.A(new_n16763), .Y(new_n16764));
  nor_5  g14416(.A(new_n16764), .B(new_n16693), .Y(new_n16765));
  nor_5  g14417(.A(new_n16765), .B(new_n16692), .Y(new_n16766));
  xor_4  g14418(.A(new_n16766), .B(new_n16686), .Y(n2853));
  nand_5 g14419(.A(new_n3007), .B(n1118), .Y(new_n16768));
  nand_5 g14420(.A(n4665), .B(new_n3042), .Y(new_n16769));
  nand_5 g14421(.A(n25974), .B(new_n3010_1), .Y(new_n16770));
  nand_5 g14422(.A(new_n3047), .B(n19005), .Y(new_n16771));
  nand_5 g14423(.A(new_n3013), .B(n1630), .Y(new_n16772));
  nand_5 g14424(.A(n4326), .B(new_n3050), .Y(new_n16773));
  nand_5 g14425(.A(n5438), .B(new_n3158), .Y(new_n16774));
  nand_5 g14426(.A(new_n16774), .B(new_n16773), .Y(new_n16775));
  nand_5 g14427(.A(new_n16775), .B(new_n16772), .Y(new_n16776));
  nand_5 g14428(.A(new_n16776), .B(new_n16771), .Y(new_n16777));
  nand_5 g14429(.A(new_n16777), .B(new_n16770), .Y(new_n16778));
  nand_5 g14430(.A(new_n16778), .B(new_n16769), .Y(new_n16779));
  nand_5 g14431(.A(new_n16779), .B(new_n16768), .Y(new_n16780));
  nand_5 g14432(.A(n12811), .B(new_n3004), .Y(new_n16781));
  nand_5 g14433(.A(new_n3039), .B(n5213), .Y(new_n16782));
  nand_5 g14434(.A(new_n16782), .B(new_n16781), .Y(new_n16783));
  xor_4  g14435(.A(new_n16783), .B(new_n16780), .Y(new_n16784));
  nand_5 g14436(.A(new_n16784), .B(new_n4806), .Y(new_n16785));
  nor_5  g14437(.A(new_n16784), .B(new_n4806), .Y(new_n16786));
  not_8  g14438(.A(new_n16786), .Y(new_n16787));
  nand_5 g14439(.A(new_n16769), .B(new_n16768), .Y(new_n16788));
  xor_4  g14440(.A(new_n16788), .B(new_n16778), .Y(new_n16789));
  nand_5 g14441(.A(new_n16789), .B(new_n4734), .Y(new_n16790));
  nor_5  g14442(.A(new_n16789), .B(new_n4734), .Y(new_n16791));
  not_8  g14443(.A(new_n16791), .Y(new_n16792));
  nand_5 g14444(.A(new_n16771), .B(new_n16770), .Y(new_n16793));
  xor_4  g14445(.A(new_n16793), .B(new_n16776), .Y(new_n16794));
  nand_5 g14446(.A(new_n16794), .B(new_n4739), .Y(new_n16795));
  nor_5  g14447(.A(new_n16794), .B(new_n4739), .Y(new_n16796));
  not_8  g14448(.A(new_n16796), .Y(new_n16797));
  nand_5 g14449(.A(new_n3015), .B(n1451), .Y(new_n16798_1));
  nand_5 g14450(.A(new_n16798_1), .B(new_n16774), .Y(new_n16799));
  nand_5 g14451(.A(new_n16799), .B(new_n4754), .Y(new_n16800));
  nand_5 g14452(.A(new_n16800), .B(new_n4750), .Y(new_n16801));
  nor_5  g14453(.A(new_n16800), .B(new_n4749), .Y(new_n16802));
  not_8  g14454(.A(new_n16802), .Y(new_n16803));
  nand_5 g14455(.A(new_n16773), .B(new_n16772), .Y(new_n16804));
  xor_4  g14456(.A(new_n16804), .B(new_n16774), .Y(new_n16805));
  nand_5 g14457(.A(new_n16805), .B(new_n16803), .Y(new_n16806));
  nand_5 g14458(.A(new_n16806), .B(new_n16801), .Y(new_n16807));
  nand_5 g14459(.A(new_n16807), .B(new_n16797), .Y(new_n16808));
  nand_5 g14460(.A(new_n16808), .B(new_n16795), .Y(new_n16809));
  nand_5 g14461(.A(new_n16809), .B(new_n16792), .Y(new_n16810));
  nand_5 g14462(.A(new_n16810), .B(new_n16790), .Y(new_n16811));
  nand_5 g14463(.A(new_n16811), .B(new_n16787), .Y(new_n16812_1));
  nand_5 g14464(.A(new_n16812_1), .B(new_n16785), .Y(new_n16813));
  nand_5 g14465(.A(new_n4803), .B(new_n4779), .Y(new_n16814));
  nand_5 g14466(.A(new_n16814), .B(new_n4801), .Y(new_n16815));
  nand_5 g14467(.A(new_n4786), .B(new_n4781), .Y(new_n16816));
  nand_5 g14468(.A(new_n16816), .B(new_n4785_1), .Y(new_n16817));
  nand_5 g14469(.A(new_n4783), .B(new_n4782), .Y(new_n16818_1));
  xor_4  g14470(.A(new_n16818_1), .B(n3570), .Y(new_n16819));
  or_5   g14471(.A(new_n16819), .B(n5337), .Y(new_n16820));
  nand_5 g14472(.A(new_n16819), .B(n5337), .Y(new_n16821));
  nand_5 g14473(.A(new_n16821), .B(new_n16820), .Y(new_n16822));
  xor_4  g14474(.A(new_n16822), .B(new_n16817), .Y(new_n16823));
  or_5   g14475(.A(new_n16823), .B(new_n12771), .Y(new_n16824_1));
  nand_5 g14476(.A(new_n16823), .B(new_n12771), .Y(new_n16825));
  nand_5 g14477(.A(new_n16825), .B(new_n16824_1), .Y(new_n16826));
  xor_4  g14478(.A(new_n16826), .B(new_n16815), .Y(new_n16827));
  nand_5 g14479(.A(new_n16782), .B(new_n16780), .Y(new_n16828));
  nand_5 g14480(.A(new_n16828), .B(new_n16781), .Y(new_n16829));
  not_8  g14481(.A(new_n16829), .Y(new_n16830));
  nand_5 g14482(.A(n7099), .B(new_n3000), .Y(new_n16831));
  nand_5 g14483(.A(new_n3034), .B(n2035), .Y(new_n16832));
  nand_5 g14484(.A(new_n16832), .B(new_n16831), .Y(new_n16833));
  xor_4  g14485(.A(new_n16833), .B(new_n16830), .Y(new_n16834_1));
  or_5   g14486(.A(new_n16834_1), .B(new_n16827), .Y(new_n16835));
  nand_5 g14487(.A(new_n16834_1), .B(new_n16827), .Y(new_n16836));
  nand_5 g14488(.A(new_n16836), .B(new_n16835), .Y(new_n16837_1));
  xor_4  g14489(.A(new_n16837_1), .B(new_n16813), .Y(n2860));
  nand_5 g14490(.A(new_n15778), .B(new_n15777), .Y(new_n16839));
  xor_4  g14491(.A(new_n16839), .B(new_n15802), .Y(n2887));
  nor_5  g14492(.A(new_n16818_1), .B(n3570), .Y(new_n16841_1));
  nand_5 g14493(.A(new_n16841_1), .B(new_n6861_1), .Y(new_n16842));
  nor_5  g14494(.A(new_n16842), .B(n20359), .Y(new_n16843));
  xor_4  g14495(.A(new_n16843), .B(n2816), .Y(new_n16844));
  nand_5 g14496(.A(new_n16844), .B(new_n6800), .Y(new_n16845));
  or_5   g14497(.A(new_n16844), .B(new_n6800), .Y(new_n16846));
  xor_4  g14498(.A(new_n16842), .B(new_n6855), .Y(new_n16847));
  nand_5 g14499(.A(new_n16847), .B(new_n6804), .Y(new_n16848));
  or_5   g14500(.A(new_n16847), .B(new_n6804), .Y(new_n16849));
  xor_4  g14501(.A(new_n16841_1), .B(new_n6861_1), .Y(new_n16850));
  or_5   g14502(.A(new_n16850), .B(n4325), .Y(new_n16851));
  nand_5 g14503(.A(new_n16850), .B(n4325), .Y(new_n16852));
  nand_5 g14504(.A(new_n16821), .B(new_n16817), .Y(new_n16853));
  nand_5 g14505(.A(new_n16853), .B(new_n16820), .Y(new_n16854));
  nand_5 g14506(.A(new_n16854), .B(new_n16852), .Y(new_n16855));
  nand_5 g14507(.A(new_n16855), .B(new_n16851), .Y(new_n16856));
  nand_5 g14508(.A(new_n16856), .B(new_n16849), .Y(new_n16857));
  nand_5 g14509(.A(new_n16857), .B(new_n16848), .Y(new_n16858));
  nand_5 g14510(.A(new_n16858), .B(new_n16846), .Y(new_n16859));
  nand_5 g14511(.A(new_n16859), .B(new_n16845), .Y(new_n16860));
  nand_5 g14512(.A(new_n16843), .B(new_n6849), .Y(new_n16861));
  xor_4  g14513(.A(new_n16861), .B(n8526), .Y(new_n16862));
  nor_5  g14514(.A(new_n16862), .B(n21784), .Y(new_n16863));
  nor_5  g14515(.A(new_n16863), .B(new_n16860), .Y(new_n16864));
  or_5   g14516(.A(new_n16861), .B(n8526), .Y(new_n16865));
  nand_5 g14517(.A(new_n16862), .B(n21784), .Y(new_n16866));
  nand_5 g14518(.A(new_n16866), .B(new_n16865), .Y(new_n16867));
  nor_5  g14519(.A(new_n16867), .B(new_n16864), .Y(new_n16868));
  nand_5 g14520(.A(new_n16868), .B(new_n12732), .Y(new_n16869));
  not_8  g14521(.A(new_n16868), .Y(new_n16870));
  nand_5 g14522(.A(new_n16870), .B(new_n12733), .Y(new_n16871));
  nand_5 g14523(.A(new_n16871), .B(new_n16869), .Y(new_n16872));
  xor_4  g14524(.A(new_n16862), .B(n21784), .Y(new_n16873));
  xor_4  g14525(.A(new_n16873), .B(new_n16860), .Y(new_n16874));
  not_8  g14526(.A(new_n16874), .Y(new_n16875));
  nand_5 g14527(.A(new_n16875), .B(new_n12742_1), .Y(new_n16876));
  nand_5 g14528(.A(new_n16874), .B(new_n12743), .Y(new_n16877));
  nand_5 g14529(.A(new_n16846), .B(new_n16845), .Y(new_n16878));
  xor_4  g14530(.A(new_n16878), .B(new_n16858), .Y(new_n16879));
  nand_5 g14531(.A(new_n16879), .B(new_n12750), .Y(new_n16880));
  not_8  g14532(.A(new_n16879), .Y(new_n16881));
  nand_5 g14533(.A(new_n16881), .B(new_n12751), .Y(new_n16882));
  nand_5 g14534(.A(new_n16849), .B(new_n16848), .Y(new_n16883));
  xor_4  g14535(.A(new_n16883), .B(new_n16856), .Y(new_n16884));
  nand_5 g14536(.A(new_n16884), .B(new_n12757), .Y(new_n16885_1));
  not_8  g14537(.A(new_n16884), .Y(new_n16886));
  nand_5 g14538(.A(new_n16886), .B(new_n12758), .Y(new_n16887));
  nand_5 g14539(.A(new_n16852), .B(new_n16851), .Y(new_n16888));
  xor_4  g14540(.A(new_n16888), .B(new_n16854), .Y(new_n16889));
  nand_5 g14541(.A(new_n16889), .B(new_n12764), .Y(new_n16890));
  or_5   g14542(.A(new_n16889), .B(new_n12764), .Y(new_n16891));
  nand_5 g14543(.A(new_n16825), .B(new_n16815), .Y(new_n16892));
  nand_5 g14544(.A(new_n16892), .B(new_n16824_1), .Y(new_n16893));
  not_8  g14545(.A(new_n16893), .Y(new_n16894));
  nand_5 g14546(.A(new_n16894), .B(new_n16891), .Y(new_n16895));
  nand_5 g14547(.A(new_n16895), .B(new_n16890), .Y(new_n16896));
  nand_5 g14548(.A(new_n16896), .B(new_n16887), .Y(new_n16897));
  nand_5 g14549(.A(new_n16897), .B(new_n16885_1), .Y(new_n16898));
  nand_5 g14550(.A(new_n16898), .B(new_n16882), .Y(new_n16899));
  nand_5 g14551(.A(new_n16899), .B(new_n16880), .Y(new_n16900));
  nand_5 g14552(.A(new_n16900), .B(new_n16877), .Y(new_n16901));
  nand_5 g14553(.A(new_n16901), .B(new_n16876), .Y(new_n16902));
  nand_5 g14554(.A(new_n16902), .B(new_n16872), .Y(new_n16903));
  nor_5  g14555(.A(new_n16902), .B(new_n16872), .Y(new_n16904));
  not_8  g14556(.A(new_n16904), .Y(new_n16905_1));
  and_5  g14557(.A(new_n16905_1), .B(new_n16903), .Y(new_n16906));
  not_8  g14558(.A(new_n16906), .Y(new_n16907));
  not_8  g14559(.A(new_n4770_1), .Y(new_n16908));
  nand_5 g14560(.A(new_n16908), .B(new_n12136), .Y(new_n16909));
  or_5   g14561(.A(new_n16909), .B(n15546), .Y(new_n16910));
  nor_5  g14562(.A(new_n16910), .B(n5077), .Y(new_n16911_1));
  nand_5 g14563(.A(new_n16911_1), .B(new_n12392), .Y(new_n16912));
  nor_5  g14564(.A(new_n16912), .B(n8827), .Y(new_n16913));
  not_8  g14565(.A(new_n16913), .Y(new_n16914));
  nand_5 g14566(.A(new_n16912), .B(n8827), .Y(new_n16915));
  nand_5 g14567(.A(new_n16915), .B(new_n16914), .Y(new_n16916));
  nand_5 g14568(.A(new_n16916), .B(new_n8431), .Y(new_n16917));
  not_8  g14569(.A(new_n16917), .Y(new_n16918));
  xor_4  g14570(.A(new_n16911_1), .B(new_n12392), .Y(new_n16919));
  or_5   g14571(.A(new_n16919), .B(n19941), .Y(new_n16920));
  nand_5 g14572(.A(new_n16919), .B(n19941), .Y(new_n16921));
  xor_4  g14573(.A(new_n16910), .B(n5077), .Y(new_n16922));
  or_5   g14574(.A(new_n16922), .B(n1099), .Y(new_n16923));
  nand_5 g14575(.A(new_n16922), .B(n1099), .Y(new_n16924));
  nand_5 g14576(.A(new_n16909), .B(n15546), .Y(new_n16925));
  and_5  g14577(.A(new_n16925), .B(new_n16910), .Y(new_n16926));
  or_5   g14578(.A(new_n16926), .B(n2113), .Y(new_n16927));
  nand_5 g14579(.A(new_n16926), .B(n2113), .Y(new_n16928));
  nand_5 g14580(.A(new_n4770_1), .B(n26452), .Y(new_n16929));
  and_5  g14581(.A(new_n16929), .B(new_n16909), .Y(new_n16930));
  or_5   g14582(.A(new_n16930), .B(n21134), .Y(new_n16931));
  nand_5 g14583(.A(new_n16930), .B(n21134), .Y(new_n16932));
  nand_5 g14584(.A(new_n4775), .B(new_n4766_1), .Y(new_n16933));
  nand_5 g14585(.A(new_n16933), .B(new_n4773), .Y(new_n16934));
  nand_5 g14586(.A(new_n16934), .B(new_n16932), .Y(new_n16935));
  nand_5 g14587(.A(new_n16935), .B(new_n16931), .Y(new_n16936));
  nand_5 g14588(.A(new_n16936), .B(new_n16928), .Y(new_n16937));
  nand_5 g14589(.A(new_n16937), .B(new_n16927), .Y(new_n16938));
  nand_5 g14590(.A(new_n16938), .B(new_n16924), .Y(new_n16939));
  nand_5 g14591(.A(new_n16939), .B(new_n16923), .Y(new_n16940));
  nand_5 g14592(.A(new_n16940), .B(new_n16921), .Y(new_n16941));
  nand_5 g14593(.A(new_n16941), .B(new_n16920), .Y(new_n16942));
  nor_5  g14594(.A(new_n16942), .B(new_n16918), .Y(new_n16943));
  nor_5  g14595(.A(new_n16916), .B(new_n8431), .Y(new_n16944));
  not_8  g14596(.A(new_n16944), .Y(new_n16945));
  nand_5 g14597(.A(new_n16945), .B(new_n16914), .Y(new_n16946));
  nor_5  g14598(.A(new_n16946), .B(new_n16943), .Y(new_n16947));
  nand_5 g14599(.A(new_n16947), .B(new_n16907), .Y(new_n16948));
  not_8  g14600(.A(new_n16947), .Y(new_n16949));
  nand_5 g14601(.A(new_n16949), .B(new_n16906), .Y(new_n16950));
  nand_5 g14602(.A(new_n16950), .B(new_n16948), .Y(new_n16951_1));
  nand_5 g14603(.A(new_n16877), .B(new_n16876), .Y(new_n16952));
  xor_4  g14604(.A(new_n16952), .B(new_n16900), .Y(new_n16953));
  nand_5 g14605(.A(new_n16945), .B(new_n16917), .Y(new_n16954_1));
  xor_4  g14606(.A(new_n16954_1), .B(new_n16942), .Y(new_n16955));
  not_8  g14607(.A(new_n16955), .Y(new_n16956));
  nand_5 g14608(.A(new_n16956), .B(new_n16953), .Y(new_n16957));
  not_8  g14609(.A(new_n16953), .Y(new_n16958));
  nand_5 g14610(.A(new_n16955), .B(new_n16958), .Y(new_n16959));
  nand_5 g14611(.A(new_n16921), .B(new_n16920), .Y(new_n16960));
  xor_4  g14612(.A(new_n16960), .B(new_n16940), .Y(new_n16961));
  not_8  g14613(.A(new_n16961), .Y(new_n16962));
  nand_5 g14614(.A(new_n16882), .B(new_n16880), .Y(new_n16963));
  xor_4  g14615(.A(new_n16963), .B(new_n16898), .Y(new_n16964));
  nand_5 g14616(.A(new_n16964), .B(new_n16962), .Y(new_n16965));
  or_5   g14617(.A(new_n16964), .B(new_n16962), .Y(new_n16966));
  nand_5 g14618(.A(new_n16887), .B(new_n16885_1), .Y(new_n16967));
  xor_4  g14619(.A(new_n16967), .B(new_n16896), .Y(new_n16968_1));
  nand_5 g14620(.A(new_n16924), .B(new_n16923), .Y(new_n16969));
  xor_4  g14621(.A(new_n16969), .B(new_n16938), .Y(new_n16970));
  not_8  g14622(.A(new_n16970), .Y(new_n16971_1));
  nand_5 g14623(.A(new_n16971_1), .B(new_n16968_1), .Y(new_n16972));
  not_8  g14624(.A(new_n16968_1), .Y(new_n16973));
  nand_5 g14625(.A(new_n16970), .B(new_n16973), .Y(new_n16974));
  nand_5 g14626(.A(new_n16928), .B(new_n16927), .Y(new_n16975));
  xor_4  g14627(.A(new_n16975), .B(new_n16936), .Y(new_n16976));
  not_8  g14628(.A(new_n16976), .Y(new_n16977));
  nand_5 g14629(.A(new_n16890), .B(new_n16891), .Y(new_n16978));
  xor_4  g14630(.A(new_n16978), .B(new_n16894), .Y(new_n16979));
  nand_5 g14631(.A(new_n16979), .B(new_n16977), .Y(new_n16980));
  or_5   g14632(.A(new_n16979), .B(new_n16977), .Y(new_n16981));
  nand_5 g14633(.A(new_n16932), .B(new_n16931), .Y(new_n16982));
  xor_4  g14634(.A(new_n16982), .B(new_n16934), .Y(new_n16983));
  or_5   g14635(.A(new_n16983), .B(new_n16827), .Y(new_n16984));
  nand_5 g14636(.A(new_n16983), .B(new_n16827), .Y(new_n16985));
  nand_5 g14637(.A(new_n4809), .B(new_n4764), .Y(new_n16986));
  nand_5 g14638(.A(new_n16986), .B(new_n4807), .Y(new_n16987));
  nand_5 g14639(.A(new_n16987), .B(new_n16985), .Y(new_n16988_1));
  nand_5 g14640(.A(new_n16988_1), .B(new_n16984), .Y(new_n16989_1));
  nand_5 g14641(.A(new_n16989_1), .B(new_n16981), .Y(new_n16990));
  nand_5 g14642(.A(new_n16990), .B(new_n16980), .Y(new_n16991));
  nand_5 g14643(.A(new_n16991), .B(new_n16974), .Y(new_n16992));
  nand_5 g14644(.A(new_n16992), .B(new_n16972), .Y(new_n16993));
  nand_5 g14645(.A(new_n16993), .B(new_n16966), .Y(new_n16994_1));
  nand_5 g14646(.A(new_n16994_1), .B(new_n16965), .Y(new_n16995));
  nand_5 g14647(.A(new_n16995), .B(new_n16959), .Y(new_n16996));
  nand_5 g14648(.A(new_n16996), .B(new_n16957), .Y(new_n16997));
  xor_4  g14649(.A(new_n16997), .B(new_n16951_1), .Y(n2929));
  nand_5 g14650(.A(n12821), .B(new_n11708), .Y(new_n16999));
  nand_5 g14651(.A(new_n2862), .B(n5579), .Y(new_n17000));
  nand_5 g14652(.A(new_n2768), .B(n3468), .Y(new_n17001));
  nand_5 g14653(.A(n23430), .B(new_n3002), .Y(new_n17002));
  nand_5 g14654(.A(new_n15555_1), .B(new_n15552), .Y(new_n17003));
  nand_5 g14655(.A(new_n17003), .B(new_n15554), .Y(new_n17004));
  nand_5 g14656(.A(new_n17004), .B(new_n17002), .Y(new_n17005));
  nand_5 g14657(.A(new_n17005), .B(new_n17001), .Y(new_n17006_1));
  nand_5 g14658(.A(new_n17006_1), .B(new_n17000), .Y(new_n17007));
  nand_5 g14659(.A(new_n17007), .B(new_n16999), .Y(new_n17008));
  nand_5 g14660(.A(new_n2767), .B(n22492), .Y(new_n17009));
  nand_5 g14661(.A(n25523), .B(new_n2798), .Y(new_n17010));
  nand_5 g14662(.A(new_n17010), .B(new_n17009), .Y(new_n17011));
  xor_4  g14663(.A(new_n17011), .B(new_n17008), .Y(new_n17012));
  nand_5 g14664(.A(new_n17012), .B(new_n8376_1), .Y(new_n17013));
  not_8  g14665(.A(new_n17012), .Y(new_n17014));
  nand_5 g14666(.A(new_n17014), .B(new_n8377), .Y(new_n17015));
  nand_5 g14667(.A(new_n17000), .B(new_n16999), .Y(new_n17016));
  xor_4  g14668(.A(new_n17016), .B(new_n17006_1), .Y(new_n17017));
  nand_5 g14669(.A(new_n17017), .B(new_n8381_1), .Y(new_n17018));
  not_8  g14670(.A(new_n17017), .Y(new_n17019));
  nand_5 g14671(.A(new_n17019), .B(new_n8383), .Y(new_n17020));
  nand_5 g14672(.A(new_n17002), .B(new_n17001), .Y(new_n17021));
  xor_4  g14673(.A(new_n17021), .B(new_n17004), .Y(new_n17022));
  nand_5 g14674(.A(new_n17022), .B(new_n8386), .Y(new_n17023));
  not_8  g14675(.A(new_n17022), .Y(new_n17024));
  nand_5 g14676(.A(new_n17024), .B(new_n8388), .Y(new_n17025));
  nand_5 g14677(.A(new_n15858), .B(new_n15855), .Y(new_n17026));
  nand_5 g14678(.A(new_n17026), .B(new_n15857), .Y(new_n17027));
  nand_5 g14679(.A(new_n17027), .B(new_n17025), .Y(new_n17028));
  nand_5 g14680(.A(new_n17028), .B(new_n17023), .Y(new_n17029));
  nand_5 g14681(.A(new_n17029), .B(new_n17020), .Y(new_n17030));
  nand_5 g14682(.A(new_n17030), .B(new_n17018), .Y(new_n17031));
  nand_5 g14683(.A(new_n17031), .B(new_n17015), .Y(new_n17032));
  nand_5 g14684(.A(new_n17032), .B(new_n17013), .Y(new_n17033));
  nand_5 g14685(.A(new_n17010), .B(new_n17008), .Y(new_n17034));
  nand_5 g14686(.A(new_n17034), .B(new_n17009), .Y(new_n17035_1));
  nand_5 g14687(.A(new_n11701), .B(n7330), .Y(new_n17036));
  nand_5 g14688(.A(n8439), .B(new_n2792), .Y(new_n17037_1));
  nand_5 g14689(.A(new_n17037_1), .B(new_n17036), .Y(new_n17038));
  xor_4  g14690(.A(new_n17038), .B(new_n17035_1), .Y(new_n17039));
  nand_5 g14691(.A(new_n17039), .B(new_n8370), .Y(new_n17040));
  not_8  g14692(.A(new_n8370), .Y(new_n17041));
  not_8  g14693(.A(new_n17039), .Y(new_n17042));
  nand_5 g14694(.A(new_n17042), .B(new_n17041), .Y(new_n17043));
  nand_5 g14695(.A(new_n17043), .B(new_n17040), .Y(new_n17044));
  xor_4  g14696(.A(new_n17044), .B(new_n17033), .Y(new_n17045));
  not_8  g14697(.A(new_n17045), .Y(new_n17046));
  nand_5 g14698(.A(new_n11706), .B(n12875), .Y(new_n17047));
  nand_5 g14699(.A(n26318), .B(new_n2997), .Y(new_n17048));
  nand_5 g14700(.A(new_n11710_1), .B(n2035), .Y(new_n17049));
  nand_5 g14701(.A(n26054), .B(new_n3000), .Y(new_n17050));
  nand_5 g14702(.A(new_n11713), .B(n5213), .Y(new_n17051));
  nand_5 g14703(.A(n19081), .B(new_n3004), .Y(new_n17052));
  nand_5 g14704(.A(new_n15865), .B(new_n15863), .Y(new_n17053));
  nand_5 g14705(.A(new_n17053), .B(new_n15864), .Y(new_n17054));
  nand_5 g14706(.A(new_n17054), .B(new_n17052), .Y(new_n17055));
  nand_5 g14707(.A(new_n17055), .B(new_n17051), .Y(new_n17056));
  nand_5 g14708(.A(new_n17056), .B(new_n17050), .Y(new_n17057));
  nand_5 g14709(.A(new_n17057), .B(new_n17049), .Y(new_n17058));
  nand_5 g14710(.A(new_n17058), .B(new_n17048), .Y(new_n17059));
  nand_5 g14711(.A(new_n17059), .B(new_n17047), .Y(new_n17060));
  nand_5 g14712(.A(new_n11703), .B(n1662), .Y(new_n17061));
  nand_5 g14713(.A(n3710), .B(new_n3030_1), .Y(new_n17062));
  nand_5 g14714(.A(new_n17062), .B(new_n17061), .Y(new_n17063));
  xor_4  g14715(.A(new_n17063), .B(new_n17060), .Y(new_n17064));
  or_5   g14716(.A(new_n17064), .B(new_n17046), .Y(new_n17065));
  nand_5 g14717(.A(new_n17064), .B(new_n17046), .Y(new_n17066));
  nand_5 g14718(.A(new_n17013), .B(new_n17015), .Y(new_n17067));
  xor_4  g14719(.A(new_n17067), .B(new_n17031), .Y(new_n17068_1));
  not_8  g14720(.A(new_n17068_1), .Y(new_n17069_1));
  nand_5 g14721(.A(new_n17048), .B(new_n17047), .Y(new_n17070_1));
  xor_4  g14722(.A(new_n17070_1), .B(new_n17058), .Y(new_n17071));
  or_5   g14723(.A(new_n17071), .B(new_n17069_1), .Y(new_n17072));
  nand_5 g14724(.A(new_n17071), .B(new_n17069_1), .Y(new_n17073));
  nand_5 g14725(.A(new_n17018), .B(new_n17020), .Y(new_n17074));
  xor_4  g14726(.A(new_n17074), .B(new_n17029), .Y(new_n17075_1));
  not_8  g14727(.A(new_n17075_1), .Y(new_n17076));
  nand_5 g14728(.A(new_n17050), .B(new_n17049), .Y(new_n17077_1));
  xor_4  g14729(.A(new_n17077_1), .B(new_n17056), .Y(new_n17078));
  or_5   g14730(.A(new_n17078), .B(new_n17076), .Y(new_n17079));
  nand_5 g14731(.A(new_n17078), .B(new_n17076), .Y(new_n17080));
  nand_5 g14732(.A(new_n17023), .B(new_n17025), .Y(new_n17081));
  xor_4  g14733(.A(new_n17081), .B(new_n17027), .Y(new_n17082));
  nand_5 g14734(.A(new_n17052), .B(new_n17051), .Y(new_n17083));
  xor_4  g14735(.A(new_n17083), .B(new_n17054), .Y(new_n17084_1));
  not_8  g14736(.A(new_n17084_1), .Y(new_n17085));
  nand_5 g14737(.A(new_n17085), .B(new_n17082), .Y(new_n17086));
  not_8  g14738(.A(new_n17086), .Y(new_n17087));
  not_8  g14739(.A(new_n17082), .Y(new_n17088));
  nand_5 g14740(.A(new_n17084_1), .B(new_n17088), .Y(new_n17089));
  not_8  g14741(.A(new_n17089), .Y(new_n17090_1));
  not_8  g14742(.A(new_n15853), .Y(new_n17091));
  nor_5  g14743(.A(new_n15870), .B(new_n17091), .Y(new_n17092));
  nor_5  g14744(.A(new_n17092), .B(new_n15869_1), .Y(new_n17093));
  nor_5  g14745(.A(new_n17093), .B(new_n17090_1), .Y(new_n17094));
  nor_5  g14746(.A(new_n17094), .B(new_n17087), .Y(new_n17095_1));
  not_8  g14747(.A(new_n17095_1), .Y(new_n17096));
  nand_5 g14748(.A(new_n17096), .B(new_n17080), .Y(new_n17097));
  nand_5 g14749(.A(new_n17097), .B(new_n17079), .Y(new_n17098));
  nand_5 g14750(.A(new_n17098), .B(new_n17073), .Y(new_n17099));
  nand_5 g14751(.A(new_n17099), .B(new_n17072), .Y(new_n17100));
  nand_5 g14752(.A(new_n17100), .B(new_n17066), .Y(new_n17101));
  nand_5 g14753(.A(new_n17101), .B(new_n17065), .Y(new_n17102));
  nand_5 g14754(.A(new_n17043), .B(new_n17033), .Y(new_n17103));
  nand_5 g14755(.A(new_n17103), .B(new_n17040), .Y(new_n17104_1));
  not_8  g14756(.A(new_n17104_1), .Y(new_n17105));
  nand_5 g14757(.A(new_n17037_1), .B(new_n17035_1), .Y(new_n17106_1));
  nand_5 g14758(.A(new_n17106_1), .B(new_n17036), .Y(new_n17107));
  not_8  g14759(.A(new_n17107), .Y(new_n17108));
  nand_5 g14760(.A(new_n2766), .B(n767), .Y(new_n17109));
  nand_5 g14761(.A(n22793), .B(new_n2785), .Y(new_n17110));
  nand_5 g14762(.A(new_n17110), .B(new_n17109), .Y(new_n17111));
  xor_4  g14763(.A(new_n17111), .B(new_n17108), .Y(new_n17112));
  not_8  g14764(.A(new_n17112), .Y(new_n17113));
  nand_5 g14765(.A(new_n17113), .B(new_n8364), .Y(new_n17114));
  not_8  g14766(.A(new_n8364), .Y(new_n17115));
  nand_5 g14767(.A(new_n17112), .B(new_n17115), .Y(new_n17116));
  nand_5 g14768(.A(new_n17116), .B(new_n17114), .Y(new_n17117));
  xor_4  g14769(.A(new_n17117), .B(new_n17105), .Y(new_n17118));
  not_8  g14770(.A(new_n17118), .Y(new_n17119_1));
  nand_5 g14771(.A(new_n17062), .B(new_n17060), .Y(new_n17120));
  nand_5 g14772(.A(new_n17120), .B(new_n17061), .Y(new_n17121));
  nand_5 g14773(.A(n22379), .B(new_n11699), .Y(new_n17122));
  nand_5 g14774(.A(new_n3276), .B(n15077), .Y(new_n17123));
  nand_5 g14775(.A(new_n17123), .B(new_n17122), .Y(new_n17124));
  xnor_4 g14776(.A(new_n17124), .B(new_n17121), .Y(new_n17125));
  nand_5 g14777(.A(new_n17125), .B(new_n17119_1), .Y(new_n17126));
  not_8  g14778(.A(new_n17126), .Y(new_n17127));
  nor_5  g14779(.A(new_n17125), .B(new_n17119_1), .Y(new_n17128));
  nor_5  g14780(.A(new_n17128), .B(new_n17127), .Y(new_n17129));
  xor_4  g14781(.A(new_n17129), .B(new_n17102), .Y(n2948));
  nand_5 g14782(.A(new_n16402), .B(new_n16400), .Y(new_n17131));
  xnor_4 g14783(.A(new_n17131), .B(new_n16427), .Y(n2961));
  nand_5 g14784(.A(new_n13091), .B(new_n13093), .Y(new_n17133));
  xnor_4 g14785(.A(new_n17133), .B(new_n13114), .Y(n2971));
  nand_5 g14786(.A(new_n2536), .B(new_n2535_1), .Y(new_n17135));
  xnor_4 g14787(.A(new_n17135), .B(new_n2559), .Y(n3010));
  nand_5 g14788(.A(new_n7691), .B(new_n7690), .Y(new_n17137));
  xor_4  g14789(.A(new_n17137), .B(new_n7702), .Y(n3017));
  nor_5  g14790(.A(new_n13507), .B(new_n13504), .Y(new_n17139));
  xor_4  g14791(.A(new_n17139), .B(new_n13501_1), .Y(n3020));
  nor_5  g14792(.A(new_n6948), .B(new_n6947), .Y(new_n17141));
  xor_4  g14793(.A(new_n17141), .B(new_n6977), .Y(n3067));
  nand_5 g14794(.A(n23541), .B(n19234), .Y(new_n17143));
  not_8  g14795(.A(new_n17143), .Y(new_n17144));
  nor_5  g14796(.A(n23541), .B(n19234), .Y(new_n17145));
  or_5   g14797(.A(new_n17145), .B(new_n17144), .Y(new_n17146));
  not_8  g14798(.A(new_n17146), .Y(new_n17147));
  nand_5 g14799(.A(n27134), .B(new_n2611), .Y(new_n17148));
  nand_5 g14800(.A(new_n11378), .B(n4588), .Y(new_n17149));
  and_5  g14801(.A(new_n17149), .B(new_n17148), .Y(new_n17150));
  not_8  g14802(.A(new_n17150), .Y(new_n17151));
  nand_5 g14803(.A(new_n17151), .B(new_n17147), .Y(new_n17152));
  not_8  g14804(.A(new_n17152), .Y(new_n17153));
  nor_5  g14805(.A(new_n17151), .B(new_n17147), .Y(new_n17154));
  nor_5  g14806(.A(new_n17154), .B(new_n17153), .Y(new_n17155));
  nand_5 g14807(.A(new_n17155), .B(new_n11498), .Y(new_n17156));
  not_8  g14808(.A(new_n17156), .Y(new_n17157));
  nor_5  g14809(.A(new_n17155), .B(new_n11498), .Y(new_n17158));
  nor_5  g14810(.A(new_n17158), .B(new_n17157), .Y(n3076));
  nand_5 g14811(.A(new_n7550), .B(new_n7558_1), .Y(new_n17160));
  nand_5 g14812(.A(n15490), .B(n18), .Y(new_n17161));
  and_5  g14813(.A(new_n17161), .B(new_n17160), .Y(new_n17162));
  or_5   g14814(.A(new_n17162), .B(n2809), .Y(new_n17163_1));
  nand_5 g14815(.A(new_n17162), .B(n2809), .Y(new_n17164));
  nand_5 g14816(.A(n15508), .B(n18), .Y(new_n17165));
  nand_5 g14817(.A(new_n17165), .B(new_n17164), .Y(new_n17166));
  nand_5 g14818(.A(new_n17166), .B(new_n17163_1), .Y(new_n17167));
  not_8  g14819(.A(new_n17160), .Y(new_n17168_1));
  nand_5 g14820(.A(new_n17168_1), .B(new_n7569_1), .Y(new_n17169));
  nand_5 g14821(.A(new_n17160), .B(n2783), .Y(new_n17170));
  and_5  g14822(.A(new_n17170), .B(new_n17169), .Y(new_n17171));
  not_8  g14823(.A(new_n17171), .Y(new_n17172));
  nand_5 g14824(.A(new_n17172), .B(new_n5391), .Y(new_n17173));
  nand_5 g14825(.A(new_n17171), .B(n19680), .Y(new_n17174));
  nand_5 g14826(.A(new_n17174), .B(new_n17173), .Y(new_n17175));
  xor_4  g14827(.A(new_n17175), .B(new_n17167), .Y(new_n17176));
  nand_5 g14828(.A(new_n17176), .B(new_n12289), .Y(new_n17177));
  not_8  g14829(.A(new_n17176), .Y(new_n17178));
  nand_5 g14830(.A(new_n17178), .B(new_n12290), .Y(new_n17179));
  nand_5 g14831(.A(new_n17164), .B(new_n17163_1), .Y(new_n17180));
  xnor_4 g14832(.A(new_n17180), .B(new_n17165), .Y(new_n17181));
  or_5   g14833(.A(new_n17181), .B(new_n6552), .Y(new_n17182));
  nand_5 g14834(.A(new_n17181), .B(new_n6552), .Y(new_n17183));
  xor_4  g14835(.A(n15508), .B(n18), .Y(new_n17184));
  nand_5 g14836(.A(new_n17184), .B(new_n6554), .Y(new_n17185));
  not_8  g14837(.A(new_n17185), .Y(new_n17186));
  nand_5 g14838(.A(new_n17186), .B(new_n17183), .Y(new_n17187));
  nand_5 g14839(.A(new_n17187), .B(new_n17182), .Y(new_n17188));
  nand_5 g14840(.A(new_n17188), .B(new_n17179), .Y(new_n17189));
  nand_5 g14841(.A(new_n17189), .B(new_n17177), .Y(new_n17190));
  nand_5 g14842(.A(new_n17174), .B(new_n17167), .Y(new_n17191));
  nand_5 g14843(.A(new_n17191), .B(new_n17173), .Y(new_n17192));
  not_8  g14844(.A(new_n17192), .Y(new_n17193));
  nor_5  g14845(.A(new_n17169), .B(n10611), .Y(new_n17194));
  not_8  g14846(.A(new_n17194), .Y(new_n17195));
  nand_5 g14847(.A(new_n17169), .B(n10611), .Y(new_n17196));
  and_5  g14848(.A(new_n17196), .B(new_n17195), .Y(new_n17197));
  not_8  g14849(.A(new_n17197), .Y(new_n17198));
  nand_5 g14850(.A(new_n17198), .B(new_n5388), .Y(new_n17199));
  nand_5 g14851(.A(new_n17197), .B(n7421), .Y(new_n17200));
  nand_5 g14852(.A(new_n17200), .B(new_n17199), .Y(new_n17201));
  xor_4  g14853(.A(new_n17201), .B(new_n17193), .Y(new_n17202_1));
  not_8  g14854(.A(new_n17202_1), .Y(new_n17203));
  nand_5 g14855(.A(new_n17203), .B(new_n12284), .Y(new_n17204));
  nand_5 g14856(.A(new_n17202_1), .B(new_n12285), .Y(new_n17205));
  nand_5 g14857(.A(new_n17205), .B(new_n17204), .Y(new_n17206));
  xnor_4 g14858(.A(new_n17206), .B(new_n17190), .Y(n3089));
  xor_4  g14859(.A(new_n5840_1), .B(new_n5839), .Y(n3125));
  nand_5 g14860(.A(new_n4813), .B(new_n8335), .Y(new_n17209));
  nand_5 g14861(.A(n21839), .B(n19282), .Y(new_n17210));
  nand_5 g14862(.A(new_n3298), .B(new_n3294), .Y(new_n17211));
  nand_5 g14863(.A(new_n17211), .B(new_n3297), .Y(new_n17212));
  nand_5 g14864(.A(new_n17212), .B(new_n17210), .Y(new_n17213));
  nand_5 g14865(.A(new_n17213), .B(new_n17209), .Y(new_n17214));
  nand_5 g14866(.A(new_n17214), .B(new_n12697), .Y(new_n17215));
  nand_5 g14867(.A(new_n17210), .B(new_n17209), .Y(new_n17216));
  xor_4  g14868(.A(new_n17216), .B(new_n17212), .Y(new_n17217));
  nand_5 g14869(.A(new_n17217), .B(new_n12700), .Y(new_n17218));
  not_8  g14870(.A(new_n17217), .Y(new_n17219_1));
  nand_5 g14871(.A(new_n17219_1), .B(new_n12699), .Y(new_n17220));
  nand_5 g14872(.A(new_n12704), .B(new_n3300), .Y(new_n17221));
  nand_5 g14873(.A(new_n12703), .B(new_n3303), .Y(new_n17222));
  nand_5 g14874(.A(new_n12708), .B(new_n3200), .Y(new_n17223));
  nand_5 g14875(.A(new_n12707_1), .B(new_n3199), .Y(new_n17224));
  nand_5 g14876(.A(new_n12712), .B(new_n3113), .Y(new_n17225));
  nand_5 g14877(.A(new_n12711), .B(new_n3112), .Y(new_n17226));
  nand_5 g14878(.A(new_n15279), .B(new_n15277), .Y(new_n17227));
  nand_5 g14879(.A(new_n17227), .B(new_n15278), .Y(new_n17228));
  nand_5 g14880(.A(new_n17228), .B(new_n17226), .Y(new_n17229));
  nand_5 g14881(.A(new_n17229), .B(new_n17225), .Y(new_n17230));
  nand_5 g14882(.A(new_n17230), .B(new_n17224), .Y(new_n17231));
  nand_5 g14883(.A(new_n17231), .B(new_n17223), .Y(new_n17232_1));
  nand_5 g14884(.A(new_n17232_1), .B(new_n17222), .Y(new_n17233));
  nand_5 g14885(.A(new_n17233), .B(new_n17221), .Y(new_n17234));
  nand_5 g14886(.A(new_n17234), .B(new_n17220), .Y(new_n17235));
  nand_5 g14887(.A(new_n17235), .B(new_n17218), .Y(new_n17236_1));
  nor_5  g14888(.A(new_n17236_1), .B(new_n17215), .Y(new_n17237));
  not_8  g14889(.A(new_n17236_1), .Y(new_n17238));
  not_8  g14890(.A(new_n17214), .Y(new_n17239));
  nand_5 g14891(.A(new_n17239), .B(new_n12698), .Y(new_n17240));
  nor_5  g14892(.A(new_n17240), .B(new_n17238), .Y(new_n17241));
  nor_5  g14893(.A(new_n17241), .B(new_n17237), .Y(new_n17242));
  nand_5 g14894(.A(new_n17242), .B(new_n13162), .Y(new_n17243_1));
  or_5   g14895(.A(new_n17242), .B(new_n13162), .Y(new_n17244));
  nand_5 g14896(.A(new_n17244), .B(new_n17243_1), .Y(new_n17245));
  nand_5 g14897(.A(new_n17240), .B(new_n17215), .Y(new_n17246));
  xor_4  g14898(.A(new_n17246), .B(new_n17238), .Y(new_n17247));
  nand_5 g14899(.A(new_n17247), .B(new_n13165), .Y(new_n17248));
  or_5   g14900(.A(new_n17247), .B(new_n13165), .Y(new_n17249));
  nand_5 g14901(.A(new_n17218), .B(new_n17220), .Y(new_n17250_1));
  xor_4  g14902(.A(new_n17250_1), .B(new_n17234), .Y(new_n17251_1));
  nand_5 g14903(.A(new_n17251_1), .B(new_n13175), .Y(new_n17252));
  or_5   g14904(.A(new_n17251_1), .B(new_n13175), .Y(new_n17253));
  nand_5 g14905(.A(new_n17221), .B(new_n17222), .Y(new_n17254));
  xor_4  g14906(.A(new_n17254), .B(new_n17232_1), .Y(new_n17255));
  nand_5 g14907(.A(new_n17255), .B(new_n13183), .Y(new_n17256));
  or_5   g14908(.A(new_n17255), .B(new_n13183), .Y(new_n17257));
  nand_5 g14909(.A(new_n17223), .B(new_n17224), .Y(new_n17258));
  xor_4  g14910(.A(new_n17258), .B(new_n17230), .Y(new_n17259));
  nand_5 g14911(.A(new_n17259), .B(new_n13189), .Y(new_n17260));
  or_5   g14912(.A(new_n17259), .B(new_n13189), .Y(new_n17261));
  nand_5 g14913(.A(new_n17225), .B(new_n17226), .Y(new_n17262));
  xor_4  g14914(.A(new_n17262), .B(new_n17228), .Y(new_n17263_1));
  nand_5 g14915(.A(new_n17263_1), .B(new_n13196), .Y(new_n17264));
  or_5   g14916(.A(new_n17263_1), .B(new_n13196), .Y(new_n17265));
  nand_5 g14917(.A(new_n15283), .B(new_n15274), .Y(new_n17266));
  nand_5 g14918(.A(new_n17266), .B(new_n15282), .Y(new_n17267));
  nand_5 g14919(.A(new_n17267), .B(new_n17265), .Y(new_n17268));
  nand_5 g14920(.A(new_n17268), .B(new_n17264), .Y(new_n17269));
  nand_5 g14921(.A(new_n17269), .B(new_n17261), .Y(new_n17270));
  nand_5 g14922(.A(new_n17270), .B(new_n17260), .Y(new_n17271));
  nand_5 g14923(.A(new_n17271), .B(new_n17257), .Y(new_n17272));
  nand_5 g14924(.A(new_n17272), .B(new_n17256), .Y(new_n17273));
  nand_5 g14925(.A(new_n17273), .B(new_n17253), .Y(new_n17274));
  nand_5 g14926(.A(new_n17274), .B(new_n17252), .Y(new_n17275));
  nand_5 g14927(.A(new_n17275), .B(new_n17249), .Y(new_n17276));
  nand_5 g14928(.A(new_n17276), .B(new_n17248), .Y(new_n17277));
  xnor_4 g14929(.A(new_n17277), .B(new_n17245), .Y(n3126));
  nand_5 g14930(.A(new_n13808), .B(new_n13807), .Y(new_n17279));
  xor_4  g14931(.A(new_n17279), .B(new_n13847), .Y(n3208));
  nand_5 g14932(.A(new_n16234), .B(new_n16233), .Y(new_n17281));
  xor_4  g14933(.A(new_n17281), .B(new_n16239), .Y(n3219));
  nor_5  g14934(.A(new_n16733_1), .B(new_n16732), .Y(new_n17283));
  xor_4  g14935(.A(new_n17283), .B(new_n16745), .Y(n3235));
  nand_5 g14936(.A(new_n12925), .B(new_n12924), .Y(new_n17285_1));
  xnor_4 g14937(.A(new_n17285_1), .B(new_n12941_1), .Y(n3244));
  nand_5 g14938(.A(new_n2973), .B(new_n2741), .Y(new_n17287));
  or_5   g14939(.A(new_n17287), .B(n8638), .Y(new_n17288));
  nor_5  g14940(.A(new_n17288), .B(n15979), .Y(new_n17289));
  nand_5 g14941(.A(new_n17289), .B(new_n2725), .Y(new_n17290));
  nor_5  g14942(.A(new_n17290), .B(n24768), .Y(new_n17291));
  not_8  g14943(.A(new_n17291), .Y(new_n17292));
  nand_5 g14944(.A(new_n17290), .B(n24768), .Y(new_n17293));
  nand_5 g14945(.A(new_n17293), .B(new_n17292), .Y(new_n17294));
  nand_5 g14946(.A(new_n17294), .B(new_n10048), .Y(new_n17295));
  nor_5  g14947(.A(new_n17294), .B(new_n10048), .Y(new_n17296));
  not_8  g14948(.A(new_n17296), .Y(new_n17297));
  xor_4  g14949(.A(new_n17289), .B(new_n2725), .Y(new_n17298));
  or_5   g14950(.A(new_n17298), .B(n5226), .Y(new_n17299));
  nand_5 g14951(.A(new_n17298), .B(n5226), .Y(new_n17300));
  xor_4  g14952(.A(new_n17288), .B(n15979), .Y(new_n17301));
  or_5   g14953(.A(new_n17301), .B(n17664), .Y(new_n17302_1));
  nand_5 g14954(.A(new_n17301), .B(n17664), .Y(new_n17303));
  nand_5 g14955(.A(new_n17287), .B(n8638), .Y(new_n17304));
  nand_5 g14956(.A(new_n17304), .B(new_n17288), .Y(new_n17305));
  nand_5 g14957(.A(new_n17305), .B(new_n2669), .Y(new_n17306));
  nor_5  g14958(.A(new_n17305), .B(new_n2669), .Y(new_n17307));
  not_8  g14959(.A(new_n17307), .Y(new_n17308));
  nand_5 g14960(.A(n23541), .B(n16247), .Y(new_n17309));
  and_5  g14961(.A(new_n17309), .B(new_n17287), .Y(new_n17310));
  or_5   g14962(.A(new_n17310), .B(n1136), .Y(new_n17311));
  nand_5 g14963(.A(new_n17310), .B(n1136), .Y(new_n17312));
  nand_5 g14964(.A(new_n17312), .B(new_n17143), .Y(new_n17313));
  nand_5 g14965(.A(new_n17313), .B(new_n17311), .Y(new_n17314));
  nand_5 g14966(.A(new_n17314), .B(new_n17308), .Y(new_n17315));
  nand_5 g14967(.A(new_n17315), .B(new_n17306), .Y(new_n17316));
  nand_5 g14968(.A(new_n17316), .B(new_n17303), .Y(new_n17317));
  nand_5 g14969(.A(new_n17317), .B(new_n17302_1), .Y(new_n17318));
  nand_5 g14970(.A(new_n17318), .B(new_n17300), .Y(new_n17319));
  nand_5 g14971(.A(new_n17319), .B(new_n17299), .Y(new_n17320_1));
  nand_5 g14972(.A(new_n17320_1), .B(new_n17297), .Y(new_n17321));
  nand_5 g14973(.A(new_n17321), .B(new_n17295), .Y(new_n17322));
  not_8  g14974(.A(new_n17322), .Y(new_n17323));
  nand_5 g14975(.A(new_n17291), .B(new_n2715), .Y(new_n17324));
  nand_5 g14976(.A(new_n17292), .B(n8687), .Y(new_n17325));
  nand_5 g14977(.A(new_n17325), .B(new_n17324), .Y(new_n17326));
  nand_5 g14978(.A(new_n17326), .B(new_n2658), .Y(new_n17327));
  nor_5  g14979(.A(new_n17326), .B(new_n2658), .Y(new_n17328));
  not_8  g14980(.A(new_n17328), .Y(new_n17329));
  nand_5 g14981(.A(new_n17329), .B(new_n17327), .Y(new_n17330));
  xor_4  g14982(.A(new_n17330), .B(new_n17323), .Y(new_n17331));
  nand_5 g14983(.A(n6427), .B(new_n9122), .Y(new_n17332));
  nand_5 g14984(.A(new_n17332), .B(new_n15549), .Y(new_n17333));
  nand_5 g14985(.A(new_n11418), .B(n1682), .Y(new_n17334));
  nand_5 g14986(.A(new_n17334), .B(new_n17333), .Y(new_n17335));
  nand_5 g14987(.A(n23513), .B(new_n9120), .Y(new_n17336));
  nand_5 g14988(.A(new_n17336), .B(new_n17335), .Y(new_n17337_1));
  nand_5 g14989(.A(new_n11415), .B(n21), .Y(new_n17338));
  nand_5 g14990(.A(new_n17338), .B(new_n17337_1), .Y(new_n17339));
  xor_4  g14991(.A(new_n17339), .B(new_n11470_1), .Y(new_n17340));
  nand_5 g14992(.A(new_n17340), .B(new_n17019), .Y(new_n17341));
  not_8  g14993(.A(new_n17340), .Y(new_n17342));
  nand_5 g14994(.A(new_n17342), .B(new_n17017), .Y(new_n17343));
  xor_4  g14995(.A(new_n17335), .B(new_n11476), .Y(new_n17344_1));
  not_8  g14996(.A(new_n17344_1), .Y(new_n17345));
  nand_5 g14997(.A(new_n17345), .B(new_n17024), .Y(new_n17346));
  nand_5 g14998(.A(new_n17344_1), .B(new_n17022), .Y(new_n17347));
  nand_5 g14999(.A(new_n15561), .B(new_n15545), .Y(new_n17348));
  nand_5 g15000(.A(new_n17348), .B(new_n15558_1), .Y(new_n17349));
  nand_5 g15001(.A(new_n17349), .B(new_n17347), .Y(new_n17350));
  nand_5 g15002(.A(new_n17350), .B(new_n17346), .Y(new_n17351_1));
  nand_5 g15003(.A(new_n17351_1), .B(new_n17343), .Y(new_n17352));
  nand_5 g15004(.A(new_n17352), .B(new_n17341), .Y(new_n17353));
  nand_5 g15005(.A(new_n9116), .B(n3962), .Y(new_n17354));
  nand_5 g15006(.A(new_n17354), .B(new_n17339), .Y(new_n17355));
  nand_5 g15007(.A(n11579), .B(new_n11412), .Y(new_n17356));
  nand_5 g15008(.A(new_n17356), .B(new_n17355), .Y(new_n17357));
  xor_4  g15009(.A(new_n17357), .B(new_n11465), .Y(new_n17358));
  nand_5 g15010(.A(new_n17358), .B(new_n17014), .Y(new_n17359_1));
  not_8  g15011(.A(new_n17358), .Y(new_n17360));
  nand_5 g15012(.A(new_n17360), .B(new_n17012), .Y(new_n17361));
  nand_5 g15013(.A(new_n17361), .B(new_n17359_1), .Y(new_n17362));
  xor_4  g15014(.A(new_n17362), .B(new_n17353), .Y(new_n17363));
  nand_5 g15015(.A(new_n17363), .B(new_n17331), .Y(new_n17364));
  not_8  g15016(.A(new_n17331), .Y(new_n17365));
  not_8  g15017(.A(new_n17363), .Y(new_n17366));
  nand_5 g15018(.A(new_n17366), .B(new_n17365), .Y(new_n17367));
  nand_5 g15019(.A(new_n17297), .B(new_n17295), .Y(new_n17368));
  xor_4  g15020(.A(new_n17368), .B(new_n17320_1), .Y(new_n17369));
  not_8  g15021(.A(new_n17369), .Y(new_n17370));
  nand_5 g15022(.A(new_n17341), .B(new_n17343), .Y(new_n17371));
  xor_4  g15023(.A(new_n17371), .B(new_n17351_1), .Y(new_n17372));
  nand_5 g15024(.A(new_n17372), .B(new_n17370), .Y(new_n17373));
  not_8  g15025(.A(new_n17372), .Y(new_n17374));
  nand_5 g15026(.A(new_n17374), .B(new_n17369), .Y(new_n17375));
  nand_5 g15027(.A(new_n17300), .B(new_n17299), .Y(new_n17376));
  xor_4  g15028(.A(new_n17376), .B(new_n17318), .Y(new_n17377));
  not_8  g15029(.A(new_n17377), .Y(new_n17378));
  nand_5 g15030(.A(new_n17346), .B(new_n17347), .Y(new_n17379));
  xor_4  g15031(.A(new_n17379), .B(new_n17349), .Y(new_n17380));
  nand_5 g15032(.A(new_n17380), .B(new_n17378), .Y(new_n17381));
  not_8  g15033(.A(new_n17380), .Y(new_n17382));
  nand_5 g15034(.A(new_n17382), .B(new_n17377), .Y(new_n17383));
  nand_5 g15035(.A(new_n17303), .B(new_n17302_1), .Y(new_n17384));
  xor_4  g15036(.A(new_n17384), .B(new_n17316), .Y(new_n17385));
  not_8  g15037(.A(new_n17385), .Y(new_n17386));
  nand_5 g15038(.A(new_n17386), .B(new_n15563), .Y(new_n17387_1));
  nand_5 g15039(.A(new_n17385), .B(new_n15574), .Y(new_n17388));
  nand_5 g15040(.A(new_n17308), .B(new_n17306), .Y(new_n17389));
  xor_4  g15041(.A(new_n17389), .B(new_n17314), .Y(new_n17390));
  not_8  g15042(.A(new_n17390), .Y(new_n17391_1));
  nand_5 g15043(.A(new_n17391_1), .B(new_n15512), .Y(new_n17392_1));
  nand_5 g15044(.A(new_n17390), .B(new_n15524), .Y(new_n17393));
  and_5  g15045(.A(new_n17312), .B(new_n17311), .Y(new_n17394));
  xor_4  g15046(.A(new_n17394), .B(new_n17144), .Y(new_n17395));
  not_8  g15047(.A(new_n17395), .Y(new_n17396));
  nand_5 g15048(.A(new_n17396), .B(new_n15539_1), .Y(new_n17397));
  or_5   g15049(.A(new_n17396), .B(new_n15539_1), .Y(new_n17398));
  nand_5 g15050(.A(new_n17147), .B(new_n15529), .Y(new_n17399));
  nand_5 g15051(.A(new_n17399), .B(new_n17398), .Y(new_n17400));
  nand_5 g15052(.A(new_n17400), .B(new_n17397), .Y(new_n17401));
  nand_5 g15053(.A(new_n17401), .B(new_n17393), .Y(new_n17402));
  nand_5 g15054(.A(new_n17402), .B(new_n17392_1), .Y(new_n17403));
  nand_5 g15055(.A(new_n17403), .B(new_n17388), .Y(new_n17404));
  nand_5 g15056(.A(new_n17404), .B(new_n17387_1), .Y(new_n17405));
  nand_5 g15057(.A(new_n17405), .B(new_n17383), .Y(new_n17406));
  nand_5 g15058(.A(new_n17406), .B(new_n17381), .Y(new_n17407));
  nand_5 g15059(.A(new_n17407), .B(new_n17375), .Y(new_n17408));
  nand_5 g15060(.A(new_n17408), .B(new_n17373), .Y(new_n17409));
  nand_5 g15061(.A(new_n17409), .B(new_n17367), .Y(new_n17410));
  nand_5 g15062(.A(new_n17410), .B(new_n17364), .Y(new_n17411));
  nand_5 g15063(.A(new_n17329), .B(new_n17322), .Y(new_n17412));
  nand_5 g15064(.A(new_n17412), .B(new_n17327), .Y(new_n17413));
  not_8  g15065(.A(new_n17413), .Y(new_n17414));
  not_8  g15066(.A(new_n17324), .Y(new_n17415));
  nand_5 g15067(.A(new_n17415), .B(new_n2709), .Y(new_n17416));
  nand_5 g15068(.A(new_n17324), .B(n19270), .Y(new_n17417));
  nand_5 g15069(.A(new_n17417), .B(new_n17416), .Y(new_n17418));
  nand_5 g15070(.A(new_n17418), .B(new_n10043), .Y(new_n17419));
  nor_5  g15071(.A(new_n17418), .B(new_n10043), .Y(new_n17420));
  not_8  g15072(.A(new_n17420), .Y(new_n17421_1));
  nand_5 g15073(.A(new_n17421_1), .B(new_n17419), .Y(new_n17422));
  xor_4  g15074(.A(new_n17422), .B(new_n17414), .Y(new_n17423));
  nand_5 g15075(.A(new_n17361), .B(new_n17353), .Y(new_n17424));
  nand_5 g15076(.A(new_n17424), .B(new_n17359_1), .Y(new_n17425));
  not_8  g15077(.A(new_n17425), .Y(new_n17426));
  nand_5 g15078(.A(new_n9113), .B(n5532), .Y(new_n17427));
  nand_5 g15079(.A(new_n17427), .B(new_n17357), .Y(new_n17428));
  nand_5 g15080(.A(n15146), .B(new_n11409), .Y(new_n17429));
  nand_5 g15081(.A(new_n17429), .B(new_n17428), .Y(new_n17430));
  not_8  g15082(.A(new_n17430), .Y(new_n17431));
  xor_4  g15083(.A(new_n17431), .B(new_n11461), .Y(new_n17432_1));
  nand_5 g15084(.A(new_n17432_1), .B(new_n17042), .Y(new_n17433));
  not_8  g15085(.A(new_n17432_1), .Y(new_n17434));
  nand_5 g15086(.A(new_n17434), .B(new_n17039), .Y(new_n17435));
  nand_5 g15087(.A(new_n17435), .B(new_n17433), .Y(new_n17436_1));
  xor_4  g15088(.A(new_n17436_1), .B(new_n17426), .Y(new_n17437));
  not_8  g15089(.A(new_n17437), .Y(new_n17438));
  nand_5 g15090(.A(new_n17438), .B(new_n17423), .Y(new_n17439));
  not_8  g15091(.A(new_n17423), .Y(new_n17440_1));
  nand_5 g15092(.A(new_n17437), .B(new_n17440_1), .Y(new_n17441));
  nand_5 g15093(.A(new_n17441), .B(new_n17439), .Y(new_n17442));
  xor_4  g15094(.A(new_n17442), .B(new_n17411), .Y(n3263));
  nand_5 g15095(.A(new_n14063), .B(new_n14064), .Y(new_n17444));
  xnor_4 g15096(.A(new_n17444), .B(new_n14078), .Y(n3289));
  nand_5 g15097(.A(new_n5719), .B(new_n5708), .Y(new_n17446));
  nand_5 g15098(.A(new_n17446), .B(new_n5718), .Y(new_n17447));
  nand_5 g15099(.A(new_n5714), .B(new_n5711), .Y(new_n17448));
  nand_5 g15100(.A(new_n17448), .B(new_n5713), .Y(new_n17449));
  nand_5 g15101(.A(new_n2496), .B(new_n3043), .Y(new_n17450_1));
  nand_5 g15102(.A(n26913), .B(n12956), .Y(new_n17451));
  nand_5 g15103(.A(new_n17451), .B(new_n17450_1), .Y(new_n17452));
  xor_4  g15104(.A(new_n17452), .B(new_n17449), .Y(new_n17453));
  nand_5 g15105(.A(new_n17453), .B(new_n9760), .Y(new_n17454));
  not_8  g15106(.A(new_n17453), .Y(new_n17455));
  nand_5 g15107(.A(new_n17455), .B(n7057), .Y(new_n17456));
  nand_5 g15108(.A(new_n17456), .B(new_n17454), .Y(new_n17457));
  xor_4  g15109(.A(new_n17457), .B(new_n17447), .Y(new_n17458_1));
  nand_5 g15110(.A(new_n10891), .B(new_n5729), .Y(new_n17459));
  nand_5 g15111(.A(new_n10892), .B(n3828), .Y(new_n17460));
  nand_5 g15112(.A(new_n10917), .B(new_n5687_1), .Y(new_n17461_1));
  nand_5 g15113(.A(new_n10859), .B(n23842), .Y(new_n17462));
  nand_5 g15114(.A(new_n10863), .B(n21654), .Y(new_n17463));
  nand_5 g15115(.A(new_n17463), .B(new_n17462), .Y(new_n17464));
  nand_5 g15116(.A(new_n17464), .B(new_n17461_1), .Y(new_n17465));
  nand_5 g15117(.A(new_n17465), .B(new_n17460), .Y(new_n17466_1));
  nand_5 g15118(.A(new_n17466_1), .B(new_n17459), .Y(new_n17467));
  nand_5 g15119(.A(new_n10939), .B(new_n5806), .Y(new_n17468));
  nand_5 g15120(.A(new_n10938), .B(n18274), .Y(new_n17469));
  nand_5 g15121(.A(new_n17469), .B(new_n17468), .Y(new_n17470));
  xor_4  g15122(.A(new_n17470), .B(new_n17467), .Y(new_n17471));
  or_5   g15123(.A(new_n17471), .B(new_n17458_1), .Y(new_n17472));
  nand_5 g15124(.A(new_n17471), .B(new_n17458_1), .Y(new_n17473));
  nand_5 g15125(.A(new_n17459), .B(new_n17460), .Y(new_n17474));
  xor_4  g15126(.A(new_n17474), .B(new_n17465), .Y(new_n17475));
  or_5   g15127(.A(new_n17475), .B(new_n5721), .Y(new_n17476));
  nand_5 g15128(.A(new_n17475), .B(new_n5721), .Y(new_n17477));
  nand_5 g15129(.A(new_n17461_1), .B(new_n17462), .Y(new_n17478));
  xor_4  g15130(.A(new_n17478), .B(new_n17463), .Y(new_n17479));
  or_5   g15131(.A(new_n17479), .B(new_n5676), .Y(new_n17480));
  nand_5 g15132(.A(new_n17479), .B(new_n5676), .Y(new_n17481));
  xor_4  g15133(.A(new_n10863), .B(n21654), .Y(new_n17482));
  nand_5 g15134(.A(new_n17482), .B(new_n5698), .Y(new_n17483));
  nand_5 g15135(.A(new_n17483), .B(new_n17481), .Y(new_n17484));
  nand_5 g15136(.A(new_n17484), .B(new_n17480), .Y(new_n17485));
  nand_5 g15137(.A(new_n17485), .B(new_n17477), .Y(new_n17486));
  nand_5 g15138(.A(new_n17486), .B(new_n17476), .Y(new_n17487));
  nand_5 g15139(.A(new_n17487), .B(new_n17473), .Y(new_n17488));
  nand_5 g15140(.A(new_n17488), .B(new_n17472), .Y(new_n17489));
  nand_5 g15141(.A(new_n17456), .B(new_n17447), .Y(new_n17490));
  nand_5 g15142(.A(new_n17490), .B(new_n17454), .Y(new_n17491));
  nand_5 g15143(.A(new_n17451), .B(new_n17449), .Y(new_n17492));
  nand_5 g15144(.A(new_n17492), .B(new_n17450_1), .Y(new_n17493_1));
  nand_5 g15145(.A(new_n2492), .B(new_n3038), .Y(new_n17494));
  nand_5 g15146(.A(n21832), .B(n5211), .Y(new_n17495));
  nand_5 g15147(.A(new_n17495), .B(new_n17494), .Y(new_n17496));
  xor_4  g15148(.A(new_n17496), .B(new_n17493_1), .Y(new_n17497));
  nand_5 g15149(.A(new_n17497), .B(new_n9757), .Y(new_n17498));
  not_8  g15150(.A(new_n17497), .Y(new_n17499));
  nand_5 g15151(.A(new_n17499), .B(n18537), .Y(new_n17500_1));
  nand_5 g15152(.A(new_n17500_1), .B(new_n17498), .Y(new_n17501));
  xor_4  g15153(.A(new_n17501), .B(new_n17491), .Y(new_n17502));
  nand_5 g15154(.A(new_n17469), .B(new_n17467), .Y(new_n17503));
  nand_5 g15155(.A(new_n17503), .B(new_n17468), .Y(new_n17504));
  nand_5 g15156(.A(new_n16329), .B(new_n5820), .Y(new_n17505));
  nand_5 g15157(.A(new_n16327_1), .B(n21649), .Y(new_n17506));
  nand_5 g15158(.A(new_n17506), .B(new_n17505), .Y(new_n17507));
  xor_4  g15159(.A(new_n17507), .B(new_n17504), .Y(new_n17508));
  or_5   g15160(.A(new_n17508), .B(new_n17502), .Y(new_n17509));
  nand_5 g15161(.A(new_n17508), .B(new_n17502), .Y(new_n17510));
  nand_5 g15162(.A(new_n17510), .B(new_n17509), .Y(new_n17511));
  xor_4  g15163(.A(new_n17511), .B(new_n17489), .Y(n3301));
  nand_5 g15164(.A(new_n12348), .B(n22588), .Y(new_n17513));
  nand_5 g15165(.A(new_n12347), .B(new_n15518), .Y(new_n17514));
  nand_5 g15166(.A(new_n15294), .B(new_n15288), .Y(new_n17515));
  and_5  g15167(.A(new_n17515), .B(new_n15295), .Y(new_n17516));
  nand_5 g15168(.A(new_n17516), .B(new_n17514), .Y(new_n17517));
  nand_5 g15169(.A(new_n17517), .B(new_n17513), .Y(new_n17518));
  nand_5 g15170(.A(new_n12437), .B(n19515), .Y(new_n17519));
  nand_5 g15171(.A(new_n12357), .B(new_n15567), .Y(new_n17520));
  nand_5 g15172(.A(new_n17520), .B(new_n17519), .Y(new_n17521));
  xor_4  g15173(.A(new_n17521), .B(new_n17518), .Y(new_n17522));
  not_8  g15174(.A(new_n17522), .Y(new_n17523));
  nand_5 g15175(.A(new_n17523), .B(new_n11578), .Y(new_n17524_1));
  nand_5 g15176(.A(new_n17522), .B(new_n11579_1), .Y(new_n17525));
  nand_5 g15177(.A(new_n17513), .B(new_n17514), .Y(new_n17526));
  xor_4  g15178(.A(new_n17526), .B(new_n17516), .Y(new_n17527));
  not_8  g15179(.A(new_n17527), .Y(new_n17528));
  nand_5 g15180(.A(new_n17528), .B(new_n11585), .Y(new_n17529_1));
  nand_5 g15181(.A(new_n17527), .B(new_n11586), .Y(new_n17530));
  nand_5 g15182(.A(new_n15300_1), .B(new_n15292), .Y(new_n17531));
  nand_5 g15183(.A(new_n17531), .B(new_n15299), .Y(new_n17532));
  nand_5 g15184(.A(new_n17532), .B(new_n17530), .Y(new_n17533));
  nand_5 g15185(.A(new_n17533), .B(new_n17529_1), .Y(new_n17534));
  nand_5 g15186(.A(new_n17534), .B(new_n17525), .Y(new_n17535));
  nand_5 g15187(.A(new_n17535), .B(new_n17524_1), .Y(new_n17536));
  nand_5 g15188(.A(new_n17520), .B(new_n17518), .Y(new_n17537));
  nand_5 g15189(.A(new_n17537), .B(new_n17519), .Y(new_n17538));
  nand_5 g15190(.A(new_n12364_1), .B(n3030), .Y(new_n17539));
  not_8  g15191(.A(n3030), .Y(new_n17540));
  not_8  g15192(.A(new_n12364_1), .Y(new_n17541));
  nand_5 g15193(.A(new_n17541), .B(new_n17540), .Y(new_n17542));
  nand_5 g15194(.A(new_n17542), .B(new_n17539), .Y(new_n17543));
  xor_4  g15195(.A(new_n17543), .B(new_n17538), .Y(new_n17544));
  or_5   g15196(.A(new_n17544), .B(new_n11572), .Y(new_n17545));
  nand_5 g15197(.A(new_n17544), .B(new_n11572), .Y(new_n17546));
  nand_5 g15198(.A(new_n17546), .B(new_n17545), .Y(new_n17547));
  xor_4  g15199(.A(new_n17547), .B(new_n17536), .Y(n3316));
  nand_5 g15200(.A(new_n15254), .B(new_n15255_1), .Y(new_n17549));
  xor_4  g15201(.A(new_n17549), .B(new_n15270), .Y(n3332));
  nand_5 g15202(.A(new_n14741), .B(new_n14738), .Y(new_n17551));
  nand_5 g15203(.A(new_n17551), .B(new_n14740), .Y(new_n17552));
  not_8  g15204(.A(new_n17552), .Y(new_n17553));
  nand_5 g15205(.A(new_n14746_1), .B(new_n14736), .Y(new_n17554));
  nand_5 g15206(.A(new_n17554), .B(new_n14745), .Y(new_n17555));
  nand_5 g15207(.A(new_n17555), .B(new_n17553), .Y(new_n17556));
  not_8  g15208(.A(new_n17556), .Y(new_n17557_1));
  nand_5 g15209(.A(new_n9153), .B(n17458), .Y(new_n17558));
  nand_5 g15210(.A(new_n9155), .B(new_n8291), .Y(new_n17559));
  nand_5 g15211(.A(new_n9159), .B(n1222), .Y(new_n17560));
  nand_5 g15212(.A(new_n9161), .B(new_n8294), .Y(new_n17561));
  nand_5 g15213(.A(new_n12193), .B(new_n12191), .Y(new_n17562));
  nand_5 g15214(.A(new_n17562), .B(new_n12192_1), .Y(new_n17563));
  nand_5 g15215(.A(new_n17563), .B(new_n17561), .Y(new_n17564));
  nand_5 g15216(.A(new_n17564), .B(new_n17560), .Y(new_n17565));
  nand_5 g15217(.A(new_n17565), .B(new_n17559), .Y(new_n17566));
  nand_5 g15218(.A(new_n17566), .B(new_n17558), .Y(new_n17567));
  nand_5 g15219(.A(new_n17567), .B(new_n9150), .Y(new_n17568));
  nand_5 g15220(.A(new_n17568), .B(new_n17557_1), .Y(new_n17569));
  or_5   g15221(.A(new_n17568), .B(new_n17557_1), .Y(new_n17570));
  nand_5 g15222(.A(new_n17570), .B(new_n17569), .Y(new_n17571));
  nor_5  g15223(.A(new_n17555), .B(new_n17553), .Y(new_n17572));
  nor_5  g15224(.A(new_n17572), .B(new_n17557_1), .Y(new_n17573));
  xor_4  g15225(.A(new_n17567), .B(new_n9149), .Y(new_n17574));
  nand_5 g15226(.A(new_n17574), .B(new_n17573), .Y(new_n17575));
  or_5   g15227(.A(new_n17574), .B(new_n17573), .Y(new_n17576));
  nand_5 g15228(.A(new_n17558), .B(new_n17559), .Y(new_n17577));
  xor_4  g15229(.A(new_n17577), .B(new_n17565), .Y(new_n17578));
  nand_5 g15230(.A(new_n17578), .B(new_n14751), .Y(new_n17579));
  or_5   g15231(.A(new_n17578), .B(new_n14751), .Y(new_n17580));
  nand_5 g15232(.A(new_n17560), .B(new_n17561), .Y(new_n17581));
  xor_4  g15233(.A(new_n17581), .B(new_n17563), .Y(new_n17582));
  nand_5 g15234(.A(new_n17582), .B(new_n14757), .Y(new_n17583_1));
  or_5   g15235(.A(new_n17582), .B(new_n14757), .Y(new_n17584));
  nand_5 g15236(.A(new_n12212), .B(new_n12189), .Y(new_n17585));
  nand_5 g15237(.A(new_n17585), .B(new_n12211), .Y(new_n17586));
  nand_5 g15238(.A(new_n17586), .B(new_n17584), .Y(new_n17587));
  nand_5 g15239(.A(new_n17587), .B(new_n17583_1), .Y(new_n17588));
  nand_5 g15240(.A(new_n17588), .B(new_n17580), .Y(new_n17589));
  nand_5 g15241(.A(new_n17589), .B(new_n17579), .Y(new_n17590));
  nand_5 g15242(.A(new_n17590), .B(new_n17576), .Y(new_n17591));
  nand_5 g15243(.A(new_n17591), .B(new_n17575), .Y(new_n17592_1));
  xor_4  g15244(.A(new_n17592_1), .B(new_n17571), .Y(n3340));
  not_8  g15245(.A(n5098), .Y(new_n17594));
  nand_5 g15246(.A(n26452), .B(new_n17594), .Y(new_n17595));
  nand_5 g15247(.A(new_n12136), .B(n5098), .Y(new_n17596));
  nand_5 g15248(.A(n19905), .B(new_n17540), .Y(new_n17597));
  nand_5 g15249(.A(new_n4768), .B(n3030), .Y(new_n17598));
  nand_5 g15250(.A(new_n15569), .B(new_n15565), .Y(new_n17599));
  nand_5 g15251(.A(new_n17599), .B(new_n15568), .Y(new_n17600));
  nand_5 g15252(.A(new_n17600), .B(new_n17598), .Y(new_n17601));
  nand_5 g15253(.A(new_n17601), .B(new_n17597), .Y(new_n17602));
  nand_5 g15254(.A(new_n17602), .B(new_n17596), .Y(new_n17603));
  nand_5 g15255(.A(new_n17603), .B(new_n17595), .Y(new_n17604));
  not_8  g15256(.A(n24937), .Y(new_n17605));
  nand_5 g15257(.A(new_n17605), .B(n15546), .Y(new_n17606));
  nand_5 g15258(.A(n24937), .B(new_n12158_1), .Y(new_n17607));
  nand_5 g15259(.A(new_n17607), .B(new_n17606), .Y(new_n17608));
  xor_4  g15260(.A(new_n17608), .B(new_n17604), .Y(new_n17609));
  nand_5 g15261(.A(new_n17609), .B(new_n17363), .Y(new_n17610));
  not_8  g15262(.A(new_n17609), .Y(new_n17611));
  nand_5 g15263(.A(new_n17611), .B(new_n17366), .Y(new_n17612));
  nand_5 g15264(.A(new_n17596), .B(new_n17595), .Y(new_n17613));
  xor_4  g15265(.A(new_n17613), .B(new_n17602), .Y(new_n17614));
  nand_5 g15266(.A(new_n17614), .B(new_n17372), .Y(new_n17615));
  not_8  g15267(.A(new_n17614), .Y(new_n17616));
  nand_5 g15268(.A(new_n17616), .B(new_n17374), .Y(new_n17617));
  nand_5 g15269(.A(new_n17598), .B(new_n17597), .Y(new_n17618));
  xor_4  g15270(.A(new_n17618), .B(new_n17600), .Y(new_n17619));
  nand_5 g15271(.A(new_n17619), .B(new_n17380), .Y(new_n17620));
  not_8  g15272(.A(new_n17619), .Y(new_n17621));
  nand_5 g15273(.A(new_n17621), .B(new_n17382), .Y(new_n17622));
  nand_5 g15274(.A(new_n15575), .B(new_n15543), .Y(new_n17623));
  nand_5 g15275(.A(new_n17623), .B(new_n15573_1), .Y(new_n17624));
  nand_5 g15276(.A(new_n17624), .B(new_n17622), .Y(new_n17625));
  nand_5 g15277(.A(new_n17625), .B(new_n17620), .Y(new_n17626));
  nand_5 g15278(.A(new_n17626), .B(new_n17617), .Y(new_n17627));
  nand_5 g15279(.A(new_n17627), .B(new_n17615), .Y(new_n17628));
  nand_5 g15280(.A(new_n17628), .B(new_n17612), .Y(new_n17629));
  nand_5 g15281(.A(new_n17629), .B(new_n17610), .Y(new_n17630));
  nand_5 g15282(.A(new_n17607), .B(new_n17604), .Y(new_n17631));
  nand_5 g15283(.A(new_n17631), .B(new_n17606), .Y(new_n17632));
  not_8  g15284(.A(new_n17632), .Y(new_n17633));
  not_8  g15285(.A(n13851), .Y(new_n17634));
  nand_5 g15286(.A(new_n17634), .B(n5077), .Y(new_n17635));
  nand_5 g15287(.A(n13851), .B(new_n12207), .Y(new_n17636));
  nand_5 g15288(.A(new_n17636), .B(new_n17635), .Y(new_n17637));
  xor_4  g15289(.A(new_n17637), .B(new_n17633), .Y(new_n17638_1));
  not_8  g15290(.A(new_n17638_1), .Y(new_n17639));
  nand_5 g15291(.A(new_n17639), .B(new_n17438), .Y(new_n17640));
  nand_5 g15292(.A(new_n17638_1), .B(new_n17437), .Y(new_n17641));
  nand_5 g15293(.A(new_n17641), .B(new_n17640), .Y(new_n17642));
  xor_4  g15294(.A(new_n17642), .B(new_n17630), .Y(n3343));
  or_5   g15295(.A(new_n17416), .B(n14704), .Y(new_n17644));
  nor_5  g15296(.A(new_n17644), .B(n25365), .Y(new_n17645));
  not_8  g15297(.A(new_n17645), .Y(new_n17646));
  nand_5 g15298(.A(new_n17644), .B(n25365), .Y(new_n17647));
  nand_5 g15299(.A(new_n17647), .B(new_n17646), .Y(new_n17648));
  nand_5 g15300(.A(new_n17648), .B(new_n2648), .Y(new_n17649));
  not_8  g15301(.A(new_n17649), .Y(new_n17650));
  nand_5 g15302(.A(new_n17416), .B(n14704), .Y(new_n17651));
  nand_5 g15303(.A(new_n17651), .B(new_n17644), .Y(new_n17652));
  nand_5 g15304(.A(new_n17652), .B(new_n2652), .Y(new_n17653));
  nor_5  g15305(.A(new_n17652), .B(new_n2652), .Y(new_n17654));
  not_8  g15306(.A(new_n17654), .Y(new_n17655));
  nand_5 g15307(.A(new_n17421_1), .B(new_n17413), .Y(new_n17656));
  nand_5 g15308(.A(new_n17656), .B(new_n17419), .Y(new_n17657));
  nand_5 g15309(.A(new_n17657), .B(new_n17655), .Y(new_n17658));
  nand_5 g15310(.A(new_n17658), .B(new_n17653), .Y(new_n17659));
  nor_5  g15311(.A(new_n17659), .B(new_n17650), .Y(new_n17660));
  nor_5  g15312(.A(new_n17648), .B(new_n2648), .Y(new_n17661));
  not_8  g15313(.A(new_n17661), .Y(new_n17662));
  nand_5 g15314(.A(new_n17662), .B(new_n17646), .Y(new_n17663));
  nor_5  g15315(.A(new_n17663), .B(new_n17660), .Y(new_n17664_1));
  nand_5 g15316(.A(new_n17662), .B(new_n17649), .Y(new_n17665));
  xor_4  g15317(.A(new_n17665), .B(new_n17659), .Y(new_n17666));
  not_8  g15318(.A(new_n17666), .Y(new_n17667));
  nand_5 g15319(.A(new_n17667), .B(new_n15881), .Y(new_n17668));
  nand_5 g15320(.A(new_n17655), .B(new_n17653), .Y(new_n17669));
  xor_4  g15321(.A(new_n17669), .B(new_n17657), .Y(new_n17670));
  not_8  g15322(.A(new_n17670), .Y(new_n17671));
  nand_5 g15323(.A(new_n17671), .B(new_n15884_1), .Y(new_n17672));
  nand_5 g15324(.A(new_n17670), .B(new_n15886), .Y(new_n17673));
  nand_5 g15325(.A(new_n17423), .B(new_n15888), .Y(new_n17674));
  nand_5 g15326(.A(new_n17440_1), .B(new_n15890), .Y(new_n17675));
  nand_5 g15327(.A(new_n17331), .B(new_n7496), .Y(new_n17676));
  nand_5 g15328(.A(new_n17365), .B(new_n7495), .Y(new_n17677));
  nand_5 g15329(.A(new_n17370), .B(new_n7421_1), .Y(new_n17678));
  nand_5 g15330(.A(new_n17369), .B(new_n7420), .Y(new_n17679));
  nand_5 g15331(.A(new_n17378), .B(new_n7365), .Y(new_n17680));
  nand_5 g15332(.A(new_n17377), .B(new_n7364), .Y(new_n17681));
  nand_5 g15333(.A(new_n17386), .B(new_n7338), .Y(new_n17682));
  nand_5 g15334(.A(new_n17385), .B(new_n7337), .Y(new_n17683));
  nand_5 g15335(.A(new_n17391_1), .B(new_n7344), .Y(new_n17684));
  nand_5 g15336(.A(new_n17390), .B(new_n7343), .Y(new_n17685));
  nand_5 g15337(.A(new_n17396), .B(new_n7350), .Y(new_n17686));
  nand_5 g15338(.A(new_n17395), .B(new_n7349_1), .Y(new_n17687_1));
  nand_5 g15339(.A(new_n17147), .B(n4939), .Y(new_n17688));
  nand_5 g15340(.A(new_n17688), .B(new_n17687_1), .Y(new_n17689));
  nand_5 g15341(.A(new_n17689), .B(new_n17686), .Y(new_n17690));
  nand_5 g15342(.A(new_n17690), .B(new_n17685), .Y(new_n17691));
  nand_5 g15343(.A(new_n17691), .B(new_n17684), .Y(new_n17692));
  nand_5 g15344(.A(new_n17692), .B(new_n17683), .Y(new_n17693));
  nand_5 g15345(.A(new_n17693), .B(new_n17682), .Y(new_n17694));
  nand_5 g15346(.A(new_n17694), .B(new_n17681), .Y(new_n17695));
  nand_5 g15347(.A(new_n17695), .B(new_n17680), .Y(new_n17696));
  nand_5 g15348(.A(new_n17696), .B(new_n17679), .Y(new_n17697));
  nand_5 g15349(.A(new_n17697), .B(new_n17678), .Y(new_n17698));
  nand_5 g15350(.A(new_n17698), .B(new_n17677), .Y(new_n17699));
  nand_5 g15351(.A(new_n17699), .B(new_n17676), .Y(new_n17700));
  nand_5 g15352(.A(new_n17700), .B(new_n17675), .Y(new_n17701));
  nand_5 g15353(.A(new_n17701), .B(new_n17674), .Y(new_n17702));
  nand_5 g15354(.A(new_n17702), .B(new_n17673), .Y(new_n17703));
  nand_5 g15355(.A(new_n17703), .B(new_n17672), .Y(new_n17704));
  not_8  g15356(.A(new_n17704), .Y(new_n17705));
  nand_5 g15357(.A(new_n17705), .B(new_n17668), .Y(new_n17706));
  nand_5 g15358(.A(new_n17666), .B(new_n15880), .Y(new_n17707));
  nand_5 g15359(.A(new_n17707), .B(new_n17706), .Y(new_n17708));
  or_5   g15360(.A(new_n17708), .B(new_n15877), .Y(new_n17709));
  xor_4  g15361(.A(new_n17709), .B(new_n17664_1), .Y(new_n17710));
  nand_5 g15362(.A(new_n14244), .B(n10250), .Y(new_n17711));
  or_5   g15363(.A(new_n14244), .B(n10250), .Y(new_n17712));
  nand_5 g15364(.A(new_n14250), .B(n7674), .Y(new_n17713));
  nand_5 g15365(.A(new_n14251), .B(new_n6991), .Y(new_n17714));
  nand_5 g15366(.A(new_n14257), .B(n6397), .Y(new_n17715));
  nand_5 g15367(.A(new_n14258), .B(new_n6997), .Y(new_n17716));
  nand_5 g15368(.A(new_n14264), .B(n19196), .Y(new_n17717));
  nand_5 g15369(.A(new_n14265), .B(new_n7003), .Y(new_n17718));
  nand_5 g15370(.A(new_n14271_1), .B(n23586), .Y(new_n17719));
  nand_5 g15371(.A(new_n14272), .B(new_n7118), .Y(new_n17720));
  nand_5 g15372(.A(new_n14278), .B(n21226), .Y(new_n17721_1));
  or_5   g15373(.A(new_n14278), .B(n21226), .Y(new_n17722));
  nand_5 g15374(.A(new_n14284), .B(n4426), .Y(new_n17723));
  nor_5  g15375(.A(new_n14284), .B(n4426), .Y(new_n17724));
  not_8  g15376(.A(new_n17724), .Y(new_n17725));
  nand_5 g15377(.A(new_n14291), .B(n20036), .Y(new_n17726));
  or_5   g15378(.A(new_n14291), .B(n20036), .Y(new_n17727));
  or_5   g15379(.A(new_n14303), .B(new_n4561), .Y(new_n17728));
  nand_5 g15380(.A(new_n14303), .B(new_n4561), .Y(new_n17729));
  or_5   g15381(.A(new_n14298), .B(n9380), .Y(new_n17730));
  nand_5 g15382(.A(new_n17730), .B(new_n17729), .Y(new_n17731));
  nand_5 g15383(.A(new_n17731), .B(new_n17728), .Y(new_n17732));
  nand_5 g15384(.A(new_n17732), .B(new_n17727), .Y(new_n17733));
  nand_5 g15385(.A(new_n17733), .B(new_n17726), .Y(new_n17734));
  nand_5 g15386(.A(new_n17734), .B(new_n17725), .Y(new_n17735_1));
  nand_5 g15387(.A(new_n17735_1), .B(new_n17723), .Y(new_n17736));
  nand_5 g15388(.A(new_n17736), .B(new_n17722), .Y(new_n17737));
  nand_5 g15389(.A(new_n17737), .B(new_n17721_1), .Y(new_n17738_1));
  nand_5 g15390(.A(new_n17738_1), .B(new_n17720), .Y(new_n17739));
  nand_5 g15391(.A(new_n17739), .B(new_n17719), .Y(new_n17740));
  nand_5 g15392(.A(new_n17740), .B(new_n17718), .Y(new_n17741));
  nand_5 g15393(.A(new_n17741), .B(new_n17717), .Y(new_n17742));
  nand_5 g15394(.A(new_n17742), .B(new_n17716), .Y(new_n17743));
  nand_5 g15395(.A(new_n17743), .B(new_n17715), .Y(new_n17744));
  nand_5 g15396(.A(new_n17744), .B(new_n17714), .Y(new_n17745));
  nand_5 g15397(.A(new_n17745), .B(new_n17713), .Y(new_n17746_1));
  nand_5 g15398(.A(new_n17746_1), .B(new_n17712), .Y(new_n17747));
  nand_5 g15399(.A(new_n17747), .B(new_n17711), .Y(new_n17748));
  xor_4  g15400(.A(new_n17748), .B(new_n14240), .Y(new_n17749_1));
  nand_5 g15401(.A(new_n17749_1), .B(new_n17710), .Y(new_n17750));
  or_5   g15402(.A(new_n17749_1), .B(new_n17710), .Y(new_n17751));
  nand_5 g15403(.A(new_n17712), .B(new_n17711), .Y(new_n17752));
  xor_4  g15404(.A(new_n17752), .B(new_n17746_1), .Y(new_n17753));
  not_8  g15405(.A(new_n17753), .Y(new_n17754));
  nand_5 g15406(.A(new_n17707), .B(new_n17668), .Y(new_n17755));
  xor_4  g15407(.A(new_n17755), .B(new_n17704), .Y(new_n17756));
  or_5   g15408(.A(new_n17756), .B(new_n17754), .Y(new_n17757));
  nand_5 g15409(.A(new_n17756), .B(new_n17754), .Y(new_n17758));
  nand_5 g15410(.A(new_n17714), .B(new_n17713), .Y(new_n17759));
  xor_4  g15411(.A(new_n17759), .B(new_n17744), .Y(new_n17760));
  not_8  g15412(.A(new_n17760), .Y(new_n17761));
  nand_5 g15413(.A(new_n17672), .B(new_n17673), .Y(new_n17762));
  xor_4  g15414(.A(new_n17762), .B(new_n17702), .Y(new_n17763));
  or_5   g15415(.A(new_n17763), .B(new_n17761), .Y(new_n17764));
  nand_5 g15416(.A(new_n17763), .B(new_n17761), .Y(new_n17765));
  nand_5 g15417(.A(new_n17716), .B(new_n17715), .Y(new_n17766));
  xor_4  g15418(.A(new_n17766), .B(new_n17742), .Y(new_n17767));
  not_8  g15419(.A(new_n17767), .Y(new_n17768));
  nand_5 g15420(.A(new_n17674), .B(new_n17675), .Y(new_n17769));
  xor_4  g15421(.A(new_n17769), .B(new_n17700), .Y(new_n17770));
  or_5   g15422(.A(new_n17770), .B(new_n17768), .Y(new_n17771));
  nand_5 g15423(.A(new_n17770), .B(new_n17768), .Y(new_n17772));
  nand_5 g15424(.A(new_n17718), .B(new_n17717), .Y(new_n17773));
  xor_4  g15425(.A(new_n17773), .B(new_n17740), .Y(new_n17774));
  not_8  g15426(.A(new_n17774), .Y(new_n17775));
  nand_5 g15427(.A(new_n17676), .B(new_n17677), .Y(new_n17776));
  xor_4  g15428(.A(new_n17776), .B(new_n17698), .Y(new_n17777));
  or_5   g15429(.A(new_n17777), .B(new_n17775), .Y(new_n17778));
  nand_5 g15430(.A(new_n17777), .B(new_n17775), .Y(new_n17779));
  nand_5 g15431(.A(new_n17720), .B(new_n17719), .Y(new_n17780));
  xor_4  g15432(.A(new_n17780), .B(new_n17738_1), .Y(new_n17781));
  nand_5 g15433(.A(new_n17678), .B(new_n17679), .Y(new_n17782));
  xor_4  g15434(.A(new_n17782), .B(new_n17696), .Y(new_n17783));
  not_8  g15435(.A(new_n17783), .Y(new_n17784_1));
  nand_5 g15436(.A(new_n17784_1), .B(new_n17781), .Y(new_n17785));
  or_5   g15437(.A(new_n17784_1), .B(new_n17781), .Y(new_n17786));
  nand_5 g15438(.A(new_n17722), .B(new_n17721_1), .Y(new_n17787));
  xor_4  g15439(.A(new_n17787), .B(new_n17736), .Y(new_n17788));
  nand_5 g15440(.A(new_n17680), .B(new_n17681), .Y(new_n17789));
  xor_4  g15441(.A(new_n17789), .B(new_n17694), .Y(new_n17790));
  not_8  g15442(.A(new_n17790), .Y(new_n17791));
  nand_5 g15443(.A(new_n17791), .B(new_n17788), .Y(new_n17792));
  or_5   g15444(.A(new_n17791), .B(new_n17788), .Y(new_n17793));
  nand_5 g15445(.A(new_n17725), .B(new_n17723), .Y(new_n17794));
  xor_4  g15446(.A(new_n17794), .B(new_n17734), .Y(new_n17795));
  nand_5 g15447(.A(new_n17682), .B(new_n17683), .Y(new_n17796));
  xor_4  g15448(.A(new_n17796), .B(new_n17692), .Y(new_n17797));
  not_8  g15449(.A(new_n17797), .Y(new_n17798));
  nand_5 g15450(.A(new_n17798), .B(new_n17795), .Y(new_n17799));
  or_5   g15451(.A(new_n17798), .B(new_n17795), .Y(new_n17800));
  nand_5 g15452(.A(new_n17727), .B(new_n17726), .Y(new_n17801));
  xor_4  g15453(.A(new_n17801), .B(new_n17732), .Y(new_n17802));
  nand_5 g15454(.A(new_n17684), .B(new_n17685), .Y(new_n17803));
  xor_4  g15455(.A(new_n17803), .B(new_n17690), .Y(new_n17804));
  not_8  g15456(.A(new_n17804), .Y(new_n17805));
  nand_5 g15457(.A(new_n17805), .B(new_n17802), .Y(new_n17806));
  nor_5  g15458(.A(new_n17805), .B(new_n17802), .Y(new_n17807));
  not_8  g15459(.A(new_n17807), .Y(new_n17808));
  nand_5 g15460(.A(new_n17729), .B(new_n17728), .Y(new_n17809));
  xor_4  g15461(.A(new_n17809), .B(new_n17730), .Y(new_n17810));
  nand_5 g15462(.A(new_n17686), .B(new_n17687_1), .Y(new_n17811));
  xor_4  g15463(.A(new_n17811), .B(new_n17688), .Y(new_n17812));
  not_8  g15464(.A(new_n17812), .Y(new_n17813));
  nand_5 g15465(.A(new_n17813), .B(new_n17810), .Y(new_n17814));
  nor_5  g15466(.A(new_n17813), .B(new_n17810), .Y(new_n17815));
  not_8  g15467(.A(new_n17815), .Y(new_n17816));
  nand_5 g15468(.A(new_n17146), .B(new_n7330_1), .Y(new_n17817));
  and_5  g15469(.A(new_n17817), .B(new_n17688), .Y(new_n17818));
  not_8  g15470(.A(new_n17818), .Y(new_n17819));
  xor_4  g15471(.A(new_n14298), .B(n9380), .Y(new_n17820_1));
  nor_5  g15472(.A(new_n17820_1), .B(new_n17819), .Y(new_n17821));
  not_8  g15473(.A(new_n17821), .Y(new_n17822));
  nand_5 g15474(.A(new_n17822), .B(new_n17816), .Y(new_n17823));
  nand_5 g15475(.A(new_n17823), .B(new_n17814), .Y(new_n17824));
  nand_5 g15476(.A(new_n17824), .B(new_n17808), .Y(new_n17825));
  nand_5 g15477(.A(new_n17825), .B(new_n17806), .Y(new_n17826));
  nand_5 g15478(.A(new_n17826), .B(new_n17800), .Y(new_n17827));
  nand_5 g15479(.A(new_n17827), .B(new_n17799), .Y(new_n17828));
  nand_5 g15480(.A(new_n17828), .B(new_n17793), .Y(new_n17829));
  nand_5 g15481(.A(new_n17829), .B(new_n17792), .Y(new_n17830));
  nand_5 g15482(.A(new_n17830), .B(new_n17786), .Y(new_n17831));
  nand_5 g15483(.A(new_n17831), .B(new_n17785), .Y(new_n17832));
  nand_5 g15484(.A(new_n17832), .B(new_n17779), .Y(new_n17833));
  nand_5 g15485(.A(new_n17833), .B(new_n17778), .Y(new_n17834));
  nand_5 g15486(.A(new_n17834), .B(new_n17772), .Y(new_n17835));
  nand_5 g15487(.A(new_n17835), .B(new_n17771), .Y(new_n17836));
  nand_5 g15488(.A(new_n17836), .B(new_n17765), .Y(new_n17837));
  nand_5 g15489(.A(new_n17837), .B(new_n17764), .Y(new_n17838));
  nand_5 g15490(.A(new_n17838), .B(new_n17758), .Y(new_n17839));
  nand_5 g15491(.A(new_n17839), .B(new_n17757), .Y(new_n17840));
  nand_5 g15492(.A(new_n17840), .B(new_n17751), .Y(new_n17841));
  nand_5 g15493(.A(new_n17841), .B(new_n17750), .Y(new_n17842));
  nor_5  g15494(.A(new_n17709), .B(new_n17664_1), .Y(new_n17843));
  nand_5 g15495(.A(new_n17748), .B(new_n14239), .Y(new_n17844));
  xor_4  g15496(.A(new_n17844), .B(new_n17843), .Y(new_n17845));
  xnor_4 g15497(.A(new_n17845), .B(new_n17842), .Y(n3390));
  nand_5 g15498(.A(new_n7451), .B(new_n7452), .Y(new_n17847));
  xor_4  g15499(.A(new_n17847), .B(new_n7455), .Y(n3426));
  nor_5  g15500(.A(new_n5268), .B(new_n5266), .Y(new_n17849));
  nor_5  g15501(.A(new_n17849), .B(new_n5270), .Y(n3451));
  nor_5  g15502(.A(new_n13942), .B(new_n13940), .Y(new_n17851));
  xor_4  g15503(.A(new_n17851), .B(new_n13963), .Y(n3459));
  nand_5 g15504(.A(n6773), .B(n583), .Y(new_n17853));
  nand_5 g15505(.A(new_n4541), .B(new_n2620), .Y(new_n17854));
  nand_5 g15506(.A(new_n17854), .B(new_n17853), .Y(new_n17855_1));
  nand_5 g15507(.A(new_n17855_1), .B(n21687), .Y(new_n17856));
  not_8  g15508(.A(new_n17856), .Y(new_n17857));
  nor_5  g15509(.A(new_n17855_1), .B(n21687), .Y(new_n17858));
  nor_5  g15510(.A(new_n17858), .B(new_n17857), .Y(new_n17859));
  nor_5  g15511(.A(new_n17859), .B(new_n15655), .Y(new_n17860));
  not_8  g15512(.A(new_n17853), .Y(new_n17861));
  nand_5 g15513(.A(new_n6171_1), .B(new_n4386), .Y(new_n17862));
  nand_5 g15514(.A(n22173), .B(n17090), .Y(new_n17863));
  nand_5 g15515(.A(new_n17863), .B(new_n17862), .Y(new_n17864));
  xor_4  g15516(.A(new_n17864), .B(new_n17861), .Y(new_n17865));
  or_5   g15517(.A(new_n17865), .B(n6729), .Y(new_n17866));
  nand_5 g15518(.A(new_n17865), .B(n6729), .Y(new_n17867));
  nand_5 g15519(.A(new_n17867), .B(new_n17866), .Y(new_n17868));
  xor_4  g15520(.A(new_n17868), .B(new_n17857), .Y(new_n17869));
  nand_5 g15521(.A(new_n17869), .B(new_n15649), .Y(new_n17870));
  or_5   g15522(.A(new_n17869), .B(new_n15649), .Y(new_n17871));
  nand_5 g15523(.A(new_n17871), .B(new_n17870), .Y(new_n17872));
  xnor_4 g15524(.A(new_n17872), .B(new_n17860), .Y(n3502));
  nand_5 g15525(.A(new_n12477), .B(new_n12476), .Y(new_n17874));
  xor_4  g15526(.A(new_n17874), .B(new_n12519), .Y(n3516));
  nand_5 g15527(.A(new_n4547), .B(new_n4559), .Y(new_n17876));
  or_5   g15528(.A(new_n17876), .B(n1689), .Y(new_n17877_1));
  xor_4  g15529(.A(new_n17877_1), .B(n19608), .Y(new_n17878));
  nand_5 g15530(.A(new_n17878), .B(new_n11995), .Y(new_n17879));
  or_5   g15531(.A(new_n17878), .B(new_n11995), .Y(new_n17880));
  xor_4  g15532(.A(new_n17876), .B(n1689), .Y(new_n17881));
  nand_5 g15533(.A(new_n17881), .B(new_n11998), .Y(new_n17882));
  or_5   g15534(.A(new_n17881), .B(new_n11998), .Y(new_n17883));
  nand_5 g15535(.A(n24129), .B(n22274), .Y(new_n17884));
  and_5  g15536(.A(new_n17884), .B(new_n17876), .Y(new_n17885));
  nand_5 g15537(.A(new_n17885), .B(new_n6602), .Y(new_n17886));
  or_5   g15538(.A(new_n17885), .B(new_n6602), .Y(new_n17887));
  nand_5 g15539(.A(new_n4547), .B(n16167), .Y(new_n17888));
  nand_5 g15540(.A(new_n17888), .B(new_n17887), .Y(new_n17889_1));
  nand_5 g15541(.A(new_n17889_1), .B(new_n17886), .Y(new_n17890));
  nand_5 g15542(.A(new_n17890), .B(new_n17883), .Y(new_n17891));
  nand_5 g15543(.A(new_n17891), .B(new_n17882), .Y(new_n17892));
  nand_5 g15544(.A(new_n17892), .B(new_n17880), .Y(new_n17893));
  nand_5 g15545(.A(new_n17893), .B(new_n17879), .Y(new_n17894));
  not_8  g15546(.A(n25126), .Y(new_n17895));
  nor_5  g15547(.A(new_n17877_1), .B(n19608), .Y(new_n17896));
  xor_4  g15548(.A(new_n17896), .B(new_n17895), .Y(new_n17897));
  nand_5 g15549(.A(new_n17897), .B(new_n11992), .Y(new_n17898));
  or_5   g15550(.A(new_n17897), .B(new_n11992), .Y(new_n17899));
  nand_5 g15551(.A(new_n17899), .B(new_n17898), .Y(new_n17900));
  xor_4  g15552(.A(new_n17900), .B(new_n17894), .Y(new_n17901));
  nand_5 g15553(.A(new_n17901), .B(new_n7853), .Y(new_n17902));
  not_8  g15554(.A(new_n17902), .Y(new_n17903));
  not_8  g15555(.A(new_n17901), .Y(new_n17904));
  nand_5 g15556(.A(new_n17904), .B(new_n7851), .Y(new_n17905));
  not_8  g15557(.A(new_n17905), .Y(new_n17906));
  nand_5 g15558(.A(new_n17880), .B(new_n17879), .Y(new_n17907));
  xor_4  g15559(.A(new_n17907), .B(new_n17892), .Y(new_n17908));
  nand_5 g15560(.A(new_n17908), .B(new_n7858), .Y(new_n17909));
  not_8  g15561(.A(new_n17909), .Y(new_n17910));
  not_8  g15562(.A(new_n17908), .Y(new_n17911_1));
  nand_5 g15563(.A(new_n17911_1), .B(new_n7856), .Y(new_n17912_1));
  not_8  g15564(.A(new_n17912_1), .Y(new_n17913));
  nand_5 g15565(.A(new_n17883), .B(new_n17882), .Y(new_n17914));
  xor_4  g15566(.A(new_n17914), .B(new_n17890), .Y(new_n17915));
  or_5   g15567(.A(new_n17915), .B(new_n4600), .Y(new_n17916));
  nand_5 g15568(.A(new_n17915), .B(new_n4600), .Y(new_n17917));
  nand_5 g15569(.A(new_n17887), .B(new_n17886), .Y(new_n17918));
  xnor_4 g15570(.A(new_n17918), .B(new_n17888), .Y(new_n17919));
  nand_5 g15571(.A(new_n17919), .B(new_n4566), .Y(new_n17920));
  nor_5  g15572(.A(new_n17919), .B(new_n4566), .Y(new_n17921));
  not_8  g15573(.A(new_n17921), .Y(new_n17922));
  xor_4  g15574(.A(n24129), .B(new_n6575), .Y(new_n17923));
  nor_5  g15575(.A(new_n17923), .B(new_n4578), .Y(new_n17924));
  nand_5 g15576(.A(new_n17924), .B(new_n17922), .Y(new_n17925));
  nand_5 g15577(.A(new_n17925), .B(new_n17920), .Y(new_n17926));
  nand_5 g15578(.A(new_n17926), .B(new_n17917), .Y(new_n17927_1));
  nand_5 g15579(.A(new_n17927_1), .B(new_n17916), .Y(new_n17928));
  nor_5  g15580(.A(new_n17928), .B(new_n17913), .Y(new_n17929));
  nor_5  g15581(.A(new_n17929), .B(new_n17910), .Y(new_n17930));
  nor_5  g15582(.A(new_n17930), .B(new_n17906), .Y(new_n17931_1));
  nor_5  g15583(.A(new_n17931_1), .B(new_n17903), .Y(new_n17932));
  not_8  g15584(.A(new_n17932), .Y(new_n17933));
  nand_5 g15585(.A(new_n17899), .B(new_n17894), .Y(new_n17934));
  nand_5 g15586(.A(new_n17934), .B(new_n17898), .Y(new_n17935));
  nand_5 g15587(.A(new_n17896), .B(new_n17895), .Y(new_n17936));
  xor_4  g15588(.A(new_n17936), .B(n10712), .Y(new_n17937));
  nand_5 g15589(.A(new_n17937), .B(new_n11989), .Y(new_n17938));
  or_5   g15590(.A(new_n17937), .B(new_n11989), .Y(new_n17939));
  nand_5 g15591(.A(new_n17939), .B(new_n17938), .Y(new_n17940));
  xor_4  g15592(.A(new_n17940), .B(new_n17935), .Y(new_n17941));
  nand_5 g15593(.A(new_n17941), .B(new_n7848), .Y(new_n17942));
  or_5   g15594(.A(new_n17941), .B(new_n7848), .Y(new_n17943));
  nand_5 g15595(.A(new_n17943), .B(new_n17942), .Y(new_n17944));
  xor_4  g15596(.A(new_n17944), .B(new_n17933), .Y(new_n17945));
  nand_5 g15597(.A(new_n17945), .B(new_n11925), .Y(new_n17946));
  or_5   g15598(.A(new_n17945), .B(new_n11925), .Y(new_n17947));
  not_8  g15599(.A(new_n11931), .Y(new_n17948_1));
  nand_5 g15600(.A(new_n17905), .B(new_n17902), .Y(new_n17949));
  xor_4  g15601(.A(new_n17949), .B(new_n17930), .Y(new_n17950));
  or_5   g15602(.A(new_n17950), .B(new_n17948_1), .Y(new_n17951));
  nand_5 g15603(.A(new_n17950), .B(new_n17948_1), .Y(new_n17952));
  nand_5 g15604(.A(new_n17912_1), .B(new_n17909), .Y(new_n17953));
  xor_4  g15605(.A(new_n17953), .B(new_n17928), .Y(new_n17954_1));
  or_5   g15606(.A(new_n17954_1), .B(new_n11938), .Y(new_n17955));
  nand_5 g15607(.A(new_n17954_1), .B(new_n11938), .Y(new_n17956_1));
  nand_5 g15608(.A(new_n17917), .B(new_n17916), .Y(new_n17957));
  xor_4  g15609(.A(new_n17957), .B(new_n17926), .Y(new_n17958));
  and_5  g15610(.A(new_n17958), .B(new_n11944), .Y(new_n17959_1));
  nor_5  g15611(.A(new_n17958), .B(new_n11944), .Y(new_n17960));
  nand_5 g15612(.A(new_n17922), .B(new_n17920), .Y(new_n17961));
  xor_4  g15613(.A(new_n17961), .B(new_n17924), .Y(new_n17962));
  not_8  g15614(.A(new_n17962), .Y(new_n17963_1));
  nand_5 g15615(.A(new_n17963_1), .B(new_n6592), .Y(new_n17964));
  nand_5 g15616(.A(new_n17962), .B(new_n6591), .Y(new_n17965));
  xor_4  g15617(.A(new_n17923), .B(new_n4578), .Y(new_n17966));
  nand_5 g15618(.A(new_n17966), .B(new_n6579), .Y(new_n17967));
  not_8  g15619(.A(new_n17967), .Y(new_n17968_1));
  nand_5 g15620(.A(new_n17968_1), .B(new_n17965), .Y(new_n17969));
  nand_5 g15621(.A(new_n17969), .B(new_n17964), .Y(new_n17970));
  nor_5  g15622(.A(new_n17970), .B(new_n17960), .Y(new_n17971));
  nor_5  g15623(.A(new_n17971), .B(new_n17959_1), .Y(new_n17972));
  nand_5 g15624(.A(new_n17972), .B(new_n17956_1), .Y(new_n17973));
  nand_5 g15625(.A(new_n17973), .B(new_n17955), .Y(new_n17974));
  nand_5 g15626(.A(new_n17974), .B(new_n17952), .Y(new_n17975));
  nand_5 g15627(.A(new_n17975), .B(new_n17951), .Y(new_n17976_1));
  nand_5 g15628(.A(new_n17976_1), .B(new_n17947), .Y(new_n17977));
  nand_5 g15629(.A(new_n17977), .B(new_n17946), .Y(new_n17978));
  not_8  g15630(.A(new_n11920), .Y(new_n17979));
  nand_5 g15631(.A(new_n17943), .B(new_n17933), .Y(new_n17980));
  nand_5 g15632(.A(new_n17980), .B(new_n17942), .Y(new_n17981));
  nand_5 g15633(.A(new_n17939), .B(new_n17935), .Y(new_n17982));
  nand_5 g15634(.A(new_n17982), .B(new_n17938), .Y(new_n17983));
  not_8  g15635(.A(n18145), .Y(new_n17984));
  nor_5  g15636(.A(new_n17936), .B(n10712), .Y(new_n17985));
  xor_4  g15637(.A(new_n17985), .B(new_n17984), .Y(new_n17986));
  nand_5 g15638(.A(new_n17986), .B(new_n11986), .Y(new_n17987));
  or_5   g15639(.A(new_n17986), .B(new_n11986), .Y(new_n17988));
  nand_5 g15640(.A(new_n17988), .B(new_n17987), .Y(new_n17989));
  xor_4  g15641(.A(new_n17989), .B(new_n17983), .Y(new_n17990));
  nand_5 g15642(.A(new_n17990), .B(new_n7841_1), .Y(new_n17991));
  or_5   g15643(.A(new_n17990), .B(new_n7841_1), .Y(new_n17992));
  nand_5 g15644(.A(new_n17992), .B(new_n17991), .Y(new_n17993));
  xnor_4 g15645(.A(new_n17993), .B(new_n17981), .Y(new_n17994));
  or_5   g15646(.A(new_n17994), .B(new_n17979), .Y(new_n17995));
  nand_5 g15647(.A(new_n17994), .B(new_n17979), .Y(new_n17996));
  nand_5 g15648(.A(new_n17996), .B(new_n17995), .Y(new_n17997));
  xnor_4 g15649(.A(new_n17997), .B(new_n17978), .Y(n3528));
  nand_5 g15650(.A(new_n10370), .B(new_n10369), .Y(new_n17999));
  xor_4  g15651(.A(new_n17999), .B(new_n10450), .Y(n3555));
  nor_5  g15652(.A(new_n2778), .B(n13951), .Y(new_n18001));
  nand_5 g15653(.A(new_n11640), .B(new_n18001), .Y(new_n18002));
  nand_5 g15654(.A(new_n2911), .B(new_n2842), .Y(new_n18003));
  not_8  g15655(.A(new_n18003), .Y(new_n18004));
  nor_5  g15656(.A(new_n18004), .B(new_n2844), .Y(new_n18005));
  not_8  g15657(.A(new_n18005), .Y(new_n18006));
  nor_5  g15658(.A(new_n18006), .B(new_n18002), .Y(new_n18007));
  or_5   g15659(.A(new_n11640), .B(new_n18001), .Y(new_n18008));
  nor_5  g15660(.A(new_n18008), .B(new_n18005), .Y(new_n18009));
  nor_5  g15661(.A(new_n18009), .B(new_n18007), .Y(new_n18010));
  or_5   g15662(.A(new_n18010), .B(new_n16643), .Y(new_n18011));
  nand_5 g15663(.A(new_n18008), .B(new_n18002), .Y(new_n18012));
  xor_4  g15664(.A(new_n18012), .B(new_n18005), .Y(new_n18013));
  nand_5 g15665(.A(new_n18013), .B(new_n16688_1), .Y(new_n18014));
  or_5   g15666(.A(new_n18013), .B(new_n16688_1), .Y(new_n18015));
  nand_5 g15667(.A(new_n2994), .B(new_n2914), .Y(new_n18016));
  nand_5 g15668(.A(new_n18016), .B(new_n2913), .Y(new_n18017));
  nand_5 g15669(.A(new_n18017), .B(new_n18015), .Y(new_n18018));
  nand_5 g15670(.A(new_n18018), .B(new_n18014), .Y(new_n18019));
  nand_5 g15671(.A(new_n18019), .B(new_n18011), .Y(new_n18020));
  nand_5 g15672(.A(new_n18010), .B(new_n16643), .Y(new_n18021));
  nand_5 g15673(.A(new_n18021), .B(new_n18020), .Y(new_n18022));
  nor_5  g15674(.A(new_n18022), .B(new_n18007), .Y(n3561));
  nand_5 g15675(.A(new_n12328), .B(new_n12302_1), .Y(new_n18024));
  nand_5 g15676(.A(new_n18024), .B(new_n12326), .Y(new_n18025_1));
  nand_5 g15677(.A(new_n12323), .B(new_n12304_1), .Y(new_n18026));
  nand_5 g15678(.A(new_n18026), .B(new_n12321), .Y(new_n18027));
  not_8  g15679(.A(new_n18027), .Y(new_n18028));
  nand_5 g15680(.A(new_n12310), .B(new_n12307), .Y(new_n18029));
  nand_5 g15681(.A(new_n18029), .B(new_n12309), .Y(new_n18030));
  nand_5 g15682(.A(new_n11164), .B(new_n8565), .Y(new_n18031));
  nand_5 g15683(.A(new_n11163), .B(n1654), .Y(new_n18032));
  nand_5 g15684(.A(new_n18032), .B(new_n18031), .Y(new_n18033));
  xor_4  g15685(.A(new_n18033), .B(new_n18030), .Y(new_n18034));
  not_8  g15686(.A(new_n18034), .Y(new_n18035_1));
  nand_5 g15687(.A(new_n12317), .B(new_n12314), .Y(new_n18036));
  nand_5 g15688(.A(new_n18036), .B(new_n12316), .Y(new_n18037));
  not_8  g15689(.A(new_n18037), .Y(new_n18038));
  nand_5 g15690(.A(new_n4862), .B(n14680), .Y(new_n18039));
  nand_5 g15691(.A(n16439), .B(new_n8804), .Y(new_n18040));
  nand_5 g15692(.A(new_n18040), .B(new_n18039), .Y(new_n18041));
  xor_4  g15693(.A(new_n18041), .B(new_n18038), .Y(new_n18042));
  not_8  g15694(.A(new_n18042), .Y(new_n18043_1));
  nand_5 g15695(.A(new_n18043_1), .B(new_n18035_1), .Y(new_n18044));
  nand_5 g15696(.A(new_n18042), .B(new_n18034), .Y(new_n18045_1));
  nand_5 g15697(.A(new_n18045_1), .B(new_n18044), .Y(new_n18046));
  xor_4  g15698(.A(new_n18046), .B(new_n18028), .Y(new_n18047));
  nand_5 g15699(.A(new_n18047), .B(new_n6291), .Y(new_n18048));
  not_8  g15700(.A(new_n18047), .Y(new_n18049));
  nand_5 g15701(.A(new_n18049), .B(new_n6292), .Y(new_n18050));
  nand_5 g15702(.A(new_n18050), .B(new_n18048), .Y(new_n18051));
  xor_4  g15703(.A(new_n18051), .B(new_n18025_1), .Y(n3563));
  nand_5 g15704(.A(new_n6968), .B(new_n6967_1), .Y(new_n18053));
  xnor_4 g15705(.A(new_n18053), .B(new_n6970), .Y(n3617));
  nand_5 g15706(.A(n22253), .B(new_n7990), .Y(new_n18055));
  nand_5 g15707(.A(new_n8015), .B(n8305), .Y(new_n18056));
  nand_5 g15708(.A(new_n18056), .B(new_n18055), .Y(new_n18057));
  nand_5 g15709(.A(new_n7994), .B(n1255), .Y(new_n18058));
  nand_5 g15710(.A(n12861), .B(new_n8020), .Y(new_n18059_1));
  nand_5 g15711(.A(new_n7997), .B(n9512), .Y(new_n18060));
  nand_5 g15712(.A(n13333), .B(new_n8024), .Y(new_n18061_1));
  nand_5 g15713(.A(n16608), .B(new_n8001), .Y(new_n18062));
  nand_5 g15714(.A(new_n8027_1), .B(n2210), .Y(new_n18063));
  nand_5 g15715(.A(new_n5318), .B(new_n5314), .Y(new_n18064));
  nand_5 g15716(.A(new_n18064), .B(new_n5316), .Y(new_n18065));
  nand_5 g15717(.A(new_n18065), .B(new_n18063), .Y(new_n18066));
  nand_5 g15718(.A(new_n18066), .B(new_n18062), .Y(new_n18067));
  nand_5 g15719(.A(new_n18067), .B(new_n18061_1), .Y(new_n18068));
  nand_5 g15720(.A(new_n18068), .B(new_n18060), .Y(new_n18069));
  nand_5 g15721(.A(new_n18069), .B(new_n18059_1), .Y(new_n18070));
  nand_5 g15722(.A(new_n18070), .B(new_n18058), .Y(new_n18071_1));
  xnor_4 g15723(.A(new_n18071_1), .B(new_n18057), .Y(new_n18072));
  nand_5 g15724(.A(new_n18072), .B(new_n13049), .Y(new_n18073));
  not_8  g15725(.A(new_n18073), .Y(new_n18074));
  nor_5  g15726(.A(new_n18072), .B(new_n13049), .Y(new_n18075));
  nor_5  g15727(.A(new_n18075), .B(new_n18074), .Y(new_n18076));
  nand_5 g15728(.A(new_n18059_1), .B(new_n18058), .Y(new_n18077));
  xor_4  g15729(.A(new_n18077), .B(new_n18069), .Y(new_n18078));
  or_5   g15730(.A(new_n18078), .B(new_n13079), .Y(new_n18079));
  nand_5 g15731(.A(new_n18078), .B(new_n13079), .Y(new_n18080));
  nand_5 g15732(.A(new_n18061_1), .B(new_n18060), .Y(new_n18081));
  xor_4  g15733(.A(new_n18081), .B(new_n18067), .Y(new_n18082));
  or_5   g15734(.A(new_n18082), .B(new_n13087), .Y(new_n18083));
  nand_5 g15735(.A(new_n18082), .B(new_n13087), .Y(new_n18084));
  nand_5 g15736(.A(new_n18063), .B(new_n18062), .Y(new_n18085));
  xor_4  g15737(.A(new_n18085), .B(new_n18065), .Y(new_n18086));
  or_5   g15738(.A(new_n18086), .B(new_n13092), .Y(new_n18087));
  nand_5 g15739(.A(new_n18086), .B(new_n13092), .Y(new_n18088));
  not_8  g15740(.A(new_n5287), .Y(new_n18089));
  nor_5  g15741(.A(new_n5323), .B(new_n18089), .Y(new_n18090));
  nor_5  g15742(.A(new_n18090), .B(new_n5322), .Y(new_n18091));
  not_8  g15743(.A(new_n18091), .Y(new_n18092));
  nand_5 g15744(.A(new_n18092), .B(new_n18088), .Y(new_n18093));
  nand_5 g15745(.A(new_n18093), .B(new_n18087), .Y(new_n18094));
  nand_5 g15746(.A(new_n18094), .B(new_n18084), .Y(new_n18095));
  nand_5 g15747(.A(new_n18095), .B(new_n18083), .Y(new_n18096));
  nand_5 g15748(.A(new_n18096), .B(new_n18080), .Y(new_n18097));
  nand_5 g15749(.A(new_n18097), .B(new_n18079), .Y(new_n18098));
  xor_4  g15750(.A(new_n18098), .B(new_n18076), .Y(n3642));
  nand_5 g15751(.A(n16544), .B(n4319), .Y(new_n18100));
  nand_5 g15752(.A(new_n10316), .B(new_n3313), .Y(new_n18101));
  nand_5 g15753(.A(new_n18101), .B(new_n18100), .Y(new_n18102));
  nand_5 g15754(.A(new_n3318), .B(new_n3286), .Y(new_n18103));
  nand_5 g15755(.A(n23463), .B(n6814), .Y(new_n18104));
  nand_5 g15756(.A(new_n3186), .B(new_n3321), .Y(new_n18105_1));
  nand_5 g15757(.A(n19701), .B(n13074), .Y(new_n18106));
  nand_5 g15758(.A(new_n3068), .B(new_n2601), .Y(new_n18107));
  nand_5 g15759(.A(n23529), .B(n10739), .Y(new_n18108));
  nand_5 g15760(.A(new_n3035), .B(new_n2518), .Y(new_n18109));
  nand_5 g15761(.A(n24620), .B(n21753), .Y(new_n18110));
  nand_5 g15762(.A(new_n17495), .B(new_n17493_1), .Y(new_n18111));
  nand_5 g15763(.A(new_n18111), .B(new_n17494), .Y(new_n18112));
  nand_5 g15764(.A(new_n18112), .B(new_n18110), .Y(new_n18113));
  nand_5 g15765(.A(new_n18113), .B(new_n18109), .Y(new_n18114));
  nand_5 g15766(.A(new_n18114), .B(new_n18108), .Y(new_n18115));
  nand_5 g15767(.A(new_n18115), .B(new_n18107), .Y(new_n18116));
  nand_5 g15768(.A(new_n18116), .B(new_n18106), .Y(new_n18117));
  nand_5 g15769(.A(new_n18117), .B(new_n18105_1), .Y(new_n18118));
  nand_5 g15770(.A(new_n18118), .B(new_n18104), .Y(new_n18119));
  nand_5 g15771(.A(new_n18119), .B(new_n18103), .Y(new_n18120));
  xor_4  g15772(.A(new_n18120), .B(new_n18102), .Y(new_n18121));
  not_8  g15773(.A(new_n18121), .Y(new_n18122));
  nand_5 g15774(.A(new_n18122), .B(n3324), .Y(new_n18123));
  not_8  g15775(.A(n3324), .Y(new_n18124));
  nand_5 g15776(.A(new_n18121), .B(new_n18124), .Y(new_n18125));
  nand_5 g15777(.A(new_n18125), .B(new_n18123), .Y(new_n18126));
  not_8  g15778(.A(n17911), .Y(new_n18127));
  nand_5 g15779(.A(new_n18104), .B(new_n18103), .Y(new_n18128));
  xor_4  g15780(.A(new_n18128), .B(new_n18118), .Y(new_n18129));
  nand_5 g15781(.A(new_n18129), .B(new_n18127), .Y(new_n18130));
  not_8  g15782(.A(new_n18129), .Y(new_n18131));
  nand_5 g15783(.A(new_n18131), .B(n17911), .Y(new_n18132));
  not_8  g15784(.A(n21997), .Y(new_n18133));
  nand_5 g15785(.A(new_n18106), .B(new_n18105_1), .Y(new_n18134));
  xor_4  g15786(.A(new_n18134), .B(new_n18116), .Y(new_n18135));
  nand_5 g15787(.A(new_n18135), .B(new_n18133), .Y(new_n18136));
  not_8  g15788(.A(new_n18135), .Y(new_n18137));
  nand_5 g15789(.A(new_n18137), .B(n21997), .Y(new_n18138));
  nand_5 g15790(.A(new_n18108), .B(new_n18107), .Y(new_n18139));
  xor_4  g15791(.A(new_n18139), .B(new_n18114), .Y(new_n18140));
  nand_5 g15792(.A(new_n18140), .B(new_n9834), .Y(new_n18141));
  not_8  g15793(.A(new_n18140), .Y(new_n18142));
  nand_5 g15794(.A(new_n18142), .B(n25119), .Y(new_n18143_1));
  nand_5 g15795(.A(new_n18110), .B(new_n18109), .Y(new_n18144));
  xor_4  g15796(.A(new_n18144), .B(new_n18112), .Y(new_n18145_1));
  nand_5 g15797(.A(new_n18145_1), .B(new_n9778_1), .Y(new_n18146));
  not_8  g15798(.A(new_n18145_1), .Y(new_n18147));
  nand_5 g15799(.A(new_n18147), .B(n1163), .Y(new_n18148));
  nand_5 g15800(.A(new_n17500_1), .B(new_n17491), .Y(new_n18149));
  nand_5 g15801(.A(new_n18149), .B(new_n17498), .Y(new_n18150));
  nand_5 g15802(.A(new_n18150), .B(new_n18148), .Y(new_n18151_1));
  nand_5 g15803(.A(new_n18151_1), .B(new_n18146), .Y(new_n18152_1));
  nand_5 g15804(.A(new_n18152_1), .B(new_n18143_1), .Y(new_n18153));
  nand_5 g15805(.A(new_n18153), .B(new_n18141), .Y(new_n18154));
  nand_5 g15806(.A(new_n18154), .B(new_n18138), .Y(new_n18155));
  nand_5 g15807(.A(new_n18155), .B(new_n18136), .Y(new_n18156));
  nand_5 g15808(.A(new_n18156), .B(new_n18132), .Y(new_n18157_1));
  nand_5 g15809(.A(new_n18157_1), .B(new_n18130), .Y(new_n18158));
  xor_4  g15810(.A(new_n18158), .B(new_n18126), .Y(new_n18159));
  not_8  g15811(.A(n13419), .Y(new_n18160));
  nand_5 g15812(.A(n6659), .B(new_n3541_1), .Y(new_n18161));
  not_8  g15813(.A(n6659), .Y(new_n18162));
  nand_5 g15814(.A(new_n18162), .B(n5101), .Y(new_n18163));
  nand_5 g15815(.A(new_n18163), .B(new_n18161), .Y(new_n18164));
  nand_5 g15816(.A(n23250), .B(new_n3587), .Y(new_n18165));
  not_8  g15817(.A(n23250), .Y(new_n18166));
  nand_5 g15818(.A(new_n18166), .B(n16507), .Y(new_n18167));
  nand_5 g15819(.A(new_n3613), .B(n11455), .Y(new_n18168));
  not_8  g15820(.A(n11455), .Y(new_n18169));
  nand_5 g15821(.A(n22470), .B(new_n18169), .Y(new_n18170));
  nand_5 g15822(.A(new_n3577), .B(n3945), .Y(new_n18171_1));
  not_8  g15823(.A(n3945), .Y(new_n18172));
  nand_5 g15824(.A(n19116), .B(new_n18172), .Y(new_n18173));
  nand_5 g15825(.A(new_n3546), .B(n5255), .Y(new_n18174));
  nand_5 g15826(.A(n6861), .B(new_n5879), .Y(new_n18175));
  not_8  g15827(.A(n19357), .Y(new_n18176));
  nand_5 g15828(.A(n21649), .B(new_n18176), .Y(new_n18177));
  nand_5 g15829(.A(new_n5820), .B(n19357), .Y(new_n18178));
  nand_5 g15830(.A(n18274), .B(new_n3547), .Y(new_n18179));
  nand_5 g15831(.A(new_n5806), .B(n2328), .Y(new_n18180));
  nand_5 g15832(.A(new_n5730), .B(new_n5726), .Y(new_n18181));
  nand_5 g15833(.A(new_n18181), .B(new_n5728), .Y(new_n18182));
  nand_5 g15834(.A(new_n18182), .B(new_n18180), .Y(new_n18183));
  nand_5 g15835(.A(new_n18183), .B(new_n18179), .Y(new_n18184));
  nand_5 g15836(.A(new_n18184), .B(new_n18178), .Y(new_n18185));
  nand_5 g15837(.A(new_n18185), .B(new_n18177), .Y(new_n18186));
  nand_5 g15838(.A(new_n18186), .B(new_n18175), .Y(new_n18187));
  nand_5 g15839(.A(new_n18187), .B(new_n18174), .Y(new_n18188));
  nand_5 g15840(.A(new_n18188), .B(new_n18173), .Y(new_n18189));
  nand_5 g15841(.A(new_n18189), .B(new_n18171_1), .Y(new_n18190));
  nand_5 g15842(.A(new_n18190), .B(new_n18170), .Y(new_n18191));
  nand_5 g15843(.A(new_n18191), .B(new_n18168), .Y(new_n18192));
  nand_5 g15844(.A(new_n18192), .B(new_n18167), .Y(new_n18193_1));
  nand_5 g15845(.A(new_n18193_1), .B(new_n18165), .Y(new_n18194));
  not_8  g15846(.A(new_n18194), .Y(new_n18195));
  xor_4  g15847(.A(new_n18195), .B(new_n18164), .Y(new_n18196));
  not_8  g15848(.A(new_n18196), .Y(new_n18197));
  nand_5 g15849(.A(new_n18197), .B(new_n18160), .Y(new_n18198));
  nand_5 g15850(.A(new_n18196), .B(n13419), .Y(new_n18199));
  nand_5 g15851(.A(new_n18199), .B(new_n18198), .Y(new_n18200));
  not_8  g15852(.A(n4967), .Y(new_n18201));
  nand_5 g15853(.A(new_n18167), .B(new_n18165), .Y(new_n18202));
  xor_4  g15854(.A(new_n18202), .B(new_n18192), .Y(new_n18203));
  nand_5 g15855(.A(new_n18203), .B(new_n18201), .Y(new_n18204));
  not_8  g15856(.A(new_n18203), .Y(new_n18205));
  nand_5 g15857(.A(new_n18205), .B(n4967), .Y(new_n18206));
  not_8  g15858(.A(n15602), .Y(new_n18207));
  nand_5 g15859(.A(new_n18170), .B(new_n18168), .Y(new_n18208));
  xor_4  g15860(.A(new_n18208), .B(new_n18190), .Y(new_n18209));
  nand_5 g15861(.A(new_n18209), .B(new_n18207), .Y(new_n18210));
  not_8  g15862(.A(new_n18209), .Y(new_n18211));
  nand_5 g15863(.A(new_n18211), .B(n15602), .Y(new_n18212));
  not_8  g15864(.A(n8255), .Y(new_n18213));
  nand_5 g15865(.A(new_n18180), .B(new_n18179), .Y(new_n18214));
  xor_4  g15866(.A(new_n18214), .B(new_n18182), .Y(new_n18215));
  nand_5 g15867(.A(new_n18215), .B(new_n18213), .Y(new_n18216));
  not_8  g15868(.A(new_n18215), .Y(new_n18217));
  nand_5 g15869(.A(new_n18217), .B(n8255), .Y(new_n18218));
  nand_5 g15870(.A(new_n5735), .B(new_n5723), .Y(new_n18219));
  nand_5 g15871(.A(new_n18219), .B(new_n5734), .Y(new_n18220));
  nand_5 g15872(.A(new_n18220), .B(new_n18218), .Y(new_n18221));
  nand_5 g15873(.A(new_n18221), .B(new_n18216), .Y(new_n18222));
  nand_5 g15874(.A(new_n18178), .B(new_n18177), .Y(new_n18223));
  xor_4  g15875(.A(new_n18223), .B(new_n18184), .Y(new_n18224));
  not_8  g15876(.A(new_n18224), .Y(new_n18225));
  nand_5 g15877(.A(new_n18225), .B(n8943), .Y(new_n18226));
  nand_5 g15878(.A(new_n18226), .B(new_n18222), .Y(new_n18227_1));
  not_8  g15879(.A(n8943), .Y(new_n18228));
  nand_5 g15880(.A(new_n18224), .B(new_n18228), .Y(new_n18229));
  nand_5 g15881(.A(new_n18229), .B(new_n18227_1), .Y(new_n18230));
  nand_5 g15882(.A(new_n18175), .B(new_n18174), .Y(new_n18231));
  xor_4  g15883(.A(new_n18231), .B(new_n18186), .Y(new_n18232_1));
  not_8  g15884(.A(new_n18232_1), .Y(new_n18233));
  nand_5 g15885(.A(new_n18233), .B(n12380), .Y(new_n18234));
  nand_5 g15886(.A(new_n18234), .B(new_n18230), .Y(new_n18235));
  not_8  g15887(.A(n12380), .Y(new_n18236));
  nand_5 g15888(.A(new_n18232_1), .B(new_n18236), .Y(new_n18237));
  nand_5 g15889(.A(new_n18237), .B(new_n18235), .Y(new_n18238_1));
  nand_5 g15890(.A(new_n18173), .B(new_n18171_1), .Y(new_n18239));
  xor_4  g15891(.A(new_n18239), .B(new_n18188), .Y(new_n18240));
  not_8  g15892(.A(new_n18240), .Y(new_n18241_1));
  nand_5 g15893(.A(new_n18241_1), .B(n8694), .Y(new_n18242));
  nand_5 g15894(.A(new_n18242), .B(new_n18238_1), .Y(new_n18243));
  not_8  g15895(.A(n8694), .Y(new_n18244));
  nand_5 g15896(.A(new_n18240), .B(new_n18244), .Y(new_n18245));
  nand_5 g15897(.A(new_n18245), .B(new_n18243), .Y(new_n18246));
  nand_5 g15898(.A(new_n18246), .B(new_n18212), .Y(new_n18247));
  nand_5 g15899(.A(new_n18247), .B(new_n18210), .Y(new_n18248));
  nand_5 g15900(.A(new_n18248), .B(new_n18206), .Y(new_n18249));
  nand_5 g15901(.A(new_n18249), .B(new_n18204), .Y(new_n18250));
  xor_4  g15902(.A(new_n18250), .B(new_n18200), .Y(new_n18251));
  nand_5 g15903(.A(new_n18251), .B(new_n18159), .Y(new_n18252));
  or_5   g15904(.A(new_n18251), .B(new_n18159), .Y(new_n18253));
  nand_5 g15905(.A(new_n18253), .B(new_n18252), .Y(new_n18254_1));
  nand_5 g15906(.A(new_n18130), .B(new_n18132), .Y(new_n18255));
  xor_4  g15907(.A(new_n18255), .B(new_n18156), .Y(new_n18256));
  not_8  g15908(.A(new_n18256), .Y(new_n18257));
  nand_5 g15909(.A(new_n18206), .B(new_n18204), .Y(new_n18258));
  xnor_4 g15910(.A(new_n18258), .B(new_n18248), .Y(new_n18259));
  or_5   g15911(.A(new_n18259), .B(new_n18257), .Y(new_n18260));
  nand_5 g15912(.A(new_n18259), .B(new_n18257), .Y(new_n18261));
  nand_5 g15913(.A(new_n18136), .B(new_n18138), .Y(new_n18262));
  xor_4  g15914(.A(new_n18262), .B(new_n18154), .Y(new_n18263));
  not_8  g15915(.A(new_n18263), .Y(new_n18264));
  nand_5 g15916(.A(new_n18212), .B(new_n18210), .Y(new_n18265));
  xnor_4 g15917(.A(new_n18265), .B(new_n18246), .Y(new_n18266));
  or_5   g15918(.A(new_n18266), .B(new_n18264), .Y(new_n18267));
  nand_5 g15919(.A(new_n18266), .B(new_n18264), .Y(new_n18268));
  nand_5 g15920(.A(new_n18141), .B(new_n18143_1), .Y(new_n18269));
  xor_4  g15921(.A(new_n18269), .B(new_n18152_1), .Y(new_n18270));
  not_8  g15922(.A(new_n18270), .Y(new_n18271));
  nand_5 g15923(.A(new_n18241_1), .B(new_n18244), .Y(new_n18272));
  nand_5 g15924(.A(new_n18240), .B(n8694), .Y(new_n18273));
  nand_5 g15925(.A(new_n18273), .B(new_n18272), .Y(new_n18274_1));
  xor_4  g15926(.A(new_n18274_1), .B(new_n18238_1), .Y(new_n18275));
  or_5   g15927(.A(new_n18275), .B(new_n18271), .Y(new_n18276));
  nand_5 g15928(.A(new_n18275), .B(new_n18271), .Y(new_n18277));
  nand_5 g15929(.A(new_n18146), .B(new_n18148), .Y(new_n18278));
  xor_4  g15930(.A(new_n18278), .B(new_n18150), .Y(new_n18279));
  not_8  g15931(.A(new_n18279), .Y(new_n18280));
  nand_5 g15932(.A(new_n18233), .B(new_n18236), .Y(new_n18281));
  nand_5 g15933(.A(new_n18232_1), .B(n12380), .Y(new_n18282));
  nand_5 g15934(.A(new_n18282), .B(new_n18281), .Y(new_n18283));
  xor_4  g15935(.A(new_n18283), .B(new_n18230), .Y(new_n18284));
  or_5   g15936(.A(new_n18284), .B(new_n18280), .Y(new_n18285));
  nand_5 g15937(.A(new_n18284), .B(new_n18280), .Y(new_n18286));
  not_8  g15938(.A(new_n17502), .Y(new_n18287));
  nand_5 g15939(.A(new_n18225), .B(new_n18228), .Y(new_n18288_1));
  nand_5 g15940(.A(new_n18224), .B(n8943), .Y(new_n18289));
  nand_5 g15941(.A(new_n18289), .B(new_n18288_1), .Y(new_n18290_1));
  xor_4  g15942(.A(new_n18290_1), .B(new_n18222), .Y(new_n18291));
  or_5   g15943(.A(new_n18291), .B(new_n18287), .Y(new_n18292));
  nand_5 g15944(.A(new_n18291), .B(new_n18287), .Y(new_n18293));
  nand_5 g15945(.A(new_n18218), .B(new_n18216), .Y(new_n18294));
  xor_4  g15946(.A(new_n18294), .B(new_n18220), .Y(new_n18295_1));
  nand_5 g15947(.A(new_n18295_1), .B(new_n17458_1), .Y(new_n18296));
  or_5   g15948(.A(new_n18295_1), .B(new_n17458_1), .Y(new_n18297));
  nand_5 g15949(.A(new_n5739), .B(new_n5706), .Y(new_n18298));
  nand_5 g15950(.A(new_n18298), .B(new_n5738), .Y(new_n18299));
  nand_5 g15951(.A(new_n18299), .B(new_n18297), .Y(new_n18300));
  nand_5 g15952(.A(new_n18300), .B(new_n18296), .Y(new_n18301_1));
  nand_5 g15953(.A(new_n18301_1), .B(new_n18293), .Y(new_n18302));
  nand_5 g15954(.A(new_n18302), .B(new_n18292), .Y(new_n18303));
  nand_5 g15955(.A(new_n18303), .B(new_n18286), .Y(new_n18304_1));
  nand_5 g15956(.A(new_n18304_1), .B(new_n18285), .Y(new_n18305));
  nand_5 g15957(.A(new_n18305), .B(new_n18277), .Y(new_n18306));
  nand_5 g15958(.A(new_n18306), .B(new_n18276), .Y(new_n18307));
  nand_5 g15959(.A(new_n18307), .B(new_n18268), .Y(new_n18308));
  nand_5 g15960(.A(new_n18308), .B(new_n18267), .Y(new_n18309));
  nand_5 g15961(.A(new_n18309), .B(new_n18261), .Y(new_n18310_1));
  nand_5 g15962(.A(new_n18310_1), .B(new_n18260), .Y(new_n18311_1));
  xnor_4 g15963(.A(new_n18311_1), .B(new_n18254_1), .Y(n3649));
  nand_5 g15964(.A(new_n10974), .B(new_n7513), .Y(new_n18313));
  or_5   g15965(.A(new_n18313), .B(n26744), .Y(new_n18314));
  nor_5  g15966(.A(new_n18314), .B(n11566), .Y(new_n18315));
  not_8  g15967(.A(new_n18315), .Y(new_n18316));
  nand_5 g15968(.A(new_n18314), .B(n11566), .Y(new_n18317));
  nand_5 g15969(.A(new_n18317), .B(new_n18316), .Y(new_n18318));
  or_5   g15970(.A(new_n18318), .B(n15378), .Y(new_n18319));
  nand_5 g15971(.A(new_n18318), .B(n15378), .Y(new_n18320));
  nand_5 g15972(.A(new_n18313), .B(n26744), .Y(new_n18321));
  nand_5 g15973(.A(new_n18321), .B(new_n18314), .Y(new_n18322));
  or_5   g15974(.A(new_n18322), .B(n17095), .Y(new_n18323_1));
  nand_5 g15975(.A(new_n18322), .B(n17095), .Y(new_n18324));
  nand_5 g15976(.A(n26625), .B(n14230), .Y(new_n18325));
  and_5  g15977(.A(new_n18325), .B(new_n18313), .Y(new_n18326));
  nand_5 g15978(.A(new_n18326), .B(new_n10998), .Y(new_n18327));
  or_5   g15979(.A(new_n18326), .B(new_n10998), .Y(new_n18328));
  nand_5 g15980(.A(n26167), .B(new_n7513), .Y(new_n18329));
  nand_5 g15981(.A(new_n18329), .B(new_n18328), .Y(new_n18330));
  nand_5 g15982(.A(new_n18330), .B(new_n18327), .Y(new_n18331));
  nand_5 g15983(.A(new_n18331), .B(new_n18324), .Y(new_n18332_1));
  nand_5 g15984(.A(new_n18332_1), .B(new_n18323_1), .Y(new_n18333));
  nand_5 g15985(.A(new_n18333), .B(new_n18320), .Y(new_n18334));
  nand_5 g15986(.A(new_n18334), .B(new_n18319), .Y(new_n18335));
  nand_5 g15987(.A(new_n18315), .B(new_n11062), .Y(new_n18336));
  not_8  g15988(.A(new_n18336), .Y(new_n18337));
  nor_5  g15989(.A(new_n18315), .B(new_n11062), .Y(new_n18338));
  or_5   g15990(.A(new_n18338), .B(new_n18337), .Y(new_n18339));
  or_5   g15991(.A(new_n18339), .B(n19575), .Y(new_n18340));
  nand_5 g15992(.A(new_n18339), .B(n19575), .Y(new_n18341));
  nand_5 g15993(.A(new_n18341), .B(new_n18340), .Y(new_n18342));
  xor_4  g15994(.A(new_n18342), .B(new_n18335), .Y(new_n18343_1));
  nand_5 g15995(.A(new_n18343_1), .B(n2013), .Y(new_n18344));
  or_5   g15996(.A(new_n18343_1), .B(n2013), .Y(new_n18345_1));
  nand_5 g15997(.A(new_n18320), .B(new_n18319), .Y(new_n18346));
  xnor_4 g15998(.A(new_n18346), .B(new_n18333), .Y(new_n18347));
  or_5   g15999(.A(new_n18347), .B(new_n16486), .Y(new_n18348));
  nand_5 g16000(.A(new_n18347), .B(new_n16486), .Y(new_n18349));
  nand_5 g16001(.A(new_n18324), .B(new_n18323_1), .Y(new_n18350_1));
  xnor_4 g16002(.A(new_n18350_1), .B(new_n18331), .Y(new_n18351));
  or_5   g16003(.A(new_n18351), .B(new_n16489), .Y(new_n18352));
  nand_5 g16004(.A(new_n18351), .B(new_n16489), .Y(new_n18353));
  nand_5 g16005(.A(new_n18328), .B(new_n18327), .Y(new_n18354));
  xnor_4 g16006(.A(new_n18354), .B(new_n18329), .Y(new_n18355));
  or_5   g16007(.A(new_n18355), .B(new_n16492), .Y(new_n18356));
  nand_5 g16008(.A(new_n18355), .B(new_n16492), .Y(new_n18357));
  nand_5 g16009(.A(new_n8284), .B(n14230), .Y(new_n18358));
  nand_5 g16010(.A(new_n18358), .B(new_n18329), .Y(new_n18359));
  not_8  g16011(.A(new_n18359), .Y(new_n18360));
  nand_5 g16012(.A(new_n18360), .B(n9646), .Y(new_n18361));
  not_8  g16013(.A(new_n18361), .Y(new_n18362_1));
  nand_5 g16014(.A(new_n18362_1), .B(new_n18357), .Y(new_n18363));
  nand_5 g16015(.A(new_n18363), .B(new_n18356), .Y(new_n18364));
  nand_5 g16016(.A(new_n18364), .B(new_n18353), .Y(new_n18365));
  nand_5 g16017(.A(new_n18365), .B(new_n18352), .Y(new_n18366));
  nand_5 g16018(.A(new_n18366), .B(new_n18349), .Y(new_n18367));
  nand_5 g16019(.A(new_n18367), .B(new_n18348), .Y(new_n18368));
  nand_5 g16020(.A(new_n18368), .B(new_n18345_1), .Y(new_n18369));
  nand_5 g16021(.A(new_n18369), .B(new_n18344), .Y(new_n18370));
  nand_5 g16022(.A(new_n18341), .B(new_n18335), .Y(new_n18371));
  nand_5 g16023(.A(new_n18371), .B(new_n18340), .Y(new_n18372));
  nand_5 g16024(.A(new_n18337), .B(new_n12540_1), .Y(new_n18373));
  not_8  g16025(.A(new_n18373), .Y(new_n18374));
  nor_5  g16026(.A(new_n18337), .B(new_n12540_1), .Y(new_n18375));
  or_5   g16027(.A(new_n18375), .B(new_n18374), .Y(new_n18376));
  or_5   g16028(.A(new_n18376), .B(n26512), .Y(new_n18377_1));
  nand_5 g16029(.A(new_n18376), .B(n26512), .Y(new_n18378));
  nand_5 g16030(.A(new_n18378), .B(new_n18377_1), .Y(new_n18379));
  xor_4  g16031(.A(new_n18379), .B(new_n18372), .Y(new_n18380));
  nand_5 g16032(.A(new_n18380), .B(n17302), .Y(new_n18381));
  or_5   g16033(.A(new_n18380), .B(n17302), .Y(new_n18382));
  nand_5 g16034(.A(new_n18382), .B(new_n18381), .Y(new_n18383));
  xor_4  g16035(.A(new_n18383), .B(new_n18370), .Y(new_n18384));
  nand_5 g16036(.A(new_n18384), .B(new_n7902), .Y(new_n18385));
  nor_5  g16037(.A(new_n18384), .B(new_n7902), .Y(new_n18386));
  not_8  g16038(.A(new_n18386), .Y(new_n18387));
  nand_5 g16039(.A(new_n18345_1), .B(new_n18344), .Y(new_n18388));
  xor_4  g16040(.A(new_n18388), .B(new_n18368), .Y(new_n18389));
  nand_5 g16041(.A(new_n18389), .B(new_n7909), .Y(new_n18390));
  nor_5  g16042(.A(new_n18389), .B(new_n7909), .Y(new_n18391));
  not_8  g16043(.A(new_n18391), .Y(new_n18392));
  nand_5 g16044(.A(new_n18349), .B(new_n18348), .Y(new_n18393));
  xor_4  g16045(.A(new_n18393), .B(new_n18366), .Y(new_n18394));
  nand_5 g16046(.A(new_n18394), .B(new_n7916), .Y(new_n18395));
  nor_5  g16047(.A(new_n18394), .B(new_n7916), .Y(new_n18396));
  not_8  g16048(.A(new_n18396), .Y(new_n18397));
  nand_5 g16049(.A(new_n18353), .B(new_n18352), .Y(new_n18398));
  xor_4  g16050(.A(new_n18398), .B(new_n18364), .Y(new_n18399));
  nand_5 g16051(.A(new_n18399), .B(new_n7922), .Y(new_n18400));
  or_5   g16052(.A(new_n18399), .B(new_n7922), .Y(new_n18401));
  not_8  g16053(.A(new_n7928), .Y(new_n18402));
  nand_5 g16054(.A(new_n18357), .B(new_n18356), .Y(new_n18403));
  xor_4  g16055(.A(new_n18403), .B(new_n18361), .Y(new_n18404));
  or_5   g16056(.A(new_n18404), .B(new_n18402), .Y(new_n18405_1));
  nand_5 g16057(.A(new_n18404), .B(new_n18402), .Y(new_n18406));
  nor_5  g16058(.A(new_n18360), .B(n9646), .Y(new_n18407));
  nor_5  g16059(.A(new_n18407), .B(new_n18362_1), .Y(new_n18408));
  nor_5  g16060(.A(new_n18408), .B(new_n13537), .Y(new_n18409_1));
  nand_5 g16061(.A(new_n18409_1), .B(new_n18406), .Y(new_n18410));
  nand_5 g16062(.A(new_n18410), .B(new_n18405_1), .Y(new_n18411));
  nand_5 g16063(.A(new_n18411), .B(new_n18401), .Y(new_n18412));
  nand_5 g16064(.A(new_n18412), .B(new_n18400), .Y(new_n18413));
  nand_5 g16065(.A(new_n18413), .B(new_n18397), .Y(new_n18414_1));
  nand_5 g16066(.A(new_n18414_1), .B(new_n18395), .Y(new_n18415));
  nand_5 g16067(.A(new_n18415), .B(new_n18392), .Y(new_n18416));
  nand_5 g16068(.A(new_n18416), .B(new_n18390), .Y(new_n18417));
  nand_5 g16069(.A(new_n18417), .B(new_n18387), .Y(new_n18418_1));
  nand_5 g16070(.A(new_n18418_1), .B(new_n18385), .Y(new_n18419));
  nand_5 g16071(.A(new_n18382), .B(new_n18370), .Y(new_n18420));
  nand_5 g16072(.A(new_n18420), .B(new_n18381), .Y(new_n18421));
  nand_5 g16073(.A(new_n18378), .B(new_n18372), .Y(new_n18422));
  nand_5 g16074(.A(new_n18422), .B(new_n18377_1), .Y(new_n18423));
  nand_5 g16075(.A(new_n18374), .B(new_n12631), .Y(new_n18424));
  not_8  g16076(.A(new_n18424), .Y(new_n18425));
  nor_5  g16077(.A(new_n18374), .B(new_n12631), .Y(new_n18426));
  or_5   g16078(.A(new_n18426), .B(new_n18425), .Y(new_n18427));
  or_5   g16079(.A(new_n18427), .B(n26191), .Y(new_n18428));
  nand_5 g16080(.A(new_n18427), .B(n26191), .Y(new_n18429));
  nand_5 g16081(.A(new_n18429), .B(new_n18428), .Y(new_n18430));
  xor_4  g16082(.A(new_n18430), .B(new_n18423), .Y(new_n18431));
  nand_5 g16083(.A(new_n18431), .B(n7917), .Y(new_n18432));
  or_5   g16084(.A(new_n18431), .B(n7917), .Y(new_n18433));
  nand_5 g16085(.A(new_n18433), .B(new_n18432), .Y(new_n18434));
  xor_4  g16086(.A(new_n18434), .B(new_n18421), .Y(new_n18435));
  nand_5 g16087(.A(new_n18435), .B(new_n7895), .Y(new_n18436));
  not_8  g16088(.A(new_n18436), .Y(new_n18437_1));
  nor_5  g16089(.A(new_n18435), .B(new_n7895), .Y(new_n18438));
  nor_5  g16090(.A(new_n18438), .B(new_n18437_1), .Y(new_n18439_1));
  xor_4  g16091(.A(new_n18439_1), .B(new_n18419), .Y(n3665));
  xor_4  g16092(.A(new_n6583), .B(new_n6576_1), .Y(n3679));
  nand_5 g16093(.A(new_n9829), .B(new_n9827), .Y(new_n18442));
  nand_5 g16094(.A(new_n18442), .B(new_n9828), .Y(new_n18443));
  nand_5 g16095(.A(new_n6857), .B(n2659), .Y(new_n18444_1));
  nand_5 g16096(.A(new_n6858), .B(new_n5508), .Y(new_n18445_1));
  nand_5 g16097(.A(new_n18445_1), .B(new_n18444_1), .Y(new_n18446));
  xor_4  g16098(.A(new_n18446), .B(new_n18443), .Y(new_n18447));
  not_8  g16099(.A(new_n18447), .Y(new_n18448));
  nand_5 g16100(.A(new_n3746), .B(new_n3748), .Y(new_n18449));
  nand_5 g16101(.A(new_n6766), .B(new_n3748), .Y(new_n18450));
  nand_5 g16102(.A(new_n18450), .B(n16521), .Y(new_n18451));
  nand_5 g16103(.A(new_n18451), .B(new_n18449), .Y(new_n18452_1));
  nand_5 g16104(.A(new_n18452_1), .B(new_n6964), .Y(new_n18453));
  not_8  g16105(.A(new_n18449), .Y(new_n18454));
  nand_5 g16106(.A(new_n18454), .B(new_n6767), .Y(new_n18455));
  nand_5 g16107(.A(new_n18455), .B(new_n18453), .Y(new_n18456));
  xor_4  g16108(.A(new_n18449), .B(n16824), .Y(new_n18457));
  nand_5 g16109(.A(new_n18457), .B(new_n6762), .Y(new_n18458));
  nand_5 g16110(.A(new_n18458), .B(new_n18456), .Y(new_n18459));
  nor_5  g16111(.A(new_n18457), .B(new_n6762), .Y(new_n18460));
  not_8  g16112(.A(new_n18460), .Y(new_n18461));
  nand_5 g16113(.A(new_n18461), .B(new_n18459), .Y(new_n18462));
  nand_5 g16114(.A(new_n18454), .B(new_n3742), .Y(new_n18463));
  xor_4  g16115(.A(new_n18463), .B(n604), .Y(new_n18464));
  nand_5 g16116(.A(new_n18464), .B(new_n6752), .Y(new_n18465));
  nand_5 g16117(.A(new_n18465), .B(new_n18462), .Y(new_n18466));
  not_8  g16118(.A(new_n18466), .Y(new_n18467_1));
  nor_5  g16119(.A(new_n18464), .B(new_n6752), .Y(new_n18468));
  nor_5  g16120(.A(new_n18468), .B(new_n18467_1), .Y(new_n18469));
  not_8  g16121(.A(new_n18469), .Y(new_n18470));
  nor_5  g16122(.A(new_n18463), .B(n604), .Y(new_n18471));
  xor_4  g16123(.A(new_n18471), .B(new_n3734), .Y(new_n18472));
  nand_5 g16124(.A(new_n18472), .B(new_n6745), .Y(new_n18473));
  nand_5 g16125(.A(new_n18473), .B(new_n18470), .Y(new_n18474));
  nor_5  g16126(.A(new_n18472), .B(new_n6745), .Y(new_n18475));
  not_8  g16127(.A(new_n18475), .Y(new_n18476));
  and_5  g16128(.A(new_n18476), .B(new_n18474), .Y(new_n18477));
  not_8  g16129(.A(new_n18477), .Y(new_n18478));
  nand_5 g16130(.A(new_n18471), .B(new_n3734), .Y(new_n18479));
  xor_4  g16131(.A(new_n18479), .B(n9172), .Y(new_n18480));
  nand_5 g16132(.A(new_n18480), .B(new_n6740), .Y(new_n18481));
  nand_5 g16133(.A(new_n18481), .B(new_n18478), .Y(new_n18482_1));
  not_8  g16134(.A(new_n18482_1), .Y(new_n18483_1));
  nor_5  g16135(.A(new_n18480), .B(new_n6740), .Y(new_n18484));
  nor_5  g16136(.A(new_n18484), .B(new_n18483_1), .Y(new_n18485));
  not_8  g16137(.A(new_n18485), .Y(new_n18486));
  nor_5  g16138(.A(new_n18479), .B(n9172), .Y(new_n18487));
  xor_4  g16139(.A(new_n18487), .B(new_n3726), .Y(new_n18488));
  nand_5 g16140(.A(new_n18488), .B(new_n6733), .Y(new_n18489));
  nand_5 g16141(.A(new_n18489), .B(new_n18486), .Y(new_n18490));
  nor_5  g16142(.A(new_n18488), .B(new_n6733), .Y(new_n18491));
  not_8  g16143(.A(new_n18491), .Y(new_n18492));
  nand_5 g16144(.A(new_n18492), .B(new_n18490), .Y(new_n18493));
  nand_5 g16145(.A(new_n18487), .B(new_n3726), .Y(new_n18494));
  xor_4  g16146(.A(new_n18494), .B(n13719), .Y(new_n18495));
  nand_5 g16147(.A(new_n18495), .B(new_n6726), .Y(new_n18496_1));
  nor_5  g16148(.A(new_n18495), .B(new_n6726), .Y(new_n18497));
  not_8  g16149(.A(new_n18497), .Y(new_n18498));
  nand_5 g16150(.A(new_n18498), .B(new_n18496_1), .Y(new_n18499));
  xor_4  g16151(.A(new_n18499), .B(new_n18493), .Y(new_n18500));
  or_5   g16152(.A(new_n18500), .B(new_n18448), .Y(new_n18501));
  not_8  g16153(.A(new_n18501), .Y(new_n18502));
  nand_5 g16154(.A(new_n18500), .B(new_n18448), .Y(new_n18503));
  not_8  g16155(.A(new_n18503), .Y(new_n18504));
  nand_5 g16156(.A(new_n18492), .B(new_n18489), .Y(new_n18505));
  xor_4  g16157(.A(new_n18505), .B(new_n18485), .Y(new_n18506));
  or_5   g16158(.A(new_n18506), .B(new_n9831), .Y(new_n18507));
  nand_5 g16159(.A(new_n18506), .B(new_n9831), .Y(new_n18508));
  not_8  g16160(.A(new_n18481), .Y(new_n18509_1));
  nor_5  g16161(.A(new_n18484), .B(new_n18509_1), .Y(new_n18510));
  xor_4  g16162(.A(new_n18510), .B(new_n18478), .Y(new_n18511));
  or_5   g16163(.A(new_n18511), .B(new_n9756), .Y(new_n18512));
  nand_5 g16164(.A(new_n18511), .B(new_n9756), .Y(new_n18513_1));
  nand_5 g16165(.A(new_n18476), .B(new_n18473), .Y(new_n18514));
  xor_4  g16166(.A(new_n18514), .B(new_n18469), .Y(new_n18515_1));
  or_5   g16167(.A(new_n18515_1), .B(new_n9786), .Y(new_n18516));
  nand_5 g16168(.A(new_n18515_1), .B(new_n9786), .Y(new_n18517));
  not_8  g16169(.A(new_n9792), .Y(new_n18518));
  not_8  g16170(.A(new_n18468), .Y(new_n18519));
  nand_5 g16171(.A(new_n18519), .B(new_n18465), .Y(new_n18520));
  xor_4  g16172(.A(new_n18520), .B(new_n18462), .Y(new_n18521));
  nand_5 g16173(.A(new_n18521), .B(new_n18518), .Y(new_n18522));
  or_5   g16174(.A(new_n18521), .B(new_n18518), .Y(new_n18523));
  not_8  g16175(.A(new_n9798), .Y(new_n18524));
  nand_5 g16176(.A(new_n18461), .B(new_n18458), .Y(new_n18525));
  xor_4  g16177(.A(new_n18525), .B(new_n18456), .Y(new_n18526));
  nand_5 g16178(.A(new_n18526), .B(new_n18524), .Y(new_n18527));
  or_5   g16179(.A(new_n18526), .B(new_n18524), .Y(new_n18528));
  nand_5 g16180(.A(new_n18455), .B(new_n18452_1), .Y(new_n18529));
  xor_4  g16181(.A(new_n18529), .B(new_n6964), .Y(new_n18530));
  nand_5 g16182(.A(new_n18530), .B(new_n9805), .Y(new_n18531));
  nor_5  g16183(.A(new_n18530), .B(new_n9805), .Y(new_n18532));
  not_8  g16184(.A(new_n18532), .Y(new_n18533));
  not_8  g16185(.A(new_n9811), .Y(new_n18534));
  nand_5 g16186(.A(new_n6767), .B(n7139), .Y(new_n18535));
  nand_5 g16187(.A(new_n18535), .B(new_n18450), .Y(new_n18536));
  nor_5  g16188(.A(new_n18536), .B(new_n18534), .Y(new_n18537_1));
  nand_5 g16189(.A(new_n18537_1), .B(new_n18533), .Y(new_n18538));
  nand_5 g16190(.A(new_n18538), .B(new_n18531), .Y(new_n18539));
  nand_5 g16191(.A(new_n18539), .B(new_n18528), .Y(new_n18540));
  nand_5 g16192(.A(new_n18540), .B(new_n18527), .Y(new_n18541));
  nand_5 g16193(.A(new_n18541), .B(new_n18523), .Y(new_n18542));
  nand_5 g16194(.A(new_n18542), .B(new_n18522), .Y(new_n18543));
  nand_5 g16195(.A(new_n18543), .B(new_n18517), .Y(new_n18544));
  nand_5 g16196(.A(new_n18544), .B(new_n18516), .Y(new_n18545));
  nand_5 g16197(.A(new_n18545), .B(new_n18513_1), .Y(new_n18546));
  nand_5 g16198(.A(new_n18546), .B(new_n18512), .Y(new_n18547));
  nand_5 g16199(.A(new_n18547), .B(new_n18508), .Y(new_n18548));
  nand_5 g16200(.A(new_n18548), .B(new_n18507), .Y(new_n18549));
  nor_5  g16201(.A(new_n18549), .B(new_n18504), .Y(new_n18550));
  nor_5  g16202(.A(new_n18550), .B(new_n18502), .Y(new_n18551));
  nand_5 g16203(.A(new_n18496_1), .B(new_n18493), .Y(new_n18552));
  nand_5 g16204(.A(new_n18552), .B(new_n18498), .Y(new_n18553));
  nor_5  g16205(.A(new_n18494), .B(n13719), .Y(new_n18554));
  nand_5 g16206(.A(new_n18554), .B(new_n3718), .Y(new_n18555));
  or_5   g16207(.A(new_n18554), .B(new_n3718), .Y(new_n18556));
  and_5  g16208(.A(new_n18556), .B(new_n18555), .Y(new_n18557));
  or_5   g16209(.A(new_n18557), .B(new_n6719), .Y(new_n18558_1));
  nand_5 g16210(.A(new_n18557), .B(new_n6719), .Y(new_n18559));
  nand_5 g16211(.A(new_n18559), .B(new_n18558_1), .Y(new_n18560));
  xor_4  g16212(.A(new_n18560), .B(new_n18553), .Y(new_n18561));
  nand_5 g16213(.A(new_n18445_1), .B(new_n18443), .Y(new_n18562));
  nand_5 g16214(.A(new_n18562), .B(new_n18444_1), .Y(new_n18563));
  nand_5 g16215(.A(new_n6851), .B(n2858), .Y(new_n18564));
  nand_5 g16216(.A(new_n6852), .B(new_n5502), .Y(new_n18565));
  nand_5 g16217(.A(new_n18565), .B(new_n18564), .Y(new_n18566));
  xor_4  g16218(.A(new_n18566), .B(new_n18563), .Y(new_n18567));
  not_8  g16219(.A(new_n18567), .Y(new_n18568));
  or_5   g16220(.A(new_n18568), .B(new_n18561), .Y(new_n18569));
  not_8  g16221(.A(new_n18569), .Y(new_n18570));
  nand_5 g16222(.A(new_n18568), .B(new_n18561), .Y(new_n18571));
  not_8  g16223(.A(new_n18571), .Y(new_n18572_1));
  nor_5  g16224(.A(new_n18572_1), .B(new_n18570), .Y(new_n18573));
  xor_4  g16225(.A(new_n18573), .B(new_n18551), .Y(n3725));
  nand_5 g16226(.A(new_n14897), .B(new_n14893), .Y(new_n18575));
  nand_5 g16227(.A(new_n18575), .B(new_n14894), .Y(new_n18576_1));
  not_8  g16228(.A(new_n18576_1), .Y(new_n18577));
  nand_5 g16229(.A(new_n14903), .B(new_n14899_1), .Y(new_n18578_1));
  nand_5 g16230(.A(new_n18578_1), .B(new_n14900), .Y(new_n18579));
  or_5   g16231(.A(new_n18579), .B(new_n18577), .Y(new_n18580));
  nand_5 g16232(.A(new_n18579), .B(new_n18577), .Y(new_n18581));
  nand_5 g16233(.A(new_n18581), .B(new_n18580), .Y(new_n18582_1));
  nand_5 g16234(.A(new_n14910), .B(new_n14907), .Y(new_n18583_1));
  nand_5 g16235(.A(new_n18583_1), .B(new_n14906), .Y(new_n18584_1));
  xor_4  g16236(.A(new_n18584_1), .B(new_n18582_1), .Y(new_n18585));
  nand_5 g16237(.A(new_n18585), .B(new_n16870), .Y(new_n18586));
  not_8  g16238(.A(new_n18585), .Y(new_n18587));
  nand_5 g16239(.A(new_n18587), .B(new_n16868), .Y(new_n18588));
  nand_5 g16240(.A(new_n18588), .B(new_n18586), .Y(new_n18589));
  nand_5 g16241(.A(new_n16875), .B(new_n14912), .Y(new_n18590));
  nand_5 g16242(.A(new_n16874), .B(new_n14911), .Y(new_n18591));
  nand_5 g16243(.A(new_n16879), .B(new_n6154), .Y(new_n18592));
  nand_5 g16244(.A(new_n16881), .B(new_n6153), .Y(new_n18593));
  nand_5 g16245(.A(new_n16884), .B(new_n6071), .Y(new_n18594));
  nand_5 g16246(.A(new_n16886), .B(new_n6070), .Y(new_n18595));
  nand_5 g16247(.A(new_n16889), .B(new_n6077), .Y(new_n18596));
  or_5   g16248(.A(new_n16889), .B(new_n6077), .Y(new_n18597));
  nand_5 g16249(.A(new_n16823), .B(new_n6083), .Y(new_n18598));
  or_5   g16250(.A(new_n16823), .B(new_n6083), .Y(new_n18599));
  nand_5 g16251(.A(new_n6090), .B(new_n4788), .Y(new_n18600));
  or_5   g16252(.A(new_n6090), .B(new_n4788), .Y(new_n18601));
  nand_5 g16253(.A(new_n6097), .B(new_n4716), .Y(new_n18602));
  nand_5 g16254(.A(new_n6096), .B(new_n4717), .Y(new_n18603));
  nand_5 g16255(.A(new_n6102), .B(new_n4669), .Y(new_n18604));
  nand_5 g16256(.A(new_n6101), .B(new_n4668), .Y(new_n18605));
  or_5   g16257(.A(new_n6110), .B(new_n4747_1), .Y(new_n18606));
  nand_5 g16258(.A(new_n6110), .B(new_n4747_1), .Y(new_n18607));
  not_8  g16259(.A(new_n4699), .Y(new_n18608));
  nor_5  g16260(.A(new_n6114), .B(new_n18608), .Y(new_n18609));
  nand_5 g16261(.A(new_n18609), .B(new_n18607), .Y(new_n18610_1));
  nand_5 g16262(.A(new_n18610_1), .B(new_n18606), .Y(new_n18611));
  nand_5 g16263(.A(new_n18611), .B(new_n18605), .Y(new_n18612));
  nand_5 g16264(.A(new_n18612), .B(new_n18604), .Y(new_n18613));
  nand_5 g16265(.A(new_n18613), .B(new_n18603), .Y(new_n18614));
  nand_5 g16266(.A(new_n18614), .B(new_n18602), .Y(new_n18615));
  nand_5 g16267(.A(new_n18615), .B(new_n18601), .Y(new_n18616));
  nand_5 g16268(.A(new_n18616), .B(new_n18600), .Y(new_n18617));
  nand_5 g16269(.A(new_n18617), .B(new_n18599), .Y(new_n18618));
  nand_5 g16270(.A(new_n18618), .B(new_n18598), .Y(new_n18619));
  nand_5 g16271(.A(new_n18619), .B(new_n18597), .Y(new_n18620));
  nand_5 g16272(.A(new_n18620), .B(new_n18596), .Y(new_n18621));
  nand_5 g16273(.A(new_n18621), .B(new_n18595), .Y(new_n18622));
  nand_5 g16274(.A(new_n18622), .B(new_n18594), .Y(new_n18623));
  nand_5 g16275(.A(new_n18623), .B(new_n18593), .Y(new_n18624));
  nand_5 g16276(.A(new_n18624), .B(new_n18592), .Y(new_n18625));
  nand_5 g16277(.A(new_n18625), .B(new_n18591), .Y(new_n18626));
  nand_5 g16278(.A(new_n18626), .B(new_n18590), .Y(new_n18627));
  not_8  g16279(.A(new_n18627), .Y(new_n18628));
  xor_4  g16280(.A(new_n18628), .B(new_n18589), .Y(n3733));
  nand_5 g16281(.A(new_n17542), .B(new_n17538), .Y(new_n18630));
  nand_5 g16282(.A(new_n18630), .B(new_n17539), .Y(new_n18631));
  nand_5 g16283(.A(new_n12372), .B(n5098), .Y(new_n18632));
  nand_5 g16284(.A(new_n12373), .B(new_n17594), .Y(new_n18633));
  nand_5 g16285(.A(new_n18633), .B(new_n18632), .Y(new_n18634));
  xor_4  g16286(.A(new_n18634), .B(new_n18631), .Y(new_n18635_1));
  or_5   g16287(.A(new_n18635_1), .B(new_n11565), .Y(new_n18636));
  nand_5 g16288(.A(new_n18635_1), .B(new_n11565), .Y(new_n18637));
  nand_5 g16289(.A(new_n17546), .B(new_n17536), .Y(new_n18638));
  nand_5 g16290(.A(new_n18638), .B(new_n17545), .Y(new_n18639));
  nand_5 g16291(.A(new_n18639), .B(new_n18637), .Y(new_n18640));
  nand_5 g16292(.A(new_n18640), .B(new_n18636), .Y(new_n18641));
  nand_5 g16293(.A(new_n18633), .B(new_n18631), .Y(new_n18642));
  nand_5 g16294(.A(new_n18642), .B(new_n18632), .Y(new_n18643));
  nand_5 g16295(.A(new_n12380_1), .B(n24937), .Y(new_n18644));
  not_8  g16296(.A(new_n12380_1), .Y(new_n18645));
  nand_5 g16297(.A(new_n18645), .B(new_n17605), .Y(new_n18646));
  nand_5 g16298(.A(new_n18646), .B(new_n18644), .Y(new_n18647));
  xor_4  g16299(.A(new_n18647), .B(new_n18643), .Y(new_n18648));
  or_5   g16300(.A(new_n18648), .B(new_n11557), .Y(new_n18649_1));
  nand_5 g16301(.A(new_n18648), .B(new_n11557), .Y(new_n18650));
  nand_5 g16302(.A(new_n18650), .B(new_n18649_1), .Y(new_n18651));
  xor_4  g16303(.A(new_n18651), .B(new_n18641), .Y(n3755));
  nand_5 g16304(.A(new_n10398), .B(new_n10397), .Y(new_n18653_1));
  xor_4  g16305(.A(new_n18653_1), .B(new_n10442), .Y(n3758));
  not_8  g16306(.A(n19033), .Y(new_n18655));
  nand_5 g16307(.A(new_n17985), .B(new_n17984), .Y(new_n18656));
  nor_5  g16308(.A(new_n18656), .B(n655), .Y(new_n18657));
  nand_5 g16309(.A(new_n18657), .B(new_n18655), .Y(new_n18658));
  nor_5  g16310(.A(new_n18658), .B(n2570), .Y(new_n18659));
  xor_4  g16311(.A(new_n18658), .B(n2570), .Y(new_n18660));
  nand_5 g16312(.A(new_n18660), .B(new_n11978), .Y(new_n18661));
  or_5   g16313(.A(new_n18660), .B(new_n11978), .Y(new_n18662));
  xor_4  g16314(.A(new_n18657), .B(new_n18655), .Y(new_n18663));
  nand_5 g16315(.A(new_n18663), .B(new_n11980_1), .Y(new_n18664));
  or_5   g16316(.A(new_n18663), .B(new_n11980_1), .Y(new_n18665));
  xor_4  g16317(.A(new_n18656), .B(n655), .Y(new_n18666));
  nand_5 g16318(.A(new_n18666), .B(new_n11983), .Y(new_n18667));
  or_5   g16319(.A(new_n18666), .B(new_n11983), .Y(new_n18668));
  nand_5 g16320(.A(new_n17988), .B(new_n17983), .Y(new_n18669));
  nand_5 g16321(.A(new_n18669), .B(new_n17987), .Y(new_n18670));
  nand_5 g16322(.A(new_n18670), .B(new_n18668), .Y(new_n18671));
  nand_5 g16323(.A(new_n18671), .B(new_n18667), .Y(new_n18672));
  nand_5 g16324(.A(new_n18672), .B(new_n18665), .Y(new_n18673));
  nand_5 g16325(.A(new_n18673), .B(new_n18664), .Y(new_n18674));
  nand_5 g16326(.A(new_n18674), .B(new_n18662), .Y(new_n18675));
  nand_5 g16327(.A(new_n18675), .B(new_n18661), .Y(new_n18676));
  and_5  g16328(.A(new_n18676), .B(new_n18659), .Y(new_n18677));
  nor_5  g16329(.A(new_n18676), .B(new_n18659), .Y(new_n18678));
  nor_5  g16330(.A(new_n18678), .B(new_n18677), .Y(new_n18679_1));
  or_5   g16331(.A(new_n18679_1), .B(new_n13748), .Y(new_n18680));
  nand_5 g16332(.A(new_n18662), .B(new_n18661), .Y(new_n18681));
  xor_4  g16333(.A(new_n18681), .B(new_n18674), .Y(new_n18682));
  nand_5 g16334(.A(new_n18682), .B(new_n13750), .Y(new_n18683));
  or_5   g16335(.A(new_n18682), .B(new_n13750), .Y(new_n18684));
  nand_5 g16336(.A(new_n18665), .B(new_n18664), .Y(new_n18685));
  xor_4  g16337(.A(new_n18685), .B(new_n18672), .Y(new_n18686));
  nand_5 g16338(.A(new_n18686), .B(new_n7978), .Y(new_n18687));
  or_5   g16339(.A(new_n18686), .B(new_n7978), .Y(new_n18688));
  nand_5 g16340(.A(new_n18668), .B(new_n18667), .Y(new_n18689));
  xor_4  g16341(.A(new_n18689), .B(new_n18670), .Y(new_n18690_1));
  nand_5 g16342(.A(new_n18690_1), .B(new_n7885), .Y(new_n18691));
  or_5   g16343(.A(new_n18690_1), .B(new_n7885), .Y(new_n18692));
  nand_5 g16344(.A(new_n17992), .B(new_n17981), .Y(new_n18693_1));
  nand_5 g16345(.A(new_n18693_1), .B(new_n17991), .Y(new_n18694));
  nand_5 g16346(.A(new_n18694), .B(new_n18692), .Y(new_n18695));
  nand_5 g16347(.A(new_n18695), .B(new_n18691), .Y(new_n18696));
  nand_5 g16348(.A(new_n18696), .B(new_n18688), .Y(new_n18697));
  nand_5 g16349(.A(new_n18697), .B(new_n18687), .Y(new_n18698));
  nand_5 g16350(.A(new_n18698), .B(new_n18684), .Y(new_n18699));
  nand_5 g16351(.A(new_n18699), .B(new_n18683), .Y(new_n18700));
  not_8  g16352(.A(new_n18700), .Y(new_n18701));
  nand_5 g16353(.A(new_n18701), .B(new_n18680), .Y(new_n18702));
  nand_5 g16354(.A(new_n18679_1), .B(new_n13748), .Y(new_n18703));
  not_8  g16355(.A(new_n18703), .Y(new_n18704));
  nor_5  g16356(.A(new_n18704), .B(new_n18677), .Y(new_n18705));
  nand_5 g16357(.A(new_n18705), .B(new_n18702), .Y(new_n18706));
  not_8  g16358(.A(new_n11973), .Y(new_n18707));
  nand_5 g16359(.A(new_n18703), .B(new_n18680), .Y(new_n18708_1));
  xor_4  g16360(.A(new_n18708_1), .B(new_n18701), .Y(new_n18709));
  or_5   g16361(.A(new_n18709), .B(new_n18707), .Y(new_n18710));
  nand_5 g16362(.A(new_n18709), .B(new_n18707), .Y(new_n18711));
  nand_5 g16363(.A(new_n18684), .B(new_n18683), .Y(new_n18712));
  xor_4  g16364(.A(new_n18712), .B(new_n18698), .Y(new_n18713));
  nand_5 g16365(.A(new_n18713), .B(new_n11965_1), .Y(new_n18714));
  or_5   g16366(.A(new_n18713), .B(new_n11965_1), .Y(new_n18715));
  nand_5 g16367(.A(new_n18688), .B(new_n18687), .Y(new_n18716));
  xor_4  g16368(.A(new_n18716), .B(new_n18696), .Y(new_n18717));
  nand_5 g16369(.A(new_n18717), .B(new_n11910), .Y(new_n18718));
  or_5   g16370(.A(new_n18717), .B(new_n11910), .Y(new_n18719));
  nand_5 g16371(.A(new_n18692), .B(new_n18691), .Y(new_n18720));
  xor_4  g16372(.A(new_n18720), .B(new_n18694), .Y(new_n18721_1));
  nand_5 g16373(.A(new_n18721_1), .B(new_n11915), .Y(new_n18722));
  or_5   g16374(.A(new_n18721_1), .B(new_n11915), .Y(new_n18723));
  nand_5 g16375(.A(new_n17996), .B(new_n17978), .Y(new_n18724));
  nand_5 g16376(.A(new_n18724), .B(new_n17995), .Y(new_n18725_1));
  nand_5 g16377(.A(new_n18725_1), .B(new_n18723), .Y(new_n18726));
  nand_5 g16378(.A(new_n18726), .B(new_n18722), .Y(new_n18727));
  nand_5 g16379(.A(new_n18727), .B(new_n18719), .Y(new_n18728));
  nand_5 g16380(.A(new_n18728), .B(new_n18718), .Y(new_n18729));
  nand_5 g16381(.A(new_n18729), .B(new_n18715), .Y(new_n18730));
  nand_5 g16382(.A(new_n18730), .B(new_n18714), .Y(new_n18731));
  nand_5 g16383(.A(new_n18731), .B(new_n18711), .Y(new_n18732));
  nand_5 g16384(.A(new_n18732), .B(new_n18710), .Y(new_n18733));
  xnor_4 g16385(.A(new_n18733), .B(new_n18706), .Y(n3760));
  nand_5 g16386(.A(new_n4244), .B(new_n4243), .Y(new_n18735));
  xnor_4 g16387(.A(new_n18735), .B(new_n4272_1), .Y(n3781));
  nand_5 g16388(.A(new_n15437), .B(new_n15438_1), .Y(new_n18737_1));
  xnor_4 g16389(.A(new_n18737_1), .B(new_n15464), .Y(n3794));
  nand_5 g16390(.A(new_n6774), .B(new_n6766), .Y(new_n18739));
  nand_5 g16391(.A(new_n6773_1), .B(new_n6767), .Y(new_n18740));
  nand_5 g16392(.A(new_n18740), .B(new_n18739), .Y(new_n18741));
  nand_5 g16393(.A(new_n18741), .B(new_n14940), .Y(new_n18742));
  not_8  g16394(.A(new_n18742), .Y(new_n18743));
  nor_5  g16395(.A(new_n18741), .B(new_n14940), .Y(new_n18744));
  nor_5  g16396(.A(new_n18744), .B(new_n18743), .Y(new_n18745_1));
  xor_4  g16397(.A(new_n18745_1), .B(new_n12530), .Y(new_n18746));
  nand_5 g16398(.A(new_n12534), .B(new_n5637), .Y(new_n18747));
  nand_5 g16399(.A(new_n12533), .B(new_n5639), .Y(new_n18748));
  nand_5 g16400(.A(new_n18748), .B(new_n18747), .Y(new_n18749));
  xnor_4 g16401(.A(new_n18749), .B(new_n18746), .Y(n3842));
  nand_5 g16402(.A(new_n14070), .B(new_n14072), .Y(new_n18751_1));
  xor_4  g16403(.A(new_n18751_1), .B(new_n10233), .Y(n3850));
  nand_5 g16404(.A(new_n16801), .B(new_n16803), .Y(new_n18753));
  xor_4  g16405(.A(new_n18753), .B(new_n16805), .Y(n3869));
  nand_5 g16406(.A(n21138), .B(n20385), .Y(new_n18755));
  nand_5 g16407(.A(new_n4535), .B(new_n10973), .Y(new_n18756));
  nand_5 g16408(.A(n25316), .B(n7769), .Y(new_n18757));
  nand_5 g16409(.A(new_n18757), .B(new_n18756), .Y(new_n18758));
  xnor_4 g16410(.A(new_n18758), .B(new_n18755), .Y(new_n18759));
  xor_4  g16411(.A(n21138), .B(n20385), .Y(new_n18760));
  not_8  g16412(.A(new_n18760), .Y(new_n18761));
  nand_5 g16413(.A(new_n18761), .B(n15332), .Y(new_n18762));
  not_8  g16414(.A(new_n18762), .Y(new_n18763));
  nand_5 g16415(.A(new_n18763), .B(n5060), .Y(new_n18764));
  or_5   g16416(.A(new_n18763), .B(n5060), .Y(new_n18765));
  nand_5 g16417(.A(new_n18765), .B(new_n18764), .Y(new_n18766));
  xor_4  g16418(.A(new_n18766), .B(new_n18759), .Y(new_n18767));
  or_5   g16419(.A(new_n18767), .B(new_n17812), .Y(new_n18768));
  nand_5 g16420(.A(new_n18767), .B(new_n17812), .Y(new_n18769));
  xor_4  g16421(.A(new_n18760), .B(n15332), .Y(new_n18770));
  nand_5 g16422(.A(new_n18770), .B(new_n17818), .Y(new_n18771));
  nand_5 g16423(.A(new_n18771), .B(new_n18769), .Y(new_n18772));
  nand_5 g16424(.A(new_n18772), .B(new_n18768), .Y(new_n18773));
  nand_5 g16425(.A(new_n18765), .B(new_n18759), .Y(new_n18774));
  nand_5 g16426(.A(new_n18774), .B(new_n18764), .Y(new_n18775));
  not_8  g16427(.A(n19584), .Y(new_n18776));
  nand_5 g16428(.A(new_n18757), .B(new_n18755), .Y(new_n18777));
  nand_5 g16429(.A(new_n18777), .B(new_n18756), .Y(new_n18778));
  not_8  g16430(.A(new_n18778), .Y(new_n18779));
  nand_5 g16431(.A(new_n10969), .B(new_n4586), .Y(new_n18780_1));
  nand_5 g16432(.A(n21749), .B(n919), .Y(new_n18781));
  nand_5 g16433(.A(new_n18781), .B(new_n18780_1), .Y(new_n18782_1));
  xor_4  g16434(.A(new_n18782_1), .B(new_n18779), .Y(new_n18783));
  not_8  g16435(.A(new_n18783), .Y(new_n18784));
  nand_5 g16436(.A(new_n18784), .B(new_n18776), .Y(new_n18785));
  nand_5 g16437(.A(new_n18783), .B(n19584), .Y(new_n18786));
  nand_5 g16438(.A(new_n18786), .B(new_n18785), .Y(new_n18787));
  xor_4  g16439(.A(new_n18787), .B(new_n18775), .Y(new_n18788));
  or_5   g16440(.A(new_n18788), .B(new_n17804), .Y(new_n18789));
  nand_5 g16441(.A(new_n18788), .B(new_n17804), .Y(new_n18790));
  nand_5 g16442(.A(new_n18790), .B(new_n18789), .Y(new_n18791));
  xor_4  g16443(.A(new_n18791), .B(new_n18773), .Y(n3871));
  nand_5 g16444(.A(new_n18528), .B(new_n18527), .Y(new_n18793));
  xnor_4 g16445(.A(new_n18793), .B(new_n18539), .Y(n3891));
  not_8  g16446(.A(n2570), .Y(new_n18795));
  nand_5 g16447(.A(n10250), .B(new_n18795), .Y(new_n18796));
  nand_5 g16448(.A(new_n7040), .B(n2570), .Y(new_n18797));
  nand_5 g16449(.A(new_n18797), .B(new_n18796), .Y(new_n18798));
  nand_5 g16450(.A(new_n18655), .B(n7674), .Y(new_n18799));
  nand_5 g16451(.A(n19033), .B(new_n6991), .Y(new_n18800));
  not_8  g16452(.A(n655), .Y(new_n18801));
  nand_5 g16453(.A(n6397), .B(new_n18801), .Y(new_n18802_1));
  nand_5 g16454(.A(new_n6997), .B(n655), .Y(new_n18803));
  nand_5 g16455(.A(n19196), .B(new_n17984), .Y(new_n18804));
  nand_5 g16456(.A(new_n7003), .B(n18145), .Y(new_n18805));
  not_8  g16457(.A(n10712), .Y(new_n18806));
  nand_5 g16458(.A(n23586), .B(new_n18806), .Y(new_n18807));
  nand_5 g16459(.A(new_n7118), .B(n10712), .Y(new_n18808));
  nand_5 g16460(.A(new_n17895), .B(n21226), .Y(new_n18809));
  nand_5 g16461(.A(n25126), .B(new_n7009), .Y(new_n18810));
  not_8  g16462(.A(n19608), .Y(new_n18811));
  nand_5 g16463(.A(new_n18811), .B(n4426), .Y(new_n18812));
  nand_5 g16464(.A(n19608), .B(new_n7012), .Y(new_n18813));
  nand_5 g16465(.A(new_n4607), .B(new_n4602), .Y(new_n18814));
  nand_5 g16466(.A(new_n18814), .B(new_n4605), .Y(new_n18815));
  nand_5 g16467(.A(new_n18815), .B(new_n18813), .Y(new_n18816));
  nand_5 g16468(.A(new_n18816), .B(new_n18812), .Y(new_n18817));
  nand_5 g16469(.A(new_n18817), .B(new_n18810), .Y(new_n18818));
  nand_5 g16470(.A(new_n18818), .B(new_n18809), .Y(new_n18819));
  nand_5 g16471(.A(new_n18819), .B(new_n18808), .Y(new_n18820));
  nand_5 g16472(.A(new_n18820), .B(new_n18807), .Y(new_n18821));
  nand_5 g16473(.A(new_n18821), .B(new_n18805), .Y(new_n18822));
  nand_5 g16474(.A(new_n18822), .B(new_n18804), .Y(new_n18823));
  nand_5 g16475(.A(new_n18823), .B(new_n18803), .Y(new_n18824));
  nand_5 g16476(.A(new_n18824), .B(new_n18802_1), .Y(new_n18825));
  nand_5 g16477(.A(new_n18825), .B(new_n18800), .Y(new_n18826));
  nand_5 g16478(.A(new_n18826), .B(new_n18799), .Y(new_n18827));
  not_8  g16479(.A(new_n18827), .Y(new_n18828));
  xor_4  g16480(.A(new_n18828), .B(new_n18798), .Y(new_n18829));
  nand_5 g16481(.A(new_n18829), .B(new_n13751), .Y(new_n18830_1));
  not_8  g16482(.A(new_n18829), .Y(new_n18831_1));
  nand_5 g16483(.A(new_n18831_1), .B(new_n13750), .Y(new_n18832));
  nand_5 g16484(.A(new_n18832), .B(new_n18830_1), .Y(new_n18833));
  nand_5 g16485(.A(new_n18800), .B(new_n18799), .Y(new_n18834));
  xor_4  g16486(.A(new_n18834), .B(new_n18825), .Y(new_n18835));
  nand_5 g16487(.A(new_n18835), .B(new_n7978), .Y(new_n18836));
  not_8  g16488(.A(new_n18835), .Y(new_n18837));
  nand_5 g16489(.A(new_n18837), .B(new_n7979), .Y(new_n18838));
  nand_5 g16490(.A(new_n18803), .B(new_n18802_1), .Y(new_n18839));
  xor_4  g16491(.A(new_n18839), .B(new_n18823), .Y(new_n18840));
  nand_5 g16492(.A(new_n18840), .B(new_n7885), .Y(new_n18841));
  not_8  g16493(.A(new_n18840), .Y(new_n18842));
  nand_5 g16494(.A(new_n18842), .B(new_n7886), .Y(new_n18843_1));
  nand_5 g16495(.A(new_n18805), .B(new_n18804), .Y(new_n18844));
  xor_4  g16496(.A(new_n18844), .B(new_n18821), .Y(new_n18845));
  nand_5 g16497(.A(new_n18845), .B(new_n7841_1), .Y(new_n18846));
  not_8  g16498(.A(new_n18845), .Y(new_n18847));
  nand_5 g16499(.A(new_n18847), .B(new_n7842), .Y(new_n18848));
  nand_5 g16500(.A(new_n18808), .B(new_n18807), .Y(new_n18849));
  xor_4  g16501(.A(new_n18849), .B(new_n18819), .Y(new_n18850));
  nand_5 g16502(.A(new_n18850), .B(new_n7848), .Y(new_n18851));
  not_8  g16503(.A(new_n18850), .Y(new_n18852));
  nand_5 g16504(.A(new_n18852), .B(new_n7846), .Y(new_n18853));
  nand_5 g16505(.A(new_n18810), .B(new_n18809), .Y(new_n18854));
  xor_4  g16506(.A(new_n18854), .B(new_n18817), .Y(new_n18855));
  nand_5 g16507(.A(new_n18855), .B(new_n7853), .Y(new_n18856));
  not_8  g16508(.A(new_n18855), .Y(new_n18857));
  nand_5 g16509(.A(new_n18857), .B(new_n7851), .Y(new_n18858_1));
  nand_5 g16510(.A(new_n18813), .B(new_n18812), .Y(new_n18859_1));
  xor_4  g16511(.A(new_n18859_1), .B(new_n18815), .Y(new_n18860));
  nand_5 g16512(.A(new_n18860), .B(new_n7858), .Y(new_n18861));
  not_8  g16513(.A(new_n18860), .Y(new_n18862));
  nand_5 g16514(.A(new_n18862), .B(new_n7856), .Y(new_n18863));
  nand_5 g16515(.A(new_n4613), .B(new_n4592), .Y(new_n18864_1));
  nand_5 g16516(.A(new_n18864_1), .B(new_n4611), .Y(new_n18865_1));
  nand_5 g16517(.A(new_n18865_1), .B(new_n18863), .Y(new_n18866));
  nand_5 g16518(.A(new_n18866), .B(new_n18861), .Y(new_n18867));
  nand_5 g16519(.A(new_n18867), .B(new_n18858_1), .Y(new_n18868));
  nand_5 g16520(.A(new_n18868), .B(new_n18856), .Y(new_n18869));
  nand_5 g16521(.A(new_n18869), .B(new_n18853), .Y(new_n18870));
  nand_5 g16522(.A(new_n18870), .B(new_n18851), .Y(new_n18871));
  nand_5 g16523(.A(new_n18871), .B(new_n18848), .Y(new_n18872));
  nand_5 g16524(.A(new_n18872), .B(new_n18846), .Y(new_n18873));
  nand_5 g16525(.A(new_n18873), .B(new_n18843_1), .Y(new_n18874));
  nand_5 g16526(.A(new_n18874), .B(new_n18841), .Y(new_n18875));
  nand_5 g16527(.A(new_n18875), .B(new_n18838), .Y(new_n18876));
  nand_5 g16528(.A(new_n18876), .B(new_n18836), .Y(new_n18877));
  xor_4  g16529(.A(new_n18877), .B(new_n18833), .Y(new_n18878));
  nand_5 g16530(.A(new_n18878), .B(new_n7211), .Y(new_n18879));
  or_5   g16531(.A(new_n18878), .B(new_n7211), .Y(new_n18880_1));
  nand_5 g16532(.A(new_n18880_1), .B(new_n18879), .Y(new_n18881));
  nand_5 g16533(.A(new_n18836), .B(new_n18838), .Y(new_n18882));
  xor_4  g16534(.A(new_n18882), .B(new_n18875), .Y(new_n18883));
  nand_5 g16535(.A(new_n18883), .B(new_n7218), .Y(new_n18884));
  or_5   g16536(.A(new_n18883), .B(new_n7218), .Y(new_n18885));
  nand_5 g16537(.A(new_n18841), .B(new_n18843_1), .Y(new_n18886_1));
  xor_4  g16538(.A(new_n18886_1), .B(new_n18873), .Y(new_n18887_1));
  nand_5 g16539(.A(new_n18887_1), .B(new_n7227), .Y(new_n18888));
  or_5   g16540(.A(new_n18887_1), .B(new_n7227), .Y(new_n18889));
  nand_5 g16541(.A(new_n18846), .B(new_n18848), .Y(new_n18890));
  xor_4  g16542(.A(new_n18890), .B(new_n18871), .Y(new_n18891));
  nand_5 g16543(.A(new_n18891), .B(new_n7236_1), .Y(new_n18892));
  or_5   g16544(.A(new_n18891), .B(new_n7236_1), .Y(new_n18893));
  nand_5 g16545(.A(new_n18851), .B(new_n18853), .Y(new_n18894));
  xor_4  g16546(.A(new_n18894), .B(new_n18869), .Y(new_n18895));
  nand_5 g16547(.A(new_n18895), .B(new_n7243), .Y(new_n18896));
  or_5   g16548(.A(new_n18895), .B(new_n7243), .Y(new_n18897));
  nand_5 g16549(.A(new_n18856), .B(new_n18858_1), .Y(new_n18898));
  xor_4  g16550(.A(new_n18898), .B(new_n18867), .Y(new_n18899));
  nand_5 g16551(.A(new_n18899), .B(new_n7251), .Y(new_n18900));
  or_5   g16552(.A(new_n18899), .B(new_n7251), .Y(new_n18901_1));
  nand_5 g16553(.A(new_n18861), .B(new_n18863), .Y(new_n18902));
  xor_4  g16554(.A(new_n18902), .B(new_n18865_1), .Y(new_n18903));
  nand_5 g16555(.A(new_n18903), .B(new_n7259), .Y(new_n18904));
  or_5   g16556(.A(new_n18903), .B(new_n7259), .Y(new_n18905));
  nand_5 g16557(.A(new_n4617), .B(new_n4583), .Y(new_n18906));
  nand_5 g16558(.A(new_n18906), .B(new_n4616), .Y(new_n18907_1));
  nand_5 g16559(.A(new_n18907_1), .B(new_n18905), .Y(new_n18908));
  nand_5 g16560(.A(new_n18908), .B(new_n18904), .Y(new_n18909));
  nand_5 g16561(.A(new_n18909), .B(new_n18901_1), .Y(new_n18910));
  nand_5 g16562(.A(new_n18910), .B(new_n18900), .Y(new_n18911));
  nand_5 g16563(.A(new_n18911), .B(new_n18897), .Y(new_n18912));
  nand_5 g16564(.A(new_n18912), .B(new_n18896), .Y(new_n18913));
  nand_5 g16565(.A(new_n18913), .B(new_n18893), .Y(new_n18914));
  nand_5 g16566(.A(new_n18914), .B(new_n18892), .Y(new_n18915));
  nand_5 g16567(.A(new_n18915), .B(new_n18889), .Y(new_n18916));
  nand_5 g16568(.A(new_n18916), .B(new_n18888), .Y(new_n18917));
  nand_5 g16569(.A(new_n18917), .B(new_n18885), .Y(new_n18918));
  nand_5 g16570(.A(new_n18918), .B(new_n18884), .Y(new_n18919_1));
  xnor_4 g16571(.A(new_n18919_1), .B(new_n18881), .Y(n3932));
  nand_5 g16572(.A(new_n4262), .B(new_n4261), .Y(new_n18921));
  xnor_4 g16573(.A(new_n18921), .B(new_n4266_1), .Y(n3934));
  nand_5 g16574(.A(new_n4477), .B(new_n4475), .Y(new_n18923));
  xor_4  g16575(.A(new_n18923), .B(new_n2642), .Y(n3971));
  nand_5 g16576(.A(new_n7526), .B(new_n7519), .Y(new_n18925));
  or_5   g16577(.A(new_n18925), .B(n12161), .Y(new_n18926_1));
  nor_5  g16578(.A(new_n18926_1), .B(n18157), .Y(new_n18927));
  nand_5 g16579(.A(new_n18927), .B(new_n8306_1), .Y(new_n18928));
  xor_4  g16580(.A(new_n18928), .B(n8067), .Y(new_n18929));
  or_5   g16581(.A(new_n18929), .B(n26054), .Y(new_n18930));
  nand_5 g16582(.A(new_n18929), .B(n26054), .Y(new_n18931));
  xor_4  g16583(.A(new_n18927), .B(n20923), .Y(new_n18932));
  nand_5 g16584(.A(new_n18932), .B(new_n11713), .Y(new_n18933));
  or_5   g16585(.A(new_n18932), .B(new_n11713), .Y(new_n18934));
  xor_4  g16586(.A(new_n18926_1), .B(n18157), .Y(new_n18935));
  or_5   g16587(.A(new_n18935), .B(n8309), .Y(new_n18936));
  nand_5 g16588(.A(new_n18935), .B(n8309), .Y(new_n18937));
  nand_5 g16589(.A(new_n18925), .B(n12161), .Y(new_n18938));
  nand_5 g16590(.A(new_n18938), .B(new_n18926_1), .Y(new_n18939));
  nand_5 g16591(.A(new_n18939), .B(new_n11720), .Y(new_n18940_1));
  nor_5  g16592(.A(new_n18939), .B(new_n11720), .Y(new_n18941));
  not_8  g16593(.A(new_n18941), .Y(new_n18942));
  nand_5 g16594(.A(n8581), .B(n5026), .Y(new_n18943));
  and_5  g16595(.A(new_n18943), .B(new_n18925), .Y(new_n18944));
  or_5   g16596(.A(new_n18944), .B(n12593), .Y(new_n18945_1));
  nand_5 g16597(.A(new_n18944), .B(n12593), .Y(new_n18946));
  nand_5 g16598(.A(n13714), .B(n8581), .Y(new_n18947));
  nand_5 g16599(.A(new_n18947), .B(new_n18946), .Y(new_n18948));
  nand_5 g16600(.A(new_n18948), .B(new_n18945_1), .Y(new_n18949));
  nand_5 g16601(.A(new_n18949), .B(new_n18942), .Y(new_n18950));
  nand_5 g16602(.A(new_n18950), .B(new_n18940_1), .Y(new_n18951));
  nand_5 g16603(.A(new_n18951), .B(new_n18937), .Y(new_n18952));
  nand_5 g16604(.A(new_n18952), .B(new_n18936), .Y(new_n18953));
  nand_5 g16605(.A(new_n18953), .B(new_n18934), .Y(new_n18954));
  nand_5 g16606(.A(new_n18954), .B(new_n18933), .Y(new_n18955));
  nand_5 g16607(.A(new_n18955), .B(new_n18931), .Y(new_n18956));
  nand_5 g16608(.A(new_n18956), .B(new_n18930), .Y(new_n18957));
  nor_5  g16609(.A(new_n18928), .B(n8067), .Y(new_n18958));
  xor_4  g16610(.A(new_n18958), .B(new_n8300), .Y(new_n18959));
  or_5   g16611(.A(new_n18959), .B(n26318), .Y(new_n18960));
  nand_5 g16612(.A(new_n18959), .B(n26318), .Y(new_n18961));
  nand_5 g16613(.A(new_n18961), .B(new_n18960), .Y(new_n18962_1));
  xor_4  g16614(.A(new_n18962_1), .B(new_n18957), .Y(new_n18963));
  not_8  g16615(.A(new_n18963), .Y(new_n18964));
  nand_5 g16616(.A(new_n18964), .B(new_n6169), .Y(new_n18965));
  nand_5 g16617(.A(new_n18963), .B(n22554), .Y(new_n18966));
  nand_5 g16618(.A(new_n18931), .B(new_n18930), .Y(new_n18967));
  xor_4  g16619(.A(new_n18967), .B(new_n18955), .Y(new_n18968));
  not_8  g16620(.A(new_n18968), .Y(new_n18969));
  nand_5 g16621(.A(new_n18969), .B(new_n9241), .Y(new_n18970_1));
  nand_5 g16622(.A(new_n18968), .B(n20429), .Y(new_n18971));
  nand_5 g16623(.A(new_n18934), .B(new_n18933), .Y(new_n18972));
  xor_4  g16624(.A(new_n18972), .B(new_n18953), .Y(new_n18973));
  not_8  g16625(.A(new_n18973), .Y(new_n18974));
  nand_5 g16626(.A(new_n18974), .B(new_n6170), .Y(new_n18975));
  nand_5 g16627(.A(new_n18973), .B(n3909), .Y(new_n18976));
  nand_5 g16628(.A(new_n18937), .B(new_n18936), .Y(new_n18977_1));
  xor_4  g16629(.A(new_n18977_1), .B(new_n18951), .Y(new_n18978));
  not_8  g16630(.A(new_n18978), .Y(new_n18979));
  nand_5 g16631(.A(new_n18979), .B(new_n9247), .Y(new_n18980));
  nand_5 g16632(.A(new_n18978), .B(n23974), .Y(new_n18981));
  nand_5 g16633(.A(new_n18942), .B(new_n18940_1), .Y(new_n18982_1));
  xor_4  g16634(.A(new_n18982_1), .B(new_n18949), .Y(new_n18983));
  not_8  g16635(.A(new_n18983), .Y(new_n18984));
  nand_5 g16636(.A(new_n18984), .B(new_n9251_1), .Y(new_n18985));
  nand_5 g16637(.A(new_n18983), .B(n2146), .Y(new_n18986));
  nand_5 g16638(.A(new_n18946), .B(new_n18945_1), .Y(new_n18987));
  not_8  g16639(.A(new_n18987), .Y(new_n18988));
  xor_4  g16640(.A(new_n18988), .B(new_n18947), .Y(new_n18989));
  nand_5 g16641(.A(new_n18989), .B(new_n6171_1), .Y(new_n18990));
  or_5   g16642(.A(new_n18989), .B(new_n6171_1), .Y(new_n18991));
  nand_5 g16643(.A(new_n10138), .B(new_n7526), .Y(new_n18992));
  and_5  g16644(.A(new_n18992), .B(new_n18947), .Y(new_n18993));
  nand_5 g16645(.A(new_n18993), .B(n583), .Y(new_n18994));
  nand_5 g16646(.A(new_n18994), .B(new_n18991), .Y(new_n18995));
  nand_5 g16647(.A(new_n18995), .B(new_n18990), .Y(new_n18996));
  nand_5 g16648(.A(new_n18996), .B(new_n18986), .Y(new_n18997));
  nand_5 g16649(.A(new_n18997), .B(new_n18985), .Y(new_n18998));
  nand_5 g16650(.A(new_n18998), .B(new_n18981), .Y(new_n18999_1));
  nand_5 g16651(.A(new_n18999_1), .B(new_n18980), .Y(new_n19000));
  nand_5 g16652(.A(new_n19000), .B(new_n18976), .Y(new_n19001));
  nand_5 g16653(.A(new_n19001), .B(new_n18975), .Y(new_n19002));
  nand_5 g16654(.A(new_n19002), .B(new_n18971), .Y(new_n19003));
  nand_5 g16655(.A(new_n19003), .B(new_n18970_1), .Y(new_n19004));
  nand_5 g16656(.A(new_n19004), .B(new_n18966), .Y(new_n19005_1));
  nand_5 g16657(.A(new_n19005_1), .B(new_n18965), .Y(new_n19006));
  nand_5 g16658(.A(new_n18961), .B(new_n18957), .Y(new_n19007));
  nand_5 g16659(.A(new_n19007), .B(new_n18960), .Y(new_n19008));
  nand_5 g16660(.A(new_n18958), .B(new_n8300), .Y(new_n19009));
  xor_4  g16661(.A(new_n19009), .B(n25240), .Y(new_n19010));
  or_5   g16662(.A(new_n19010), .B(n3710), .Y(new_n19011));
  nand_5 g16663(.A(new_n19010), .B(n3710), .Y(new_n19012));
  nand_5 g16664(.A(new_n19012), .B(new_n19011), .Y(new_n19013));
  xor_4  g16665(.A(new_n19013), .B(new_n19008), .Y(new_n19014));
  not_8  g16666(.A(new_n19014), .Y(new_n19015));
  nand_5 g16667(.A(new_n19015), .B(new_n9235), .Y(new_n19016));
  nand_5 g16668(.A(new_n19014), .B(n23913), .Y(new_n19017));
  nand_5 g16669(.A(new_n19017), .B(new_n19016), .Y(new_n19018));
  xor_4  g16670(.A(new_n19018), .B(new_n19006), .Y(new_n19019));
  or_5   g16671(.A(new_n19019), .B(new_n9366), .Y(new_n19020));
  nand_5 g16672(.A(new_n19019), .B(new_n9366), .Y(new_n19021));
  nand_5 g16673(.A(new_n18965), .B(new_n18966), .Y(new_n19022));
  xor_4  g16674(.A(new_n19022), .B(new_n19004), .Y(new_n19023));
  or_5   g16675(.A(new_n19023), .B(new_n9372_1), .Y(new_n19024));
  nand_5 g16676(.A(new_n19023), .B(new_n9372_1), .Y(new_n19025));
  nand_5 g16677(.A(new_n18970_1), .B(new_n18971), .Y(new_n19026));
  xor_4  g16678(.A(new_n19026), .B(new_n19002), .Y(new_n19027));
  or_5   g16679(.A(new_n19027), .B(new_n9378), .Y(new_n19028));
  nand_5 g16680(.A(new_n19027), .B(new_n9378), .Y(new_n19029));
  nand_5 g16681(.A(new_n18975), .B(new_n18976), .Y(new_n19030));
  xor_4  g16682(.A(new_n19030), .B(new_n19000), .Y(new_n19031));
  or_5   g16683(.A(new_n19031), .B(new_n9384), .Y(new_n19032));
  nand_5 g16684(.A(new_n19031), .B(new_n9384), .Y(new_n19033_1));
  nand_5 g16685(.A(new_n18980), .B(new_n18981), .Y(new_n19034));
  xor_4  g16686(.A(new_n19034), .B(new_n18998), .Y(new_n19035));
  or_5   g16687(.A(new_n19035), .B(new_n9390), .Y(new_n19036));
  nand_5 g16688(.A(new_n19035), .B(new_n9390), .Y(new_n19037));
  nand_5 g16689(.A(new_n18985), .B(new_n18986), .Y(new_n19038));
  xor_4  g16690(.A(new_n19038), .B(new_n18996), .Y(new_n19039));
  or_5   g16691(.A(new_n19039), .B(new_n9396_1), .Y(new_n19040));
  nand_5 g16692(.A(new_n19039), .B(new_n9396_1), .Y(new_n19041));
  nand_5 g16693(.A(new_n18990), .B(new_n18991), .Y(new_n19042_1));
  xor_4  g16694(.A(new_n19042_1), .B(new_n18994), .Y(new_n19043));
  or_5   g16695(.A(new_n19043), .B(new_n9403_1), .Y(new_n19044_1));
  nand_5 g16696(.A(new_n19043), .B(new_n9403_1), .Y(new_n19045));
  xor_4  g16697(.A(new_n18993), .B(n583), .Y(new_n19046));
  nand_5 g16698(.A(new_n19046), .B(new_n2618), .Y(new_n19047));
  nand_5 g16699(.A(new_n19047), .B(new_n19045), .Y(new_n19048));
  nand_5 g16700(.A(new_n19048), .B(new_n19044_1), .Y(new_n19049));
  nand_5 g16701(.A(new_n19049), .B(new_n19041), .Y(new_n19050));
  nand_5 g16702(.A(new_n19050), .B(new_n19040), .Y(new_n19051));
  nand_5 g16703(.A(new_n19051), .B(new_n19037), .Y(new_n19052));
  nand_5 g16704(.A(new_n19052), .B(new_n19036), .Y(new_n19053));
  nand_5 g16705(.A(new_n19053), .B(new_n19033_1), .Y(new_n19054));
  nand_5 g16706(.A(new_n19054), .B(new_n19032), .Y(new_n19055));
  nand_5 g16707(.A(new_n19055), .B(new_n19029), .Y(new_n19056));
  nand_5 g16708(.A(new_n19056), .B(new_n19028), .Y(new_n19057));
  nand_5 g16709(.A(new_n19057), .B(new_n19025), .Y(new_n19058));
  nand_5 g16710(.A(new_n19058), .B(new_n19024), .Y(new_n19059));
  nand_5 g16711(.A(new_n19059), .B(new_n19021), .Y(new_n19060));
  nand_5 g16712(.A(new_n19060), .B(new_n19020), .Y(new_n19061));
  nand_5 g16713(.A(new_n19017), .B(new_n19006), .Y(new_n19062));
  nand_5 g16714(.A(new_n19062), .B(new_n19016), .Y(new_n19063));
  nor_5  g16715(.A(new_n19009), .B(n25240), .Y(new_n19064));
  xor_4  g16716(.A(new_n19064), .B(new_n8294), .Y(new_n19065));
  nand_5 g16717(.A(new_n19065), .B(n15077), .Y(new_n19066));
  or_5   g16718(.A(new_n19065), .B(n15077), .Y(new_n19067));
  nand_5 g16719(.A(new_n19067), .B(new_n19066), .Y(new_n19068));
  nand_5 g16720(.A(new_n19012), .B(new_n19008), .Y(new_n19069));
  nand_5 g16721(.A(new_n19069), .B(new_n19011), .Y(new_n19070));
  xor_4  g16722(.A(new_n19070), .B(new_n19068), .Y(new_n19071));
  not_8  g16723(.A(new_n19071), .Y(new_n19072));
  nand_5 g16724(.A(new_n19072), .B(new_n6168), .Y(new_n19073));
  nand_5 g16725(.A(new_n19071), .B(n26797), .Y(new_n19074));
  nand_5 g16726(.A(new_n19074), .B(new_n19073), .Y(new_n19075));
  xnor_4 g16727(.A(new_n19075), .B(new_n19063), .Y(new_n19076));
  not_8  g16728(.A(new_n19076), .Y(new_n19077));
  nand_5 g16729(.A(new_n19077), .B(new_n9360), .Y(new_n19078));
  not_8  g16730(.A(new_n19078), .Y(new_n19079));
  nor_5  g16731(.A(new_n19077), .B(new_n9360), .Y(new_n19080));
  or_5   g16732(.A(new_n19080), .B(new_n19079), .Y(new_n19081_1));
  xor_4  g16733(.A(new_n19081_1), .B(new_n19061), .Y(n3983));
  not_8  g16734(.A(new_n7590), .Y(new_n19083));
  nand_5 g16735(.A(n13714), .B(n583), .Y(new_n19084));
  nand_5 g16736(.A(new_n10138), .B(new_n2620), .Y(new_n19085));
  nand_5 g16737(.A(new_n19085), .B(new_n19084), .Y(new_n19086));
  xor_4  g16738(.A(new_n19086), .B(new_n6339_1), .Y(new_n19087));
  nor_5  g16739(.A(new_n19087), .B(new_n19083), .Y(new_n19088));
  not_8  g16740(.A(new_n19088), .Y(new_n19089));
  nor_5  g16741(.A(new_n19086), .B(new_n6339_1), .Y(new_n19090));
  not_8  g16742(.A(new_n19084), .Y(new_n19091));
  nand_5 g16743(.A(new_n6171_1), .B(new_n11723), .Y(new_n19092));
  nand_5 g16744(.A(n22173), .B(n12593), .Y(new_n19093));
  nand_5 g16745(.A(new_n19093), .B(new_n19092), .Y(new_n19094));
  xor_4  g16746(.A(new_n19094), .B(new_n19091), .Y(new_n19095));
  or_5   g16747(.A(new_n19095), .B(new_n10338), .Y(new_n19096));
  nand_5 g16748(.A(new_n19095), .B(new_n10338), .Y(new_n19097));
  nand_5 g16749(.A(new_n19097), .B(new_n19096), .Y(new_n19098));
  xnor_4 g16750(.A(new_n19098), .B(new_n19090), .Y(new_n19099));
  nand_5 g16751(.A(new_n19099), .B(new_n19089), .Y(new_n19100));
  nor_5  g16752(.A(new_n19099), .B(new_n19089), .Y(new_n19101));
  not_8  g16753(.A(new_n19101), .Y(new_n19102));
  nand_5 g16754(.A(new_n19102), .B(new_n19100), .Y(new_n19103));
  xor_4  g16755(.A(new_n19103), .B(new_n7582), .Y(n4000));
  nand_5 g16756(.A(n24278), .B(new_n7735), .Y(new_n19105));
  nand_5 g16757(.A(new_n2350), .B(n15539), .Y(new_n19106));
  nand_5 g16758(.A(n24618), .B(new_n7738), .Y(new_n19107_1));
  nand_5 g16759(.A(new_n2354), .B(n8052), .Y(new_n19108));
  nand_5 g16760(.A(new_n12965), .B(new_n12963), .Y(new_n19109));
  nand_5 g16761(.A(new_n19109), .B(new_n12964), .Y(new_n19110));
  nand_5 g16762(.A(new_n19110), .B(new_n19108), .Y(new_n19111));
  nand_5 g16763(.A(new_n19111), .B(new_n19107_1), .Y(new_n19112));
  nand_5 g16764(.A(new_n19112), .B(new_n19106), .Y(new_n19113));
  nand_5 g16765(.A(new_n19113), .B(new_n19105), .Y(new_n19114));
  nand_5 g16766(.A(new_n7732), .B(n4812), .Y(new_n19115));
  nand_5 g16767(.A(n19228), .B(new_n2371), .Y(new_n19116_1));
  nand_5 g16768(.A(new_n19116_1), .B(new_n19115), .Y(new_n19117));
  xor_4  g16769(.A(new_n19117), .B(new_n19114), .Y(new_n19118));
  or_5   g16770(.A(new_n19118), .B(new_n8514), .Y(new_n19119));
  nand_5 g16771(.A(new_n19118), .B(new_n8514), .Y(new_n19120));
  nand_5 g16772(.A(new_n19106), .B(new_n19105), .Y(new_n19121));
  xor_4  g16773(.A(new_n19121), .B(new_n19112), .Y(new_n19122));
  or_5   g16774(.A(new_n19122), .B(new_n8521), .Y(new_n19123));
  nand_5 g16775(.A(new_n19122), .B(new_n8521), .Y(new_n19124));
  nand_5 g16776(.A(new_n19108), .B(new_n19107_1), .Y(new_n19125_1));
  xor_4  g16777(.A(new_n19125_1), .B(new_n19110), .Y(new_n19126));
  or_5   g16778(.A(new_n19126), .B(new_n8528), .Y(new_n19127));
  nand_5 g16779(.A(new_n19126), .B(new_n8528), .Y(new_n19128));
  not_8  g16780(.A(new_n8543), .Y(new_n19129));
  nand_5 g16781(.A(new_n12970), .B(new_n19129), .Y(new_n19130));
  nand_5 g16782(.A(new_n19130), .B(new_n12968), .Y(new_n19131));
  nand_5 g16783(.A(new_n19131), .B(new_n19128), .Y(new_n19132));
  nand_5 g16784(.A(new_n19132), .B(new_n19127), .Y(new_n19133));
  nand_5 g16785(.A(new_n19133), .B(new_n19124), .Y(new_n19134));
  nand_5 g16786(.A(new_n19134), .B(new_n19123), .Y(new_n19135));
  nand_5 g16787(.A(new_n19135), .B(new_n19120), .Y(new_n19136));
  nand_5 g16788(.A(new_n19136), .B(new_n19119), .Y(new_n19137));
  nand_5 g16789(.A(new_n19116_1), .B(new_n19114), .Y(new_n19138));
  nand_5 g16790(.A(new_n19138), .B(new_n19115), .Y(new_n19139));
  nand_5 g16791(.A(n26823), .B(new_n7729), .Y(new_n19140));
  nand_5 g16792(.A(new_n2468), .B(n20179), .Y(new_n19141_1));
  nand_5 g16793(.A(new_n19141_1), .B(new_n19140), .Y(new_n19142));
  xnor_4 g16794(.A(new_n19142), .B(new_n19139), .Y(new_n19143));
  nand_5 g16795(.A(new_n19143), .B(new_n8506), .Y(new_n19144_1));
  not_8  g16796(.A(new_n19144_1), .Y(new_n19145));
  nor_5  g16797(.A(new_n19143), .B(new_n8506), .Y(new_n19146));
  nor_5  g16798(.A(new_n19146), .B(new_n19145), .Y(new_n19147));
  xor_4  g16799(.A(new_n19147), .B(new_n19137), .Y(n4010));
  nand_5 g16800(.A(n11220), .B(new_n13565), .Y(new_n19149));
  nand_5 g16801(.A(new_n11623), .B(n2160), .Y(new_n19150));
  nand_5 g16802(.A(new_n19150), .B(new_n19149), .Y(new_n19151));
  nand_5 g16803(.A(new_n3276), .B(n10763), .Y(new_n19152));
  nand_5 g16804(.A(n22379), .B(new_n3287), .Y(new_n19153));
  nand_5 g16805(.A(n7437), .B(new_n3030_1), .Y(new_n19154));
  nand_5 g16806(.A(new_n3185), .B(n1662), .Y(new_n19155));
  nand_5 g16807(.A(n20700), .B(new_n2997), .Y(new_n19156));
  nand_5 g16808(.A(new_n3067_1), .B(n12875), .Y(new_n19157));
  nand_5 g16809(.A(new_n16832), .B(new_n16829), .Y(new_n19158));
  nand_5 g16810(.A(new_n19158), .B(new_n16831), .Y(new_n19159));
  nand_5 g16811(.A(new_n19159), .B(new_n19157), .Y(new_n19160));
  nand_5 g16812(.A(new_n19160), .B(new_n19156), .Y(new_n19161));
  nand_5 g16813(.A(new_n19161), .B(new_n19155), .Y(new_n19162));
  nand_5 g16814(.A(new_n19162), .B(new_n19154), .Y(new_n19163_1));
  nand_5 g16815(.A(new_n19163_1), .B(new_n19153), .Y(new_n19164_1));
  nand_5 g16816(.A(new_n19164_1), .B(new_n19152), .Y(new_n19165));
  xnor_4 g16817(.A(new_n19165), .B(new_n19151), .Y(new_n19166));
  nand_5 g16818(.A(new_n19166), .B(new_n16958), .Y(new_n19167));
  or_5   g16819(.A(new_n19166), .B(new_n16958), .Y(new_n19168));
  nand_5 g16820(.A(new_n19168), .B(new_n19167), .Y(new_n19169));
  nand_5 g16821(.A(new_n19153), .B(new_n19152), .Y(new_n19170));
  xor_4  g16822(.A(new_n19170), .B(new_n19163_1), .Y(new_n19171));
  nand_5 g16823(.A(new_n19171), .B(new_n16964), .Y(new_n19172));
  or_5   g16824(.A(new_n19171), .B(new_n16964), .Y(new_n19173));
  nand_5 g16825(.A(new_n19155), .B(new_n19154), .Y(new_n19174_1));
  xor_4  g16826(.A(new_n19174_1), .B(new_n19161), .Y(new_n19175));
  nand_5 g16827(.A(new_n19175), .B(new_n16968_1), .Y(new_n19176_1));
  or_5   g16828(.A(new_n19175), .B(new_n16968_1), .Y(new_n19177));
  nand_5 g16829(.A(new_n19157), .B(new_n19156), .Y(new_n19178));
  xor_4  g16830(.A(new_n19178), .B(new_n19159), .Y(new_n19179));
  nand_5 g16831(.A(new_n19179), .B(new_n16979), .Y(new_n19180));
  or_5   g16832(.A(new_n19179), .B(new_n16979), .Y(new_n19181));
  nand_5 g16833(.A(new_n16836), .B(new_n16813), .Y(new_n19182));
  nand_5 g16834(.A(new_n19182), .B(new_n16835), .Y(new_n19183));
  nand_5 g16835(.A(new_n19183), .B(new_n19181), .Y(new_n19184));
  nand_5 g16836(.A(new_n19184), .B(new_n19180), .Y(new_n19185));
  nand_5 g16837(.A(new_n19185), .B(new_n19177), .Y(new_n19186));
  nand_5 g16838(.A(new_n19186), .B(new_n19176_1), .Y(new_n19187));
  nand_5 g16839(.A(new_n19187), .B(new_n19173), .Y(new_n19188));
  nand_5 g16840(.A(new_n19188), .B(new_n19172), .Y(new_n19189));
  xor_4  g16841(.A(new_n19189), .B(new_n19169), .Y(n4014));
  nand_5 g16842(.A(new_n4308), .B(new_n4292), .Y(new_n19191));
  nand_5 g16843(.A(new_n19191), .B(new_n4307), .Y(new_n19192));
  nand_5 g16844(.A(new_n4304), .B(new_n4295), .Y(new_n19193));
  nand_5 g16845(.A(new_n19193), .B(new_n4303), .Y(new_n19194));
  nand_5 g16846(.A(new_n16125), .B(new_n5588), .Y(new_n19195));
  nand_5 g16847(.A(new_n16124), .B(n26224), .Y(new_n19196_1));
  nand_5 g16848(.A(new_n19196_1), .B(new_n19195), .Y(new_n19197));
  xor_4  g16849(.A(new_n19197), .B(new_n19194), .Y(new_n19198));
  not_8  g16850(.A(new_n19198), .Y(new_n19199));
  nand_5 g16851(.A(new_n19199), .B(new_n5375), .Y(new_n19200));
  nand_5 g16852(.A(new_n19198), .B(n20409), .Y(new_n19201));
  nand_5 g16853(.A(new_n19201), .B(new_n19200), .Y(new_n19202_1));
  xor_4  g16854(.A(new_n19202_1), .B(new_n19192), .Y(new_n19203));
  nand_5 g16855(.A(new_n19203), .B(new_n13678), .Y(new_n19204));
  or_5   g16856(.A(new_n19203), .B(new_n13678), .Y(new_n19205));
  nand_5 g16857(.A(new_n4311), .B(new_n4276), .Y(new_n19206));
  nand_5 g16858(.A(new_n19206), .B(new_n4312), .Y(new_n19207));
  nand_5 g16859(.A(new_n19207), .B(new_n19205), .Y(new_n19208));
  nand_5 g16860(.A(new_n19208), .B(new_n19204), .Y(new_n19209));
  nand_5 g16861(.A(new_n19201), .B(new_n19192), .Y(new_n19210));
  nand_5 g16862(.A(new_n19210), .B(new_n19200), .Y(new_n19211));
  nand_5 g16863(.A(new_n19196_1), .B(new_n19194), .Y(new_n19212));
  nand_5 g16864(.A(new_n19212), .B(new_n19195), .Y(new_n19213));
  not_8  g16865(.A(new_n19213), .Y(new_n19214));
  nand_5 g16866(.A(new_n16121), .B(new_n5363), .Y(new_n19215));
  nand_5 g16867(.A(new_n16120), .B(n18496), .Y(new_n19216));
  nand_5 g16868(.A(new_n19216), .B(new_n19215), .Y(new_n19217));
  xor_4  g16869(.A(new_n19217), .B(new_n19214), .Y(new_n19218));
  nand_5 g16870(.A(new_n19218), .B(new_n5370), .Y(new_n19219));
  or_5   g16871(.A(new_n19218), .B(new_n5370), .Y(new_n19220_1));
  nand_5 g16872(.A(new_n19220_1), .B(new_n19219), .Y(new_n19221_1));
  xor_4  g16873(.A(new_n19221_1), .B(new_n19211), .Y(new_n19222));
  or_5   g16874(.A(new_n19222), .B(new_n13671), .Y(new_n19223_1));
  nand_5 g16875(.A(new_n19222), .B(new_n13671), .Y(new_n19224_1));
  nand_5 g16876(.A(new_n19224_1), .B(new_n19223_1), .Y(new_n19225));
  xnor_4 g16877(.A(new_n19225), .B(new_n19209), .Y(n4071));
  nand_5 g16878(.A(new_n14776), .B(new_n14775), .Y(new_n19227));
  xor_4  g16879(.A(new_n19227), .B(new_n14782), .Y(n4088));
  nor_5  g16880(.A(new_n14919), .B(new_n14915), .Y(new_n19229));
  nor_5  g16881(.A(new_n6157), .B(n7593), .Y(new_n19230));
  not_8  g16882(.A(new_n19230), .Y(new_n19231));
  nand_5 g16883(.A(new_n14914), .B(new_n19231), .Y(new_n19232));
  nor_5  g16884(.A(new_n19232), .B(new_n19229), .Y(new_n19233_1));
  not_8  g16885(.A(new_n19233_1), .Y(new_n19234_1));
  nand_5 g16886(.A(new_n19234_1), .B(new_n18585), .Y(new_n19235));
  not_8  g16887(.A(new_n19235), .Y(new_n19236));
  nand_5 g16888(.A(new_n19233_1), .B(new_n18587), .Y(new_n19237));
  not_8  g16889(.A(new_n19237), .Y(new_n19238));
  nor_5  g16890(.A(new_n14926), .B(new_n14922), .Y(new_n19239));
  nor_5  g16891(.A(new_n19239), .B(new_n14923), .Y(new_n19240));
  nor_5  g16892(.A(new_n19240), .B(new_n19238), .Y(new_n19241));
  nor_5  g16893(.A(new_n19241), .B(new_n19236), .Y(new_n19242));
  nand_5 g16894(.A(new_n18584_1), .B(new_n18581), .Y(new_n19243));
  nand_5 g16895(.A(new_n19243), .B(new_n18580), .Y(new_n19244_1));
  not_8  g16896(.A(new_n19244_1), .Y(new_n19245));
  nor_5  g16897(.A(new_n19245), .B(new_n19234_1), .Y(new_n19246));
  nor_5  g16898(.A(new_n19246), .B(new_n19242), .Y(new_n19247));
  nor_5  g16899(.A(new_n19244_1), .B(new_n19233_1), .Y(new_n19248));
  nor_5  g16900(.A(new_n19248), .B(new_n19241), .Y(new_n19249));
  nor_5  g16901(.A(new_n19249), .B(new_n19247), .Y(n4089));
  nand_5 g16902(.A(new_n9932), .B(new_n9925), .Y(new_n19251));
  nand_5 g16903(.A(new_n19251), .B(new_n9931), .Y(new_n19252));
  not_8  g16904(.A(new_n19252), .Y(new_n19253));
  nand_5 g16905(.A(new_n13919), .B(new_n3626), .Y(new_n19254));
  nand_5 g16906(.A(new_n13918), .B(n25738), .Y(new_n19255));
  nand_5 g16907(.A(new_n19255), .B(new_n19254), .Y(new_n19256));
  xor_4  g16908(.A(new_n19256), .B(new_n19253), .Y(new_n19257));
  nand_5 g16909(.A(new_n19257), .B(new_n7819), .Y(new_n19258));
  or_5   g16910(.A(new_n19257), .B(new_n7819), .Y(new_n19259));
  nand_5 g16911(.A(new_n9936), .B(new_n9923), .Y(new_n19260));
  nand_5 g16912(.A(new_n19260), .B(new_n9935), .Y(new_n19261));
  nand_5 g16913(.A(new_n19261), .B(new_n19259), .Y(new_n19262));
  nand_5 g16914(.A(new_n19262), .B(new_n19258), .Y(new_n19263));
  nand_5 g16915(.A(new_n19255), .B(new_n19252), .Y(new_n19264));
  nand_5 g16916(.A(new_n19264), .B(new_n19254), .Y(new_n19265));
  not_8  g16917(.A(new_n19265), .Y(new_n19266));
  nand_5 g16918(.A(new_n13986), .B(new_n5889), .Y(new_n19267));
  nand_5 g16919(.A(new_n13985), .B(n5302), .Y(new_n19268));
  nand_5 g16920(.A(new_n19268), .B(new_n19267), .Y(new_n19269));
  xor_4  g16921(.A(new_n19269), .B(new_n19266), .Y(new_n19270_1));
  nand_5 g16922(.A(new_n19270_1), .B(new_n7838), .Y(new_n19271));
  or_5   g16923(.A(new_n19270_1), .B(new_n7838), .Y(new_n19272));
  nand_5 g16924(.A(new_n19272), .B(new_n19271), .Y(new_n19273));
  xor_4  g16925(.A(new_n19273), .B(new_n19263), .Y(new_n19274));
  nand_5 g16926(.A(new_n2472), .B(new_n6399), .Y(new_n19275));
  nand_5 g16927(.A(new_n2471), .B(n17959), .Y(new_n19276));
  nand_5 g16928(.A(new_n7713), .B(new_n7710), .Y(new_n19277));
  nand_5 g16929(.A(new_n19277), .B(new_n7712), .Y(new_n19278));
  nand_5 g16930(.A(new_n19278), .B(new_n19276), .Y(new_n19279));
  nand_5 g16931(.A(new_n19279), .B(new_n19275), .Y(new_n19280));
  nand_5 g16932(.A(new_n2590), .B(new_n6396), .Y(new_n19281));
  nand_5 g16933(.A(new_n2589), .B(n23200), .Y(new_n19282_1));
  nand_5 g16934(.A(new_n19282_1), .B(new_n19281), .Y(new_n19283));
  xor_4  g16935(.A(new_n19283), .B(new_n19280), .Y(new_n19284));
  or_5   g16936(.A(new_n19284), .B(new_n19274), .Y(new_n19285));
  nand_5 g16937(.A(new_n19284), .B(new_n19274), .Y(new_n19286));
  nand_5 g16938(.A(new_n19275), .B(new_n19276), .Y(new_n19287));
  xor_4  g16939(.A(new_n19287), .B(new_n19278), .Y(new_n19288));
  nand_5 g16940(.A(new_n19258), .B(new_n19259), .Y(new_n19289));
  xor_4  g16941(.A(new_n19289), .B(new_n19261), .Y(new_n19290));
  or_5   g16942(.A(new_n19290), .B(new_n19288), .Y(new_n19291));
  nand_5 g16943(.A(new_n19290), .B(new_n19288), .Y(new_n19292));
  nand_5 g16944(.A(new_n9940), .B(new_n9920), .Y(new_n19293));
  nand_5 g16945(.A(new_n19293), .B(new_n9939), .Y(new_n19294));
  nand_5 g16946(.A(new_n19294), .B(new_n19292), .Y(new_n19295));
  nand_5 g16947(.A(new_n19295), .B(new_n19291), .Y(new_n19296));
  nand_5 g16948(.A(new_n19296), .B(new_n19286), .Y(new_n19297));
  nand_5 g16949(.A(new_n19297), .B(new_n19285), .Y(new_n19298));
  nand_5 g16950(.A(new_n19272), .B(new_n19263), .Y(new_n19299));
  nand_5 g16951(.A(new_n19299), .B(new_n19271), .Y(new_n19300));
  nand_5 g16952(.A(new_n19268), .B(new_n19265), .Y(new_n19301));
  nand_5 g16953(.A(new_n19301), .B(new_n19267), .Y(new_n19302));
  not_8  g16954(.A(new_n19302), .Y(new_n19303));
  nor_5  g16955(.A(new_n13983), .B(n2289), .Y(new_n19304));
  not_8  g16956(.A(new_n19304), .Y(new_n19305));
  nand_5 g16957(.A(new_n13983), .B(n2289), .Y(new_n19306));
  and_5  g16958(.A(new_n19306), .B(new_n19305), .Y(new_n19307));
  not_8  g16959(.A(new_n19307), .Y(new_n19308));
  nand_5 g16960(.A(new_n19308), .B(new_n3545), .Y(new_n19309));
  nand_5 g16961(.A(new_n19307), .B(n3228), .Y(new_n19310));
  nand_5 g16962(.A(new_n19310), .B(new_n19309), .Y(new_n19311));
  xor_4  g16963(.A(new_n19311), .B(new_n19303), .Y(new_n19312));
  nand_5 g16964(.A(new_n19312), .B(new_n7882), .Y(new_n19313));
  or_5   g16965(.A(new_n19312), .B(new_n7882), .Y(new_n19314_1));
  nand_5 g16966(.A(new_n19314_1), .B(new_n19313), .Y(new_n19315_1));
  xor_4  g16967(.A(new_n19315_1), .B(new_n19300), .Y(new_n19316));
  nand_5 g16968(.A(new_n19282_1), .B(new_n19280), .Y(new_n19317));
  nand_5 g16969(.A(new_n19317), .B(new_n19281), .Y(new_n19318));
  not_8  g16970(.A(new_n19318), .Y(new_n19319));
  nand_5 g16971(.A(new_n8632), .B(new_n6392), .Y(new_n19320));
  or_5   g16972(.A(new_n8632), .B(new_n6392), .Y(new_n19321));
  nand_5 g16973(.A(new_n19321), .B(new_n19320), .Y(new_n19322));
  xor_4  g16974(.A(new_n19322), .B(new_n19319), .Y(new_n19323_1));
  not_8  g16975(.A(new_n19323_1), .Y(new_n19324));
  or_5   g16976(.A(new_n19324), .B(new_n19316), .Y(new_n19325));
  nand_5 g16977(.A(new_n19324), .B(new_n19316), .Y(new_n19326));
  nand_5 g16978(.A(new_n19326), .B(new_n19325), .Y(new_n19327_1));
  xor_4  g16979(.A(new_n19327_1), .B(new_n19298), .Y(n4103));
  xor_4  g16980(.A(new_n16868), .B(new_n14428), .Y(new_n19329));
  nand_5 g16981(.A(new_n16874), .B(new_n14430), .Y(new_n19330));
  nand_5 g16982(.A(new_n16875), .B(new_n14507), .Y(new_n19331));
  or_5   g16983(.A(new_n16879), .B(new_n14443), .Y(new_n19332));
  nand_5 g16984(.A(new_n16879), .B(new_n14443), .Y(new_n19333_1));
  or_5   g16985(.A(new_n16884), .B(new_n14448), .Y(new_n19334));
  nand_5 g16986(.A(new_n16884), .B(new_n14448), .Y(new_n19335));
  or_5   g16987(.A(new_n16889), .B(new_n14453), .Y(new_n19336));
  nand_5 g16988(.A(new_n16889), .B(new_n14453), .Y(new_n19337));
  or_5   g16989(.A(new_n16823), .B(new_n14458), .Y(new_n19338));
  nand_5 g16990(.A(new_n16823), .B(new_n14458), .Y(new_n19339));
  or_5   g16991(.A(new_n14463), .B(new_n4788), .Y(new_n19340));
  nand_5 g16992(.A(new_n14463), .B(new_n4788), .Y(new_n19341));
  or_5   g16993(.A(new_n14468), .B(new_n4716), .Y(new_n19342));
  nand_5 g16994(.A(new_n14468), .B(new_n4716), .Y(new_n19343));
  nand_5 g16995(.A(new_n14473), .B(new_n4669), .Y(new_n19344));
  nor_5  g16996(.A(new_n14473), .B(new_n4669), .Y(new_n19345));
  not_8  g16997(.A(new_n19345), .Y(new_n19346));
  nand_5 g16998(.A(new_n14479), .B(new_n4692), .Y(new_n19347));
  nand_5 g16999(.A(new_n14478), .B(new_n4747_1), .Y(new_n19348_1));
  nand_5 g17000(.A(new_n14486), .B(new_n4699), .Y(new_n19349));
  not_8  g17001(.A(new_n19349), .Y(new_n19350));
  nand_5 g17002(.A(new_n19350), .B(new_n19348_1), .Y(new_n19351));
  nand_5 g17003(.A(new_n19351), .B(new_n19347), .Y(new_n19352));
  nand_5 g17004(.A(new_n19352), .B(new_n19346), .Y(new_n19353));
  nand_5 g17005(.A(new_n19353), .B(new_n19344), .Y(new_n19354_1));
  not_8  g17006(.A(new_n19354_1), .Y(new_n19355));
  nand_5 g17007(.A(new_n19355), .B(new_n19343), .Y(new_n19356));
  nand_5 g17008(.A(new_n19356), .B(new_n19342), .Y(new_n19357_1));
  nand_5 g17009(.A(new_n19357_1), .B(new_n19341), .Y(new_n19358));
  nand_5 g17010(.A(new_n19358), .B(new_n19340), .Y(new_n19359));
  nand_5 g17011(.A(new_n19359), .B(new_n19339), .Y(new_n19360));
  nand_5 g17012(.A(new_n19360), .B(new_n19338), .Y(new_n19361_1));
  nand_5 g17013(.A(new_n19361_1), .B(new_n19337), .Y(new_n19362));
  nand_5 g17014(.A(new_n19362), .B(new_n19336), .Y(new_n19363));
  nand_5 g17015(.A(new_n19363), .B(new_n19335), .Y(new_n19364));
  nand_5 g17016(.A(new_n19364), .B(new_n19334), .Y(new_n19365));
  nand_5 g17017(.A(new_n19365), .B(new_n19333_1), .Y(new_n19366));
  nand_5 g17018(.A(new_n19366), .B(new_n19332), .Y(new_n19367_1));
  nand_5 g17019(.A(new_n19367_1), .B(new_n19331), .Y(new_n19368));
  nand_5 g17020(.A(new_n19368), .B(new_n19330), .Y(new_n19369));
  not_8  g17021(.A(new_n19369), .Y(new_n19370));
  nand_5 g17022(.A(new_n19370), .B(new_n19329), .Y(new_n19371));
  not_8  g17023(.A(new_n19371), .Y(new_n19372));
  nor_5  g17024(.A(new_n19370), .B(new_n19329), .Y(new_n19373));
  or_5   g17025(.A(new_n19373), .B(new_n19372), .Y(new_n19374));
  nand_5 g17026(.A(new_n6711), .B(new_n6663), .Y(new_n19375));
  not_8  g17027(.A(new_n19375), .Y(new_n19376));
  nand_5 g17028(.A(new_n6715), .B(new_n6666), .Y(new_n19377));
  nand_5 g17029(.A(new_n6714), .B(n4085), .Y(new_n19378));
  nand_5 g17030(.A(new_n6722), .B(new_n6669_1), .Y(new_n19379));
  nand_5 g17031(.A(new_n6721), .B(n26725), .Y(new_n19380));
  nand_5 g17032(.A(new_n6729_1), .B(new_n6672), .Y(new_n19381));
  nand_5 g17033(.A(new_n6728), .B(n11980), .Y(new_n19382));
  nand_5 g17034(.A(new_n6736_1), .B(new_n6675), .Y(new_n19383));
  nand_5 g17035(.A(new_n6735), .B(n3253), .Y(new_n19384));
  nand_5 g17036(.A(new_n6743), .B(new_n6679), .Y(new_n19385_1));
  nand_5 g17037(.A(new_n6742), .B(n7759), .Y(new_n19386));
  nand_5 g17038(.A(new_n6750), .B(new_n6681), .Y(new_n19387));
  nand_5 g17039(.A(new_n6749), .B(n12562), .Y(new_n19388));
  nand_5 g17040(.A(new_n6758), .B(new_n6682), .Y(new_n19389_1));
  nand_5 g17041(.A(new_n6757), .B(n7949), .Y(new_n19390));
  nand_5 g17042(.A(new_n14935), .B(new_n6685), .Y(new_n19391));
  nand_5 g17043(.A(new_n6770), .B(n24374), .Y(new_n19392));
  nand_5 g17044(.A(n20658), .B(n14575), .Y(new_n19393));
  nand_5 g17045(.A(new_n19393), .B(new_n19392), .Y(new_n19394));
  nand_5 g17046(.A(new_n19394), .B(new_n19391), .Y(new_n19395));
  nand_5 g17047(.A(new_n19395), .B(new_n19390), .Y(new_n19396));
  nand_5 g17048(.A(new_n19396), .B(new_n19389_1), .Y(new_n19397));
  nand_5 g17049(.A(new_n19397), .B(new_n19388), .Y(new_n19398));
  nand_5 g17050(.A(new_n19398), .B(new_n19387), .Y(new_n19399));
  nand_5 g17051(.A(new_n19399), .B(new_n19386), .Y(new_n19400));
  nand_5 g17052(.A(new_n19400), .B(new_n19385_1), .Y(new_n19401_1));
  nand_5 g17053(.A(new_n19401_1), .B(new_n19384), .Y(new_n19402));
  nand_5 g17054(.A(new_n19402), .B(new_n19383), .Y(new_n19403));
  nand_5 g17055(.A(new_n19403), .B(new_n19382), .Y(new_n19404));
  nand_5 g17056(.A(new_n19404), .B(new_n19381), .Y(new_n19405));
  nand_5 g17057(.A(new_n19405), .B(new_n19380), .Y(new_n19406));
  nand_5 g17058(.A(new_n19406), .B(new_n19379), .Y(new_n19407));
  nand_5 g17059(.A(new_n19407), .B(new_n19378), .Y(new_n19408));
  nand_5 g17060(.A(new_n19408), .B(new_n19377), .Y(new_n19409));
  nor_5  g17061(.A(new_n19409), .B(new_n19376), .Y(new_n19410));
  nand_5 g17062(.A(new_n6661), .B(n6456), .Y(new_n19411));
  nand_5 g17063(.A(new_n19411), .B(new_n6660), .Y(new_n19412));
  nor_5  g17064(.A(new_n19412), .B(new_n19410), .Y(new_n19413));
  not_8  g17065(.A(new_n19413), .Y(new_n19414_1));
  nor_5  g17066(.A(new_n19414_1), .B(new_n19374), .Y(new_n19415));
  nand_5 g17067(.A(new_n19414_1), .B(new_n19374), .Y(new_n19416));
  nand_5 g17068(.A(new_n19330), .B(new_n19331), .Y(new_n19417));
  xor_4  g17069(.A(new_n19417), .B(new_n19367_1), .Y(new_n19418));
  nand_5 g17070(.A(new_n19411), .B(new_n19375), .Y(new_n19419));
  xor_4  g17071(.A(new_n19419), .B(new_n19409), .Y(new_n19420));
  nand_5 g17072(.A(new_n19420), .B(new_n19418), .Y(new_n19421));
  nor_5  g17073(.A(new_n19420), .B(new_n19418), .Y(new_n19422));
  not_8  g17074(.A(new_n19422), .Y(new_n19423));
  nand_5 g17075(.A(new_n19332), .B(new_n19333_1), .Y(new_n19424_1));
  xor_4  g17076(.A(new_n19424_1), .B(new_n19365), .Y(new_n19425));
  nand_5 g17077(.A(new_n19378), .B(new_n19377), .Y(new_n19426));
  xor_4  g17078(.A(new_n19426), .B(new_n19407), .Y(new_n19427));
  nand_5 g17079(.A(new_n19427), .B(new_n19425), .Y(new_n19428));
  nor_5  g17080(.A(new_n19427), .B(new_n19425), .Y(new_n19429));
  not_8  g17081(.A(new_n19429), .Y(new_n19430));
  nand_5 g17082(.A(new_n19334), .B(new_n19335), .Y(new_n19431));
  xor_4  g17083(.A(new_n19431), .B(new_n19363), .Y(new_n19432));
  nand_5 g17084(.A(new_n19380), .B(new_n19379), .Y(new_n19433));
  xor_4  g17085(.A(new_n19433), .B(new_n19405), .Y(new_n19434));
  nand_5 g17086(.A(new_n19434), .B(new_n19432), .Y(new_n19435));
  nor_5  g17087(.A(new_n19434), .B(new_n19432), .Y(new_n19436));
  not_8  g17088(.A(new_n19436), .Y(new_n19437));
  nand_5 g17089(.A(new_n19336), .B(new_n19337), .Y(new_n19438));
  xor_4  g17090(.A(new_n19438), .B(new_n19361_1), .Y(new_n19439));
  nand_5 g17091(.A(new_n19382), .B(new_n19381), .Y(new_n19440));
  xor_4  g17092(.A(new_n19440), .B(new_n19403), .Y(new_n19441));
  nand_5 g17093(.A(new_n19441), .B(new_n19439), .Y(new_n19442));
  nor_5  g17094(.A(new_n19441), .B(new_n19439), .Y(new_n19443));
  not_8  g17095(.A(new_n19443), .Y(new_n19444));
  nand_5 g17096(.A(new_n19338), .B(new_n19339), .Y(new_n19445));
  xor_4  g17097(.A(new_n19445), .B(new_n19359), .Y(new_n19446));
  nand_5 g17098(.A(new_n19384), .B(new_n19383), .Y(new_n19447));
  xor_4  g17099(.A(new_n19447), .B(new_n19401_1), .Y(new_n19448));
  nand_5 g17100(.A(new_n19448), .B(new_n19446), .Y(new_n19449));
  nor_5  g17101(.A(new_n19448), .B(new_n19446), .Y(new_n19450_1));
  not_8  g17102(.A(new_n19450_1), .Y(new_n19451));
  nand_5 g17103(.A(new_n19340), .B(new_n19341), .Y(new_n19452));
  xor_4  g17104(.A(new_n19452), .B(new_n19357_1), .Y(new_n19453));
  nand_5 g17105(.A(new_n19386), .B(new_n19385_1), .Y(new_n19454_1));
  xor_4  g17106(.A(new_n19454_1), .B(new_n19399), .Y(new_n19455));
  nand_5 g17107(.A(new_n19455), .B(new_n19453), .Y(new_n19456));
  nor_5  g17108(.A(new_n19455), .B(new_n19453), .Y(new_n19457));
  not_8  g17109(.A(new_n19457), .Y(new_n19458_1));
  nand_5 g17110(.A(new_n19342), .B(new_n19343), .Y(new_n19459));
  xor_4  g17111(.A(new_n19459), .B(new_n19355), .Y(new_n19460));
  nand_5 g17112(.A(new_n19388), .B(new_n19387), .Y(new_n19461));
  xor_4  g17113(.A(new_n19461), .B(new_n19397), .Y(new_n19462));
  nand_5 g17114(.A(new_n19462), .B(new_n19460), .Y(new_n19463));
  or_5   g17115(.A(new_n19462), .B(new_n19460), .Y(new_n19464));
  nand_5 g17116(.A(new_n19346), .B(new_n19344), .Y(new_n19465));
  xor_4  g17117(.A(new_n19465), .B(new_n19352), .Y(new_n19466));
  not_8  g17118(.A(new_n19466), .Y(new_n19467_1));
  nand_5 g17119(.A(new_n19390), .B(new_n19389_1), .Y(new_n19468));
  xor_4  g17120(.A(new_n19468), .B(new_n19395), .Y(new_n19469));
  or_5   g17121(.A(new_n19469), .B(new_n19467_1), .Y(new_n19470));
  nand_5 g17122(.A(new_n19469), .B(new_n19467_1), .Y(new_n19471));
  nand_5 g17123(.A(new_n19392), .B(new_n19391), .Y(new_n19472_1));
  not_8  g17124(.A(new_n19472_1), .Y(new_n19473));
  nand_5 g17125(.A(new_n19473), .B(new_n19393), .Y(new_n19474));
  nor_5  g17126(.A(new_n14486), .B(new_n4699), .Y(new_n19475));
  nor_5  g17127(.A(new_n19475), .B(new_n19350), .Y(new_n19476));
  xor_4  g17128(.A(n20658), .B(n14575), .Y(new_n19477_1));
  nand_5 g17129(.A(new_n19477_1), .B(new_n19476), .Y(new_n19478));
  not_8  g17130(.A(new_n19478), .Y(new_n19479));
  nor_5  g17131(.A(new_n19473), .B(new_n19393), .Y(new_n19480));
  nor_5  g17132(.A(new_n19480), .B(new_n19479), .Y(new_n19481));
  nand_5 g17133(.A(new_n19481), .B(new_n19474), .Y(new_n19482));
  xor_4  g17134(.A(new_n14479), .B(new_n4692), .Y(new_n19483));
  xor_4  g17135(.A(new_n19483), .B(new_n19350), .Y(new_n19484));
  not_8  g17136(.A(new_n19484), .Y(new_n19485));
  nand_5 g17137(.A(new_n19473), .B(new_n19479), .Y(new_n19486));
  nand_5 g17138(.A(new_n19486), .B(new_n19485), .Y(new_n19487));
  nand_5 g17139(.A(new_n19487), .B(new_n19482), .Y(new_n19488));
  nand_5 g17140(.A(new_n19488), .B(new_n19471), .Y(new_n19489));
  and_5  g17141(.A(new_n19489), .B(new_n19470), .Y(new_n19490));
  nand_5 g17142(.A(new_n19490), .B(new_n19464), .Y(new_n19491));
  nand_5 g17143(.A(new_n19491), .B(new_n19463), .Y(new_n19492));
  nand_5 g17144(.A(new_n19492), .B(new_n19458_1), .Y(new_n19493));
  nand_5 g17145(.A(new_n19493), .B(new_n19456), .Y(new_n19494_1));
  nand_5 g17146(.A(new_n19494_1), .B(new_n19451), .Y(new_n19495));
  nand_5 g17147(.A(new_n19495), .B(new_n19449), .Y(new_n19496_1));
  nand_5 g17148(.A(new_n19496_1), .B(new_n19444), .Y(new_n19497));
  nand_5 g17149(.A(new_n19497), .B(new_n19442), .Y(new_n19498));
  nand_5 g17150(.A(new_n19498), .B(new_n19437), .Y(new_n19499));
  nand_5 g17151(.A(new_n19499), .B(new_n19435), .Y(new_n19500));
  nand_5 g17152(.A(new_n19500), .B(new_n19430), .Y(new_n19501));
  nand_5 g17153(.A(new_n19501), .B(new_n19428), .Y(new_n19502));
  nand_5 g17154(.A(new_n19502), .B(new_n19423), .Y(new_n19503));
  nand_5 g17155(.A(new_n19503), .B(new_n19421), .Y(new_n19504));
  and_5  g17156(.A(new_n19504), .B(new_n19416), .Y(new_n19505));
  nor_5  g17157(.A(new_n19505), .B(new_n19415), .Y(new_n19506));
  or_5   g17158(.A(new_n16868), .B(new_n14428), .Y(new_n19507));
  nand_5 g17159(.A(new_n19371), .B(new_n19507), .Y(new_n19508));
  nor_5  g17160(.A(new_n19508), .B(new_n19413), .Y(new_n19509));
  nor_5  g17161(.A(new_n19509), .B(new_n19506), .Y(new_n19510));
  not_8  g17162(.A(new_n19508), .Y(new_n19511));
  nor_5  g17163(.A(new_n19511), .B(new_n19414_1), .Y(new_n19512));
  nor_5  g17164(.A(new_n19512), .B(new_n19505), .Y(new_n19513));
  nor_5  g17165(.A(new_n19513), .B(new_n19510), .Y(n4123));
  nand_5 g17166(.A(new_n15177), .B(new_n9063), .Y(new_n19515_1));
  nand_5 g17167(.A(new_n15176_1), .B(new_n9062), .Y(new_n19516));
  nand_5 g17168(.A(new_n15184), .B(new_n9086), .Y(new_n19517));
  nand_5 g17169(.A(new_n15183), .B(new_n9085), .Y(new_n19518));
  nand_5 g17170(.A(new_n15194), .B(new_n9076), .Y(new_n19519));
  or_5   g17171(.A(new_n15194), .B(new_n9076), .Y(new_n19520));
  nand_5 g17172(.A(new_n11255), .B(new_n9071), .Y(new_n19521));
  nand_5 g17173(.A(new_n19521), .B(new_n19520), .Y(new_n19522));
  nand_5 g17174(.A(new_n19522), .B(new_n19519), .Y(new_n19523_1));
  nand_5 g17175(.A(new_n19523_1), .B(new_n19518), .Y(new_n19524));
  nand_5 g17176(.A(new_n19524), .B(new_n19517), .Y(new_n19525));
  nand_5 g17177(.A(new_n19525), .B(new_n19516), .Y(new_n19526));
  nand_5 g17178(.A(new_n19526), .B(new_n19515_1), .Y(new_n19527));
  nand_5 g17179(.A(new_n15156), .B(new_n9055), .Y(new_n19528));
  nand_5 g17180(.A(new_n15155), .B(new_n9054), .Y(new_n19529));
  nand_5 g17181(.A(new_n19529), .B(new_n19528), .Y(new_n19530));
  xor_4  g17182(.A(new_n19530), .B(new_n19527), .Y(n4134));
  nand_5 g17183(.A(new_n10377), .B(new_n10376), .Y(new_n19532));
  xor_4  g17184(.A(new_n19532), .B(new_n10448), .Y(n4146));
  nand_5 g17185(.A(new_n17527), .B(new_n16222), .Y(new_n19534));
  nand_5 g17186(.A(new_n17528), .B(new_n16223_1), .Y(new_n19535));
  nand_5 g17187(.A(new_n16229), .B(new_n15298), .Y(new_n19536));
  nand_5 g17188(.A(new_n16230_1), .B(new_n15297), .Y(new_n19537));
  nand_5 g17189(.A(new_n16237), .B(new_n15290), .Y(new_n19538));
  nand_5 g17190(.A(new_n19538), .B(new_n19537), .Y(new_n19539_1));
  nand_5 g17191(.A(new_n19539_1), .B(new_n19536), .Y(new_n19540));
  nand_5 g17192(.A(new_n19540), .B(new_n19535), .Y(new_n19541));
  nand_5 g17193(.A(new_n19541), .B(new_n19534), .Y(new_n19542));
  nand_5 g17194(.A(new_n17522), .B(new_n16215_1), .Y(new_n19543));
  nand_5 g17195(.A(new_n17523), .B(new_n16216), .Y(new_n19544));
  nand_5 g17196(.A(new_n19544), .B(new_n19543), .Y(new_n19545));
  xnor_4 g17197(.A(new_n19545), .B(new_n19542), .Y(n4150));
  nand_5 g17198(.A(new_n14347), .B(new_n14346), .Y(new_n19547));
  xor_4  g17199(.A(new_n19547), .B(new_n14356), .Y(n4151));
  nor_5  g17200(.A(new_n14634), .B(new_n14633_1), .Y(new_n19549));
  xor_4  g17201(.A(new_n19549), .B(new_n14711), .Y(n4152));
  nand_5 g17202(.A(new_n6935), .B(new_n6933), .Y(new_n19551));
  xnor_4 g17203(.A(new_n19551), .B(new_n6982), .Y(n4153));
  nand_5 g17204(.A(new_n9979), .B(new_n9944), .Y(new_n19553));
  nand_5 g17205(.A(new_n19553), .B(new_n9945), .Y(new_n19554));
  not_8  g17206(.A(new_n19554), .Y(new_n19555));
  xor_4  g17207(.A(new_n19555), .B(new_n14045), .Y(new_n19556));
  nand_5 g17208(.A(new_n19554), .B(new_n14049), .Y(new_n19557));
  nand_5 g17209(.A(new_n19555), .B(new_n14051), .Y(new_n19558));
  nand_5 g17210(.A(new_n10251), .B(new_n10168), .Y(new_n19559));
  nand_5 g17211(.A(new_n19559), .B(new_n10169), .Y(new_n19560));
  nand_5 g17212(.A(new_n19560), .B(new_n19558), .Y(new_n19561));
  and_5  g17213(.A(new_n19561), .B(new_n19557), .Y(new_n19562));
  xor_4  g17214(.A(new_n19562), .B(new_n19556), .Y(n4165));
  nand_5 g17215(.A(new_n13248), .B(new_n13247), .Y(new_n19564));
  xor_4  g17216(.A(new_n19564), .B(new_n13280), .Y(n4172));
  nand_5 g17217(.A(new_n13103), .B(new_n13104), .Y(new_n19566));
  xor_4  g17218(.A(new_n19566), .B(new_n5277), .Y(n4173));
  nand_5 g17219(.A(new_n7436), .B(new_n7438), .Y(new_n19568));
  xor_4  g17220(.A(new_n19568), .B(new_n7461), .Y(n4176));
  nor_5  g17221(.A(new_n10433), .B(new_n10429), .Y(new_n19570_1));
  xor_4  g17222(.A(new_n19570_1), .B(new_n10431), .Y(n4186));
  nand_5 g17223(.A(new_n19028), .B(new_n19029), .Y(new_n19572));
  xor_4  g17224(.A(new_n19572), .B(new_n19055), .Y(n4204));
  nand_5 g17225(.A(new_n18425), .B(new_n13228), .Y(new_n19574));
  xor_4  g17226(.A(new_n19574), .B(n3984), .Y(new_n19575_1));
  nand_5 g17227(.A(new_n19575_1), .B(new_n13166), .Y(new_n19576));
  not_8  g17228(.A(new_n19576), .Y(new_n19577));
  nor_5  g17229(.A(new_n19575_1), .B(new_n13166), .Y(new_n19578));
  not_8  g17230(.A(new_n19574), .Y(new_n19579));
  nor_5  g17231(.A(new_n18425), .B(new_n13228), .Y(new_n19580));
  or_5   g17232(.A(new_n19580), .B(new_n19579), .Y(new_n19581));
  or_5   g17233(.A(new_n19581), .B(n5386), .Y(new_n19582));
  nand_5 g17234(.A(new_n19581), .B(n5386), .Y(new_n19583));
  nand_5 g17235(.A(new_n18429), .B(new_n18423), .Y(new_n19584_1));
  nand_5 g17236(.A(new_n19584_1), .B(new_n18428), .Y(new_n19585));
  nand_5 g17237(.A(new_n19585), .B(new_n19583), .Y(new_n19586));
  nand_5 g17238(.A(new_n19586), .B(new_n19582), .Y(new_n19587));
  not_8  g17239(.A(new_n19587), .Y(new_n19588));
  nor_5  g17240(.A(new_n19588), .B(new_n19578), .Y(new_n19589));
  nor_5  g17241(.A(new_n19589), .B(new_n19577), .Y(new_n19590));
  not_8  g17242(.A(new_n19590), .Y(new_n19591));
  not_8  g17243(.A(n7569), .Y(new_n19592));
  nand_5 g17244(.A(new_n19579), .B(new_n13223), .Y(new_n19593));
  nor_5  g17245(.A(new_n19593), .B(n4514), .Y(new_n19594));
  not_8  g17246(.A(new_n19594), .Y(new_n19595));
  nand_5 g17247(.A(new_n19593), .B(n4514), .Y(new_n19596));
  and_5  g17248(.A(new_n19596), .B(new_n19595), .Y(new_n19597));
  or_5   g17249(.A(new_n19597), .B(new_n19592), .Y(new_n19598));
  nand_5 g17250(.A(new_n19597), .B(new_n19592), .Y(new_n19599));
  nand_5 g17251(.A(new_n19599), .B(new_n19598), .Y(new_n19600));
  xor_4  g17252(.A(new_n19600), .B(new_n19591), .Y(new_n19601));
  nand_5 g17253(.A(new_n19601), .B(n25586), .Y(new_n19602_1));
  or_5   g17254(.A(new_n19601), .B(n25586), .Y(new_n19603));
  nor_5  g17255(.A(new_n19578), .B(new_n19577), .Y(new_n19604));
  xor_4  g17256(.A(new_n19604), .B(new_n19587), .Y(new_n19605));
  or_5   g17257(.A(new_n19605), .B(new_n16471), .Y(new_n19606));
  nand_5 g17258(.A(new_n19605), .B(new_n16471), .Y(new_n19607));
  nand_5 g17259(.A(new_n19583), .B(new_n19582), .Y(new_n19608_1));
  xnor_4 g17260(.A(new_n19608_1), .B(new_n19585), .Y(new_n19609));
  or_5   g17261(.A(new_n19609), .B(new_n16474), .Y(new_n19610));
  nand_5 g17262(.A(new_n19609), .B(new_n16474), .Y(new_n19611));
  nand_5 g17263(.A(new_n18433), .B(new_n18421), .Y(new_n19612));
  nand_5 g17264(.A(new_n19612), .B(new_n18432), .Y(new_n19613));
  nand_5 g17265(.A(new_n19613), .B(new_n19611), .Y(new_n19614));
  nand_5 g17266(.A(new_n19614), .B(new_n19610), .Y(new_n19615));
  nand_5 g17267(.A(new_n19615), .B(new_n19607), .Y(new_n19616));
  nand_5 g17268(.A(new_n19616), .B(new_n19606), .Y(new_n19617_1));
  nand_5 g17269(.A(new_n19617_1), .B(new_n19603), .Y(new_n19618_1));
  nand_5 g17270(.A(new_n19618_1), .B(new_n19602_1), .Y(new_n19619));
  nand_5 g17271(.A(new_n19598), .B(new_n19591), .Y(new_n19620));
  not_8  g17272(.A(new_n19620), .Y(new_n19621));
  nand_5 g17273(.A(new_n19621), .B(new_n19594), .Y(new_n19622));
  or_5   g17274(.A(new_n19622), .B(new_n19619), .Y(new_n19623_1));
  nand_5 g17275(.A(new_n13140), .B(n13494), .Y(new_n19624));
  nand_5 g17276(.A(new_n13138), .B(new_n6233_1), .Y(new_n19625));
  nand_5 g17277(.A(new_n7965), .B(new_n7954), .Y(new_n19626));
  nand_5 g17278(.A(new_n19626), .B(new_n7964), .Y(new_n19627));
  nand_5 g17279(.A(new_n19627), .B(new_n19625), .Y(new_n19628));
  nand_5 g17280(.A(new_n19628), .B(new_n19624), .Y(new_n19629));
  nand_5 g17281(.A(new_n19629), .B(new_n13135), .Y(new_n19630));
  not_8  g17282(.A(new_n19630), .Y(new_n19631));
  nand_5 g17283(.A(new_n19599), .B(new_n19595), .Y(new_n19632));
  nor_5  g17284(.A(new_n19632), .B(new_n19621), .Y(new_n19633));
  nand_5 g17285(.A(new_n19633), .B(new_n19619), .Y(new_n19634));
  nand_5 g17286(.A(new_n19634), .B(new_n19631), .Y(new_n19635));
  nand_5 g17287(.A(new_n19635), .B(new_n19623_1), .Y(new_n19636));
  or_5   g17288(.A(new_n19629), .B(new_n13135), .Y(new_n19637));
  and_5  g17289(.A(new_n19637), .B(new_n19630), .Y(new_n19638));
  not_8  g17290(.A(new_n19622), .Y(new_n19639));
  nor_5  g17291(.A(new_n19633), .B(new_n19639), .Y(new_n19640));
  xor_4  g17292(.A(new_n19640), .B(new_n19619), .Y(new_n19641_1));
  nand_5 g17293(.A(new_n19641_1), .B(new_n19638), .Y(new_n19642));
  not_8  g17294(.A(new_n19642), .Y(new_n19643));
  nor_5  g17295(.A(new_n19641_1), .B(new_n19638), .Y(new_n19644));
  nand_5 g17296(.A(new_n19624), .B(new_n19625), .Y(new_n19645));
  xor_4  g17297(.A(new_n19645), .B(new_n19627), .Y(new_n19646));
  not_8  g17298(.A(new_n19646), .Y(new_n19647));
  nand_5 g17299(.A(new_n19603), .B(new_n19602_1), .Y(new_n19648_1));
  xor_4  g17300(.A(new_n19648_1), .B(new_n19617_1), .Y(new_n19649));
  nand_5 g17301(.A(new_n19649), .B(new_n19647), .Y(new_n19650));
  nor_5  g17302(.A(new_n19649), .B(new_n19647), .Y(new_n19651));
  not_8  g17303(.A(new_n19651), .Y(new_n19652_1));
  nand_5 g17304(.A(new_n19607), .B(new_n19606), .Y(new_n19653));
  xor_4  g17305(.A(new_n19653), .B(new_n19615), .Y(new_n19654));
  nand_5 g17306(.A(new_n19654), .B(new_n7968_1), .Y(new_n19655));
  nor_5  g17307(.A(new_n19654), .B(new_n7968_1), .Y(new_n19656));
  not_8  g17308(.A(new_n19656), .Y(new_n19657));
  nand_5 g17309(.A(new_n19611), .B(new_n19610), .Y(new_n19658));
  xor_4  g17310(.A(new_n19658), .B(new_n19613), .Y(new_n19659));
  nand_5 g17311(.A(new_n19659), .B(new_n7818), .Y(new_n19660));
  nor_5  g17312(.A(new_n19659), .B(new_n7818), .Y(new_n19661));
  not_8  g17313(.A(new_n18419), .Y(new_n19662));
  nor_5  g17314(.A(new_n18438), .B(new_n19662), .Y(new_n19663));
  nor_5  g17315(.A(new_n19663), .B(new_n18437_1), .Y(new_n19664_1));
  or_5   g17316(.A(new_n19664_1), .B(new_n19661), .Y(new_n19665));
  nand_5 g17317(.A(new_n19665), .B(new_n19660), .Y(new_n19666));
  nand_5 g17318(.A(new_n19666), .B(new_n19657), .Y(new_n19667));
  nand_5 g17319(.A(new_n19667), .B(new_n19655), .Y(new_n19668));
  nand_5 g17320(.A(new_n19668), .B(new_n19652_1), .Y(new_n19669));
  nand_5 g17321(.A(new_n19669), .B(new_n19650), .Y(new_n19670));
  not_8  g17322(.A(new_n19670), .Y(new_n19671));
  nor_5  g17323(.A(new_n19671), .B(new_n19644), .Y(new_n19672));
  nor_5  g17324(.A(new_n19672), .B(new_n19643), .Y(new_n19673));
  nor_5  g17325(.A(new_n19634), .B(new_n19631), .Y(new_n19674));
  nor_5  g17326(.A(new_n19674), .B(new_n19673), .Y(new_n19675));
  nor_5  g17327(.A(new_n19675), .B(new_n19636), .Y(n4205));
  nand_5 g17328(.A(new_n15216), .B(new_n15206), .Y(new_n19677));
  nand_5 g17329(.A(new_n19677), .B(new_n15215), .Y(new_n19678));
  nand_5 g17330(.A(new_n15212), .B(new_n15208), .Y(new_n19679));
  nand_5 g17331(.A(new_n19679), .B(new_n15211), .Y(new_n19680_1));
  nor_5  g17332(.A(new_n15209), .B(n22198), .Y(new_n19681));
  xor_4  g17333(.A(new_n19681), .B(new_n5514), .Y(new_n19682));
  nand_5 g17334(.A(new_n19682), .B(n24638), .Y(new_n19683));
  or_5   g17335(.A(new_n19682), .B(n24638), .Y(new_n19684));
  nand_5 g17336(.A(new_n19684), .B(new_n19683), .Y(new_n19685));
  xor_4  g17337(.A(new_n19685), .B(new_n19680_1), .Y(new_n19686));
  or_5   g17338(.A(new_n19686), .B(new_n8874), .Y(new_n19687));
  nand_5 g17339(.A(new_n19686), .B(new_n8874), .Y(new_n19688));
  nand_5 g17340(.A(new_n19688), .B(new_n19687), .Y(new_n19689));
  xor_4  g17341(.A(new_n19689), .B(new_n19678), .Y(new_n19690));
  nand_5 g17342(.A(new_n15223), .B(new_n15220), .Y(new_n19691));
  nand_5 g17343(.A(new_n19691), .B(new_n15222), .Y(new_n19692));
  not_8  g17344(.A(new_n19692), .Y(new_n19693));
  nand_5 g17345(.A(new_n9834), .B(n23923), .Y(new_n19694));
  nand_5 g17346(.A(n25119), .B(new_n8028), .Y(new_n19695));
  nand_5 g17347(.A(new_n19695), .B(new_n19694), .Y(new_n19696));
  xor_4  g17348(.A(new_n19696), .B(new_n19693), .Y(new_n19697));
  nand_5 g17349(.A(new_n19697), .B(new_n19690), .Y(new_n19698));
  or_5   g17350(.A(new_n19697), .B(new_n19690), .Y(new_n19699));
  nand_5 g17351(.A(new_n15229), .B(new_n15204), .Y(new_n19700));
  nand_5 g17352(.A(new_n19700), .B(new_n15226), .Y(new_n19701_1));
  nand_5 g17353(.A(new_n19701_1), .B(new_n19699), .Y(new_n19702));
  nand_5 g17354(.A(new_n19702), .B(new_n19698), .Y(new_n19703));
  nand_5 g17355(.A(new_n19688), .B(new_n19678), .Y(new_n19704));
  nand_5 g17356(.A(new_n19704), .B(new_n19687), .Y(new_n19705));
  nand_5 g17357(.A(new_n19683), .B(new_n19680_1), .Y(new_n19706));
  nand_5 g17358(.A(new_n19706), .B(new_n19684), .Y(new_n19707));
  nand_5 g17359(.A(new_n19681), .B(new_n5514), .Y(new_n19708));
  xor_4  g17360(.A(new_n19708), .B(n2659), .Y(new_n19709));
  or_5   g17361(.A(new_n19709), .B(n18444), .Y(new_n19710));
  nand_5 g17362(.A(new_n19709), .B(n18444), .Y(new_n19711));
  nand_5 g17363(.A(new_n19711), .B(new_n19710), .Y(new_n19712));
  xor_4  g17364(.A(new_n19712), .B(new_n19707), .Y(new_n19713));
  or_5   g17365(.A(new_n19713), .B(new_n8866), .Y(new_n19714));
  nand_5 g17366(.A(new_n19713), .B(new_n8866), .Y(new_n19715));
  nand_5 g17367(.A(new_n19715), .B(new_n19714), .Y(new_n19716));
  xor_4  g17368(.A(new_n19716), .B(new_n19705), .Y(new_n19717));
  nand_5 g17369(.A(new_n19695), .B(new_n19692), .Y(new_n19718));
  nand_5 g17370(.A(new_n19718), .B(new_n19694), .Y(new_n19719));
  nand_5 g17371(.A(new_n18133), .B(n5400), .Y(new_n19720));
  nand_5 g17372(.A(n21997), .B(new_n8023), .Y(new_n19721));
  nand_5 g17373(.A(new_n19721), .B(new_n19720), .Y(new_n19722));
  xnor_4 g17374(.A(new_n19722), .B(new_n19719), .Y(new_n19723));
  nand_5 g17375(.A(new_n19723), .B(new_n19717), .Y(new_n19724));
  not_8  g17376(.A(new_n19724), .Y(new_n19725));
  nor_5  g17377(.A(new_n19723), .B(new_n19717), .Y(new_n19726));
  nor_5  g17378(.A(new_n19726), .B(new_n19725), .Y(new_n19727));
  xor_4  g17379(.A(new_n19727), .B(new_n19703), .Y(n4215));
  nand_5 g17380(.A(new_n17194), .B(new_n10485), .Y(new_n19729));
  nor_5  g17381(.A(new_n19729), .B(n11356), .Y(new_n19730));
  nand_5 g17382(.A(new_n19730), .B(new_n10479), .Y(new_n19731));
  nor_5  g17383(.A(new_n19731), .B(n6381), .Y(new_n19732));
  nand_5 g17384(.A(new_n19732), .B(new_n10473), .Y(new_n19733));
  nand_5 g17385(.A(new_n19733), .B(n23166), .Y(new_n19734));
  nor_5  g17386(.A(new_n19733), .B(n23166), .Y(new_n19735));
  not_8  g17387(.A(new_n19735), .Y(new_n19736_1));
  and_5  g17388(.A(new_n19736_1), .B(new_n19734), .Y(new_n19737));
  nand_5 g17389(.A(new_n19737), .B(n9554), .Y(new_n19738));
  not_8  g17390(.A(new_n19737), .Y(new_n19739));
  nand_5 g17391(.A(new_n19739), .B(new_n5420), .Y(new_n19740));
  nand_5 g17392(.A(new_n19740), .B(new_n19738), .Y(new_n19741));
  xor_4  g17393(.A(new_n19732), .B(new_n10473), .Y(new_n19742));
  not_8  g17394(.A(new_n19742), .Y(new_n19743));
  nand_5 g17395(.A(new_n19743), .B(new_n5371), .Y(new_n19744));
  nand_5 g17396(.A(new_n19742), .B(n26408), .Y(new_n19745));
  xor_4  g17397(.A(new_n19731), .B(n6381), .Y(new_n19746));
  not_8  g17398(.A(new_n19746), .Y(new_n19747));
  nand_5 g17399(.A(new_n19747), .B(new_n5374), .Y(new_n19748));
  nand_5 g17400(.A(new_n19746), .B(n18227), .Y(new_n19749_1));
  xor_4  g17401(.A(new_n19730), .B(new_n10479), .Y(new_n19750));
  not_8  g17402(.A(new_n19750), .Y(new_n19751));
  nand_5 g17403(.A(new_n19751), .B(new_n5378), .Y(new_n19752));
  nand_5 g17404(.A(new_n19750), .B(n7377), .Y(new_n19753));
  xor_4  g17405(.A(new_n19729), .B(n11356), .Y(new_n19754));
  not_8  g17406(.A(new_n19754), .Y(new_n19755));
  nand_5 g17407(.A(new_n19755), .B(new_n5381), .Y(new_n19756_1));
  nand_5 g17408(.A(new_n19754), .B(n11630), .Y(new_n19757));
  nand_5 g17409(.A(new_n17195), .B(n3164), .Y(new_n19758));
  and_5  g17410(.A(new_n19758), .B(new_n19729), .Y(new_n19759));
  not_8  g17411(.A(new_n19759), .Y(new_n19760));
  nand_5 g17412(.A(new_n19760), .B(new_n5385), .Y(new_n19761));
  nand_5 g17413(.A(new_n19759), .B(n13453), .Y(new_n19762));
  nand_5 g17414(.A(new_n17200), .B(new_n17192), .Y(new_n19763));
  nand_5 g17415(.A(new_n19763), .B(new_n17199), .Y(new_n19764));
  nand_5 g17416(.A(new_n19764), .B(new_n19762), .Y(new_n19765));
  nand_5 g17417(.A(new_n19765), .B(new_n19761), .Y(new_n19766));
  nand_5 g17418(.A(new_n19766), .B(new_n19757), .Y(new_n19767_1));
  nand_5 g17419(.A(new_n19767_1), .B(new_n19756_1), .Y(new_n19768));
  nand_5 g17420(.A(new_n19768), .B(new_n19753), .Y(new_n19769));
  nand_5 g17421(.A(new_n19769), .B(new_n19752), .Y(new_n19770_1));
  nand_5 g17422(.A(new_n19770_1), .B(new_n19749_1), .Y(new_n19771));
  nand_5 g17423(.A(new_n19771), .B(new_n19748), .Y(new_n19772));
  nand_5 g17424(.A(new_n19772), .B(new_n19745), .Y(new_n19773));
  nand_5 g17425(.A(new_n19773), .B(new_n19744), .Y(new_n19774));
  xor_4  g17426(.A(new_n19774), .B(new_n19741), .Y(new_n19775));
  nand_5 g17427(.A(new_n16442), .B(n3582), .Y(new_n19776));
  nor_5  g17428(.A(new_n16442), .B(n3582), .Y(new_n19777));
  not_8  g17429(.A(new_n19777), .Y(new_n19778));
  and_5  g17430(.A(new_n19778), .B(new_n19776), .Y(new_n19779));
  or_5   g17431(.A(new_n19779), .B(n3740), .Y(new_n19780_1));
  nand_5 g17432(.A(new_n19779), .B(n3740), .Y(new_n19781));
  nand_5 g17433(.A(new_n19781), .B(new_n19780_1), .Y(new_n19782));
  nand_5 g17434(.A(new_n16446), .B(new_n16441), .Y(new_n19783));
  nand_5 g17435(.A(new_n19783), .B(new_n16445_1), .Y(new_n19784));
  not_8  g17436(.A(new_n19784), .Y(new_n19785));
  xor_4  g17437(.A(new_n19785), .B(new_n19782), .Y(new_n19786));
  not_8  g17438(.A(new_n19786), .Y(new_n19787));
  nand_5 g17439(.A(new_n11235), .B(n21839), .Y(new_n19788));
  nor_5  g17440(.A(new_n11235), .B(n21839), .Y(new_n19789_1));
  not_8  g17441(.A(new_n19789_1), .Y(new_n19790));
  and_5  g17442(.A(new_n19790), .B(new_n19788), .Y(new_n19791));
  nand_5 g17443(.A(new_n19791), .B(n22626), .Y(new_n19792_1));
  not_8  g17444(.A(new_n19791), .Y(new_n19793));
  nand_5 g17445(.A(new_n19793), .B(new_n8584), .Y(new_n19794));
  nand_5 g17446(.A(new_n19794), .B(new_n19792_1), .Y(new_n19795));
  nand_5 g17447(.A(new_n11238), .B(new_n8574), .Y(new_n19796));
  nand_5 g17448(.A(new_n11237), .B(n14440), .Y(new_n19797));
  nand_5 g17449(.A(new_n18032), .B(new_n18030), .Y(new_n19798_1));
  nand_5 g17450(.A(new_n19798_1), .B(new_n18031), .Y(new_n19799));
  nand_5 g17451(.A(new_n19799), .B(new_n19797), .Y(new_n19800));
  nand_5 g17452(.A(new_n19800), .B(new_n19796), .Y(new_n19801));
  xor_4  g17453(.A(new_n19801), .B(new_n19795), .Y(new_n19802));
  nand_5 g17454(.A(new_n19802), .B(new_n19787), .Y(new_n19803_1));
  not_8  g17455(.A(new_n19802), .Y(new_n19804));
  nand_5 g17456(.A(new_n19804), .B(new_n19786), .Y(new_n19805));
  nand_5 g17457(.A(new_n19805), .B(new_n19803_1), .Y(new_n19806));
  nand_5 g17458(.A(new_n19797), .B(new_n19796), .Y(new_n19807));
  xor_4  g17459(.A(new_n19807), .B(new_n19799), .Y(new_n19808));
  not_8  g17460(.A(new_n19808), .Y(new_n19809));
  nand_5 g17461(.A(new_n19809), .B(new_n16450), .Y(new_n19810));
  nand_5 g17462(.A(new_n19808), .B(new_n16448), .Y(new_n19811));
  nand_5 g17463(.A(new_n18035_1), .B(new_n16362), .Y(new_n19812));
  nand_5 g17464(.A(new_n18034), .B(new_n16360), .Y(new_n19813));
  nand_5 g17465(.A(new_n16319), .B(new_n12312), .Y(new_n19814));
  nand_5 g17466(.A(new_n16317), .B(new_n12322), .Y(new_n19815));
  nand_5 g17467(.A(new_n16324), .B(new_n12263), .Y(new_n19816));
  nand_5 g17468(.A(new_n16322_1), .B(new_n12262), .Y(new_n19817));
  nand_5 g17469(.A(new_n16329), .B(new_n12221), .Y(new_n19818));
  nand_5 g17470(.A(new_n16327_1), .B(new_n12220), .Y(new_n19819));
  nand_5 g17471(.A(new_n10954), .B(new_n10928), .Y(new_n19820));
  nand_5 g17472(.A(new_n19820), .B(new_n10952), .Y(new_n19821));
  nand_5 g17473(.A(new_n19821), .B(new_n19819), .Y(new_n19822));
  nand_5 g17474(.A(new_n19822), .B(new_n19818), .Y(new_n19823));
  nand_5 g17475(.A(new_n19823), .B(new_n19817), .Y(new_n19824));
  nand_5 g17476(.A(new_n19824), .B(new_n19816), .Y(new_n19825));
  nand_5 g17477(.A(new_n19825), .B(new_n19815), .Y(new_n19826));
  nand_5 g17478(.A(new_n19826), .B(new_n19814), .Y(new_n19827));
  nand_5 g17479(.A(new_n19827), .B(new_n19813), .Y(new_n19828));
  nand_5 g17480(.A(new_n19828), .B(new_n19812), .Y(new_n19829));
  nand_5 g17481(.A(new_n19829), .B(new_n19811), .Y(new_n19830));
  nand_5 g17482(.A(new_n19830), .B(new_n19810), .Y(new_n19831));
  xor_4  g17483(.A(new_n19831), .B(new_n19806), .Y(new_n19832));
  nand_5 g17484(.A(new_n19832), .B(new_n19775), .Y(new_n19833));
  not_8  g17485(.A(new_n19775), .Y(new_n19834));
  not_8  g17486(.A(new_n19832), .Y(new_n19835));
  nand_5 g17487(.A(new_n19835), .B(new_n19834), .Y(new_n19836));
  nand_5 g17488(.A(new_n19836), .B(new_n19833), .Y(new_n19837));
  nand_5 g17489(.A(new_n19745), .B(new_n19744), .Y(new_n19838));
  xor_4  g17490(.A(new_n19838), .B(new_n19772), .Y(new_n19839));
  not_8  g17491(.A(new_n19839), .Y(new_n19840));
  nand_5 g17492(.A(new_n19810), .B(new_n19811), .Y(new_n19841));
  xor_4  g17493(.A(new_n19841), .B(new_n19829), .Y(new_n19842));
  not_8  g17494(.A(new_n19842), .Y(new_n19843));
  nand_5 g17495(.A(new_n19843), .B(new_n19840), .Y(new_n19844));
  nand_5 g17496(.A(new_n19842), .B(new_n19839), .Y(new_n19845));
  nand_5 g17497(.A(new_n19749_1), .B(new_n19748), .Y(new_n19846));
  xor_4  g17498(.A(new_n19846), .B(new_n19770_1), .Y(new_n19847));
  not_8  g17499(.A(new_n19847), .Y(new_n19848));
  nand_5 g17500(.A(new_n19812), .B(new_n19813), .Y(new_n19849));
  xor_4  g17501(.A(new_n19849), .B(new_n19827), .Y(new_n19850));
  not_8  g17502(.A(new_n19850), .Y(new_n19851));
  nand_5 g17503(.A(new_n19851), .B(new_n19848), .Y(new_n19852));
  nand_5 g17504(.A(new_n19850), .B(new_n19847), .Y(new_n19853));
  nand_5 g17505(.A(new_n19753), .B(new_n19752), .Y(new_n19854));
  xor_4  g17506(.A(new_n19854), .B(new_n19768), .Y(new_n19855));
  not_8  g17507(.A(new_n19855), .Y(new_n19856));
  nand_5 g17508(.A(new_n19814), .B(new_n19815), .Y(new_n19857));
  xor_4  g17509(.A(new_n19857), .B(new_n19825), .Y(new_n19858));
  not_8  g17510(.A(new_n19858), .Y(new_n19859));
  nand_5 g17511(.A(new_n19859), .B(new_n19856), .Y(new_n19860));
  nand_5 g17512(.A(new_n19858), .B(new_n19855), .Y(new_n19861));
  nand_5 g17513(.A(new_n19757), .B(new_n19756_1), .Y(new_n19862));
  xor_4  g17514(.A(new_n19862), .B(new_n19766), .Y(new_n19863));
  not_8  g17515(.A(new_n19863), .Y(new_n19864));
  nand_5 g17516(.A(new_n19816), .B(new_n19817), .Y(new_n19865));
  xor_4  g17517(.A(new_n19865), .B(new_n19823), .Y(new_n19866));
  not_8  g17518(.A(new_n19866), .Y(new_n19867));
  nand_5 g17519(.A(new_n19867), .B(new_n19864), .Y(new_n19868));
  nand_5 g17520(.A(new_n19866), .B(new_n19863), .Y(new_n19869));
  nand_5 g17521(.A(new_n19762), .B(new_n19761), .Y(new_n19870));
  xor_4  g17522(.A(new_n19870), .B(new_n19764), .Y(new_n19871));
  not_8  g17523(.A(new_n19871), .Y(new_n19872));
  nand_5 g17524(.A(new_n19818), .B(new_n19819), .Y(new_n19873_1));
  xor_4  g17525(.A(new_n19873_1), .B(new_n19821), .Y(new_n19874));
  not_8  g17526(.A(new_n19874), .Y(new_n19875));
  nand_5 g17527(.A(new_n19875), .B(new_n19872), .Y(new_n19876));
  nand_5 g17528(.A(new_n19874), .B(new_n19871), .Y(new_n19877));
  or_5   g17529(.A(new_n17203), .B(new_n10956), .Y(new_n19878));
  nand_5 g17530(.A(new_n17203), .B(new_n10956), .Y(new_n19879));
  nand_5 g17531(.A(new_n17178), .B(new_n10896), .Y(new_n19880));
  or_5   g17532(.A(new_n17178), .B(new_n10896), .Y(new_n19881));
  not_8  g17533(.A(new_n10920), .Y(new_n19882));
  nand_5 g17534(.A(new_n17181), .B(new_n19882), .Y(new_n19883));
  or_5   g17535(.A(new_n17181), .B(new_n19882), .Y(new_n19884));
  nand_5 g17536(.A(new_n17184), .B(new_n10910), .Y(new_n19885));
  nand_5 g17537(.A(new_n19885), .B(new_n19884), .Y(new_n19886));
  nand_5 g17538(.A(new_n19886), .B(new_n19883), .Y(new_n19887));
  nand_5 g17539(.A(new_n19887), .B(new_n19881), .Y(new_n19888));
  nand_5 g17540(.A(new_n19888), .B(new_n19880), .Y(new_n19889));
  nand_5 g17541(.A(new_n19889), .B(new_n19879), .Y(new_n19890));
  nand_5 g17542(.A(new_n19890), .B(new_n19878), .Y(new_n19891));
  nand_5 g17543(.A(new_n19891), .B(new_n19877), .Y(new_n19892));
  nand_5 g17544(.A(new_n19892), .B(new_n19876), .Y(new_n19893));
  nand_5 g17545(.A(new_n19893), .B(new_n19869), .Y(new_n19894));
  nand_5 g17546(.A(new_n19894), .B(new_n19868), .Y(new_n19895));
  nand_5 g17547(.A(new_n19895), .B(new_n19861), .Y(new_n19896));
  nand_5 g17548(.A(new_n19896), .B(new_n19860), .Y(new_n19897));
  nand_5 g17549(.A(new_n19897), .B(new_n19853), .Y(new_n19898));
  nand_5 g17550(.A(new_n19898), .B(new_n19852), .Y(new_n19899));
  nand_5 g17551(.A(new_n19899), .B(new_n19845), .Y(new_n19900));
  nand_5 g17552(.A(new_n19900), .B(new_n19844), .Y(new_n19901));
  xor_4  g17553(.A(new_n19901), .B(new_n19837), .Y(n4221));
  nand_5 g17554(.A(new_n12134), .B(n11630), .Y(new_n19903));
  nand_5 g17555(.A(new_n12133), .B(new_n5381), .Y(new_n19904));
  nand_5 g17556(.A(new_n14844), .B(new_n14842), .Y(new_n19905_1));
  nand_5 g17557(.A(new_n19905_1), .B(new_n14843), .Y(new_n19906));
  nand_5 g17558(.A(new_n19906), .B(new_n19904), .Y(new_n19907));
  nand_5 g17559(.A(new_n19907), .B(new_n19903), .Y(new_n19908));
  nand_5 g17560(.A(new_n12156), .B(n7377), .Y(new_n19909_1));
  nand_5 g17561(.A(new_n12155), .B(new_n5378), .Y(new_n19910));
  nand_5 g17562(.A(new_n19910), .B(new_n19909_1), .Y(new_n19911_1));
  xor_4  g17563(.A(new_n19911_1), .B(new_n19908), .Y(new_n19912));
  not_8  g17564(.A(new_n19912), .Y(new_n19913));
  nand_5 g17565(.A(new_n19913), .B(new_n9831), .Y(new_n19914));
  or_5   g17566(.A(new_n19913), .B(new_n9831), .Y(new_n19915));
  nand_5 g17567(.A(new_n19903), .B(new_n19904), .Y(new_n19916_1));
  xor_4  g17568(.A(new_n19916_1), .B(new_n19906), .Y(new_n19917));
  not_8  g17569(.A(new_n19917), .Y(new_n19918));
  nand_5 g17570(.A(new_n19918), .B(new_n9756), .Y(new_n19919));
  or_5   g17571(.A(new_n19918), .B(new_n9756), .Y(new_n19920));
  nand_5 g17572(.A(new_n14849_1), .B(new_n9786), .Y(new_n19921));
  or_5   g17573(.A(new_n14849_1), .B(new_n9786), .Y(new_n19922_1));
  nand_5 g17574(.A(new_n9792), .B(new_n7632), .Y(new_n19923_1));
  nand_5 g17575(.A(new_n18518), .B(new_n7629), .Y(new_n19924));
  nand_5 g17576(.A(new_n9798), .B(new_n7578), .Y(new_n19925));
  nand_5 g17577(.A(new_n18524), .B(new_n7577), .Y(new_n19926));
  nand_5 g17578(.A(new_n9804), .B(new_n7586), .Y(new_n19927));
  nand_5 g17579(.A(new_n9805), .B(new_n7585_1), .Y(new_n19928));
  nor_5  g17580(.A(new_n9811), .B(new_n7593_1), .Y(new_n19929));
  nand_5 g17581(.A(new_n19929), .B(new_n19928), .Y(new_n19930_1));
  nand_5 g17582(.A(new_n19930_1), .B(new_n19927), .Y(new_n19931));
  nand_5 g17583(.A(new_n19931), .B(new_n19926), .Y(new_n19932));
  nand_5 g17584(.A(new_n19932), .B(new_n19925), .Y(new_n19933));
  nand_5 g17585(.A(new_n19933), .B(new_n19924), .Y(new_n19934));
  nand_5 g17586(.A(new_n19934), .B(new_n19923_1), .Y(new_n19935));
  nand_5 g17587(.A(new_n19935), .B(new_n19922_1), .Y(new_n19936));
  nand_5 g17588(.A(new_n19936), .B(new_n19921), .Y(new_n19937));
  nand_5 g17589(.A(new_n19937), .B(new_n19920), .Y(new_n19938));
  nand_5 g17590(.A(new_n19938), .B(new_n19919), .Y(new_n19939));
  nand_5 g17591(.A(new_n19939), .B(new_n19915), .Y(new_n19940));
  nand_5 g17592(.A(new_n19940), .B(new_n19914), .Y(new_n19941_1));
  nand_5 g17593(.A(new_n19910), .B(new_n19908), .Y(new_n19942));
  nand_5 g17594(.A(new_n19942), .B(new_n19909_1), .Y(new_n19943));
  nand_5 g17595(.A(new_n12205), .B(n18227), .Y(new_n19944));
  nand_5 g17596(.A(new_n12204), .B(new_n5374), .Y(new_n19945));
  nand_5 g17597(.A(new_n19945), .B(new_n19944), .Y(new_n19946));
  xor_4  g17598(.A(new_n19946), .B(new_n19943), .Y(new_n19947));
  nand_5 g17599(.A(new_n19947), .B(new_n18448), .Y(new_n19948));
  not_8  g17600(.A(new_n19947), .Y(new_n19949));
  nand_5 g17601(.A(new_n19949), .B(new_n18447), .Y(new_n19950));
  nand_5 g17602(.A(new_n19950), .B(new_n19948), .Y(new_n19951));
  xor_4  g17603(.A(new_n19951), .B(new_n19941_1), .Y(n4224));
  nand_5 g17604(.A(new_n12291), .B(new_n12292), .Y(new_n19953));
  xor_4  g17605(.A(new_n19953), .B(new_n12294), .Y(n4231));
  nand_5 g17606(.A(new_n16116), .B(n9934), .Y(new_n19955));
  nand_5 g17607(.A(new_n16117), .B(new_n5326), .Y(new_n19956));
  nand_5 g17608(.A(new_n19956), .B(new_n19955), .Y(new_n19957));
  nand_5 g17609(.A(new_n19216), .B(new_n19213), .Y(new_n19958));
  nand_5 g17610(.A(new_n19958), .B(new_n19215), .Y(new_n19959));
  xor_4  g17611(.A(new_n19959), .B(new_n19957), .Y(new_n19960));
  nand_5 g17612(.A(new_n19960), .B(n2979), .Y(new_n19961));
  not_8  g17613(.A(new_n19960), .Y(new_n19962));
  nand_5 g17614(.A(new_n19962), .B(new_n5369), .Y(new_n19963));
  nand_5 g17615(.A(new_n19963), .B(new_n19961), .Y(new_n19964));
  nand_5 g17616(.A(new_n19220_1), .B(new_n19211), .Y(new_n19965));
  nand_5 g17617(.A(new_n19965), .B(new_n19219), .Y(new_n19966));
  xor_4  g17618(.A(new_n19966), .B(new_n19964), .Y(new_n19967));
  nand_5 g17619(.A(new_n19967), .B(new_n13564), .Y(new_n19968_1));
  or_5   g17620(.A(new_n19967), .B(new_n13564), .Y(new_n19969));
  nand_5 g17621(.A(new_n19969), .B(new_n19968_1), .Y(new_n19970));
  nand_5 g17622(.A(new_n19223_1), .B(new_n19209), .Y(new_n19971));
  nand_5 g17623(.A(new_n19971), .B(new_n19224_1), .Y(new_n19972));
  xnor_4 g17624(.A(new_n19972), .B(new_n19970), .Y(n4266));
  nand_5 g17625(.A(new_n7913), .B(new_n7912), .Y(new_n19974));
  xnor_4 g17626(.A(new_n19974), .B(new_n7944), .Y(n4340));
  nand_5 g17627(.A(new_n18748), .B(new_n18746), .Y(new_n19976));
  nand_5 g17628(.A(new_n19976), .B(new_n18747), .Y(new_n19977));
  not_8  g17629(.A(new_n5625), .Y(new_n19978));
  nor_5  g17630(.A(new_n18744), .B(new_n12530), .Y(new_n19979));
  nor_5  g17631(.A(new_n19979), .B(new_n18743), .Y(new_n19980));
  xor_4  g17632(.A(new_n18739), .B(new_n6760), .Y(new_n19981));
  or_5   g17633(.A(new_n19981), .B(new_n14951), .Y(new_n19982));
  nand_5 g17634(.A(new_n19981), .B(new_n14951), .Y(new_n19983));
  nand_5 g17635(.A(new_n19983), .B(new_n19982), .Y(new_n19984));
  xor_4  g17636(.A(new_n19984), .B(new_n19980), .Y(new_n19985));
  or_5   g17637(.A(new_n19985), .B(new_n19978), .Y(new_n19986));
  nand_5 g17638(.A(new_n19985), .B(new_n19978), .Y(new_n19987));
  nand_5 g17639(.A(new_n19987), .B(new_n19986), .Y(new_n19988_1));
  xnor_4 g17640(.A(new_n19988_1), .B(new_n19977), .Y(n4374));
  nand_5 g17641(.A(new_n12828), .B(new_n12827), .Y(new_n19990));
  xor_4  g17642(.A(new_n19990), .B(new_n12887), .Y(n4401));
  nand_5 g17643(.A(new_n14870), .B(new_n14869), .Y(new_n19992));
  xnor_4 g17644(.A(new_n19992), .B(new_n14872), .Y(n4424));
  nand_5 g17645(.A(new_n12407), .B(new_n12401), .Y(new_n19994));
  nand_5 g17646(.A(new_n19994), .B(new_n12404), .Y(new_n19995));
  not_8  g17647(.A(new_n19995), .Y(new_n19996));
  nand_5 g17648(.A(new_n12408_1), .B(n1881), .Y(new_n19997));
  not_8  g17649(.A(n1881), .Y(new_n19998));
  not_8  g17650(.A(new_n12408_1), .Y(new_n19999));
  nand_5 g17651(.A(new_n19999), .B(new_n19998), .Y(new_n20000));
  nand_5 g17652(.A(new_n12398_1), .B(n5834), .Y(new_n20001));
  not_8  g17653(.A(n5834), .Y(new_n20002));
  nand_5 g17654(.A(new_n12399), .B(new_n20002), .Y(new_n20003));
  nand_5 g17655(.A(new_n12388), .B(n13851), .Y(new_n20004_1));
  nand_5 g17656(.A(new_n12389), .B(new_n17634), .Y(new_n20005));
  nand_5 g17657(.A(new_n18646), .B(new_n18643), .Y(new_n20006));
  nand_5 g17658(.A(new_n20006), .B(new_n18644), .Y(new_n20007));
  nand_5 g17659(.A(new_n20007), .B(new_n20005), .Y(new_n20008));
  nand_5 g17660(.A(new_n20008), .B(new_n20004_1), .Y(new_n20009));
  nand_5 g17661(.A(new_n20009), .B(new_n20003), .Y(new_n20010));
  nand_5 g17662(.A(new_n20010), .B(new_n20001), .Y(new_n20011));
  nand_5 g17663(.A(new_n20011), .B(new_n20000), .Y(new_n20012));
  nand_5 g17664(.A(new_n20012), .B(new_n19997), .Y(new_n20013_1));
  nand_5 g17665(.A(new_n20013_1), .B(new_n19996), .Y(new_n20014));
  or_5   g17666(.A(new_n20013_1), .B(new_n19996), .Y(new_n20015));
  and_5  g17667(.A(new_n20015), .B(new_n20014), .Y(new_n20016));
  not_8  g17668(.A(new_n20016), .Y(new_n20017_1));
  nand_5 g17669(.A(new_n20017_1), .B(new_n11528), .Y(new_n20018));
  nand_5 g17670(.A(new_n20016), .B(new_n11529), .Y(new_n20019));
  nand_5 g17671(.A(new_n20019), .B(new_n20018), .Y(new_n20020));
  nand_5 g17672(.A(new_n19997), .B(new_n20000), .Y(new_n20021));
  xor_4  g17673(.A(new_n20021), .B(new_n20011), .Y(new_n20022));
  not_8  g17674(.A(new_n20022), .Y(new_n20023));
  nand_5 g17675(.A(new_n20023), .B(new_n11535), .Y(new_n20024));
  or_5   g17676(.A(new_n20023), .B(new_n11535), .Y(new_n20025));
  nand_5 g17677(.A(new_n20001), .B(new_n20003), .Y(new_n20026));
  xor_4  g17678(.A(new_n20026), .B(new_n20009), .Y(new_n20027));
  or_5   g17679(.A(new_n20027), .B(new_n11542), .Y(new_n20028));
  nand_5 g17680(.A(new_n20027), .B(new_n11542), .Y(new_n20029));
  nand_5 g17681(.A(new_n20004_1), .B(new_n20005), .Y(new_n20030));
  xor_4  g17682(.A(new_n20030), .B(new_n20007), .Y(new_n20031));
  or_5   g17683(.A(new_n20031), .B(new_n11549), .Y(new_n20032));
  nand_5 g17684(.A(new_n20031), .B(new_n11549), .Y(new_n20033_1));
  nand_5 g17685(.A(new_n18650), .B(new_n18641), .Y(new_n20034));
  nand_5 g17686(.A(new_n20034), .B(new_n18649_1), .Y(new_n20035));
  nand_5 g17687(.A(new_n20035), .B(new_n20033_1), .Y(new_n20036_1));
  nand_5 g17688(.A(new_n20036_1), .B(new_n20032), .Y(new_n20037));
  nand_5 g17689(.A(new_n20037), .B(new_n20029), .Y(new_n20038));
  nand_5 g17690(.A(new_n20038), .B(new_n20028), .Y(new_n20039));
  nand_5 g17691(.A(new_n20039), .B(new_n20025), .Y(new_n20040_1));
  nand_5 g17692(.A(new_n20040_1), .B(new_n20024), .Y(new_n20041));
  xor_4  g17693(.A(new_n20041), .B(new_n20020), .Y(n4432));
  nand_5 g17694(.A(new_n16787), .B(new_n16785), .Y(new_n20043));
  xor_4  g17695(.A(new_n20043), .B(new_n16811), .Y(n4441));
  nand_5 g17696(.A(new_n4553), .B(new_n4542), .Y(new_n20045));
  or_5   g17697(.A(new_n20045), .B(n24786), .Y(new_n20046));
  nor_5  g17698(.A(new_n20046), .B(n25370), .Y(new_n20047));
  nand_5 g17699(.A(new_n20047), .B(new_n7822), .Y(new_n20048));
  xor_4  g17700(.A(new_n20048), .B(new_n7819), .Y(new_n20049));
  or_5   g17701(.A(new_n20049), .B(new_n19257), .Y(new_n20050));
  nand_5 g17702(.A(new_n20049), .B(new_n19257), .Y(new_n20051));
  xor_4  g17703(.A(new_n20047), .B(n19472), .Y(new_n20052));
  or_5   g17704(.A(new_n20052), .B(new_n9934_1), .Y(new_n20053));
  nand_5 g17705(.A(new_n20052), .B(new_n9934_1), .Y(new_n20054));
  xor_4  g17706(.A(new_n20046), .B(new_n7825), .Y(new_n20055));
  or_5   g17707(.A(new_n20055), .B(new_n9891), .Y(new_n20056));
  nand_5 g17708(.A(new_n20055), .B(new_n9891), .Y(new_n20057));
  nand_5 g17709(.A(new_n20045), .B(n24786), .Y(new_n20058));
  nand_5 g17710(.A(new_n20058), .B(new_n20046), .Y(new_n20059));
  or_5   g17711(.A(new_n20059), .B(new_n9860), .Y(new_n20060));
  nand_5 g17712(.A(new_n20059), .B(new_n9860), .Y(new_n20061_1));
  xor_4  g17713(.A(n27120), .B(n23065), .Y(new_n20062));
  nand_5 g17714(.A(new_n20062), .B(new_n9874), .Y(new_n20063));
  nand_5 g17715(.A(new_n20063), .B(new_n9870), .Y(new_n20064));
  nand_5 g17716(.A(new_n20064), .B(new_n20061_1), .Y(new_n20065));
  nand_5 g17717(.A(new_n20065), .B(new_n20060), .Y(new_n20066));
  nand_5 g17718(.A(new_n20066), .B(new_n20057), .Y(new_n20067));
  nand_5 g17719(.A(new_n20067), .B(new_n20056), .Y(new_n20068));
  nand_5 g17720(.A(new_n20068), .B(new_n20054), .Y(new_n20069_1));
  nand_5 g17721(.A(new_n20069_1), .B(new_n20053), .Y(new_n20070));
  nand_5 g17722(.A(new_n20070), .B(new_n20051), .Y(new_n20071));
  nand_5 g17723(.A(new_n20071), .B(new_n20050), .Y(new_n20072));
  nor_5  g17724(.A(new_n20048), .B(n19042), .Y(new_n20073));
  xor_4  g17725(.A(new_n20073), .B(n1293), .Y(new_n20074));
  or_5   g17726(.A(new_n20074), .B(new_n19270_1), .Y(new_n20075));
  nand_5 g17727(.A(new_n20074), .B(new_n19270_1), .Y(new_n20076));
  nand_5 g17728(.A(new_n20076), .B(new_n20075), .Y(new_n20077_1));
  xor_4  g17729(.A(new_n20077_1), .B(new_n20072), .Y(new_n20078));
  nand_5 g17730(.A(new_n20078), .B(new_n13979), .Y(new_n20079));
  or_5   g17731(.A(new_n20078), .B(new_n13979), .Y(new_n20080));
  nand_5 g17732(.A(new_n20050), .B(new_n20051), .Y(new_n20081));
  xor_4  g17733(.A(new_n20081), .B(new_n20070), .Y(new_n20082));
  nand_5 g17734(.A(new_n20082), .B(new_n13896), .Y(new_n20083));
  or_5   g17735(.A(new_n20082), .B(new_n13896), .Y(new_n20084));
  nand_5 g17736(.A(new_n20053), .B(new_n20054), .Y(new_n20085));
  xor_4  g17737(.A(new_n20085), .B(new_n20068), .Y(new_n20086_1));
  nand_5 g17738(.A(new_n20086_1), .B(new_n13928), .Y(new_n20087));
  or_5   g17739(.A(new_n20086_1), .B(new_n13928), .Y(new_n20088));
  nand_5 g17740(.A(new_n20057), .B(new_n20056), .Y(new_n20089));
  xor_4  g17741(.A(new_n20089), .B(new_n20066), .Y(new_n20090));
  nand_5 g17742(.A(new_n20090), .B(new_n13935), .Y(new_n20091));
  or_5   g17743(.A(new_n20090), .B(new_n13935), .Y(new_n20092));
  nand_5 g17744(.A(new_n20061_1), .B(new_n20060), .Y(new_n20093));
  xnor_4 g17745(.A(new_n20093), .B(new_n20064), .Y(new_n20094));
  or_5   g17746(.A(new_n20094), .B(new_n13945), .Y(new_n20095));
  nand_5 g17747(.A(new_n20094), .B(new_n13945), .Y(new_n20096_1));
  xor_4  g17748(.A(new_n9902), .B(n23065), .Y(new_n20097));
  not_8  g17749(.A(new_n20097), .Y(new_n20098));
  or_5   g17750(.A(new_n20098), .B(new_n13951_1), .Y(new_n20099));
  nand_5 g17751(.A(new_n20098), .B(new_n13951_1), .Y(new_n20100));
  nand_5 g17752(.A(new_n13957), .B(new_n9906), .Y(new_n20101));
  nand_5 g17753(.A(new_n20101), .B(new_n20100), .Y(new_n20102));
  nand_5 g17754(.A(new_n20102), .B(new_n20099), .Y(new_n20103_1));
  nand_5 g17755(.A(new_n20103_1), .B(new_n20096_1), .Y(new_n20104));
  nand_5 g17756(.A(new_n20104), .B(new_n20095), .Y(new_n20105));
  nand_5 g17757(.A(new_n20105), .B(new_n20092), .Y(new_n20106));
  nand_5 g17758(.A(new_n20106), .B(new_n20091), .Y(new_n20107));
  nand_5 g17759(.A(new_n20107), .B(new_n20088), .Y(new_n20108));
  nand_5 g17760(.A(new_n20108), .B(new_n20087), .Y(new_n20109));
  nand_5 g17761(.A(new_n20109), .B(new_n20084), .Y(new_n20110));
  nand_5 g17762(.A(new_n20110), .B(new_n20083), .Y(new_n20111));
  nand_5 g17763(.A(new_n20111), .B(new_n20080), .Y(new_n20112));
  nand_5 g17764(.A(new_n20112), .B(new_n20079), .Y(new_n20113));
  nand_5 g17765(.A(new_n13977), .B(new_n13974), .Y(new_n20114));
  nand_5 g17766(.A(new_n20114), .B(new_n13976), .Y(new_n20115));
  nand_5 g17767(.A(new_n13890), .B(new_n11706), .Y(new_n20116));
  xor_4  g17768(.A(new_n20116), .B(n3710), .Y(new_n20117));
  nand_5 g17769(.A(new_n20117), .B(new_n6066), .Y(new_n20118));
  or_5   g17770(.A(new_n20117), .B(new_n6066), .Y(new_n20119));
  nand_5 g17771(.A(new_n20119), .B(new_n20118), .Y(new_n20120));
  xor_4  g17772(.A(new_n20120), .B(new_n20115), .Y(new_n20121));
  nand_5 g17773(.A(new_n20076), .B(new_n20072), .Y(new_n20122));
  nand_5 g17774(.A(new_n20122), .B(new_n20075), .Y(new_n20123));
  nand_5 g17775(.A(new_n20073), .B(new_n7838), .Y(new_n20124));
  not_8  g17776(.A(new_n20124), .Y(new_n20125));
  nand_5 g17777(.A(new_n20125), .B(new_n7882), .Y(new_n20126_1));
  nand_5 g17778(.A(new_n20124), .B(n13775), .Y(new_n20127));
  nand_5 g17779(.A(new_n20127), .B(new_n20126_1), .Y(new_n20128));
  or_5   g17780(.A(new_n20128), .B(new_n19312), .Y(new_n20129));
  nand_5 g17781(.A(new_n20128), .B(new_n19312), .Y(new_n20130));
  nand_5 g17782(.A(new_n20130), .B(new_n20129), .Y(new_n20131));
  xor_4  g17783(.A(new_n20131), .B(new_n20123), .Y(new_n20132));
  nand_5 g17784(.A(new_n20132), .B(new_n20121), .Y(new_n20133));
  or_5   g17785(.A(new_n20132), .B(new_n20121), .Y(new_n20134));
  nand_5 g17786(.A(new_n20134), .B(new_n20133), .Y(new_n20135));
  xor_4  g17787(.A(new_n20135), .B(new_n20113), .Y(n4451));
  not_8  g17788(.A(new_n15066), .Y(new_n20137));
  nand_5 g17789(.A(new_n12993), .B(n6659), .Y(new_n20138_1));
  nand_5 g17790(.A(n25494), .B(new_n18162), .Y(new_n20139));
  nand_5 g17791(.A(new_n20139), .B(new_n20138_1), .Y(new_n20140));
  nand_5 g17792(.A(n23250), .B(new_n12973), .Y(new_n20141));
  nand_5 g17793(.A(new_n18166), .B(n10117), .Y(new_n20142));
  nand_5 g17794(.A(new_n12976), .B(n11455), .Y(new_n20143));
  nand_5 g17795(.A(n13460), .B(new_n18169), .Y(new_n20144));
  nand_5 g17796(.A(new_n12980_1), .B(n3945), .Y(new_n20145));
  nand_5 g17797(.A(n6104), .B(new_n18172), .Y(new_n20146));
  nand_5 g17798(.A(new_n5880), .B(new_n5876), .Y(new_n20147));
  nand_5 g17799(.A(new_n20147), .B(new_n5878), .Y(new_n20148));
  nand_5 g17800(.A(new_n20148), .B(new_n20146), .Y(new_n20149_1));
  nand_5 g17801(.A(new_n20149_1), .B(new_n20145), .Y(new_n20150));
  nand_5 g17802(.A(new_n20150), .B(new_n20144), .Y(new_n20151_1));
  nand_5 g17803(.A(new_n20151_1), .B(new_n20143), .Y(new_n20152));
  nand_5 g17804(.A(new_n20152), .B(new_n20142), .Y(new_n20153));
  nand_5 g17805(.A(new_n20153), .B(new_n20141), .Y(new_n20154));
  not_8  g17806(.A(new_n20154), .Y(new_n20155));
  xor_4  g17807(.A(new_n20155), .B(new_n20140), .Y(new_n20156));
  or_5   g17808(.A(new_n20156), .B(new_n20137), .Y(new_n20157));
  nand_5 g17809(.A(new_n20156), .B(new_n20137), .Y(new_n20158));
  nand_5 g17810(.A(new_n20158), .B(new_n20157), .Y(new_n20159));
  nand_5 g17811(.A(new_n20142), .B(new_n20141), .Y(new_n20160));
  xor_4  g17812(.A(new_n20160), .B(new_n20152), .Y(new_n20161));
  nand_5 g17813(.A(new_n20161), .B(new_n15072), .Y(new_n20162));
  or_5   g17814(.A(new_n20161), .B(new_n15072), .Y(new_n20163));
  nand_5 g17815(.A(new_n20144), .B(new_n20143), .Y(new_n20164));
  xor_4  g17816(.A(new_n20164), .B(new_n20150), .Y(new_n20165));
  nand_5 g17817(.A(new_n20165), .B(new_n15078), .Y(new_n20166));
  or_5   g17818(.A(new_n20165), .B(new_n15078), .Y(new_n20167));
  nand_5 g17819(.A(new_n20146), .B(new_n20145), .Y(new_n20168));
  xor_4  g17820(.A(new_n20168), .B(new_n20148), .Y(new_n20169_1));
  nand_5 g17821(.A(new_n20169_1), .B(new_n15084), .Y(new_n20170));
  not_8  g17822(.A(new_n20170), .Y(new_n20171));
  nor_5  g17823(.A(new_n20169_1), .B(new_n15084), .Y(new_n20172));
  nor_5  g17824(.A(new_n5886), .B(new_n5858), .Y(new_n20173));
  nor_5  g17825(.A(new_n20173), .B(new_n5884), .Y(new_n20174));
  nor_5  g17826(.A(new_n20174), .B(new_n20172), .Y(new_n20175));
  nor_5  g17827(.A(new_n20175), .B(new_n20171), .Y(new_n20176));
  not_8  g17828(.A(new_n20176), .Y(new_n20177));
  nand_5 g17829(.A(new_n20177), .B(new_n20167), .Y(new_n20178));
  nand_5 g17830(.A(new_n20178), .B(new_n20166), .Y(new_n20179_1));
  nand_5 g17831(.A(new_n20179_1), .B(new_n20163), .Y(new_n20180));
  nand_5 g17832(.A(new_n20180), .B(new_n20162), .Y(new_n20181));
  xor_4  g17833(.A(new_n20181), .B(new_n20159), .Y(n4476));
  not_8  g17834(.A(new_n13413), .Y(new_n20183));
  nor_5  g17835(.A(new_n4524), .B(n12398), .Y(new_n20184));
  nand_5 g17836(.A(new_n20184), .B(new_n7004), .Y(new_n20185));
  nor_5  g17837(.A(new_n20185), .B(n18452), .Y(new_n20186));
  nand_5 g17838(.A(new_n20186), .B(new_n6992), .Y(new_n20187_1));
  nor_5  g17839(.A(new_n20187_1), .B(n1831), .Y(new_n20188));
  xor_4  g17840(.A(new_n20187_1), .B(n1831), .Y(new_n20189));
  or_5   g17841(.A(new_n20189), .B(new_n7089), .Y(new_n20190));
  xor_4  g17842(.A(new_n20186), .B(n13137), .Y(new_n20191));
  or_5   g17843(.A(new_n20191), .B(new_n7098), .Y(new_n20192));
  nand_5 g17844(.A(new_n20191), .B(new_n7098), .Y(new_n20193));
  xor_4  g17845(.A(new_n20185), .B(new_n6998_1), .Y(new_n20194));
  or_5   g17846(.A(new_n20194), .B(new_n7106), .Y(new_n20195));
  nand_5 g17847(.A(new_n20194), .B(new_n7106), .Y(new_n20196));
  xor_4  g17848(.A(new_n20184), .B(n21317), .Y(new_n20197));
  or_5   g17849(.A(new_n20197), .B(new_n7114), .Y(new_n20198));
  nand_5 g17850(.A(new_n20197), .B(new_n7114), .Y(new_n20199));
  nand_5 g17851(.A(new_n4527), .B(new_n4509), .Y(new_n20200));
  nand_5 g17852(.A(new_n20200), .B(new_n4526), .Y(new_n20201));
  nand_5 g17853(.A(new_n20201), .B(new_n20199), .Y(new_n20202));
  nand_5 g17854(.A(new_n20202), .B(new_n20198), .Y(new_n20203));
  nand_5 g17855(.A(new_n20203), .B(new_n20196), .Y(new_n20204));
  nand_5 g17856(.A(new_n20204), .B(new_n20195), .Y(new_n20205));
  nand_5 g17857(.A(new_n20205), .B(new_n20193), .Y(new_n20206));
  nand_5 g17858(.A(new_n20206), .B(new_n20192), .Y(new_n20207));
  nand_5 g17859(.A(new_n20207), .B(new_n20190), .Y(new_n20208));
  nand_5 g17860(.A(new_n20189), .B(new_n7089), .Y(new_n20209));
  nand_5 g17861(.A(new_n20209), .B(new_n20208), .Y(new_n20210));
  or_5   g17862(.A(new_n20210), .B(new_n20188), .Y(new_n20211));
  xor_4  g17863(.A(new_n20211), .B(new_n7082), .Y(new_n20212));
  nand_5 g17864(.A(new_n20212), .B(new_n20183), .Y(new_n20213_1));
  nor_5  g17865(.A(new_n20212), .B(new_n20183), .Y(new_n20214));
  not_8  g17866(.A(new_n20214), .Y(new_n20215));
  nand_5 g17867(.A(new_n20215), .B(new_n20213_1), .Y(new_n20216));
  nand_5 g17868(.A(new_n20209), .B(new_n20190), .Y(new_n20217));
  xor_4  g17869(.A(new_n20217), .B(new_n20207), .Y(new_n20218));
  nand_5 g17870(.A(new_n20218), .B(new_n13421), .Y(new_n20219));
  or_5   g17871(.A(new_n20218), .B(new_n13421), .Y(new_n20220));
  nand_5 g17872(.A(new_n20193), .B(new_n20192), .Y(new_n20221));
  xor_4  g17873(.A(new_n20221), .B(new_n20205), .Y(new_n20222));
  nand_5 g17874(.A(new_n20222), .B(new_n13429), .Y(new_n20223));
  or_5   g17875(.A(new_n20222), .B(new_n13429), .Y(new_n20224));
  nand_5 g17876(.A(new_n20196), .B(new_n20195), .Y(new_n20225));
  xor_4  g17877(.A(new_n20225), .B(new_n20203), .Y(new_n20226));
  nand_5 g17878(.A(new_n20226), .B(new_n13436), .Y(new_n20227));
  or_5   g17879(.A(new_n20226), .B(new_n13436), .Y(new_n20228));
  nand_5 g17880(.A(new_n20199), .B(new_n20198), .Y(new_n20229));
  xor_4  g17881(.A(new_n20229), .B(new_n20201), .Y(new_n20230));
  nand_5 g17882(.A(new_n20230), .B(new_n13441), .Y(new_n20231));
  or_5   g17883(.A(new_n20230), .B(new_n13441), .Y(new_n20232));
  nand_5 g17884(.A(new_n4531), .B(new_n4486), .Y(new_n20233));
  nand_5 g17885(.A(new_n20233), .B(new_n4530), .Y(new_n20234));
  nand_5 g17886(.A(new_n20234), .B(new_n20232), .Y(new_n20235_1));
  nand_5 g17887(.A(new_n20235_1), .B(new_n20231), .Y(new_n20236));
  nand_5 g17888(.A(new_n20236), .B(new_n20228), .Y(new_n20237));
  nand_5 g17889(.A(new_n20237), .B(new_n20227), .Y(new_n20238));
  nand_5 g17890(.A(new_n20238), .B(new_n20224), .Y(new_n20239));
  nand_5 g17891(.A(new_n20239), .B(new_n20223), .Y(new_n20240));
  nand_5 g17892(.A(new_n20240), .B(new_n20220), .Y(new_n20241));
  nand_5 g17893(.A(new_n20241), .B(new_n20219), .Y(new_n20242));
  xor_4  g17894(.A(new_n20242), .B(new_n20216), .Y(n4478));
  nand_5 g17895(.A(new_n14275_1), .B(new_n14276), .Y(new_n20244));
  xor_4  g17896(.A(new_n20244), .B(new_n14317), .Y(n4529));
  nand_5 g17897(.A(new_n6928), .B(new_n6926), .Y(new_n20246));
  xnor_4 g17898(.A(new_n20246), .B(new_n6984), .Y(n4552));
  not_8  g17899(.A(new_n6941), .Y(new_n20248));
  nand_5 g17900(.A(new_n20248), .B(new_n6940), .Y(new_n20249));
  xor_4  g17901(.A(new_n20249), .B(new_n6980), .Y(n4595));
  nand_5 g17902(.A(new_n16201), .B(new_n16200), .Y(new_n20251));
  xor_4  g17903(.A(new_n20251), .B(new_n16249), .Y(n4624));
  nor_5  g17904(.A(new_n19708), .B(n2659), .Y(new_n20253));
  nand_5 g17905(.A(new_n20253), .B(new_n5502), .Y(new_n20254));
  xor_4  g17906(.A(new_n20254), .B(n3740), .Y(new_n20255));
  nor_5  g17907(.A(new_n20255), .B(n3506), .Y(new_n20256));
  xor_4  g17908(.A(new_n20253), .B(new_n5502), .Y(new_n20257));
  or_5   g17909(.A(new_n20257), .B(n14899), .Y(new_n20258));
  nand_5 g17910(.A(new_n20257), .B(n14899), .Y(new_n20259_1));
  nand_5 g17911(.A(new_n19711), .B(new_n19707), .Y(new_n20260));
  nand_5 g17912(.A(new_n20260), .B(new_n19710), .Y(new_n20261));
  nand_5 g17913(.A(new_n20261), .B(new_n20259_1), .Y(new_n20262));
  nand_5 g17914(.A(new_n20262), .B(new_n20258), .Y(new_n20263));
  nor_5  g17915(.A(new_n20263), .B(new_n20256), .Y(new_n20264));
  or_5   g17916(.A(new_n20254), .B(n3740), .Y(new_n20265));
  nand_5 g17917(.A(new_n20255), .B(n3506), .Y(new_n20266));
  nand_5 g17918(.A(new_n20266), .B(new_n20265), .Y(new_n20267));
  nor_5  g17919(.A(new_n20267), .B(new_n20264), .Y(new_n20268));
  nor_5  g17920(.A(new_n20268), .B(new_n8796), .Y(new_n20269));
  nand_5 g17921(.A(new_n20268), .B(new_n8796), .Y(new_n20270));
  not_8  g17922(.A(new_n20270), .Y(new_n20271));
  nor_5  g17923(.A(new_n20271), .B(new_n20269), .Y(new_n20272));
  xor_4  g17924(.A(new_n20255), .B(n3506), .Y(new_n20273));
  xor_4  g17925(.A(new_n20273), .B(new_n20263), .Y(new_n20274));
  nand_5 g17926(.A(new_n20274), .B(new_n8849_1), .Y(new_n20275));
  or_5   g17927(.A(new_n20274), .B(new_n8849_1), .Y(new_n20276));
  nand_5 g17928(.A(new_n20259_1), .B(new_n20258), .Y(new_n20277));
  xor_4  g17929(.A(new_n20277), .B(new_n20261), .Y(new_n20278));
  or_5   g17930(.A(new_n20278), .B(new_n8858), .Y(new_n20279_1));
  nand_5 g17931(.A(new_n20278), .B(new_n8858), .Y(new_n20280));
  nand_5 g17932(.A(new_n19715), .B(new_n19705), .Y(new_n20281));
  nand_5 g17933(.A(new_n20281), .B(new_n19714), .Y(new_n20282));
  nand_5 g17934(.A(new_n20282), .B(new_n20280), .Y(new_n20283));
  nand_5 g17935(.A(new_n20283), .B(new_n20279_1), .Y(new_n20284));
  nand_5 g17936(.A(new_n20284), .B(new_n20276), .Y(new_n20285));
  nand_5 g17937(.A(new_n20285), .B(new_n20275), .Y(new_n20286));
  xor_4  g17938(.A(new_n20286), .B(new_n20272), .Y(new_n20287_1));
  not_8  g17939(.A(new_n20287_1), .Y(new_n20288));
  nand_5 g17940(.A(new_n20288), .B(new_n9011), .Y(new_n20289));
  nand_5 g17941(.A(new_n20287_1), .B(new_n9009), .Y(new_n20290));
  nand_5 g17942(.A(new_n20290), .B(new_n20289), .Y(new_n20291));
  nand_5 g17943(.A(new_n20276), .B(new_n20275), .Y(new_n20292));
  xor_4  g17944(.A(new_n20292), .B(new_n20284), .Y(new_n20293));
  not_8  g17945(.A(new_n20293), .Y(new_n20294));
  nand_5 g17946(.A(new_n20294), .B(new_n9019), .Y(new_n20295));
  nand_5 g17947(.A(new_n20293), .B(new_n9018), .Y(new_n20296));
  nand_5 g17948(.A(new_n20280), .B(new_n20279_1), .Y(new_n20297));
  xor_4  g17949(.A(new_n20297), .B(new_n20282), .Y(new_n20298));
  or_5   g17950(.A(new_n20298), .B(new_n9025), .Y(new_n20299));
  nand_5 g17951(.A(new_n20298), .B(new_n9025), .Y(new_n20300));
  or_5   g17952(.A(new_n19717), .B(new_n9031), .Y(new_n20301_1));
  nand_5 g17953(.A(new_n19717), .B(new_n9031), .Y(new_n20302));
  or_5   g17954(.A(new_n19690), .B(new_n9038), .Y(new_n20303));
  nand_5 g17955(.A(new_n19690), .B(new_n9038), .Y(new_n20304));
  nand_5 g17956(.A(new_n15227), .B(new_n9047_1), .Y(new_n20305));
  nand_5 g17957(.A(new_n15218), .B(new_n9046_1), .Y(new_n20306));
  nand_5 g17958(.A(new_n19529), .B(new_n19527), .Y(new_n20307));
  nand_5 g17959(.A(new_n20307), .B(new_n19528), .Y(new_n20308));
  nand_5 g17960(.A(new_n20308), .B(new_n20306), .Y(new_n20309));
  nand_5 g17961(.A(new_n20309), .B(new_n20305), .Y(new_n20310));
  nand_5 g17962(.A(new_n20310), .B(new_n20304), .Y(new_n20311));
  nand_5 g17963(.A(new_n20311), .B(new_n20303), .Y(new_n20312));
  nand_5 g17964(.A(new_n20312), .B(new_n20302), .Y(new_n20313));
  nand_5 g17965(.A(new_n20313), .B(new_n20301_1), .Y(new_n20314));
  nand_5 g17966(.A(new_n20314), .B(new_n20300), .Y(new_n20315));
  nand_5 g17967(.A(new_n20315), .B(new_n20299), .Y(new_n20316));
  nand_5 g17968(.A(new_n20316), .B(new_n20296), .Y(new_n20317));
  nand_5 g17969(.A(new_n20317), .B(new_n20295), .Y(new_n20318));
  xor_4  g17970(.A(new_n20318), .B(new_n20291), .Y(n4646));
  nand_5 g17971(.A(new_n16177), .B(new_n16176), .Y(new_n20320));
  xor_4  g17972(.A(new_n20320), .B(new_n16257), .Y(n4674));
  nand_5 g17973(.A(n20235), .B(new_n2383), .Y(new_n20322));
  nand_5 g17974(.A(new_n9765), .B(n11486), .Y(new_n20323));
  nand_5 g17975(.A(n13781), .B(new_n5669), .Y(new_n20324));
  nand_5 g17976(.A(new_n20324), .B(new_n20323), .Y(new_n20325));
  nand_5 g17977(.A(new_n20325), .B(new_n20322), .Y(new_n20326));
  nand_5 g17978(.A(new_n2394), .B(n8381), .Y(new_n20327));
  nand_5 g17979(.A(n16722), .B(new_n5709), .Y(new_n20328));
  nand_5 g17980(.A(new_n20328), .B(new_n20327), .Y(new_n20329));
  xor_4  g17981(.A(new_n20329), .B(new_n20326), .Y(new_n20330_1));
  nand_5 g17982(.A(new_n20330_1), .B(new_n3241), .Y(new_n20331));
  not_8  g17983(.A(new_n20331), .Y(new_n20332));
  or_5   g17984(.A(new_n20330_1), .B(new_n3241), .Y(new_n20333_1));
  not_8  g17985(.A(new_n20333_1), .Y(new_n20334));
  xor_4  g17986(.A(n13781), .B(new_n5669), .Y(new_n20335));
  nor_5  g17987(.A(new_n20335), .B(new_n3246), .Y(new_n20336));
  nand_5 g17988(.A(new_n20336), .B(new_n3258), .Y(new_n20337));
  or_5   g17989(.A(new_n20336), .B(new_n3258), .Y(new_n20338));
  nand_5 g17990(.A(new_n20323), .B(new_n20322), .Y(new_n20339));
  xnor_4 g17991(.A(new_n20339), .B(new_n20324), .Y(new_n20340));
  nand_5 g17992(.A(new_n20340), .B(new_n20338), .Y(new_n20341));
  nand_5 g17993(.A(new_n20341), .B(new_n20337), .Y(new_n20342));
  nor_5  g17994(.A(new_n20342), .B(new_n20334), .Y(new_n20343));
  nor_5  g17995(.A(new_n20343), .B(new_n20332), .Y(new_n20344));
  nand_5 g17996(.A(new_n20328), .B(new_n20326), .Y(new_n20345));
  nand_5 g17997(.A(new_n20345), .B(new_n20327), .Y(new_n20346));
  not_8  g17998(.A(new_n20346), .Y(new_n20347));
  nand_5 g17999(.A(n7057), .B(new_n2401), .Y(new_n20348));
  nand_5 g18000(.A(new_n9760), .B(n3480), .Y(new_n20349_1));
  nand_5 g18001(.A(new_n20349_1), .B(new_n20348), .Y(new_n20350));
  xor_4  g18002(.A(new_n20350), .B(new_n20347), .Y(new_n20351));
  or_5   g18003(.A(new_n20351), .B(new_n3233), .Y(new_n20352));
  not_8  g18004(.A(new_n20352), .Y(new_n20353));
  nand_5 g18005(.A(new_n20351), .B(new_n3233), .Y(new_n20354));
  not_8  g18006(.A(new_n20354), .Y(new_n20355_1));
  nor_5  g18007(.A(new_n20355_1), .B(new_n20353), .Y(new_n20356));
  xor_4  g18008(.A(new_n20356), .B(new_n20344), .Y(n4693));
  nand_5 g18009(.A(new_n12286), .B(new_n12287), .Y(new_n20358));
  xor_4  g18010(.A(new_n20358), .B(new_n12296), .Y(n4731));
  nand_5 g18011(.A(new_n6841), .B(new_n6794_1), .Y(new_n20360));
  nand_5 g18012(.A(new_n20360), .B(new_n6797), .Y(new_n20361));
  nand_5 g18013(.A(new_n6910), .B(new_n6845), .Y(new_n20362));
  nand_5 g18014(.A(new_n20362), .B(new_n6847), .Y(new_n20363));
  nor_5  g18015(.A(new_n20363), .B(new_n20361), .Y(new_n20364));
  not_8  g18016(.A(new_n20364), .Y(new_n20365));
  nand_5 g18017(.A(new_n20365), .B(new_n17557_1), .Y(new_n20366_1));
  nand_5 g18018(.A(new_n20364), .B(new_n17556), .Y(new_n20367));
  nand_5 g18019(.A(new_n20367), .B(new_n20366_1), .Y(new_n20368));
  nand_5 g18020(.A(new_n20363), .B(new_n20361), .Y(new_n20369));
  and_5  g18021(.A(new_n20369), .B(new_n20365), .Y(new_n20370));
  not_8  g18022(.A(new_n20370), .Y(new_n20371));
  nand_5 g18023(.A(new_n20371), .B(new_n17573), .Y(new_n20372));
  or_5   g18024(.A(new_n20371), .B(new_n17573), .Y(new_n20373));
  nand_5 g18025(.A(new_n14796), .B(new_n14749), .Y(new_n20374));
  nand_5 g18026(.A(new_n20374), .B(new_n14752), .Y(new_n20375));
  nand_5 g18027(.A(new_n20375), .B(new_n20373), .Y(new_n20376));
  nand_5 g18028(.A(new_n20376), .B(new_n20372), .Y(new_n20377));
  xor_4  g18029(.A(new_n20377), .B(new_n20368), .Y(n4745));
  xor_4  g18030(.A(new_n7142), .B(n6773), .Y(new_n20379));
  nor_5  g18031(.A(new_n20379), .B(new_n12609), .Y(new_n20380));
  not_8  g18032(.A(new_n20380), .Y(new_n20381));
  nand_5 g18033(.A(new_n20379), .B(new_n12609), .Y(new_n20382));
  nand_5 g18034(.A(new_n20382), .B(new_n20381), .Y(n4747));
  nand_5 g18035(.A(new_n6492), .B(new_n6491), .Y(new_n20384));
  xor_4  g18036(.A(new_n20384), .B(new_n6494), .Y(n4766));
  nand_5 g18037(.A(new_n15639), .B(new_n15638), .Y(new_n20386));
  xnor_4 g18038(.A(new_n20386), .B(new_n15660), .Y(n4770));
  xor_4  g18039(.A(new_n18770), .B(new_n17818), .Y(n4777));
  nand_5 g18040(.A(new_n6405), .B(n2328), .Y(new_n20389));
  nand_5 g18041(.A(n7731), .B(new_n3547), .Y(new_n20390));
  nand_5 g18042(.A(n15053), .B(new_n6408), .Y(new_n20391));
  nand_5 g18043(.A(new_n3549), .B(n12341), .Y(new_n20392));
  nand_5 g18044(.A(n25471), .B(new_n6411), .Y(new_n20393));
  nand_5 g18045(.A(new_n3553), .B(n20986), .Y(new_n20394));
  nand_5 g18046(.A(new_n3653), .B(n12384), .Y(new_n20395));
  nand_5 g18047(.A(new_n20395), .B(new_n20394), .Y(new_n20396));
  nand_5 g18048(.A(new_n20396), .B(new_n20393), .Y(new_n20397));
  nand_5 g18049(.A(new_n20397), .B(new_n20392), .Y(new_n20398));
  nand_5 g18050(.A(new_n20398), .B(new_n20391), .Y(new_n20399));
  nand_5 g18051(.A(new_n20399), .B(new_n20390), .Y(new_n20400));
  nand_5 g18052(.A(new_n20400), .B(new_n20389), .Y(new_n20401));
  nand_5 g18053(.A(n19357), .B(new_n6402), .Y(new_n20402_1));
  nand_5 g18054(.A(new_n18176), .B(n7566), .Y(new_n20403_1));
  nand_5 g18055(.A(new_n20403_1), .B(new_n20402_1), .Y(new_n20404));
  xor_4  g18056(.A(new_n20404), .B(new_n20401), .Y(new_n20405));
  nand_5 g18057(.A(new_n2358), .B(new_n2442), .Y(new_n20406));
  xor_4  g18058(.A(new_n20406), .B(n15636), .Y(new_n20407));
  nand_5 g18059(.A(new_n20407), .B(new_n6205), .Y(new_n20408));
  or_5   g18060(.A(new_n20407), .B(new_n6205), .Y(new_n20409_1));
  nand_5 g18061(.A(n20077), .B(n6794), .Y(new_n20410));
  and_5  g18062(.A(new_n20410), .B(new_n20406), .Y(new_n20411_1));
  nand_5 g18063(.A(new_n20411_1), .B(new_n10338), .Y(new_n20412));
  or_5   g18064(.A(new_n20411_1), .B(new_n10338), .Y(new_n20413));
  nand_5 g18065(.A(new_n2442), .B(n6611), .Y(new_n20414));
  nand_5 g18066(.A(new_n20414), .B(new_n20413), .Y(new_n20415));
  nand_5 g18067(.A(new_n20415), .B(new_n20412), .Y(new_n20416));
  nand_5 g18068(.A(new_n20416), .B(new_n20409_1), .Y(new_n20417));
  nand_5 g18069(.A(new_n20417), .B(new_n20408), .Y(new_n20418));
  or_5   g18070(.A(new_n20406), .B(n15636), .Y(new_n20419));
  xor_4  g18071(.A(new_n20419), .B(n8745), .Y(new_n20420));
  nand_5 g18072(.A(new_n20420), .B(new_n10333), .Y(new_n20421));
  or_5   g18073(.A(new_n20420), .B(new_n10333), .Y(new_n20422));
  nand_5 g18074(.A(new_n20422), .B(new_n20421), .Y(new_n20423));
  xor_4  g18075(.A(new_n20423), .B(new_n20418), .Y(new_n20424_1));
  nand_5 g18076(.A(new_n20424_1), .B(new_n17455), .Y(new_n20425));
  nor_5  g18077(.A(new_n20424_1), .B(new_n17455), .Y(new_n20426));
  nand_5 g18078(.A(new_n20409_1), .B(new_n20408), .Y(new_n20427));
  xor_4  g18079(.A(new_n20427), .B(new_n20416), .Y(new_n20428));
  nand_5 g18080(.A(new_n20428), .B(new_n5716), .Y(new_n20429_1));
  not_8  g18081(.A(new_n20429_1), .Y(new_n20430));
  not_8  g18082(.A(new_n20428), .Y(new_n20431));
  nand_5 g18083(.A(new_n20431), .B(new_n5717), .Y(new_n20432));
  not_8  g18084(.A(new_n20432), .Y(new_n20433));
  nand_5 g18085(.A(new_n20413), .B(new_n20412), .Y(new_n20434));
  xnor_4 g18086(.A(new_n20434), .B(new_n20414), .Y(new_n20435));
  nand_5 g18087(.A(new_n20435), .B(new_n5668), .Y(new_n20436_1));
  nor_5  g18088(.A(new_n20435), .B(new_n5668), .Y(new_n20437));
  not_8  g18089(.A(new_n20437), .Y(new_n20438));
  nand_5 g18090(.A(n6794), .B(new_n6339_1), .Y(new_n20439));
  and_5  g18091(.A(new_n20439), .B(new_n20414), .Y(new_n20440));
  not_8  g18092(.A(new_n20440), .Y(new_n20441_1));
  nand_5 g18093(.A(new_n20441_1), .B(new_n5671), .Y(new_n20442));
  not_8  g18094(.A(new_n20442), .Y(new_n20443));
  nand_5 g18095(.A(new_n20443), .B(new_n20438), .Y(new_n20444));
  nand_5 g18096(.A(new_n20444), .B(new_n20436_1), .Y(new_n20445_1));
  nor_5  g18097(.A(new_n20445_1), .B(new_n20433), .Y(new_n20446));
  nor_5  g18098(.A(new_n20446), .B(new_n20430), .Y(new_n20447));
  or_5   g18099(.A(new_n20447), .B(new_n20426), .Y(new_n20448));
  nand_5 g18100(.A(new_n20448), .B(new_n20425), .Y(new_n20449));
  nand_5 g18101(.A(new_n20422), .B(new_n20418), .Y(new_n20450_1));
  nand_5 g18102(.A(new_n20450_1), .B(new_n20421), .Y(new_n20451));
  nor_5  g18103(.A(new_n20419), .B(n8745), .Y(new_n20452));
  xor_4  g18104(.A(new_n20452), .B(n1777), .Y(new_n20453));
  or_5   g18105(.A(new_n20453), .B(n15884), .Y(new_n20454));
  nand_5 g18106(.A(new_n20453), .B(n15884), .Y(new_n20455_1));
  nand_5 g18107(.A(new_n20455_1), .B(new_n20454), .Y(new_n20456));
  xor_4  g18108(.A(new_n20456), .B(new_n20451), .Y(new_n20457));
  nand_5 g18109(.A(new_n20457), .B(new_n17499), .Y(new_n20458));
  or_5   g18110(.A(new_n20457), .B(new_n17499), .Y(new_n20459));
  nand_5 g18111(.A(new_n20459), .B(new_n20458), .Y(new_n20460));
  xor_4  g18112(.A(new_n20460), .B(new_n20449), .Y(new_n20461));
  not_8  g18113(.A(new_n20461), .Y(new_n20462));
  or_5   g18114(.A(new_n20462), .B(new_n20405), .Y(new_n20463));
  nand_5 g18115(.A(new_n20462), .B(new_n20405), .Y(new_n20464));
  nand_5 g18116(.A(new_n20390), .B(new_n20389), .Y(new_n20465));
  xor_4  g18117(.A(new_n20465), .B(new_n20399), .Y(new_n20466));
  xor_4  g18118(.A(new_n20424_1), .B(new_n17455), .Y(new_n20467));
  xor_4  g18119(.A(new_n20467), .B(new_n20447), .Y(new_n20468));
  not_8  g18120(.A(new_n20468), .Y(new_n20469));
  or_5   g18121(.A(new_n20469), .B(new_n20466), .Y(new_n20470_1));
  nand_5 g18122(.A(new_n20469), .B(new_n20466), .Y(new_n20471));
  nand_5 g18123(.A(new_n20392), .B(new_n20391), .Y(new_n20472));
  xor_4  g18124(.A(new_n20472), .B(new_n20397), .Y(new_n20473));
  nand_5 g18125(.A(new_n20432), .B(new_n20429_1), .Y(new_n20474));
  xor_4  g18126(.A(new_n20474), .B(new_n20445_1), .Y(new_n20475));
  or_5   g18127(.A(new_n20475), .B(new_n20473), .Y(new_n20476));
  nand_5 g18128(.A(new_n20475), .B(new_n20473), .Y(new_n20477));
  nor_5  g18129(.A(new_n20441_1), .B(new_n5671), .Y(new_n20478_1));
  nor_5  g18130(.A(new_n20478_1), .B(new_n20443), .Y(new_n20479));
  nand_5 g18131(.A(n16502), .B(new_n6413), .Y(new_n20480));
  nand_5 g18132(.A(new_n20480), .B(new_n20395), .Y(new_n20481));
  nand_5 g18133(.A(new_n20481), .B(new_n20479), .Y(new_n20482));
  not_8  g18134(.A(new_n20395), .Y(new_n20483));
  and_5  g18135(.A(new_n20394), .B(new_n20393), .Y(new_n20484));
  xor_4  g18136(.A(new_n20484), .B(new_n20483), .Y(new_n20485));
  or_5   g18137(.A(new_n20485), .B(new_n20482), .Y(new_n20486));
  nand_5 g18138(.A(new_n20485), .B(new_n20482), .Y(new_n20487));
  nand_5 g18139(.A(new_n20438), .B(new_n20436_1), .Y(new_n20488));
  xor_4  g18140(.A(new_n20488), .B(new_n20443), .Y(new_n20489_1));
  not_8  g18141(.A(new_n20489_1), .Y(new_n20490_1));
  nand_5 g18142(.A(new_n20490_1), .B(new_n20487), .Y(new_n20491));
  nand_5 g18143(.A(new_n20491), .B(new_n20486), .Y(new_n20492));
  nand_5 g18144(.A(new_n20492), .B(new_n20477), .Y(new_n20493));
  nand_5 g18145(.A(new_n20493), .B(new_n20476), .Y(new_n20494));
  nand_5 g18146(.A(new_n20494), .B(new_n20471), .Y(new_n20495_1));
  nand_5 g18147(.A(new_n20495_1), .B(new_n20470_1), .Y(new_n20496));
  nand_5 g18148(.A(new_n20496), .B(new_n20464), .Y(new_n20497));
  nand_5 g18149(.A(new_n20497), .B(new_n20463), .Y(new_n20498));
  nand_5 g18150(.A(new_n20459), .B(new_n20449), .Y(new_n20499));
  nand_5 g18151(.A(new_n20499), .B(new_n20458), .Y(new_n20500));
  nand_5 g18152(.A(new_n20455_1), .B(new_n20451), .Y(new_n20501));
  nand_5 g18153(.A(new_n20501), .B(new_n20454), .Y(new_n20502));
  nand_5 g18154(.A(new_n20452), .B(new_n2370), .Y(new_n20503));
  not_8  g18155(.A(new_n20503), .Y(new_n20504));
  nand_5 g18156(.A(new_n20504), .B(new_n2467), .Y(new_n20505));
  nand_5 g18157(.A(new_n20503), .B(n22660), .Y(new_n20506));
  nand_5 g18158(.A(new_n20506), .B(new_n20505), .Y(new_n20507));
  or_5   g18159(.A(new_n20507), .B(n11580), .Y(new_n20508));
  nand_5 g18160(.A(new_n20507), .B(n11580), .Y(new_n20509));
  nand_5 g18161(.A(new_n20509), .B(new_n20508), .Y(new_n20510));
  xor_4  g18162(.A(new_n20510), .B(new_n20502), .Y(new_n20511));
  nand_5 g18163(.A(new_n20511), .B(new_n18147), .Y(new_n20512));
  or_5   g18164(.A(new_n20511), .B(new_n18147), .Y(new_n20513));
  nand_5 g18165(.A(new_n20513), .B(new_n20512), .Y(new_n20514));
  xor_4  g18166(.A(new_n20514), .B(new_n20500), .Y(new_n20515_1));
  nand_5 g18167(.A(new_n20403_1), .B(new_n20401), .Y(new_n20516));
  nand_5 g18168(.A(new_n20516), .B(new_n20402_1), .Y(new_n20517));
  nand_5 g18169(.A(new_n6399), .B(n6861), .Y(new_n20518));
  nand_5 g18170(.A(n17959), .B(new_n3546), .Y(new_n20519));
  nand_5 g18171(.A(new_n20519), .B(new_n20518), .Y(new_n20520));
  xnor_4 g18172(.A(new_n20520), .B(new_n20517), .Y(new_n20521));
  nand_5 g18173(.A(new_n20521), .B(new_n20515_1), .Y(new_n20522));
  or_5   g18174(.A(new_n20521), .B(new_n20515_1), .Y(new_n20523));
  nand_5 g18175(.A(new_n20523), .B(new_n20522), .Y(new_n20524));
  xnor_4 g18176(.A(new_n20524), .B(new_n20498), .Y(n4785));
  nor_5  g18177(.A(new_n15972), .B(new_n15971), .Y(new_n20526));
  xor_4  g18178(.A(new_n20526), .B(new_n16011), .Y(n4804));
  nand_5 g18179(.A(new_n17800), .B(new_n17799), .Y(new_n20528));
  xor_4  g18180(.A(new_n20528), .B(new_n17826), .Y(n4810));
  xor_4  g18181(.A(new_n19995), .B(new_n12409), .Y(new_n20530));
  xor_4  g18182(.A(new_n20530), .B(new_n9149), .Y(new_n20531));
  nand_5 g18183(.A(new_n12465), .B(new_n12413), .Y(new_n20532));
  nand_5 g18184(.A(new_n20532), .B(new_n12412), .Y(new_n20533_1));
  xor_4  g18185(.A(new_n20533_1), .B(new_n20531), .Y(new_n20534));
  nand_5 g18186(.A(new_n10509), .B(new_n10469), .Y(new_n20535));
  nand_5 g18187(.A(new_n20535), .B(new_n10470), .Y(new_n20536));
  or_5   g18188(.A(new_n20536), .B(new_n20534), .Y(new_n20537));
  nand_5 g18189(.A(new_n20536), .B(new_n20534), .Y(new_n20538));
  nand_5 g18190(.A(new_n12523), .B(new_n12468), .Y(new_n20539));
  nand_5 g18191(.A(new_n20539), .B(new_n12467_1), .Y(new_n20540));
  nand_5 g18192(.A(new_n20540), .B(new_n20538), .Y(new_n20541));
  nand_5 g18193(.A(new_n20541), .B(new_n20537), .Y(new_n20542));
  not_8  g18194(.A(new_n20542), .Y(new_n20543));
  nand_5 g18195(.A(new_n20530), .B(new_n9149), .Y(new_n20544));
  nand_5 g18196(.A(new_n20533_1), .B(new_n20544), .Y(new_n20545));
  nor_5  g18197(.A(new_n19996), .B(new_n12409), .Y(new_n20546));
  nor_5  g18198(.A(new_n20530), .B(new_n9149), .Y(new_n20547));
  nor_5  g18199(.A(new_n20547), .B(new_n20546), .Y(new_n20548));
  nand_5 g18200(.A(new_n20548), .B(new_n20545), .Y(new_n20549));
  nand_5 g18201(.A(new_n20549), .B(new_n20543), .Y(n4814));
  nand_5 g18202(.A(new_n18533), .B(new_n18531), .Y(new_n20551));
  xnor_4 g18203(.A(new_n20551), .B(new_n18537_1), .Y(n4850));
  nand_5 g18204(.A(new_n19444), .B(new_n19442), .Y(new_n20553));
  xnor_4 g18205(.A(new_n20553), .B(new_n19496_1), .Y(n4891));
  nor_5  g18206(.A(new_n19644), .B(new_n19643), .Y(new_n20555));
  xor_4  g18207(.A(new_n20555), .B(new_n19670), .Y(n4925));
  nand_5 g18208(.A(new_n18517), .B(new_n18516), .Y(new_n20557));
  xnor_4 g18209(.A(new_n20557), .B(new_n18543), .Y(n4947));
  not_8  g18210(.A(new_n10803), .Y(new_n20559));
  xor_4  g18211(.A(new_n10806), .B(new_n20559), .Y(n4952));
  or_5   g18212(.A(new_n9193), .B(n5882), .Y(new_n20561));
  nand_5 g18213(.A(new_n9193), .B(n5882), .Y(new_n20562));
  or_5   g18214(.A(new_n9981), .B(n11775), .Y(new_n20563));
  nand_5 g18215(.A(new_n9981), .B(n11775), .Y(new_n20564));
  nand_5 g18216(.A(new_n20564), .B(new_n17148), .Y(new_n20565));
  nand_5 g18217(.A(new_n20565), .B(new_n20563), .Y(new_n20566));
  nand_5 g18218(.A(new_n20566), .B(new_n20562), .Y(new_n20567));
  nand_5 g18219(.A(new_n20567), .B(new_n20561), .Y(new_n20568));
  nand_5 g18220(.A(n22631), .B(new_n11365), .Y(new_n20569));
  nand_5 g18221(.A(new_n9187), .B(n2117), .Y(new_n20570));
  nand_5 g18222(.A(new_n20570), .B(new_n20569), .Y(new_n20571));
  xor_4  g18223(.A(new_n20571), .B(new_n20568), .Y(new_n20572));
  or_5   g18224(.A(new_n20572), .B(new_n17386), .Y(new_n20573));
  nand_5 g18225(.A(new_n20572), .B(new_n17386), .Y(new_n20574));
  nand_5 g18226(.A(new_n20562), .B(new_n20561), .Y(new_n20575));
  xor_4  g18227(.A(new_n20575), .B(new_n20566), .Y(new_n20576));
  or_5   g18228(.A(new_n20576), .B(new_n17391_1), .Y(new_n20577));
  nand_5 g18229(.A(new_n20576), .B(new_n17391_1), .Y(new_n20578));
  nand_5 g18230(.A(new_n20564), .B(new_n20563), .Y(new_n20579));
  xnor_4 g18231(.A(new_n20579), .B(new_n17148), .Y(new_n20580));
  nand_5 g18232(.A(new_n20580), .B(new_n17395), .Y(new_n20581));
  nor_5  g18233(.A(new_n20580), .B(new_n17395), .Y(new_n20582_1));
  not_8  g18234(.A(new_n20582_1), .Y(new_n20583));
  nand_5 g18235(.A(new_n20583), .B(new_n17153), .Y(new_n20584));
  nand_5 g18236(.A(new_n20584), .B(new_n20581), .Y(new_n20585));
  nand_5 g18237(.A(new_n20585), .B(new_n20578), .Y(new_n20586));
  nand_5 g18238(.A(new_n20586), .B(new_n20577), .Y(new_n20587));
  nand_5 g18239(.A(new_n20587), .B(new_n20574), .Y(new_n20588));
  nand_5 g18240(.A(new_n20588), .B(new_n20573), .Y(new_n20589));
  nand_5 g18241(.A(new_n20570), .B(new_n20568), .Y(new_n20590_1));
  nand_5 g18242(.A(new_n20590_1), .B(new_n20569), .Y(new_n20591));
  nand_5 g18243(.A(new_n11360), .B(n2331), .Y(new_n20592));
  nand_5 g18244(.A(n22879), .B(new_n9181), .Y(new_n20593));
  nand_5 g18245(.A(new_n20593), .B(new_n20592), .Y(new_n20594));
  xor_4  g18246(.A(new_n20594), .B(new_n20591), .Y(new_n20595));
  or_5   g18247(.A(new_n20595), .B(new_n17378), .Y(new_n20596));
  nand_5 g18248(.A(new_n20595), .B(new_n17378), .Y(new_n20597));
  nand_5 g18249(.A(new_n20597), .B(new_n20596), .Y(new_n20598));
  xor_4  g18250(.A(new_n20598), .B(new_n20589), .Y(new_n20599));
  or_5   g18251(.A(new_n20599), .B(new_n17344_1), .Y(new_n20600));
  nand_5 g18252(.A(new_n20599), .B(new_n17344_1), .Y(new_n20601));
  nand_5 g18253(.A(new_n20574), .B(new_n20573), .Y(new_n20602_1));
  xor_4  g18254(.A(new_n20602_1), .B(new_n20587), .Y(new_n20603));
  or_5   g18255(.A(new_n20603), .B(new_n15559_1), .Y(new_n20604_1));
  nand_5 g18256(.A(new_n20603), .B(new_n15559_1), .Y(new_n20605));
  nand_5 g18257(.A(new_n20578), .B(new_n20577), .Y(new_n20606));
  xor_4  g18258(.A(new_n20606), .B(new_n20585), .Y(new_n20607));
  not_8  g18259(.A(new_n20607), .Y(new_n20608));
  nand_5 g18260(.A(new_n20608), .B(new_n15500), .Y(new_n20609_1));
  nand_5 g18261(.A(new_n20607), .B(new_n15509), .Y(new_n20610));
  nand_5 g18262(.A(new_n17157), .B(new_n15493), .Y(new_n20611));
  or_5   g18263(.A(new_n17157), .B(new_n15493), .Y(new_n20612));
  nand_5 g18264(.A(new_n20583), .B(new_n20581), .Y(new_n20613));
  xor_4  g18265(.A(new_n20613), .B(new_n17153), .Y(new_n20614));
  not_8  g18266(.A(new_n20614), .Y(new_n20615));
  nand_5 g18267(.A(new_n20615), .B(new_n20612), .Y(new_n20616));
  nand_5 g18268(.A(new_n20616), .B(new_n20611), .Y(new_n20617));
  nand_5 g18269(.A(new_n20617), .B(new_n20610), .Y(new_n20618));
  nand_5 g18270(.A(new_n20618), .B(new_n20609_1), .Y(new_n20619));
  nand_5 g18271(.A(new_n20619), .B(new_n20605), .Y(new_n20620));
  nand_5 g18272(.A(new_n20620), .B(new_n20604_1), .Y(new_n20621));
  nand_5 g18273(.A(new_n20621), .B(new_n20601), .Y(new_n20622));
  nand_5 g18274(.A(new_n20622), .B(new_n20600), .Y(new_n20623_1));
  nand_5 g18275(.A(new_n20597), .B(new_n20589), .Y(new_n20624));
  nand_5 g18276(.A(new_n20624), .B(new_n20596), .Y(new_n20625));
  nand_5 g18277(.A(new_n20593), .B(new_n20591), .Y(new_n20626));
  nand_5 g18278(.A(new_n20626), .B(new_n20592), .Y(new_n20627));
  nand_5 g18279(.A(n25068), .B(new_n11355), .Y(new_n20628));
  nand_5 g18280(.A(new_n9175), .B(n6790), .Y(new_n20629_1));
  nand_5 g18281(.A(new_n20629_1), .B(new_n20628), .Y(new_n20630));
  xnor_4 g18282(.A(new_n20630), .B(new_n20627), .Y(new_n20631));
  nand_5 g18283(.A(new_n20631), .B(new_n17369), .Y(new_n20632));
  or_5   g18284(.A(new_n20631), .B(new_n17369), .Y(new_n20633));
  nand_5 g18285(.A(new_n20633), .B(new_n20632), .Y(new_n20634));
  xor_4  g18286(.A(new_n20634), .B(new_n20625), .Y(new_n20635));
  not_8  g18287(.A(new_n20635), .Y(new_n20636));
  nand_5 g18288(.A(new_n20636), .B(new_n17340), .Y(new_n20637));
  nand_5 g18289(.A(new_n20635), .B(new_n17342), .Y(new_n20638));
  nand_5 g18290(.A(new_n20638), .B(new_n20637), .Y(new_n20639));
  xnor_4 g18291(.A(new_n20639), .B(new_n20623_1), .Y(n4966));
  nand_5 g18292(.A(new_n20029), .B(new_n20028), .Y(new_n20641));
  xor_4  g18293(.A(new_n20641), .B(new_n20037), .Y(n4972));
  nand_5 g18294(.A(new_n8619), .B(new_n6384), .Y(new_n20643));
  or_5   g18295(.A(new_n8619), .B(new_n6384), .Y(new_n20644));
  nand_5 g18296(.A(new_n8625), .B(new_n6388), .Y(new_n20645));
  or_5   g18297(.A(new_n8625), .B(new_n6388), .Y(new_n20646));
  nand_5 g18298(.A(new_n19321), .B(new_n19318), .Y(new_n20647));
  nand_5 g18299(.A(new_n20647), .B(new_n19320), .Y(new_n20648));
  nand_5 g18300(.A(new_n20648), .B(new_n20646), .Y(new_n20649));
  nand_5 g18301(.A(new_n20649), .B(new_n20645), .Y(new_n20650));
  nand_5 g18302(.A(new_n20650), .B(new_n20644), .Y(new_n20651));
  nand_5 g18303(.A(new_n20651), .B(new_n20643), .Y(new_n20652));
  not_8  g18304(.A(new_n20652), .Y(new_n20653));
  nand_5 g18305(.A(new_n20653), .B(new_n8611), .Y(new_n20654));
  nand_5 g18306(.A(new_n19304), .B(new_n7958), .Y(new_n20655));
  nand_5 g18307(.A(new_n20655), .B(n2978), .Y(new_n20656));
  nor_5  g18308(.A(new_n20655), .B(n2978), .Y(new_n20657));
  not_8  g18309(.A(new_n20657), .Y(new_n20658_1));
  and_5  g18310(.A(new_n20658_1), .B(new_n20656), .Y(new_n20659));
  not_8  g18311(.A(new_n20659), .Y(new_n20660));
  nand_5 g18312(.A(new_n20660), .B(new_n3542), .Y(new_n20661_1));
  not_8  g18313(.A(new_n20661_1), .Y(new_n20662));
  nand_5 g18314(.A(new_n19305), .B(n23697), .Y(new_n20663));
  and_5  g18315(.A(new_n20663), .B(new_n20655), .Y(new_n20664));
  or_5   g18316(.A(new_n20664), .B(n337), .Y(new_n20665));
  nand_5 g18317(.A(new_n20664), .B(n337), .Y(new_n20666));
  nand_5 g18318(.A(new_n19310), .B(new_n19302), .Y(new_n20667));
  nand_5 g18319(.A(new_n20667), .B(new_n19309), .Y(new_n20668));
  nand_5 g18320(.A(new_n20668), .B(new_n20666), .Y(new_n20669));
  nand_5 g18321(.A(new_n20669), .B(new_n20665), .Y(new_n20670));
  nor_5  g18322(.A(new_n20670), .B(new_n20662), .Y(new_n20671));
  nand_5 g18323(.A(new_n20659), .B(n7593), .Y(new_n20672));
  nand_5 g18324(.A(new_n20672), .B(new_n20658_1), .Y(new_n20673_1));
  nor_5  g18325(.A(new_n20673_1), .B(new_n20671), .Y(new_n20674));
  not_8  g18326(.A(new_n20674), .Y(new_n20675));
  nand_5 g18327(.A(new_n20672), .B(new_n20661_1), .Y(new_n20676));
  xor_4  g18328(.A(new_n20676), .B(new_n20670), .Y(new_n20677));
  not_8  g18329(.A(new_n20677), .Y(new_n20678_1));
  nand_5 g18330(.A(new_n20678_1), .B(new_n9943), .Y(new_n20679));
  nand_5 g18331(.A(new_n20677), .B(n25972), .Y(new_n20680_1));
  nand_5 g18332(.A(new_n20666), .B(new_n20665), .Y(new_n20681));
  xor_4  g18333(.A(new_n20681), .B(new_n20668), .Y(new_n20682));
  not_8  g18334(.A(new_n20682), .Y(new_n20683));
  nand_5 g18335(.A(new_n20683), .B(new_n7974), .Y(new_n20684));
  nand_5 g18336(.A(new_n20682), .B(n21915), .Y(new_n20685_1));
  nand_5 g18337(.A(new_n19314_1), .B(new_n19300), .Y(new_n20686));
  nand_5 g18338(.A(new_n20686), .B(new_n19313), .Y(new_n20687));
  nand_5 g18339(.A(new_n20687), .B(new_n20685_1), .Y(new_n20688));
  nand_5 g18340(.A(new_n20688), .B(new_n20684), .Y(new_n20689));
  nand_5 g18341(.A(new_n20689), .B(new_n20680_1), .Y(new_n20690));
  nand_5 g18342(.A(new_n20690), .B(new_n20679), .Y(new_n20691_1));
  or_5   g18343(.A(new_n20691_1), .B(new_n20675), .Y(new_n20692));
  nand_5 g18344(.A(new_n20691_1), .B(new_n20675), .Y(new_n20693));
  and_5  g18345(.A(new_n20693), .B(new_n20692), .Y(new_n20694));
  nand_5 g18346(.A(new_n20652), .B(new_n8612), .Y(new_n20695));
  and_5  g18347(.A(new_n20695), .B(new_n20654), .Y(new_n20696_1));
  or_5   g18348(.A(new_n20696_1), .B(new_n20694), .Y(new_n20697));
  nand_5 g18349(.A(new_n20643), .B(new_n20644), .Y(new_n20698));
  xor_4  g18350(.A(new_n20698), .B(new_n20650), .Y(new_n20699));
  nand_5 g18351(.A(new_n20679), .B(new_n20680_1), .Y(new_n20700_1));
  xor_4  g18352(.A(new_n20700_1), .B(new_n20689), .Y(new_n20701));
  or_5   g18353(.A(new_n20701), .B(new_n20699), .Y(new_n20702));
  nand_5 g18354(.A(new_n20701), .B(new_n20699), .Y(new_n20703));
  nand_5 g18355(.A(new_n20645), .B(new_n20646), .Y(new_n20704_1));
  xor_4  g18356(.A(new_n20704_1), .B(new_n20648), .Y(new_n20705_1));
  nand_5 g18357(.A(new_n20684), .B(new_n20685_1), .Y(new_n20706));
  xor_4  g18358(.A(new_n20706), .B(new_n20687), .Y(new_n20707));
  or_5   g18359(.A(new_n20707), .B(new_n20705_1), .Y(new_n20708));
  nand_5 g18360(.A(new_n20707), .B(new_n20705_1), .Y(new_n20709_1));
  nand_5 g18361(.A(new_n19326), .B(new_n19298), .Y(new_n20710));
  nand_5 g18362(.A(new_n20710), .B(new_n19325), .Y(new_n20711));
  nand_5 g18363(.A(new_n20711), .B(new_n20709_1), .Y(new_n20712));
  nand_5 g18364(.A(new_n20712), .B(new_n20708), .Y(new_n20713_1));
  nand_5 g18365(.A(new_n20713_1), .B(new_n20703), .Y(new_n20714));
  nand_5 g18366(.A(new_n20714), .B(new_n20702), .Y(new_n20715));
  not_8  g18367(.A(new_n20715), .Y(new_n20716));
  nand_5 g18368(.A(new_n20716), .B(new_n20697), .Y(new_n20717));
  nor_5  g18369(.A(new_n20717), .B(new_n20692), .Y(new_n20718));
  not_8  g18370(.A(new_n20717), .Y(new_n20719));
  nand_5 g18371(.A(new_n20696_1), .B(new_n20694), .Y(new_n20720));
  nand_5 g18372(.A(new_n20720), .B(new_n20692), .Y(new_n20721));
  nor_5  g18373(.A(new_n20721), .B(new_n20719), .Y(new_n20722_1));
  nor_5  g18374(.A(new_n20722_1), .B(new_n20718), .Y(new_n20723_1));
  xor_4  g18375(.A(new_n20723_1), .B(new_n20654), .Y(n5011));
  nand_5 g18376(.A(new_n3289_1), .B(new_n3284), .Y(new_n20725));
  nand_5 g18377(.A(new_n20725), .B(new_n3288), .Y(new_n20726));
  or_5   g18378(.A(new_n20726), .B(new_n13565), .Y(new_n20727));
  nand_5 g18379(.A(new_n20727), .B(new_n10316), .Y(new_n20728));
  nand_5 g18380(.A(new_n20726), .B(new_n13565), .Y(new_n20729));
  nand_5 g18381(.A(new_n20729), .B(new_n20728), .Y(new_n20730));
  or_5   g18382(.A(new_n20730), .B(new_n17239), .Y(new_n20731));
  nand_5 g18383(.A(new_n20730), .B(new_n17239), .Y(new_n20732));
  nand_5 g18384(.A(new_n20732), .B(new_n20731), .Y(new_n20733));
  and_5  g18385(.A(new_n20729), .B(new_n20727), .Y(new_n20734));
  xor_4  g18386(.A(new_n20734), .B(new_n10316), .Y(new_n20735));
  nand_5 g18387(.A(new_n20735), .B(new_n17217), .Y(new_n20736));
  not_8  g18388(.A(new_n20735), .Y(new_n20737));
  nand_5 g18389(.A(new_n20737), .B(new_n17219_1), .Y(new_n20738));
  nand_5 g18390(.A(new_n3304), .B(new_n3281), .Y(new_n20739));
  nand_5 g18391(.A(new_n20739), .B(new_n3301_1), .Y(new_n20740));
  nand_5 g18392(.A(new_n20740), .B(new_n20738), .Y(new_n20741));
  nand_5 g18393(.A(new_n20741), .B(new_n20736), .Y(new_n20742));
  xor_4  g18394(.A(new_n20742), .B(new_n20733), .Y(new_n20743));
  nand_5 g18395(.A(n11220), .B(new_n2781), .Y(new_n20744));
  nand_5 g18396(.A(new_n11623), .B(n2944), .Y(new_n20745));
  nand_5 g18397(.A(new_n3277), .B(new_n3274), .Y(new_n20746));
  nand_5 g18398(.A(new_n20746), .B(new_n3275), .Y(new_n20747));
  nand_5 g18399(.A(new_n20747), .B(new_n20745), .Y(new_n20748_1));
  nand_5 g18400(.A(new_n20748_1), .B(new_n20744), .Y(new_n20749));
  not_8  g18401(.A(new_n20749), .Y(new_n20750));
  nand_5 g18402(.A(new_n20750), .B(new_n20743), .Y(new_n20751));
  or_5   g18403(.A(new_n20750), .B(new_n20743), .Y(new_n20752));
  nand_5 g18404(.A(new_n20745), .B(new_n20744), .Y(new_n20753));
  xor_4  g18405(.A(new_n20753), .B(new_n20747), .Y(new_n20754));
  nand_5 g18406(.A(new_n20736), .B(new_n20738), .Y(new_n20755));
  xor_4  g18407(.A(new_n20755), .B(new_n20740), .Y(new_n20756));
  not_8  g18408(.A(new_n20756), .Y(new_n20757));
  or_5   g18409(.A(new_n20757), .B(new_n20754), .Y(new_n20758));
  nand_5 g18410(.A(new_n20757), .B(new_n20754), .Y(new_n20759));
  not_8  g18411(.A(new_n3272), .Y(new_n20760));
  nor_5  g18412(.A(new_n3310), .B(new_n20760), .Y(new_n20761_1));
  nor_5  g18413(.A(new_n20761_1), .B(new_n3309), .Y(new_n20762));
  not_8  g18414(.A(new_n20762), .Y(new_n20763));
  nand_5 g18415(.A(new_n20763), .B(new_n20759), .Y(new_n20764));
  nand_5 g18416(.A(new_n20764), .B(new_n20758), .Y(new_n20765));
  nand_5 g18417(.A(new_n20765), .B(new_n20752), .Y(new_n20766));
  nand_5 g18418(.A(new_n20766), .B(new_n20751), .Y(new_n20767));
  nand_5 g18419(.A(new_n20742), .B(new_n20731), .Y(new_n20768));
  nand_5 g18420(.A(new_n20768), .B(new_n20732), .Y(new_n20769));
  nand_5 g18421(.A(new_n20769), .B(new_n20749), .Y(new_n20770));
  nand_5 g18422(.A(new_n20770), .B(new_n20767), .Y(new_n20771));
  not_8  g18423(.A(new_n20769), .Y(new_n20772));
  nand_5 g18424(.A(new_n20772), .B(new_n20750), .Y(new_n20773));
  nand_5 g18425(.A(new_n20773), .B(new_n20766), .Y(new_n20774_1));
  and_5  g18426(.A(new_n20774_1), .B(new_n20771), .Y(n5020));
  nand_5 g18427(.A(new_n2378), .B(new_n2383), .Y(new_n20776));
  or_5   g18428(.A(new_n20776), .B(n16722), .Y(new_n20777));
  nand_5 g18429(.A(new_n20776), .B(n16722), .Y(new_n20778));
  and_5  g18430(.A(new_n20778), .B(new_n20777), .Y(new_n20779));
  or_5   g18431(.A(new_n20779), .B(new_n3148), .Y(new_n20780));
  nand_5 g18432(.A(new_n20779), .B(new_n3148), .Y(new_n20781));
  nand_5 g18433(.A(n13781), .B(n11486), .Y(new_n20782));
  and_5  g18434(.A(new_n20782), .B(new_n20776), .Y(new_n20783));
  or_5   g18435(.A(new_n20783), .B(new_n3156), .Y(new_n20784));
  nand_5 g18436(.A(new_n20783), .B(new_n3156), .Y(new_n20785));
  nand_5 g18437(.A(new_n3166), .B(new_n2378), .Y(new_n20786));
  not_8  g18438(.A(new_n20786), .Y(new_n20787));
  nand_5 g18439(.A(new_n20787), .B(new_n20785), .Y(new_n20788_1));
  nand_5 g18440(.A(new_n20788_1), .B(new_n20784), .Y(new_n20789));
  nand_5 g18441(.A(new_n20789), .B(new_n20781), .Y(new_n20790));
  nand_5 g18442(.A(new_n20790), .B(new_n20780), .Y(new_n20791));
  nor_5  g18443(.A(new_n20777), .B(n3480), .Y(new_n20792));
  not_8  g18444(.A(new_n20792), .Y(new_n20793));
  nand_5 g18445(.A(new_n20777), .B(n3480), .Y(new_n20794_1));
  and_5  g18446(.A(new_n20794_1), .B(new_n20793), .Y(new_n20795_1));
  or_5   g18447(.A(new_n20795_1), .B(new_n3138), .Y(new_n20796));
  nand_5 g18448(.A(new_n20795_1), .B(new_n3138), .Y(new_n20797));
  nand_5 g18449(.A(new_n20797), .B(new_n20796), .Y(new_n20798));
  xor_4  g18450(.A(new_n20798), .B(new_n20791), .Y(new_n20799));
  nand_5 g18451(.A(new_n20799), .B(new_n7916), .Y(new_n20800));
  or_5   g18452(.A(new_n20799), .B(new_n7916), .Y(new_n20801));
  nand_5 g18453(.A(new_n20781), .B(new_n20780), .Y(new_n20802));
  xor_4  g18454(.A(new_n20802), .B(new_n20789), .Y(new_n20803_1));
  nand_5 g18455(.A(new_n20803_1), .B(new_n7922), .Y(new_n20804));
  or_5   g18456(.A(new_n20803_1), .B(new_n7922), .Y(new_n20805));
  nand_5 g18457(.A(new_n20785), .B(new_n20784), .Y(new_n20806));
  xor_4  g18458(.A(new_n20806), .B(new_n20787), .Y(new_n20807));
  or_5   g18459(.A(new_n20807), .B(new_n7928), .Y(new_n20808));
  nand_5 g18460(.A(new_n20807), .B(new_n7928), .Y(new_n20809));
  nor_5  g18461(.A(new_n3166), .B(new_n2378), .Y(new_n20810));
  nor_5  g18462(.A(new_n20810), .B(new_n20787), .Y(new_n20811));
  nor_5  g18463(.A(new_n20811), .B(new_n13537), .Y(new_n20812));
  not_8  g18464(.A(new_n20812), .Y(new_n20813));
  nand_5 g18465(.A(new_n20813), .B(new_n20809), .Y(new_n20814));
  nand_5 g18466(.A(new_n20814), .B(new_n20808), .Y(new_n20815));
  not_8  g18467(.A(new_n20815), .Y(new_n20816));
  nand_5 g18468(.A(new_n20816), .B(new_n20805), .Y(new_n20817));
  nand_5 g18469(.A(new_n20817), .B(new_n20804), .Y(new_n20818));
  nand_5 g18470(.A(new_n20818), .B(new_n20801), .Y(new_n20819));
  nand_5 g18471(.A(new_n20819), .B(new_n20800), .Y(new_n20820));
  nand_5 g18472(.A(new_n20797), .B(new_n20791), .Y(new_n20821));
  nand_5 g18473(.A(new_n20821), .B(new_n20796), .Y(new_n20822));
  nand_5 g18474(.A(new_n20792), .B(new_n2412), .Y(new_n20823));
  nand_5 g18475(.A(new_n20793), .B(n3018), .Y(new_n20824));
  and_5  g18476(.A(new_n20824), .B(new_n20823), .Y(new_n20825));
  or_5   g18477(.A(new_n20825), .B(new_n3129), .Y(new_n20826_1));
  nand_5 g18478(.A(new_n20825), .B(new_n3129), .Y(new_n20827));
  nand_5 g18479(.A(new_n20827), .B(new_n20826_1), .Y(new_n20828));
  xor_4  g18480(.A(new_n20828), .B(new_n20822), .Y(new_n20829));
  nand_5 g18481(.A(new_n20829), .B(new_n7909), .Y(new_n20830));
  not_8  g18482(.A(new_n20830), .Y(new_n20831));
  nor_5  g18483(.A(new_n20829), .B(new_n7909), .Y(new_n20832));
  nor_5  g18484(.A(new_n20832), .B(new_n20831), .Y(new_n20833));
  xor_4  g18485(.A(new_n20833), .B(new_n20820), .Y(n5024));
  nand_5 g18486(.A(new_n4013), .B(new_n4012), .Y(new_n20835));
  xnor_4 g18487(.A(new_n20835), .B(new_n4054), .Y(n5046));
  xor_4  g18488(.A(new_n6626), .B(new_n6625), .Y(n5062));
  nand_5 g18489(.A(new_n14339), .B(new_n14338), .Y(new_n20838));
  xor_4  g18490(.A(new_n20838), .B(new_n14364_1), .Y(n5064));
  nand_5 g18491(.A(n12495), .B(n11479), .Y(new_n20840));
  nand_5 g18492(.A(new_n5669), .B(new_n8170), .Y(new_n20841));
  and_5  g18493(.A(new_n20841), .B(new_n20840), .Y(new_n20842));
  or_5   g18494(.A(new_n20842), .B(new_n2380), .Y(new_n20843));
  not_8  g18495(.A(new_n2387_1), .Y(new_n20844));
  nand_5 g18496(.A(new_n9765), .B(new_n8168), .Y(new_n20845));
  nand_5 g18497(.A(n20235), .B(n8259), .Y(new_n20846));
  nand_5 g18498(.A(new_n20846), .B(new_n20845), .Y(new_n20847));
  xnor_4 g18499(.A(new_n20847), .B(new_n20840), .Y(new_n20848));
  or_5   g18500(.A(new_n20848), .B(new_n20844), .Y(new_n20849));
  nand_5 g18501(.A(new_n20848), .B(new_n20844), .Y(new_n20850));
  nand_5 g18502(.A(new_n20850), .B(new_n20849), .Y(new_n20851));
  xor_4  g18503(.A(new_n20851), .B(new_n20843), .Y(new_n20852));
  nand_5 g18504(.A(new_n20842), .B(new_n2380), .Y(new_n20853));
  nand_5 g18505(.A(new_n20853), .B(new_n20843), .Y(new_n20854));
  nand_5 g18506(.A(n9251), .B(new_n11256), .Y(new_n20855));
  nand_5 g18507(.A(new_n3850_1), .B(n7428), .Y(new_n20856));
  nand_5 g18508(.A(new_n20856), .B(new_n20855), .Y(new_n20857));
  nand_5 g18509(.A(new_n20857), .B(new_n20854), .Y(new_n20858));
  not_8  g18510(.A(new_n20858), .Y(new_n20859));
  nand_5 g18511(.A(new_n2502), .B(n10372), .Y(new_n20860));
  nand_5 g18512(.A(n20138), .B(new_n8038), .Y(new_n20861));
  nand_5 g18513(.A(new_n20861), .B(new_n20860), .Y(new_n20862));
  xnor_4 g18514(.A(new_n20862), .B(new_n20855), .Y(new_n20863));
  nand_5 g18515(.A(new_n20863), .B(new_n20859), .Y(new_n20864));
  or_5   g18516(.A(new_n20863), .B(new_n20859), .Y(new_n20865));
  nand_5 g18517(.A(new_n20865), .B(new_n20864), .Y(new_n20866));
  xor_4  g18518(.A(new_n20866), .B(new_n20852), .Y(n5082));
  xor_4  g18519(.A(new_n15655), .B(new_n15653), .Y(n5120));
  nand_5 g18520(.A(new_n16980), .B(new_n16981), .Y(new_n20869_1));
  xor_4  g18521(.A(new_n20869_1), .B(new_n16989_1), .Y(n5158));
  nand_5 g18522(.A(new_n18523), .B(new_n18522), .Y(new_n20871));
  xnor_4 g18523(.A(new_n20871), .B(new_n18541), .Y(n5168));
  nand_5 g18524(.A(new_n19787), .B(n6659), .Y(new_n20873));
  nand_5 g18525(.A(new_n19786), .B(new_n18162), .Y(new_n20874));
  nand_5 g18526(.A(new_n20874), .B(new_n20873), .Y(new_n20875));
  nand_5 g18527(.A(new_n16450), .B(new_n18166), .Y(new_n20876));
  nand_5 g18528(.A(new_n16448), .B(n23250), .Y(new_n20877));
  nand_5 g18529(.A(new_n16362), .B(new_n18169), .Y(new_n20878));
  nand_5 g18530(.A(new_n16360), .B(n11455), .Y(new_n20879_1));
  nand_5 g18531(.A(new_n16319), .B(new_n18172), .Y(new_n20880));
  nand_5 g18532(.A(new_n16317), .B(n3945), .Y(new_n20881));
  nand_5 g18533(.A(new_n16324), .B(new_n5879), .Y(new_n20882));
  nand_5 g18534(.A(new_n16322_1), .B(n5255), .Y(new_n20883));
  nand_5 g18535(.A(new_n17506), .B(new_n17504), .Y(new_n20884));
  nand_5 g18536(.A(new_n20884), .B(new_n17505), .Y(new_n20885));
  nand_5 g18537(.A(new_n20885), .B(new_n20883), .Y(new_n20886));
  nand_5 g18538(.A(new_n20886), .B(new_n20882), .Y(new_n20887));
  nand_5 g18539(.A(new_n20887), .B(new_n20881), .Y(new_n20888));
  nand_5 g18540(.A(new_n20888), .B(new_n20880), .Y(new_n20889));
  nand_5 g18541(.A(new_n20889), .B(new_n20879_1), .Y(new_n20890));
  nand_5 g18542(.A(new_n20890), .B(new_n20878), .Y(new_n20891));
  nand_5 g18543(.A(new_n20891), .B(new_n20877), .Y(new_n20892));
  nand_5 g18544(.A(new_n20892), .B(new_n20876), .Y(new_n20893));
  xor_4  g18545(.A(new_n20893), .B(new_n20875), .Y(new_n20894));
  nand_5 g18546(.A(new_n20894), .B(new_n18159), .Y(new_n20895));
  or_5   g18547(.A(new_n20894), .B(new_n18159), .Y(new_n20896));
  nand_5 g18548(.A(new_n20896), .B(new_n20895), .Y(new_n20897));
  nand_5 g18549(.A(new_n20876), .B(new_n20877), .Y(new_n20898));
  xor_4  g18550(.A(new_n20898), .B(new_n20891), .Y(new_n20899));
  or_5   g18551(.A(new_n20899), .B(new_n18256), .Y(new_n20900));
  nand_5 g18552(.A(new_n20899), .B(new_n18256), .Y(new_n20901));
  nand_5 g18553(.A(new_n20878), .B(new_n20879_1), .Y(new_n20902));
  xor_4  g18554(.A(new_n20902), .B(new_n20889), .Y(new_n20903));
  or_5   g18555(.A(new_n20903), .B(new_n18263), .Y(new_n20904));
  nand_5 g18556(.A(new_n20903), .B(new_n18263), .Y(new_n20905));
  nand_5 g18557(.A(new_n20880), .B(new_n20881), .Y(new_n20906));
  xor_4  g18558(.A(new_n20906), .B(new_n20887), .Y(new_n20907));
  or_5   g18559(.A(new_n20907), .B(new_n18270), .Y(new_n20908));
  nand_5 g18560(.A(new_n20907), .B(new_n18270), .Y(new_n20909));
  nand_5 g18561(.A(new_n20882), .B(new_n20883), .Y(new_n20910));
  xor_4  g18562(.A(new_n20910), .B(new_n20885), .Y(new_n20911));
  or_5   g18563(.A(new_n20911), .B(new_n18279), .Y(new_n20912));
  nand_5 g18564(.A(new_n20911), .B(new_n18279), .Y(new_n20913));
  nand_5 g18565(.A(new_n17510), .B(new_n17489), .Y(new_n20914));
  nand_5 g18566(.A(new_n20914), .B(new_n17509), .Y(new_n20915_1));
  nand_5 g18567(.A(new_n20915_1), .B(new_n20913), .Y(new_n20916));
  nand_5 g18568(.A(new_n20916), .B(new_n20912), .Y(new_n20917));
  nand_5 g18569(.A(new_n20917), .B(new_n20909), .Y(new_n20918));
  nand_5 g18570(.A(new_n20918), .B(new_n20908), .Y(new_n20919));
  nand_5 g18571(.A(new_n20919), .B(new_n20905), .Y(new_n20920));
  nand_5 g18572(.A(new_n20920), .B(new_n20904), .Y(new_n20921));
  nand_5 g18573(.A(new_n20921), .B(new_n20901), .Y(new_n20922));
  nand_5 g18574(.A(new_n20922), .B(new_n20900), .Y(new_n20923_1));
  xor_4  g18575(.A(new_n20923_1), .B(new_n20897), .Y(n5184));
  nor_5  g18576(.A(new_n5133), .B(new_n5041), .Y(new_n20925));
  nor_5  g18577(.A(new_n5134), .B(new_n5040), .Y(new_n20926));
  nor_5  g18578(.A(new_n20926), .B(new_n20925), .Y(n5228));
  nand_5 g18579(.A(new_n12995), .B(new_n12991), .Y(new_n20928));
  nand_5 g18580(.A(new_n20928), .B(new_n12994), .Y(new_n20929_1));
  not_8  g18581(.A(new_n20929_1), .Y(new_n20930));
  nand_5 g18582(.A(new_n20930), .B(new_n8139_1), .Y(new_n20931));
  nand_5 g18583(.A(new_n20929_1), .B(new_n8138), .Y(new_n20932));
  nand_5 g18584(.A(new_n20932), .B(new_n20931), .Y(new_n20933));
  nand_5 g18585(.A(new_n13018), .B(new_n8197), .Y(new_n20934));
  or_5   g18586(.A(new_n13018), .B(new_n8197), .Y(new_n20935_1));
  nand_5 g18587(.A(new_n14367), .B(new_n14366), .Y(new_n20936_1));
  nand_5 g18588(.A(new_n20936_1), .B(new_n14368), .Y(new_n20937));
  nand_5 g18589(.A(new_n20937), .B(new_n20935_1), .Y(new_n20938));
  nand_5 g18590(.A(new_n20938), .B(new_n20934), .Y(new_n20939));
  xor_4  g18591(.A(new_n20939), .B(new_n20933), .Y(n5256));
  nand_5 g18592(.A(new_n7580), .B(new_n7579), .Y(new_n20941));
  xor_4  g18593(.A(new_n20941), .B(new_n7596), .Y(n5265));
  nand_5 g18594(.A(new_n19437), .B(new_n19435), .Y(new_n20943));
  xnor_4 g18595(.A(new_n20943), .B(new_n19498), .Y(n5273));
  nand_5 g18596(.A(new_n19141_1), .B(new_n19139), .Y(new_n20945));
  nand_5 g18597(.A(new_n20945), .B(new_n19140), .Y(new_n20946_1));
  not_8  g18598(.A(new_n20946_1), .Y(new_n20947));
  nand_5 g18599(.A(n7751), .B(new_n7757), .Y(new_n20948));
  nand_5 g18600(.A(new_n2584), .B(n1112), .Y(new_n20949));
  nand_5 g18601(.A(new_n20949), .B(new_n20948), .Y(new_n20950));
  xor_4  g18602(.A(new_n20950), .B(new_n20947), .Y(new_n20951));
  nand_5 g18603(.A(new_n20951), .B(new_n8499), .Y(new_n20952));
  or_5   g18604(.A(new_n20951), .B(new_n8499), .Y(new_n20953));
  not_8  g18605(.A(new_n19137), .Y(new_n20954));
  nor_5  g18606(.A(new_n19146), .B(new_n20954), .Y(new_n20955));
  nor_5  g18607(.A(new_n20955), .B(new_n19145), .Y(new_n20956));
  not_8  g18608(.A(new_n20956), .Y(new_n20957));
  nand_5 g18609(.A(new_n20957), .B(new_n20953), .Y(new_n20958));
  nand_5 g18610(.A(new_n20958), .B(new_n20952), .Y(new_n20959));
  nand_5 g18611(.A(new_n20949), .B(new_n20946_1), .Y(new_n20960));
  nand_5 g18612(.A(new_n20960), .B(new_n20948), .Y(new_n20961));
  nand_5 g18613(.A(n20946), .B(new_n7810), .Y(new_n20962));
  nand_5 g18614(.A(new_n6062), .B(n2289), .Y(new_n20963));
  nand_5 g18615(.A(new_n20963), .B(new_n20962), .Y(new_n20964));
  xnor_4 g18616(.A(new_n20964), .B(new_n20961), .Y(new_n20965));
  nand_5 g18617(.A(new_n20965), .B(new_n8492), .Y(new_n20966));
  not_8  g18618(.A(new_n20966), .Y(new_n20967));
  nor_5  g18619(.A(new_n20965), .B(new_n8492), .Y(new_n20968));
  nor_5  g18620(.A(new_n20968), .B(new_n20967), .Y(new_n20969));
  xor_4  g18621(.A(new_n20969), .B(new_n20959), .Y(n5274));
  nand_5 g18622(.A(new_n4535), .B(new_n4573), .Y(new_n20971));
  not_8  g18623(.A(new_n20971), .Y(new_n20972));
  nand_5 g18624(.A(new_n20972), .B(new_n4586), .Y(new_n20973));
  nand_5 g18625(.A(new_n20971), .B(n919), .Y(new_n20974));
  and_5  g18626(.A(new_n20974), .B(new_n20973), .Y(new_n20975));
  or_5   g18627(.A(new_n20975), .B(new_n10130), .Y(new_n20976));
  nand_5 g18628(.A(new_n20975), .B(new_n10130), .Y(new_n20977));
  nand_5 g18629(.A(n25316), .B(n20385), .Y(new_n20978));
  nand_5 g18630(.A(new_n20978), .B(new_n20971), .Y(new_n20979));
  nand_5 g18631(.A(new_n20979), .B(new_n10144), .Y(new_n20980));
  nor_5  g18632(.A(new_n20979), .B(new_n10144), .Y(new_n20981));
  not_8  g18633(.A(new_n20981), .Y(new_n20982));
  nand_5 g18634(.A(new_n20982), .B(new_n10253), .Y(new_n20983));
  nand_5 g18635(.A(new_n20983), .B(new_n20980), .Y(new_n20984));
  nand_5 g18636(.A(new_n20984), .B(new_n20977), .Y(new_n20985));
  nand_5 g18637(.A(new_n20985), .B(new_n20976), .Y(new_n20986_1));
  xor_4  g18638(.A(new_n20973), .B(n3918), .Y(new_n20987));
  or_5   g18639(.A(new_n20987), .B(new_n10123), .Y(new_n20988));
  nand_5 g18640(.A(new_n20987), .B(new_n10123), .Y(new_n20989));
  nand_5 g18641(.A(new_n20989), .B(new_n20988), .Y(new_n20990));
  xor_4  g18642(.A(new_n20990), .B(new_n20986_1), .Y(new_n20991));
  not_8  g18643(.A(new_n20991), .Y(new_n20992));
  nand_5 g18644(.A(new_n4610), .B(n24786), .Y(new_n20993));
  nand_5 g18645(.A(new_n4609), .B(new_n4596), .Y(new_n20994));
  nand_5 g18646(.A(new_n4564), .B(n27120), .Y(new_n20995));
  nand_5 g18647(.A(new_n4567), .B(new_n4553), .Y(new_n20996));
  nand_5 g18648(.A(new_n4550), .B(new_n4542), .Y(new_n20997));
  nand_5 g18649(.A(new_n20997), .B(new_n20996), .Y(new_n20998));
  nand_5 g18650(.A(new_n20998), .B(new_n20995), .Y(new_n20999));
  nand_5 g18651(.A(new_n20999), .B(new_n20994), .Y(new_n21000));
  nand_5 g18652(.A(new_n21000), .B(new_n20993), .Y(new_n21001));
  nand_5 g18653(.A(new_n18860), .B(n25370), .Y(new_n21002));
  nand_5 g18654(.A(new_n18862), .B(new_n7825), .Y(new_n21003));
  nand_5 g18655(.A(new_n21003), .B(new_n21002), .Y(new_n21004));
  xor_4  g18656(.A(new_n21004), .B(new_n21001), .Y(new_n21005));
  or_5   g18657(.A(new_n21005), .B(new_n20992), .Y(new_n21006));
  nand_5 g18658(.A(new_n21005), .B(new_n20992), .Y(new_n21007));
  nand_5 g18659(.A(new_n20977), .B(new_n20976), .Y(new_n21008_1));
  xor_4  g18660(.A(new_n21008_1), .B(new_n20984), .Y(new_n21009));
  not_8  g18661(.A(new_n21009), .Y(new_n21010));
  nand_5 g18662(.A(new_n20994), .B(new_n20993), .Y(new_n21011));
  xor_4  g18663(.A(new_n21011), .B(new_n20999), .Y(new_n21012));
  or_5   g18664(.A(new_n21012), .B(new_n21010), .Y(new_n21013));
  nand_5 g18665(.A(new_n21012), .B(new_n21010), .Y(new_n21014));
  nand_5 g18666(.A(new_n20982), .B(new_n20980), .Y(new_n21015));
  xor_4  g18667(.A(new_n21015), .B(new_n10254), .Y(new_n21016));
  nand_5 g18668(.A(new_n20996), .B(new_n20995), .Y(new_n21017_1));
  xor_4  g18669(.A(new_n21017_1), .B(new_n20997), .Y(new_n21018));
  nand_5 g18670(.A(new_n21018), .B(new_n21016), .Y(new_n21019));
  nor_5  g18671(.A(new_n21018), .B(new_n21016), .Y(new_n21020));
  not_8  g18672(.A(new_n21020), .Y(new_n21021));
  xor_4  g18673(.A(new_n4549), .B(n23065), .Y(new_n21022));
  nor_5  g18674(.A(new_n21022), .B(new_n10256), .Y(new_n21023));
  not_8  g18675(.A(new_n21023), .Y(new_n21024));
  nand_5 g18676(.A(new_n21024), .B(new_n21021), .Y(new_n21025));
  and_5  g18677(.A(new_n21025), .B(new_n21019), .Y(new_n21026));
  nand_5 g18678(.A(new_n21026), .B(new_n21014), .Y(new_n21027));
  nand_5 g18679(.A(new_n21027), .B(new_n21013), .Y(new_n21028));
  nand_5 g18680(.A(new_n21028), .B(new_n21007), .Y(new_n21029));
  nand_5 g18681(.A(new_n21029), .B(new_n21006), .Y(new_n21030));
  nand_5 g18682(.A(new_n20989), .B(new_n20986_1), .Y(new_n21031));
  nand_5 g18683(.A(new_n21031), .B(new_n20988), .Y(new_n21032));
  nor_5  g18684(.A(new_n20973), .B(n3918), .Y(new_n21033));
  nand_5 g18685(.A(new_n21033), .B(new_n7185), .Y(new_n21034_1));
  or_5   g18686(.A(new_n21033), .B(new_n7185), .Y(new_n21035));
  and_5  g18687(.A(new_n21035), .B(new_n21034_1), .Y(new_n21036));
  or_5   g18688(.A(new_n21036), .B(new_n10116), .Y(new_n21037));
  nand_5 g18689(.A(new_n21036), .B(new_n10116), .Y(new_n21038));
  nand_5 g18690(.A(new_n21038), .B(new_n21037), .Y(new_n21039));
  xor_4  g18691(.A(new_n21039), .B(new_n21032), .Y(new_n21040));
  not_8  g18692(.A(new_n21040), .Y(new_n21041));
  nand_5 g18693(.A(new_n21003), .B(new_n21001), .Y(new_n21042));
  nand_5 g18694(.A(new_n21042), .B(new_n21002), .Y(new_n21043));
  nand_5 g18695(.A(new_n18855), .B(n19472), .Y(new_n21044));
  nand_5 g18696(.A(new_n18857), .B(new_n7822), .Y(new_n21045));
  nand_5 g18697(.A(new_n21045), .B(new_n21044), .Y(new_n21046_1));
  xor_4  g18698(.A(new_n21046_1), .B(new_n21043), .Y(new_n21047));
  or_5   g18699(.A(new_n21047), .B(new_n21041), .Y(new_n21048));
  nand_5 g18700(.A(new_n21047), .B(new_n21041), .Y(new_n21049));
  nand_5 g18701(.A(new_n21049), .B(new_n21048), .Y(new_n21050));
  xnor_4 g18702(.A(new_n21050), .B(new_n21030), .Y(n5300));
  nand_5 g18703(.A(new_n8137), .B(new_n8066), .Y(new_n21052));
  nand_5 g18704(.A(new_n21052), .B(new_n8068), .Y(new_n21053));
  and_5  g18705(.A(new_n21053), .B(new_n20929_1), .Y(new_n21054));
  xor_4  g18706(.A(new_n21053), .B(new_n20930), .Y(new_n21055));
  nand_5 g18707(.A(new_n20939), .B(new_n20931), .Y(new_n21056));
  nand_5 g18708(.A(new_n21056), .B(new_n20932), .Y(new_n21057));
  nor_5  g18709(.A(new_n21057), .B(new_n21055), .Y(new_n21058));
  nor_5  g18710(.A(new_n21058), .B(new_n21054), .Y(n5325));
  nand_5 g18711(.A(new_n8798), .B(new_n8291), .Y(new_n21060));
  nand_5 g18712(.A(n25120), .B(n17458), .Y(new_n21061));
  nand_5 g18713(.A(new_n21061), .B(new_n21060), .Y(new_n21062_1));
  nand_5 g18714(.A(new_n8801), .B(new_n8294), .Y(new_n21063));
  nand_5 g18715(.A(n8363), .B(n1222), .Y(new_n21064));
  nand_5 g18716(.A(new_n8297), .B(new_n8804), .Y(new_n21065));
  nand_5 g18717(.A(n25240), .B(n14680), .Y(new_n21066));
  nand_5 g18718(.A(new_n8807), .B(new_n8300), .Y(new_n21067));
  nand_5 g18719(.A(n17250), .B(n10125), .Y(new_n21068));
  nand_5 g18720(.A(new_n8810), .B(new_n8303), .Y(new_n21069));
  nand_5 g18721(.A(n23160), .B(n8067), .Y(new_n21070));
  nand_5 g18722(.A(new_n14834), .B(new_n14831), .Y(new_n21071));
  nand_5 g18723(.A(new_n21071), .B(new_n14833), .Y(new_n21072));
  nand_5 g18724(.A(new_n21072), .B(new_n21070), .Y(new_n21073));
  nand_5 g18725(.A(new_n21073), .B(new_n21069), .Y(new_n21074));
  nand_5 g18726(.A(new_n21074), .B(new_n21068), .Y(new_n21075));
  nand_5 g18727(.A(new_n21075), .B(new_n21067), .Y(new_n21076));
  nand_5 g18728(.A(new_n21076), .B(new_n21066), .Y(new_n21077));
  nand_5 g18729(.A(new_n21077), .B(new_n21065), .Y(new_n21078_1));
  nand_5 g18730(.A(new_n21078_1), .B(new_n21064), .Y(new_n21079));
  nand_5 g18731(.A(new_n21079), .B(new_n21063), .Y(new_n21080));
  xor_4  g18732(.A(new_n21080), .B(new_n21062_1), .Y(new_n21081));
  nand_5 g18733(.A(new_n21081), .B(n23272), .Y(new_n21082));
  or_5   g18734(.A(new_n21081), .B(n23272), .Y(new_n21083));
  nand_5 g18735(.A(new_n21064), .B(new_n21063), .Y(new_n21084));
  xor_4  g18736(.A(new_n21084), .B(new_n21078_1), .Y(new_n21085));
  nand_5 g18737(.A(new_n21085), .B(n11481), .Y(new_n21086));
  or_5   g18738(.A(new_n21085), .B(n11481), .Y(new_n21087));
  nand_5 g18739(.A(new_n21066), .B(new_n21065), .Y(new_n21088));
  xor_4  g18740(.A(new_n21088), .B(new_n21076), .Y(new_n21089));
  nand_5 g18741(.A(new_n21089), .B(n16439), .Y(new_n21090));
  or_5   g18742(.A(new_n21089), .B(n16439), .Y(new_n21091));
  nand_5 g18743(.A(new_n21068), .B(new_n21067), .Y(new_n21092));
  xor_4  g18744(.A(new_n21092), .B(new_n21074), .Y(new_n21093_1));
  nand_5 g18745(.A(new_n21093_1), .B(n15241), .Y(new_n21094_1));
  or_5   g18746(.A(new_n21093_1), .B(n15241), .Y(new_n21095_1));
  nand_5 g18747(.A(new_n21070), .B(new_n21069), .Y(new_n21096));
  xor_4  g18748(.A(new_n21096), .B(new_n21072), .Y(new_n21097));
  nand_5 g18749(.A(new_n21097), .B(n7678), .Y(new_n21098));
  or_5   g18750(.A(new_n21097), .B(n7678), .Y(new_n21099));
  nand_5 g18751(.A(new_n14838), .B(new_n14828), .Y(new_n21100));
  nand_5 g18752(.A(new_n21100), .B(new_n14837), .Y(new_n21101));
  nand_5 g18753(.A(new_n21101), .B(new_n21099), .Y(new_n21102));
  nand_5 g18754(.A(new_n21102), .B(new_n21098), .Y(new_n21103));
  nand_5 g18755(.A(new_n21103), .B(new_n21095_1), .Y(new_n21104));
  nand_5 g18756(.A(new_n21104), .B(new_n21094_1), .Y(new_n21105));
  nand_5 g18757(.A(new_n21105), .B(new_n21091), .Y(new_n21106));
  nand_5 g18758(.A(new_n21106), .B(new_n21090), .Y(new_n21107));
  nand_5 g18759(.A(new_n21107), .B(new_n21087), .Y(new_n21108));
  nand_5 g18760(.A(new_n21108), .B(new_n21086), .Y(new_n21109));
  nand_5 g18761(.A(new_n21109), .B(new_n21083), .Y(new_n21110));
  nand_5 g18762(.A(new_n21110), .B(new_n21082), .Y(new_n21111));
  nand_5 g18763(.A(new_n21080), .B(new_n21061), .Y(new_n21112));
  nand_5 g18764(.A(new_n21112), .B(new_n21060), .Y(new_n21113));
  not_8  g18765(.A(new_n21113), .Y(new_n21114));
  nand_5 g18766(.A(new_n21114), .B(new_n21111), .Y(new_n21115));
  not_8  g18767(.A(new_n21115), .Y(new_n21116));
  nand_5 g18768(.A(new_n9271), .B(new_n11696), .Y(new_n21117));
  nand_5 g18769(.A(n12702), .B(n12507), .Y(new_n21118));
  nand_5 g18770(.A(new_n21118), .B(new_n21117), .Y(new_n21119));
  nand_5 g18771(.A(new_n6168), .B(new_n11699), .Y(new_n21120));
  nand_5 g18772(.A(n26797), .B(n15077), .Y(new_n21121));
  nand_5 g18773(.A(new_n9235), .B(new_n11703), .Y(new_n21122));
  nand_5 g18774(.A(n23913), .B(n3710), .Y(new_n21123_1));
  nand_5 g18775(.A(new_n11706), .B(new_n6169), .Y(new_n21124));
  nand_5 g18776(.A(n26318), .B(n22554), .Y(new_n21125));
  nand_5 g18777(.A(new_n11710_1), .B(new_n9241), .Y(new_n21126));
  nand_5 g18778(.A(n26054), .B(n20429), .Y(new_n21127));
  nand_5 g18779(.A(new_n11713), .B(new_n6170), .Y(new_n21128));
  nand_5 g18780(.A(n19081), .B(n3909), .Y(new_n21129));
  nand_5 g18781(.A(new_n9247), .B(new_n11716), .Y(new_n21130));
  nand_5 g18782(.A(n23974), .B(n8309), .Y(new_n21131));
  nand_5 g18783(.A(new_n11720), .B(new_n9251_1), .Y(new_n21132));
  nand_5 g18784(.A(n19144), .B(n2146), .Y(new_n21133));
  nand_5 g18785(.A(new_n19093), .B(new_n19084), .Y(new_n21134_1));
  nand_5 g18786(.A(new_n21134_1), .B(new_n19092), .Y(new_n21135));
  nand_5 g18787(.A(new_n21135), .B(new_n21133), .Y(new_n21136));
  nand_5 g18788(.A(new_n21136), .B(new_n21132), .Y(new_n21137));
  nand_5 g18789(.A(new_n21137), .B(new_n21131), .Y(new_n21138_1));
  nand_5 g18790(.A(new_n21138_1), .B(new_n21130), .Y(new_n21139));
  nand_5 g18791(.A(new_n21139), .B(new_n21129), .Y(new_n21140));
  nand_5 g18792(.A(new_n21140), .B(new_n21128), .Y(new_n21141));
  nand_5 g18793(.A(new_n21141), .B(new_n21127), .Y(new_n21142));
  nand_5 g18794(.A(new_n21142), .B(new_n21126), .Y(new_n21143));
  nand_5 g18795(.A(new_n21143), .B(new_n21125), .Y(new_n21144));
  nand_5 g18796(.A(new_n21144), .B(new_n21124), .Y(new_n21145));
  nand_5 g18797(.A(new_n21145), .B(new_n21123_1), .Y(new_n21146));
  nand_5 g18798(.A(new_n21146), .B(new_n21122), .Y(new_n21147));
  nand_5 g18799(.A(new_n21147), .B(new_n21121), .Y(new_n21148));
  nand_5 g18800(.A(new_n21148), .B(new_n21120), .Y(new_n21149));
  xor_4  g18801(.A(new_n21149), .B(new_n21119), .Y(new_n21150));
  nand_5 g18802(.A(new_n21150), .B(n12650), .Y(new_n21151));
  or_5   g18803(.A(new_n21150), .B(n12650), .Y(new_n21152));
  nand_5 g18804(.A(new_n21121), .B(new_n21120), .Y(new_n21153));
  xor_4  g18805(.A(new_n21153), .B(new_n21147), .Y(new_n21154_1));
  nand_5 g18806(.A(new_n21154_1), .B(n10201), .Y(new_n21155));
  or_5   g18807(.A(new_n21154_1), .B(n10201), .Y(new_n21156));
  nand_5 g18808(.A(new_n21123_1), .B(new_n21122), .Y(new_n21157_1));
  xor_4  g18809(.A(new_n21157_1), .B(new_n21145), .Y(new_n21158));
  nand_5 g18810(.A(new_n21158), .B(n10593), .Y(new_n21159));
  or_5   g18811(.A(new_n21158), .B(n10593), .Y(new_n21160));
  nand_5 g18812(.A(new_n21125), .B(new_n21124), .Y(new_n21161));
  xor_4  g18813(.A(new_n21161), .B(new_n21143), .Y(new_n21162));
  nand_5 g18814(.A(new_n21162), .B(n18290), .Y(new_n21163));
  or_5   g18815(.A(new_n21162), .B(n18290), .Y(new_n21164));
  nand_5 g18816(.A(new_n21127), .B(new_n21126), .Y(new_n21165));
  xor_4  g18817(.A(new_n21165), .B(new_n21141), .Y(new_n21166));
  nand_5 g18818(.A(new_n21166), .B(n11580), .Y(new_n21167));
  or_5   g18819(.A(new_n21166), .B(n11580), .Y(new_n21168_1));
  nand_5 g18820(.A(new_n21129), .B(new_n21128), .Y(new_n21169));
  xor_4  g18821(.A(new_n21169), .B(new_n21139), .Y(new_n21170));
  nand_5 g18822(.A(new_n21170), .B(n15884), .Y(new_n21171));
  or_5   g18823(.A(new_n21170), .B(n15884), .Y(new_n21172));
  nand_5 g18824(.A(new_n21131), .B(new_n21130), .Y(new_n21173_1));
  xor_4  g18825(.A(new_n21173_1), .B(new_n21137), .Y(new_n21174));
  nand_5 g18826(.A(new_n21174), .B(n6356), .Y(new_n21175));
  or_5   g18827(.A(new_n21174), .B(n6356), .Y(new_n21176_1));
  nand_5 g18828(.A(new_n21133), .B(new_n21132), .Y(new_n21177));
  xor_4  g18829(.A(new_n21177), .B(new_n21135), .Y(new_n21178));
  nand_5 g18830(.A(new_n21178), .B(n27104), .Y(new_n21179));
  or_5   g18831(.A(new_n21178), .B(n27104), .Y(new_n21180));
  nand_5 g18832(.A(new_n19097), .B(new_n19090), .Y(new_n21181));
  nand_5 g18833(.A(new_n21181), .B(new_n19096), .Y(new_n21182_1));
  nand_5 g18834(.A(new_n21182_1), .B(new_n21180), .Y(new_n21183));
  nand_5 g18835(.A(new_n21183), .B(new_n21179), .Y(new_n21184));
  nand_5 g18836(.A(new_n21184), .B(new_n21176_1), .Y(new_n21185));
  nand_5 g18837(.A(new_n21185), .B(new_n21175), .Y(new_n21186));
  nand_5 g18838(.A(new_n21186), .B(new_n21172), .Y(new_n21187));
  nand_5 g18839(.A(new_n21187), .B(new_n21171), .Y(new_n21188));
  nand_5 g18840(.A(new_n21188), .B(new_n21168_1), .Y(new_n21189));
  nand_5 g18841(.A(new_n21189), .B(new_n21167), .Y(new_n21190));
  nand_5 g18842(.A(new_n21190), .B(new_n21164), .Y(new_n21191));
  nand_5 g18843(.A(new_n21191), .B(new_n21163), .Y(new_n21192));
  nand_5 g18844(.A(new_n21192), .B(new_n21160), .Y(new_n21193_1));
  nand_5 g18845(.A(new_n21193_1), .B(new_n21159), .Y(new_n21194));
  nand_5 g18846(.A(new_n21194), .B(new_n21156), .Y(new_n21195));
  nand_5 g18847(.A(new_n21195), .B(new_n21155), .Y(new_n21196));
  nand_5 g18848(.A(new_n21196), .B(new_n21152), .Y(new_n21197));
  nand_5 g18849(.A(new_n21197), .B(new_n21151), .Y(new_n21198));
  nand_5 g18850(.A(new_n21149), .B(new_n21118), .Y(new_n21199));
  nand_5 g18851(.A(new_n21199), .B(new_n21117), .Y(new_n21200));
  not_8  g18852(.A(new_n21200), .Y(new_n21201));
  nand_5 g18853(.A(new_n21201), .B(new_n21198), .Y(new_n21202));
  or_5   g18854(.A(new_n21202), .B(new_n21116), .Y(new_n21203_1));
  nand_5 g18855(.A(new_n21202), .B(new_n21116), .Y(new_n21204));
  nand_5 g18856(.A(new_n21204), .B(new_n21203_1), .Y(new_n21205));
  nor_5  g18857(.A(new_n21114), .B(new_n21111), .Y(new_n21206));
  nor_5  g18858(.A(new_n21206), .B(new_n21116), .Y(new_n21207));
  xor_4  g18859(.A(new_n21200), .B(new_n21198), .Y(new_n21208));
  or_5   g18860(.A(new_n21208), .B(new_n21207), .Y(new_n21209));
  nand_5 g18861(.A(new_n21208), .B(new_n21207), .Y(new_n21210));
  nand_5 g18862(.A(new_n21083), .B(new_n21082), .Y(new_n21211));
  xor_4  g18863(.A(new_n21211), .B(new_n21109), .Y(new_n21212));
  not_8  g18864(.A(new_n21212), .Y(new_n21213));
  nand_5 g18865(.A(new_n21152), .B(new_n21151), .Y(new_n21214));
  xor_4  g18866(.A(new_n21214), .B(new_n21196), .Y(new_n21215));
  or_5   g18867(.A(new_n21215), .B(new_n21213), .Y(new_n21216));
  nand_5 g18868(.A(new_n21215), .B(new_n21213), .Y(new_n21217));
  nand_5 g18869(.A(new_n21087), .B(new_n21086), .Y(new_n21218));
  xor_4  g18870(.A(new_n21218), .B(new_n21107), .Y(new_n21219));
  not_8  g18871(.A(new_n21219), .Y(new_n21220));
  nand_5 g18872(.A(new_n21156), .B(new_n21155), .Y(new_n21221));
  xor_4  g18873(.A(new_n21221), .B(new_n21194), .Y(new_n21222_1));
  or_5   g18874(.A(new_n21222_1), .B(new_n21220), .Y(new_n21223));
  nand_5 g18875(.A(new_n21222_1), .B(new_n21220), .Y(new_n21224));
  nand_5 g18876(.A(new_n21091), .B(new_n21090), .Y(new_n21225_1));
  xor_4  g18877(.A(new_n21225_1), .B(new_n21105), .Y(new_n21226_1));
  not_8  g18878(.A(new_n21226_1), .Y(new_n21227));
  nand_5 g18879(.A(new_n21160), .B(new_n21159), .Y(new_n21228));
  xor_4  g18880(.A(new_n21228), .B(new_n21192), .Y(new_n21229));
  or_5   g18881(.A(new_n21229), .B(new_n21227), .Y(new_n21230));
  nand_5 g18882(.A(new_n21229), .B(new_n21227), .Y(new_n21231));
  nand_5 g18883(.A(new_n21095_1), .B(new_n21094_1), .Y(new_n21232));
  xor_4  g18884(.A(new_n21232), .B(new_n21103), .Y(new_n21233));
  not_8  g18885(.A(new_n21233), .Y(new_n21234));
  nand_5 g18886(.A(new_n21164), .B(new_n21163), .Y(new_n21235));
  xor_4  g18887(.A(new_n21235), .B(new_n21190), .Y(new_n21236));
  or_5   g18888(.A(new_n21236), .B(new_n21234), .Y(new_n21237));
  nand_5 g18889(.A(new_n21236), .B(new_n21234), .Y(new_n21238_1));
  nand_5 g18890(.A(new_n21099), .B(new_n21098), .Y(new_n21239));
  xor_4  g18891(.A(new_n21239), .B(new_n21101), .Y(new_n21240));
  not_8  g18892(.A(new_n21240), .Y(new_n21241));
  nand_5 g18893(.A(new_n21168_1), .B(new_n21167), .Y(new_n21242));
  xor_4  g18894(.A(new_n21242), .B(new_n21188), .Y(new_n21243));
  or_5   g18895(.A(new_n21243), .B(new_n21241), .Y(new_n21244));
  nand_5 g18896(.A(new_n21243), .B(new_n21241), .Y(new_n21245));
  nand_5 g18897(.A(new_n21172), .B(new_n21171), .Y(new_n21246));
  xor_4  g18898(.A(new_n21246), .B(new_n21186), .Y(new_n21247));
  or_5   g18899(.A(new_n21247), .B(new_n14840), .Y(new_n21248));
  nand_5 g18900(.A(new_n21247), .B(new_n14840), .Y(new_n21249));
  nand_5 g18901(.A(new_n21176_1), .B(new_n21175), .Y(new_n21250));
  xor_4  g18902(.A(new_n21250), .B(new_n21184), .Y(new_n21251));
  or_5   g18903(.A(new_n21251), .B(new_n7614), .Y(new_n21252));
  nand_5 g18904(.A(new_n21251), .B(new_n7614), .Y(new_n21253));
  nand_5 g18905(.A(new_n21180), .B(new_n21179), .Y(new_n21254_1));
  xor_4  g18906(.A(new_n21254_1), .B(new_n21182_1), .Y(new_n21255));
  or_5   g18907(.A(new_n21255), .B(new_n7546), .Y(new_n21256));
  nand_5 g18908(.A(new_n21255), .B(new_n7546), .Y(new_n21257));
  nand_5 g18909(.A(new_n19102), .B(new_n7583), .Y(new_n21258));
  nand_5 g18910(.A(new_n21258), .B(new_n19100), .Y(new_n21259));
  nand_5 g18911(.A(new_n21259), .B(new_n21257), .Y(new_n21260));
  nand_5 g18912(.A(new_n21260), .B(new_n21256), .Y(new_n21261));
  nand_5 g18913(.A(new_n21261), .B(new_n21253), .Y(new_n21262));
  nand_5 g18914(.A(new_n21262), .B(new_n21252), .Y(new_n21263));
  nand_5 g18915(.A(new_n21263), .B(new_n21249), .Y(new_n21264));
  nand_5 g18916(.A(new_n21264), .B(new_n21248), .Y(new_n21265));
  nand_5 g18917(.A(new_n21265), .B(new_n21245), .Y(new_n21266));
  nand_5 g18918(.A(new_n21266), .B(new_n21244), .Y(new_n21267));
  nand_5 g18919(.A(new_n21267), .B(new_n21238_1), .Y(new_n21268));
  nand_5 g18920(.A(new_n21268), .B(new_n21237), .Y(new_n21269));
  nand_5 g18921(.A(new_n21269), .B(new_n21231), .Y(new_n21270));
  nand_5 g18922(.A(new_n21270), .B(new_n21230), .Y(new_n21271));
  nand_5 g18923(.A(new_n21271), .B(new_n21224), .Y(new_n21272));
  nand_5 g18924(.A(new_n21272), .B(new_n21223), .Y(new_n21273));
  nand_5 g18925(.A(new_n21273), .B(new_n21217), .Y(new_n21274));
  nand_5 g18926(.A(new_n21274), .B(new_n21216), .Y(new_n21275));
  nand_5 g18927(.A(new_n21275), .B(new_n21210), .Y(new_n21276_1));
  nand_5 g18928(.A(new_n21276_1), .B(new_n21209), .Y(new_n21277));
  not_8  g18929(.A(new_n21277), .Y(new_n21278));
  xor_4  g18930(.A(new_n21278), .B(new_n21205), .Y(n5351));
  nor_5  g18931(.A(new_n18733), .B(new_n18706), .Y(n5353));
  not_8  g18932(.A(new_n13605), .Y(new_n21281));
  not_8  g18933(.A(new_n13606), .Y(new_n21282));
  nor_5  g18934(.A(new_n13665), .B(new_n21282), .Y(new_n21283));
  nor_5  g18935(.A(new_n21283), .B(new_n21281), .Y(new_n21284));
  nand_5 g18936(.A(new_n13601), .B(new_n13566), .Y(new_n21285));
  nand_5 g18937(.A(new_n21285), .B(new_n13567), .Y(new_n21286));
  nand_5 g18938(.A(new_n21286), .B(new_n21284), .Y(new_n21287_1));
  nand_5 g18939(.A(new_n13543), .B(new_n8349), .Y(new_n21288));
  nand_5 g18940(.A(new_n13563), .B(new_n13546), .Y(new_n21289));
  nand_5 g18941(.A(new_n21289), .B(new_n13547), .Y(new_n21290));
  not_8  g18942(.A(new_n21290), .Y(new_n21291));
  nor_5  g18943(.A(new_n21291), .B(new_n21288), .Y(new_n21292));
  xor_4  g18944(.A(new_n21292), .B(new_n21287_1), .Y(new_n21293));
  not_8  g18945(.A(new_n21287_1), .Y(new_n21294));
  nor_5  g18946(.A(new_n21286), .B(new_n21284), .Y(new_n21295));
  nor_5  g18947(.A(new_n21295), .B(new_n21294), .Y(new_n21296));
  xor_4  g18948(.A(new_n13543), .B(new_n8349), .Y(new_n21297));
  xor_4  g18949(.A(new_n21297), .B(new_n21291), .Y(new_n21298_1));
  nand_5 g18950(.A(new_n21298_1), .B(new_n21296), .Y(new_n21299));
  or_5   g18951(.A(new_n21298_1), .B(new_n21296), .Y(new_n21300));
  nand_5 g18952(.A(new_n13738), .B(new_n13667), .Y(new_n21301));
  nand_5 g18953(.A(new_n21301), .B(new_n13668_1), .Y(new_n21302_1));
  nand_5 g18954(.A(new_n21302_1), .B(new_n21300), .Y(new_n21303));
  nand_5 g18955(.A(new_n21303), .B(new_n21299), .Y(new_n21304));
  xor_4  g18956(.A(new_n21304), .B(new_n21293), .Y(n5399));
  not_8  g18957(.A(new_n19956), .Y(new_n21306));
  nor_5  g18958(.A(new_n19959), .B(new_n21306), .Y(new_n21307));
  nand_5 g18959(.A(new_n19955), .B(new_n16114), .Y(new_n21308));
  nor_5  g18960(.A(new_n21308), .B(new_n21307), .Y(new_n21309));
  not_8  g18961(.A(new_n21309), .Y(new_n21310));
  nand_5 g18962(.A(new_n19966), .B(new_n19961), .Y(new_n21311));
  nand_5 g18963(.A(new_n21311), .B(new_n19963), .Y(new_n21312));
  nor_5  g18964(.A(new_n21312), .B(new_n21310), .Y(new_n21313));
  or_5   g18965(.A(new_n21313), .B(new_n21292), .Y(new_n21314));
  nand_5 g18966(.A(new_n21313), .B(new_n21292), .Y(new_n21315));
  nand_5 g18967(.A(new_n21315), .B(new_n21314), .Y(new_n21316));
  xor_4  g18968(.A(new_n21312), .B(new_n21310), .Y(new_n21317_1));
  not_8  g18969(.A(new_n21317_1), .Y(new_n21318));
  or_5   g18970(.A(new_n21318), .B(new_n21298_1), .Y(new_n21319));
  nand_5 g18971(.A(new_n21318), .B(new_n21298_1), .Y(new_n21320));
  nand_5 g18972(.A(new_n19972), .B(new_n19969), .Y(new_n21321));
  nand_5 g18973(.A(new_n21321), .B(new_n19968_1), .Y(new_n21322));
  nand_5 g18974(.A(new_n21322), .B(new_n21320), .Y(new_n21323));
  nand_5 g18975(.A(new_n21323), .B(new_n21319), .Y(new_n21324));
  xnor_4 g18976(.A(new_n21324), .B(new_n21316), .Y(n5403));
  nand_5 g18977(.A(new_n17786), .B(new_n17785), .Y(new_n21326));
  xor_4  g18978(.A(new_n21326), .B(new_n17830), .Y(n5430));
  not_8  g18979(.A(new_n16631), .Y(new_n21328));
  nand_5 g18980(.A(new_n16633), .B(new_n21328), .Y(new_n21329));
  not_8  g18981(.A(new_n21329), .Y(new_n21330));
  nand_5 g18982(.A(new_n16635), .B(new_n16624), .Y(new_n21331));
  nor_5  g18983(.A(new_n16626), .B(new_n12022), .Y(new_n21332));
  nand_5 g18984(.A(new_n21332), .B(new_n21331), .Y(new_n21333));
  nor_5  g18985(.A(new_n21333), .B(new_n21330), .Y(n5439));
  nand_5 g18986(.A(new_n14061), .B(new_n14062), .Y(new_n21335));
  xnor_4 g18987(.A(new_n21335), .B(new_n14080), .Y(n5472));
  nand_5 g18988(.A(new_n9582), .B(new_n9581), .Y(new_n21337));
  xor_4  g18989(.A(new_n21337), .B(new_n9623), .Y(n5485));
  nand_5 g18990(.A(new_n20720), .B(new_n20697), .Y(new_n21339));
  xor_4  g18991(.A(new_n21339), .B(new_n20715), .Y(n5524));
  nor_5  g18992(.A(new_n18739), .B(new_n6760), .Y(new_n21341));
  nand_5 g18993(.A(new_n21341), .B(new_n6752), .Y(new_n21342));
  nor_5  g18994(.A(new_n21342), .B(new_n6746), .Y(new_n21343));
  nand_5 g18995(.A(new_n21343), .B(new_n6740), .Y(new_n21344));
  nor_5  g18996(.A(new_n21344), .B(new_n6731), .Y(new_n21345));
  nand_5 g18997(.A(new_n21345), .B(new_n6726), .Y(new_n21346));
  nor_5  g18998(.A(new_n21346), .B(new_n6717), .Y(new_n21347));
  nand_5 g18999(.A(new_n21347), .B(new_n6709), .Y(new_n21348));
  xor_4  g19000(.A(new_n21348), .B(new_n15343), .Y(new_n21349_1));
  nor_5  g19001(.A(new_n21349_1), .B(new_n15712), .Y(new_n21350));
  not_8  g19002(.A(new_n21350), .Y(new_n21351));
  nand_5 g19003(.A(new_n21349_1), .B(new_n15712), .Y(new_n21352));
  nand_5 g19004(.A(new_n21352), .B(new_n21351), .Y(new_n21353));
  xor_4  g19005(.A(new_n21347), .B(new_n6708), .Y(new_n21354));
  or_5   g19006(.A(new_n21354), .B(new_n15715), .Y(new_n21355));
  nand_5 g19007(.A(new_n21354), .B(new_n15715), .Y(new_n21356));
  xor_4  g19008(.A(new_n21346), .B(new_n6719), .Y(new_n21357));
  or_5   g19009(.A(new_n21357), .B(new_n15720), .Y(new_n21358));
  nand_5 g19010(.A(new_n21357), .B(new_n15720), .Y(new_n21359));
  not_8  g19011(.A(new_n21345), .Y(new_n21360));
  nand_5 g19012(.A(new_n21360), .B(new_n6724), .Y(new_n21361));
  and_5  g19013(.A(new_n21361), .B(new_n21346), .Y(new_n21362));
  nand_5 g19014(.A(new_n21362), .B(new_n15724), .Y(new_n21363));
  or_5   g19015(.A(new_n21362), .B(new_n15724), .Y(new_n21364));
  nand_5 g19016(.A(new_n21344), .B(new_n6731), .Y(new_n21365_1));
  and_5  g19017(.A(new_n21365_1), .B(new_n21360), .Y(new_n21366));
  nand_5 g19018(.A(new_n21366), .B(new_n15729), .Y(new_n21367_1));
  or_5   g19019(.A(new_n21366), .B(new_n15729), .Y(new_n21368));
  not_8  g19020(.A(new_n21343), .Y(new_n21369));
  nand_5 g19021(.A(new_n21369), .B(new_n6738), .Y(new_n21370));
  and_5  g19022(.A(new_n21370), .B(new_n21344), .Y(new_n21371));
  nand_5 g19023(.A(new_n21371), .B(new_n15734), .Y(new_n21372));
  or_5   g19024(.A(new_n21371), .B(new_n15734), .Y(new_n21373));
  nand_5 g19025(.A(new_n21342), .B(new_n6746), .Y(new_n21374));
  and_5  g19026(.A(new_n21374), .B(new_n21369), .Y(new_n21375));
  nand_5 g19027(.A(new_n21375), .B(new_n15739), .Y(new_n21376));
  or_5   g19028(.A(new_n21375), .B(new_n15739), .Y(new_n21377));
  or_5   g19029(.A(new_n21341), .B(new_n6752), .Y(new_n21378));
  nand_5 g19030(.A(new_n21378), .B(new_n21342), .Y(new_n21379));
  not_8  g19031(.A(new_n19980), .Y(new_n21380));
  nand_5 g19032(.A(new_n19983), .B(new_n21380), .Y(new_n21381));
  nand_5 g19033(.A(new_n21381), .B(new_n19982), .Y(new_n21382));
  or_5   g19034(.A(new_n21382), .B(new_n21379), .Y(new_n21383));
  nand_5 g19035(.A(new_n21382), .B(new_n21379), .Y(new_n21384));
  nand_5 g19036(.A(new_n21384), .B(new_n14979), .Y(new_n21385));
  nand_5 g19037(.A(new_n21385), .B(new_n21383), .Y(new_n21386));
  nand_5 g19038(.A(new_n21386), .B(new_n21377), .Y(new_n21387));
  nand_5 g19039(.A(new_n21387), .B(new_n21376), .Y(new_n21388));
  nand_5 g19040(.A(new_n21388), .B(new_n21373), .Y(new_n21389));
  nand_5 g19041(.A(new_n21389), .B(new_n21372), .Y(new_n21390));
  nand_5 g19042(.A(new_n21390), .B(new_n21368), .Y(new_n21391));
  nand_5 g19043(.A(new_n21391), .B(new_n21367_1), .Y(new_n21392));
  nand_5 g19044(.A(new_n21392), .B(new_n21364), .Y(new_n21393));
  nand_5 g19045(.A(new_n21393), .B(new_n21363), .Y(new_n21394));
  nand_5 g19046(.A(new_n21394), .B(new_n21359), .Y(new_n21395));
  nand_5 g19047(.A(new_n21395), .B(new_n21358), .Y(new_n21396_1));
  nand_5 g19048(.A(new_n21396_1), .B(new_n21356), .Y(new_n21397));
  nand_5 g19049(.A(new_n21397), .B(new_n21355), .Y(new_n21398_1));
  xor_4  g19050(.A(new_n21398_1), .B(new_n21353), .Y(new_n21399_1));
  nand_5 g19051(.A(new_n21399_1), .B(new_n5368), .Y(new_n21400));
  or_5   g19052(.A(new_n21399_1), .B(new_n5368), .Y(new_n21401));
  nand_5 g19053(.A(new_n21356), .B(new_n21355), .Y(new_n21402));
  xor_4  g19054(.A(new_n21402), .B(new_n21396_1), .Y(new_n21403));
  not_8  g19055(.A(new_n21403), .Y(new_n21404_1));
  or_5   g19056(.A(new_n21404_1), .B(new_n5576), .Y(new_n21405));
  nand_5 g19057(.A(new_n21404_1), .B(new_n5576), .Y(new_n21406));
  nand_5 g19058(.A(new_n21359), .B(new_n21358), .Y(new_n21407));
  xor_4  g19059(.A(new_n21407), .B(new_n21394), .Y(new_n21408));
  nand_5 g19060(.A(new_n21408), .B(new_n5582), .Y(new_n21409));
  not_8  g19061(.A(new_n21409), .Y(new_n21410));
  nor_5  g19062(.A(new_n21408), .B(new_n5582), .Y(new_n21411));
  nand_5 g19063(.A(new_n21364), .B(new_n21363), .Y(new_n21412));
  xor_4  g19064(.A(new_n21412), .B(new_n21392), .Y(new_n21413));
  nand_5 g19065(.A(new_n21413), .B(new_n5590), .Y(new_n21414));
  not_8  g19066(.A(new_n21414), .Y(new_n21415));
  nor_5  g19067(.A(new_n21413), .B(new_n5590), .Y(new_n21416));
  nand_5 g19068(.A(new_n21368), .B(new_n21367_1), .Y(new_n21417));
  xor_4  g19069(.A(new_n21417), .B(new_n21390), .Y(new_n21418));
  nand_5 g19070(.A(new_n21418), .B(new_n5597), .Y(new_n21419));
  not_8  g19071(.A(new_n21419), .Y(new_n21420));
  nor_5  g19072(.A(new_n21418), .B(new_n5597), .Y(new_n21421));
  nand_5 g19073(.A(new_n21373), .B(new_n21372), .Y(new_n21422));
  xor_4  g19074(.A(new_n21422), .B(new_n21388), .Y(new_n21423));
  nand_5 g19075(.A(new_n21423), .B(new_n5604), .Y(new_n21424));
  not_8  g19076(.A(new_n21424), .Y(new_n21425));
  nor_5  g19077(.A(new_n21423), .B(new_n5604), .Y(new_n21426));
  nand_5 g19078(.A(new_n21377), .B(new_n21376), .Y(new_n21427));
  xor_4  g19079(.A(new_n21427), .B(new_n21386), .Y(new_n21428));
  nand_5 g19080(.A(new_n21428), .B(new_n5611), .Y(new_n21429));
  not_8  g19081(.A(new_n21429), .Y(new_n21430));
  nor_5  g19082(.A(new_n21428), .B(new_n5611), .Y(new_n21431));
  nand_5 g19083(.A(new_n21384), .B(new_n21383), .Y(new_n21432));
  xor_4  g19084(.A(new_n21432), .B(new_n14977_1), .Y(new_n21433));
  nand_5 g19085(.A(new_n21433), .B(new_n5619), .Y(new_n21434));
  or_5   g19086(.A(new_n21433), .B(new_n5619), .Y(new_n21435));
  nand_5 g19087(.A(new_n19987), .B(new_n19977), .Y(new_n21436));
  nand_5 g19088(.A(new_n21436), .B(new_n19986), .Y(new_n21437));
  nand_5 g19089(.A(new_n21437), .B(new_n21435), .Y(new_n21438));
  nand_5 g19090(.A(new_n21438), .B(new_n21434), .Y(new_n21439));
  nor_5  g19091(.A(new_n21439), .B(new_n21431), .Y(new_n21440));
  nor_5  g19092(.A(new_n21440), .B(new_n21430), .Y(new_n21441));
  nor_5  g19093(.A(new_n21441), .B(new_n21426), .Y(new_n21442));
  nor_5  g19094(.A(new_n21442), .B(new_n21425), .Y(new_n21443));
  nor_5  g19095(.A(new_n21443), .B(new_n21421), .Y(new_n21444));
  nor_5  g19096(.A(new_n21444), .B(new_n21420), .Y(new_n21445));
  nor_5  g19097(.A(new_n21445), .B(new_n21416), .Y(new_n21446_1));
  nor_5  g19098(.A(new_n21446_1), .B(new_n21415), .Y(new_n21447));
  nor_5  g19099(.A(new_n21447), .B(new_n21411), .Y(new_n21448));
  nor_5  g19100(.A(new_n21448), .B(new_n21410), .Y(new_n21449));
  not_8  g19101(.A(new_n21449), .Y(new_n21450));
  nand_5 g19102(.A(new_n21450), .B(new_n21406), .Y(new_n21451));
  nand_5 g19103(.A(new_n21451), .B(new_n21405), .Y(new_n21452));
  nand_5 g19104(.A(new_n21452), .B(new_n21401), .Y(new_n21453));
  nand_5 g19105(.A(new_n21453), .B(new_n21400), .Y(new_n21454));
  nor_5  g19106(.A(new_n21348), .B(new_n15344), .Y(new_n21455));
  nand_5 g19107(.A(new_n21398_1), .B(new_n21352), .Y(new_n21456));
  nand_5 g19108(.A(new_n21456), .B(new_n21351), .Y(new_n21457));
  nor_5  g19109(.A(new_n21457), .B(new_n21455), .Y(new_n21458));
  and_5  g19110(.A(new_n21458), .B(new_n21454), .Y(n23066));
  nor_5  g19111(.A(new_n21458), .B(new_n21454), .Y(new_n21460));
  or_5   g19112(.A(new_n21460), .B(n23066), .Y(n5564));
  nand_5 g19113(.A(new_n7925), .B(new_n7926), .Y(new_n21462));
  xnor_4 g19114(.A(new_n21462), .B(new_n7940), .Y(n5593));
  nand_5 g19115(.A(new_n18648), .B(new_n16197), .Y(new_n21464));
  or_5   g19116(.A(new_n18648), .B(new_n16197), .Y(new_n21465));
  nand_5 g19117(.A(new_n18635_1), .B(new_n16203), .Y(new_n21466));
  or_5   g19118(.A(new_n18635_1), .B(new_n16203), .Y(new_n21467));
  nand_5 g19119(.A(new_n17544), .B(new_n16209), .Y(new_n21468));
  or_5   g19120(.A(new_n17544), .B(new_n16209), .Y(new_n21469));
  nand_5 g19121(.A(new_n19544), .B(new_n19542), .Y(new_n21470));
  nand_5 g19122(.A(new_n21470), .B(new_n19543), .Y(new_n21471_1));
  nand_5 g19123(.A(new_n21471_1), .B(new_n21469), .Y(new_n21472_1));
  nand_5 g19124(.A(new_n21472_1), .B(new_n21468), .Y(new_n21473));
  nand_5 g19125(.A(new_n21473), .B(new_n21467), .Y(new_n21474));
  nand_5 g19126(.A(new_n21474), .B(new_n21466), .Y(new_n21475));
  nand_5 g19127(.A(new_n21475), .B(new_n21465), .Y(new_n21476));
  nand_5 g19128(.A(new_n21476), .B(new_n21464), .Y(new_n21477));
  nand_5 g19129(.A(new_n20031), .B(new_n16191), .Y(new_n21478));
  not_8  g19130(.A(new_n21478), .Y(new_n21479));
  nor_5  g19131(.A(new_n20031), .B(new_n16191), .Y(new_n21480));
  nor_5  g19132(.A(new_n21480), .B(new_n21479), .Y(new_n21481));
  xor_4  g19133(.A(new_n21481), .B(new_n21477), .Y(n5603));
  nand_5 g19134(.A(n25119), .B(new_n2568), .Y(new_n21483));
  nand_5 g19135(.A(new_n9834), .B(n13783), .Y(new_n21484));
  nand_5 g19136(.A(new_n2475), .B(n1163), .Y(new_n21485));
  nand_5 g19137(.A(n26660), .B(new_n9778_1), .Y(new_n21486));
  nand_5 g19138(.A(n18537), .B(new_n2412), .Y(new_n21487));
  nand_5 g19139(.A(new_n9757), .B(n3018), .Y(new_n21488));
  nand_5 g19140(.A(new_n20349_1), .B(new_n20346), .Y(new_n21489_1));
  nand_5 g19141(.A(new_n21489_1), .B(new_n20348), .Y(new_n21490));
  nand_5 g19142(.A(new_n21490), .B(new_n21488), .Y(new_n21491));
  nand_5 g19143(.A(new_n21491), .B(new_n21487), .Y(new_n21492));
  nand_5 g19144(.A(new_n21492), .B(new_n21486), .Y(new_n21493));
  nand_5 g19145(.A(new_n21493), .B(new_n21485), .Y(new_n21494));
  nand_5 g19146(.A(new_n21494), .B(new_n21484), .Y(new_n21495));
  nand_5 g19147(.A(new_n21495), .B(new_n21483), .Y(new_n21496));
  nand_5 g19148(.A(n21997), .B(new_n8565), .Y(new_n21497));
  nand_5 g19149(.A(new_n18133), .B(n1654), .Y(new_n21498));
  nand_5 g19150(.A(new_n21498), .B(new_n21497), .Y(new_n21499));
  xor_4  g19151(.A(new_n21499), .B(new_n21496), .Y(new_n21500));
  nand_5 g19152(.A(new_n21500), .B(new_n3206), .Y(new_n21501));
  not_8  g19153(.A(new_n21501), .Y(new_n21502));
  nor_5  g19154(.A(new_n21500), .B(new_n3206), .Y(new_n21503));
  nand_5 g19155(.A(new_n21484), .B(new_n21483), .Y(new_n21504));
  xor_4  g19156(.A(new_n21504), .B(new_n21494), .Y(new_n21505));
  nand_5 g19157(.A(new_n21505), .B(new_n3213), .Y(new_n21506));
  not_8  g19158(.A(new_n21506), .Y(new_n21507));
  nor_5  g19159(.A(new_n21505), .B(new_n3213), .Y(new_n21508));
  nand_5 g19160(.A(new_n21486), .B(new_n21485), .Y(new_n21509));
  xor_4  g19161(.A(new_n21509), .B(new_n21492), .Y(new_n21510));
  nand_5 g19162(.A(new_n21510), .B(new_n3220), .Y(new_n21511));
  not_8  g19163(.A(new_n21511), .Y(new_n21512));
  nor_5  g19164(.A(new_n21510), .B(new_n3220), .Y(new_n21513));
  nand_5 g19165(.A(new_n21488), .B(new_n21487), .Y(new_n21514));
  xor_4  g19166(.A(new_n21514), .B(new_n21490), .Y(new_n21515));
  nand_5 g19167(.A(new_n21515), .B(new_n3227), .Y(new_n21516));
  not_8  g19168(.A(new_n21516), .Y(new_n21517));
  nor_5  g19169(.A(new_n21515), .B(new_n3227), .Y(new_n21518));
  nor_5  g19170(.A(new_n20355_1), .B(new_n20344), .Y(new_n21519));
  nor_5  g19171(.A(new_n21519), .B(new_n20353), .Y(new_n21520));
  nor_5  g19172(.A(new_n21520), .B(new_n21518), .Y(new_n21521));
  nor_5  g19173(.A(new_n21521), .B(new_n21517), .Y(new_n21522));
  nor_5  g19174(.A(new_n21522), .B(new_n21513), .Y(new_n21523));
  nor_5  g19175(.A(new_n21523), .B(new_n21512), .Y(new_n21524));
  nor_5  g19176(.A(new_n21524), .B(new_n21508), .Y(new_n21525_1));
  nor_5  g19177(.A(new_n21525_1), .B(new_n21507), .Y(new_n21526));
  nor_5  g19178(.A(new_n21526), .B(new_n21503), .Y(new_n21527));
  nor_5  g19179(.A(new_n21527), .B(new_n21502), .Y(new_n21528));
  nand_5 g19180(.A(new_n21498), .B(new_n21496), .Y(new_n21529));
  nand_5 g19181(.A(new_n21529), .B(new_n21497), .Y(new_n21530));
  not_8  g19182(.A(new_n21530), .Y(new_n21531));
  nand_5 g19183(.A(n17911), .B(new_n8574), .Y(new_n21532));
  nand_5 g19184(.A(new_n18127), .B(n14440), .Y(new_n21533));
  nand_5 g19185(.A(new_n21533), .B(new_n21532), .Y(new_n21534));
  xor_4  g19186(.A(new_n21534), .B(new_n21531), .Y(new_n21535));
  or_5   g19187(.A(new_n21535), .B(new_n3307), .Y(new_n21536));
  not_8  g19188(.A(new_n21536), .Y(new_n21537));
  nand_5 g19189(.A(new_n21535), .B(new_n3307), .Y(new_n21538_1));
  not_8  g19190(.A(new_n21538_1), .Y(new_n21539));
  nor_5  g19191(.A(new_n21539), .B(new_n21537), .Y(new_n21540));
  xor_4  g19192(.A(new_n21540), .B(new_n21528), .Y(n5609));
  nand_5 g19193(.A(new_n15251), .B(new_n15250), .Y(new_n21542));
  xnor_4 g19194(.A(new_n21542), .B(new_n15272), .Y(n5634));
  nand_5 g19195(.A(n3425), .B(new_n8648), .Y(new_n21544));
  nand_5 g19196(.A(new_n8597), .B(n2978), .Y(new_n21545));
  nand_5 g19197(.A(new_n7958), .B(n9967), .Y(new_n21546));
  nand_5 g19198(.A(n23697), .B(new_n3442), .Y(new_n21547));
  nand_5 g19199(.A(new_n20963), .B(new_n20961), .Y(new_n21548));
  nand_5 g19200(.A(new_n21548), .B(new_n20962), .Y(new_n21549_1));
  nand_5 g19201(.A(new_n21549_1), .B(new_n21547), .Y(new_n21550));
  nand_5 g19202(.A(new_n21550), .B(new_n21546), .Y(new_n21551));
  nand_5 g19203(.A(new_n21551), .B(new_n21545), .Y(new_n21552));
  nand_5 g19204(.A(new_n21552), .B(new_n21544), .Y(new_n21553));
  not_8  g19205(.A(new_n21553), .Y(new_n21554));
  nand_5 g19206(.A(new_n21554), .B(new_n8473), .Y(new_n21555));
  nand_5 g19207(.A(new_n21553), .B(new_n8430), .Y(new_n21556));
  nand_5 g19208(.A(new_n21545), .B(new_n21544), .Y(new_n21557));
  xor_4  g19209(.A(new_n21557), .B(new_n21551), .Y(new_n21558));
  or_5   g19210(.A(new_n21558), .B(new_n8479), .Y(new_n21559));
  nand_5 g19211(.A(new_n21558), .B(new_n8479), .Y(new_n21560));
  nand_5 g19212(.A(new_n21547), .B(new_n21546), .Y(new_n21561));
  xor_4  g19213(.A(new_n21561), .B(new_n21549_1), .Y(new_n21562));
  or_5   g19214(.A(new_n21562), .B(new_n8486), .Y(new_n21563));
  nand_5 g19215(.A(new_n21562), .B(new_n8486), .Y(new_n21564));
  not_8  g19216(.A(new_n20959), .Y(new_n21565));
  nor_5  g19217(.A(new_n20968), .B(new_n21565), .Y(new_n21566));
  nor_5  g19218(.A(new_n21566), .B(new_n20967), .Y(new_n21567));
  not_8  g19219(.A(new_n21567), .Y(new_n21568));
  nand_5 g19220(.A(new_n21568), .B(new_n21564), .Y(new_n21569));
  nand_5 g19221(.A(new_n21569), .B(new_n21563), .Y(new_n21570));
  nand_5 g19222(.A(new_n21570), .B(new_n21560), .Y(new_n21571));
  nand_5 g19223(.A(new_n21571), .B(new_n21559), .Y(new_n21572));
  nand_5 g19224(.A(new_n21572), .B(new_n21556), .Y(new_n21573));
  nand_5 g19225(.A(new_n21573), .B(new_n21555), .Y(new_n21574));
  nand_5 g19226(.A(new_n8428), .B(new_n8351), .Y(new_n21575));
  not_8  g19227(.A(new_n21575), .Y(new_n21576));
  nand_5 g19228(.A(new_n21576), .B(new_n21553), .Y(new_n21577));
  nand_5 g19229(.A(new_n21575), .B(new_n21554), .Y(new_n21578));
  nand_5 g19230(.A(new_n21578), .B(new_n21577), .Y(new_n21579));
  xnor_4 g19231(.A(new_n21579), .B(new_n21574), .Y(n5643));
  nand_5 g19232(.A(new_n17639), .B(new_n17046), .Y(new_n21581));
  nand_5 g19233(.A(new_n17638_1), .B(new_n17045), .Y(new_n21582));
  nand_5 g19234(.A(new_n17609), .B(new_n17069_1), .Y(new_n21583));
  nand_5 g19235(.A(new_n17611), .B(new_n17068_1), .Y(new_n21584));
  nand_5 g19236(.A(new_n17614), .B(new_n17076), .Y(new_n21585));
  nand_5 g19237(.A(new_n17616), .B(new_n17075_1), .Y(new_n21586));
  nand_5 g19238(.A(new_n17619), .B(new_n17088), .Y(new_n21587));
  nand_5 g19239(.A(new_n17621), .B(new_n17082), .Y(new_n21588));
  nand_5 g19240(.A(new_n15860), .B(new_n15572), .Y(new_n21589));
  nand_5 g19241(.A(new_n15861), .B(new_n15571), .Y(new_n21590));
  nand_5 g19242(.A(new_n15826), .B(new_n15522), .Y(new_n21591));
  or_5   g19243(.A(new_n15826), .B(new_n15522), .Y(new_n21592));
  not_8  g19244(.A(new_n15532), .Y(new_n21593));
  nor_5  g19245(.A(new_n15839), .B(new_n21593), .Y(new_n21594));
  not_8  g19246(.A(new_n21594), .Y(new_n21595));
  nand_5 g19247(.A(new_n21595), .B(new_n15535), .Y(new_n21596));
  or_5   g19248(.A(new_n21595), .B(new_n15535), .Y(new_n21597));
  nand_5 g19249(.A(new_n21597), .B(new_n15847), .Y(new_n21598));
  nand_5 g19250(.A(new_n21598), .B(new_n21596), .Y(new_n21599_1));
  nand_5 g19251(.A(new_n21599_1), .B(new_n21592), .Y(new_n21600));
  nand_5 g19252(.A(new_n21600), .B(new_n21591), .Y(new_n21601));
  nand_5 g19253(.A(new_n21601), .B(new_n21590), .Y(new_n21602));
  nand_5 g19254(.A(new_n21602), .B(new_n21589), .Y(new_n21603));
  nand_5 g19255(.A(new_n21603), .B(new_n21588), .Y(new_n21604));
  nand_5 g19256(.A(new_n21604), .B(new_n21587), .Y(new_n21605));
  nand_5 g19257(.A(new_n21605), .B(new_n21586), .Y(new_n21606));
  nand_5 g19258(.A(new_n21606), .B(new_n21585), .Y(new_n21607));
  nand_5 g19259(.A(new_n21607), .B(new_n21584), .Y(new_n21608));
  nand_5 g19260(.A(new_n21608), .B(new_n21583), .Y(new_n21609));
  nand_5 g19261(.A(new_n21609), .B(new_n21582), .Y(new_n21610));
  nand_5 g19262(.A(new_n21610), .B(new_n21581), .Y(new_n21611));
  nand_5 g19263(.A(new_n17636), .B(new_n17632), .Y(new_n21612));
  nand_5 g19264(.A(new_n21612), .B(new_n17635), .Y(new_n21613));
  not_8  g19265(.A(new_n21613), .Y(new_n21614));
  nand_5 g19266(.A(n18035), .B(new_n20002), .Y(new_n21615_1));
  nand_5 g19267(.A(new_n12392), .B(n5834), .Y(new_n21616));
  nand_5 g19268(.A(new_n21616), .B(new_n21615_1), .Y(new_n21617));
  xor_4  g19269(.A(new_n21617), .B(new_n21614), .Y(new_n21618));
  not_8  g19270(.A(new_n21618), .Y(new_n21619));
  nand_5 g19271(.A(new_n21619), .B(new_n17118), .Y(new_n21620));
  nand_5 g19272(.A(new_n21618), .B(new_n17119_1), .Y(new_n21621));
  nand_5 g19273(.A(new_n21621), .B(new_n21620), .Y(new_n21622));
  xor_4  g19274(.A(new_n21622), .B(new_n21611), .Y(n5680));
  nand_5 g19275(.A(new_n16737), .B(new_n2968), .Y(new_n21624));
  nand_5 g19276(.A(new_n21624), .B(new_n16736), .Y(new_n21625));
  xor_4  g19277(.A(new_n21625), .B(new_n16742), .Y(n5687));
  nor_5  g19278(.A(new_n17960), .B(new_n17959_1), .Y(new_n21627));
  xor_4  g19279(.A(new_n21627), .B(new_n17970), .Y(n5700));
  nand_5 g19280(.A(new_n12037), .B(new_n12036), .Y(new_n21629));
  xor_4  g19281(.A(new_n21629), .B(new_n12103), .Y(n5732));
  not_8  g19282(.A(new_n20852), .Y(new_n21631));
  nand_5 g19283(.A(new_n20865), .B(new_n21631), .Y(new_n21632));
  nand_5 g19284(.A(new_n21632), .B(new_n20864), .Y(new_n21633));
  nand_5 g19285(.A(new_n20850), .B(new_n20843), .Y(new_n21634));
  nand_5 g19286(.A(new_n21634), .B(new_n20849), .Y(new_n21635));
  nand_5 g19287(.A(new_n20846), .B(new_n20840), .Y(new_n21636));
  nand_5 g19288(.A(new_n21636), .B(new_n20845), .Y(new_n21637_1));
  nand_5 g19289(.A(new_n8165), .B(new_n5709), .Y(new_n21638));
  nand_5 g19290(.A(n23775), .B(n8381), .Y(new_n21639));
  nand_5 g19291(.A(new_n21639), .B(new_n21638), .Y(new_n21640));
  xor_4  g19292(.A(new_n21640), .B(new_n21637_1), .Y(new_n21641));
  nand_5 g19293(.A(new_n21641), .B(new_n2397), .Y(new_n21642));
  or_5   g19294(.A(new_n21641), .B(new_n2397), .Y(new_n21643));
  nand_5 g19295(.A(new_n21643), .B(new_n21642), .Y(new_n21644));
  xor_4  g19296(.A(new_n21644), .B(new_n21635), .Y(new_n21645_1));
  not_8  g19297(.A(new_n21645_1), .Y(new_n21646));
  nand_5 g19298(.A(new_n20861), .B(new_n20855), .Y(new_n21647));
  nand_5 g19299(.A(new_n21647), .B(new_n20860), .Y(new_n21648));
  nand_5 g19300(.A(n8869), .B(new_n2498), .Y(new_n21649_1));
  nand_5 g19301(.A(new_n8035), .B(n6385), .Y(new_n21650));
  nand_5 g19302(.A(new_n21650), .B(new_n21649_1), .Y(new_n21651));
  xnor_4 g19303(.A(new_n21651), .B(new_n21648), .Y(new_n21652));
  nand_5 g19304(.A(new_n21652), .B(new_n21646), .Y(new_n21653));
  or_5   g19305(.A(new_n21652), .B(new_n21646), .Y(new_n21654_1));
  nand_5 g19306(.A(new_n21654_1), .B(new_n21653), .Y(new_n21655));
  xnor_4 g19307(.A(new_n21655), .B(new_n21633), .Y(n5742));
  nand_5 g19308(.A(new_n15523), .B(new_n15526), .Y(new_n21657));
  xor_4  g19309(.A(new_n21657), .B(new_n15541), .Y(n5765));
  nand_5 g19310(.A(new_n14268), .B(new_n14269), .Y(new_n21659));
  xor_4  g19311(.A(new_n21659), .B(new_n14319), .Y(n5776));
  nand_5 g19312(.A(new_n2936), .B(new_n2935), .Y(new_n21661));
  xnor_4 g19313(.A(new_n21661), .B(new_n2988), .Y(n5782));
  nand_5 g19314(.A(new_n21639), .B(new_n21637_1), .Y(new_n21663));
  nand_5 g19315(.A(new_n21663), .B(new_n21638), .Y(new_n21664));
  not_8  g19316(.A(new_n21664), .Y(new_n21665_1));
  nand_5 g19317(.A(new_n21665_1), .B(n7057), .Y(new_n21666));
  nand_5 g19318(.A(new_n21664), .B(new_n9760), .Y(new_n21667));
  nand_5 g19319(.A(new_n21667), .B(new_n21666), .Y(new_n21668));
  xor_4  g19320(.A(new_n21668), .B(new_n8162), .Y(new_n21669));
  nand_5 g19321(.A(new_n21643), .B(new_n21635), .Y(new_n21670));
  nand_5 g19322(.A(new_n21670), .B(new_n21642), .Y(new_n21671));
  nand_5 g19323(.A(new_n21671), .B(new_n21669), .Y(new_n21672));
  or_5   g19324(.A(new_n21671), .B(new_n21669), .Y(new_n21673));
  nand_5 g19325(.A(new_n21673), .B(new_n2408), .Y(new_n21674_1));
  nand_5 g19326(.A(new_n21674_1), .B(new_n21672), .Y(new_n21675));
  nand_5 g19327(.A(new_n21666), .B(new_n8162), .Y(new_n21676));
  nand_5 g19328(.A(new_n21676), .B(new_n21667), .Y(new_n21677));
  xor_4  g19329(.A(new_n21677), .B(new_n8159_1), .Y(new_n21678));
  xor_4  g19330(.A(new_n21678), .B(new_n9757), .Y(new_n21679));
  or_5   g19331(.A(new_n21679), .B(new_n2419), .Y(new_n21680_1));
  nand_5 g19332(.A(new_n21679), .B(new_n2419), .Y(new_n21681));
  nand_5 g19333(.A(new_n21681), .B(new_n21680_1), .Y(new_n21682));
  xor_4  g19334(.A(new_n21682), .B(new_n21675), .Y(new_n21683));
  nand_5 g19335(.A(new_n3084), .B(n1118), .Y(new_n21684));
  nand_5 g19336(.A(n10053), .B(new_n3042), .Y(new_n21685_1));
  nand_5 g19337(.A(n25974), .B(new_n3085), .Y(new_n21686));
  nand_5 g19338(.A(new_n3047), .B(n8399), .Y(new_n21687_1));
  nand_5 g19339(.A(new_n3090), .B(n1630), .Y(new_n21688));
  nand_5 g19340(.A(n9507), .B(new_n3050), .Y(new_n21689));
  nand_5 g19341(.A(n26979), .B(new_n3158), .Y(new_n21690));
  nand_5 g19342(.A(new_n21690), .B(new_n21689), .Y(new_n21691));
  nand_5 g19343(.A(new_n21691), .B(new_n21688), .Y(new_n21692));
  nand_5 g19344(.A(new_n21692), .B(new_n21687_1), .Y(new_n21693));
  nand_5 g19345(.A(new_n21693), .B(new_n21686), .Y(new_n21694));
  nand_5 g19346(.A(new_n21694), .B(new_n21685_1), .Y(new_n21695));
  nand_5 g19347(.A(new_n21695), .B(new_n21684), .Y(new_n21696));
  nand_5 g19348(.A(new_n3079), .B(n12811), .Y(new_n21697));
  nand_5 g19349(.A(n19514), .B(new_n3039), .Y(new_n21698));
  nand_5 g19350(.A(new_n21698), .B(new_n21697), .Y(new_n21699));
  xor_4  g19351(.A(new_n21699), .B(new_n21696), .Y(new_n21700));
  nand_5 g19352(.A(new_n21700), .B(new_n21683), .Y(new_n21701));
  not_8  g19353(.A(new_n21701), .Y(new_n21702));
  nor_5  g19354(.A(new_n21700), .B(new_n21683), .Y(new_n21703));
  nand_5 g19355(.A(new_n21673), .B(new_n21672), .Y(new_n21704));
  xor_4  g19356(.A(new_n21704), .B(new_n2427), .Y(new_n21705));
  not_8  g19357(.A(new_n21705), .Y(new_n21706));
  nand_5 g19358(.A(new_n21685_1), .B(new_n21684), .Y(new_n21707));
  xor_4  g19359(.A(new_n21707), .B(new_n21694), .Y(new_n21708));
  or_5   g19360(.A(new_n21708), .B(new_n21706), .Y(new_n21709));
  nand_5 g19361(.A(new_n21708), .B(new_n21706), .Y(new_n21710));
  nand_5 g19362(.A(new_n21687_1), .B(new_n21686), .Y(new_n21711));
  xor_4  g19363(.A(new_n21711), .B(new_n21692), .Y(new_n21712));
  or_5   g19364(.A(new_n21712), .B(new_n21645_1), .Y(new_n21713));
  nand_5 g19365(.A(new_n21712), .B(new_n21645_1), .Y(new_n21714));
  not_8  g19366(.A(new_n20854), .Y(new_n21715));
  xor_4  g19367(.A(n26979), .B(new_n3158), .Y(new_n21716));
  nor_5  g19368(.A(new_n21716), .B(new_n21715), .Y(new_n21717_1));
  nand_5 g19369(.A(new_n21689), .B(new_n21688), .Y(new_n21718));
  xnor_4 g19370(.A(new_n21718), .B(new_n21690), .Y(new_n21719_1));
  nand_5 g19371(.A(new_n21719_1), .B(new_n21717_1), .Y(new_n21720));
  not_8  g19372(.A(new_n21720), .Y(new_n21721));
  nor_5  g19373(.A(new_n21719_1), .B(new_n21717_1), .Y(new_n21722));
  nor_5  g19374(.A(new_n21722), .B(new_n20852), .Y(new_n21723));
  nor_5  g19375(.A(new_n21723), .B(new_n21721), .Y(new_n21724));
  not_8  g19376(.A(new_n21724), .Y(new_n21725));
  nand_5 g19377(.A(new_n21725), .B(new_n21714), .Y(new_n21726));
  nand_5 g19378(.A(new_n21726), .B(new_n21713), .Y(new_n21727));
  nand_5 g19379(.A(new_n21727), .B(new_n21710), .Y(new_n21728));
  nand_5 g19380(.A(new_n21728), .B(new_n21709), .Y(new_n21729));
  nor_5  g19381(.A(new_n21729), .B(new_n21703), .Y(new_n21730));
  nor_5  g19382(.A(new_n21730), .B(new_n21702), .Y(new_n21731));
  nand_5 g19383(.A(new_n21681), .B(new_n21675), .Y(new_n21732));
  nand_5 g19384(.A(new_n21732), .B(new_n21680_1), .Y(new_n21733));
  nand_5 g19385(.A(n18537), .B(n4376), .Y(new_n21734));
  nor_5  g19386(.A(n18537), .B(n4376), .Y(new_n21735_1));
  or_5   g19387(.A(new_n21735_1), .B(new_n21677), .Y(new_n21736));
  nand_5 g19388(.A(new_n21736), .B(new_n21734), .Y(new_n21737));
  nand_5 g19389(.A(new_n8156), .B(new_n9778_1), .Y(new_n21738));
  nand_5 g19390(.A(n18901), .B(n1163), .Y(new_n21739));
  nand_5 g19391(.A(new_n21739), .B(new_n21738), .Y(new_n21740));
  xor_4  g19392(.A(new_n21740), .B(new_n21737), .Y(new_n21741));
  or_5   g19393(.A(new_n21741), .B(new_n2483), .Y(new_n21742));
  nand_5 g19394(.A(new_n21741), .B(new_n2483), .Y(new_n21743));
  nand_5 g19395(.A(new_n21743), .B(new_n21742), .Y(new_n21744));
  xor_4  g19396(.A(new_n21744), .B(new_n21733), .Y(new_n21745));
  not_8  g19397(.A(new_n21745), .Y(new_n21746));
  nand_5 g19398(.A(new_n21698), .B(new_n21696), .Y(new_n21747));
  nand_5 g19399(.A(new_n21747), .B(new_n21697), .Y(new_n21748));
  not_8  g19400(.A(new_n21748), .Y(new_n21749_1));
  nand_5 g19401(.A(new_n3073), .B(n7099), .Y(new_n21750_1));
  nand_5 g19402(.A(n23068), .B(new_n3034), .Y(new_n21751));
  nand_5 g19403(.A(new_n21751), .B(new_n21750_1), .Y(new_n21752));
  xor_4  g19404(.A(new_n21752), .B(new_n21749_1), .Y(new_n21753_1));
  or_5   g19405(.A(new_n21753_1), .B(new_n21746), .Y(new_n21754));
  not_8  g19406(.A(new_n21754), .Y(new_n21755));
  nand_5 g19407(.A(new_n21753_1), .B(new_n21746), .Y(new_n21756));
  not_8  g19408(.A(new_n21756), .Y(new_n21757));
  nor_5  g19409(.A(new_n21757), .B(new_n21755), .Y(new_n21758));
  xor_4  g19410(.A(new_n21758), .B(new_n21731), .Y(n5833));
  nand_5 g19411(.A(new_n14281), .B(new_n14282), .Y(new_n21760));
  xor_4  g19412(.A(new_n21760), .B(new_n14315), .Y(n5840));
  nor_5  g19413(.A(new_n21518), .B(new_n21517), .Y(new_n21762));
  xor_4  g19414(.A(new_n21762), .B(new_n21520), .Y(n5841));
  nand_5 g19415(.A(new_n14807), .B(new_n14808), .Y(new_n21764));
  xor_4  g19416(.A(new_n21764), .B(new_n14809), .Y(n5850));
  nand_5 g19417(.A(new_n21589), .B(new_n21590), .Y(new_n21766));
  xor_4  g19418(.A(new_n21766), .B(new_n21601), .Y(n5903));
  nand_5 g19419(.A(new_n21049), .B(new_n21030), .Y(new_n21768));
  nand_5 g19420(.A(new_n21768), .B(new_n21048), .Y(new_n21769));
  nand_5 g19421(.A(new_n21038), .B(new_n21032), .Y(new_n21770));
  nand_5 g19422(.A(new_n21770), .B(new_n21037), .Y(new_n21771));
  nor_5  g19423(.A(new_n21034_1), .B(n26752), .Y(new_n21772));
  not_8  g19424(.A(new_n21772), .Y(new_n21773));
  nand_5 g19425(.A(new_n21034_1), .B(n26752), .Y(new_n21774));
  and_5  g19426(.A(new_n21774), .B(new_n21773), .Y(new_n21775));
  or_5   g19427(.A(new_n21775), .B(new_n10108), .Y(new_n21776));
  nand_5 g19428(.A(new_n21775), .B(new_n10108), .Y(new_n21777));
  nand_5 g19429(.A(new_n21777), .B(new_n21776), .Y(new_n21778));
  xor_4  g19430(.A(new_n21778), .B(new_n21771), .Y(new_n21779_1));
  not_8  g19431(.A(new_n21779_1), .Y(new_n21780));
  nand_5 g19432(.A(new_n21045), .B(new_n21043), .Y(new_n21781));
  nand_5 g19433(.A(new_n21781), .B(new_n21044), .Y(new_n21782));
  nand_5 g19434(.A(new_n18850), .B(n19042), .Y(new_n21783));
  nand_5 g19435(.A(new_n18852), .B(new_n7819), .Y(new_n21784_1));
  nand_5 g19436(.A(new_n21784_1), .B(new_n21783), .Y(new_n21785));
  xor_4  g19437(.A(new_n21785), .B(new_n21782), .Y(new_n21786));
  or_5   g19438(.A(new_n21786), .B(new_n21780), .Y(new_n21787));
  nand_5 g19439(.A(new_n21786), .B(new_n21780), .Y(new_n21788));
  nand_5 g19440(.A(new_n21788), .B(new_n21787), .Y(new_n21789));
  xnor_4 g19441(.A(new_n21789), .B(new_n21769), .Y(n5904));
  nand_5 g19442(.A(n23529), .B(new_n3108), .Y(new_n21791));
  nand_5 g19443(.A(new_n3068), .B(n10710), .Y(new_n21792));
  nand_5 g19444(.A(n24620), .B(new_n3072), .Y(new_n21793));
  nand_5 g19445(.A(new_n3035), .B(n20929), .Y(new_n21794));
  nand_5 g19446(.A(new_n3078), .B(n5211), .Y(new_n21795));
  nand_5 g19447(.A(n8006), .B(new_n3038), .Y(new_n21796));
  nand_5 g19448(.A(new_n3136_1), .B(n12956), .Y(new_n21797));
  nand_5 g19449(.A(n25074), .B(new_n3043), .Y(new_n21798));
  nand_5 g19450(.A(n18295), .B(new_n3086), .Y(new_n21799));
  nand_5 g19451(.A(new_n3046), .B(n16396), .Y(new_n21800_1));
  nand_5 g19452(.A(new_n3089_1), .B(n6502), .Y(new_n21801));
  nand_5 g19453(.A(n9399), .B(new_n3051), .Y(new_n21802));
  nand_5 g19454(.A(new_n3159), .B(n2088), .Y(new_n21803));
  nand_5 g19455(.A(new_n21803), .B(new_n21802), .Y(new_n21804));
  nand_5 g19456(.A(new_n21804), .B(new_n21801), .Y(new_n21805));
  nand_5 g19457(.A(new_n21805), .B(new_n21800_1), .Y(new_n21806));
  nand_5 g19458(.A(new_n21806), .B(new_n21799), .Y(new_n21807));
  nand_5 g19459(.A(new_n21807), .B(new_n21798), .Y(new_n21808));
  nand_5 g19460(.A(new_n21808), .B(new_n21797), .Y(new_n21809));
  nand_5 g19461(.A(new_n21809), .B(new_n21796), .Y(new_n21810));
  nand_5 g19462(.A(new_n21810), .B(new_n21795), .Y(new_n21811));
  nand_5 g19463(.A(new_n21811), .B(new_n21794), .Y(new_n21812));
  nand_5 g19464(.A(new_n21812), .B(new_n21793), .Y(new_n21813));
  nand_5 g19465(.A(new_n21813), .B(new_n21792), .Y(new_n21814));
  nand_5 g19466(.A(new_n21814), .B(new_n21791), .Y(new_n21815));
  nand_5 g19467(.A(n19701), .B(new_n3194), .Y(new_n21816));
  nand_5 g19468(.A(new_n3186), .B(n11841), .Y(new_n21817));
  nand_5 g19469(.A(new_n21817), .B(new_n21816), .Y(new_n21818));
  xor_4  g19470(.A(new_n21818), .B(new_n21815), .Y(new_n21819));
  or_5   g19471(.A(new_n21819), .B(new_n11766), .Y(new_n21820_1));
  nand_5 g19472(.A(new_n21819), .B(new_n11766), .Y(new_n21821));
  nand_5 g19473(.A(new_n21792), .B(new_n21791), .Y(new_n21822));
  xor_4  g19474(.A(new_n21822), .B(new_n21813), .Y(new_n21823));
  or_5   g19475(.A(new_n21823), .B(new_n11773), .Y(new_n21824));
  nand_5 g19476(.A(new_n21823), .B(new_n11773), .Y(new_n21825));
  nand_5 g19477(.A(new_n21794), .B(new_n21793), .Y(new_n21826));
  xor_4  g19478(.A(new_n21826), .B(new_n21811), .Y(new_n21827));
  or_5   g19479(.A(new_n21827), .B(new_n11780), .Y(new_n21828));
  nand_5 g19480(.A(new_n21827), .B(new_n11780), .Y(new_n21829));
  nand_5 g19481(.A(new_n21796), .B(new_n21795), .Y(new_n21830));
  xor_4  g19482(.A(new_n21830), .B(new_n21809), .Y(new_n21831));
  or_5   g19483(.A(new_n21831), .B(new_n11787), .Y(new_n21832_1));
  nand_5 g19484(.A(new_n21831), .B(new_n11787), .Y(new_n21833));
  nand_5 g19485(.A(new_n21798), .B(new_n21797), .Y(new_n21834));
  xor_4  g19486(.A(new_n21834), .B(new_n21807), .Y(new_n21835));
  or_5   g19487(.A(new_n21835), .B(new_n11794), .Y(new_n21836));
  nand_5 g19488(.A(new_n21835), .B(new_n11794), .Y(new_n21837));
  nand_5 g19489(.A(new_n21800_1), .B(new_n21799), .Y(new_n21838));
  xor_4  g19490(.A(new_n21838), .B(new_n21805), .Y(new_n21839_1));
  or_5   g19491(.A(new_n21839_1), .B(new_n11802), .Y(new_n21840));
  nand_5 g19492(.A(new_n21839_1), .B(new_n11802), .Y(new_n21841));
  nand_5 g19493(.A(n15780), .B(new_n3163), .Y(new_n21842));
  nand_5 g19494(.A(new_n21842), .B(new_n21803), .Y(new_n21843));
  nand_5 g19495(.A(new_n21843), .B(new_n11805), .Y(new_n21844));
  not_8  g19496(.A(new_n21803), .Y(new_n21845));
  and_5  g19497(.A(new_n21802), .B(new_n21801), .Y(new_n21846));
  xor_4  g19498(.A(new_n21846), .B(new_n21845), .Y(new_n21847));
  or_5   g19499(.A(new_n21847), .B(new_n21844), .Y(new_n21848));
  nand_5 g19500(.A(new_n21847), .B(new_n21844), .Y(new_n21849));
  nand_5 g19501(.A(new_n21849), .B(new_n11815), .Y(new_n21850));
  nand_5 g19502(.A(new_n21850), .B(new_n21848), .Y(new_n21851));
  nand_5 g19503(.A(new_n21851), .B(new_n21841), .Y(new_n21852));
  nand_5 g19504(.A(new_n21852), .B(new_n21840), .Y(new_n21853));
  nand_5 g19505(.A(new_n21853), .B(new_n21837), .Y(new_n21854));
  nand_5 g19506(.A(new_n21854), .B(new_n21836), .Y(new_n21855));
  nand_5 g19507(.A(new_n21855), .B(new_n21833), .Y(new_n21856));
  nand_5 g19508(.A(new_n21856), .B(new_n21832_1), .Y(new_n21857));
  nand_5 g19509(.A(new_n21857), .B(new_n21829), .Y(new_n21858));
  nand_5 g19510(.A(new_n21858), .B(new_n21828), .Y(new_n21859));
  nand_5 g19511(.A(new_n21859), .B(new_n21825), .Y(new_n21860));
  nand_5 g19512(.A(new_n21860), .B(new_n21824), .Y(new_n21861));
  nand_5 g19513(.A(new_n21861), .B(new_n21821), .Y(new_n21862));
  nand_5 g19514(.A(new_n21862), .B(new_n21820_1), .Y(new_n21863));
  nand_5 g19515(.A(new_n21817), .B(new_n21815), .Y(new_n21864));
  nand_5 g19516(.A(new_n21864), .B(new_n21816), .Y(new_n21865));
  nand_5 g19517(.A(new_n3296), .B(n6814), .Y(new_n21866));
  nand_5 g19518(.A(n27089), .B(new_n3286), .Y(new_n21867));
  nand_5 g19519(.A(new_n21867), .B(new_n21866), .Y(new_n21868));
  xnor_4 g19520(.A(new_n21868), .B(new_n21865), .Y(new_n21869));
  nand_5 g19521(.A(new_n21869), .B(new_n11758), .Y(new_n21870));
  not_8  g19522(.A(new_n21870), .Y(new_n21871));
  nor_5  g19523(.A(new_n21869), .B(new_n11758), .Y(new_n21872));
  nor_5  g19524(.A(new_n21872), .B(new_n21871), .Y(new_n21873));
  xor_4  g19525(.A(new_n21873), .B(new_n21863), .Y(n5911));
  xor_4  g19526(.A(new_n13713), .B(new_n13712), .Y(n5936));
  nand_5 g19527(.A(new_n11560), .B(new_n11558), .Y(new_n21876));
  xor_4  g19528(.A(new_n21876), .B(new_n11611), .Y(n5943));
  nand_5 g19529(.A(new_n16207), .B(new_n16206_1), .Y(new_n21878));
  xor_4  g19530(.A(new_n21878), .B(new_n16247_1), .Y(n5964));
  nand_5 g19531(.A(new_n18215), .B(n8255), .Y(new_n21880));
  not_8  g19532(.A(new_n5700_1), .Y(new_n21881));
  nand_5 g19533(.A(new_n21881), .B(new_n5684), .Y(new_n21882));
  nand_5 g19534(.A(new_n21882), .B(new_n5690), .Y(new_n21883));
  nand_5 g19535(.A(new_n5700_1), .B(n23146), .Y(new_n21884));
  nand_5 g19536(.A(new_n21884), .B(new_n21883), .Y(new_n21885));
  nand_5 g19537(.A(new_n5732_1), .B(new_n5724), .Y(new_n21886));
  nand_5 g19538(.A(new_n21886), .B(new_n21885), .Y(new_n21887));
  nand_5 g19539(.A(new_n5733), .B(n11184), .Y(new_n21888));
  nand_5 g19540(.A(new_n21888), .B(new_n21887), .Y(new_n21889));
  nand_5 g19541(.A(new_n18217), .B(new_n18213), .Y(new_n21890));
  nand_5 g19542(.A(new_n21890), .B(new_n21889), .Y(new_n21891));
  nand_5 g19543(.A(new_n21891), .B(new_n21880), .Y(new_n21892));
  nand_5 g19544(.A(new_n21892), .B(new_n18288_1), .Y(new_n21893));
  nand_5 g19545(.A(new_n21893), .B(new_n18289), .Y(new_n21894));
  nand_5 g19546(.A(new_n21894), .B(new_n18281), .Y(new_n21895));
  nand_5 g19547(.A(new_n21895), .B(new_n18282), .Y(new_n21896));
  nand_5 g19548(.A(new_n21896), .B(new_n18272), .Y(new_n21897));
  nand_5 g19549(.A(new_n21897), .B(new_n18273), .Y(new_n21898_1));
  xor_4  g19550(.A(new_n21898_1), .B(new_n18265), .Y(new_n21899));
  or_5   g19551(.A(new_n21899), .B(new_n3469), .Y(new_n21900));
  nand_5 g19552(.A(new_n21899), .B(new_n3469), .Y(new_n21901));
  xor_4  g19553(.A(new_n21896), .B(new_n18274_1), .Y(new_n21902));
  nand_5 g19554(.A(new_n21902), .B(new_n3479), .Y(new_n21903));
  nor_5  g19555(.A(new_n21902), .B(new_n3479), .Y(new_n21904));
  not_8  g19556(.A(new_n21904), .Y(new_n21905_1));
  xor_4  g19557(.A(new_n21894), .B(new_n18283), .Y(new_n21906));
  nand_5 g19558(.A(new_n21906), .B(new_n3486), .Y(new_n21907));
  nor_5  g19559(.A(new_n21906), .B(new_n3486), .Y(new_n21908));
  not_8  g19560(.A(new_n21908), .Y(new_n21909));
  xor_4  g19561(.A(new_n21892), .B(new_n18290_1), .Y(new_n21910));
  nand_5 g19562(.A(new_n21910), .B(new_n3493), .Y(new_n21911));
  not_8  g19563(.A(new_n21911), .Y(new_n21912));
  nor_5  g19564(.A(new_n21910), .B(new_n3493), .Y(new_n21913));
  xor_4  g19565(.A(new_n21889), .B(new_n18294), .Y(new_n21914));
  nand_5 g19566(.A(new_n21914), .B(new_n3497), .Y(new_n21915_1));
  or_5   g19567(.A(new_n21914), .B(new_n3497), .Y(new_n21916));
  xor_4  g19568(.A(new_n21885), .B(new_n5736), .Y(new_n21917));
  nand_5 g19569(.A(new_n21917), .B(new_n3503), .Y(new_n21918));
  or_5   g19570(.A(new_n21917), .B(new_n3503), .Y(new_n21919));
  xor_4  g19571(.A(new_n21881), .B(new_n5693), .Y(new_n21920));
  or_5   g19572(.A(new_n21920), .B(new_n3517), .Y(new_n21921));
  nand_5 g19573(.A(new_n21920), .B(new_n3517), .Y(new_n21922));
  nand_5 g19574(.A(new_n21922), .B(new_n14931_1), .Y(new_n21923));
  nand_5 g19575(.A(new_n21923), .B(new_n21921), .Y(new_n21924));
  nand_5 g19576(.A(new_n21924), .B(new_n21919), .Y(new_n21925));
  nand_5 g19577(.A(new_n21925), .B(new_n21918), .Y(new_n21926));
  nand_5 g19578(.A(new_n21926), .B(new_n21916), .Y(new_n21927));
  nand_5 g19579(.A(new_n21927), .B(new_n21915_1), .Y(new_n21928));
  nor_5  g19580(.A(new_n21928), .B(new_n21913), .Y(new_n21929));
  nor_5  g19581(.A(new_n21929), .B(new_n21912), .Y(new_n21930));
  not_8  g19582(.A(new_n21930), .Y(new_n21931));
  nand_5 g19583(.A(new_n21931), .B(new_n21909), .Y(new_n21932));
  nand_5 g19584(.A(new_n21932), .B(new_n21907), .Y(new_n21933));
  nand_5 g19585(.A(new_n21933), .B(new_n21905_1), .Y(new_n21934_1));
  nand_5 g19586(.A(new_n21934_1), .B(new_n21903), .Y(new_n21935));
  nand_5 g19587(.A(new_n21935), .B(new_n21901), .Y(new_n21936));
  nand_5 g19588(.A(new_n21936), .B(new_n21900), .Y(new_n21937));
  nor_5  g19589(.A(new_n21898_1), .B(new_n18209), .Y(new_n21938));
  nor_5  g19590(.A(new_n21938), .B(new_n18207), .Y(new_n21939));
  and_5  g19591(.A(new_n21898_1), .B(new_n18209), .Y(new_n21940));
  nor_5  g19592(.A(new_n21940), .B(new_n21939), .Y(new_n21941));
  xor_4  g19593(.A(new_n21941), .B(new_n18258), .Y(new_n21942));
  nand_5 g19594(.A(new_n21942), .B(new_n3465), .Y(new_n21943_1));
  nor_5  g19595(.A(new_n21942), .B(new_n3465), .Y(new_n21944));
  not_8  g19596(.A(new_n21944), .Y(new_n21945));
  nand_5 g19597(.A(new_n21945), .B(new_n21943_1), .Y(new_n21946));
  xor_4  g19598(.A(new_n21946), .B(new_n21937), .Y(n5980));
  nand_5 g19599(.A(new_n12916), .B(new_n12917_1), .Y(new_n21948));
  xnor_4 g19600(.A(new_n21948), .B(new_n12945), .Y(n6012));
  nand_5 g19601(.A(new_n11646), .B(n16544), .Y(new_n21950));
  nand_5 g19602(.A(new_n11647_1), .B(new_n10316), .Y(new_n21951));
  nand_5 g19603(.A(new_n11651), .B(n6814), .Y(new_n21952));
  nand_5 g19604(.A(new_n11652), .B(new_n3286), .Y(new_n21953));
  nand_5 g19605(.A(new_n11656), .B(n19701), .Y(new_n21954));
  nand_5 g19606(.A(new_n11657), .B(new_n3186), .Y(new_n21955));
  nand_5 g19607(.A(new_n10829), .B(new_n10819), .Y(new_n21956));
  nand_5 g19608(.A(new_n21956), .B(new_n10827), .Y(new_n21957_1));
  nand_5 g19609(.A(new_n21957_1), .B(new_n21955), .Y(new_n21958));
  nand_5 g19610(.A(new_n21958), .B(new_n21954), .Y(new_n21959));
  nand_5 g19611(.A(new_n21959), .B(new_n21953), .Y(new_n21960_1));
  nand_5 g19612(.A(new_n21960_1), .B(new_n21952), .Y(new_n21961));
  nand_5 g19613(.A(new_n21961), .B(new_n21951), .Y(new_n21962));
  nand_5 g19614(.A(new_n21962), .B(new_n21950), .Y(new_n21963));
  xor_4  g19615(.A(new_n21963), .B(new_n11638), .Y(new_n21964));
  nand_5 g19616(.A(new_n16065), .B(new_n6795), .Y(new_n21965));
  nand_5 g19617(.A(new_n16064), .B(n3582), .Y(new_n21966));
  nand_5 g19618(.A(new_n16070), .B(new_n6799), .Y(new_n21967));
  nand_5 g19619(.A(new_n16069), .B(n2145), .Y(new_n21968));
  nand_5 g19620(.A(new_n16075), .B(new_n6803), .Y(new_n21969));
  nand_5 g19621(.A(new_n16074), .B(n5031), .Y(new_n21970));
  nand_5 g19622(.A(new_n10843), .B(new_n10833), .Y(new_n21971));
  nand_5 g19623(.A(new_n21971), .B(new_n10841), .Y(new_n21972));
  nand_5 g19624(.A(new_n21972), .B(new_n21970), .Y(new_n21973));
  nand_5 g19625(.A(new_n21973), .B(new_n21969), .Y(new_n21974));
  nand_5 g19626(.A(new_n21974), .B(new_n21968), .Y(new_n21975));
  nand_5 g19627(.A(new_n21975), .B(new_n21967), .Y(new_n21976_1));
  nand_5 g19628(.A(new_n21976_1), .B(new_n21966), .Y(new_n21977));
  nand_5 g19629(.A(new_n21977), .B(new_n21965), .Y(new_n21978));
  nor_5  g19630(.A(new_n21978), .B(new_n16062_1), .Y(new_n21979));
  not_8  g19631(.A(new_n21979), .Y(new_n21980));
  nand_5 g19632(.A(new_n21978), .B(new_n16062_1), .Y(new_n21981_1));
  and_5  g19633(.A(new_n21981_1), .B(new_n21980), .Y(new_n21982));
  not_8  g19634(.A(new_n21982), .Y(new_n21983));
  or_5   g19635(.A(new_n21983), .B(new_n21964), .Y(new_n21984));
  nand_5 g19636(.A(new_n21983), .B(new_n21964), .Y(new_n21985));
  nand_5 g19637(.A(new_n21950), .B(new_n21951), .Y(new_n21986_1));
  xor_4  g19638(.A(new_n21986_1), .B(new_n21961), .Y(new_n21987));
  nand_5 g19639(.A(new_n21965), .B(new_n21966), .Y(new_n21988));
  xor_4  g19640(.A(new_n21988), .B(new_n21976_1), .Y(new_n21989));
  nand_5 g19641(.A(new_n21989), .B(new_n21987), .Y(new_n21990));
  nand_5 g19642(.A(new_n21952), .B(new_n21953), .Y(new_n21991));
  xor_4  g19643(.A(new_n21991), .B(new_n21959), .Y(new_n21992));
  nand_5 g19644(.A(new_n21967), .B(new_n21968), .Y(new_n21993_1));
  xor_4  g19645(.A(new_n21993_1), .B(new_n21974), .Y(new_n21994));
  nand_5 g19646(.A(new_n21994), .B(new_n21992), .Y(new_n21995));
  or_5   g19647(.A(new_n21994), .B(new_n21992), .Y(new_n21996));
  nand_5 g19648(.A(new_n21954), .B(new_n21955), .Y(new_n21997_1));
  xor_4  g19649(.A(new_n21997_1), .B(new_n21957_1), .Y(new_n21998));
  nand_5 g19650(.A(new_n21969), .B(new_n21970), .Y(new_n21999));
  xor_4  g19651(.A(new_n21999), .B(new_n21972), .Y(new_n22000));
  nand_5 g19652(.A(new_n22000), .B(new_n21998), .Y(new_n22001));
  or_5   g19653(.A(new_n22000), .B(new_n21998), .Y(new_n22002));
  nand_5 g19654(.A(new_n10849), .B(new_n10817_1), .Y(new_n22003));
  nand_5 g19655(.A(new_n22003), .B(new_n10847), .Y(new_n22004));
  not_8  g19656(.A(new_n22004), .Y(new_n22005));
  nand_5 g19657(.A(new_n22005), .B(new_n22002), .Y(new_n22006));
  nand_5 g19658(.A(new_n22006), .B(new_n22001), .Y(new_n22007));
  nand_5 g19659(.A(new_n22007), .B(new_n21996), .Y(new_n22008));
  nand_5 g19660(.A(new_n22008), .B(new_n21995), .Y(new_n22009));
  or_5   g19661(.A(new_n21989), .B(new_n21987), .Y(new_n22010));
  nand_5 g19662(.A(new_n22010), .B(new_n22009), .Y(new_n22011));
  nand_5 g19663(.A(new_n22011), .B(new_n21990), .Y(new_n22012));
  nand_5 g19664(.A(new_n22012), .B(new_n21985), .Y(new_n22013));
  nand_5 g19665(.A(new_n22013), .B(new_n21984), .Y(new_n22014));
  nand_5 g19666(.A(new_n21963), .B(new_n11638), .Y(new_n22015));
  or_5   g19667(.A(new_n21979), .B(new_n22015), .Y(new_n22016_1));
  nand_5 g19668(.A(new_n21979), .B(new_n22015), .Y(new_n22017));
  nand_5 g19669(.A(new_n22017), .B(new_n22016_1), .Y(new_n22018));
  xor_4  g19670(.A(new_n22018), .B(new_n22014), .Y(n6022));
  nand_5 g19671(.A(new_n21585), .B(new_n21586), .Y(new_n22020));
  xor_4  g19672(.A(new_n22020), .B(new_n21605), .Y(n6031));
  nand_5 g19673(.A(new_n19064), .B(new_n8294), .Y(new_n22022));
  xor_4  g19674(.A(new_n22022), .B(n17458), .Y(new_n22023));
  xor_4  g19675(.A(new_n22023), .B(n12507), .Y(new_n22024));
  nand_5 g19676(.A(new_n19070), .B(new_n19066), .Y(new_n22025));
  nand_5 g19677(.A(new_n22025), .B(new_n19067), .Y(new_n22026));
  xor_4  g19678(.A(new_n22026), .B(new_n22024), .Y(new_n22027_1));
  not_8  g19679(.A(new_n22027_1), .Y(new_n22028));
  nand_5 g19680(.A(new_n22028), .B(n12702), .Y(new_n22029));
  nand_5 g19681(.A(new_n22027_1), .B(new_n9271), .Y(new_n22030));
  nand_5 g19682(.A(new_n22030), .B(new_n22029), .Y(new_n22031));
  nand_5 g19683(.A(new_n19074), .B(new_n19063), .Y(new_n22032));
  nand_5 g19684(.A(new_n22032), .B(new_n19073), .Y(new_n22033));
  xor_4  g19685(.A(new_n22033), .B(new_n22031), .Y(new_n22034));
  nand_5 g19686(.A(new_n22034), .B(new_n9354), .Y(new_n22035));
  not_8  g19687(.A(new_n22035), .Y(new_n22036));
  nor_5  g19688(.A(new_n22034), .B(new_n9354), .Y(new_n22037));
  or_5   g19689(.A(new_n22037), .B(new_n22036), .Y(new_n22038));
  nor_5  g19690(.A(new_n19080), .B(new_n19061), .Y(new_n22039));
  nor_5  g19691(.A(new_n22039), .B(new_n19079), .Y(new_n22040));
  xor_4  g19692(.A(new_n22040), .B(new_n22038), .Y(n6044));
  nor_5  g19693(.A(new_n10466), .B(n4306), .Y(new_n22042));
  not_8  g19694(.A(new_n22042), .Y(new_n22043_1));
  nand_5 g19695(.A(new_n20536), .B(new_n22043_1), .Y(new_n22044));
  nand_5 g19696(.A(new_n10584), .B(new_n10513), .Y(new_n22045));
  nand_5 g19697(.A(new_n22045), .B(new_n10512), .Y(new_n22046));
  nor_5  g19698(.A(new_n22046), .B(new_n22044), .Y(new_n22047));
  and_5  g19699(.A(new_n22047), .B(new_n4927), .Y(new_n22048));
  or_5   g19700(.A(new_n22046), .B(new_n22042), .Y(new_n22049));
  xor_4  g19701(.A(new_n22049), .B(new_n20536), .Y(new_n22050_1));
  or_5   g19702(.A(new_n22050_1), .B(new_n5044), .Y(new_n22051));
  nand_5 g19703(.A(new_n10647_1), .B(new_n10587), .Y(new_n22052));
  nand_5 g19704(.A(new_n22052), .B(new_n10588_1), .Y(new_n22053));
  and_5  g19705(.A(new_n22053), .B(new_n22051), .Y(new_n22054));
  nor_5  g19706(.A(new_n22054), .B(new_n22048), .Y(new_n22055));
  nor_5  g19707(.A(new_n22047), .B(new_n4927), .Y(new_n22056));
  nand_5 g19708(.A(new_n22050_1), .B(new_n5044), .Y(new_n22057));
  not_8  g19709(.A(new_n22057), .Y(new_n22058));
  nor_5  g19710(.A(new_n22058), .B(new_n22054), .Y(new_n22059));
  nor_5  g19711(.A(new_n22059), .B(new_n22056), .Y(new_n22060));
  nor_5  g19712(.A(new_n22060), .B(new_n22055), .Y(n6046));
  nand_5 g19713(.A(new_n21743), .B(new_n21733), .Y(new_n22062));
  nand_5 g19714(.A(new_n22062), .B(new_n21742), .Y(new_n22063_1));
  not_8  g19715(.A(new_n21738), .Y(new_n22064));
  not_8  g19716(.A(new_n21739), .Y(new_n22065));
  nor_5  g19717(.A(new_n22065), .B(new_n21737), .Y(new_n22066));
  nor_5  g19718(.A(new_n22066), .B(new_n22064), .Y(new_n22067));
  nand_5 g19719(.A(new_n9834), .B(new_n8153), .Y(new_n22068_1));
  nand_5 g19720(.A(n25119), .B(n21934), .Y(new_n22069));
  nand_5 g19721(.A(new_n22069), .B(new_n22068_1), .Y(new_n22070));
  xor_4  g19722(.A(new_n22070), .B(new_n22067), .Y(new_n22071));
  or_5   g19723(.A(new_n22071), .B(new_n2576), .Y(new_n22072_1));
  nand_5 g19724(.A(new_n22071), .B(new_n2576), .Y(new_n22073));
  nand_5 g19725(.A(new_n22073), .B(new_n22072_1), .Y(new_n22074));
  xor_4  g19726(.A(new_n22074), .B(new_n22063_1), .Y(new_n22075));
  not_8  g19727(.A(new_n22075), .Y(new_n22076_1));
  nand_5 g19728(.A(new_n21751), .B(new_n21748), .Y(new_n22077));
  nand_5 g19729(.A(new_n22077), .B(new_n21750_1), .Y(new_n22078));
  not_8  g19730(.A(new_n22078), .Y(new_n22079));
  nand_5 g19731(.A(new_n3109), .B(n20700), .Y(new_n22080));
  nand_5 g19732(.A(n26510), .B(new_n3067_1), .Y(new_n22081));
  nand_5 g19733(.A(new_n22081), .B(new_n22080), .Y(new_n22082));
  xor_4  g19734(.A(new_n22082), .B(new_n22079), .Y(new_n22083));
  or_5   g19735(.A(new_n22083), .B(new_n22076_1), .Y(new_n22084));
  nand_5 g19736(.A(new_n22083), .B(new_n22076_1), .Y(new_n22085));
  nor_5  g19737(.A(new_n21757), .B(new_n21731), .Y(new_n22086));
  nor_5  g19738(.A(new_n22086), .B(new_n21755), .Y(new_n22087));
  not_8  g19739(.A(new_n22087), .Y(new_n22088));
  nand_5 g19740(.A(new_n22088), .B(new_n22085), .Y(new_n22089));
  nand_5 g19741(.A(new_n22089), .B(new_n22084), .Y(new_n22090_1));
  nand_5 g19742(.A(new_n22073), .B(new_n22063_1), .Y(new_n22091));
  nand_5 g19743(.A(new_n22091), .B(new_n22072_1), .Y(new_n22092));
  not_8  g19744(.A(new_n22068_1), .Y(new_n22093));
  not_8  g19745(.A(new_n22069), .Y(new_n22094));
  nor_5  g19746(.A(new_n22094), .B(new_n22067), .Y(new_n22095));
  nor_5  g19747(.A(new_n22095), .B(new_n22093), .Y(new_n22096));
  nand_5 g19748(.A(new_n18133), .B(new_n8150), .Y(new_n22097));
  nand_5 g19749(.A(n21997), .B(n18483), .Y(new_n22098));
  nand_5 g19750(.A(new_n22098), .B(new_n22097), .Y(new_n22099));
  xor_4  g19751(.A(new_n22099), .B(new_n22096), .Y(new_n22100));
  or_5   g19752(.A(new_n22100), .B(new_n8628), .Y(new_n22101));
  nand_5 g19753(.A(new_n22100), .B(new_n8628), .Y(new_n22102));
  nand_5 g19754(.A(new_n22102), .B(new_n22101), .Y(new_n22103));
  xor_4  g19755(.A(new_n22103), .B(new_n22092), .Y(new_n22104));
  not_8  g19756(.A(new_n22104), .Y(new_n22105));
  nand_5 g19757(.A(new_n22081), .B(new_n22078), .Y(new_n22106));
  nand_5 g19758(.A(new_n22106), .B(new_n22080), .Y(new_n22107_1));
  not_8  g19759(.A(new_n22107_1), .Y(new_n22108));
  nand_5 g19760(.A(new_n3195), .B(n7437), .Y(new_n22109));
  nand_5 g19761(.A(n17077), .B(new_n3185), .Y(new_n22110));
  nand_5 g19762(.A(new_n22110), .B(new_n22109), .Y(new_n22111));
  xor_4  g19763(.A(new_n22111), .B(new_n22108), .Y(new_n22112));
  or_5   g19764(.A(new_n22112), .B(new_n22105), .Y(new_n22113_1));
  nand_5 g19765(.A(new_n22112), .B(new_n22105), .Y(new_n22114));
  nand_5 g19766(.A(new_n22114), .B(new_n22113_1), .Y(new_n22115));
  xor_4  g19767(.A(new_n22115), .B(new_n22090_1), .Y(n6084));
  nand_5 g19768(.A(new_n21849), .B(new_n21848), .Y(new_n22117));
  xnor_4 g19769(.A(new_n22117), .B(new_n11815), .Y(n6160));
  nand_5 g19770(.A(new_n21837), .B(new_n21836), .Y(new_n22119));
  xnor_4 g19771(.A(new_n22119), .B(new_n21853), .Y(n6171));
  nand_5 g19772(.A(new_n20629_1), .B(new_n20627), .Y(new_n22121));
  nand_5 g19773(.A(new_n22121), .B(new_n20628), .Y(new_n22122));
  nand_5 g19774(.A(new_n11350), .B(n16812), .Y(new_n22123));
  nand_5 g19775(.A(n25923), .B(new_n9169), .Y(new_n22124_1));
  nand_5 g19776(.A(new_n22124_1), .B(new_n22123), .Y(new_n22125));
  xnor_4 g19777(.A(new_n22125), .B(new_n22122), .Y(new_n22126_1));
  nand_5 g19778(.A(new_n22126_1), .B(new_n17365), .Y(new_n22127));
  or_5   g19779(.A(new_n22126_1), .B(new_n17365), .Y(new_n22128));
  nand_5 g19780(.A(new_n20633), .B(new_n20625), .Y(new_n22129));
  nand_5 g19781(.A(new_n22129), .B(new_n20632), .Y(new_n22130_1));
  nand_5 g19782(.A(new_n22130_1), .B(new_n22128), .Y(new_n22131));
  nand_5 g19783(.A(new_n22131), .B(new_n22127), .Y(new_n22132));
  nand_5 g19784(.A(new_n22124_1), .B(new_n22122), .Y(new_n22133));
  nand_5 g19785(.A(new_n22133), .B(new_n22123), .Y(new_n22134));
  nand_5 g19786(.A(new_n11345), .B(n7841), .Y(new_n22135));
  nand_5 g19787(.A(n22918), .B(new_n9163), .Y(new_n22136));
  nand_5 g19788(.A(new_n22136), .B(new_n22135), .Y(new_n22137));
  xor_4  g19789(.A(new_n22137), .B(new_n22134), .Y(new_n22138));
  or_5   g19790(.A(new_n22138), .B(new_n17423), .Y(new_n22139));
  nand_5 g19791(.A(new_n22138), .B(new_n17423), .Y(new_n22140));
  nand_5 g19792(.A(new_n22140), .B(new_n22139), .Y(new_n22141));
  xor_4  g19793(.A(new_n22141), .B(new_n22132), .Y(new_n22142));
  nand_5 g19794(.A(new_n22142), .B(new_n17434), .Y(new_n22143));
  or_5   g19795(.A(new_n22142), .B(new_n17434), .Y(new_n22144_1));
  nand_5 g19796(.A(new_n22128), .B(new_n22127), .Y(new_n22145));
  xor_4  g19797(.A(new_n22145), .B(new_n22130_1), .Y(new_n22146));
  not_8  g19798(.A(new_n22146), .Y(new_n22147));
  nand_5 g19799(.A(new_n22147), .B(new_n17358), .Y(new_n22148));
  nand_5 g19800(.A(new_n22146), .B(new_n17360), .Y(new_n22149));
  nand_5 g19801(.A(new_n20638), .B(new_n20623_1), .Y(new_n22150_1));
  nand_5 g19802(.A(new_n22150_1), .B(new_n20637), .Y(new_n22151));
  nand_5 g19803(.A(new_n22151), .B(new_n22149), .Y(new_n22152));
  nand_5 g19804(.A(new_n22152), .B(new_n22148), .Y(new_n22153));
  not_8  g19805(.A(new_n22153), .Y(new_n22154));
  nand_5 g19806(.A(new_n22154), .B(new_n22144_1), .Y(new_n22155));
  nand_5 g19807(.A(new_n22155), .B(new_n22143), .Y(new_n22156));
  nand_5 g19808(.A(new_n22140), .B(new_n22132), .Y(new_n22157_1));
  nand_5 g19809(.A(new_n22157_1), .B(new_n22139), .Y(new_n22158));
  nand_5 g19810(.A(new_n22136), .B(new_n22134), .Y(new_n22159));
  nand_5 g19811(.A(new_n22159), .B(new_n22135), .Y(new_n22160));
  nand_5 g19812(.A(n26264), .B(new_n11340), .Y(new_n22161));
  nand_5 g19813(.A(new_n9157), .B(n21905), .Y(new_n22162));
  nand_5 g19814(.A(new_n22162), .B(new_n22161), .Y(new_n22163));
  xnor_4 g19815(.A(new_n22163), .B(new_n22160), .Y(new_n22164));
  nand_5 g19816(.A(new_n22164), .B(new_n17670), .Y(new_n22165));
  or_5   g19817(.A(new_n22164), .B(new_n17670), .Y(new_n22166));
  nand_5 g19818(.A(new_n22166), .B(new_n22165), .Y(new_n22167));
  xor_4  g19819(.A(new_n22167), .B(new_n22158), .Y(new_n22168));
  nand_5 g19820(.A(new_n17430), .B(new_n11460), .Y(new_n22169));
  nand_5 g19821(.A(new_n22169), .B(new_n11459), .Y(new_n22170));
  not_8  g19822(.A(new_n22170), .Y(new_n22171));
  xor_4  g19823(.A(new_n22171), .B(new_n11455_1), .Y(new_n22172));
  not_8  g19824(.A(new_n22172), .Y(new_n22173_1));
  nand_5 g19825(.A(new_n22173_1), .B(new_n22168), .Y(new_n22174));
  or_5   g19826(.A(new_n22173_1), .B(new_n22168), .Y(new_n22175));
  nand_5 g19827(.A(new_n22175), .B(new_n22174), .Y(new_n22176));
  xor_4  g19828(.A(new_n22176), .B(new_n22156), .Y(n6183));
  nand_5 g19829(.A(n3164), .B(new_n10456), .Y(new_n22178));
  nand_5 g19830(.A(new_n10485), .B(n2547), .Y(new_n22179));
  nand_5 g19831(.A(new_n16042), .B(new_n16040), .Y(new_n22180));
  nand_5 g19832(.A(new_n22180), .B(new_n16041), .Y(new_n22181));
  nand_5 g19833(.A(new_n22181), .B(new_n22179), .Y(new_n22182));
  nand_5 g19834(.A(new_n22182), .B(new_n22178), .Y(new_n22183));
  nand_5 g19835(.A(n11356), .B(new_n12366), .Y(new_n22184));
  nand_5 g19836(.A(new_n10482), .B(n2999), .Y(new_n22185));
  nand_5 g19837(.A(new_n22185), .B(new_n22184), .Y(new_n22186));
  xor_4  g19838(.A(new_n22186), .B(new_n22183), .Y(new_n22187));
  nand_5 g19839(.A(new_n22187), .B(new_n10394), .Y(new_n22188));
  or_5   g19840(.A(new_n22187), .B(new_n10394), .Y(new_n22189));
  nand_5 g19841(.A(new_n22179), .B(new_n22178), .Y(new_n22190));
  xor_4  g19842(.A(new_n22190), .B(new_n22181), .Y(new_n22191));
  nand_5 g19843(.A(new_n22191), .B(new_n10401), .Y(new_n22192));
  or_5   g19844(.A(new_n22191), .B(new_n10401), .Y(new_n22193));
  nand_5 g19845(.A(new_n16045), .B(new_n16038), .Y(new_n22194));
  nand_5 g19846(.A(new_n22194), .B(new_n16046), .Y(new_n22195));
  nand_5 g19847(.A(new_n22195), .B(new_n22193), .Y(new_n22196));
  nand_5 g19848(.A(new_n22196), .B(new_n22192), .Y(new_n22197));
  nand_5 g19849(.A(new_n22197), .B(new_n22189), .Y(new_n22198_1));
  nand_5 g19850(.A(new_n22198_1), .B(new_n22188), .Y(new_n22199));
  nand_5 g19851(.A(new_n22185), .B(new_n22183), .Y(new_n22200));
  nand_5 g19852(.A(new_n22200), .B(new_n22184), .Y(new_n22201_1));
  nand_5 g19853(.A(new_n10455), .B(n14345), .Y(new_n22202));
  nand_5 g19854(.A(n14702), .B(new_n10479), .Y(new_n22203));
  nand_5 g19855(.A(new_n22203), .B(new_n22202), .Y(new_n22204));
  xnor_4 g19856(.A(new_n22204), .B(new_n22201_1), .Y(new_n22205));
  or_5   g19857(.A(new_n22205), .B(new_n10386), .Y(new_n22206));
  nand_5 g19858(.A(new_n22205), .B(new_n10386), .Y(new_n22207));
  nand_5 g19859(.A(new_n22207), .B(new_n22206), .Y(new_n22208));
  xor_4  g19860(.A(new_n22208), .B(new_n22199), .Y(n6189));
  xor_4  g19861(.A(n9380), .B(n8656), .Y(new_n22210));
  nand_5 g19862(.A(new_n22210), .B(new_n17155), .Y(new_n22211));
  nand_5 g19863(.A(new_n4545), .B(n8656), .Y(new_n22212));
  not_8  g19864(.A(new_n22212), .Y(new_n22213_1));
  nand_5 g19865(.A(new_n7347), .B(n11192), .Y(new_n22214));
  nand_5 g19866(.A(n21095), .B(new_n4561), .Y(new_n22215));
  and_5  g19867(.A(new_n22215), .B(new_n22214), .Y(new_n22216));
  xor_4  g19868(.A(new_n22216), .B(new_n22213_1), .Y(new_n22217));
  or_5   g19869(.A(new_n22217), .B(new_n22211), .Y(new_n22218));
  nand_5 g19870(.A(new_n22217), .B(new_n22211), .Y(new_n22219));
  nand_5 g19871(.A(new_n22219), .B(new_n20615), .Y(new_n22220));
  nand_5 g19872(.A(new_n22220), .B(new_n22218), .Y(new_n22221));
  nand_5 g19873(.A(new_n22215), .B(new_n22212), .Y(new_n22222));
  nand_5 g19874(.A(new_n22222), .B(new_n22214), .Y(new_n22223));
  nand_5 g19875(.A(n20036), .B(new_n7341), .Y(new_n22224));
  nand_5 g19876(.A(new_n4606), .B(n15167), .Y(new_n22225));
  nand_5 g19877(.A(new_n22225), .B(new_n22224), .Y(new_n22226));
  xnor_4 g19878(.A(new_n22226), .B(new_n22223), .Y(new_n22227));
  nand_5 g19879(.A(new_n22227), .B(new_n20608), .Y(new_n22228));
  or_5   g19880(.A(new_n22227), .B(new_n20608), .Y(new_n22229));
  nand_5 g19881(.A(new_n22229), .B(new_n22228), .Y(new_n22230));
  xnor_4 g19882(.A(new_n22230), .B(new_n22221), .Y(n6223));
  nand_5 g19883(.A(new_n16028), .B(new_n16027), .Y(new_n22232));
  xor_4  g19884(.A(new_n22232), .B(new_n16036), .Y(n6233));
  nand_5 g19885(.A(new_n21299), .B(new_n21300), .Y(new_n22234));
  xor_4  g19886(.A(new_n22234), .B(new_n21302_1), .Y(n6245));
  nand_5 g19887(.A(new_n11803), .B(new_n11804), .Y(new_n22236));
  xnor_4 g19888(.A(new_n22236), .B(new_n11817), .Y(n6248));
  nand_5 g19889(.A(new_n4813), .B(n16544), .Y(new_n22238));
  nand_5 g19890(.A(n21839), .B(new_n10316), .Y(new_n22239));
  nand_5 g19891(.A(new_n22239), .B(new_n22238), .Y(new_n22240));
  nand_5 g19892(.A(new_n21867), .B(new_n21865), .Y(new_n22241));
  nand_5 g19893(.A(new_n22241), .B(new_n21866), .Y(new_n22242));
  xnor_4 g19894(.A(new_n22242), .B(new_n22240), .Y(new_n22243));
  nand_5 g19895(.A(new_n22243), .B(new_n11751), .Y(new_n22244));
  not_8  g19896(.A(new_n22244), .Y(new_n22245));
  nor_5  g19897(.A(new_n22243), .B(new_n11751), .Y(new_n22246));
  or_5   g19898(.A(new_n22246), .B(new_n22245), .Y(new_n22247));
  not_8  g19899(.A(new_n21863), .Y(new_n22248));
  nor_5  g19900(.A(new_n21872), .B(new_n22248), .Y(new_n22249));
  nor_5  g19901(.A(new_n22249), .B(new_n21871), .Y(new_n22250));
  xor_4  g19902(.A(new_n22250), .B(new_n22247), .Y(n6256));
  nand_5 g19903(.A(new_n16972), .B(new_n16974), .Y(new_n22252));
  xor_4  g19904(.A(new_n22252), .B(new_n16991), .Y(n6271));
  nand_5 g19905(.A(new_n22170), .B(new_n11454), .Y(new_n22254));
  nand_5 g19906(.A(new_n22254), .B(new_n11453), .Y(new_n22255));
  nand_5 g19907(.A(new_n9104_1), .B(n13549), .Y(new_n22256));
  nand_5 g19908(.A(new_n22256), .B(new_n22255), .Y(new_n22257));
  nand_5 g19909(.A(n14826), .B(new_n11404), .Y(new_n22258));
  nand_5 g19910(.A(new_n22258), .B(new_n22257), .Y(new_n22259));
  not_8  g19911(.A(new_n22259), .Y(new_n22260));
  nand_5 g19912(.A(new_n11694), .B(n2944), .Y(new_n22261));
  nand_5 g19913(.A(new_n17110), .B(new_n17107), .Y(new_n22262));
  nand_5 g19914(.A(new_n22262), .B(new_n17109), .Y(new_n22263));
  nand_5 g19915(.A(n13951), .B(new_n2781), .Y(new_n22264));
  nand_5 g19916(.A(new_n22264), .B(new_n22263), .Y(new_n22265));
  nand_5 g19917(.A(new_n22265), .B(new_n22261), .Y(new_n22266));
  not_8  g19918(.A(new_n22266), .Y(new_n22267));
  nand_5 g19919(.A(new_n22267), .B(new_n22260), .Y(new_n22268));
  xor_4  g19920(.A(new_n22255), .B(new_n11408), .Y(new_n22269));
  not_8  g19921(.A(new_n22269), .Y(new_n22270_1));
  nand_5 g19922(.A(new_n22264), .B(new_n22261), .Y(new_n22271));
  xor_4  g19923(.A(new_n22271), .B(new_n22263), .Y(new_n22272));
  not_8  g19924(.A(new_n22272), .Y(new_n22273));
  nand_5 g19925(.A(new_n22273), .B(new_n22270_1), .Y(new_n22274_1));
  nand_5 g19926(.A(new_n22272), .B(new_n22269), .Y(new_n22275));
  nand_5 g19927(.A(new_n22172), .B(new_n17112), .Y(new_n22276));
  nand_5 g19928(.A(new_n22173_1), .B(new_n17113), .Y(new_n22277));
  nand_5 g19929(.A(new_n17435), .B(new_n17425), .Y(new_n22278));
  nand_5 g19930(.A(new_n22278), .B(new_n17433), .Y(new_n22279));
  nand_5 g19931(.A(new_n22279), .B(new_n22277), .Y(new_n22280));
  nand_5 g19932(.A(new_n22280), .B(new_n22276), .Y(new_n22281));
  nand_5 g19933(.A(new_n22281), .B(new_n22275), .Y(new_n22282));
  nand_5 g19934(.A(new_n22282), .B(new_n22274_1), .Y(new_n22283_1));
  not_8  g19935(.A(new_n22268), .Y(new_n22284));
  nor_5  g19936(.A(new_n22267), .B(new_n22260), .Y(new_n22285));
  nor_5  g19937(.A(new_n22285), .B(new_n22284), .Y(new_n22286));
  not_8  g19938(.A(new_n22286), .Y(new_n22287));
  or_5   g19939(.A(new_n22287), .B(new_n22283_1), .Y(new_n22288));
  nand_5 g19940(.A(new_n22288), .B(new_n22268), .Y(new_n22289));
  nand_5 g19941(.A(n8827), .B(new_n19998), .Y(new_n22290_1));
  nand_5 g19942(.A(new_n12403), .B(n1881), .Y(new_n22291));
  nand_5 g19943(.A(new_n21616), .B(new_n21613), .Y(new_n22292));
  nand_5 g19944(.A(new_n22292), .B(new_n21615_1), .Y(new_n22293));
  nand_5 g19945(.A(new_n22293), .B(new_n22291), .Y(new_n22294));
  nand_5 g19946(.A(new_n22294), .B(new_n22290_1), .Y(new_n22295));
  xor_4  g19947(.A(new_n22295), .B(new_n22289), .Y(new_n22296));
  nand_5 g19948(.A(new_n22287), .B(new_n22283_1), .Y(new_n22297));
  and_5  g19949(.A(new_n22297), .B(new_n22288), .Y(new_n22298));
  nand_5 g19950(.A(new_n22298), .B(new_n22295), .Y(new_n22299));
  not_8  g19951(.A(new_n22295), .Y(new_n22300));
  not_8  g19952(.A(new_n22298), .Y(new_n22301));
  nand_5 g19953(.A(new_n22301), .B(new_n22300), .Y(new_n22302));
  nand_5 g19954(.A(new_n22274_1), .B(new_n22275), .Y(new_n22303));
  xor_4  g19955(.A(new_n22303), .B(new_n22281), .Y(new_n22304));
  nand_5 g19956(.A(new_n22291), .B(new_n22290_1), .Y(new_n22305));
  xor_4  g19957(.A(new_n22305), .B(new_n22293), .Y(new_n22306));
  nand_5 g19958(.A(new_n22306), .B(new_n22304), .Y(new_n22307));
  not_8  g19959(.A(new_n22304), .Y(new_n22308));
  not_8  g19960(.A(new_n22306), .Y(new_n22309_1));
  nand_5 g19961(.A(new_n22309_1), .B(new_n22308), .Y(new_n22310));
  nand_5 g19962(.A(new_n22276), .B(new_n22277), .Y(new_n22311_1));
  xor_4  g19963(.A(new_n22311_1), .B(new_n22279), .Y(new_n22312));
  nand_5 g19964(.A(new_n22312), .B(new_n21619), .Y(new_n22313));
  not_8  g19965(.A(new_n22312), .Y(new_n22314));
  nand_5 g19966(.A(new_n22314), .B(new_n21618), .Y(new_n22315));
  nand_5 g19967(.A(new_n17641), .B(new_n17630), .Y(new_n22316));
  nand_5 g19968(.A(new_n22316), .B(new_n17640), .Y(new_n22317_1));
  nand_5 g19969(.A(new_n22317_1), .B(new_n22315), .Y(new_n22318));
  nand_5 g19970(.A(new_n22318), .B(new_n22313), .Y(new_n22319));
  nand_5 g19971(.A(new_n22319), .B(new_n22310), .Y(new_n22320));
  nand_5 g19972(.A(new_n22320), .B(new_n22307), .Y(new_n22321));
  nand_5 g19973(.A(new_n22321), .B(new_n22302), .Y(new_n22322));
  nand_5 g19974(.A(new_n22322), .B(new_n22299), .Y(new_n22323));
  xor_4  g19975(.A(new_n22323), .B(new_n22296), .Y(n6276));
  nand_5 g19976(.A(new_n21253), .B(new_n21252), .Y(new_n22325));
  xnor_4 g19977(.A(new_n22325), .B(new_n21261), .Y(n6308));
  nand_5 g19978(.A(new_n19173), .B(new_n19172), .Y(new_n22327));
  xor_4  g19979(.A(new_n22327), .B(new_n19187), .Y(n6311));
  nand_5 g19980(.A(new_n18897), .B(new_n18896), .Y(new_n22329));
  xnor_4 g19981(.A(new_n22329), .B(new_n18911), .Y(n6323));
  nand_5 g19982(.A(new_n6792), .B(new_n6710), .Y(new_n22331));
  nand_5 g19983(.A(new_n22331), .B(new_n6712), .Y(new_n22332_1));
  nand_5 g19984(.A(new_n15343), .B(new_n6659_1), .Y(new_n22333));
  nor_5  g19985(.A(new_n22333), .B(new_n22332_1), .Y(new_n22334));
  not_8  g19986(.A(new_n22332_1), .Y(new_n22335_1));
  nand_5 g19987(.A(new_n15344), .B(new_n6660), .Y(new_n22336));
  nor_5  g19988(.A(new_n22336), .B(new_n22335_1), .Y(new_n22337));
  nor_5  g19989(.A(new_n22337), .B(new_n22334), .Y(new_n22338));
  and_5  g19990(.A(new_n22336), .B(new_n22333), .Y(new_n22339));
  xor_4  g19991(.A(new_n22339), .B(new_n22332_1), .Y(new_n22340));
  or_5   g19992(.A(new_n22340), .B(new_n20370), .Y(new_n22341_1));
  nand_5 g19993(.A(new_n6989), .B(new_n6912), .Y(new_n22342));
  nand_5 g19994(.A(new_n22342), .B(new_n6913), .Y(new_n22343));
  not_8  g19995(.A(new_n22343), .Y(new_n22344));
  nand_5 g19996(.A(new_n22344), .B(new_n22341_1), .Y(new_n22345));
  nand_5 g19997(.A(new_n22340), .B(new_n20370), .Y(new_n22346));
  nand_5 g19998(.A(new_n22346), .B(new_n22345), .Y(new_n22347));
  or_5   g19999(.A(new_n22347), .B(new_n20364), .Y(new_n22348));
  nand_5 g20000(.A(new_n22348), .B(new_n22338), .Y(new_n22349));
  nand_5 g20001(.A(new_n22347), .B(new_n20364), .Y(new_n22350));
  nand_5 g20002(.A(new_n22350), .B(new_n22349), .Y(new_n22351));
  nor_5  g20003(.A(new_n22351), .B(new_n22334), .Y(n6330));
  nand_5 g20004(.A(new_n9783_1), .B(new_n9784), .Y(new_n22353_1));
  xnor_4 g20005(.A(new_n22353_1), .B(new_n9822), .Y(n6339));
  nor_5  g20006(.A(new_n15979_1), .B(new_n15978), .Y(new_n22355));
  xor_4  g20007(.A(new_n22355), .B(new_n16009), .Y(n6354));
  nand_5 g20008(.A(new_n3455), .B(new_n3314), .Y(new_n22357));
  not_8  g20009(.A(new_n22357), .Y(new_n22358_1));
  nand_5 g20010(.A(new_n3464), .B(new_n3317), .Y(new_n22359_1));
  nand_5 g20011(.A(new_n3460_1), .B(n5696), .Y(new_n22360));
  nand_5 g20012(.A(new_n3471), .B(new_n3322), .Y(new_n22361));
  nand_5 g20013(.A(new_n3467), .B(n13367), .Y(new_n22362));
  nand_5 g20014(.A(new_n3478), .B(new_n3325), .Y(new_n22363));
  nand_5 g20015(.A(new_n3474), .B(n932), .Y(new_n22364));
  nand_5 g20016(.A(new_n3485), .B(new_n3328), .Y(new_n22365));
  nand_5 g20017(.A(new_n3481), .B(n6691), .Y(new_n22366));
  nand_5 g20018(.A(new_n3492), .B(new_n3331), .Y(new_n22367));
  nand_5 g20019(.A(new_n3488), .B(n3260), .Y(new_n22368));
  or_5   g20020(.A(new_n3495), .B(n20489), .Y(new_n22369));
  nand_5 g20021(.A(new_n3495), .B(n20489), .Y(new_n22370));
  or_5   g20022(.A(new_n3501), .B(n2355), .Y(new_n22371));
  nand_5 g20023(.A(new_n3501), .B(n2355), .Y(new_n22372));
  nand_5 g20024(.A(new_n3512), .B(new_n3340_1), .Y(new_n22373));
  nand_5 g20025(.A(new_n3511), .B(n11121), .Y(new_n22374));
  nand_5 g20026(.A(n16217), .B(n12315), .Y(new_n22375));
  nand_5 g20027(.A(new_n22375), .B(new_n22374), .Y(new_n22376));
  nand_5 g20028(.A(new_n22376), .B(new_n22373), .Y(new_n22377));
  nand_5 g20029(.A(new_n22377), .B(new_n22372), .Y(new_n22378));
  nand_5 g20030(.A(new_n22378), .B(new_n22371), .Y(new_n22379_1));
  nand_5 g20031(.A(new_n22379_1), .B(new_n22370), .Y(new_n22380));
  nand_5 g20032(.A(new_n22380), .B(new_n22369), .Y(new_n22381));
  nand_5 g20033(.A(new_n22381), .B(new_n22368), .Y(new_n22382));
  nand_5 g20034(.A(new_n22382), .B(new_n22367), .Y(new_n22383));
  nand_5 g20035(.A(new_n22383), .B(new_n22366), .Y(new_n22384));
  nand_5 g20036(.A(new_n22384), .B(new_n22365), .Y(new_n22385));
  nand_5 g20037(.A(new_n22385), .B(new_n22364), .Y(new_n22386));
  nand_5 g20038(.A(new_n22386), .B(new_n22363), .Y(new_n22387));
  nand_5 g20039(.A(new_n22387), .B(new_n22362), .Y(new_n22388));
  nand_5 g20040(.A(new_n22388), .B(new_n22361), .Y(new_n22389));
  nand_5 g20041(.A(new_n22389), .B(new_n22360), .Y(new_n22390));
  nand_5 g20042(.A(new_n22390), .B(new_n22359_1), .Y(new_n22391));
  nor_5  g20043(.A(new_n22391), .B(new_n22358_1), .Y(new_n22392));
  nand_5 g20044(.A(new_n3454), .B(n7335), .Y(new_n22393));
  nand_5 g20045(.A(new_n22393), .B(new_n3452), .Y(new_n22394));
  nor_5  g20046(.A(new_n22394), .B(new_n22392), .Y(new_n22395));
  not_8  g20047(.A(new_n22395), .Y(new_n22396));
  nor_5  g20048(.A(new_n22396), .B(new_n19374), .Y(new_n22397));
  and_5  g20049(.A(new_n22396), .B(new_n19374), .Y(new_n22398));
  nand_5 g20050(.A(new_n22393), .B(new_n22357), .Y(new_n22399));
  xor_4  g20051(.A(new_n22399), .B(new_n22391), .Y(new_n22400));
  or_5   g20052(.A(new_n22400), .B(new_n19418), .Y(new_n22401));
  nand_5 g20053(.A(new_n22400), .B(new_n19418), .Y(new_n22402));
  nand_5 g20054(.A(new_n22360), .B(new_n22359_1), .Y(new_n22403));
  xor_4  g20055(.A(new_n22403), .B(new_n22389), .Y(new_n22404));
  nand_5 g20056(.A(new_n22404), .B(new_n19425), .Y(new_n22405));
  or_5   g20057(.A(new_n22404), .B(new_n19425), .Y(new_n22406));
  nand_5 g20058(.A(new_n22362), .B(new_n22361), .Y(new_n22407));
  xor_4  g20059(.A(new_n22407), .B(new_n22387), .Y(new_n22408));
  nand_5 g20060(.A(new_n22408), .B(new_n19432), .Y(new_n22409));
  or_5   g20061(.A(new_n22408), .B(new_n19432), .Y(new_n22410));
  nand_5 g20062(.A(new_n22364), .B(new_n22363), .Y(new_n22411));
  xor_4  g20063(.A(new_n22411), .B(new_n22385), .Y(new_n22412));
  nand_5 g20064(.A(new_n22412), .B(new_n19439), .Y(new_n22413));
  or_5   g20065(.A(new_n22412), .B(new_n19439), .Y(new_n22414));
  nand_5 g20066(.A(new_n22366), .B(new_n22365), .Y(new_n22415));
  xor_4  g20067(.A(new_n22415), .B(new_n22383), .Y(new_n22416));
  nand_5 g20068(.A(new_n22416), .B(new_n19446), .Y(new_n22417));
  or_5   g20069(.A(new_n22416), .B(new_n19446), .Y(new_n22418));
  nand_5 g20070(.A(new_n22368), .B(new_n22367), .Y(new_n22419));
  xor_4  g20071(.A(new_n22419), .B(new_n22381), .Y(new_n22420));
  nand_5 g20072(.A(new_n22420), .B(new_n19453), .Y(new_n22421));
  or_5   g20073(.A(new_n22420), .B(new_n19453), .Y(new_n22422));
  nand_5 g20074(.A(new_n22370), .B(new_n22369), .Y(new_n22423));
  xor_4  g20075(.A(new_n22423), .B(new_n22379_1), .Y(new_n22424));
  nand_5 g20076(.A(new_n22424), .B(new_n19460), .Y(new_n22425));
  or_5   g20077(.A(new_n22424), .B(new_n19460), .Y(new_n22426));
  nand_5 g20078(.A(new_n22372), .B(new_n22371), .Y(new_n22427));
  xor_4  g20079(.A(new_n22427), .B(new_n22377), .Y(new_n22428));
  or_5   g20080(.A(new_n22428), .B(new_n19467_1), .Y(new_n22429));
  nand_5 g20081(.A(new_n22428), .B(new_n19467_1), .Y(new_n22430));
  nand_5 g20082(.A(new_n22374), .B(new_n22373), .Y(new_n22431));
  not_8  g20083(.A(new_n22431), .Y(new_n22432));
  nand_5 g20084(.A(new_n22432), .B(new_n22375), .Y(new_n22433_1));
  xor_4  g20085(.A(n16217), .B(n12315), .Y(new_n22434));
  nand_5 g20086(.A(new_n22434), .B(new_n19476), .Y(new_n22435));
  not_8  g20087(.A(new_n22435), .Y(new_n22436));
  nor_5  g20088(.A(new_n22432), .B(new_n22375), .Y(new_n22437));
  nor_5  g20089(.A(new_n22437), .B(new_n22436), .Y(new_n22438));
  nand_5 g20090(.A(new_n22438), .B(new_n22433_1), .Y(new_n22439));
  nand_5 g20091(.A(new_n22432), .B(new_n22436), .Y(new_n22440));
  nand_5 g20092(.A(new_n22440), .B(new_n19485), .Y(new_n22441));
  nand_5 g20093(.A(new_n22441), .B(new_n22439), .Y(new_n22442_1));
  nand_5 g20094(.A(new_n22442_1), .B(new_n22430), .Y(new_n22443));
  and_5  g20095(.A(new_n22443), .B(new_n22429), .Y(new_n22444_1));
  nand_5 g20096(.A(new_n22444_1), .B(new_n22426), .Y(new_n22445));
  nand_5 g20097(.A(new_n22445), .B(new_n22425), .Y(new_n22446));
  nand_5 g20098(.A(new_n22446), .B(new_n22422), .Y(new_n22447));
  nand_5 g20099(.A(new_n22447), .B(new_n22421), .Y(new_n22448));
  nand_5 g20100(.A(new_n22448), .B(new_n22418), .Y(new_n22449));
  nand_5 g20101(.A(new_n22449), .B(new_n22417), .Y(new_n22450));
  nand_5 g20102(.A(new_n22450), .B(new_n22414), .Y(new_n22451));
  nand_5 g20103(.A(new_n22451), .B(new_n22413), .Y(new_n22452));
  nand_5 g20104(.A(new_n22452), .B(new_n22410), .Y(new_n22453));
  nand_5 g20105(.A(new_n22453), .B(new_n22409), .Y(new_n22454));
  nand_5 g20106(.A(new_n22454), .B(new_n22406), .Y(new_n22455));
  nand_5 g20107(.A(new_n22455), .B(new_n22405), .Y(new_n22456));
  not_8  g20108(.A(new_n22456), .Y(new_n22457));
  nand_5 g20109(.A(new_n22457), .B(new_n22402), .Y(new_n22458));
  nand_5 g20110(.A(new_n22458), .B(new_n22401), .Y(new_n22459));
  nor_5  g20111(.A(new_n22459), .B(new_n22398), .Y(new_n22460));
  nor_5  g20112(.A(new_n22460), .B(new_n22397), .Y(new_n22461));
  nor_5  g20113(.A(new_n22395), .B(new_n19508), .Y(new_n22462));
  nor_5  g20114(.A(new_n22462), .B(new_n22461), .Y(new_n22463));
  nor_5  g20115(.A(new_n22396), .B(new_n19511), .Y(new_n22464));
  nor_5  g20116(.A(new_n22464), .B(new_n22460), .Y(new_n22465));
  nor_5  g20117(.A(new_n22465), .B(new_n22463), .Y(n6375));
  nor_5  g20118(.A(new_n21426), .B(new_n21425), .Y(new_n22467_1));
  xor_4  g20119(.A(new_n22467_1), .B(new_n21441), .Y(n6383));
  nor_5  g20120(.A(new_n16379_1), .B(new_n16377), .Y(new_n22469));
  xor_4  g20121(.A(new_n22469), .B(new_n16433_1), .Y(n6407));
  nand_5 g20122(.A(new_n9809), .B(new_n9808), .Y(new_n22471));
  xnor_4 g20123(.A(new_n22471), .B(new_n9814), .Y(n6431));
  nand_5 g20124(.A(new_n18723), .B(new_n18722), .Y(new_n22473));
  xnor_4 g20125(.A(new_n22473), .B(new_n18725_1), .Y(n6437));
  nand_5 g20126(.A(new_n4572), .B(new_n4571), .Y(new_n22475));
  xnor_4 g20127(.A(new_n22475), .B(new_n4581), .Y(n6457));
  nand_5 g20128(.A(new_n14056), .B(new_n14055), .Y(new_n22477));
  xor_4  g20129(.A(new_n22477), .B(new_n14086), .Y(n6465));
  not_8  g20130(.A(new_n9561), .Y(new_n22479));
  nand_5 g20131(.A(new_n19785), .B(new_n19780_1), .Y(new_n22480));
  not_8  g20132(.A(new_n22480), .Y(new_n22481));
  nand_5 g20133(.A(new_n19781), .B(new_n19778), .Y(new_n22482));
  nor_5  g20134(.A(new_n22482), .B(new_n22481), .Y(new_n22483));
  not_8  g20135(.A(new_n22483), .Y(new_n22484_1));
  nand_5 g20136(.A(new_n22484_1), .B(new_n22479), .Y(new_n22485));
  nand_5 g20137(.A(new_n22483), .B(new_n9561), .Y(new_n22486));
  nand_5 g20138(.A(new_n22486), .B(new_n22485), .Y(new_n22487));
  not_8  g20139(.A(new_n22487), .Y(new_n22488));
  nand_5 g20140(.A(new_n19787), .B(new_n3907), .Y(new_n22489_1));
  nand_5 g20141(.A(new_n19786), .B(new_n3906), .Y(new_n22490));
  nand_5 g20142(.A(new_n16451), .B(new_n16439_1), .Y(new_n22491));
  nand_5 g20143(.A(new_n22491), .B(new_n16449), .Y(new_n22492_1));
  nand_5 g20144(.A(new_n22492_1), .B(new_n22490), .Y(new_n22493));
  nand_5 g20145(.A(new_n22493), .B(new_n22489_1), .Y(new_n22494_1));
  nand_5 g20146(.A(new_n22494_1), .B(new_n22488), .Y(new_n22495));
  not_8  g20147(.A(new_n22495), .Y(new_n22496));
  nor_5  g20148(.A(new_n22494_1), .B(new_n22488), .Y(new_n22497));
  nor_5  g20149(.A(new_n22497), .B(new_n22496), .Y(new_n22498));
  nand_5 g20150(.A(new_n3769), .B(new_n3713), .Y(new_n22499));
  not_8  g20151(.A(new_n22499), .Y(new_n22500));
  nand_5 g20152(.A(new_n16458), .B(new_n16456), .Y(new_n22501));
  nand_5 g20153(.A(new_n22501), .B(new_n16457), .Y(new_n22502));
  nor_5  g20154(.A(new_n22502), .B(new_n22500), .Y(new_n22503));
  nand_5 g20155(.A(new_n3710_1), .B(n2743), .Y(new_n22504));
  nand_5 g20156(.A(new_n22504), .B(new_n3708), .Y(new_n22505));
  nor_5  g20157(.A(new_n22505), .B(new_n22503), .Y(new_n22506));
  nand_5 g20158(.A(new_n22506), .B(new_n22498), .Y(new_n22507));
  not_8  g20159(.A(new_n22498), .Y(new_n22508));
  not_8  g20160(.A(new_n22506), .Y(new_n22509));
  nand_5 g20161(.A(new_n22509), .B(new_n22508), .Y(new_n22510));
  nand_5 g20162(.A(new_n22510), .B(new_n22507), .Y(new_n22511));
  nand_5 g20163(.A(new_n22504), .B(new_n22499), .Y(new_n22512));
  xor_4  g20164(.A(new_n22512), .B(new_n22502), .Y(new_n22513));
  nand_5 g20165(.A(new_n22489_1), .B(new_n22490), .Y(new_n22514));
  xor_4  g20166(.A(new_n22514), .B(new_n22492_1), .Y(new_n22515));
  not_8  g20167(.A(new_n22515), .Y(new_n22516));
  or_5   g20168(.A(new_n22516), .B(new_n22513), .Y(new_n22517));
  nand_5 g20169(.A(new_n22516), .B(new_n22513), .Y(new_n22518));
  nor_5  g20170(.A(new_n16464), .B(new_n16437), .Y(new_n22519));
  nor_5  g20171(.A(new_n22519), .B(new_n16462), .Y(new_n22520));
  not_8  g20172(.A(new_n22520), .Y(new_n22521));
  nand_5 g20173(.A(new_n22521), .B(new_n22518), .Y(new_n22522));
  nand_5 g20174(.A(new_n22522), .B(new_n22517), .Y(new_n22523));
  xor_4  g20175(.A(new_n22523), .B(new_n22511), .Y(n6470));
  nand_5 g20176(.A(new_n13254), .B(new_n13253), .Y(new_n22525));
  xor_4  g20177(.A(new_n22525), .B(new_n13278), .Y(n6476));
  nand_5 g20178(.A(new_n20908), .B(new_n20909), .Y(new_n22527));
  xor_4  g20179(.A(new_n22527), .B(new_n20917), .Y(n6506));
  nand_5 g20180(.A(new_n10753), .B(new_n10748), .Y(new_n22529));
  nor_5  g20181(.A(new_n22529), .B(new_n10742), .Y(new_n22530));
  nand_5 g20182(.A(new_n22530), .B(new_n10738), .Y(new_n22531));
  nor_5  g20183(.A(new_n22531), .B(new_n10734), .Y(new_n22532));
  nand_5 g20184(.A(new_n22532), .B(new_n10770), .Y(new_n22533_1));
  xor_4  g20185(.A(new_n22533_1), .B(new_n10840), .Y(new_n22534));
  or_5   g20186(.A(new_n22534), .B(new_n10828), .Y(new_n22535));
  nand_5 g20187(.A(new_n22534), .B(new_n10828), .Y(new_n22536));
  xor_4  g20188(.A(new_n22532), .B(new_n10772), .Y(new_n22537));
  or_5   g20189(.A(new_n22537), .B(new_n10709), .Y(new_n22538));
  nand_5 g20190(.A(new_n22537), .B(new_n10709), .Y(new_n22539));
  xor_4  g20191(.A(new_n22531), .B(new_n10732), .Y(new_n22540));
  or_5   g20192(.A(new_n22540), .B(new_n10672), .Y(new_n22541));
  nand_5 g20193(.A(new_n22540), .B(new_n10672), .Y(new_n22542));
  xor_4  g20194(.A(new_n22530), .B(new_n10737), .Y(new_n22543));
  or_5   g20195(.A(new_n22543), .B(new_n10679), .Y(new_n22544));
  nand_5 g20196(.A(new_n22543), .B(new_n10679), .Y(new_n22545));
  xor_4  g20197(.A(new_n22529), .B(new_n10743), .Y(new_n22546));
  or_5   g20198(.A(new_n22546), .B(new_n10684), .Y(new_n22547));
  nand_5 g20199(.A(new_n22546), .B(new_n10684), .Y(new_n22548));
  nand_5 g20200(.A(new_n10754), .B(new_n10692_1), .Y(new_n22549));
  nor_5  g20201(.A(new_n22549), .B(new_n10686), .Y(new_n22550));
  not_8  g20202(.A(new_n22550), .Y(new_n22551));
  nand_5 g20203(.A(new_n22549), .B(new_n10689), .Y(new_n22552));
  xor_4  g20204(.A(new_n10754), .B(new_n10748), .Y(new_n22553));
  not_8  g20205(.A(new_n22553), .Y(new_n22554_1));
  nand_5 g20206(.A(new_n22554_1), .B(new_n22552), .Y(new_n22555));
  nand_5 g20207(.A(new_n22555), .B(new_n22551), .Y(new_n22556));
  nand_5 g20208(.A(new_n22556), .B(new_n22548), .Y(new_n22557));
  nand_5 g20209(.A(new_n22557), .B(new_n22547), .Y(new_n22558));
  nand_5 g20210(.A(new_n22558), .B(new_n22545), .Y(new_n22559));
  nand_5 g20211(.A(new_n22559), .B(new_n22544), .Y(new_n22560));
  nand_5 g20212(.A(new_n22560), .B(new_n22542), .Y(new_n22561));
  nand_5 g20213(.A(new_n22561), .B(new_n22541), .Y(new_n22562));
  nand_5 g20214(.A(new_n22562), .B(new_n22539), .Y(new_n22563));
  nand_5 g20215(.A(new_n22563), .B(new_n22538), .Y(new_n22564));
  nand_5 g20216(.A(new_n22564), .B(new_n22536), .Y(new_n22565));
  nand_5 g20217(.A(new_n22565), .B(new_n22535), .Y(new_n22566));
  nor_5  g20218(.A(new_n22533_1), .B(new_n10842), .Y(new_n22567));
  xor_4  g20219(.A(new_n22567), .B(new_n16074), .Y(new_n22568));
  or_5   g20220(.A(new_n22568), .B(new_n11657), .Y(new_n22569));
  nand_5 g20221(.A(new_n22568), .B(new_n11657), .Y(new_n22570));
  nand_5 g20222(.A(new_n22570), .B(new_n22569), .Y(new_n22571));
  xor_4  g20223(.A(new_n22571), .B(new_n22566), .Y(new_n22572));
  nand_5 g20224(.A(new_n22572), .B(new_n19015), .Y(new_n22573));
  or_5   g20225(.A(new_n22572), .B(new_n19015), .Y(new_n22574));
  nand_5 g20226(.A(new_n22536), .B(new_n22535), .Y(new_n22575));
  xor_4  g20227(.A(new_n22575), .B(new_n22564), .Y(new_n22576));
  nand_5 g20228(.A(new_n22576), .B(new_n18964), .Y(new_n22577));
  or_5   g20229(.A(new_n22576), .B(new_n18964), .Y(new_n22578));
  nand_5 g20230(.A(new_n22539), .B(new_n22538), .Y(new_n22579));
  xor_4  g20231(.A(new_n22579), .B(new_n22562), .Y(new_n22580));
  nand_5 g20232(.A(new_n22580), .B(new_n18969), .Y(new_n22581));
  or_5   g20233(.A(new_n22580), .B(new_n18969), .Y(new_n22582));
  nand_5 g20234(.A(new_n22542), .B(new_n22541), .Y(new_n22583));
  xor_4  g20235(.A(new_n22583), .B(new_n22560), .Y(new_n22584_1));
  nand_5 g20236(.A(new_n22584_1), .B(new_n18974), .Y(new_n22585));
  or_5   g20237(.A(new_n22584_1), .B(new_n18974), .Y(new_n22586));
  nand_5 g20238(.A(new_n22545), .B(new_n22544), .Y(new_n22587));
  xor_4  g20239(.A(new_n22587), .B(new_n22558), .Y(new_n22588_1));
  nand_5 g20240(.A(new_n22588_1), .B(new_n18979), .Y(new_n22589_1));
  or_5   g20241(.A(new_n22588_1), .B(new_n18979), .Y(new_n22590));
  nand_5 g20242(.A(new_n22548), .B(new_n22547), .Y(new_n22591_1));
  xor_4  g20243(.A(new_n22591_1), .B(new_n22556), .Y(new_n22592));
  nand_5 g20244(.A(new_n22592), .B(new_n18984), .Y(new_n22593));
  not_8  g20245(.A(new_n22593), .Y(new_n22594));
  nor_5  g20246(.A(new_n22592), .B(new_n18984), .Y(new_n22595));
  xor_4  g20247(.A(new_n10754), .B(new_n10692_1), .Y(new_n22596));
  nand_5 g20248(.A(new_n22596), .B(new_n18993), .Y(new_n22597_1));
  not_8  g20249(.A(new_n22597_1), .Y(new_n22598));
  nand_5 g20250(.A(new_n22598), .B(new_n18988), .Y(new_n22599));
  nand_5 g20251(.A(new_n22597_1), .B(new_n18989), .Y(new_n22600));
  nand_5 g20252(.A(new_n22552), .B(new_n22551), .Y(new_n22601));
  xor_4  g20253(.A(new_n22601), .B(new_n22553), .Y(new_n22602));
  nand_5 g20254(.A(new_n22602), .B(new_n22600), .Y(new_n22603));
  nand_5 g20255(.A(new_n22603), .B(new_n22599), .Y(new_n22604));
  nor_5  g20256(.A(new_n22604), .B(new_n22595), .Y(new_n22605));
  nor_5  g20257(.A(new_n22605), .B(new_n22594), .Y(new_n22606));
  not_8  g20258(.A(new_n22606), .Y(new_n22607));
  nand_5 g20259(.A(new_n22607), .B(new_n22590), .Y(new_n22608));
  nand_5 g20260(.A(new_n22608), .B(new_n22589_1), .Y(new_n22609));
  nand_5 g20261(.A(new_n22609), .B(new_n22586), .Y(new_n22610));
  nand_5 g20262(.A(new_n22610), .B(new_n22585), .Y(new_n22611));
  nand_5 g20263(.A(new_n22611), .B(new_n22582), .Y(new_n22612));
  nand_5 g20264(.A(new_n22612), .B(new_n22581), .Y(new_n22613));
  nand_5 g20265(.A(new_n22613), .B(new_n22578), .Y(new_n22614));
  nand_5 g20266(.A(new_n22614), .B(new_n22577), .Y(new_n22615));
  nand_5 g20267(.A(new_n22615), .B(new_n22574), .Y(new_n22616));
  nand_5 g20268(.A(new_n22616), .B(new_n22573), .Y(new_n22617));
  nand_5 g20269(.A(new_n22567), .B(new_n16075), .Y(new_n22618));
  nand_5 g20270(.A(new_n22618), .B(new_n16069), .Y(new_n22619_1));
  not_8  g20271(.A(new_n22618), .Y(new_n22620_1));
  nand_5 g20272(.A(new_n22620_1), .B(new_n16070), .Y(new_n22621));
  and_5  g20273(.A(new_n22621), .B(new_n22619_1), .Y(new_n22622));
  nand_5 g20274(.A(new_n22622), .B(new_n11651), .Y(new_n22623_1));
  or_5   g20275(.A(new_n22622), .B(new_n11651), .Y(new_n22624));
  nand_5 g20276(.A(new_n22624), .B(new_n22623_1), .Y(new_n22625));
  nand_5 g20277(.A(new_n22570), .B(new_n22566), .Y(new_n22626_1));
  nand_5 g20278(.A(new_n22626_1), .B(new_n22569), .Y(new_n22627));
  xor_4  g20279(.A(new_n22627), .B(new_n22625), .Y(new_n22628));
  nand_5 g20280(.A(new_n22628), .B(new_n19072), .Y(new_n22629));
  or_5   g20281(.A(new_n22628), .B(new_n19072), .Y(new_n22630));
  nand_5 g20282(.A(new_n22630), .B(new_n22629), .Y(new_n22631_1));
  xor_4  g20283(.A(new_n22631_1), .B(new_n22617), .Y(n6514));
  xor_4  g20284(.A(new_n13177), .B(new_n13162), .Y(new_n22633));
  nor_5  g20285(.A(new_n13172), .B(new_n13793), .Y(new_n22634));
  nor_5  g20286(.A(new_n13217), .B(new_n22634), .Y(new_n22635));
  xor_4  g20287(.A(new_n22635), .B(new_n22633), .Y(new_n22636));
  nand_5 g20288(.A(new_n13282), .B(new_n13240), .Y(new_n22637));
  nand_5 g20289(.A(new_n22637), .B(new_n13241), .Y(new_n22638));
  or_5   g20290(.A(new_n22638), .B(new_n22636), .Y(new_n22639));
  nand_5 g20291(.A(new_n22638), .B(new_n22636), .Y(new_n22640));
  nand_5 g20292(.A(new_n22640), .B(new_n22639), .Y(n6542));
  nand_5 g20293(.A(new_n17472), .B(new_n17473), .Y(new_n22642));
  xor_4  g20294(.A(new_n22642), .B(new_n17487), .Y(n6558));
  nand_5 g20295(.A(new_n20337), .B(new_n20338), .Y(new_n22644));
  xnor_4 g20296(.A(new_n22644), .B(new_n20340), .Y(n6560));
  nand_5 g20297(.A(new_n7137), .B(new_n4386), .Y(new_n22646));
  nand_5 g20298(.A(new_n7142), .B(n6773), .Y(new_n22647));
  nand_5 g20299(.A(new_n7138), .B(n17090), .Y(new_n22648));
  nand_5 g20300(.A(new_n22648), .B(new_n22647), .Y(new_n22649));
  nand_5 g20301(.A(new_n22649), .B(new_n22646), .Y(new_n22650));
  nand_5 g20302(.A(new_n14168), .B(new_n4376_1), .Y(new_n22651));
  nand_5 g20303(.A(new_n7132), .B(n11302), .Y(new_n22652));
  nand_5 g20304(.A(new_n22652), .B(new_n22651), .Y(new_n22653));
  xor_4  g20305(.A(new_n22653), .B(new_n22650), .Y(new_n22654));
  nand_5 g20306(.A(new_n22654), .B(new_n12567), .Y(new_n22655));
  or_5   g20307(.A(new_n22654), .B(new_n12567), .Y(new_n22656));
  not_8  g20308(.A(new_n11204), .Y(new_n22657));
  nand_5 g20309(.A(new_n22646), .B(new_n22648), .Y(new_n22658));
  xor_4  g20310(.A(new_n22658), .B(new_n22647), .Y(new_n22659));
  nand_5 g20311(.A(new_n22659), .B(new_n22657), .Y(new_n22660_1));
  or_5   g20312(.A(new_n22659), .B(new_n22657), .Y(new_n22661));
  nand_5 g20313(.A(new_n22661), .B(new_n20381), .Y(new_n22662));
  nand_5 g20314(.A(new_n22662), .B(new_n22660_1), .Y(new_n22663));
  nand_5 g20315(.A(new_n22663), .B(new_n22656), .Y(new_n22664));
  nand_5 g20316(.A(new_n22664), .B(new_n22655), .Y(new_n22665));
  nand_5 g20317(.A(new_n22652), .B(new_n22650), .Y(new_n22666));
  nand_5 g20318(.A(new_n22666), .B(new_n22651), .Y(new_n22667));
  nand_5 g20319(.A(new_n7128), .B(new_n4396), .Y(new_n22668));
  nand_5 g20320(.A(new_n7127), .B(n10405), .Y(new_n22669));
  nand_5 g20321(.A(new_n22669), .B(new_n22668), .Y(new_n22670));
  xnor_4 g20322(.A(new_n22670), .B(new_n22667), .Y(new_n22671));
  or_5   g20323(.A(new_n22671), .B(new_n11192_1), .Y(new_n22672));
  nand_5 g20324(.A(new_n22671), .B(new_n11192_1), .Y(new_n22673));
  nand_5 g20325(.A(new_n22673), .B(new_n22672), .Y(new_n22674));
  xnor_4 g20326(.A(new_n22674), .B(new_n22665), .Y(n6567));
  nor_5  g20327(.A(new_n15667), .B(n8324), .Y(new_n22676));
  nand_5 g20328(.A(new_n22676), .B(new_n9293), .Y(new_n22677));
  nor_5  g20329(.A(new_n22677), .B(n9445), .Y(new_n22678));
  nand_5 g20330(.A(new_n22678), .B(new_n9281), .Y(new_n22679));
  xor_4  g20331(.A(new_n22679), .B(n1536), .Y(new_n22680));
  nand_5 g20332(.A(new_n22680), .B(new_n4984), .Y(new_n22681));
  nor_5  g20333(.A(new_n22680), .B(new_n4984), .Y(new_n22682));
  not_8  g20334(.A(new_n22682), .Y(new_n22683));
  nand_5 g20335(.A(new_n22683), .B(new_n22681), .Y(new_n22684));
  xor_4  g20336(.A(new_n22678), .B(new_n9281), .Y(new_n22685));
  or_5   g20337(.A(new_n22685), .B(new_n4989), .Y(new_n22686));
  nand_5 g20338(.A(new_n22685), .B(new_n4989), .Y(new_n22687));
  xor_4  g20339(.A(new_n22677), .B(n9445), .Y(new_n22688));
  or_5   g20340(.A(new_n22688), .B(new_n4994), .Y(new_n22689));
  nand_5 g20341(.A(new_n22688), .B(new_n4994), .Y(new_n22690));
  xor_4  g20342(.A(new_n22676), .B(new_n9293), .Y(new_n22691));
  or_5   g20343(.A(new_n22691), .B(new_n4999), .Y(new_n22692));
  nand_5 g20344(.A(new_n22691), .B(new_n4999), .Y(new_n22693));
  nand_5 g20345(.A(new_n15670), .B(new_n15666), .Y(new_n22694));
  nand_5 g20346(.A(new_n22694), .B(new_n15669), .Y(new_n22695));
  nand_5 g20347(.A(new_n22695), .B(new_n22693), .Y(new_n22696));
  nand_5 g20348(.A(new_n22696), .B(new_n22692), .Y(new_n22697_1));
  nand_5 g20349(.A(new_n22697_1), .B(new_n22690), .Y(new_n22698));
  nand_5 g20350(.A(new_n22698), .B(new_n22689), .Y(new_n22699));
  nand_5 g20351(.A(new_n22699), .B(new_n22687), .Y(new_n22700));
  nand_5 g20352(.A(new_n22700), .B(new_n22686), .Y(new_n22701));
  xor_4  g20353(.A(new_n22701), .B(new_n22684), .Y(new_n22702));
  not_8  g20354(.A(new_n22702), .Y(new_n22703));
  nand_5 g20355(.A(new_n9279), .B(n23272), .Y(new_n22704));
  nand_5 g20356(.A(new_n9277), .B(new_n4850_1), .Y(new_n22705));
  nand_5 g20357(.A(new_n22705), .B(new_n22704), .Y(new_n22706));
  nand_5 g20358(.A(new_n9283), .B(new_n4856), .Y(new_n22707));
  nand_5 g20359(.A(new_n9285), .B(n11481), .Y(new_n22708));
  nand_5 g20360(.A(new_n9289), .B(new_n4862), .Y(new_n22709));
  nand_5 g20361(.A(new_n9291), .B(n16439), .Y(new_n22710));
  nand_5 g20362(.A(new_n9295), .B(new_n4868), .Y(new_n22711));
  nand_5 g20363(.A(new_n9297), .B(n15241), .Y(new_n22712));
  nand_5 g20364(.A(new_n15677), .B(new_n15675), .Y(new_n22713));
  nand_5 g20365(.A(new_n22713), .B(new_n15676), .Y(new_n22714_1));
  nand_5 g20366(.A(new_n22714_1), .B(new_n22712), .Y(new_n22715));
  nand_5 g20367(.A(new_n22715), .B(new_n22711), .Y(new_n22716));
  nand_5 g20368(.A(new_n22716), .B(new_n22710), .Y(new_n22717));
  nand_5 g20369(.A(new_n22717), .B(new_n22709), .Y(new_n22718));
  nand_5 g20370(.A(new_n22718), .B(new_n22708), .Y(new_n22719));
  nand_5 g20371(.A(new_n22719), .B(new_n22707), .Y(new_n22720));
  xnor_4 g20372(.A(new_n22720), .B(new_n22706), .Y(new_n22721));
  or_5   g20373(.A(new_n22721), .B(new_n22703), .Y(new_n22722));
  nand_5 g20374(.A(new_n22721), .B(new_n22703), .Y(new_n22723));
  nand_5 g20375(.A(new_n22723), .B(new_n22722), .Y(new_n22724));
  nand_5 g20376(.A(new_n22708), .B(new_n22707), .Y(new_n22725));
  xor_4  g20377(.A(new_n22725), .B(new_n22718), .Y(new_n22726));
  nand_5 g20378(.A(new_n22687), .B(new_n22686), .Y(new_n22727));
  xor_4  g20379(.A(new_n22727), .B(new_n22699), .Y(new_n22728));
  nand_5 g20380(.A(new_n22728), .B(new_n22726), .Y(new_n22729));
  or_5   g20381(.A(new_n22728), .B(new_n22726), .Y(new_n22730));
  nand_5 g20382(.A(new_n22710), .B(new_n22709), .Y(new_n22731));
  xor_4  g20383(.A(new_n22731), .B(new_n22716), .Y(new_n22732));
  nand_5 g20384(.A(new_n22690), .B(new_n22689), .Y(new_n22733));
  xor_4  g20385(.A(new_n22733), .B(new_n22697_1), .Y(new_n22734));
  nand_5 g20386(.A(new_n22734), .B(new_n22732), .Y(new_n22735));
  or_5   g20387(.A(new_n22734), .B(new_n22732), .Y(new_n22736));
  nand_5 g20388(.A(new_n22712), .B(new_n22711), .Y(new_n22737));
  xnor_4 g20389(.A(new_n22737), .B(new_n22714_1), .Y(new_n22738));
  nand_5 g20390(.A(new_n22693), .B(new_n22692), .Y(new_n22739));
  xor_4  g20391(.A(new_n22739), .B(new_n22695), .Y(new_n22740));
  not_8  g20392(.A(new_n22740), .Y(new_n22741));
  or_5   g20393(.A(new_n22741), .B(new_n22738), .Y(new_n22742));
  nand_5 g20394(.A(new_n22741), .B(new_n22738), .Y(new_n22743));
  nand_5 g20395(.A(new_n15681), .B(new_n15664), .Y(new_n22744));
  nand_5 g20396(.A(new_n22744), .B(new_n15680), .Y(new_n22745));
  nand_5 g20397(.A(new_n22745), .B(new_n22743), .Y(new_n22746));
  nand_5 g20398(.A(new_n22746), .B(new_n22742), .Y(new_n22747));
  nand_5 g20399(.A(new_n22747), .B(new_n22736), .Y(new_n22748));
  nand_5 g20400(.A(new_n22748), .B(new_n22735), .Y(new_n22749));
  nand_5 g20401(.A(new_n22749), .B(new_n22730), .Y(new_n22750));
  nand_5 g20402(.A(new_n22750), .B(new_n22729), .Y(new_n22751));
  xnor_4 g20403(.A(new_n22751), .B(new_n22724), .Y(n6576));
  nand_5 g20404(.A(new_n22439), .B(new_n22440), .Y(new_n22753));
  xor_4  g20405(.A(new_n22753), .B(new_n19485), .Y(n6587));
  nand_5 g20406(.A(new_n21217), .B(new_n21216), .Y(new_n22755));
  xnor_4 g20407(.A(new_n22755), .B(new_n21273), .Y(n6612));
  nand_5 g20408(.A(new_n19995), .B(new_n19735), .Y(new_n22757));
  nand_5 g20409(.A(new_n19739), .B(new_n12408_1), .Y(new_n22758));
  nand_5 g20410(.A(new_n19737), .B(new_n19999), .Y(new_n22759));
  nand_5 g20411(.A(new_n19743), .B(new_n12398_1), .Y(new_n22760));
  nand_5 g20412(.A(new_n19742), .B(new_n12399), .Y(new_n22761_1));
  nand_5 g20413(.A(new_n19747), .B(new_n12388), .Y(new_n22762));
  nand_5 g20414(.A(new_n19746), .B(new_n12389), .Y(new_n22763));
  nand_5 g20415(.A(new_n19751), .B(new_n12380_1), .Y(new_n22764_1));
  nand_5 g20416(.A(new_n19750), .B(new_n18645), .Y(new_n22765));
  nand_5 g20417(.A(new_n19755), .B(new_n12372), .Y(new_n22766));
  nand_5 g20418(.A(new_n19754), .B(new_n12373), .Y(new_n22767));
  nand_5 g20419(.A(new_n19760), .B(new_n12364_1), .Y(new_n22768));
  nand_5 g20420(.A(new_n19759), .B(new_n17541), .Y(new_n22769));
  nand_5 g20421(.A(new_n17198), .B(new_n12437), .Y(new_n22770));
  nand_5 g20422(.A(new_n17197), .B(new_n12357), .Y(new_n22771));
  nand_5 g20423(.A(new_n17172), .B(new_n12348), .Y(new_n22772));
  nand_5 g20424(.A(new_n17171), .B(new_n12347), .Y(new_n22773));
  nand_5 g20425(.A(new_n12444), .B(new_n7558_1), .Y(new_n22774));
  nand_5 g20426(.A(new_n22774), .B(new_n17162), .Y(new_n22775));
  nand_5 g20427(.A(new_n17168_1), .B(new_n12444), .Y(new_n22776));
  nand_5 g20428(.A(new_n22776), .B(new_n12338), .Y(new_n22777));
  nand_5 g20429(.A(new_n22777), .B(new_n22775), .Y(new_n22778));
  not_8  g20430(.A(new_n22778), .Y(new_n22779_1));
  nand_5 g20431(.A(new_n22779_1), .B(new_n22773), .Y(new_n22780));
  nand_5 g20432(.A(new_n22780), .B(new_n22772), .Y(new_n22781));
  nand_5 g20433(.A(new_n22781), .B(new_n22771), .Y(new_n22782));
  nand_5 g20434(.A(new_n22782), .B(new_n22770), .Y(new_n22783));
  nand_5 g20435(.A(new_n22783), .B(new_n22769), .Y(new_n22784));
  nand_5 g20436(.A(new_n22784), .B(new_n22768), .Y(new_n22785));
  nand_5 g20437(.A(new_n22785), .B(new_n22767), .Y(new_n22786));
  nand_5 g20438(.A(new_n22786), .B(new_n22766), .Y(new_n22787_1));
  nand_5 g20439(.A(new_n22787_1), .B(new_n22765), .Y(new_n22788));
  nand_5 g20440(.A(new_n22788), .B(new_n22764_1), .Y(new_n22789));
  nand_5 g20441(.A(new_n22789), .B(new_n22763), .Y(new_n22790));
  nand_5 g20442(.A(new_n22790), .B(new_n22762), .Y(new_n22791));
  nand_5 g20443(.A(new_n22791), .B(new_n22761_1), .Y(new_n22792));
  nand_5 g20444(.A(new_n22792), .B(new_n22760), .Y(new_n22793_1));
  nand_5 g20445(.A(new_n22793_1), .B(new_n22759), .Y(new_n22794));
  nand_5 g20446(.A(new_n22794), .B(new_n22758), .Y(new_n22795));
  nor_5  g20447(.A(new_n22795), .B(new_n22757), .Y(new_n22796));
  not_8  g20448(.A(new_n22795), .Y(new_n22797));
  nand_5 g20449(.A(new_n19996), .B(new_n19736_1), .Y(new_n22798));
  nor_5  g20450(.A(new_n22798), .B(new_n22797), .Y(new_n22799));
  nor_5  g20451(.A(new_n22799), .B(new_n22796), .Y(new_n22800));
  and_5  g20452(.A(new_n22798), .B(new_n22757), .Y(new_n22801));
  xor_4  g20453(.A(new_n22801), .B(new_n22795), .Y(new_n22802));
  or_5   g20454(.A(new_n22802), .B(new_n21982), .Y(new_n22803));
  nand_5 g20455(.A(new_n22759), .B(new_n22758), .Y(new_n22804));
  xor_4  g20456(.A(new_n22804), .B(new_n22793_1), .Y(new_n22805));
  nand_5 g20457(.A(new_n22805), .B(new_n21989), .Y(new_n22806));
  nor_5  g20458(.A(new_n22805), .B(new_n21989), .Y(new_n22807));
  not_8  g20459(.A(new_n22807), .Y(new_n22808));
  nand_5 g20460(.A(new_n22761_1), .B(new_n22760), .Y(new_n22809));
  xor_4  g20461(.A(new_n22809), .B(new_n22791), .Y(new_n22810));
  nand_5 g20462(.A(new_n22810), .B(new_n21994), .Y(new_n22811));
  nor_5  g20463(.A(new_n22810), .B(new_n21994), .Y(new_n22812));
  not_8  g20464(.A(new_n22812), .Y(new_n22813));
  nand_5 g20465(.A(new_n22763), .B(new_n22762), .Y(new_n22814));
  xor_4  g20466(.A(new_n22814), .B(new_n22789), .Y(new_n22815));
  nand_5 g20467(.A(new_n22815), .B(new_n22000), .Y(new_n22816));
  nor_5  g20468(.A(new_n22815), .B(new_n22000), .Y(new_n22817));
  not_8  g20469(.A(new_n22817), .Y(new_n22818));
  nand_5 g20470(.A(new_n22765), .B(new_n22764_1), .Y(new_n22819_1));
  xor_4  g20471(.A(new_n22819_1), .B(new_n22787_1), .Y(new_n22820));
  nand_5 g20472(.A(new_n22820), .B(new_n10845), .Y(new_n22821));
  nor_5  g20473(.A(new_n22820), .B(new_n10845), .Y(new_n22822));
  not_8  g20474(.A(new_n22822), .Y(new_n22823));
  nand_5 g20475(.A(new_n22767), .B(new_n22766), .Y(new_n22824));
  xor_4  g20476(.A(new_n22824), .B(new_n22785), .Y(new_n22825));
  nand_5 g20477(.A(new_n22825), .B(new_n10775_1), .Y(new_n22826));
  nor_5  g20478(.A(new_n22825), .B(new_n10775_1), .Y(new_n22827));
  not_8  g20479(.A(new_n22827), .Y(new_n22828));
  nand_5 g20480(.A(new_n22769), .B(new_n22768), .Y(new_n22829));
  xor_4  g20481(.A(new_n22829), .B(new_n22783), .Y(new_n22830));
  nand_5 g20482(.A(new_n22830), .B(new_n10779), .Y(new_n22831));
  nor_5  g20483(.A(new_n22830), .B(new_n10779), .Y(new_n22832));
  not_8  g20484(.A(new_n22832), .Y(new_n22833));
  nand_5 g20485(.A(new_n22771), .B(new_n22770), .Y(new_n22834));
  xor_4  g20486(.A(new_n22834), .B(new_n22781), .Y(new_n22835));
  nand_5 g20487(.A(new_n22835), .B(new_n10787), .Y(new_n22836));
  or_5   g20488(.A(new_n22835), .B(new_n10787), .Y(new_n22837));
  nand_5 g20489(.A(new_n22773), .B(new_n22772), .Y(new_n22838));
  xor_4  g20490(.A(new_n22838), .B(new_n22779_1), .Y(new_n22839));
  nor_5  g20491(.A(new_n22839), .B(new_n10793), .Y(new_n22840));
  and_5  g20492(.A(new_n22839), .B(new_n10793), .Y(new_n22841));
  and_5  g20493(.A(new_n22776), .B(new_n22775), .Y(new_n22842));
  xor_4  g20494(.A(new_n22842), .B(new_n12338), .Y(new_n22843_1));
  or_5   g20495(.A(new_n22843_1), .B(new_n10797), .Y(new_n22844));
  nand_5 g20496(.A(new_n22843_1), .B(new_n10797), .Y(new_n22845));
  xor_4  g20497(.A(new_n12333), .B(n18), .Y(new_n22846));
  nor_5  g20498(.A(new_n22846), .B(new_n20559), .Y(new_n22847));
  not_8  g20499(.A(new_n22847), .Y(new_n22848));
  nand_5 g20500(.A(new_n22848), .B(new_n22845), .Y(new_n22849));
  and_5  g20501(.A(new_n22849), .B(new_n22844), .Y(new_n22850));
  nor_5  g20502(.A(new_n22850), .B(new_n22841), .Y(new_n22851));
  nor_5  g20503(.A(new_n22851), .B(new_n22840), .Y(new_n22852));
  nand_5 g20504(.A(new_n22852), .B(new_n22837), .Y(new_n22853));
  nand_5 g20505(.A(new_n22853), .B(new_n22836), .Y(new_n22854));
  nand_5 g20506(.A(new_n22854), .B(new_n22833), .Y(new_n22855));
  nand_5 g20507(.A(new_n22855), .B(new_n22831), .Y(new_n22856));
  nand_5 g20508(.A(new_n22856), .B(new_n22828), .Y(new_n22857));
  nand_5 g20509(.A(new_n22857), .B(new_n22826), .Y(new_n22858_1));
  nand_5 g20510(.A(new_n22858_1), .B(new_n22823), .Y(new_n22859));
  nand_5 g20511(.A(new_n22859), .B(new_n22821), .Y(new_n22860));
  nand_5 g20512(.A(new_n22860), .B(new_n22818), .Y(new_n22861));
  nand_5 g20513(.A(new_n22861), .B(new_n22816), .Y(new_n22862));
  nand_5 g20514(.A(new_n22862), .B(new_n22813), .Y(new_n22863));
  nand_5 g20515(.A(new_n22863), .B(new_n22811), .Y(new_n22864));
  nand_5 g20516(.A(new_n22864), .B(new_n22808), .Y(new_n22865));
  nand_5 g20517(.A(new_n22865), .B(new_n22806), .Y(new_n22866));
  nand_5 g20518(.A(new_n22866), .B(new_n22803), .Y(new_n22867));
  nand_5 g20519(.A(new_n22802), .B(new_n21982), .Y(new_n22868));
  nand_5 g20520(.A(new_n22868), .B(new_n22867), .Y(new_n22869));
  nand_5 g20521(.A(new_n22869), .B(new_n21979), .Y(new_n22870_1));
  or_5   g20522(.A(new_n22869), .B(new_n21979), .Y(new_n22871_1));
  nand_5 g20523(.A(new_n22871_1), .B(new_n22870_1), .Y(new_n22872));
  xnor_4 g20524(.A(new_n22872), .B(new_n22800), .Y(n6628));
  nand_5 g20525(.A(new_n2957), .B(new_n2956), .Y(new_n22874));
  xnor_4 g20526(.A(new_n22874), .B(new_n2982), .Y(n6630));
  nand_5 g20527(.A(n23923), .B(new_n2599), .Y(new_n22876));
  nand_5 g20528(.A(new_n8028), .B(n9942), .Y(new_n22877));
  nand_5 g20529(.A(new_n2516), .B(n329), .Y(new_n22878));
  nand_5 g20530(.A(n25643), .B(new_n8031_1), .Y(new_n22879_1));
  nand_5 g20531(.A(n24170), .B(new_n2490), .Y(new_n22880));
  nand_5 g20532(.A(new_n8052_1), .B(n9557), .Y(new_n22881));
  nand_5 g20533(.A(new_n2494), .B(n2409), .Y(new_n22882));
  nand_5 g20534(.A(n3136), .B(new_n8034), .Y(new_n22883));
  nand_5 g20535(.A(new_n21650), .B(new_n21648), .Y(new_n22884));
  nand_5 g20536(.A(new_n22884), .B(new_n21649_1), .Y(new_n22885));
  nand_5 g20537(.A(new_n22885), .B(new_n22883), .Y(new_n22886));
  nand_5 g20538(.A(new_n22886), .B(new_n22882), .Y(new_n22887));
  nand_5 g20539(.A(new_n22887), .B(new_n22881), .Y(new_n22888));
  nand_5 g20540(.A(new_n22888), .B(new_n22880), .Y(new_n22889));
  nand_5 g20541(.A(new_n22889), .B(new_n22879_1), .Y(new_n22890));
  nand_5 g20542(.A(new_n22890), .B(new_n22878), .Y(new_n22891_1));
  nand_5 g20543(.A(new_n22891_1), .B(new_n22877), .Y(new_n22892));
  nand_5 g20544(.A(new_n22892), .B(new_n22876), .Y(new_n22893));
  nand_5 g20545(.A(new_n7998), .B(n5400), .Y(new_n22894));
  nand_5 g20546(.A(n16482), .B(new_n8023), .Y(new_n22895));
  nand_5 g20547(.A(new_n22895), .B(new_n22894), .Y(new_n22896));
  xor_4  g20548(.A(new_n22896), .B(new_n22893), .Y(new_n22897_1));
  or_5   g20549(.A(new_n22897_1), .B(new_n22104), .Y(new_n22898));
  nand_5 g20550(.A(new_n22897_1), .B(new_n22104), .Y(new_n22899));
  nand_5 g20551(.A(new_n22877), .B(new_n22876), .Y(new_n22900));
  xor_4  g20552(.A(new_n22900), .B(new_n22891_1), .Y(new_n22901));
  or_5   g20553(.A(new_n22901), .B(new_n22075), .Y(new_n22902));
  nand_5 g20554(.A(new_n22901), .B(new_n22075), .Y(new_n22903_1));
  nand_5 g20555(.A(new_n22879_1), .B(new_n22878), .Y(new_n22904));
  xor_4  g20556(.A(new_n22904), .B(new_n22889), .Y(new_n22905));
  or_5   g20557(.A(new_n22905), .B(new_n21745), .Y(new_n22906));
  nand_5 g20558(.A(new_n22905), .B(new_n21745), .Y(new_n22907_1));
  nand_5 g20559(.A(new_n22881), .B(new_n22880), .Y(new_n22908));
  xor_4  g20560(.A(new_n22908), .B(new_n22887), .Y(new_n22909));
  or_5   g20561(.A(new_n22909), .B(new_n21683), .Y(new_n22910_1));
  nand_5 g20562(.A(new_n22909), .B(new_n21683), .Y(new_n22911));
  nand_5 g20563(.A(new_n22883), .B(new_n22882), .Y(new_n22912));
  xor_4  g20564(.A(new_n22912), .B(new_n22885), .Y(new_n22913));
  or_5   g20565(.A(new_n22913), .B(new_n21706), .Y(new_n22914_1));
  nand_5 g20566(.A(new_n22913), .B(new_n21706), .Y(new_n22915));
  nand_5 g20567(.A(new_n21654_1), .B(new_n21633), .Y(new_n22916));
  nand_5 g20568(.A(new_n22916), .B(new_n21653), .Y(new_n22917));
  nand_5 g20569(.A(new_n22917), .B(new_n22915), .Y(new_n22918_1));
  nand_5 g20570(.A(new_n22918_1), .B(new_n22914_1), .Y(new_n22919));
  nand_5 g20571(.A(new_n22919), .B(new_n22911), .Y(new_n22920));
  nand_5 g20572(.A(new_n22920), .B(new_n22910_1), .Y(new_n22921));
  nand_5 g20573(.A(new_n22921), .B(new_n22907_1), .Y(new_n22922));
  nand_5 g20574(.A(new_n22922), .B(new_n22906), .Y(new_n22923));
  nand_5 g20575(.A(new_n22923), .B(new_n22903_1), .Y(new_n22924));
  nand_5 g20576(.A(new_n22924), .B(new_n22902), .Y(new_n22925));
  nand_5 g20577(.A(new_n22925), .B(new_n22899), .Y(new_n22926));
  nand_5 g20578(.A(new_n22926), .B(new_n22898), .Y(new_n22927));
  nand_5 g20579(.A(new_n22102), .B(new_n22092), .Y(new_n22928));
  nand_5 g20580(.A(new_n22928), .B(new_n22101), .Y(new_n22929));
  not_8  g20581(.A(new_n22097), .Y(new_n22930));
  not_8  g20582(.A(new_n22098), .Y(new_n22931));
  nor_5  g20583(.A(new_n22931), .B(new_n22096), .Y(new_n22932));
  nor_5  g20584(.A(new_n22932), .B(new_n22930), .Y(new_n22933));
  nand_5 g20585(.A(new_n8146), .B(new_n18127), .Y(new_n22934));
  nand_5 g20586(.A(n25331), .B(n17911), .Y(new_n22935));
  nand_5 g20587(.A(new_n22935), .B(new_n22934), .Y(new_n22936));
  xor_4  g20588(.A(new_n22936), .B(new_n22933), .Y(new_n22937));
  or_5   g20589(.A(new_n22937), .B(new_n8581_1), .Y(new_n22938));
  nand_5 g20590(.A(new_n22937), .B(new_n8581_1), .Y(new_n22939_1));
  nand_5 g20591(.A(new_n22939_1), .B(new_n22938), .Y(new_n22940));
  xor_4  g20592(.A(new_n22940), .B(new_n22929), .Y(new_n22941));
  not_8  g20593(.A(new_n22941), .Y(new_n22942));
  nand_5 g20594(.A(new_n22895), .B(new_n22893), .Y(new_n22943));
  nand_5 g20595(.A(new_n22943), .B(new_n22894), .Y(new_n22944));
  nand_5 g20596(.A(new_n3849), .B(n468), .Y(new_n22945));
  nand_5 g20597(.A(n14130), .B(new_n8019), .Y(new_n22946));
  nand_5 g20598(.A(new_n22946), .B(new_n22945), .Y(new_n22947));
  xnor_4 g20599(.A(new_n22947), .B(new_n22944), .Y(new_n22948));
  nand_5 g20600(.A(new_n22948), .B(new_n22942), .Y(new_n22949));
  not_8  g20601(.A(new_n22949), .Y(new_n22950));
  nor_5  g20602(.A(new_n22948), .B(new_n22942), .Y(new_n22951));
  nor_5  g20603(.A(new_n22951), .B(new_n22950), .Y(new_n22952));
  xor_4  g20604(.A(new_n22952), .B(new_n22927), .Y(n6634));
  nand_5 g20605(.A(new_n7441), .B(new_n7443), .Y(new_n22954));
  xor_4  g20606(.A(new_n22954), .B(new_n7459), .Y(n6652));
  nand_5 g20607(.A(new_n14345_1), .B(new_n14344), .Y(new_n22956));
  xor_4  g20608(.A(new_n22956), .B(new_n14358), .Y(n6655));
  nand_5 g20609(.A(new_n13820), .B(new_n13819), .Y(new_n22958));
  xor_4  g20610(.A(new_n22958), .B(new_n13841), .Y(n6669));
  nand_5 g20611(.A(new_n10788), .B(new_n10789), .Y(new_n22960));
  xnor_4 g20612(.A(new_n22960), .B(new_n10811), .Y(n6671));
  nand_5 g20613(.A(new_n15442), .B(new_n15441), .Y(new_n22962));
  xnor_4 g20614(.A(new_n22962), .B(new_n15462), .Y(n6673));
  nor_5  g20615(.A(new_n13172), .B(new_n13162), .Y(new_n22964));
  nand_5 g20616(.A(new_n22635), .B(new_n22964), .Y(new_n22965));
  nand_5 g20617(.A(new_n22965), .B(new_n22640), .Y(n6674));
  nand_5 g20618(.A(new_n18901_1), .B(new_n18900), .Y(new_n22967));
  xnor_4 g20619(.A(new_n22967), .B(new_n18909), .Y(n6684));
  xor_4  g20620(.A(new_n14092), .B(new_n14047), .Y(n6706));
  nor_5  g20621(.A(new_n22701), .B(new_n22682), .Y(new_n22970));
  or_5   g20622(.A(new_n22679), .B(n1536), .Y(new_n22971));
  nand_5 g20623(.A(new_n22681), .B(new_n22971), .Y(new_n22972));
  nor_5  g20624(.A(new_n22972), .B(new_n22970), .Y(new_n22973));
  nor_5  g20625(.A(new_n22973), .B(new_n4979), .Y(new_n22974));
  nand_5 g20626(.A(new_n22973), .B(new_n4979), .Y(new_n22975));
  not_8  g20627(.A(new_n22975), .Y(new_n22976));
  nor_5  g20628(.A(new_n22976), .B(new_n22974), .Y(new_n22977));
  not_8  g20629(.A(new_n22977), .Y(new_n22978));
  nand_5 g20630(.A(new_n9271), .B(new_n6382), .Y(new_n22979));
  nand_5 g20631(.A(n12702), .B(n8614), .Y(new_n22980));
  nand_5 g20632(.A(new_n22980), .B(new_n22979), .Y(new_n22981));
  nand_5 g20633(.A(new_n6168), .B(new_n6386), .Y(new_n22982));
  nand_5 g20634(.A(n26797), .B(n15182), .Y(new_n22983));
  nand_5 g20635(.A(new_n6390), .B(new_n9235), .Y(new_n22984));
  nand_5 g20636(.A(n27037), .B(n23913), .Y(new_n22985));
  nand_5 g20637(.A(new_n6169), .B(new_n6394), .Y(new_n22986));
  nand_5 g20638(.A(n22554), .B(n8964), .Y(new_n22987));
  nand_5 g20639(.A(new_n9241), .B(new_n4512), .Y(new_n22988));
  nand_5 g20640(.A(n20429), .B(n20151), .Y(new_n22989));
  nand_5 g20641(.A(new_n4438), .B(new_n6170), .Y(new_n22990));
  nand_5 g20642(.A(n7693), .B(n3909), .Y(new_n22991));
  nand_5 g20643(.A(new_n9247), .B(new_n4396), .Y(new_n22992));
  nand_5 g20644(.A(n23974), .B(n10405), .Y(new_n22993));
  nand_5 g20645(.A(new_n4376_1), .B(new_n9251_1), .Y(new_n22994));
  nand_5 g20646(.A(n11302), .B(n2146), .Y(new_n22995));
  nand_5 g20647(.A(new_n17863), .B(new_n17853), .Y(new_n22996));
  nand_5 g20648(.A(new_n22996), .B(new_n17862), .Y(new_n22997));
  nand_5 g20649(.A(new_n22997), .B(new_n22995), .Y(new_n22998_1));
  nand_5 g20650(.A(new_n22998_1), .B(new_n22994), .Y(new_n22999));
  nand_5 g20651(.A(new_n22999), .B(new_n22993), .Y(new_n23000));
  nand_5 g20652(.A(new_n23000), .B(new_n22992), .Y(new_n23001));
  nand_5 g20653(.A(new_n23001), .B(new_n22991), .Y(new_n23002));
  nand_5 g20654(.A(new_n23002), .B(new_n22990), .Y(new_n23003));
  nand_5 g20655(.A(new_n23003), .B(new_n22989), .Y(new_n23004));
  nand_5 g20656(.A(new_n23004), .B(new_n22988), .Y(new_n23005));
  nand_5 g20657(.A(new_n23005), .B(new_n22987), .Y(new_n23006_1));
  nand_5 g20658(.A(new_n23006_1), .B(new_n22986), .Y(new_n23007_1));
  nand_5 g20659(.A(new_n23007_1), .B(new_n22985), .Y(new_n23008));
  nand_5 g20660(.A(new_n23008), .B(new_n22984), .Y(new_n23009_1));
  nand_5 g20661(.A(new_n23009_1), .B(new_n22983), .Y(new_n23010));
  nand_5 g20662(.A(new_n23010), .B(new_n22982), .Y(new_n23011));
  xor_4  g20663(.A(new_n23011), .B(new_n22981), .Y(new_n23012));
  nand_5 g20664(.A(new_n23012), .B(new_n15931), .Y(new_n23013));
  or_5   g20665(.A(new_n23012), .B(new_n15931), .Y(new_n23014_1));
  nand_5 g20666(.A(new_n22983), .B(new_n22982), .Y(new_n23015));
  xor_4  g20667(.A(new_n23015), .B(new_n23009_1), .Y(new_n23016));
  nand_5 g20668(.A(new_n23016), .B(new_n6992), .Y(new_n23017));
  or_5   g20669(.A(new_n23016), .B(new_n6992), .Y(new_n23018));
  nand_5 g20670(.A(new_n22985), .B(new_n22984), .Y(new_n23019));
  xor_4  g20671(.A(new_n23019), .B(new_n23007_1), .Y(new_n23020));
  nand_5 g20672(.A(new_n23020), .B(new_n6998_1), .Y(new_n23021));
  or_5   g20673(.A(new_n23020), .B(new_n6998_1), .Y(new_n23022));
  nand_5 g20674(.A(new_n22987), .B(new_n22986), .Y(new_n23023));
  xor_4  g20675(.A(new_n23023), .B(new_n23005), .Y(new_n23024));
  nand_5 g20676(.A(new_n23024), .B(new_n7004), .Y(new_n23025));
  or_5   g20677(.A(new_n23024), .B(new_n7004), .Y(new_n23026));
  nand_5 g20678(.A(new_n22989), .B(new_n22988), .Y(new_n23027));
  xor_4  g20679(.A(new_n23027), .B(new_n23003), .Y(new_n23028));
  nand_5 g20680(.A(new_n23028), .B(new_n4522), .Y(new_n23029));
  or_5   g20681(.A(new_n23028), .B(new_n4522), .Y(new_n23030));
  nand_5 g20682(.A(new_n22991), .B(new_n22990), .Y(new_n23031));
  xor_4  g20683(.A(new_n23031), .B(new_n23001), .Y(new_n23032));
  nand_5 g20684(.A(new_n23032), .B(new_n4523), .Y(new_n23033));
  or_5   g20685(.A(new_n23032), .B(new_n4523), .Y(new_n23034));
  nand_5 g20686(.A(new_n22993), .B(new_n22992), .Y(new_n23035_1));
  xor_4  g20687(.A(new_n23035_1), .B(new_n22999), .Y(new_n23036));
  nand_5 g20688(.A(new_n23036), .B(new_n4407), .Y(new_n23037));
  or_5   g20689(.A(new_n23036), .B(new_n4407), .Y(new_n23038));
  nand_5 g20690(.A(new_n22995), .B(new_n22994), .Y(new_n23039_1));
  xor_4  g20691(.A(new_n23039_1), .B(new_n22997), .Y(new_n23040));
  nand_5 g20692(.A(new_n23040), .B(new_n4408), .Y(new_n23041));
  or_5   g20693(.A(new_n23040), .B(new_n4408), .Y(new_n23042));
  nand_5 g20694(.A(new_n17867), .B(new_n17856), .Y(new_n23043));
  nand_5 g20695(.A(new_n23043), .B(new_n17866), .Y(new_n23044));
  nand_5 g20696(.A(new_n23044), .B(new_n23042), .Y(new_n23045));
  nand_5 g20697(.A(new_n23045), .B(new_n23041), .Y(new_n23046));
  nand_5 g20698(.A(new_n23046), .B(new_n23038), .Y(new_n23047_1));
  nand_5 g20699(.A(new_n23047_1), .B(new_n23037), .Y(new_n23048));
  nand_5 g20700(.A(new_n23048), .B(new_n23034), .Y(new_n23049));
  nand_5 g20701(.A(new_n23049), .B(new_n23033), .Y(new_n23050));
  nand_5 g20702(.A(new_n23050), .B(new_n23030), .Y(new_n23051));
  nand_5 g20703(.A(new_n23051), .B(new_n23029), .Y(new_n23052));
  nand_5 g20704(.A(new_n23052), .B(new_n23026), .Y(new_n23053));
  nand_5 g20705(.A(new_n23053), .B(new_n23025), .Y(new_n23054));
  nand_5 g20706(.A(new_n23054), .B(new_n23022), .Y(new_n23055));
  nand_5 g20707(.A(new_n23055), .B(new_n23021), .Y(new_n23056));
  nand_5 g20708(.A(new_n23056), .B(new_n23018), .Y(new_n23057));
  nand_5 g20709(.A(new_n23057), .B(new_n23017), .Y(new_n23058_1));
  nand_5 g20710(.A(new_n23058_1), .B(new_n23014_1), .Y(new_n23059));
  nand_5 g20711(.A(new_n23059), .B(new_n23013), .Y(new_n23060));
  nand_5 g20712(.A(new_n23011), .B(new_n22980), .Y(new_n23061));
  nand_5 g20713(.A(new_n23061), .B(new_n22979), .Y(new_n23062));
  not_8  g20714(.A(new_n23062), .Y(new_n23063));
  nor_5  g20715(.A(new_n23063), .B(new_n23060), .Y(new_n23064));
  not_8  g20716(.A(new_n23064), .Y(new_n23065_1));
  nand_5 g20717(.A(new_n23063), .B(new_n23060), .Y(new_n23066_1));
  nand_5 g20718(.A(new_n23066_1), .B(new_n23065_1), .Y(new_n23067_1));
  nor_5  g20719(.A(new_n23067_1), .B(new_n22978), .Y(new_n23068_1));
  and_5  g20720(.A(new_n23067_1), .B(new_n22978), .Y(new_n23069));
  nor_5  g20721(.A(new_n23069), .B(new_n23068_1), .Y(new_n23070));
  nand_5 g20722(.A(new_n23014_1), .B(new_n23013), .Y(new_n23071));
  xor_4  g20723(.A(new_n23071), .B(new_n23058_1), .Y(new_n23072));
  and_5  g20724(.A(new_n23072), .B(new_n22703), .Y(new_n23073));
  nor_5  g20725(.A(new_n23072), .B(new_n22703), .Y(new_n23074));
  not_8  g20726(.A(new_n22728), .Y(new_n23075));
  nand_5 g20727(.A(new_n23018), .B(new_n23017), .Y(new_n23076));
  xor_4  g20728(.A(new_n23076), .B(new_n23056), .Y(new_n23077));
  or_5   g20729(.A(new_n23077), .B(new_n23075), .Y(new_n23078));
  nand_5 g20730(.A(new_n23077), .B(new_n23075), .Y(new_n23079));
  not_8  g20731(.A(new_n22734), .Y(new_n23080));
  nand_5 g20732(.A(new_n23022), .B(new_n23021), .Y(new_n23081));
  xor_4  g20733(.A(new_n23081), .B(new_n23054), .Y(new_n23082));
  or_5   g20734(.A(new_n23082), .B(new_n23080), .Y(new_n23083));
  nand_5 g20735(.A(new_n23082), .B(new_n23080), .Y(new_n23084));
  nand_5 g20736(.A(new_n23026), .B(new_n23025), .Y(new_n23085));
  xor_4  g20737(.A(new_n23085), .B(new_n23052), .Y(new_n23086));
  or_5   g20738(.A(new_n23086), .B(new_n22741), .Y(new_n23087));
  nand_5 g20739(.A(new_n23086), .B(new_n22741), .Y(new_n23088));
  nand_5 g20740(.A(new_n23030), .B(new_n23029), .Y(new_n23089));
  xor_4  g20741(.A(new_n23089), .B(new_n23050), .Y(new_n23090));
  or_5   g20742(.A(new_n23090), .B(new_n15673), .Y(new_n23091));
  nand_5 g20743(.A(new_n23090), .B(new_n15673), .Y(new_n23092));
  nand_5 g20744(.A(new_n23034), .B(new_n23033), .Y(new_n23093));
  xor_4  g20745(.A(new_n23093), .B(new_n23048), .Y(new_n23094));
  or_5   g20746(.A(new_n23094), .B(new_n15631), .Y(new_n23095));
  nand_5 g20747(.A(new_n23094), .B(new_n15631), .Y(new_n23096));
  not_8  g20748(.A(new_n15637), .Y(new_n23097));
  nand_5 g20749(.A(new_n23038), .B(new_n23037), .Y(new_n23098));
  xor_4  g20750(.A(new_n23098), .B(new_n23046), .Y(new_n23099));
  or_5   g20751(.A(new_n23099), .B(new_n23097), .Y(new_n23100));
  nand_5 g20752(.A(new_n23099), .B(new_n23097), .Y(new_n23101));
  not_8  g20753(.A(new_n15643), .Y(new_n23102));
  nand_5 g20754(.A(new_n23042), .B(new_n23041), .Y(new_n23103));
  xor_4  g20755(.A(new_n23103), .B(new_n23044), .Y(new_n23104));
  or_5   g20756(.A(new_n23104), .B(new_n23102), .Y(new_n23105));
  nand_5 g20757(.A(new_n23104), .B(new_n23102), .Y(new_n23106));
  nand_5 g20758(.A(new_n17871), .B(new_n17860), .Y(new_n23107));
  nand_5 g20759(.A(new_n23107), .B(new_n17870), .Y(new_n23108));
  nand_5 g20760(.A(new_n23108), .B(new_n23106), .Y(new_n23109));
  nand_5 g20761(.A(new_n23109), .B(new_n23105), .Y(new_n23110));
  nand_5 g20762(.A(new_n23110), .B(new_n23101), .Y(new_n23111));
  nand_5 g20763(.A(new_n23111), .B(new_n23100), .Y(new_n23112));
  nand_5 g20764(.A(new_n23112), .B(new_n23096), .Y(new_n23113));
  nand_5 g20765(.A(new_n23113), .B(new_n23095), .Y(new_n23114));
  nand_5 g20766(.A(new_n23114), .B(new_n23092), .Y(new_n23115));
  nand_5 g20767(.A(new_n23115), .B(new_n23091), .Y(new_n23116));
  nand_5 g20768(.A(new_n23116), .B(new_n23088), .Y(new_n23117));
  nand_5 g20769(.A(new_n23117), .B(new_n23087), .Y(new_n23118));
  nand_5 g20770(.A(new_n23118), .B(new_n23084), .Y(new_n23119));
  nand_5 g20771(.A(new_n23119), .B(new_n23083), .Y(new_n23120_1));
  nand_5 g20772(.A(new_n23120_1), .B(new_n23079), .Y(new_n23121));
  nand_5 g20773(.A(new_n23121), .B(new_n23078), .Y(new_n23122));
  nor_5  g20774(.A(new_n23122), .B(new_n23074), .Y(new_n23123));
  nor_5  g20775(.A(new_n23123), .B(new_n23073), .Y(new_n23124));
  xor_4  g20776(.A(new_n23124), .B(new_n23070), .Y(n6707));
  xor_4  g20777(.A(new_n14962), .B(new_n14693), .Y(n6736));
  or_5   g20778(.A(new_n20505), .B(n13490), .Y(new_n23127));
  nor_5  g20779(.A(new_n23127), .B(n9655), .Y(new_n23128));
  nand_5 g20780(.A(new_n23128), .B(new_n6238), .Y(new_n23129));
  nor_5  g20781(.A(new_n23129), .B(n13494), .Y(new_n23130));
  not_8  g20782(.A(new_n23130), .Y(new_n23131));
  nand_5 g20783(.A(new_n23129), .B(n13494), .Y(new_n23132));
  nand_5 g20784(.A(new_n23132), .B(new_n23131), .Y(new_n23133));
  nand_5 g20785(.A(new_n23133), .B(n12650), .Y(new_n23134));
  or_5   g20786(.A(new_n23133), .B(n12650), .Y(new_n23135));
  nand_5 g20787(.A(new_n23135), .B(new_n23134), .Y(new_n23136));
  xor_4  g20788(.A(new_n23128), .B(n25345), .Y(new_n23137));
  or_5   g20789(.A(new_n23137), .B(n10201), .Y(new_n23138));
  nand_5 g20790(.A(new_n23137), .B(n10201), .Y(new_n23139));
  xor_4  g20791(.A(new_n23127), .B(new_n6242), .Y(new_n23140));
  or_5   g20792(.A(new_n23140), .B(n10593), .Y(new_n23141));
  nand_5 g20793(.A(new_n23140), .B(n10593), .Y(new_n23142));
  nand_5 g20794(.A(new_n20505), .B(n13490), .Y(new_n23143));
  nand_5 g20795(.A(new_n23143), .B(new_n23127), .Y(new_n23144));
  or_5   g20796(.A(new_n23144), .B(n18290), .Y(new_n23145));
  nand_5 g20797(.A(new_n23144), .B(n18290), .Y(new_n23146_1));
  nand_5 g20798(.A(new_n20509), .B(new_n20502), .Y(new_n23147));
  nand_5 g20799(.A(new_n23147), .B(new_n20508), .Y(new_n23148));
  nand_5 g20800(.A(new_n23148), .B(new_n23146_1), .Y(new_n23149));
  nand_5 g20801(.A(new_n23149), .B(new_n23145), .Y(new_n23150));
  nand_5 g20802(.A(new_n23150), .B(new_n23142), .Y(new_n23151));
  nand_5 g20803(.A(new_n23151), .B(new_n23141), .Y(new_n23152));
  nand_5 g20804(.A(new_n23152), .B(new_n23139), .Y(new_n23153));
  nand_5 g20805(.A(new_n23153), .B(new_n23138), .Y(new_n23154));
  xor_4  g20806(.A(new_n23154), .B(new_n23136), .Y(new_n23155));
  nand_5 g20807(.A(new_n23155), .B(new_n18122), .Y(new_n23156));
  or_5   g20808(.A(new_n23155), .B(new_n18122), .Y(new_n23157));
  nand_5 g20809(.A(new_n23157), .B(new_n23156), .Y(new_n23158));
  nand_5 g20810(.A(new_n23139), .B(new_n23138), .Y(new_n23159));
  xor_4  g20811(.A(new_n23159), .B(new_n23152), .Y(new_n23160_1));
  nand_5 g20812(.A(new_n23160_1), .B(new_n18131), .Y(new_n23161));
  or_5   g20813(.A(new_n23160_1), .B(new_n18131), .Y(new_n23162));
  nand_5 g20814(.A(new_n23142), .B(new_n23141), .Y(new_n23163));
  xor_4  g20815(.A(new_n23163), .B(new_n23150), .Y(new_n23164));
  nand_5 g20816(.A(new_n23164), .B(new_n18137), .Y(new_n23165));
  or_5   g20817(.A(new_n23164), .B(new_n18137), .Y(new_n23166_1));
  nand_5 g20818(.A(new_n23146_1), .B(new_n23145), .Y(new_n23167));
  xor_4  g20819(.A(new_n23167), .B(new_n23148), .Y(new_n23168));
  nand_5 g20820(.A(new_n23168), .B(new_n18142), .Y(new_n23169));
  or_5   g20821(.A(new_n23168), .B(new_n18142), .Y(new_n23170));
  nand_5 g20822(.A(new_n20513), .B(new_n20500), .Y(new_n23171));
  nand_5 g20823(.A(new_n23171), .B(new_n20512), .Y(new_n23172));
  nand_5 g20824(.A(new_n23172), .B(new_n23170), .Y(new_n23173));
  nand_5 g20825(.A(new_n23173), .B(new_n23169), .Y(new_n23174));
  nand_5 g20826(.A(new_n23174), .B(new_n23166_1), .Y(new_n23175));
  nand_5 g20827(.A(new_n23175), .B(new_n23165), .Y(new_n23176));
  nand_5 g20828(.A(new_n23176), .B(new_n23162), .Y(new_n23177));
  nand_5 g20829(.A(new_n23177), .B(new_n23161), .Y(new_n23178));
  xor_4  g20830(.A(new_n23178), .B(new_n23158), .Y(new_n23179));
  nand_5 g20831(.A(new_n6384), .B(n5101), .Y(new_n23180));
  nand_5 g20832(.A(n23895), .B(new_n3541_1), .Y(new_n23181));
  nand_5 g20833(.A(new_n23181), .B(new_n23180), .Y(new_n23182));
  nand_5 g20834(.A(new_n6388), .B(n16507), .Y(new_n23183));
  nand_5 g20835(.A(n17351), .B(new_n3587), .Y(new_n23184));
  nand_5 g20836(.A(n22470), .B(new_n6392), .Y(new_n23185));
  nand_5 g20837(.A(new_n3613), .B(n11736), .Y(new_n23186));
  nand_5 g20838(.A(new_n6396), .B(n19116), .Y(new_n23187));
  nand_5 g20839(.A(n23200), .B(new_n3577), .Y(new_n23188));
  nand_5 g20840(.A(new_n20519), .B(new_n20517), .Y(new_n23189));
  nand_5 g20841(.A(new_n23189), .B(new_n20518), .Y(new_n23190));
  nand_5 g20842(.A(new_n23190), .B(new_n23188), .Y(new_n23191));
  nand_5 g20843(.A(new_n23191), .B(new_n23187), .Y(new_n23192));
  nand_5 g20844(.A(new_n23192), .B(new_n23186), .Y(new_n23193));
  nand_5 g20845(.A(new_n23193), .B(new_n23185), .Y(new_n23194));
  nand_5 g20846(.A(new_n23194), .B(new_n23184), .Y(new_n23195));
  nand_5 g20847(.A(new_n23195), .B(new_n23183), .Y(new_n23196));
  xnor_4 g20848(.A(new_n23196), .B(new_n23182), .Y(new_n23197));
  nand_5 g20849(.A(new_n23197), .B(new_n23179), .Y(new_n23198));
  or_5   g20850(.A(new_n23197), .B(new_n23179), .Y(new_n23199));
  nand_5 g20851(.A(new_n23199), .B(new_n23198), .Y(new_n23200_1));
  nand_5 g20852(.A(new_n23184), .B(new_n23183), .Y(new_n23201));
  xor_4  g20853(.A(new_n23201), .B(new_n23194), .Y(new_n23202));
  nand_5 g20854(.A(new_n23162), .B(new_n23161), .Y(new_n23203));
  xor_4  g20855(.A(new_n23203), .B(new_n23176), .Y(new_n23204));
  not_8  g20856(.A(new_n23204), .Y(new_n23205));
  or_5   g20857(.A(new_n23205), .B(new_n23202), .Y(new_n23206));
  nand_5 g20858(.A(new_n23205), .B(new_n23202), .Y(new_n23207));
  nand_5 g20859(.A(new_n23186), .B(new_n23185), .Y(new_n23208));
  xor_4  g20860(.A(new_n23208), .B(new_n23192), .Y(new_n23209));
  nand_5 g20861(.A(new_n23166_1), .B(new_n23165), .Y(new_n23210));
  xor_4  g20862(.A(new_n23210), .B(new_n23174), .Y(new_n23211));
  not_8  g20863(.A(new_n23211), .Y(new_n23212));
  or_5   g20864(.A(new_n23212), .B(new_n23209), .Y(new_n23213));
  nand_5 g20865(.A(new_n23212), .B(new_n23209), .Y(new_n23214));
  nand_5 g20866(.A(new_n23188), .B(new_n23187), .Y(new_n23215));
  xor_4  g20867(.A(new_n23215), .B(new_n23190), .Y(new_n23216));
  nand_5 g20868(.A(new_n23170), .B(new_n23169), .Y(new_n23217));
  xor_4  g20869(.A(new_n23217), .B(new_n23172), .Y(new_n23218));
  not_8  g20870(.A(new_n23218), .Y(new_n23219));
  or_5   g20871(.A(new_n23219), .B(new_n23216), .Y(new_n23220));
  nand_5 g20872(.A(new_n23219), .B(new_n23216), .Y(new_n23221));
  nand_5 g20873(.A(new_n20523), .B(new_n20498), .Y(new_n23222));
  nand_5 g20874(.A(new_n23222), .B(new_n20522), .Y(new_n23223));
  nand_5 g20875(.A(new_n23223), .B(new_n23221), .Y(new_n23224));
  nand_5 g20876(.A(new_n23224), .B(new_n23220), .Y(new_n23225));
  nand_5 g20877(.A(new_n23225), .B(new_n23214), .Y(new_n23226));
  nand_5 g20878(.A(new_n23226), .B(new_n23213), .Y(new_n23227));
  nand_5 g20879(.A(new_n23227), .B(new_n23207), .Y(new_n23228));
  nand_5 g20880(.A(new_n23228), .B(new_n23206), .Y(new_n23229));
  xnor_4 g20881(.A(new_n23229), .B(new_n23200_1), .Y(n6791));
  nand_5 g20882(.A(new_n4034), .B(new_n4033), .Y(new_n23231));
  xnor_4 g20883(.A(new_n23231), .B(new_n4048), .Y(n6802));
  nand_5 g20884(.A(new_n18513_1), .B(new_n18512), .Y(new_n23233));
  xnor_4 g20885(.A(new_n23233), .B(new_n18545), .Y(n6826));
  nand_5 g20886(.A(new_n11574), .B(new_n11573), .Y(new_n23235));
  xor_4  g20887(.A(new_n23235), .B(new_n11607_1), .Y(n6835));
  nand_5 g20888(.A(new_n20735), .B(new_n11623), .Y(new_n23237));
  nand_5 g20889(.A(new_n20737), .B(n11220), .Y(new_n23238_1));
  nand_5 g20890(.A(new_n3291), .B(new_n3276), .Y(new_n23239));
  nand_5 g20891(.A(new_n3302), .B(n22379), .Y(new_n23240));
  nand_5 g20892(.A(new_n3189), .B(new_n3030_1), .Y(new_n23241));
  nand_5 g20893(.A(new_n3202), .B(n1662), .Y(new_n23242));
  nand_5 g20894(.A(new_n3071), .B(new_n2997), .Y(new_n23243));
  nand_5 g20895(.A(new_n3115), .B(n12875), .Y(new_n23244));
  nand_5 g20896(.A(new_n3119), .B(new_n3000), .Y(new_n23245));
  nand_5 g20897(.A(new_n3118), .B(n2035), .Y(new_n23246));
  nand_5 g20898(.A(new_n3127), .B(new_n3004), .Y(new_n23247_1));
  nand_5 g20899(.A(new_n3126_1), .B(n5213), .Y(new_n23248_1));
  nand_5 g20900(.A(new_n3135), .B(new_n3007), .Y(new_n23249));
  nand_5 g20901(.A(new_n3134), .B(n4665), .Y(new_n23250_1));
  nand_5 g20902(.A(new_n3144), .B(new_n3010_1), .Y(new_n23251));
  nand_5 g20903(.A(new_n3143), .B(n19005), .Y(new_n23252));
  nand_5 g20904(.A(new_n6569), .B(new_n3013), .Y(new_n23253));
  or_5   g20905(.A(new_n6569), .B(new_n3013), .Y(new_n23254));
  nand_5 g20906(.A(new_n23254), .B(new_n3152), .Y(new_n23255));
  nand_5 g20907(.A(new_n23255), .B(new_n23253), .Y(new_n23256));
  nand_5 g20908(.A(new_n23256), .B(new_n23252), .Y(new_n23257));
  nand_5 g20909(.A(new_n23257), .B(new_n23251), .Y(new_n23258));
  nand_5 g20910(.A(new_n23258), .B(new_n23250_1), .Y(new_n23259));
  nand_5 g20911(.A(new_n23259), .B(new_n23249), .Y(new_n23260));
  nand_5 g20912(.A(new_n23260), .B(new_n23248_1), .Y(new_n23261));
  nand_5 g20913(.A(new_n23261), .B(new_n23247_1), .Y(new_n23262));
  nand_5 g20914(.A(new_n23262), .B(new_n23246), .Y(new_n23263));
  nand_5 g20915(.A(new_n23263), .B(new_n23245), .Y(new_n23264));
  nand_5 g20916(.A(new_n23264), .B(new_n23244), .Y(new_n23265));
  nand_5 g20917(.A(new_n23265), .B(new_n23243), .Y(new_n23266));
  nand_5 g20918(.A(new_n23266), .B(new_n23242), .Y(new_n23267));
  nand_5 g20919(.A(new_n23267), .B(new_n23241), .Y(new_n23268));
  nand_5 g20920(.A(new_n23268), .B(new_n23240), .Y(new_n23269));
  nand_5 g20921(.A(new_n23269), .B(new_n23239), .Y(new_n23270_1));
  nand_5 g20922(.A(new_n23270_1), .B(new_n23238_1), .Y(new_n23271));
  nand_5 g20923(.A(new_n23271), .B(new_n23237), .Y(new_n23272_1));
  nor_5  g20924(.A(new_n23272_1), .B(new_n20730), .Y(new_n23273));
  or_5   g20925(.A(new_n23273), .B(new_n20365), .Y(new_n23274));
  nand_5 g20926(.A(new_n23273), .B(new_n20365), .Y(new_n23275));
  nand_5 g20927(.A(new_n23275), .B(new_n23274), .Y(new_n23276));
  xor_4  g20928(.A(new_n23272_1), .B(new_n20730), .Y(new_n23277));
  and_5  g20929(.A(new_n23277), .B(new_n20371), .Y(new_n23278));
  nor_5  g20930(.A(new_n23277), .B(new_n20371), .Y(new_n23279));
  nand_5 g20931(.A(new_n23237), .B(new_n23238_1), .Y(new_n23280));
  xor_4  g20932(.A(new_n23280), .B(new_n23270_1), .Y(new_n23281));
  nand_5 g20933(.A(new_n23281), .B(new_n14750), .Y(new_n23282));
  not_8  g20934(.A(new_n23282), .Y(new_n23283));
  nor_5  g20935(.A(new_n23281), .B(new_n14750), .Y(new_n23284));
  nand_5 g20936(.A(new_n23239), .B(new_n23240), .Y(new_n23285));
  xor_4  g20937(.A(new_n23285), .B(new_n23268), .Y(new_n23286));
  nand_5 g20938(.A(new_n23286), .B(new_n14754), .Y(new_n23287));
  not_8  g20939(.A(new_n23287), .Y(new_n23288));
  nor_5  g20940(.A(new_n23286), .B(new_n14754), .Y(new_n23289_1));
  not_8  g20941(.A(new_n6923), .Y(new_n23290));
  nand_5 g20942(.A(new_n23241), .B(new_n23242), .Y(new_n23291));
  xor_4  g20943(.A(new_n23291), .B(new_n23266), .Y(new_n23292));
  nand_5 g20944(.A(new_n23292), .B(new_n23290), .Y(new_n23293));
  not_8  g20945(.A(new_n23293), .Y(new_n23294));
  nor_5  g20946(.A(new_n23292), .B(new_n23290), .Y(new_n23295));
  nand_5 g20947(.A(new_n23243), .B(new_n23244), .Y(new_n23296));
  xor_4  g20948(.A(new_n23296), .B(new_n23264), .Y(new_n23297));
  or_5   g20949(.A(new_n23297), .B(new_n14762), .Y(new_n23298));
  nand_5 g20950(.A(new_n23297), .B(new_n14762), .Y(new_n23299));
  nand_5 g20951(.A(new_n23245), .B(new_n23246), .Y(new_n23300));
  xor_4  g20952(.A(new_n23300), .B(new_n23262), .Y(new_n23301));
  or_5   g20953(.A(new_n23301), .B(new_n14765), .Y(new_n23302));
  nand_5 g20954(.A(new_n23301), .B(new_n14765), .Y(new_n23303));
  nand_5 g20955(.A(new_n23247_1), .B(new_n23248_1), .Y(new_n23304_1));
  xor_4  g20956(.A(new_n23304_1), .B(new_n23260), .Y(new_n23305_1));
  or_5   g20957(.A(new_n23305_1), .B(new_n14768), .Y(new_n23306));
  nand_5 g20958(.A(new_n23305_1), .B(new_n14768), .Y(new_n23307));
  nand_5 g20959(.A(new_n23249), .B(new_n23250_1), .Y(new_n23308));
  xor_4  g20960(.A(new_n23308), .B(new_n23258), .Y(new_n23309));
  or_5   g20961(.A(new_n23309), .B(new_n14771), .Y(new_n23310));
  not_8  g20962(.A(new_n23310), .Y(new_n23311));
  nand_5 g20963(.A(new_n23309), .B(new_n14771), .Y(new_n23312));
  not_8  g20964(.A(new_n23312), .Y(new_n23313));
  nand_5 g20965(.A(new_n23251), .B(new_n23252), .Y(new_n23314));
  xor_4  g20966(.A(new_n23314), .B(new_n23256), .Y(new_n23315));
  nand_5 g20967(.A(new_n23315), .B(new_n14774), .Y(new_n23316));
  or_5   g20968(.A(new_n23315), .B(new_n14774), .Y(new_n23317));
  nand_5 g20969(.A(new_n23253), .B(new_n23254), .Y(new_n23318));
  xor_4  g20970(.A(new_n23318), .B(new_n3151), .Y(new_n23319));
  or_5   g20971(.A(new_n23319), .B(new_n6962), .Y(new_n23320));
  nand_5 g20972(.A(new_n6571), .B(new_n6567_1), .Y(new_n23321));
  nand_5 g20973(.A(new_n23319), .B(new_n6962), .Y(new_n23322));
  nand_5 g20974(.A(new_n23322), .B(new_n23321), .Y(new_n23323));
  nand_5 g20975(.A(new_n23323), .B(new_n23320), .Y(new_n23324));
  nand_5 g20976(.A(new_n23324), .B(new_n23317), .Y(new_n23325));
  nand_5 g20977(.A(new_n23325), .B(new_n23316), .Y(new_n23326));
  nor_5  g20978(.A(new_n23326), .B(new_n23313), .Y(new_n23327));
  nor_5  g20979(.A(new_n23327), .B(new_n23311), .Y(new_n23328));
  not_8  g20980(.A(new_n23328), .Y(new_n23329));
  nand_5 g20981(.A(new_n23329), .B(new_n23307), .Y(new_n23330));
  nand_5 g20982(.A(new_n23330), .B(new_n23306), .Y(new_n23331));
  nand_5 g20983(.A(new_n23331), .B(new_n23303), .Y(new_n23332));
  nand_5 g20984(.A(new_n23332), .B(new_n23302), .Y(new_n23333_1));
  nand_5 g20985(.A(new_n23333_1), .B(new_n23299), .Y(new_n23334));
  nand_5 g20986(.A(new_n23334), .B(new_n23298), .Y(new_n23335));
  nor_5  g20987(.A(new_n23335), .B(new_n23295), .Y(new_n23336));
  nor_5  g20988(.A(new_n23336), .B(new_n23294), .Y(new_n23337));
  nor_5  g20989(.A(new_n23337), .B(new_n23289_1), .Y(new_n23338));
  nor_5  g20990(.A(new_n23338), .B(new_n23288), .Y(new_n23339));
  nor_5  g20991(.A(new_n23339), .B(new_n23284), .Y(new_n23340));
  nor_5  g20992(.A(new_n23340), .B(new_n23283), .Y(new_n23341_1));
  nor_5  g20993(.A(new_n23341_1), .B(new_n23279), .Y(new_n23342_1));
  nor_5  g20994(.A(new_n23342_1), .B(new_n23278), .Y(new_n23343));
  xor_4  g20995(.A(new_n23343), .B(new_n23276), .Y(n6853));
  nand_5 g20996(.A(new_n16983), .B(new_n12845), .Y(new_n23345));
  or_5   g20997(.A(new_n16983), .B(new_n12845), .Y(new_n23346));
  nand_5 g20998(.A(new_n14818), .B(new_n14816), .Y(new_n23347));
  nand_5 g20999(.A(new_n23347), .B(new_n14817), .Y(new_n23348));
  nand_5 g21000(.A(new_n23348), .B(new_n23346), .Y(new_n23349));
  nand_5 g21001(.A(new_n23349), .B(new_n23345), .Y(new_n23350));
  nand_5 g21002(.A(new_n16976), .B(new_n12840), .Y(new_n23351));
  nand_5 g21003(.A(new_n16977), .B(new_n12841), .Y(new_n23352));
  nand_5 g21004(.A(new_n23352), .B(new_n23351), .Y(new_n23353));
  xnor_4 g21005(.A(new_n23353), .B(new_n23350), .Y(n6862));
  not_8  g21006(.A(new_n18098), .Y(new_n23355_1));
  nor_5  g21007(.A(new_n23355_1), .B(new_n18075), .Y(new_n23356));
  nor_5  g21008(.A(new_n23356), .B(new_n18074), .Y(new_n23357));
  not_8  g21009(.A(new_n23357), .Y(new_n23358));
  nand_5 g21010(.A(new_n13014), .B(new_n12999), .Y(new_n23359));
  nand_5 g21011(.A(new_n23359), .B(new_n13000), .Y(new_n23360));
  not_8  g21012(.A(new_n23360), .Y(new_n23361));
  nand_5 g21013(.A(new_n23361), .B(new_n20930), .Y(new_n23362));
  nand_5 g21014(.A(new_n23360), .B(new_n20929_1), .Y(new_n23363));
  nand_5 g21015(.A(new_n13048_1), .B(new_n13017), .Y(new_n23364));
  nand_5 g21016(.A(new_n23364), .B(new_n13020), .Y(new_n23365));
  nand_5 g21017(.A(new_n23365), .B(new_n23363), .Y(new_n23366));
  nand_5 g21018(.A(new_n23366), .B(new_n23362), .Y(new_n23367));
  nor_5  g21019(.A(new_n23367), .B(new_n23358), .Y(new_n23368));
  nand_5 g21020(.A(new_n18071_1), .B(new_n18056), .Y(new_n23369_1));
  nand_5 g21021(.A(new_n23369_1), .B(new_n18055), .Y(new_n23370));
  and_5  g21022(.A(new_n23370), .B(new_n23367), .Y(new_n23371_1));
  nor_5  g21023(.A(new_n23371_1), .B(new_n23368), .Y(new_n23372));
  nand_5 g21024(.A(new_n23362), .B(new_n23363), .Y(new_n23373));
  xor_4  g21025(.A(new_n23373), .B(new_n23365), .Y(new_n23374));
  not_8  g21026(.A(new_n23374), .Y(new_n23375));
  nand_5 g21027(.A(new_n23375), .B(new_n23370), .Y(new_n23376));
  nand_5 g21028(.A(new_n23374), .B(new_n23357), .Y(new_n23377));
  nand_5 g21029(.A(new_n23377), .B(new_n23376), .Y(new_n23378));
  nor_5  g21030(.A(new_n23378), .B(new_n23372), .Y(n6863));
  nand_5 g21031(.A(new_n6921), .B(new_n6919), .Y(new_n23380));
  xnor_4 g21032(.A(new_n23380), .B(new_n6986), .Y(n6867));
  nand_5 g21033(.A(new_n20303), .B(new_n20304), .Y(new_n23382));
  xor_4  g21034(.A(new_n23382), .B(new_n20310), .Y(n6965));
  nand_5 g21035(.A(new_n8504), .B(new_n8503), .Y(new_n23384));
  xnor_4 g21036(.A(new_n23384), .B(new_n8555), .Y(n6967));
  nor_5  g21037(.A(new_n16370), .B(new_n16368), .Y(new_n23386));
  xor_4  g21038(.A(new_n23386), .B(new_n16435), .Y(n6975));
  nand_5 g21039(.A(new_n22600), .B(new_n22599), .Y(new_n23388));
  xnor_4 g21040(.A(new_n23388), .B(new_n22602), .Y(n6983));
  nand_5 g21041(.A(new_n16949), .B(new_n12820), .Y(new_n23390));
  nand_5 g21042(.A(new_n16947), .B(new_n12819), .Y(new_n23391));
  nand_5 g21043(.A(new_n23391), .B(new_n23390), .Y(new_n23392));
  nand_5 g21044(.A(new_n16956), .B(new_n12826), .Y(new_n23393));
  nand_5 g21045(.A(new_n16955), .B(new_n12825), .Y(new_n23394));
  nand_5 g21046(.A(new_n16962), .B(new_n12831), .Y(new_n23395));
  nand_5 g21047(.A(new_n16961), .B(new_n12830), .Y(new_n23396));
  nand_5 g21048(.A(new_n16970), .B(new_n12835), .Y(new_n23397));
  nand_5 g21049(.A(new_n16971_1), .B(new_n12836), .Y(new_n23398));
  nand_5 g21050(.A(new_n23352), .B(new_n23350), .Y(new_n23399));
  nand_5 g21051(.A(new_n23399), .B(new_n23351), .Y(new_n23400));
  nand_5 g21052(.A(new_n23400), .B(new_n23398), .Y(new_n23401_1));
  and_5  g21053(.A(new_n23401_1), .B(new_n23397), .Y(new_n23402));
  nand_5 g21054(.A(new_n23402), .B(new_n23396), .Y(new_n23403));
  nand_5 g21055(.A(new_n23403), .B(new_n23395), .Y(new_n23404));
  nand_5 g21056(.A(new_n23404), .B(new_n23394), .Y(new_n23405));
  nand_5 g21057(.A(new_n23405), .B(new_n23393), .Y(new_n23406));
  xor_4  g21058(.A(new_n23406), .B(new_n23392), .Y(n6985));
  nand_5 g21059(.A(new_n16702), .B(new_n16701), .Y(new_n23408));
  xor_4  g21060(.A(new_n23408), .B(new_n16758), .Y(n6998));
  xor_4  g21061(.A(new_n12794), .B(new_n10224), .Y(n7032));
  nand_5 g21062(.A(new_n22409), .B(new_n22410), .Y(new_n23411));
  xnor_4 g21063(.A(new_n23411), .B(new_n22452), .Y(n7038));
  nand_5 g21064(.A(new_n20100), .B(new_n20099), .Y(new_n23413));
  xor_4  g21065(.A(new_n23413), .B(new_n20101), .Y(n7079));
  nor_5  g21066(.A(new_n8544), .B(new_n8541), .Y(new_n23415));
  xor_4  g21067(.A(new_n23415), .B(new_n19129), .Y(n7190));
  nand_5 g21068(.A(new_n18015), .B(new_n18014), .Y(new_n23417));
  xnor_4 g21069(.A(new_n23417), .B(new_n18017), .Y(n7229));
  nand_5 g21070(.A(new_n9801), .B(new_n9802), .Y(new_n23419));
  xnor_4 g21071(.A(new_n23419), .B(new_n9816), .Y(n7230));
  nand_5 g21072(.A(new_n21587), .B(new_n21588), .Y(new_n23421));
  xor_4  g21073(.A(new_n23421), .B(new_n21603), .Y(n7233));
  nand_5 g21074(.A(new_n15086), .B(new_n15085), .Y(new_n23423));
  xor_4  g21075(.A(new_n23423), .B(new_n15094_1), .Y(n7236));
  xor_4  g21076(.A(new_n18408), .B(new_n13537), .Y(n7253));
  nor_5  g21077(.A(new_n22023), .B(n12507), .Y(new_n23426));
  nor_5  g21078(.A(new_n22026), .B(new_n23426), .Y(new_n23427));
  or_5   g21079(.A(new_n22022), .B(n17458), .Y(new_n23428));
  nand_5 g21080(.A(new_n22023), .B(n12507), .Y(new_n23429_1));
  nand_5 g21081(.A(new_n23429_1), .B(new_n23428), .Y(new_n23430_1));
  nor_5  g21082(.A(new_n23430_1), .B(new_n23427), .Y(new_n23431));
  not_8  g21083(.A(new_n23431), .Y(new_n23432));
  or_5   g21084(.A(new_n22621), .B(new_n16064), .Y(new_n23433_1));
  xor_4  g21085(.A(new_n23433_1), .B(new_n16062_1), .Y(new_n23434_1));
  nand_5 g21086(.A(new_n23434_1), .B(new_n11637), .Y(new_n23435));
  nor_5  g21087(.A(new_n23434_1), .B(new_n11637), .Y(new_n23436));
  not_8  g21088(.A(new_n23436), .Y(new_n23437));
  nand_5 g21089(.A(new_n23437), .B(new_n23435), .Y(new_n23438));
  nand_5 g21090(.A(new_n22621), .B(new_n16064), .Y(new_n23439));
  nand_5 g21091(.A(new_n23439), .B(new_n23433_1), .Y(new_n23440));
  or_5   g21092(.A(new_n23440), .B(new_n11647_1), .Y(new_n23441));
  nand_5 g21093(.A(new_n22627), .B(new_n22624), .Y(new_n23442));
  nand_5 g21094(.A(new_n23442), .B(new_n22623_1), .Y(new_n23443));
  nand_5 g21095(.A(new_n23440), .B(new_n11647_1), .Y(new_n23444));
  nand_5 g21096(.A(new_n23444), .B(new_n23443), .Y(new_n23445));
  nand_5 g21097(.A(new_n23445), .B(new_n23441), .Y(new_n23446));
  xor_4  g21098(.A(new_n23446), .B(new_n23438), .Y(new_n23447));
  nand_5 g21099(.A(new_n23447), .B(new_n23432), .Y(new_n23448));
  nand_5 g21100(.A(new_n23444), .B(new_n23441), .Y(new_n23449));
  xor_4  g21101(.A(new_n23449), .B(new_n23443), .Y(new_n23450_1));
  nand_5 g21102(.A(new_n23450_1), .B(new_n22027_1), .Y(new_n23451));
  nand_5 g21103(.A(new_n22630), .B(new_n22617), .Y(new_n23452));
  nand_5 g21104(.A(new_n23452), .B(new_n22629), .Y(new_n23453));
  or_5   g21105(.A(new_n23450_1), .B(new_n22027_1), .Y(new_n23454));
  nand_5 g21106(.A(new_n23454), .B(new_n23453), .Y(new_n23455));
  nand_5 g21107(.A(new_n23455), .B(new_n23451), .Y(new_n23456));
  or_5   g21108(.A(new_n23447), .B(new_n23432), .Y(new_n23457));
  nand_5 g21109(.A(new_n23457), .B(new_n23456), .Y(new_n23458));
  nand_5 g21110(.A(new_n23458), .B(new_n23448), .Y(new_n23459));
  not_8  g21111(.A(new_n16062_1), .Y(new_n23460));
  nor_5  g21112(.A(new_n23433_1), .B(new_n23460), .Y(new_n23461));
  nand_5 g21113(.A(new_n23446), .B(new_n23435), .Y(new_n23462));
  nand_5 g21114(.A(new_n23462), .B(new_n23437), .Y(new_n23463_1));
  nor_5  g21115(.A(new_n23463_1), .B(new_n23461), .Y(new_n23464));
  and_5  g21116(.A(new_n23464), .B(new_n23459), .Y(n24172));
  nor_5  g21117(.A(new_n23464), .B(new_n23459), .Y(new_n23466));
  or_5   g21118(.A(new_n23466), .B(n24172), .Y(n7256));
  nand_5 g21119(.A(new_n22162), .B(new_n22160), .Y(new_n23468));
  nand_5 g21120(.A(new_n23468), .B(new_n22161), .Y(new_n23469));
  or_5   g21121(.A(new_n9151), .B(n2416), .Y(new_n23470));
  nand_5 g21122(.A(new_n9151), .B(n2416), .Y(new_n23471_1));
  nand_5 g21123(.A(new_n23471_1), .B(new_n23470), .Y(new_n23472));
  xor_4  g21124(.A(new_n23472), .B(new_n23469), .Y(new_n23473));
  or_5   g21125(.A(new_n23473), .B(new_n17667), .Y(new_n23474));
  nand_5 g21126(.A(new_n23473), .B(new_n17667), .Y(new_n23475));
  nand_5 g21127(.A(new_n22166), .B(new_n22158), .Y(new_n23476));
  nand_5 g21128(.A(new_n23476), .B(new_n22165), .Y(new_n23477));
  nand_5 g21129(.A(new_n23477), .B(new_n23475), .Y(new_n23478));
  nand_5 g21130(.A(new_n23478), .B(new_n23474), .Y(new_n23479));
  not_8  g21131(.A(new_n17664_1), .Y(new_n23480_1));
  nand_5 g21132(.A(new_n23471_1), .B(new_n23469), .Y(new_n23481));
  nand_5 g21133(.A(new_n23481), .B(new_n23470), .Y(new_n23482));
  nand_5 g21134(.A(new_n23482), .B(new_n23480_1), .Y(new_n23483));
  not_8  g21135(.A(new_n23482), .Y(new_n23484));
  nand_5 g21136(.A(new_n23484), .B(new_n17664_1), .Y(new_n23485));
  nand_5 g21137(.A(new_n23485), .B(new_n23483), .Y(new_n23486));
  xor_4  g21138(.A(new_n23486), .B(new_n23479), .Y(new_n23487));
  not_8  g21139(.A(new_n23487), .Y(new_n23488));
  nand_5 g21140(.A(new_n23488), .B(new_n22260), .Y(new_n23489));
  nand_5 g21141(.A(new_n23487), .B(new_n22259), .Y(new_n23490));
  nand_5 g21142(.A(new_n23490), .B(new_n23489), .Y(new_n23491));
  nand_5 g21143(.A(new_n23475), .B(new_n23474), .Y(new_n23492));
  xor_4  g21144(.A(new_n23492), .B(new_n23477), .Y(new_n23493_1));
  nand_5 g21145(.A(new_n23493_1), .B(new_n22269), .Y(new_n23494));
  or_5   g21146(.A(new_n23493_1), .B(new_n22269), .Y(new_n23495));
  nand_5 g21147(.A(new_n22175), .B(new_n22156), .Y(new_n23496));
  nand_5 g21148(.A(new_n23496), .B(new_n22174), .Y(new_n23497));
  nand_5 g21149(.A(new_n23497), .B(new_n23495), .Y(new_n23498));
  nand_5 g21150(.A(new_n23498), .B(new_n23494), .Y(new_n23499));
  xor_4  g21151(.A(new_n23499), .B(new_n23491), .Y(n7268));
  not_8  g21152(.A(n13026), .Y(new_n23501));
  nor_5  g21153(.A(new_n12639), .B(n2175), .Y(new_n23502));
  nand_5 g21154(.A(new_n23502), .B(new_n23501), .Y(new_n23503));
  nor_5  g21155(.A(new_n23503), .B(n23912), .Y(new_n23504));
  not_8  g21156(.A(new_n23504), .Y(new_n23505));
  nand_5 g21157(.A(new_n23503), .B(n23912), .Y(new_n23506));
  and_5  g21158(.A(new_n23506), .B(new_n23505), .Y(new_n23507));
  not_8  g21159(.A(new_n23507), .Y(new_n23508));
  nand_5 g21160(.A(new_n23508), .B(n10514), .Y(new_n23509));
  xor_4  g21161(.A(new_n23502), .B(new_n23501), .Y(new_n23510));
  nand_5 g21162(.A(new_n23510), .B(new_n13224), .Y(new_n23511));
  not_8  g21163(.A(new_n23510), .Y(new_n23512));
  nand_5 g21164(.A(new_n23512), .B(n18649), .Y(new_n23513_1));
  xor_4  g21165(.A(new_n12639), .B(n2175), .Y(new_n23514));
  nand_5 g21166(.A(new_n23514), .B(new_n13227), .Y(new_n23515));
  not_8  g21167(.A(new_n23514), .Y(new_n23516));
  nand_5 g21168(.A(new_n23516), .B(n6218), .Y(new_n23517));
  nand_5 g21169(.A(new_n12641), .B(new_n12632), .Y(new_n23518));
  nand_5 g21170(.A(new_n12644), .B(n20470), .Y(new_n23519));
  nand_5 g21171(.A(new_n12587_1), .B(new_n12539), .Y(new_n23520));
  nand_5 g21172(.A(new_n12590), .B(n21222), .Y(new_n23521));
  nand_5 g21173(.A(new_n12554), .B(new_n11063_1), .Y(new_n23522));
  nand_5 g21174(.A(new_n12557), .B(n9832), .Y(new_n23523));
  nand_5 g21175(.A(new_n12561), .B(new_n10982), .Y(new_n23524));
  nand_5 g21176(.A(new_n12560), .B(n1558), .Y(new_n23525));
  nand_5 g21177(.A(new_n12565), .B(new_n10969), .Y(new_n23526));
  nand_5 g21178(.A(new_n12568), .B(n21749), .Y(new_n23527));
  nand_5 g21179(.A(new_n12573), .B(new_n10973), .Y(new_n23528));
  nand_5 g21180(.A(new_n12574), .B(n7769), .Y(new_n23529_1));
  nand_5 g21181(.A(n21138), .B(new_n12547), .Y(new_n23530));
  nand_5 g21182(.A(new_n23530), .B(new_n23529_1), .Y(new_n23531));
  nand_5 g21183(.A(new_n23531), .B(new_n23528), .Y(new_n23532));
  nand_5 g21184(.A(new_n23532), .B(new_n23527), .Y(new_n23533));
  nand_5 g21185(.A(new_n23533), .B(new_n23526), .Y(new_n23534));
  nand_5 g21186(.A(new_n23534), .B(new_n23525), .Y(new_n23535));
  nand_5 g21187(.A(new_n23535), .B(new_n23524), .Y(new_n23536));
  nand_5 g21188(.A(new_n23536), .B(new_n23523), .Y(new_n23537));
  nand_5 g21189(.A(new_n23537), .B(new_n23522), .Y(new_n23538));
  nand_5 g21190(.A(new_n23538), .B(new_n23521), .Y(new_n23539));
  nand_5 g21191(.A(new_n23539), .B(new_n23520), .Y(new_n23540));
  nand_5 g21192(.A(new_n23540), .B(new_n23519), .Y(new_n23541_1));
  nand_5 g21193(.A(new_n23541_1), .B(new_n23518), .Y(new_n23542));
  nand_5 g21194(.A(new_n23542), .B(new_n23517), .Y(new_n23543));
  nand_5 g21195(.A(new_n23543), .B(new_n23515), .Y(new_n23544));
  nand_5 g21196(.A(new_n23544), .B(new_n23513_1), .Y(new_n23545));
  nand_5 g21197(.A(new_n23545), .B(new_n23511), .Y(new_n23546_1));
  nand_5 g21198(.A(new_n23546_1), .B(new_n23509), .Y(new_n23547));
  not_8  g21199(.A(new_n23547), .Y(new_n23548));
  nand_5 g21200(.A(new_n23548), .B(new_n23504), .Y(new_n23549));
  not_8  g21201(.A(new_n23549), .Y(new_n23550_1));
  nand_5 g21202(.A(new_n23507), .B(new_n13220), .Y(new_n23551));
  nand_5 g21203(.A(new_n23551), .B(new_n23509), .Y(new_n23552));
  xor_4  g21204(.A(new_n23552), .B(new_n23546_1), .Y(new_n23553));
  nand_5 g21205(.A(new_n23553), .B(n9872), .Y(new_n23554));
  or_5   g21206(.A(new_n23553), .B(n9872), .Y(new_n23555));
  nand_5 g21207(.A(new_n23511), .B(new_n23513_1), .Y(new_n23556));
  xor_4  g21208(.A(new_n23556), .B(new_n23544), .Y(new_n23557));
  nand_5 g21209(.A(new_n23557), .B(n5842), .Y(new_n23558));
  or_5   g21210(.A(new_n23557), .B(n5842), .Y(new_n23559));
  nand_5 g21211(.A(new_n23515), .B(new_n23517), .Y(new_n23560));
  xor_4  g21212(.A(new_n23560), .B(new_n23542), .Y(new_n23561));
  nand_5 g21213(.A(new_n23561), .B(n6379), .Y(new_n23562));
  or_5   g21214(.A(new_n23561), .B(n6379), .Y(new_n23563));
  nand_5 g21215(.A(new_n23518), .B(new_n23519), .Y(new_n23564));
  xor_4  g21216(.A(new_n23564), .B(new_n23540), .Y(new_n23565));
  nand_5 g21217(.A(new_n23565), .B(n2102), .Y(new_n23566));
  or_5   g21218(.A(new_n23565), .B(n2102), .Y(new_n23567));
  nand_5 g21219(.A(new_n23520), .B(new_n23521), .Y(new_n23568));
  xor_4  g21220(.A(new_n23568), .B(new_n23538), .Y(new_n23569));
  nand_5 g21221(.A(new_n23569), .B(n17954), .Y(new_n23570));
  or_5   g21222(.A(new_n23569), .B(n17954), .Y(new_n23571));
  nand_5 g21223(.A(new_n23522), .B(new_n23523), .Y(new_n23572));
  xor_4  g21224(.A(new_n23572), .B(new_n23536), .Y(new_n23573));
  nand_5 g21225(.A(new_n23573), .B(n8256), .Y(new_n23574));
  or_5   g21226(.A(new_n23573), .B(n8256), .Y(new_n23575));
  nand_5 g21227(.A(new_n23524), .B(new_n23525), .Y(new_n23576));
  xor_4  g21228(.A(new_n23576), .B(new_n23534), .Y(new_n23577));
  nand_5 g21229(.A(new_n23577), .B(n24150), .Y(new_n23578));
  or_5   g21230(.A(new_n23577), .B(n24150), .Y(new_n23579));
  nand_5 g21231(.A(new_n23526), .B(new_n23527), .Y(new_n23580));
  xor_4  g21232(.A(new_n23580), .B(new_n23532), .Y(new_n23581));
  nand_5 g21233(.A(new_n23581), .B(n19584), .Y(new_n23582));
  or_5   g21234(.A(new_n23581), .B(n19584), .Y(new_n23583));
  nand_5 g21235(.A(new_n23528), .B(new_n23529_1), .Y(new_n23584));
  xor_4  g21236(.A(new_n23584), .B(new_n23530), .Y(new_n23585_1));
  nand_5 g21237(.A(new_n23585_1), .B(n5060), .Y(new_n23586_1));
  or_5   g21238(.A(new_n23585_1), .B(n5060), .Y(new_n23587));
  xor_4  g21239(.A(n21138), .B(new_n12547), .Y(new_n23588_1));
  nand_5 g21240(.A(new_n23588_1), .B(n15332), .Y(new_n23589));
  not_8  g21241(.A(new_n23589), .Y(new_n23590));
  nand_5 g21242(.A(new_n23590), .B(new_n23587), .Y(new_n23591));
  nand_5 g21243(.A(new_n23591), .B(new_n23586_1), .Y(new_n23592));
  nand_5 g21244(.A(new_n23592), .B(new_n23583), .Y(new_n23593));
  nand_5 g21245(.A(new_n23593), .B(new_n23582), .Y(new_n23594));
  nand_5 g21246(.A(new_n23594), .B(new_n23579), .Y(new_n23595));
  nand_5 g21247(.A(new_n23595), .B(new_n23578), .Y(new_n23596));
  nand_5 g21248(.A(new_n23596), .B(new_n23575), .Y(new_n23597));
  nand_5 g21249(.A(new_n23597), .B(new_n23574), .Y(new_n23598));
  nand_5 g21250(.A(new_n23598), .B(new_n23571), .Y(new_n23599));
  nand_5 g21251(.A(new_n23599), .B(new_n23570), .Y(new_n23600));
  nand_5 g21252(.A(new_n23600), .B(new_n23567), .Y(new_n23601));
  nand_5 g21253(.A(new_n23601), .B(new_n23566), .Y(new_n23602));
  nand_5 g21254(.A(new_n23602), .B(new_n23563), .Y(new_n23603));
  nand_5 g21255(.A(new_n23603), .B(new_n23562), .Y(new_n23604));
  nand_5 g21256(.A(new_n23604), .B(new_n23559), .Y(new_n23605));
  nand_5 g21257(.A(new_n23605), .B(new_n23558), .Y(new_n23606));
  nand_5 g21258(.A(new_n23606), .B(new_n23555), .Y(new_n23607));
  nand_5 g21259(.A(new_n23607), .B(new_n23554), .Y(new_n23608));
  not_8  g21260(.A(new_n23608), .Y(new_n23609));
  nand_5 g21261(.A(new_n23609), .B(new_n23550_1), .Y(new_n23610));
  nand_5 g21262(.A(new_n23551), .B(new_n23505), .Y(new_n23611));
  nor_5  g21263(.A(new_n23611), .B(new_n23548), .Y(new_n23612));
  nand_5 g21264(.A(new_n23612), .B(new_n23608), .Y(new_n23613));
  nand_5 g21265(.A(new_n23613), .B(new_n23610), .Y(new_n23614));
  not_8  g21266(.A(new_n23614), .Y(new_n23615));
  nand_5 g21267(.A(new_n23615), .B(new_n16643), .Y(new_n23616));
  nand_5 g21268(.A(new_n23614), .B(new_n16642), .Y(new_n23617));
  nand_5 g21269(.A(new_n23617), .B(new_n23616), .Y(new_n23618));
  nor_5  g21270(.A(new_n23612), .B(new_n23550_1), .Y(new_n23619_1));
  xor_4  g21271(.A(new_n23619_1), .B(new_n23609), .Y(new_n23620));
  nand_5 g21272(.A(new_n23620), .B(new_n16689), .Y(new_n23621));
  or_5   g21273(.A(new_n23620), .B(new_n16689), .Y(new_n23622));
  nand_5 g21274(.A(new_n23554), .B(new_n23555), .Y(new_n23623));
  xor_4  g21275(.A(new_n23623), .B(new_n23606), .Y(new_n23624_1));
  or_5   g21276(.A(new_n23624_1), .B(new_n16694), .Y(new_n23625));
  nand_5 g21277(.A(new_n23624_1), .B(new_n16694), .Y(new_n23626));
  nand_5 g21278(.A(new_n23558), .B(new_n23559), .Y(new_n23627));
  xor_4  g21279(.A(new_n23627), .B(new_n23604), .Y(new_n23628_1));
  or_5   g21280(.A(new_n23628_1), .B(new_n2918), .Y(new_n23629));
  nand_5 g21281(.A(new_n23628_1), .B(new_n2918), .Y(new_n23630));
  nand_5 g21282(.A(new_n23562), .B(new_n23563), .Y(new_n23631));
  xor_4  g21283(.A(new_n23631), .B(new_n23602), .Y(new_n23632));
  or_5   g21284(.A(new_n23632), .B(new_n2925), .Y(new_n23633));
  nand_5 g21285(.A(new_n23632), .B(new_n2925), .Y(new_n23634));
  nand_5 g21286(.A(new_n23566), .B(new_n23567), .Y(new_n23635));
  xor_4  g21287(.A(new_n23635), .B(new_n23600), .Y(new_n23636));
  or_5   g21288(.A(new_n23636), .B(new_n2932), .Y(new_n23637_1));
  nand_5 g21289(.A(new_n23636), .B(new_n2932), .Y(new_n23638));
  nand_5 g21290(.A(new_n23570), .B(new_n23571), .Y(new_n23639));
  xor_4  g21291(.A(new_n23639), .B(new_n23598), .Y(new_n23640));
  or_5   g21292(.A(new_n23640), .B(new_n2939), .Y(new_n23641));
  nand_5 g21293(.A(new_n23640), .B(new_n2939), .Y(new_n23642));
  nand_5 g21294(.A(new_n23574), .B(new_n23575), .Y(new_n23643));
  xor_4  g21295(.A(new_n23643), .B(new_n23596), .Y(new_n23644));
  or_5   g21296(.A(new_n23644), .B(new_n2946), .Y(new_n23645));
  nand_5 g21297(.A(new_n23644), .B(new_n2946), .Y(new_n23646));
  nand_5 g21298(.A(new_n23578), .B(new_n23579), .Y(new_n23647));
  xor_4  g21299(.A(new_n23647), .B(new_n23594), .Y(new_n23648));
  or_5   g21300(.A(new_n23648), .B(new_n2953), .Y(new_n23649));
  nand_5 g21301(.A(new_n23648), .B(new_n2953), .Y(new_n23650));
  nand_5 g21302(.A(new_n23582), .B(new_n23583), .Y(new_n23651));
  xor_4  g21303(.A(new_n23651), .B(new_n23592), .Y(new_n23652));
  or_5   g21304(.A(new_n23652), .B(new_n2960), .Y(new_n23653));
  nand_5 g21305(.A(new_n23652), .B(new_n2960), .Y(new_n23654));
  nand_5 g21306(.A(new_n23586_1), .B(new_n23587), .Y(new_n23655));
  xor_4  g21307(.A(new_n23655), .B(new_n23590), .Y(new_n23656));
  or_5   g21308(.A(new_n23656), .B(new_n2969), .Y(new_n23657_1));
  nand_5 g21309(.A(new_n23656), .B(new_n2969), .Y(new_n23658));
  not_8  g21310(.A(new_n2976), .Y(new_n23659));
  nor_5  g21311(.A(new_n23588_1), .B(n15332), .Y(new_n23660));
  nor_5  g21312(.A(new_n23660), .B(new_n23590), .Y(new_n23661));
  or_5   g21313(.A(new_n23661), .B(new_n23659), .Y(new_n23662));
  nand_5 g21314(.A(new_n23662), .B(new_n23658), .Y(new_n23663_1));
  nand_5 g21315(.A(new_n23663_1), .B(new_n23657_1), .Y(new_n23664));
  nand_5 g21316(.A(new_n23664), .B(new_n23654), .Y(new_n23665));
  nand_5 g21317(.A(new_n23665), .B(new_n23653), .Y(new_n23666));
  nand_5 g21318(.A(new_n23666), .B(new_n23650), .Y(new_n23667));
  nand_5 g21319(.A(new_n23667), .B(new_n23649), .Y(new_n23668));
  nand_5 g21320(.A(new_n23668), .B(new_n23646), .Y(new_n23669_1));
  nand_5 g21321(.A(new_n23669_1), .B(new_n23645), .Y(new_n23670));
  nand_5 g21322(.A(new_n23670), .B(new_n23642), .Y(new_n23671));
  nand_5 g21323(.A(new_n23671), .B(new_n23641), .Y(new_n23672));
  nand_5 g21324(.A(new_n23672), .B(new_n23638), .Y(new_n23673));
  nand_5 g21325(.A(new_n23673), .B(new_n23637_1), .Y(new_n23674));
  nand_5 g21326(.A(new_n23674), .B(new_n23634), .Y(new_n23675));
  nand_5 g21327(.A(new_n23675), .B(new_n23633), .Y(new_n23676));
  nand_5 g21328(.A(new_n23676), .B(new_n23630), .Y(new_n23677));
  nand_5 g21329(.A(new_n23677), .B(new_n23629), .Y(new_n23678));
  nand_5 g21330(.A(new_n23678), .B(new_n23626), .Y(new_n23679));
  nand_5 g21331(.A(new_n23679), .B(new_n23625), .Y(new_n23680));
  nand_5 g21332(.A(new_n23680), .B(new_n23622), .Y(new_n23681));
  nand_5 g21333(.A(new_n23681), .B(new_n23621), .Y(new_n23682));
  xor_4  g21334(.A(new_n23682), .B(new_n23618), .Y(n7277));
  nand_5 g21335(.A(new_n15258_1), .B(new_n15259), .Y(new_n23684_1));
  xor_4  g21336(.A(new_n23684_1), .B(new_n15268), .Y(n7280));
  nand_5 g21337(.A(new_n6469), .B(new_n6468), .Y(new_n23686));
  xnor_4 g21338(.A(new_n23686), .B(new_n6501), .Y(n7298));
  nand_5 g21339(.A(new_n21996), .B(new_n21995), .Y(new_n23688));
  xor_4  g21340(.A(new_n23688), .B(new_n22007), .Y(n7308));
  nand_5 g21341(.A(new_n22266), .B(new_n8333), .Y(new_n23690_1));
  nand_5 g21342(.A(new_n22267), .B(new_n8334), .Y(new_n23691));
  nand_5 g21343(.A(new_n23691), .B(new_n23690_1), .Y(new_n23692));
  nand_5 g21344(.A(new_n22272), .B(new_n8356), .Y(new_n23693));
  nand_5 g21345(.A(new_n22273), .B(new_n8360), .Y(new_n23694));
  nand_5 g21346(.A(new_n17116), .B(new_n17104_1), .Y(new_n23695));
  nand_5 g21347(.A(new_n23695), .B(new_n17114), .Y(new_n23696));
  nand_5 g21348(.A(new_n23696), .B(new_n23694), .Y(new_n23697_1));
  nand_5 g21349(.A(new_n23697_1), .B(new_n23693), .Y(new_n23698));
  not_8  g21350(.A(new_n23698), .Y(new_n23699));
  nor_5  g21351(.A(new_n23699), .B(new_n23692), .Y(new_n23700));
  not_8  g21352(.A(new_n23700), .Y(new_n23701));
  nand_5 g21353(.A(new_n23699), .B(new_n23692), .Y(new_n23702));
  and_5  g21354(.A(new_n23702), .B(new_n23701), .Y(new_n23703));
  not_8  g21355(.A(new_n23703), .Y(new_n23704));
  nand_5 g21356(.A(new_n23704), .B(new_n22300), .Y(new_n23705));
  nand_5 g21357(.A(new_n23703), .B(new_n22295), .Y(new_n23706));
  nand_5 g21358(.A(new_n23706), .B(new_n23705), .Y(new_n23707));
  nand_5 g21359(.A(new_n23693), .B(new_n23694), .Y(new_n23708));
  xor_4  g21360(.A(new_n23708), .B(new_n23696), .Y(new_n23709));
  not_8  g21361(.A(new_n23709), .Y(new_n23710));
  nand_5 g21362(.A(new_n23710), .B(new_n22306), .Y(new_n23711));
  nand_5 g21363(.A(new_n23709), .B(new_n22309_1), .Y(new_n23712));
  nand_5 g21364(.A(new_n21621), .B(new_n21611), .Y(new_n23713));
  nand_5 g21365(.A(new_n23713), .B(new_n21620), .Y(new_n23714_1));
  nand_5 g21366(.A(new_n23714_1), .B(new_n23712), .Y(new_n23715));
  nand_5 g21367(.A(new_n23715), .B(new_n23711), .Y(new_n23716));
  xor_4  g21368(.A(new_n23716), .B(new_n23707), .Y(n7313));
  nand_5 g21369(.A(new_n4020), .B(new_n4019), .Y(new_n23718));
  xnor_4 g21370(.A(new_n23718), .B(new_n4052), .Y(n7346));
  xor_4  g21371(.A(new_n23360), .B(new_n15930), .Y(new_n23720));
  nand_5 g21372(.A(new_n23360), .B(new_n15963), .Y(new_n23721));
  nand_5 g21373(.A(new_n23361), .B(new_n15962), .Y(new_n23722));
  nand_5 g21374(.A(new_n15969), .B(new_n13019), .Y(new_n23723));
  or_5   g21375(.A(new_n15969), .B(new_n13019), .Y(new_n23724));
  nand_5 g21376(.A(new_n15976), .B(new_n13025), .Y(new_n23725));
  or_5   g21377(.A(new_n15976), .B(new_n13025), .Y(new_n23726));
  nand_5 g21378(.A(new_n15981), .B(new_n13033), .Y(new_n23727));
  or_5   g21379(.A(new_n15981), .B(new_n13033), .Y(new_n23728));
  nand_5 g21380(.A(new_n7507_1), .B(new_n7465), .Y(new_n23729));
  nand_5 g21381(.A(new_n23729), .B(new_n7506), .Y(new_n23730));
  nand_5 g21382(.A(new_n23730), .B(new_n23728), .Y(new_n23731));
  nand_5 g21383(.A(new_n23731), .B(new_n23727), .Y(new_n23732));
  nand_5 g21384(.A(new_n23732), .B(new_n23726), .Y(new_n23733));
  nand_5 g21385(.A(new_n23733), .B(new_n23725), .Y(new_n23734));
  nand_5 g21386(.A(new_n23734), .B(new_n23724), .Y(new_n23735));
  nand_5 g21387(.A(new_n23735), .B(new_n23723), .Y(new_n23736));
  nand_5 g21388(.A(new_n23736), .B(new_n23722), .Y(new_n23737));
  nand_5 g21389(.A(new_n23737), .B(new_n23721), .Y(new_n23738));
  xor_4  g21390(.A(new_n23738), .B(new_n23720), .Y(n7349));
  nand_5 g21391(.A(new_n23626), .B(new_n23625), .Y(new_n23740));
  xor_4  g21392(.A(new_n23740), .B(new_n23678), .Y(n7363));
  nand_5 g21393(.A(new_n22242), .B(new_n22239), .Y(new_n23742));
  nand_5 g21394(.A(new_n23742), .B(new_n22238), .Y(new_n23743));
  not_8  g21395(.A(new_n23743), .Y(new_n23744));
  nand_5 g21396(.A(new_n23744), .B(new_n11692), .Y(new_n23745));
  nand_5 g21397(.A(new_n23743), .B(new_n11693), .Y(new_n23746));
  nand_5 g21398(.A(new_n23746), .B(new_n23745), .Y(new_n23747));
  nor_5  g21399(.A(new_n22250), .B(new_n22246), .Y(new_n23748_1));
  nor_5  g21400(.A(new_n23748_1), .B(new_n22245), .Y(new_n23749));
  xor_4  g21401(.A(new_n23749), .B(new_n23747), .Y(n7390));
  nand_5 g21402(.A(new_n10412), .B(new_n10411_1), .Y(new_n23751));
  xor_4  g21403(.A(new_n23751), .B(new_n10438), .Y(n7403));
  nand_5 g21404(.A(new_n10594), .B(new_n10592), .Y(new_n23753));
  xnor_4 g21405(.A(new_n23753), .B(new_n10645), .Y(n7408));
  nand_5 g21406(.A(new_n22582), .B(new_n22581), .Y(new_n23755_1));
  xor_4  g21407(.A(new_n23755_1), .B(new_n22611), .Y(n7432));
  nand_5 g21408(.A(new_n20377), .B(new_n20367), .Y(new_n23757));
  nand_5 g21409(.A(new_n23757), .B(new_n20366_1), .Y(n7475));
  nor_5  g21410(.A(new_n5849), .B(new_n5845), .Y(new_n23759));
  xor_4  g21411(.A(new_n23759), .B(new_n5847), .Y(n7477));
  nor_5  g21412(.A(new_n10207), .B(new_n10206), .Y(new_n23761));
  xor_4  g21413(.A(new_n23761), .B(new_n10240), .Y(n7507));
  not_8  g21414(.A(new_n19638), .Y(new_n23763));
  nand_5 g21415(.A(new_n13751), .B(n23895), .Y(new_n23764));
  nand_5 g21416(.A(new_n13750), .B(new_n6384), .Y(new_n23765));
  nand_5 g21417(.A(new_n7981), .B(new_n7970), .Y(new_n23766));
  nand_5 g21418(.A(new_n23766), .B(new_n7980), .Y(new_n23767));
  nand_5 g21419(.A(new_n23767), .B(new_n23765), .Y(new_n23768));
  nand_5 g21420(.A(new_n23768), .B(new_n23764), .Y(new_n23769));
  xor_4  g21421(.A(new_n23769), .B(new_n13748), .Y(new_n23770));
  nand_5 g21422(.A(new_n23770), .B(new_n23763), .Y(new_n23771));
  or_5   g21423(.A(new_n23770), .B(new_n23763), .Y(new_n23772));
  nand_5 g21424(.A(new_n23772), .B(new_n23771), .Y(new_n23773));
  nand_5 g21425(.A(new_n23764), .B(new_n23765), .Y(new_n23774));
  xor_4  g21426(.A(new_n23774), .B(new_n23767), .Y(new_n23775_1));
  or_5   g21427(.A(new_n23775_1), .B(new_n19647), .Y(new_n23776));
  nand_5 g21428(.A(new_n23775_1), .B(new_n19647), .Y(new_n23777));
  nor_5  g21429(.A(new_n7987), .B(new_n7952), .Y(new_n23778));
  nor_5  g21430(.A(new_n23778), .B(new_n7985), .Y(new_n23779));
  nand_5 g21431(.A(new_n23779), .B(new_n23777), .Y(new_n23780));
  nand_5 g21432(.A(new_n23780), .B(new_n23776), .Y(new_n23781));
  xnor_4 g21433(.A(new_n23781), .B(new_n23773), .Y(n7514));
  nand_5 g21434(.A(new_n12485), .B(new_n12484), .Y(new_n23783));
  xor_4  g21435(.A(new_n23783), .B(new_n12515_1), .Y(n7558));
  nand_5 g21436(.A(new_n13832), .B(new_n13831), .Y(new_n23785));
  xor_4  g21437(.A(new_n23785), .B(new_n13835_1), .Y(n7572));
  nand_5 g21438(.A(new_n22673), .B(new_n22665), .Y(new_n23787));
  nand_5 g21439(.A(new_n23787), .B(new_n22672), .Y(new_n23788));
  nand_5 g21440(.A(new_n22669), .B(new_n22667), .Y(new_n23789));
  nand_5 g21441(.A(new_n23789), .B(new_n22668), .Y(new_n23790));
  not_8  g21442(.A(new_n23790), .Y(new_n23791));
  nand_5 g21443(.A(new_n7125), .B(new_n4438), .Y(new_n23792));
  nand_5 g21444(.A(new_n7124), .B(n7693), .Y(new_n23793));
  nand_5 g21445(.A(new_n23793), .B(new_n23792), .Y(new_n23794));
  xor_4  g21446(.A(new_n23794), .B(new_n23791), .Y(new_n23795));
  or_5   g21447(.A(new_n23795), .B(new_n11184_1), .Y(new_n23796));
  nand_5 g21448(.A(new_n23795), .B(new_n11184_1), .Y(new_n23797));
  nand_5 g21449(.A(new_n23797), .B(new_n23796), .Y(new_n23798));
  xnor_4 g21450(.A(new_n23798), .B(new_n23788), .Y(n7575));
  not_8  g21451(.A(new_n13256), .Y(new_n23800));
  nand_5 g21452(.A(new_n12645), .B(new_n12638), .Y(new_n23801));
  nand_5 g21453(.A(new_n23801), .B(new_n12642), .Y(new_n23802));
  nand_5 g21454(.A(new_n23514), .B(new_n11118), .Y(new_n23803));
  not_8  g21455(.A(new_n11118), .Y(new_n23804));
  nand_5 g21456(.A(new_n23516), .B(new_n23804), .Y(new_n23805));
  nand_5 g21457(.A(new_n23805), .B(new_n23803), .Y(new_n23806));
  xnor_4 g21458(.A(new_n23806), .B(new_n23802), .Y(new_n23807));
  or_5   g21459(.A(new_n23807), .B(new_n23800), .Y(new_n23808));
  nand_5 g21460(.A(new_n23807), .B(new_n23800), .Y(new_n23809));
  not_8  g21461(.A(new_n12627), .Y(new_n23810));
  nor_5  g21462(.A(new_n12650_1), .B(new_n23810), .Y(new_n23811));
  nor_5  g21463(.A(new_n23811), .B(new_n12649), .Y(new_n23812));
  nand_5 g21464(.A(new_n23812), .B(new_n23809), .Y(new_n23813));
  nand_5 g21465(.A(new_n23813), .B(new_n23808), .Y(new_n23814));
  nand_5 g21466(.A(new_n23805), .B(new_n23802), .Y(new_n23815));
  nand_5 g21467(.A(new_n23815), .B(new_n23803), .Y(new_n23816));
  nand_5 g21468(.A(new_n23510), .B(new_n11230), .Y(new_n23817));
  nand_5 g21469(.A(new_n23512), .B(new_n11245_1), .Y(new_n23818));
  nand_5 g21470(.A(new_n23818), .B(new_n23817), .Y(new_n23819));
  xor_4  g21471(.A(new_n23819), .B(new_n23816), .Y(new_n23820));
  nand_5 g21472(.A(new_n23820), .B(new_n13250), .Y(new_n23821));
  or_5   g21473(.A(new_n23820), .B(new_n13250), .Y(new_n23822));
  nand_5 g21474(.A(new_n23822), .B(new_n23821), .Y(new_n23823));
  xor_4  g21475(.A(new_n23823), .B(new_n23814), .Y(n7585));
  or_5   g21476(.A(new_n23179), .B(new_n10272), .Y(new_n23825));
  nand_5 g21477(.A(new_n23179), .B(new_n10272), .Y(new_n23826));
  nand_5 g21478(.A(new_n23826), .B(new_n23825), .Y(new_n23827));
  nand_5 g21479(.A(new_n23204), .B(new_n8857), .Y(new_n23828));
  nand_5 g21480(.A(new_n23205), .B(new_n8853), .Y(new_n23829));
  nand_5 g21481(.A(new_n23211), .B(new_n8865), .Y(new_n23830));
  nand_5 g21482(.A(new_n23212), .B(new_n8861_1), .Y(new_n23831_1));
  nand_5 g21483(.A(new_n23218), .B(new_n8873), .Y(new_n23832));
  nand_5 g21484(.A(new_n23219), .B(new_n8869_1), .Y(new_n23833));
  nand_5 g21485(.A(new_n20515_1), .B(new_n8881), .Y(new_n23834));
  or_5   g21486(.A(new_n20515_1), .B(new_n8881), .Y(new_n23835));
  nand_5 g21487(.A(new_n20461), .B(new_n8889), .Y(new_n23836));
  nand_5 g21488(.A(new_n20462), .B(new_n8885), .Y(new_n23837));
  nand_5 g21489(.A(new_n20468), .B(new_n8897), .Y(new_n23838));
  nand_5 g21490(.A(new_n20469), .B(new_n8893), .Y(new_n23839));
  or_5   g21491(.A(new_n20475), .B(new_n8901), .Y(new_n23840));
  nand_5 g21492(.A(new_n20475), .B(new_n8901), .Y(new_n23841));
  nand_5 g21493(.A(new_n20479), .B(new_n8917), .Y(new_n23842_1));
  or_5   g21494(.A(new_n23842_1), .B(new_n8910), .Y(new_n23843));
  nand_5 g21495(.A(new_n23842_1), .B(new_n8910), .Y(new_n23844));
  nand_5 g21496(.A(new_n23844), .B(new_n20490_1), .Y(new_n23845));
  nand_5 g21497(.A(new_n23845), .B(new_n23843), .Y(new_n23846));
  nand_5 g21498(.A(new_n23846), .B(new_n23841), .Y(new_n23847));
  nand_5 g21499(.A(new_n23847), .B(new_n23840), .Y(new_n23848));
  nand_5 g21500(.A(new_n23848), .B(new_n23839), .Y(new_n23849_1));
  nand_5 g21501(.A(new_n23849_1), .B(new_n23838), .Y(new_n23850));
  nand_5 g21502(.A(new_n23850), .B(new_n23837), .Y(new_n23851));
  nand_5 g21503(.A(new_n23851), .B(new_n23836), .Y(new_n23852));
  nand_5 g21504(.A(new_n23852), .B(new_n23835), .Y(new_n23853));
  nand_5 g21505(.A(new_n23853), .B(new_n23834), .Y(new_n23854));
  nand_5 g21506(.A(new_n23854), .B(new_n23833), .Y(new_n23855));
  nand_5 g21507(.A(new_n23855), .B(new_n23832), .Y(new_n23856_1));
  nand_5 g21508(.A(new_n23856_1), .B(new_n23831_1), .Y(new_n23857));
  nand_5 g21509(.A(new_n23857), .B(new_n23830), .Y(new_n23858));
  nand_5 g21510(.A(new_n23858), .B(new_n23829), .Y(new_n23859));
  nand_5 g21511(.A(new_n23859), .B(new_n23828), .Y(new_n23860));
  xnor_4 g21512(.A(new_n23860), .B(new_n23827), .Y(n7588));
  nor_5  g21513(.A(new_n7717), .B(n21753), .Y(new_n23862));
  nand_5 g21514(.A(new_n23862), .B(new_n2601), .Y(new_n23863));
  not_8  g21515(.A(new_n23863), .Y(new_n23864));
  nor_5  g21516(.A(new_n23862), .B(new_n2601), .Y(new_n23865));
  nor_5  g21517(.A(new_n23865), .B(new_n23864), .Y(new_n23866));
  or_5   g21518(.A(new_n23866), .B(n3945), .Y(new_n23867));
  nand_5 g21519(.A(new_n23866), .B(n3945), .Y(new_n23868));
  xor_4  g21520(.A(new_n7717), .B(n21753), .Y(new_n23869));
  or_5   g21521(.A(new_n23869), .B(n5255), .Y(new_n23870));
  nand_5 g21522(.A(new_n23869), .B(n5255), .Y(new_n23871));
  nand_5 g21523(.A(new_n7721_1), .B(new_n5820), .Y(new_n23872));
  nand_5 g21524(.A(new_n7719), .B(n21649), .Y(new_n23873));
  nand_5 g21525(.A(new_n7682), .B(new_n5806), .Y(new_n23874));
  nand_5 g21526(.A(new_n7679_1), .B(n18274), .Y(new_n23875));
  nand_5 g21527(.A(new_n7652), .B(new_n5729), .Y(new_n23876));
  nand_5 g21528(.A(new_n7649), .B(n3828), .Y(new_n23877));
  nand_5 g21529(.A(new_n7660), .B(new_n5687_1), .Y(new_n23878));
  nand_5 g21530(.A(new_n7659), .B(n23842), .Y(new_n23879));
  nand_5 g21531(.A(n21654), .B(n2387), .Y(new_n23880));
  nand_5 g21532(.A(new_n23880), .B(new_n23879), .Y(new_n23881));
  nand_5 g21533(.A(new_n23881), .B(new_n23878), .Y(new_n23882));
  nand_5 g21534(.A(new_n23882), .B(new_n23877), .Y(new_n23883_1));
  nand_5 g21535(.A(new_n23883_1), .B(new_n23876), .Y(new_n23884));
  nand_5 g21536(.A(new_n23884), .B(new_n23875), .Y(new_n23885));
  nand_5 g21537(.A(new_n23885), .B(new_n23874), .Y(new_n23886));
  nand_5 g21538(.A(new_n23886), .B(new_n23873), .Y(new_n23887));
  nand_5 g21539(.A(new_n23887), .B(new_n23872), .Y(new_n23888_1));
  nand_5 g21540(.A(new_n23888_1), .B(new_n23871), .Y(new_n23889));
  nand_5 g21541(.A(new_n23889), .B(new_n23870), .Y(new_n23890));
  nand_5 g21542(.A(new_n23890), .B(new_n23868), .Y(new_n23891));
  nand_5 g21543(.A(new_n23891), .B(new_n23867), .Y(new_n23892));
  nand_5 g21544(.A(new_n23864), .B(new_n3321), .Y(new_n23893));
  nand_5 g21545(.A(new_n23863), .B(n13074), .Y(new_n23894));
  and_5  g21546(.A(new_n23894), .B(new_n23893), .Y(new_n23895_1));
  not_8  g21547(.A(new_n23895_1), .Y(new_n23896));
  nand_5 g21548(.A(new_n23896), .B(new_n18169), .Y(new_n23897));
  nand_5 g21549(.A(new_n23895_1), .B(n11455), .Y(new_n23898));
  nand_5 g21550(.A(new_n23898), .B(new_n23897), .Y(new_n23899_1));
  xor_4  g21551(.A(new_n23899_1), .B(new_n23892), .Y(new_n23900));
  nand_5 g21552(.A(new_n23900), .B(new_n16366), .Y(new_n23901));
  or_5   g21553(.A(new_n23900), .B(new_n16366), .Y(new_n23902));
  nand_5 g21554(.A(new_n23868), .B(new_n23867), .Y(new_n23903_1));
  xor_4  g21555(.A(new_n23903_1), .B(new_n23890), .Y(new_n23904));
  nand_5 g21556(.A(new_n23904), .B(new_n16375), .Y(new_n23905));
  or_5   g21557(.A(new_n23904), .B(new_n16375), .Y(new_n23906));
  nand_5 g21558(.A(new_n23871), .B(new_n23870), .Y(new_n23907));
  xor_4  g21559(.A(new_n23907), .B(new_n23888_1), .Y(new_n23908));
  nand_5 g21560(.A(new_n23908), .B(new_n16384), .Y(new_n23909));
  or_5   g21561(.A(new_n23908), .B(new_n16384), .Y(new_n23910));
  nand_5 g21562(.A(new_n23873), .B(new_n23872), .Y(new_n23911));
  xor_4  g21563(.A(new_n23911), .B(new_n23886), .Y(new_n23912_1));
  nand_5 g21564(.A(new_n23912_1), .B(new_n16391), .Y(new_n23913_1));
  nor_5  g21565(.A(new_n23912_1), .B(new_n16391), .Y(new_n23914));
  not_8  g21566(.A(new_n23914), .Y(new_n23915));
  nand_5 g21567(.A(new_n23875), .B(new_n23874), .Y(new_n23916));
  xor_4  g21568(.A(new_n23916), .B(new_n23884), .Y(new_n23917));
  nand_5 g21569(.A(new_n23917), .B(new_n16399), .Y(new_n23918));
  nor_5  g21570(.A(new_n23917), .B(new_n16399), .Y(new_n23919));
  not_8  g21571(.A(new_n23919), .Y(new_n23920));
  nand_5 g21572(.A(new_n23877), .B(new_n23876), .Y(new_n23921));
  xor_4  g21573(.A(new_n23921), .B(new_n23882), .Y(new_n23922));
  nand_5 g21574(.A(new_n23922), .B(new_n16405), .Y(new_n23923_1));
  or_5   g21575(.A(new_n23922), .B(new_n16405), .Y(new_n23924_1));
  nand_5 g21576(.A(new_n5678), .B(new_n2506), .Y(new_n23925));
  nand_5 g21577(.A(new_n23925), .B(new_n23880), .Y(new_n23926));
  nor_5  g21578(.A(new_n23926), .B(new_n16412), .Y(new_n23927));
  nand_5 g21579(.A(new_n23879), .B(new_n23878), .Y(new_n23928));
  nand_5 g21580(.A(new_n23928), .B(new_n16420), .Y(new_n23929));
  nand_5 g21581(.A(new_n23929), .B(new_n23927), .Y(new_n23930));
  xor_4  g21582(.A(new_n23928), .B(new_n23880), .Y(new_n23931));
  nand_5 g21583(.A(new_n23931), .B(new_n16419_1), .Y(new_n23932));
  nand_5 g21584(.A(new_n23932), .B(new_n23930), .Y(new_n23933));
  nand_5 g21585(.A(new_n23933), .B(new_n23924_1), .Y(new_n23934));
  nand_5 g21586(.A(new_n23934), .B(new_n23923_1), .Y(new_n23935_1));
  nand_5 g21587(.A(new_n23935_1), .B(new_n23920), .Y(new_n23936));
  nand_5 g21588(.A(new_n23936), .B(new_n23918), .Y(new_n23937));
  nand_5 g21589(.A(new_n23937), .B(new_n23915), .Y(new_n23938));
  nand_5 g21590(.A(new_n23938), .B(new_n23913_1), .Y(new_n23939));
  nand_5 g21591(.A(new_n23939), .B(new_n23910), .Y(new_n23940));
  nand_5 g21592(.A(new_n23940), .B(new_n23909), .Y(new_n23941));
  nand_5 g21593(.A(new_n23941), .B(new_n23906), .Y(new_n23942_1));
  nand_5 g21594(.A(new_n23942_1), .B(new_n23905), .Y(new_n23943));
  nand_5 g21595(.A(new_n23943), .B(new_n23902), .Y(new_n23944));
  nand_5 g21596(.A(new_n23944), .B(new_n23901), .Y(new_n23945));
  nand_5 g21597(.A(new_n23898), .B(new_n23892), .Y(new_n23946));
  nand_5 g21598(.A(new_n23946), .B(new_n23897), .Y(new_n23947));
  or_5   g21599(.A(new_n23893), .B(n23463), .Y(new_n23948));
  nand_5 g21600(.A(new_n23893), .B(n23463), .Y(new_n23949));
  and_5  g21601(.A(new_n23949), .B(new_n23948), .Y(new_n23950));
  or_5   g21602(.A(new_n23950), .B(n23250), .Y(new_n23951));
  nand_5 g21603(.A(new_n23950), .B(n23250), .Y(new_n23952));
  nand_5 g21604(.A(new_n23952), .B(new_n23951), .Y(new_n23953));
  xnor_4 g21605(.A(new_n23953), .B(new_n23947), .Y(new_n23954_1));
  nand_5 g21606(.A(new_n23954_1), .B(new_n16453), .Y(new_n23955));
  not_8  g21607(.A(new_n23955), .Y(new_n23956));
  nor_5  g21608(.A(new_n23954_1), .B(new_n16453), .Y(new_n23957));
  nor_5  g21609(.A(new_n23957), .B(new_n23956), .Y(new_n23958_1));
  xor_4  g21610(.A(new_n23958_1), .B(new_n23945), .Y(n7598));
  nand_5 g21611(.A(new_n20373), .B(new_n20372), .Y(new_n23960));
  xor_4  g21612(.A(new_n23960), .B(new_n20375), .Y(n7607));
  nand_5 g21613(.A(new_n5616), .B(new_n5615), .Y(new_n23962));
  xor_4  g21614(.A(new_n23962), .B(new_n5649), .Y(n7610));
  nand_5 g21615(.A(new_n3651), .B(new_n3652), .Y(new_n23964));
  xnor_4 g21616(.A(new_n23964), .B(new_n3669), .Y(n7616));
  nand_5 g21617(.A(new_n13220), .B(new_n7166), .Y(new_n23966));
  nand_5 g21618(.A(n10514), .B(n6105), .Y(new_n23967));
  nand_5 g21619(.A(new_n13224), .B(new_n7170), .Y(new_n23968));
  nand_5 g21620(.A(n18649), .B(n3795), .Y(new_n23969));
  nand_5 g21621(.A(new_n7175), .B(new_n13227), .Y(new_n23970));
  nand_5 g21622(.A(n25464), .B(n6218), .Y(new_n23971));
  nand_5 g21623(.A(new_n12632), .B(new_n7178), .Y(new_n23972));
  nand_5 g21624(.A(n20470), .B(n4590), .Y(new_n23973));
  nand_5 g21625(.A(new_n7182), .B(new_n12539), .Y(new_n23974_1));
  nand_5 g21626(.A(n26752), .B(n21222), .Y(new_n23975));
  nand_5 g21627(.A(new_n11063_1), .B(new_n7185), .Y(new_n23976));
  nand_5 g21628(.A(n9832), .B(n6513), .Y(new_n23977));
  nand_5 g21629(.A(new_n7188), .B(new_n10982), .Y(new_n23978));
  nand_5 g21630(.A(n3918), .B(n1558), .Y(new_n23979));
  nand_5 g21631(.A(new_n18781), .B(new_n18778), .Y(new_n23980));
  nand_5 g21632(.A(new_n23980), .B(new_n18780_1), .Y(new_n23981));
  nand_5 g21633(.A(new_n23981), .B(new_n23979), .Y(new_n23982));
  nand_5 g21634(.A(new_n23982), .B(new_n23978), .Y(new_n23983));
  nand_5 g21635(.A(new_n23983), .B(new_n23977), .Y(new_n23984));
  nand_5 g21636(.A(new_n23984), .B(new_n23976), .Y(new_n23985));
  nand_5 g21637(.A(new_n23985), .B(new_n23975), .Y(new_n23986_1));
  nand_5 g21638(.A(new_n23986_1), .B(new_n23974_1), .Y(new_n23987));
  nand_5 g21639(.A(new_n23987), .B(new_n23973), .Y(new_n23988));
  nand_5 g21640(.A(new_n23988), .B(new_n23972), .Y(new_n23989));
  nand_5 g21641(.A(new_n23989), .B(new_n23971), .Y(new_n23990));
  nand_5 g21642(.A(new_n23990), .B(new_n23970), .Y(new_n23991));
  nand_5 g21643(.A(new_n23991), .B(new_n23969), .Y(new_n23992));
  nand_5 g21644(.A(new_n23992), .B(new_n23968), .Y(new_n23993));
  nand_5 g21645(.A(new_n23993), .B(new_n23967), .Y(new_n23994));
  nand_5 g21646(.A(new_n23994), .B(new_n23966), .Y(new_n23995));
  not_8  g21647(.A(new_n23995), .Y(new_n23996));
  nand_5 g21648(.A(new_n23967), .B(new_n23966), .Y(new_n23997));
  xor_4  g21649(.A(new_n23997), .B(new_n23993), .Y(new_n23998));
  not_8  g21650(.A(new_n23998), .Y(new_n23999));
  or_5   g21651(.A(new_n23999), .B(n9872), .Y(new_n24000));
  nand_5 g21652(.A(new_n23999), .B(n9872), .Y(new_n24001));
  nand_5 g21653(.A(new_n23969), .B(new_n23968), .Y(new_n24002_1));
  xor_4  g21654(.A(new_n24002_1), .B(new_n23991), .Y(new_n24003));
  not_8  g21655(.A(new_n24003), .Y(new_n24004_1));
  or_5   g21656(.A(new_n24004_1), .B(n5842), .Y(new_n24005));
  nand_5 g21657(.A(new_n24004_1), .B(n5842), .Y(new_n24006));
  nand_5 g21658(.A(new_n23971), .B(new_n23970), .Y(new_n24007));
  xor_4  g21659(.A(new_n24007), .B(new_n23989), .Y(new_n24008));
  not_8  g21660(.A(new_n24008), .Y(new_n24009));
  or_5   g21661(.A(new_n24009), .B(n6379), .Y(new_n24010));
  nand_5 g21662(.A(new_n24009), .B(n6379), .Y(new_n24011));
  nand_5 g21663(.A(new_n23973), .B(new_n23972), .Y(new_n24012));
  xor_4  g21664(.A(new_n24012), .B(new_n23987), .Y(new_n24013));
  not_8  g21665(.A(new_n24013), .Y(new_n24014));
  or_5   g21666(.A(new_n24014), .B(n2102), .Y(new_n24015));
  nand_5 g21667(.A(new_n24014), .B(n2102), .Y(new_n24016));
  not_8  g21668(.A(n17954), .Y(new_n24017));
  nand_5 g21669(.A(new_n23975), .B(new_n23974_1), .Y(new_n24018));
  xor_4  g21670(.A(new_n24018), .B(new_n23985), .Y(new_n24019));
  nand_5 g21671(.A(new_n24019), .B(new_n24017), .Y(new_n24020));
  nor_5  g21672(.A(new_n24019), .B(new_n24017), .Y(new_n24021));
  not_8  g21673(.A(new_n24021), .Y(new_n24022));
  not_8  g21674(.A(n8256), .Y(new_n24023));
  nand_5 g21675(.A(new_n23977), .B(new_n23976), .Y(new_n24024));
  xor_4  g21676(.A(new_n24024), .B(new_n23983), .Y(new_n24025));
  nand_5 g21677(.A(new_n24025), .B(new_n24023), .Y(new_n24026));
  nor_5  g21678(.A(new_n24025), .B(new_n24023), .Y(new_n24027));
  not_8  g21679(.A(new_n24027), .Y(new_n24028));
  not_8  g21680(.A(n24150), .Y(new_n24029));
  nand_5 g21681(.A(new_n23979), .B(new_n23978), .Y(new_n24030));
  xor_4  g21682(.A(new_n24030), .B(new_n23981), .Y(new_n24031));
  nand_5 g21683(.A(new_n24031), .B(new_n24029), .Y(new_n24032_1));
  nor_5  g21684(.A(new_n24031), .B(new_n24029), .Y(new_n24033));
  not_8  g21685(.A(new_n18785), .Y(new_n24034));
  not_8  g21686(.A(new_n18786), .Y(new_n24035));
  nor_5  g21687(.A(new_n24035), .B(new_n18775), .Y(new_n24036));
  nor_5  g21688(.A(new_n24036), .B(new_n24034), .Y(new_n24037));
  or_5   g21689(.A(new_n24037), .B(new_n24033), .Y(new_n24038));
  nand_5 g21690(.A(new_n24038), .B(new_n24032_1), .Y(new_n24039_1));
  nand_5 g21691(.A(new_n24039_1), .B(new_n24028), .Y(new_n24040));
  nand_5 g21692(.A(new_n24040), .B(new_n24026), .Y(new_n24041));
  nand_5 g21693(.A(new_n24041), .B(new_n24022), .Y(new_n24042));
  nand_5 g21694(.A(new_n24042), .B(new_n24020), .Y(new_n24043));
  nand_5 g21695(.A(new_n24043), .B(new_n24016), .Y(new_n24044));
  nand_5 g21696(.A(new_n24044), .B(new_n24015), .Y(new_n24045));
  nand_5 g21697(.A(new_n24045), .B(new_n24011), .Y(new_n24046));
  nand_5 g21698(.A(new_n24046), .B(new_n24010), .Y(new_n24047));
  nand_5 g21699(.A(new_n24047), .B(new_n24006), .Y(new_n24048_1));
  nand_5 g21700(.A(new_n24048_1), .B(new_n24005), .Y(new_n24049));
  nand_5 g21701(.A(new_n24049), .B(new_n24001), .Y(new_n24050));
  nand_5 g21702(.A(new_n24050), .B(new_n24000), .Y(new_n24051));
  nor_5  g21703(.A(new_n24051), .B(new_n23996), .Y(new_n24052_1));
  xor_4  g21704(.A(new_n24052_1), .B(new_n17843), .Y(new_n24053));
  not_8  g21705(.A(new_n17710), .Y(new_n24054));
  xor_4  g21706(.A(new_n24051), .B(new_n23995), .Y(new_n24055));
  or_5   g21707(.A(new_n24055), .B(new_n24054), .Y(new_n24056));
  nand_5 g21708(.A(new_n24055), .B(new_n24054), .Y(new_n24057));
  nand_5 g21709(.A(new_n24001), .B(new_n24000), .Y(new_n24058));
  xnor_4 g21710(.A(new_n24058), .B(new_n24049), .Y(new_n24059));
  or_5   g21711(.A(new_n24059), .B(new_n17756), .Y(new_n24060));
  nand_5 g21712(.A(new_n24059), .B(new_n17756), .Y(new_n24061));
  nand_5 g21713(.A(new_n24006), .B(new_n24005), .Y(new_n24062));
  xnor_4 g21714(.A(new_n24062), .B(new_n24047), .Y(new_n24063));
  or_5   g21715(.A(new_n24063), .B(new_n17763), .Y(new_n24064));
  nand_5 g21716(.A(new_n24063), .B(new_n17763), .Y(new_n24065));
  nand_5 g21717(.A(new_n24011), .B(new_n24010), .Y(new_n24066));
  xnor_4 g21718(.A(new_n24066), .B(new_n24045), .Y(new_n24067));
  or_5   g21719(.A(new_n24067), .B(new_n17770), .Y(new_n24068));
  nand_5 g21720(.A(new_n24067), .B(new_n17770), .Y(new_n24069));
  nand_5 g21721(.A(new_n24016), .B(new_n24015), .Y(new_n24070));
  xnor_4 g21722(.A(new_n24070), .B(new_n24043), .Y(new_n24071));
  or_5   g21723(.A(new_n24071), .B(new_n17777), .Y(new_n24072));
  nand_5 g21724(.A(new_n24071), .B(new_n17777), .Y(new_n24073));
  nand_5 g21725(.A(new_n24022), .B(new_n24020), .Y(new_n24074));
  xor_4  g21726(.A(new_n24074), .B(new_n24041), .Y(new_n24075));
  nand_5 g21727(.A(new_n24075), .B(new_n17784_1), .Y(new_n24076));
  or_5   g21728(.A(new_n24075), .B(new_n17784_1), .Y(new_n24077));
  nand_5 g21729(.A(new_n24028), .B(new_n24026), .Y(new_n24078));
  xor_4  g21730(.A(new_n24078), .B(new_n24039_1), .Y(new_n24079));
  nand_5 g21731(.A(new_n24079), .B(new_n17791), .Y(new_n24080));
  or_5   g21732(.A(new_n24079), .B(new_n17791), .Y(new_n24081));
  not_8  g21733(.A(new_n24033), .Y(new_n24082));
  nand_5 g21734(.A(new_n24082), .B(new_n24032_1), .Y(new_n24083));
  xor_4  g21735(.A(new_n24083), .B(new_n24037), .Y(new_n24084));
  or_5   g21736(.A(new_n24084), .B(new_n17797), .Y(new_n24085_1));
  nand_5 g21737(.A(new_n24084), .B(new_n17797), .Y(new_n24086));
  nand_5 g21738(.A(new_n18790), .B(new_n18773), .Y(new_n24087));
  nand_5 g21739(.A(new_n24087), .B(new_n18789), .Y(new_n24088));
  nand_5 g21740(.A(new_n24088), .B(new_n24086), .Y(new_n24089));
  nand_5 g21741(.A(new_n24089), .B(new_n24085_1), .Y(new_n24090));
  nand_5 g21742(.A(new_n24090), .B(new_n24081), .Y(new_n24091));
  nand_5 g21743(.A(new_n24091), .B(new_n24080), .Y(new_n24092_1));
  nand_5 g21744(.A(new_n24092_1), .B(new_n24077), .Y(new_n24093_1));
  nand_5 g21745(.A(new_n24093_1), .B(new_n24076), .Y(new_n24094));
  nand_5 g21746(.A(new_n24094), .B(new_n24073), .Y(new_n24095));
  nand_5 g21747(.A(new_n24095), .B(new_n24072), .Y(new_n24096_1));
  nand_5 g21748(.A(new_n24096_1), .B(new_n24069), .Y(new_n24097_1));
  nand_5 g21749(.A(new_n24097_1), .B(new_n24068), .Y(new_n24098));
  nand_5 g21750(.A(new_n24098), .B(new_n24065), .Y(new_n24099));
  nand_5 g21751(.A(new_n24099), .B(new_n24064), .Y(new_n24100));
  nand_5 g21752(.A(new_n24100), .B(new_n24061), .Y(new_n24101));
  nand_5 g21753(.A(new_n24101), .B(new_n24060), .Y(new_n24102));
  nand_5 g21754(.A(new_n24102), .B(new_n24057), .Y(new_n24103));
  nand_5 g21755(.A(new_n24103), .B(new_n24056), .Y(new_n24104));
  xnor_4 g21756(.A(new_n24104), .B(new_n24053), .Y(n7630));
  nand_5 g21757(.A(new_n21324), .B(new_n21314), .Y(new_n24106));
  nand_5 g21758(.A(new_n24106), .B(new_n21315), .Y(n7643));
  nand_5 g21759(.A(new_n13933), .B(new_n13932), .Y(new_n24108));
  xor_4  g21760(.A(new_n24108), .B(new_n13966), .Y(n7647));
  nand_5 g21761(.A(new_n11567), .B(new_n11566_1), .Y(new_n24110));
  xor_4  g21762(.A(new_n24110), .B(new_n11609), .Y(n7679));
  nand_5 g21763(.A(new_n22828), .B(new_n22826), .Y(new_n24112));
  xnor_4 g21764(.A(new_n24112), .B(new_n22856), .Y(n7686));
  nand_5 g21765(.A(new_n20773), .B(new_n20770), .Y(new_n24114));
  xor_4  g21766(.A(new_n24114), .B(new_n20767), .Y(n7698));
  nand_5 g21767(.A(new_n22010), .B(new_n21990), .Y(new_n24116));
  xor_4  g21768(.A(new_n24116), .B(new_n22009), .Y(n7708));
  nand_5 g21769(.A(new_n18565), .B(new_n18563), .Y(new_n24118));
  nand_5 g21770(.A(new_n24118), .B(new_n18564), .Y(new_n24119_1));
  nand_5 g21771(.A(new_n6844), .B(n3740), .Y(new_n24120));
  nand_5 g21772(.A(new_n6843), .B(new_n5496), .Y(new_n24121));
  nand_5 g21773(.A(new_n24121), .B(new_n24120), .Y(new_n24122));
  xor_4  g21774(.A(new_n24122), .B(new_n24119_1), .Y(new_n24123));
  not_8  g21775(.A(new_n24123), .Y(new_n24124));
  nand_5 g21776(.A(new_n20737), .B(n3324), .Y(new_n24125));
  nand_5 g21777(.A(new_n20735), .B(new_n18124), .Y(new_n24126));
  nand_5 g21778(.A(new_n24126), .B(new_n24125), .Y(new_n24127));
  nand_5 g21779(.A(new_n3291), .B(new_n18127), .Y(new_n24128));
  nand_5 g21780(.A(new_n3302), .B(n17911), .Y(new_n24129_1));
  nand_5 g21781(.A(new_n3189), .B(new_n18133), .Y(new_n24130));
  nand_5 g21782(.A(new_n3202), .B(n21997), .Y(new_n24131));
  nand_5 g21783(.A(new_n9836), .B(new_n9833_1), .Y(new_n24132));
  nand_5 g21784(.A(new_n24132), .B(new_n9835), .Y(new_n24133_1));
  nand_5 g21785(.A(new_n24133_1), .B(new_n24131), .Y(new_n24134));
  nand_5 g21786(.A(new_n24134), .B(new_n24130), .Y(new_n24135));
  nand_5 g21787(.A(new_n24135), .B(new_n24129_1), .Y(new_n24136));
  nand_5 g21788(.A(new_n24136), .B(new_n24128), .Y(new_n24137));
  xnor_4 g21789(.A(new_n24137), .B(new_n24127), .Y(new_n24138));
  or_5   g21790(.A(new_n24138), .B(new_n24124), .Y(new_n24139));
  nand_5 g21791(.A(new_n24138), .B(new_n24124), .Y(new_n24140));
  nand_5 g21792(.A(new_n24140), .B(new_n24139), .Y(new_n24141_1));
  nand_5 g21793(.A(new_n24128), .B(new_n24129_1), .Y(new_n24142));
  xor_4  g21794(.A(new_n24142), .B(new_n24135), .Y(new_n24143));
  or_5   g21795(.A(new_n24143), .B(new_n18567), .Y(new_n24144));
  nand_5 g21796(.A(new_n24143), .B(new_n18567), .Y(new_n24145_1));
  nand_5 g21797(.A(new_n24130), .B(new_n24131), .Y(new_n24146_1));
  xor_4  g21798(.A(new_n24146_1), .B(new_n24133_1), .Y(new_n24147));
  or_5   g21799(.A(new_n24147), .B(new_n18447), .Y(new_n24148));
  nand_5 g21800(.A(new_n24147), .B(new_n18447), .Y(new_n24149));
  nand_5 g21801(.A(new_n9840), .B(new_n9825), .Y(new_n24150_1));
  nand_5 g21802(.A(new_n24150_1), .B(new_n9839), .Y(new_n24151));
  nand_5 g21803(.A(new_n24151), .B(new_n24149), .Y(new_n24152));
  nand_5 g21804(.A(new_n24152), .B(new_n24148), .Y(new_n24153));
  nand_5 g21805(.A(new_n24153), .B(new_n24145_1), .Y(new_n24154));
  nand_5 g21806(.A(new_n24154), .B(new_n24144), .Y(new_n24155_1));
  xor_4  g21807(.A(new_n24155_1), .B(new_n24141_1), .Y(n7780));
  nand_5 g21808(.A(new_n2695), .B(new_n4966_1), .Y(new_n24157));
  nand_5 g21809(.A(new_n2696), .B(n18880), .Y(new_n24158));
  nand_5 g21810(.A(new_n11228), .B(new_n11226), .Y(new_n24159));
  nand_5 g21811(.A(new_n24159), .B(new_n11227), .Y(new_n24160_1));
  nand_5 g21812(.A(new_n24160_1), .B(new_n24158), .Y(new_n24161));
  nand_5 g21813(.A(new_n24161), .B(new_n24157), .Y(new_n24162));
  nor_5  g21814(.A(new_n24162), .B(new_n16638), .Y(new_n24163));
  not_8  g21815(.A(new_n24163), .Y(new_n24164));
  nand_5 g21816(.A(new_n24162), .B(new_n16638), .Y(new_n24165));
  and_5  g21817(.A(new_n24165), .B(new_n24164), .Y(new_n24166));
  nand_5 g21818(.A(new_n19790), .B(new_n11642), .Y(new_n24167_1));
  nand_5 g21819(.A(new_n19789_1), .B(new_n11640), .Y(new_n24168));
  nand_5 g21820(.A(new_n24168), .B(new_n24167_1), .Y(new_n24169));
  nand_5 g21821(.A(new_n19793), .B(new_n2840), .Y(new_n24170_1));
  nand_5 g21822(.A(new_n19791), .B(new_n2841), .Y(new_n24171));
  nand_5 g21823(.A(new_n11240), .B(new_n11232), .Y(new_n24172_1));
  nand_5 g21824(.A(new_n24172_1), .B(new_n11239), .Y(new_n24173));
  nand_5 g21825(.A(new_n24173), .B(new_n24171), .Y(new_n24174));
  nand_5 g21826(.A(new_n24174), .B(new_n24170_1), .Y(new_n24175));
  not_8  g21827(.A(new_n24175), .Y(new_n24176));
  xor_4  g21828(.A(new_n24176), .B(new_n24169), .Y(new_n24177_1));
  nand_5 g21829(.A(new_n24177_1), .B(new_n24166), .Y(new_n24178));
  or_5   g21830(.A(new_n24177_1), .B(new_n24166), .Y(new_n24179));
  nand_5 g21831(.A(new_n24179), .B(new_n24178), .Y(new_n24180));
  nand_5 g21832(.A(new_n24157), .B(new_n24158), .Y(new_n24181));
  xor_4  g21833(.A(new_n24181), .B(new_n24160_1), .Y(new_n24182));
  nand_5 g21834(.A(new_n24170_1), .B(new_n24171), .Y(new_n24183));
  xor_4  g21835(.A(new_n24183), .B(new_n24173), .Y(new_n24184));
  or_5   g21836(.A(new_n24184), .B(new_n24182), .Y(new_n24185));
  nand_5 g21837(.A(new_n24184), .B(new_n24182), .Y(new_n24186));
  not_8  g21838(.A(new_n11244), .Y(new_n24187));
  not_8  g21839(.A(new_n11246), .Y(new_n24188));
  nor_5  g21840(.A(new_n24188), .B(new_n11224), .Y(new_n24189));
  nor_5  g21841(.A(new_n24189), .B(new_n24187), .Y(new_n24190));
  nand_5 g21842(.A(new_n24190), .B(new_n24186), .Y(new_n24191));
  nand_5 g21843(.A(new_n24191), .B(new_n24185), .Y(new_n24192));
  xor_4  g21844(.A(new_n24192), .B(new_n24180), .Y(n7794));
  nand_5 g21845(.A(new_n19926), .B(new_n19925), .Y(new_n24194));
  xor_4  g21846(.A(new_n24194), .B(new_n19931), .Y(n7811));
  nand_5 g21847(.A(new_n19880), .B(new_n19881), .Y(new_n24196_1));
  xor_4  g21848(.A(new_n24196_1), .B(new_n19887), .Y(n7830));
  nand_5 g21849(.A(new_n23830), .B(new_n23831_1), .Y(new_n24198));
  xnor_4 g21850(.A(new_n24198), .B(new_n23856_1), .Y(n7834));
  nand_5 g21851(.A(new_n12602), .B(new_n12603), .Y(new_n24200));
  xnor_4 g21852(.A(new_n24200), .B(new_n12621_1), .Y(n7884));
  nand_5 g21853(.A(new_n3256), .B(new_n3255), .Y(new_n24202));
  xnor_4 g21854(.A(new_n24202), .B(new_n3258), .Y(n7937));
  nand_5 g21855(.A(new_n3208_1), .B(new_n3207), .Y(new_n24204));
  xnor_4 g21856(.A(new_n24204), .B(new_n3270), .Y(n7943));
  nand_5 g21857(.A(new_n11181), .B(new_n11182_1), .Y(new_n24206));
  xor_4  g21858(.A(new_n24206), .B(new_n11218), .Y(n7950));
  nand_5 g21859(.A(new_n22301), .B(new_n17664_1), .Y(new_n24208));
  nand_5 g21860(.A(new_n22298), .B(new_n23480_1), .Y(new_n24209));
  nand_5 g21861(.A(new_n24209), .B(new_n24208), .Y(new_n24210));
  nand_5 g21862(.A(new_n22304), .B(new_n17667), .Y(new_n24211));
  nand_5 g21863(.A(new_n22308), .B(new_n17666), .Y(new_n24212));
  nand_5 g21864(.A(new_n22312), .B(new_n17671), .Y(new_n24213));
  nand_5 g21865(.A(new_n22314), .B(new_n17670), .Y(new_n24214));
  nand_5 g21866(.A(new_n17441), .B(new_n17411), .Y(new_n24215));
  nand_5 g21867(.A(new_n24215), .B(new_n17439), .Y(new_n24216));
  nand_5 g21868(.A(new_n24216), .B(new_n24214), .Y(new_n24217));
  nand_5 g21869(.A(new_n24217), .B(new_n24213), .Y(new_n24218));
  nand_5 g21870(.A(new_n24218), .B(new_n24212), .Y(new_n24219));
  nand_5 g21871(.A(new_n24219), .B(new_n24211), .Y(new_n24220));
  xor_4  g21872(.A(new_n24220), .B(new_n24210), .Y(n7959));
  nand_5 g21873(.A(new_n19922_1), .B(new_n19921), .Y(new_n24222));
  xor_4  g21874(.A(new_n24222), .B(new_n19935), .Y(n7968));
  nand_5 g21875(.A(new_n21021), .B(new_n21019), .Y(new_n24224));
  xor_4  g21876(.A(new_n24224), .B(new_n21024), .Y(n7992));
  nand_5 g21877(.A(new_n14744), .B(n9554), .Y(new_n24226));
  nand_5 g21878(.A(new_n14743), .B(new_n5420), .Y(new_n24227));
  nand_5 g21879(.A(new_n24227), .B(new_n24226), .Y(new_n24228_1));
  nand_5 g21880(.A(new_n14730), .B(n26408), .Y(new_n24229));
  nand_5 g21881(.A(new_n14729), .B(new_n5371), .Y(new_n24230));
  nand_5 g21882(.A(new_n19945), .B(new_n19943), .Y(new_n24231));
  nand_5 g21883(.A(new_n24231), .B(new_n19944), .Y(new_n24232));
  nand_5 g21884(.A(new_n24232), .B(new_n24230), .Y(new_n24233));
  nand_5 g21885(.A(new_n24233), .B(new_n24229), .Y(new_n24234));
  xor_4  g21886(.A(new_n24234), .B(new_n24228_1), .Y(new_n24235));
  nand_5 g21887(.A(new_n24235), .B(new_n21213), .Y(new_n24236));
  not_8  g21888(.A(new_n24235), .Y(new_n24237));
  nand_5 g21889(.A(new_n24237), .B(new_n21212), .Y(new_n24238));
  nand_5 g21890(.A(new_n24238), .B(new_n24236), .Y(new_n24239));
  nand_5 g21891(.A(new_n24229), .B(new_n24230), .Y(new_n24240));
  xor_4  g21892(.A(new_n24240), .B(new_n24232), .Y(new_n24241));
  not_8  g21893(.A(new_n24241), .Y(new_n24242));
  nand_5 g21894(.A(new_n24242), .B(new_n21219), .Y(new_n24243));
  nand_5 g21895(.A(new_n24241), .B(new_n21220), .Y(new_n24244));
  nand_5 g21896(.A(new_n21226_1), .B(new_n19949), .Y(new_n24245));
  nand_5 g21897(.A(new_n21227), .B(new_n19947), .Y(new_n24246));
  nand_5 g21898(.A(new_n21233), .B(new_n19913), .Y(new_n24247));
  nand_5 g21899(.A(new_n21234), .B(new_n19912), .Y(new_n24248));
  nand_5 g21900(.A(new_n21240), .B(new_n19918), .Y(new_n24249));
  nand_5 g21901(.A(new_n21241), .B(new_n19917), .Y(new_n24250));
  nand_5 g21902(.A(new_n14847), .B(new_n14826_1), .Y(new_n24251));
  nand_5 g21903(.A(new_n24251), .B(new_n14850), .Y(new_n24252));
  nand_5 g21904(.A(new_n24252), .B(new_n24250), .Y(new_n24253));
  nand_5 g21905(.A(new_n24253), .B(new_n24249), .Y(new_n24254));
  nand_5 g21906(.A(new_n24254), .B(new_n24248), .Y(new_n24255));
  nand_5 g21907(.A(new_n24255), .B(new_n24247), .Y(new_n24256));
  nand_5 g21908(.A(new_n24256), .B(new_n24246), .Y(new_n24257));
  nand_5 g21909(.A(new_n24257), .B(new_n24245), .Y(new_n24258_1));
  nand_5 g21910(.A(new_n24258_1), .B(new_n24244), .Y(new_n24259));
  nand_5 g21911(.A(new_n24259), .B(new_n24243), .Y(new_n24260_1));
  xor_4  g21912(.A(new_n24260_1), .B(new_n24239), .Y(n7999));
  nand_5 g21913(.A(new_n20604_1), .B(new_n20605), .Y(new_n24262));
  xnor_4 g21914(.A(new_n24262), .B(new_n20619), .Y(n8027));
  nand_5 g21915(.A(new_n7087), .B(new_n6382), .Y(new_n24264));
  nand_5 g21916(.A(new_n7092), .B(n8614), .Y(new_n24265));
  nand_5 g21917(.A(new_n7095), .B(new_n6386), .Y(new_n24266));
  nand_5 g21918(.A(new_n7100), .B(n15182), .Y(new_n24267));
  nand_5 g21919(.A(new_n7103), .B(new_n6390), .Y(new_n24268));
  nand_5 g21920(.A(new_n7108), .B(n27037), .Y(new_n24269));
  nand_5 g21921(.A(new_n7111), .B(new_n6394), .Y(new_n24270));
  nand_5 g21922(.A(new_n7116), .B(n8964), .Y(new_n24271));
  nand_5 g21923(.A(new_n7120), .B(new_n4512), .Y(new_n24272));
  nand_5 g21924(.A(new_n16652), .B(n20151), .Y(new_n24273));
  nand_5 g21925(.A(new_n23793), .B(new_n23790), .Y(new_n24274));
  nand_5 g21926(.A(new_n24274), .B(new_n23792), .Y(new_n24275));
  nand_5 g21927(.A(new_n24275), .B(new_n24273), .Y(new_n24276));
  nand_5 g21928(.A(new_n24276), .B(new_n24272), .Y(new_n24277));
  nand_5 g21929(.A(new_n24277), .B(new_n24271), .Y(new_n24278_1));
  nand_5 g21930(.A(new_n24278_1), .B(new_n24270), .Y(new_n24279));
  nand_5 g21931(.A(new_n24279), .B(new_n24269), .Y(new_n24280));
  nand_5 g21932(.A(new_n24280), .B(new_n24268), .Y(new_n24281));
  nand_5 g21933(.A(new_n24281), .B(new_n24267), .Y(new_n24282));
  nand_5 g21934(.A(new_n24282), .B(new_n24266), .Y(new_n24283));
  nand_5 g21935(.A(new_n24283), .B(new_n24265), .Y(new_n24284));
  nand_5 g21936(.A(new_n24284), .B(new_n24264), .Y(new_n24285));
  nor_5  g21937(.A(new_n24285), .B(new_n7043), .Y(new_n24286));
  or_5   g21938(.A(new_n24286), .B(new_n24164), .Y(new_n24287));
  nand_5 g21939(.A(new_n24286), .B(new_n24164), .Y(new_n24288));
  xor_4  g21940(.A(new_n24285), .B(new_n7044), .Y(new_n24289_1));
  nor_5  g21941(.A(new_n24289_1), .B(new_n24166), .Y(new_n24290));
  and_5  g21942(.A(new_n24289_1), .B(new_n24166), .Y(new_n24291));
  not_8  g21943(.A(new_n24182), .Y(new_n24292));
  nand_5 g21944(.A(new_n24264), .B(new_n24265), .Y(new_n24293));
  xor_4  g21945(.A(new_n24293), .B(new_n24283), .Y(new_n24294));
  nand_5 g21946(.A(new_n24294), .B(new_n24292), .Y(new_n24295));
  not_8  g21947(.A(new_n24295), .Y(new_n24296));
  nor_5  g21948(.A(new_n24294), .B(new_n24292), .Y(new_n24297_1));
  nand_5 g21949(.A(new_n24266), .B(new_n24267), .Y(new_n24298));
  xor_4  g21950(.A(new_n24298), .B(new_n24281), .Y(new_n24299));
  nand_5 g21951(.A(new_n24299), .B(new_n11245_1), .Y(new_n24300));
  not_8  g21952(.A(new_n24300), .Y(new_n24301));
  nor_5  g21953(.A(new_n24299), .B(new_n11245_1), .Y(new_n24302));
  nand_5 g21954(.A(new_n24268), .B(new_n24269), .Y(new_n24303));
  xor_4  g21955(.A(new_n24303), .B(new_n24279), .Y(new_n24304));
  nand_5 g21956(.A(new_n24304), .B(new_n23804), .Y(new_n24305));
  not_8  g21957(.A(new_n24305), .Y(new_n24306));
  nor_5  g21958(.A(new_n24304), .B(new_n23804), .Y(new_n24307_1));
  nand_5 g21959(.A(new_n24270), .B(new_n24271), .Y(new_n24308));
  xor_4  g21960(.A(new_n24308), .B(new_n24277), .Y(new_n24309));
  nand_5 g21961(.A(new_n24309), .B(new_n12643), .Y(new_n24310));
  not_8  g21962(.A(new_n24310), .Y(new_n24311));
  nor_5  g21963(.A(new_n24309), .B(new_n12643), .Y(new_n24312));
  nand_5 g21964(.A(new_n24272), .B(new_n24273), .Y(new_n24313));
  xor_4  g21965(.A(new_n24313), .B(new_n24275), .Y(new_n24314));
  nand_5 g21966(.A(new_n24314), .B(new_n12589), .Y(new_n24315));
  or_5   g21967(.A(new_n24314), .B(new_n12589), .Y(new_n24316));
  nand_5 g21968(.A(new_n23797), .B(new_n23788), .Y(new_n24317));
  nand_5 g21969(.A(new_n24317), .B(new_n23796), .Y(new_n24318));
  nand_5 g21970(.A(new_n24318), .B(new_n24316), .Y(new_n24319_1));
  nand_5 g21971(.A(new_n24319_1), .B(new_n24315), .Y(new_n24320));
  not_8  g21972(.A(new_n24320), .Y(new_n24321));
  nor_5  g21973(.A(new_n24321), .B(new_n24312), .Y(new_n24322));
  nor_5  g21974(.A(new_n24322), .B(new_n24311), .Y(new_n24323_1));
  nor_5  g21975(.A(new_n24323_1), .B(new_n24307_1), .Y(new_n24324));
  nor_5  g21976(.A(new_n24324), .B(new_n24306), .Y(new_n24325));
  nor_5  g21977(.A(new_n24325), .B(new_n24302), .Y(new_n24326));
  nor_5  g21978(.A(new_n24326), .B(new_n24301), .Y(new_n24327_1));
  nor_5  g21979(.A(new_n24327_1), .B(new_n24297_1), .Y(new_n24328));
  nor_5  g21980(.A(new_n24328), .B(new_n24296), .Y(new_n24329));
  nor_5  g21981(.A(new_n24329), .B(new_n24291), .Y(new_n24330));
  nor_5  g21982(.A(new_n24330), .B(new_n24290), .Y(new_n24331));
  nand_5 g21983(.A(new_n24331), .B(new_n24288), .Y(new_n24332));
  nand_5 g21984(.A(new_n24332), .B(new_n24287), .Y(n8031));
  not_8  g21985(.A(new_n19740), .Y(new_n24334));
  nor_5  g21986(.A(new_n19774), .B(new_n24334), .Y(new_n24335));
  nand_5 g21987(.A(new_n19738), .B(new_n19736_1), .Y(new_n24336));
  nor_5  g21988(.A(new_n24336), .B(new_n24335), .Y(new_n24337));
  not_8  g21989(.A(new_n19794), .Y(new_n24338));
  nor_5  g21990(.A(new_n19801), .B(new_n24338), .Y(new_n24339));
  nand_5 g21991(.A(new_n19792_1), .B(new_n19790), .Y(new_n24340));
  nor_5  g21992(.A(new_n24340), .B(new_n24339), .Y(new_n24341));
  nand_5 g21993(.A(new_n24341), .B(new_n22483), .Y(new_n24342_1));
  not_8  g21994(.A(new_n24342_1), .Y(new_n24343));
  nand_5 g21995(.A(new_n19831), .B(new_n19803_1), .Y(new_n24344));
  nand_5 g21996(.A(new_n24344), .B(new_n19805), .Y(new_n24345_1));
  nor_5  g21997(.A(new_n24341), .B(new_n22483), .Y(new_n24346));
  not_8  g21998(.A(new_n24346), .Y(new_n24347_1));
  nand_5 g21999(.A(new_n24347_1), .B(new_n24342_1), .Y(new_n24348));
  not_8  g22000(.A(new_n24348), .Y(new_n24349));
  and_5  g22001(.A(new_n24349), .B(new_n24345_1), .Y(new_n24350));
  nor_5  g22002(.A(new_n24350), .B(new_n24343), .Y(new_n24351));
  not_8  g22003(.A(new_n24351), .Y(new_n24352));
  nor_5  g22004(.A(new_n24352), .B(new_n24337), .Y(new_n24353));
  xor_4  g22005(.A(new_n24351), .B(new_n24337), .Y(new_n24354));
  not_8  g22006(.A(new_n24337), .Y(new_n24355));
  nor_5  g22007(.A(new_n24349), .B(new_n24345_1), .Y(new_n24356));
  or_5   g22008(.A(new_n24356), .B(new_n24350), .Y(new_n24357));
  not_8  g22009(.A(new_n24357), .Y(new_n24358));
  nand_5 g22010(.A(new_n24358), .B(new_n24355), .Y(new_n24359));
  nand_5 g22011(.A(new_n24357), .B(new_n24337), .Y(new_n24360));
  nand_5 g22012(.A(new_n19901), .B(new_n19833), .Y(new_n24361));
  nand_5 g22013(.A(new_n24361), .B(new_n19836), .Y(new_n24362));
  nand_5 g22014(.A(new_n24362), .B(new_n24360), .Y(new_n24363));
  nand_5 g22015(.A(new_n24363), .B(new_n24359), .Y(new_n24364));
  nor_5  g22016(.A(new_n24364), .B(new_n24354), .Y(new_n24365));
  nor_5  g22017(.A(new_n24365), .B(new_n24353), .Y(n8042));
  nand_5 g22018(.A(new_n11621), .B(new_n11524), .Y(new_n24367));
  nand_5 g22019(.A(new_n24367), .B(new_n11523), .Y(n8095));
  nand_5 g22020(.A(n23166), .B(new_n12402), .Y(new_n24369));
  nand_5 g22021(.A(new_n10468), .B(n4306), .Y(new_n24370));
  nand_5 g22022(.A(n10577), .B(new_n10454), .Y(new_n24371));
  nand_5 g22023(.A(new_n10473), .B(n3279), .Y(new_n24372));
  nand_5 g22024(.A(new_n12382), .B(n6381), .Y(new_n24373_1));
  nand_5 g22025(.A(n13914), .B(new_n10476), .Y(new_n24374_1));
  nand_5 g22026(.A(new_n22203), .B(new_n22201_1), .Y(new_n24375));
  nand_5 g22027(.A(new_n24375), .B(new_n22202), .Y(new_n24376));
  nand_5 g22028(.A(new_n24376), .B(new_n24374_1), .Y(new_n24377));
  nand_5 g22029(.A(new_n24377), .B(new_n24373_1), .Y(new_n24378));
  nand_5 g22030(.A(new_n24378), .B(new_n24372), .Y(new_n24379));
  nand_5 g22031(.A(new_n24379), .B(new_n24371), .Y(new_n24380));
  nand_5 g22032(.A(new_n24380), .B(new_n24370), .Y(new_n24381));
  nand_5 g22033(.A(new_n24381), .B(new_n24369), .Y(new_n24382));
  nor_5  g22034(.A(new_n24382), .B(new_n10313), .Y(new_n24383));
  not_8  g22035(.A(new_n24382), .Y(new_n24384));
  nor_5  g22036(.A(new_n24384), .B(new_n10312), .Y(new_n24385));
  or_5   g22037(.A(new_n24385), .B(new_n24383), .Y(new_n24386));
  nand_5 g22038(.A(new_n24370), .B(new_n24369), .Y(new_n24387));
  xor_4  g22039(.A(new_n24387), .B(new_n24380), .Y(new_n24388));
  nand_5 g22040(.A(new_n24388), .B(new_n10366), .Y(new_n24389));
  or_5   g22041(.A(new_n24388), .B(new_n10366), .Y(new_n24390));
  nand_5 g22042(.A(new_n24372), .B(new_n24371), .Y(new_n24391));
  xor_4  g22043(.A(new_n24391), .B(new_n24378), .Y(new_n24392));
  nand_5 g22044(.A(new_n24392), .B(new_n10373), .Y(new_n24393));
  or_5   g22045(.A(new_n24392), .B(new_n10373), .Y(new_n24394));
  nand_5 g22046(.A(new_n24374_1), .B(new_n24373_1), .Y(new_n24395));
  xor_4  g22047(.A(new_n24395), .B(new_n24376), .Y(new_n24396));
  nand_5 g22048(.A(new_n24396), .B(new_n10380), .Y(new_n24397));
  or_5   g22049(.A(new_n24396), .B(new_n10380), .Y(new_n24398));
  nand_5 g22050(.A(new_n22207), .B(new_n22199), .Y(new_n24399));
  nand_5 g22051(.A(new_n24399), .B(new_n22206), .Y(new_n24400));
  nand_5 g22052(.A(new_n24400), .B(new_n24398), .Y(new_n24401));
  nand_5 g22053(.A(new_n24401), .B(new_n24397), .Y(new_n24402));
  nand_5 g22054(.A(new_n24402), .B(new_n24394), .Y(new_n24403));
  nand_5 g22055(.A(new_n24403), .B(new_n24393), .Y(new_n24404));
  nand_5 g22056(.A(new_n24404), .B(new_n24390), .Y(new_n24405));
  nand_5 g22057(.A(new_n24405), .B(new_n24389), .Y(new_n24406_1));
  xor_4  g22058(.A(new_n24406_1), .B(new_n24386), .Y(n8103));
  nand_5 g22059(.A(new_n21464), .B(new_n21465), .Y(new_n24408));
  xnor_4 g22060(.A(new_n24408), .B(new_n21475), .Y(n8109));
  nand_5 g22061(.A(new_n22016_1), .B(new_n22014), .Y(new_n24410));
  nand_5 g22062(.A(new_n24410), .B(new_n22017), .Y(n8127));
  nand_5 g22063(.A(new_n19205), .B(new_n19204), .Y(new_n24412));
  xnor_4 g22064(.A(new_n24412), .B(new_n19207), .Y(n8130));
  nand_5 g22065(.A(new_n7991), .B(n4319), .Y(new_n24414));
  nand_5 g22066(.A(n8856), .B(new_n3313), .Y(new_n24415_1));
  nand_5 g22067(.A(n23463), .B(new_n3849), .Y(new_n24416));
  nand_5 g22068(.A(new_n3318), .B(n14130), .Y(new_n24417));
  nand_5 g22069(.A(new_n7998), .B(n13074), .Y(new_n24418));
  nand_5 g22070(.A(n16482), .B(new_n3321), .Y(new_n24419));
  nand_5 g22071(.A(new_n2602_1), .B(new_n2597), .Y(new_n24420));
  nand_5 g22072(.A(new_n24420), .B(new_n2600), .Y(new_n24421_1));
  nand_5 g22073(.A(new_n24421_1), .B(new_n24419), .Y(new_n24422));
  nand_5 g22074(.A(new_n24422), .B(new_n24418), .Y(new_n24423));
  nand_5 g22075(.A(new_n24423), .B(new_n24417), .Y(new_n24424));
  nand_5 g22076(.A(new_n24424), .B(new_n24416), .Y(new_n24425));
  nand_5 g22077(.A(new_n24425), .B(new_n24415_1), .Y(new_n24426));
  nand_5 g22078(.A(new_n24426), .B(new_n24414), .Y(new_n24427));
  nor_5  g22079(.A(new_n24427), .B(new_n8646), .Y(new_n24428));
  not_8  g22080(.A(new_n24427), .Y(new_n24429));
  nor_5  g22081(.A(new_n24429), .B(new_n8686), .Y(new_n24430));
  nor_5  g22082(.A(new_n24430), .B(new_n24428), .Y(new_n24431_1));
  nor_5  g22083(.A(new_n24427), .B(new_n8691), .Y(new_n24432));
  nor_5  g22084(.A(new_n24429), .B(new_n8693), .Y(new_n24433));
  nand_5 g22085(.A(new_n24415_1), .B(new_n24414), .Y(new_n24434));
  xor_4  g22086(.A(new_n24434), .B(new_n24425), .Y(new_n24435));
  nand_5 g22087(.A(new_n24435), .B(new_n8698), .Y(new_n24436));
  or_5   g22088(.A(new_n24435), .B(new_n8698), .Y(new_n24437));
  nand_5 g22089(.A(new_n24417), .B(new_n24416), .Y(new_n24438));
  xor_4  g22090(.A(new_n24438), .B(new_n24423), .Y(new_n24439));
  nand_5 g22091(.A(new_n24439), .B(new_n8704), .Y(new_n24440));
  or_5   g22092(.A(new_n24439), .B(new_n8704), .Y(new_n24441));
  nand_5 g22093(.A(new_n24419), .B(new_n24418), .Y(new_n24442));
  xor_4  g22094(.A(new_n24442), .B(new_n24421_1), .Y(new_n24443));
  nand_5 g22095(.A(new_n24443), .B(new_n8710), .Y(new_n24444));
  not_8  g22096(.A(new_n24444), .Y(new_n24445));
  nor_5  g22097(.A(new_n24443), .B(new_n8710), .Y(new_n24446));
  nor_5  g22098(.A(new_n2608), .B(new_n2565), .Y(new_n24447));
  nor_5  g22099(.A(new_n24447), .B(new_n2606), .Y(new_n24448));
  nor_5  g22100(.A(new_n24448), .B(new_n24446), .Y(new_n24449));
  nor_5  g22101(.A(new_n24449), .B(new_n24445), .Y(new_n24450));
  not_8  g22102(.A(new_n24450), .Y(new_n24451));
  nand_5 g22103(.A(new_n24451), .B(new_n24441), .Y(new_n24452));
  nand_5 g22104(.A(new_n24452), .B(new_n24440), .Y(new_n24453));
  nand_5 g22105(.A(new_n24453), .B(new_n24437), .Y(new_n24454));
  nand_5 g22106(.A(new_n24454), .B(new_n24436), .Y(new_n24455));
  nor_5  g22107(.A(new_n24455), .B(new_n24433), .Y(new_n24456));
  nor_5  g22108(.A(new_n24456), .B(new_n24432), .Y(new_n24457));
  xor_4  g22109(.A(new_n24457), .B(new_n24431_1), .Y(n8135));
  nand_5 g22110(.A(new_n8738), .B(new_n8737), .Y(new_n24459));
  xor_4  g22111(.A(new_n24459), .B(new_n2553_1), .Y(n8139));
  nand_5 g22112(.A(new_n20827), .B(new_n20822), .Y(new_n24461));
  nand_5 g22113(.A(new_n24461), .B(new_n20826_1), .Y(new_n24462));
  nor_5  g22114(.A(new_n20823), .B(n26660), .Y(new_n24463));
  not_8  g22115(.A(new_n24463), .Y(new_n24464));
  nand_5 g22116(.A(new_n20823), .B(n26660), .Y(new_n24465));
  and_5  g22117(.A(new_n24465), .B(new_n24464), .Y(new_n24466));
  or_5   g22118(.A(new_n24466), .B(new_n3121), .Y(new_n24467));
  nand_5 g22119(.A(new_n24466), .B(new_n3121), .Y(new_n24468));
  nand_5 g22120(.A(new_n24468), .B(new_n24467), .Y(new_n24469));
  xor_4  g22121(.A(new_n24469), .B(new_n24462), .Y(new_n24470));
  or_5   g22122(.A(new_n24470), .B(new_n7902), .Y(new_n24471));
  nand_5 g22123(.A(new_n24470), .B(new_n7902), .Y(new_n24472_1));
  not_8  g22124(.A(new_n20820), .Y(new_n24473));
  nor_5  g22125(.A(new_n20832), .B(new_n24473), .Y(new_n24474));
  nor_5  g22126(.A(new_n24474), .B(new_n20831), .Y(new_n24475));
  nand_5 g22127(.A(new_n24475), .B(new_n24472_1), .Y(new_n24476_1));
  nand_5 g22128(.A(new_n24476_1), .B(new_n24471), .Y(new_n24477));
  nand_5 g22129(.A(new_n24468), .B(new_n24462), .Y(new_n24478));
  nand_5 g22130(.A(new_n24478), .B(new_n24467), .Y(new_n24479));
  nand_5 g22131(.A(new_n24463), .B(new_n2568), .Y(new_n24480));
  nand_5 g22132(.A(new_n24464), .B(n13783), .Y(new_n24481));
  and_5  g22133(.A(new_n24481), .B(new_n24480), .Y(new_n24482));
  or_5   g22134(.A(new_n24482), .B(new_n3112), .Y(new_n24483_1));
  nand_5 g22135(.A(new_n24482), .B(new_n3112), .Y(new_n24484));
  nand_5 g22136(.A(new_n24484), .B(new_n24483_1), .Y(new_n24485_1));
  xor_4  g22137(.A(new_n24485_1), .B(new_n24479), .Y(new_n24486));
  or_5   g22138(.A(new_n24486), .B(new_n7895), .Y(new_n24487));
  nand_5 g22139(.A(new_n24486), .B(new_n7895), .Y(new_n24488));
  nand_5 g22140(.A(new_n24488), .B(new_n24487), .Y(new_n24489));
  xor_4  g22141(.A(new_n24489), .B(new_n24477), .Y(n8148));
  nand_5 g22142(.A(new_n20088), .B(new_n20087), .Y(new_n24491));
  xor_4  g22143(.A(new_n24491), .B(new_n20107), .Y(n8149));
  nand_5 g22144(.A(new_n4250), .B(new_n4249), .Y(new_n24493));
  xnor_4 g22145(.A(new_n24493), .B(new_n4270), .Y(n8159));
  xor_4  g22146(.A(new_n13470), .B(new_n2635), .Y(n8179));
  nand_5 g22147(.A(new_n16984), .B(new_n16985), .Y(new_n24496));
  xor_4  g22148(.A(new_n24496), .B(new_n16987), .Y(n8215));
  nand_5 g22149(.A(new_n21466), .B(new_n21467), .Y(new_n24498));
  xnor_4 g22150(.A(new_n24498), .B(new_n21473), .Y(n8267));
  nand_5 g22151(.A(new_n22661), .B(new_n22660_1), .Y(new_n24500));
  xor_4  g22152(.A(new_n24500), .B(new_n20380), .Y(n8276));
  nor_5  g22153(.A(new_n24480), .B(n1654), .Y(new_n24502));
  nand_5 g22154(.A(new_n24502), .B(new_n8574), .Y(new_n24503));
  nor_5  g22155(.A(new_n24503), .B(n22626), .Y(new_n24504));
  nand_5 g22156(.A(new_n24504), .B(new_n17214), .Y(new_n24505));
  not_8  g22157(.A(new_n24504), .Y(new_n24506));
  nand_5 g22158(.A(new_n24503), .B(n22626), .Y(new_n24507));
  and_5  g22159(.A(new_n24507), .B(new_n24506), .Y(new_n24508));
  or_5   g22160(.A(new_n24508), .B(new_n17219_1), .Y(new_n24509));
  nand_5 g22161(.A(new_n24508), .B(new_n17219_1), .Y(new_n24510));
  xor_4  g22162(.A(new_n24502), .B(new_n8574), .Y(new_n24511));
  or_5   g22163(.A(new_n24511), .B(new_n3303), .Y(new_n24512_1));
  nand_5 g22164(.A(new_n24511), .B(new_n3303), .Y(new_n24513));
  xor_4  g22165(.A(new_n24480), .B(n1654), .Y(new_n24514));
  or_5   g22166(.A(new_n24514), .B(new_n3199), .Y(new_n24515));
  nand_5 g22167(.A(new_n24514), .B(new_n3199), .Y(new_n24516));
  nand_5 g22168(.A(new_n24484), .B(new_n24479), .Y(new_n24517));
  nand_5 g22169(.A(new_n24517), .B(new_n24483_1), .Y(new_n24518));
  nand_5 g22170(.A(new_n24518), .B(new_n24516), .Y(new_n24519));
  nand_5 g22171(.A(new_n24519), .B(new_n24515), .Y(new_n24520));
  nand_5 g22172(.A(new_n24520), .B(new_n24513), .Y(new_n24521));
  nand_5 g22173(.A(new_n24521), .B(new_n24512_1), .Y(new_n24522));
  nand_5 g22174(.A(new_n24522), .B(new_n24510), .Y(new_n24523));
  nand_5 g22175(.A(new_n24523), .B(new_n24509), .Y(new_n24524));
  nor_5  g22176(.A(new_n24524), .B(new_n24505), .Y(new_n24525));
  not_8  g22177(.A(new_n24524), .Y(new_n24526));
  nand_5 g22178(.A(new_n24506), .B(new_n17239), .Y(new_n24527));
  nor_5  g22179(.A(new_n24527), .B(new_n24526), .Y(new_n24528));
  nor_5  g22180(.A(new_n24528), .B(new_n24525), .Y(new_n24529));
  and_5  g22181(.A(new_n24527), .B(new_n24505), .Y(new_n24530));
  xor_4  g22182(.A(new_n24530), .B(new_n24524), .Y(new_n24531));
  not_8  g22183(.A(new_n24531), .Y(new_n24532));
  nand_5 g22184(.A(new_n24532), .B(new_n23763), .Y(new_n24533));
  nand_5 g22185(.A(new_n24510), .B(new_n24509), .Y(new_n24534));
  xor_4  g22186(.A(new_n24534), .B(new_n24522), .Y(new_n24535));
  nand_5 g22187(.A(new_n24535), .B(new_n19647), .Y(new_n24536));
  or_5   g22188(.A(new_n24535), .B(new_n19647), .Y(new_n24537));
  nand_5 g22189(.A(new_n24513), .B(new_n24512_1), .Y(new_n24538));
  xor_4  g22190(.A(new_n24538), .B(new_n24520), .Y(new_n24539));
  nand_5 g22191(.A(new_n24539), .B(new_n7968_1), .Y(new_n24540));
  nor_5  g22192(.A(new_n24539), .B(new_n7968_1), .Y(new_n24541));
  not_8  g22193(.A(new_n24541), .Y(new_n24542));
  nand_5 g22194(.A(new_n24516), .B(new_n24515), .Y(new_n24543));
  xor_4  g22195(.A(new_n24543), .B(new_n24518), .Y(new_n24544));
  nand_5 g22196(.A(new_n24544), .B(new_n7818), .Y(new_n24545));
  nor_5  g22197(.A(new_n24544), .B(new_n7818), .Y(new_n24546));
  nand_5 g22198(.A(new_n24488), .B(new_n24477), .Y(new_n24547));
  nand_5 g22199(.A(new_n24547), .B(new_n24487), .Y(new_n24548));
  or_5   g22200(.A(new_n24548), .B(new_n24546), .Y(new_n24549));
  nand_5 g22201(.A(new_n24549), .B(new_n24545), .Y(new_n24550));
  nand_5 g22202(.A(new_n24550), .B(new_n24542), .Y(new_n24551));
  nand_5 g22203(.A(new_n24551), .B(new_n24540), .Y(new_n24552));
  nand_5 g22204(.A(new_n24552), .B(new_n24537), .Y(new_n24553));
  nand_5 g22205(.A(new_n24553), .B(new_n24536), .Y(new_n24554));
  nand_5 g22206(.A(new_n24554), .B(new_n24533), .Y(new_n24555));
  nand_5 g22207(.A(new_n24531), .B(new_n19638), .Y(new_n24556));
  and_5  g22208(.A(new_n24556), .B(new_n19630), .Y(new_n24557));
  nand_5 g22209(.A(new_n24557), .B(new_n24555), .Y(new_n24558_1));
  nand_5 g22210(.A(new_n24558_1), .B(new_n24529), .Y(new_n24559));
  or_5   g22211(.A(new_n24555), .B(new_n19630), .Y(new_n24560));
  nand_5 g22212(.A(new_n24560), .B(new_n24559), .Y(new_n24561));
  nor_5  g22213(.A(new_n24561), .B(new_n24525), .Y(n8288));
  nor_5  g22214(.A(new_n12960), .B(new_n12958), .Y(new_n24563));
  nor_5  g22215(.A(new_n24563), .B(new_n12962), .Y(n8306));
  nand_5 g22216(.A(new_n9033), .B(new_n9032_1), .Y(new_n24565));
  xor_4  g22217(.A(new_n24565), .B(new_n9096), .Y(n8320));
  nand_5 g22218(.A(new_n14289), .B(new_n14287), .Y(new_n24567));
  xor_4  g22219(.A(new_n24567), .B(new_n14313), .Y(n8321));
  nand_5 g22220(.A(new_n18715), .B(new_n18714), .Y(new_n24569));
  xnor_4 g22221(.A(new_n24569), .B(new_n18729), .Y(n8339));
  nand_5 g22222(.A(new_n10384), .B(new_n10383), .Y(new_n24571));
  xor_4  g22223(.A(new_n24571), .B(new_n10446), .Y(n8376));
  xor_4  g22224(.A(new_n21843), .B(new_n11805), .Y(n8408));
  xor_4  g22225(.A(new_n16414), .B(new_n16412), .Y(n8417));
  nand_5 g22226(.A(new_n14770), .B(new_n14769), .Y(new_n24575));
  xor_4  g22227(.A(new_n24575), .B(new_n14786), .Y(n8432));
  nor_5  g22228(.A(new_n11834), .B(new_n11746), .Y(new_n24577));
  nor_5  g22229(.A(new_n24577), .B(new_n11744), .Y(new_n24578));
  nand_5 g22230(.A(new_n11691), .B(new_n11641), .Y(new_n24579_1));
  nand_5 g22231(.A(new_n24579_1), .B(new_n11643), .Y(new_n24580));
  not_8  g22232(.A(new_n24580), .Y(new_n24581));
  nor_5  g22233(.A(new_n24581), .B(new_n11745), .Y(new_n24582));
  nor_5  g22234(.A(new_n24582), .B(new_n24578), .Y(new_n24583));
  nor_5  g22235(.A(new_n24580), .B(new_n11743), .Y(new_n24584));
  nor_5  g22236(.A(new_n24584), .B(new_n24577), .Y(new_n24585));
  nor_5  g22237(.A(new_n24585), .B(new_n24583), .Y(n8453));
  xor_4  g22238(.A(new_n17859), .B(new_n15655), .Y(n8480));
  nand_5 g22239(.A(new_n18893), .B(new_n18892), .Y(new_n24588));
  xnor_4 g22240(.A(new_n24588), .B(new_n18913), .Y(n8489));
  nand_5 g22241(.A(new_n24437), .B(new_n24436), .Y(new_n24590));
  xor_4  g22242(.A(new_n24590), .B(new_n24453), .Y(n8505));
  nand_5 g22243(.A(new_n22299), .B(new_n22302), .Y(new_n24592));
  xor_4  g22244(.A(new_n24592), .B(new_n22321), .Y(n8510));
  xor_4  g22245(.A(new_n13957), .B(new_n9906), .Y(n8519));
  nand_5 g22246(.A(new_n11205), .B(new_n11206), .Y(new_n24595));
  xor_4  g22247(.A(new_n24595), .B(new_n11210), .Y(n8535));
  nand_5 g22248(.A(new_n22002), .B(new_n22001), .Y(new_n24597));
  xor_4  g22249(.A(new_n24597), .B(new_n22005), .Y(n8550));
  nand_5 g22250(.A(new_n23316), .B(new_n23317), .Y(new_n24599));
  xnor_4 g22251(.A(new_n24599), .B(new_n23324), .Y(n8563));
  nand_5 g22252(.A(new_n15262), .B(new_n15263), .Y(new_n24601));
  xor_4  g22253(.A(new_n24601), .B(new_n15266), .Y(n8594));
  nand_5 g22254(.A(new_n7920), .B(new_n7919), .Y(new_n24603));
  xnor_4 g22255(.A(new_n24603), .B(new_n7942), .Y(n8608));
  xor_4  g22256(.A(new_n5112), .B(new_n5110), .Y(n8620));
  nand_5 g22257(.A(new_n8490), .B(new_n8489_1), .Y(new_n24606));
  xnor_4 g22258(.A(new_n24606), .B(new_n8559), .Y(n8637));
  not_8  g22259(.A(new_n19661), .Y(new_n24608));
  nand_5 g22260(.A(new_n24608), .B(new_n19660), .Y(new_n24609));
  xor_4  g22261(.A(new_n24609), .B(new_n19664_1), .Y(n8662));
  nor_5  g22262(.A(new_n21513), .B(new_n21512), .Y(new_n24611));
  xor_4  g22263(.A(new_n24611), .B(new_n21522), .Y(n8716));
  nand_5 g22264(.A(new_n9041), .B(new_n9040), .Y(new_n24613));
  xor_4  g22265(.A(new_n24613), .B(new_n9094), .Y(n8744));
  nand_5 g22266(.A(new_n24121), .B(new_n24119_1), .Y(new_n24615));
  nand_5 g22267(.A(new_n24615), .B(new_n24120), .Y(new_n24616));
  not_8  g22268(.A(new_n24616), .Y(new_n24617));
  nor_5  g22269(.A(new_n24617), .B(new_n20361), .Y(new_n24618_1));
  not_8  g22270(.A(new_n24618_1), .Y(new_n24619));
  nand_5 g22271(.A(new_n24617), .B(new_n20361), .Y(new_n24620_1));
  and_5  g22272(.A(new_n24620_1), .B(new_n24619), .Y(new_n24621));
  nand_5 g22273(.A(new_n24234), .B(new_n24227), .Y(new_n24622));
  nand_5 g22274(.A(new_n24622), .B(new_n24226), .Y(new_n24623));
  nand_5 g22275(.A(new_n24623), .B(new_n17553), .Y(new_n24624));
  or_5   g22276(.A(new_n24623), .B(new_n17553), .Y(new_n24625));
  and_5  g22277(.A(new_n24625), .B(new_n24624), .Y(new_n24626_1));
  not_8  g22278(.A(new_n24626_1), .Y(new_n24627));
  nand_5 g22279(.A(new_n24627), .B(new_n24621), .Y(new_n24628));
  not_8  g22280(.A(new_n24621), .Y(new_n24629_1));
  nand_5 g22281(.A(new_n24626_1), .B(new_n24629_1), .Y(new_n24630));
  nand_5 g22282(.A(new_n24630), .B(new_n24628), .Y(new_n24631));
  nand_5 g22283(.A(new_n24237), .B(new_n24123), .Y(new_n24632));
  nand_5 g22284(.A(new_n24235), .B(new_n24124), .Y(new_n24633));
  nand_5 g22285(.A(new_n24242), .B(new_n18567), .Y(new_n24634));
  nand_5 g22286(.A(new_n24241), .B(new_n18568), .Y(new_n24635));
  nand_5 g22287(.A(new_n19948), .B(new_n19941_1), .Y(new_n24636_1));
  nand_5 g22288(.A(new_n24636_1), .B(new_n19950), .Y(new_n24637));
  nand_5 g22289(.A(new_n24637), .B(new_n24635), .Y(new_n24638_1));
  nand_5 g22290(.A(new_n24638_1), .B(new_n24634), .Y(new_n24639));
  nand_5 g22291(.A(new_n24639), .B(new_n24633), .Y(new_n24640));
  nand_5 g22292(.A(new_n24640), .B(new_n24632), .Y(new_n24641));
  xor_4  g22293(.A(new_n24641), .B(new_n24631), .Y(n8803));
  nand_5 g22294(.A(new_n23154), .B(new_n23134), .Y(new_n24643));
  nand_5 g22295(.A(new_n24643), .B(new_n23135), .Y(new_n24644));
  xor_4  g22296(.A(new_n24644), .B(new_n23131), .Y(new_n24645));
  nand_5 g22297(.A(new_n18120), .B(new_n18100), .Y(new_n24646));
  nand_5 g22298(.A(new_n24646), .B(new_n18101), .Y(new_n24647));
  nand_5 g22299(.A(new_n24647), .B(new_n24645), .Y(new_n24648));
  or_5   g22300(.A(new_n24647), .B(new_n24645), .Y(new_n24649));
  and_5  g22301(.A(new_n24649), .B(new_n24648), .Y(new_n24650));
  nand_5 g22302(.A(new_n23178), .B(new_n23157), .Y(new_n24651));
  nand_5 g22303(.A(new_n24651), .B(new_n23156), .Y(new_n24652));
  xor_4  g22304(.A(new_n24652), .B(new_n24650), .Y(new_n24653));
  not_8  g22305(.A(new_n24653), .Y(new_n24654));
  nand_5 g22306(.A(new_n24654), .B(new_n8841), .Y(new_n24655));
  nand_5 g22307(.A(new_n24653), .B(new_n8840), .Y(new_n24656));
  nand_5 g22308(.A(new_n24656), .B(new_n24655), .Y(new_n24657));
  nand_5 g22309(.A(new_n23860), .B(new_n23825), .Y(new_n24658));
  nand_5 g22310(.A(new_n24658), .B(new_n23826), .Y(new_n24659));
  not_8  g22311(.A(new_n24659), .Y(new_n24660));
  xor_4  g22312(.A(new_n24660), .B(new_n24657), .Y(n8809));
  nand_5 g22313(.A(new_n24137), .B(new_n24125), .Y(new_n24662));
  nand_5 g22314(.A(new_n24662), .B(new_n24126), .Y(new_n24663));
  nor_5  g22315(.A(new_n24663), .B(new_n20730), .Y(new_n24664));
  or_5   g22316(.A(new_n24664), .B(new_n24619), .Y(new_n24665));
  nand_5 g22317(.A(new_n24664), .B(new_n24619), .Y(new_n24666));
  nand_5 g22318(.A(new_n24666), .B(new_n24665), .Y(new_n24667));
  xor_4  g22319(.A(new_n24663), .B(new_n20730), .Y(new_n24668));
  or_5   g22320(.A(new_n24668), .B(new_n24629_1), .Y(new_n24669));
  nand_5 g22321(.A(new_n24668), .B(new_n24629_1), .Y(new_n24670));
  nand_5 g22322(.A(new_n24155_1), .B(new_n24139), .Y(new_n24671));
  nand_5 g22323(.A(new_n24671), .B(new_n24140), .Y(new_n24672));
  nand_5 g22324(.A(new_n24672), .B(new_n24670), .Y(new_n24673));
  nand_5 g22325(.A(new_n24673), .B(new_n24669), .Y(new_n24674));
  xor_4  g22326(.A(new_n24674), .B(new_n24667), .Y(n8821));
  nand_5 g22327(.A(new_n17808), .B(new_n17806), .Y(new_n24676));
  xor_4  g22328(.A(new_n24676), .B(new_n17824), .Y(n8824));
  nand_5 g22329(.A(new_n20305), .B(new_n20306), .Y(new_n24678));
  xor_4  g22330(.A(new_n24678), .B(new_n20308), .Y(n8849));
  nand_5 g22331(.A(new_n15788), .B(new_n15787), .Y(new_n24680));
  xor_4  g22332(.A(new_n24680), .B(new_n15798), .Y(n8861));
  not_8  g22333(.A(new_n22934), .Y(new_n24682));
  not_8  g22334(.A(new_n22935), .Y(new_n24683));
  nor_5  g22335(.A(new_n24683), .B(new_n22933), .Y(new_n24684));
  nor_5  g22336(.A(new_n24684), .B(new_n24682), .Y(new_n24685));
  nand_5 g22337(.A(n3324), .B(n2272), .Y(new_n24686));
  nand_5 g22338(.A(new_n18124), .B(new_n8142), .Y(new_n24687));
  nand_5 g22339(.A(new_n24687), .B(new_n24686), .Y(new_n24688));
  xor_4  g22340(.A(new_n24688), .B(new_n24685), .Y(new_n24689));
  or_5   g22341(.A(new_n24689), .B(new_n8615), .Y(new_n24690));
  nand_5 g22342(.A(new_n24689), .B(new_n8615), .Y(new_n24691));
  nand_5 g22343(.A(new_n24691), .B(new_n24690), .Y(new_n24692));
  nand_5 g22344(.A(new_n22939_1), .B(new_n22929), .Y(new_n24693));
  nand_5 g22345(.A(new_n24693), .B(new_n22938), .Y(new_n24694));
  xor_4  g22346(.A(new_n24694), .B(new_n24692), .Y(new_n24695));
  not_8  g22347(.A(new_n24695), .Y(new_n24696));
  nand_5 g22348(.A(n22442), .B(new_n7991), .Y(new_n24697));
  nand_5 g22349(.A(new_n8016), .B(n8856), .Y(new_n24698));
  nand_5 g22350(.A(new_n24698), .B(new_n24697), .Y(new_n24699));
  nand_5 g22351(.A(new_n22946), .B(new_n22944), .Y(new_n24700));
  nand_5 g22352(.A(new_n24700), .B(new_n22945), .Y(new_n24701));
  xnor_4 g22353(.A(new_n24701), .B(new_n24699), .Y(new_n24702));
  nand_5 g22354(.A(new_n24702), .B(new_n24696), .Y(new_n24703));
  not_8  g22355(.A(new_n24703), .Y(new_n24704));
  nor_5  g22356(.A(new_n24702), .B(new_n24696), .Y(new_n24705));
  or_5   g22357(.A(new_n24705), .B(new_n24704), .Y(new_n24706));
  not_8  g22358(.A(new_n22927), .Y(new_n24707));
  nor_5  g22359(.A(new_n22951), .B(new_n24707), .Y(new_n24708));
  nor_5  g22360(.A(new_n24708), .B(new_n22950), .Y(new_n24709));
  xor_4  g22361(.A(new_n24709), .B(new_n24706), .Y(n8862));
  nand_5 g22362(.A(new_n15645), .B(new_n15644), .Y(new_n24711));
  xnor_4 g22363(.A(new_n24711), .B(new_n15658), .Y(n8884));
  xor_4  g22364(.A(new_n21716), .B(new_n21715), .Y(n8909));
  nand_5 g22365(.A(new_n13431), .B(new_n13430), .Y(new_n24714));
  xor_4  g22366(.A(new_n24714), .B(new_n13485), .Y(n8911));
  nand_5 g22367(.A(new_n12823), .B(new_n12821_1), .Y(new_n24716));
  xor_4  g22368(.A(new_n24716), .B(new_n12889), .Y(n8971));
  or_5   g22369(.A(new_n24297_1), .B(new_n24296), .Y(new_n24718));
  xor_4  g22370(.A(new_n24718), .B(new_n24327_1), .Y(n8982));
  nand_5 g22371(.A(new_n6099), .B(new_n6098), .Y(new_n24720));
  xor_4  g22372(.A(new_n24720), .B(new_n6122), .Y(n8993));
  nand_5 g22373(.A(new_n16394), .B(new_n16392), .Y(new_n24722));
  xnor_4 g22374(.A(new_n24722), .B(new_n16429), .Y(n9012));
  nand_5 g22375(.A(new_n23064), .B(new_n22976), .Y(new_n24724));
  nand_5 g22376(.A(new_n23065_1), .B(new_n22975), .Y(new_n24725));
  nand_5 g22377(.A(new_n24725), .B(new_n24724), .Y(new_n24726));
  nor_5  g22378(.A(new_n23124), .B(new_n23069), .Y(new_n24727));
  nor_5  g22379(.A(new_n24727), .B(new_n23068_1), .Y(new_n24728));
  xnor_4 g22380(.A(new_n24728), .B(new_n24726), .Y(n9032));
  nand_5 g22381(.A(new_n18406), .B(new_n18405_1), .Y(new_n24730));
  xnor_4 g22382(.A(new_n24730), .B(new_n18409_1), .Y(n9042));
  nand_5 g22383(.A(new_n19861), .B(new_n19860), .Y(new_n24732_1));
  xor_4  g22384(.A(new_n24732_1), .B(new_n19895), .Y(n9046));
  nand_5 g22385(.A(new_n9356), .B(new_n9355), .Y(new_n24734));
  xnor_4 g22386(.A(new_n24734), .B(new_n9421), .Y(n9047));
  nand_5 g22387(.A(new_n17480), .B(new_n17481), .Y(new_n24736));
  xor_4  g22388(.A(new_n24736), .B(new_n17483), .Y(n9104));
  nand_5 g22389(.A(new_n23483), .B(new_n23479), .Y(new_n24738));
  nand_5 g22390(.A(new_n24738), .B(new_n23485), .Y(new_n24739));
  xor_4  g22391(.A(new_n24739), .B(new_n23484), .Y(new_n24740));
  xor_4  g22392(.A(new_n24740), .B(new_n22259), .Y(new_n24741));
  nand_5 g22393(.A(new_n23499), .B(new_n23489), .Y(new_n24742));
  nand_5 g22394(.A(new_n24742), .B(new_n23490), .Y(new_n24743));
  xor_4  g22395(.A(new_n24743), .B(new_n24741), .Y(n9129));
  nand_5 g22396(.A(new_n21901), .B(new_n21900), .Y(new_n24745));
  xor_4  g22397(.A(new_n24745), .B(new_n21935), .Y(n9146));
  xor_4  g22398(.A(new_n9906), .B(new_n7656), .Y(n9164));
  nand_5 g22399(.A(new_n14689), .B(new_n14688), .Y(new_n24748));
  xor_4  g22400(.A(new_n24748), .B(new_n14694), .Y(n9166));
  nand_5 g22401(.A(new_n20752), .B(new_n20751), .Y(new_n24750));
  xnor_4 g22402(.A(new_n24750), .B(new_n20765), .Y(n9182));
  nand_5 g22403(.A(new_n8223), .B(new_n8222), .Y(new_n24752));
  xor_4  g22404(.A(new_n24752), .B(new_n8263), .Y(n9191));
  nand_5 g22405(.A(new_n13415), .B(new_n13416), .Y(new_n24754));
  xor_4  g22406(.A(new_n24754), .B(new_n13491), .Y(n9217));
  nand_5 g22407(.A(new_n18594), .B(new_n18595), .Y(new_n24756));
  xnor_4 g22408(.A(new_n24756), .B(new_n18621), .Y(n9220));
  nand_5 g22409(.A(new_n21918), .B(new_n21919), .Y(new_n24758_1));
  xnor_4 g22410(.A(new_n24758_1), .B(new_n21924), .Y(n9261));
  nand_5 g22411(.A(new_n8584), .B(n3324), .Y(new_n24760));
  nand_5 g22412(.A(n22626), .B(new_n18124), .Y(new_n24761));
  nand_5 g22413(.A(new_n21533), .B(new_n21530), .Y(new_n24762));
  nand_5 g22414(.A(new_n24762), .B(new_n21532), .Y(new_n24763));
  nand_5 g22415(.A(new_n24763), .B(new_n24761), .Y(new_n24764));
  nand_5 g22416(.A(new_n24764), .B(new_n24760), .Y(new_n24765));
  nand_5 g22417(.A(new_n24765), .B(new_n20743), .Y(new_n24766));
  or_5   g22418(.A(new_n24765), .B(new_n20743), .Y(new_n24767));
  nand_5 g22419(.A(new_n24767), .B(new_n24766), .Y(new_n24768_1));
  nand_5 g22420(.A(new_n24761), .B(new_n24760), .Y(new_n24769));
  xor_4  g22421(.A(new_n24769), .B(new_n24763), .Y(new_n24770));
  nand_5 g22422(.A(new_n24770), .B(new_n20757), .Y(new_n24771));
  not_8  g22423(.A(new_n24771), .Y(new_n24772));
  or_5   g22424(.A(new_n24770), .B(new_n20757), .Y(new_n24773));
  not_8  g22425(.A(new_n24773), .Y(new_n24774));
  nor_5  g22426(.A(new_n21539), .B(new_n21528), .Y(new_n24775));
  nor_5  g22427(.A(new_n24775), .B(new_n21537), .Y(new_n24776));
  nor_5  g22428(.A(new_n24776), .B(new_n24774), .Y(new_n24777));
  nor_5  g22429(.A(new_n24777), .B(new_n24772), .Y(new_n24778));
  xor_4  g22430(.A(new_n24778), .B(new_n24768_1), .Y(n9287));
  nand_5 g22431(.A(new_n16227), .B(new_n16226), .Y(new_n24780));
  xor_4  g22432(.A(new_n24780), .B(new_n16241), .Y(n9308));
  nand_5 g22433(.A(new_n5602), .B(new_n5601), .Y(new_n24782));
  xor_4  g22434(.A(new_n24782), .B(new_n5653), .Y(n9344));
  nand_5 g22435(.A(new_n4027), .B(new_n4026), .Y(new_n24784_1));
  xnor_4 g22436(.A(new_n24784_1), .B(new_n4050), .Y(n9364));
  nand_5 g22437(.A(new_n24778), .B(new_n24766), .Y(new_n24786_1));
  not_8  g22438(.A(new_n24778), .Y(new_n24787));
  nand_5 g22439(.A(new_n24787), .B(new_n24767), .Y(new_n24788));
  nand_5 g22440(.A(new_n24788), .B(new_n24786_1), .Y(new_n24789));
  xor_4  g22441(.A(new_n24765), .B(new_n20769), .Y(new_n24790));
  nor_5  g22442(.A(new_n24790), .B(new_n24789), .Y(n9371));
  xor_4  g22443(.A(new_n11807), .B(new_n11805), .Y(n9382));
  xor_4  g22444(.A(new_n24364), .B(new_n24354), .Y(n9403));
  nand_5 g22445(.A(new_n14668), .B(new_n14667), .Y(new_n24794));
  xor_4  g22446(.A(new_n24794), .B(new_n14700), .Y(n9419));
  nand_5 g22447(.A(new_n24068), .B(new_n24069), .Y(new_n24796));
  xor_4  g22448(.A(new_n24796), .B(new_n24096_1), .Y(n9423));
  nor_5  g22449(.A(new_n21508), .B(new_n21507), .Y(new_n24798));
  xor_4  g22450(.A(new_n24798), .B(new_n21524), .Y(n9430));
  nand_5 g22451(.A(new_n8798), .B(n23272), .Y(new_n24800));
  nand_5 g22452(.A(n25120), .B(new_n4850_1), .Y(new_n24801));
  nand_5 g22453(.A(new_n24801), .B(new_n24800), .Y(new_n24802));
  nand_5 g22454(.A(new_n4856), .B(n8363), .Y(new_n24803));
  nand_5 g22455(.A(n11481), .B(new_n8801), .Y(new_n24804));
  nand_5 g22456(.A(new_n18040), .B(new_n18037), .Y(new_n24805));
  nand_5 g22457(.A(new_n24805), .B(new_n18039), .Y(new_n24806));
  nand_5 g22458(.A(new_n24806), .B(new_n24804), .Y(new_n24807_1));
  nand_5 g22459(.A(new_n24807_1), .B(new_n24803), .Y(new_n24808));
  not_8  g22460(.A(new_n24808), .Y(new_n24809));
  xor_4  g22461(.A(new_n24809), .B(new_n24802), .Y(new_n24810));
  nand_5 g22462(.A(new_n24810), .B(new_n19802), .Y(new_n24811));
  not_8  g22463(.A(new_n24810), .Y(new_n24812));
  nand_5 g22464(.A(new_n24812), .B(new_n19804), .Y(new_n24813));
  nand_5 g22465(.A(new_n24813), .B(new_n24811), .Y(new_n24814));
  nand_5 g22466(.A(new_n24804), .B(new_n24803), .Y(new_n24815));
  xor_4  g22467(.A(new_n24815), .B(new_n24806), .Y(new_n24816));
  nand_5 g22468(.A(new_n24816), .B(new_n19809), .Y(new_n24817));
  not_8  g22469(.A(new_n24816), .Y(new_n24818));
  nand_5 g22470(.A(new_n24818), .B(new_n19808), .Y(new_n24819));
  nand_5 g22471(.A(new_n18045_1), .B(new_n18027), .Y(new_n24820));
  nand_5 g22472(.A(new_n24820), .B(new_n18044), .Y(new_n24821));
  nand_5 g22473(.A(new_n24821), .B(new_n24819), .Y(new_n24822));
  nand_5 g22474(.A(new_n24822), .B(new_n24817), .Y(new_n24823));
  xor_4  g22475(.A(new_n24823), .B(new_n24814), .Y(new_n24824));
  nand_5 g22476(.A(new_n24824), .B(new_n19775), .Y(new_n24825));
  not_8  g22477(.A(new_n24824), .Y(new_n24826_1));
  nand_5 g22478(.A(new_n24826_1), .B(new_n19834), .Y(new_n24827));
  nand_5 g22479(.A(new_n24827), .B(new_n24825), .Y(new_n24828));
  nand_5 g22480(.A(new_n24817), .B(new_n24819), .Y(new_n24829));
  xor_4  g22481(.A(new_n24829), .B(new_n24821), .Y(new_n24830));
  not_8  g22482(.A(new_n24830), .Y(new_n24831));
  nand_5 g22483(.A(new_n24831), .B(new_n19840), .Y(new_n24832));
  nand_5 g22484(.A(new_n24830), .B(new_n19839), .Y(new_n24833));
  nand_5 g22485(.A(new_n19848), .B(new_n18047), .Y(new_n24834));
  nand_5 g22486(.A(new_n19847), .B(new_n18049), .Y(new_n24835));
  nand_5 g22487(.A(new_n19856), .B(new_n12325_1), .Y(new_n24836));
  nand_5 g22488(.A(new_n19855), .B(new_n12327), .Y(new_n24837));
  nand_5 g22489(.A(new_n19864), .B(new_n12275), .Y(new_n24838));
  nand_5 g22490(.A(new_n19863), .B(new_n12274), .Y(new_n24839));
  nand_5 g22491(.A(new_n19871), .B(new_n12279), .Y(new_n24840_1));
  nand_5 g22492(.A(new_n19872), .B(new_n12280), .Y(new_n24841_1));
  nand_5 g22493(.A(new_n17205), .B(new_n17190), .Y(new_n24842));
  nand_5 g22494(.A(new_n24842), .B(new_n17204), .Y(new_n24843));
  nand_5 g22495(.A(new_n24843), .B(new_n24841_1), .Y(new_n24844));
  and_5  g22496(.A(new_n24844), .B(new_n24840_1), .Y(new_n24845));
  nand_5 g22497(.A(new_n24845), .B(new_n24839), .Y(new_n24846));
  nand_5 g22498(.A(new_n24846), .B(new_n24838), .Y(new_n24847));
  nand_5 g22499(.A(new_n24847), .B(new_n24837), .Y(new_n24848));
  nand_5 g22500(.A(new_n24848), .B(new_n24836), .Y(new_n24849));
  nand_5 g22501(.A(new_n24849), .B(new_n24835), .Y(new_n24850));
  nand_5 g22502(.A(new_n24850), .B(new_n24834), .Y(new_n24851));
  nand_5 g22503(.A(new_n24851), .B(new_n24833), .Y(new_n24852));
  nand_5 g22504(.A(new_n24852), .B(new_n24832), .Y(new_n24853_1));
  xor_4  g22505(.A(new_n24853_1), .B(new_n24828), .Y(n9435));
  nand_5 g22506(.A(new_n18508), .B(new_n18507), .Y(new_n24855));
  xnor_4 g22507(.A(new_n24855), .B(new_n18547), .Y(n9451));
  nand_5 g22508(.A(new_n22114), .B(new_n22090_1), .Y(new_n24857_1));
  nand_5 g22509(.A(new_n24857_1), .B(new_n22113_1), .Y(new_n24858));
  nand_5 g22510(.A(new_n22110), .B(new_n22107_1), .Y(new_n24859));
  nand_5 g22511(.A(new_n24859), .B(new_n22109), .Y(new_n24860));
  not_8  g22512(.A(new_n24860), .Y(new_n24861));
  nand_5 g22513(.A(new_n3295), .B(n10763), .Y(new_n24862));
  nand_5 g22514(.A(n12657), .B(new_n3287), .Y(new_n24863));
  nand_5 g22515(.A(new_n24863), .B(new_n24862), .Y(new_n24864));
  xor_4  g22516(.A(new_n24864), .B(new_n24861), .Y(new_n24865));
  or_5   g22517(.A(new_n24865), .B(new_n22942), .Y(new_n24866));
  nand_5 g22518(.A(new_n24865), .B(new_n22942), .Y(new_n24867));
  nand_5 g22519(.A(new_n24867), .B(new_n24866), .Y(new_n24868));
  xor_4  g22520(.A(new_n24868), .B(new_n24858), .Y(n9458));
  nand_5 g22521(.A(new_n11696), .B(n11220), .Y(new_n24870));
  nand_5 g22522(.A(n12507), .B(new_n11623), .Y(new_n24871));
  nand_5 g22523(.A(new_n17123), .B(new_n17121), .Y(new_n24872));
  nand_5 g22524(.A(new_n24872), .B(new_n17122), .Y(new_n24873));
  nand_5 g22525(.A(new_n24873), .B(new_n24871), .Y(new_n24874));
  nand_5 g22526(.A(new_n24874), .B(new_n24870), .Y(new_n24875));
  not_8  g22527(.A(new_n24875), .Y(new_n24876));
  nand_5 g22528(.A(new_n24876), .B(new_n23704), .Y(new_n24877));
  nand_5 g22529(.A(new_n24875), .B(new_n23703), .Y(new_n24878));
  nand_5 g22530(.A(new_n24878), .B(new_n24877), .Y(new_n24879_1));
  nand_5 g22531(.A(new_n24871), .B(new_n24870), .Y(new_n24880));
  xor_4  g22532(.A(new_n24880), .B(new_n24873), .Y(new_n24881));
  or_5   g22533(.A(new_n24881), .B(new_n23710), .Y(new_n24882));
  nand_5 g22534(.A(new_n24881), .B(new_n23710), .Y(new_n24883));
  not_8  g22535(.A(new_n17102), .Y(new_n24884));
  nor_5  g22536(.A(new_n17128), .B(new_n24884), .Y(new_n24885));
  nor_5  g22537(.A(new_n24885), .B(new_n17127), .Y(new_n24886));
  not_8  g22538(.A(new_n24886), .Y(new_n24887_1));
  nand_5 g22539(.A(new_n24887_1), .B(new_n24883), .Y(new_n24888));
  nand_5 g22540(.A(new_n24888), .B(new_n24882), .Y(new_n24889));
  xnor_4 g22541(.A(new_n24889), .B(new_n24879_1), .Y(n9459));
  nand_5 g22542(.A(new_n17364), .B(new_n17367), .Y(new_n24891));
  xor_4  g22543(.A(new_n24891), .B(new_n17409), .Y(n9508));
  nor_5  g22544(.A(new_n14655), .B(new_n14654), .Y(new_n24893));
  xor_4  g22545(.A(new_n24893), .B(new_n14705), .Y(n9552));
  nand_5 g22546(.A(new_n5106), .B(new_n5107), .Y(new_n24895));
  xor_4  g22547(.A(new_n24895), .B(new_n5113), .Y(n9556));
  xor_4  g22548(.A(new_n12866), .B(new_n10137), .Y(n9558));
  xor_4  g22549(.A(new_n23926), .B(new_n16412), .Y(n9616));
  nand_5 g22550(.A(new_n9789), .B(new_n9790), .Y(new_n24899));
  xnor_4 g22551(.A(new_n24899), .B(new_n9820), .Y(n9622));
  nand_5 g22552(.A(new_n19120), .B(new_n19119), .Y(new_n24901));
  xnor_4 g22553(.A(new_n24901), .B(new_n19135), .Y(n9626));
  nand_5 g22554(.A(new_n5095), .B(new_n5094), .Y(new_n24903));
  xnor_4 g22555(.A(new_n24903), .B(new_n5117), .Y(n9633));
  nand_5 g22556(.A(new_n24808), .B(new_n24800), .Y(new_n24905));
  nand_5 g22557(.A(new_n24905), .B(new_n24801), .Y(new_n24906));
  not_8  g22558(.A(new_n24906), .Y(new_n24907));
  nand_5 g22559(.A(new_n24907), .B(new_n24341), .Y(new_n24908));
  xor_4  g22560(.A(new_n24907), .B(new_n24341), .Y(new_n24909));
  nand_5 g22561(.A(new_n24823), .B(new_n24811), .Y(new_n24910));
  nand_5 g22562(.A(new_n24910), .B(new_n24813), .Y(new_n24911));
  nand_5 g22563(.A(new_n24911), .B(new_n24909), .Y(new_n24912));
  nand_5 g22564(.A(new_n24912), .B(new_n24908), .Y(new_n24913));
  nor_5  g22565(.A(new_n24913), .B(new_n11976), .Y(new_n24914));
  xor_4  g22566(.A(new_n24913), .B(new_n6379_1), .Y(new_n24915));
  or_5   g22567(.A(new_n24911), .B(new_n24909), .Y(new_n24916));
  and_5  g22568(.A(new_n24916), .B(new_n24912), .Y(new_n24917));
  nand_5 g22569(.A(new_n24917), .B(new_n6379_1), .Y(new_n24918));
  not_8  g22570(.A(new_n24917), .Y(new_n24919));
  nand_5 g22571(.A(new_n24919), .B(new_n11976), .Y(new_n24920));
  nand_5 g22572(.A(new_n24826_1), .B(new_n6280), .Y(new_n24921));
  nand_5 g22573(.A(new_n24824), .B(new_n6279), .Y(new_n24922));
  nand_5 g22574(.A(new_n24831), .B(new_n6284), .Y(new_n24923));
  nand_5 g22575(.A(new_n24830), .B(new_n6285), .Y(new_n24924));
  nand_5 g22576(.A(new_n18050), .B(new_n18025_1), .Y(new_n24925));
  nand_5 g22577(.A(new_n24925), .B(new_n18048), .Y(new_n24926));
  nand_5 g22578(.A(new_n24926), .B(new_n24924), .Y(new_n24927));
  nand_5 g22579(.A(new_n24927), .B(new_n24923), .Y(new_n24928));
  nand_5 g22580(.A(new_n24928), .B(new_n24922), .Y(new_n24929));
  nand_5 g22581(.A(new_n24929), .B(new_n24921), .Y(new_n24930));
  nand_5 g22582(.A(new_n24930), .B(new_n24920), .Y(new_n24931));
  nand_5 g22583(.A(new_n24931), .B(new_n24918), .Y(new_n24932));
  nor_5  g22584(.A(new_n24932), .B(new_n24915), .Y(new_n24933));
  nor_5  g22585(.A(new_n24933), .B(new_n24914), .Y(n9635));
  nand_5 g22586(.A(new_n22346), .B(new_n22341_1), .Y(new_n24935));
  xor_4  g22587(.A(new_n24935), .B(new_n22343), .Y(n9648));
  nor_5  g22588(.A(new_n5633), .B(new_n5630), .Y(new_n24937_1));
  nor_5  g22589(.A(new_n24937_1), .B(new_n5635), .Y(n9689));
  nand_5 g22590(.A(new_n12489), .B(new_n12488), .Y(new_n24939));
  xor_4  g22591(.A(new_n24939), .B(new_n12513), .Y(n9695));
  nand_5 g22592(.A(new_n8706), .B(new_n8705), .Y(new_n24941));
  xor_4  g22593(.A(new_n24941), .B(new_n8752), .Y(n9699));
  xor_4  g22594(.A(new_n19244_1), .B(new_n16868), .Y(new_n24943));
  nand_5 g22595(.A(new_n18628), .B(new_n18588), .Y(new_n24944));
  nand_5 g22596(.A(new_n24944), .B(new_n18586), .Y(new_n24945));
  xor_4  g22597(.A(new_n24945), .B(new_n24943), .Y(n9726));
  not_8  g22598(.A(new_n15290), .Y(new_n24947));
  nand_5 g22599(.A(new_n24947), .B(new_n11599), .Y(new_n24948));
  nand_5 g22600(.A(new_n24948), .B(new_n15291), .Y(n9753));
  nand_5 g22601(.A(new_n3644), .B(new_n3645), .Y(new_n24950));
  xnor_4 g22602(.A(new_n24950), .B(new_n3671), .Y(n9761));
  nand_5 g22603(.A(new_n11552), .B(new_n11550), .Y(new_n24952));
  xor_4  g22604(.A(new_n24952), .B(new_n11613), .Y(n9763));
  nand_5 g22605(.A(new_n15651), .B(new_n15650), .Y(new_n24954));
  xnor_4 g22606(.A(new_n24954), .B(new_n15656), .Y(n9767));
  xor_4  g22607(.A(new_n15839), .B(new_n21593), .Y(n9771));
  nor_5  g22608(.A(new_n24446), .B(new_n24445), .Y(new_n24957));
  xor_4  g22609(.A(new_n24957), .B(new_n24448), .Y(n9778));
  nand_5 g22610(.A(new_n18293), .B(new_n18292), .Y(new_n24959));
  xnor_4 g22611(.A(new_n24959), .B(new_n18301_1), .Y(n9783));
  or_5   g22612(.A(new_n7697), .B(new_n7696), .Y(new_n24961));
  xor_4  g22613(.A(new_n24961), .B(new_n7700), .Y(n9803));
  not_8  g22614(.A(new_n20654), .Y(new_n24963));
  nor_5  g22615(.A(new_n23948), .B(n4319), .Y(new_n24964));
  not_8  g22616(.A(new_n24964), .Y(new_n24965));
  nand_5 g22617(.A(new_n24965), .B(new_n24963), .Y(new_n24966));
  nand_5 g22618(.A(new_n24964), .B(new_n20654), .Y(new_n24967));
  nand_5 g22619(.A(new_n24967), .B(new_n24966), .Y(new_n24968));
  nand_5 g22620(.A(new_n23948), .B(n4319), .Y(new_n24969));
  and_5  g22621(.A(new_n24969), .B(new_n24965), .Y(new_n24970));
  nand_5 g22622(.A(new_n24970), .B(new_n20699), .Y(new_n24971));
  or_5   g22623(.A(new_n24970), .B(new_n20699), .Y(new_n24972));
  nand_5 g22624(.A(new_n23950), .B(new_n20705_1), .Y(new_n24973));
  or_5   g22625(.A(new_n23950), .B(new_n20705_1), .Y(new_n24974));
  nand_5 g22626(.A(new_n23895_1), .B(new_n19324), .Y(new_n24975));
  nand_5 g22627(.A(new_n23896), .B(new_n19323_1), .Y(new_n24976));
  nand_5 g22628(.A(new_n23866), .B(new_n19284), .Y(new_n24977));
  or_5   g22629(.A(new_n23866), .B(new_n19284), .Y(new_n24978));
  nand_5 g22630(.A(new_n23869), .B(new_n19288), .Y(new_n24979));
  or_5   g22631(.A(new_n23869), .B(new_n19288), .Y(new_n24980));
  nand_5 g22632(.A(new_n7722), .B(new_n7708_1), .Y(new_n24981));
  nand_5 g22633(.A(new_n24981), .B(new_n7720), .Y(new_n24982));
  nand_5 g22634(.A(new_n24982), .B(new_n24980), .Y(new_n24983));
  nand_5 g22635(.A(new_n24983), .B(new_n24979), .Y(new_n24984));
  nand_5 g22636(.A(new_n24984), .B(new_n24978), .Y(new_n24985));
  nand_5 g22637(.A(new_n24985), .B(new_n24977), .Y(new_n24986));
  nand_5 g22638(.A(new_n24986), .B(new_n24976), .Y(new_n24987));
  nand_5 g22639(.A(new_n24987), .B(new_n24975), .Y(new_n24988));
  nand_5 g22640(.A(new_n24988), .B(new_n24974), .Y(new_n24989));
  nand_5 g22641(.A(new_n24989), .B(new_n24973), .Y(new_n24990));
  nand_5 g22642(.A(new_n24990), .B(new_n24972), .Y(new_n24991));
  nand_5 g22643(.A(new_n24991), .B(new_n24971), .Y(new_n24992));
  not_8  g22644(.A(new_n24992), .Y(new_n24993));
  nand_5 g22645(.A(new_n24965), .B(new_n20696_1), .Y(new_n24994));
  nand_5 g22646(.A(new_n24994), .B(new_n24993), .Y(new_n24995));
  xor_4  g22647(.A(new_n24995), .B(new_n24968), .Y(new_n24996));
  xor_4  g22648(.A(new_n24964), .B(new_n20696_1), .Y(new_n24997));
  xor_4  g22649(.A(new_n24997), .B(new_n24992), .Y(new_n24998_1));
  or_5   g22650(.A(new_n24998_1), .B(new_n3592), .Y(new_n24999));
  nand_5 g22651(.A(new_n24998_1), .B(new_n3592), .Y(new_n25000));
  nand_5 g22652(.A(new_n24971), .B(new_n24972), .Y(new_n25001));
  xor_4  g22653(.A(new_n25001), .B(new_n24990), .Y(new_n25002));
  or_5   g22654(.A(new_n25002), .B(new_n3602), .Y(new_n25003));
  nand_5 g22655(.A(new_n25002), .B(new_n3602), .Y(new_n25004));
  nand_5 g22656(.A(new_n24973), .B(new_n24974), .Y(new_n25005));
  xor_4  g22657(.A(new_n25005), .B(new_n24988), .Y(new_n25006_1));
  or_5   g22658(.A(new_n25006_1), .B(new_n3608), .Y(new_n25007));
  nand_5 g22659(.A(new_n25006_1), .B(new_n3608), .Y(new_n25008));
  nand_5 g22660(.A(new_n24975), .B(new_n24976), .Y(new_n25009));
  xor_4  g22661(.A(new_n25009), .B(new_n24986), .Y(new_n25010));
  or_5   g22662(.A(new_n25010), .B(new_n3615), .Y(new_n25011));
  nand_5 g22663(.A(new_n25010), .B(new_n3615), .Y(new_n25012));
  nand_5 g22664(.A(new_n24977), .B(new_n24978), .Y(new_n25013));
  xor_4  g22665(.A(new_n25013), .B(new_n24984), .Y(new_n25014));
  or_5   g22666(.A(new_n25014), .B(new_n3621), .Y(new_n25015));
  nand_5 g22667(.A(new_n25014), .B(new_n3621), .Y(new_n25016));
  nand_5 g22668(.A(new_n24979), .B(new_n24980), .Y(new_n25017));
  xor_4  g22669(.A(new_n25017), .B(new_n24982), .Y(new_n25018));
  or_5   g22670(.A(new_n25018), .B(new_n3628), .Y(new_n25019));
  nand_5 g22671(.A(new_n25018), .B(new_n3628), .Y(new_n25020));
  nand_5 g22672(.A(new_n7726), .B(new_n7706), .Y(new_n25021));
  nand_5 g22673(.A(new_n25021), .B(new_n7725), .Y(new_n25022));
  nand_5 g22674(.A(new_n25022), .B(new_n25020), .Y(new_n25023_1));
  nand_5 g22675(.A(new_n25023_1), .B(new_n25019), .Y(new_n25024));
  nand_5 g22676(.A(new_n25024), .B(new_n25016), .Y(new_n25025));
  nand_5 g22677(.A(new_n25025), .B(new_n25015), .Y(new_n25026));
  nand_5 g22678(.A(new_n25026), .B(new_n25012), .Y(new_n25027));
  nand_5 g22679(.A(new_n25027), .B(new_n25011), .Y(new_n25028));
  nand_5 g22680(.A(new_n25028), .B(new_n25008), .Y(new_n25029));
  nand_5 g22681(.A(new_n25029), .B(new_n25007), .Y(new_n25030));
  nand_5 g22682(.A(new_n25030), .B(new_n25004), .Y(new_n25031));
  nand_5 g22683(.A(new_n25031), .B(new_n25003), .Y(new_n25032_1));
  nand_5 g22684(.A(new_n25032_1), .B(new_n25000), .Y(new_n25033));
  nand_5 g22685(.A(new_n25033), .B(new_n24999), .Y(new_n25034));
  nand_5 g22686(.A(new_n25034), .B(new_n24996), .Y(new_n25035));
  or_5   g22687(.A(new_n24992), .B(new_n24966), .Y(new_n25036));
  xor_4  g22688(.A(new_n25036), .B(new_n25035), .Y(n9833));
  or_5   g22689(.A(new_n20126_1), .B(n21915), .Y(new_n25038));
  nor_5  g22690(.A(new_n25038), .B(n25972), .Y(new_n25039));
  not_8  g22691(.A(new_n25039), .Y(new_n25040));
  nand_5 g22692(.A(new_n25038), .B(n25972), .Y(new_n25041));
  and_5  g22693(.A(new_n25041), .B(new_n25040), .Y(new_n25042));
  or_5   g22694(.A(new_n25042), .B(new_n20677), .Y(new_n25043));
  nand_5 g22695(.A(new_n20126_1), .B(n21915), .Y(new_n25044));
  nand_5 g22696(.A(new_n25044), .B(new_n25038), .Y(new_n25045));
  or_5   g22697(.A(new_n25045), .B(new_n20683), .Y(new_n25046));
  nand_5 g22698(.A(new_n25045), .B(new_n20683), .Y(new_n25047));
  nand_5 g22699(.A(new_n20130), .B(new_n20123), .Y(new_n25048));
  nand_5 g22700(.A(new_n25048), .B(new_n20129), .Y(new_n25049));
  nand_5 g22701(.A(new_n25049), .B(new_n25047), .Y(new_n25050));
  nand_5 g22702(.A(new_n25050), .B(new_n25046), .Y(new_n25051));
  nand_5 g22703(.A(new_n25051), .B(new_n25043), .Y(new_n25052));
  not_8  g22704(.A(new_n25052), .Y(new_n25053));
  nand_5 g22705(.A(new_n25042), .B(new_n20677), .Y(new_n25054));
  nand_5 g22706(.A(new_n25054), .B(new_n25040), .Y(new_n25055));
  nor_5  g22707(.A(new_n25055), .B(new_n25053), .Y(new_n25056));
  nand_5 g22708(.A(new_n25056), .B(new_n20675), .Y(new_n25057));
  not_8  g22709(.A(new_n25057), .Y(new_n25058));
  nor_5  g22710(.A(new_n25056), .B(new_n20675), .Y(new_n25059));
  or_5   g22711(.A(new_n25059), .B(new_n25058), .Y(new_n25060));
  nor_5  g22712(.A(new_n20116), .B(n3710), .Y(new_n25061));
  nand_5 g22713(.A(new_n25061), .B(new_n11699), .Y(new_n25062_1));
  nor_5  g22714(.A(new_n25062_1), .B(n12507), .Y(new_n25063));
  not_8  g22715(.A(new_n25063), .Y(new_n25064));
  xor_4  g22716(.A(new_n25064), .B(new_n18576_1), .Y(new_n25065));
  not_8  g22717(.A(new_n14898), .Y(new_n25066));
  nand_5 g22718(.A(new_n25062_1), .B(n12507), .Y(new_n25067));
  nand_5 g22719(.A(new_n25067), .B(new_n25064), .Y(new_n25068_1));
  or_5   g22720(.A(new_n25068_1), .B(new_n25066), .Y(new_n25069));
  nand_5 g22721(.A(new_n25068_1), .B(new_n25066), .Y(new_n25070));
  xor_4  g22722(.A(new_n25061), .B(n15077), .Y(new_n25071));
  or_5   g22723(.A(new_n25071), .B(new_n6141), .Y(new_n25072));
  nand_5 g22724(.A(new_n25071), .B(new_n6141), .Y(new_n25073_1));
  nand_5 g22725(.A(new_n20119), .B(new_n20115), .Y(new_n25074_1));
  nand_5 g22726(.A(new_n25074_1), .B(new_n20118), .Y(new_n25075));
  nand_5 g22727(.A(new_n25075), .B(new_n25073_1), .Y(new_n25076));
  nand_5 g22728(.A(new_n25076), .B(new_n25072), .Y(new_n25077));
  nand_5 g22729(.A(new_n25077), .B(new_n25070), .Y(new_n25078));
  nand_5 g22730(.A(new_n25078), .B(new_n25069), .Y(new_n25079));
  xor_4  g22731(.A(new_n25079), .B(new_n25065), .Y(new_n25080));
  not_8  g22732(.A(new_n25080), .Y(new_n25081));
  nand_5 g22733(.A(new_n25081), .B(new_n25060), .Y(new_n25082));
  nand_5 g22734(.A(new_n25054), .B(new_n25043), .Y(new_n25083_1));
  xnor_4 g22735(.A(new_n25083_1), .B(new_n25051), .Y(new_n25084));
  nand_5 g22736(.A(new_n25070), .B(new_n25069), .Y(new_n25085));
  xor_4  g22737(.A(new_n25085), .B(new_n25077), .Y(new_n25086));
  not_8  g22738(.A(new_n25086), .Y(new_n25087));
  or_5   g22739(.A(new_n25087), .B(new_n25084), .Y(new_n25088));
  nand_5 g22740(.A(new_n25087), .B(new_n25084), .Y(new_n25089));
  nand_5 g22741(.A(new_n25073_1), .B(new_n25072), .Y(new_n25090));
  xor_4  g22742(.A(new_n25090), .B(new_n25075), .Y(new_n25091));
  not_8  g22743(.A(new_n25091), .Y(new_n25092));
  nand_5 g22744(.A(new_n25047), .B(new_n25046), .Y(new_n25093));
  xnor_4 g22745(.A(new_n25093), .B(new_n25049), .Y(new_n25094_1));
  or_5   g22746(.A(new_n25094_1), .B(new_n25092), .Y(new_n25095));
  nand_5 g22747(.A(new_n25094_1), .B(new_n25092), .Y(new_n25096));
  nand_5 g22748(.A(new_n20134), .B(new_n20113), .Y(new_n25097_1));
  nand_5 g22749(.A(new_n25097_1), .B(new_n20133), .Y(new_n25098));
  nand_5 g22750(.A(new_n25098), .B(new_n25096), .Y(new_n25099));
  nand_5 g22751(.A(new_n25099), .B(new_n25095), .Y(new_n25100));
  nand_5 g22752(.A(new_n25100), .B(new_n25089), .Y(new_n25101));
  nand_5 g22753(.A(new_n25101), .B(new_n25088), .Y(new_n25102));
  nand_5 g22754(.A(new_n25102), .B(new_n25082), .Y(new_n25103));
  or_5   g22755(.A(new_n25081), .B(new_n25060), .Y(new_n25104));
  nand_5 g22756(.A(new_n25104), .B(new_n25103), .Y(new_n25105));
  nand_5 g22757(.A(new_n25064), .B(new_n18576_1), .Y(new_n25106));
  nor_5  g22758(.A(new_n25079), .B(new_n25106), .Y(new_n25107));
  nor_5  g22759(.A(new_n25107), .B(new_n25058), .Y(new_n25108));
  nor_5  g22760(.A(new_n25108), .B(new_n25105), .Y(new_n25109));
  xor_4  g22761(.A(new_n25109), .B(new_n25058), .Y(n9838));
  nand_5 g22762(.A(new_n22517), .B(new_n22518), .Y(new_n25111));
  xor_4  g22763(.A(new_n25111), .B(new_n22521), .Y(n9867));
  nand_5 g22764(.A(new_n22033), .B(new_n22029), .Y(new_n25113));
  nand_5 g22765(.A(new_n25113), .B(new_n22030), .Y(new_n25114));
  nor_5  g22766(.A(new_n25114), .B(new_n23432), .Y(new_n25115));
  not_8  g22767(.A(new_n25115), .Y(new_n25116));
  nand_5 g22768(.A(new_n25114), .B(new_n23432), .Y(new_n25117));
  and_5  g22769(.A(new_n25117), .B(new_n25116), .Y(new_n25118));
  or_5   g22770(.A(new_n25118), .B(new_n9227), .Y(new_n25119_1));
  nor_5  g22771(.A(new_n22040), .B(new_n22037), .Y(new_n25120_1));
  nor_5  g22772(.A(new_n25120_1), .B(new_n22036), .Y(new_n25121));
  not_8  g22773(.A(new_n25121), .Y(new_n25122));
  nand_5 g22774(.A(new_n25122), .B(new_n25119_1), .Y(new_n25123));
  nand_5 g22775(.A(new_n25118), .B(new_n9227), .Y(new_n25124));
  nand_5 g22776(.A(new_n25124), .B(new_n25123), .Y(new_n25125));
  nor_5  g22777(.A(new_n25125), .B(new_n25115), .Y(new_n25126_1));
  nor_5  g22778(.A(new_n25126_1), .B(new_n9224), .Y(n9890));
  nand_5 g22779(.A(new_n20702), .B(new_n20703), .Y(new_n25128));
  xor_4  g22780(.A(new_n25128), .B(new_n20713_1), .Y(n9917));
  nand_5 g22781(.A(new_n23726), .B(new_n23725), .Y(new_n25130));
  xor_4  g22782(.A(new_n25130), .B(new_n23732), .Y(n9919));
  nand_5 g22783(.A(new_n20904), .B(new_n20905), .Y(new_n25132));
  xor_4  g22784(.A(new_n25132), .B(new_n20919), .Y(n9938));
  nand_5 g22785(.A(new_n20487), .B(new_n20486), .Y(new_n25134));
  xor_4  g22786(.A(new_n25134), .B(new_n20489_1), .Y(n9946));
  nand_5 g22787(.A(n21784), .B(n3740), .Y(new_n25136));
  nand_5 g22788(.A(new_n6796), .B(new_n5496), .Y(new_n25137));
  nand_5 g22789(.A(new_n25137), .B(new_n25136), .Y(new_n25138));
  nand_5 g22790(.A(new_n6800), .B(new_n5502), .Y(new_n25139));
  not_8  g22791(.A(new_n25139), .Y(new_n25140));
  nand_5 g22792(.A(n5521), .B(n2858), .Y(new_n25141));
  not_8  g22793(.A(new_n25141), .Y(new_n25142));
  nand_5 g22794(.A(new_n6804), .B(new_n5508), .Y(new_n25143));
  not_8  g22795(.A(new_n25143), .Y(new_n25144));
  nand_5 g22796(.A(n11926), .B(n2659), .Y(new_n25145));
  not_8  g22797(.A(new_n25145), .Y(new_n25146));
  nand_5 g22798(.A(new_n5514), .B(new_n6807), .Y(new_n25147));
  not_8  g22799(.A(new_n25147), .Y(new_n25148));
  nand_5 g22800(.A(n24327), .B(n4325), .Y(new_n25149));
  not_8  g22801(.A(new_n25149), .Y(new_n25150));
  nand_5 g22802(.A(new_n14879), .B(new_n5526), .Y(new_n25151));
  nand_5 g22803(.A(new_n25151), .B(new_n14878), .Y(new_n25152));
  nand_5 g22804(.A(new_n25152), .B(new_n4137), .Y(new_n25153));
  not_8  g22805(.A(new_n25153), .Y(new_n25154));
  nor_5  g22806(.A(new_n25152), .B(new_n4137), .Y(new_n25155_1));
  nor_5  g22807(.A(new_n25155_1), .B(n22198), .Y(new_n25156));
  nor_5  g22808(.A(new_n25156), .B(new_n25154), .Y(new_n25157));
  nor_5  g22809(.A(new_n25157), .B(new_n25150), .Y(new_n25158));
  nor_5  g22810(.A(new_n25158), .B(new_n25148), .Y(new_n25159));
  nor_5  g22811(.A(new_n25159), .B(new_n25146), .Y(new_n25160));
  nor_5  g22812(.A(new_n25160), .B(new_n25144), .Y(new_n25161));
  nor_5  g22813(.A(new_n25161), .B(new_n25142), .Y(new_n25162));
  nor_5  g22814(.A(new_n25162), .B(new_n25140), .Y(new_n25163));
  xor_4  g22815(.A(new_n25163), .B(new_n25138), .Y(new_n25164));
  or_5   g22816(.A(new_n25164), .B(new_n5424), .Y(new_n25165));
  nand_5 g22817(.A(new_n25164), .B(new_n5424), .Y(new_n25166));
  nand_5 g22818(.A(new_n25166), .B(new_n25165), .Y(new_n25167));
  nand_5 g22819(.A(new_n25141), .B(new_n25139), .Y(new_n25168_1));
  xor_4  g22820(.A(new_n25168_1), .B(new_n25161), .Y(new_n25169));
  or_5   g22821(.A(new_n25169), .B(new_n5427), .Y(new_n25170));
  nand_5 g22822(.A(new_n25169), .B(new_n5427), .Y(new_n25171));
  nand_5 g22823(.A(new_n25145), .B(new_n25143), .Y(new_n25172));
  xor_4  g22824(.A(new_n25172), .B(new_n25159), .Y(new_n25173));
  or_5   g22825(.A(new_n25173), .B(new_n5432), .Y(new_n25174));
  nand_5 g22826(.A(new_n25173), .B(new_n5432), .Y(new_n25175));
  nand_5 g22827(.A(new_n25149), .B(new_n25147), .Y(new_n25176));
  xor_4  g22828(.A(new_n25176), .B(new_n25157), .Y(new_n25177));
  or_5   g22829(.A(new_n25177), .B(new_n5437), .Y(new_n25178));
  nand_5 g22830(.A(new_n25177), .B(new_n5437), .Y(new_n25179));
  nor_5  g22831(.A(new_n25155_1), .B(new_n25154), .Y(new_n25180));
  xor_4  g22832(.A(new_n25180), .B(new_n5520), .Y(new_n25181_1));
  or_5   g22833(.A(new_n25181_1), .B(new_n5442), .Y(new_n25182));
  nand_5 g22834(.A(new_n25181_1), .B(new_n5442), .Y(new_n25183));
  nand_5 g22835(.A(new_n14886), .B(new_n5448), .Y(new_n25184));
  nand_5 g22836(.A(new_n25184), .B(new_n14885), .Y(new_n25185));
  nand_5 g22837(.A(new_n25185), .B(new_n25183), .Y(new_n25186));
  nand_5 g22838(.A(new_n25186), .B(new_n25182), .Y(new_n25187));
  nand_5 g22839(.A(new_n25187), .B(new_n25179), .Y(new_n25188));
  nand_5 g22840(.A(new_n25188), .B(new_n25178), .Y(new_n25189));
  nand_5 g22841(.A(new_n25189), .B(new_n25175), .Y(new_n25190));
  nand_5 g22842(.A(new_n25190), .B(new_n25174), .Y(new_n25191));
  nand_5 g22843(.A(new_n25191), .B(new_n25171), .Y(new_n25192));
  nand_5 g22844(.A(new_n25192), .B(new_n25170), .Y(new_n25193));
  xor_4  g22845(.A(new_n25193), .B(new_n25167), .Y(new_n25194));
  or_5   g22846(.A(new_n25194), .B(new_n19962), .Y(new_n25195));
  nand_5 g22847(.A(new_n25194), .B(new_n19962), .Y(new_n25196));
  nand_5 g22848(.A(new_n25196), .B(new_n25195), .Y(new_n25197));
  nand_5 g22849(.A(new_n25171), .B(new_n25170), .Y(new_n25198));
  xor_4  g22850(.A(new_n25198), .B(new_n25191), .Y(new_n25199));
  or_5   g22851(.A(new_n25199), .B(new_n19218), .Y(new_n25200_1));
  nand_5 g22852(.A(new_n25199), .B(new_n19218), .Y(new_n25201));
  nand_5 g22853(.A(new_n25175), .B(new_n25174), .Y(new_n25202));
  xor_4  g22854(.A(new_n25202), .B(new_n25189), .Y(new_n25203));
  or_5   g22855(.A(new_n25203), .B(new_n19199), .Y(new_n25204));
  nand_5 g22856(.A(new_n25203), .B(new_n19199), .Y(new_n25205));
  nand_5 g22857(.A(new_n25179), .B(new_n25178), .Y(new_n25206));
  xor_4  g22858(.A(new_n25206), .B(new_n25187), .Y(new_n25207));
  or_5   g22859(.A(new_n25207), .B(new_n4306_1), .Y(new_n25208));
  nand_5 g22860(.A(new_n25207), .B(new_n4306_1), .Y(new_n25209_1));
  nand_5 g22861(.A(new_n25183), .B(new_n25182), .Y(new_n25210));
  xor_4  g22862(.A(new_n25210), .B(new_n25185), .Y(new_n25211));
  or_5   g22863(.A(new_n25211), .B(new_n4232), .Y(new_n25212));
  nand_5 g22864(.A(new_n25211), .B(new_n4232), .Y(new_n25213));
  nand_5 g22865(.A(new_n14890), .B(new_n14874), .Y(new_n25214));
  nand_5 g22866(.A(new_n25214), .B(new_n14889), .Y(new_n25215_1));
  nand_5 g22867(.A(new_n25215_1), .B(new_n25213), .Y(new_n25216));
  nand_5 g22868(.A(new_n25216), .B(new_n25212), .Y(new_n25217));
  nand_5 g22869(.A(new_n25217), .B(new_n25209_1), .Y(new_n25218));
  nand_5 g22870(.A(new_n25218), .B(new_n25208), .Y(new_n25219));
  nand_5 g22871(.A(new_n25219), .B(new_n25205), .Y(new_n25220));
  nand_5 g22872(.A(new_n25220), .B(new_n25204), .Y(new_n25221));
  nand_5 g22873(.A(new_n25221), .B(new_n25201), .Y(new_n25222));
  nand_5 g22874(.A(new_n25222), .B(new_n25200_1), .Y(new_n25223));
  xnor_4 g22875(.A(new_n25223), .B(new_n25197), .Y(n9968));
  nor_5  g22876(.A(new_n23367), .B(new_n15904), .Y(new_n25225));
  xor_4  g22877(.A(new_n23367), .B(new_n15903), .Y(new_n25226));
  nand_5 g22878(.A(new_n23375), .B(new_n15903), .Y(new_n25227));
  nand_5 g22879(.A(new_n23374), .B(new_n15904), .Y(new_n25228));
  nand_5 g22880(.A(new_n13121), .B(new_n13070), .Y(new_n25229));
  nand_5 g22881(.A(new_n25229), .B(new_n13071), .Y(new_n25230));
  nand_5 g22882(.A(new_n25230), .B(new_n25228), .Y(new_n25231));
  nand_5 g22883(.A(new_n25231), .B(new_n25227), .Y(new_n25232));
  nor_5  g22884(.A(new_n25232), .B(new_n25226), .Y(new_n25233));
  nor_5  g22885(.A(new_n25233), .B(new_n25225), .Y(n10009));
  nand_5 g22886(.A(new_n24185), .B(new_n24186), .Y(new_n25235));
  xor_4  g22887(.A(new_n25235), .B(new_n24190), .Y(n10010));
  nand_5 g22888(.A(new_n16905_1), .B(new_n16869), .Y(new_n25237));
  nor_5  g22889(.A(new_n25237), .B(new_n16947), .Y(new_n25238));
  xor_4  g22890(.A(new_n25237), .B(new_n16949), .Y(new_n25239));
  nand_5 g22891(.A(new_n16997), .B(new_n16948), .Y(new_n25240_1));
  nand_5 g22892(.A(new_n25240_1), .B(new_n16950), .Y(new_n25241));
  nor_5  g22893(.A(new_n25241), .B(new_n25239), .Y(new_n25242));
  nor_5  g22894(.A(new_n25242), .B(new_n25238), .Y(n10019));
  nor_5  g22895(.A(new_n16693), .B(new_n16692), .Y(new_n25244_1));
  xor_4  g22896(.A(new_n25244_1), .B(new_n16763), .Y(n10021));
  nand_5 g22897(.A(new_n11044_1), .B(new_n11043), .Y(new_n25246));
  xor_4  g22898(.A(new_n25246), .B(new_n11055), .Y(n10055));
  nand_5 g22899(.A(new_n12276), .B(new_n12277), .Y(new_n25248));
  xor_4  g22900(.A(new_n25248), .B(new_n12300), .Y(n10101));
  nand_5 g22901(.A(new_n5071), .B(new_n5069), .Y(new_n25250));
  xnor_4 g22902(.A(new_n25250), .B(new_n5125), .Y(n10111));
  nand_5 g22903(.A(new_n10316), .B(n3324), .Y(new_n25252));
  nand_5 g22904(.A(n16544), .B(new_n18124), .Y(new_n25253));
  nand_5 g22905(.A(n17911), .B(new_n3286), .Y(new_n25254_1));
  nand_5 g22906(.A(new_n18127), .B(n6814), .Y(new_n25255));
  nand_5 g22907(.A(n21997), .B(new_n3186), .Y(new_n25256_1));
  nand_5 g22908(.A(new_n18133), .B(n19701), .Y(new_n25257));
  nand_5 g22909(.A(n25119), .B(new_n3068), .Y(new_n25258));
  nand_5 g22910(.A(new_n9834), .B(n23529), .Y(new_n25259));
  nand_5 g22911(.A(new_n3035), .B(n1163), .Y(new_n25260));
  nand_5 g22912(.A(n24620), .B(new_n9778_1), .Y(new_n25261));
  nand_5 g22913(.A(n18537), .B(new_n3038), .Y(new_n25262));
  nand_5 g22914(.A(new_n9757), .B(n5211), .Y(new_n25263));
  nand_5 g22915(.A(new_n10960), .B(new_n10958), .Y(new_n25264));
  nand_5 g22916(.A(new_n25264), .B(new_n10959), .Y(new_n25265));
  nand_5 g22917(.A(new_n25265), .B(new_n25263), .Y(new_n25266));
  nand_5 g22918(.A(new_n25266), .B(new_n25262), .Y(new_n25267));
  nand_5 g22919(.A(new_n25267), .B(new_n25261), .Y(new_n25268));
  nand_5 g22920(.A(new_n25268), .B(new_n25260), .Y(new_n25269));
  nand_5 g22921(.A(new_n25269), .B(new_n25259), .Y(new_n25270));
  nand_5 g22922(.A(new_n25270), .B(new_n25258), .Y(new_n25271));
  nand_5 g22923(.A(new_n25271), .B(new_n25257), .Y(new_n25272));
  nand_5 g22924(.A(new_n25272), .B(new_n25256_1), .Y(new_n25273));
  nand_5 g22925(.A(new_n25273), .B(new_n25255), .Y(new_n25274));
  nand_5 g22926(.A(new_n25274), .B(new_n25254_1), .Y(new_n25275));
  nand_5 g22927(.A(new_n25275), .B(new_n25253), .Y(new_n25276));
  nand_5 g22928(.A(new_n25276), .B(new_n25252), .Y(new_n25277));
  not_8  g22929(.A(new_n25277), .Y(new_n25278));
  nand_5 g22930(.A(new_n25278), .B(new_n24352), .Y(new_n25279));
  nand_5 g22931(.A(new_n25277), .B(new_n24351), .Y(new_n25280));
  nand_5 g22932(.A(new_n25280), .B(new_n25279), .Y(new_n25281));
  nand_5 g22933(.A(new_n25278), .B(new_n24357), .Y(new_n25282));
  nand_5 g22934(.A(new_n25277), .B(new_n24358), .Y(new_n25283));
  nand_5 g22935(.A(new_n25253), .B(new_n25252), .Y(new_n25284));
  xor_4  g22936(.A(new_n25284), .B(new_n25275), .Y(new_n25285));
  or_5   g22937(.A(new_n25285), .B(new_n19835), .Y(new_n25286));
  nand_5 g22938(.A(new_n25285), .B(new_n19835), .Y(new_n25287));
  nand_5 g22939(.A(new_n25255), .B(new_n25254_1), .Y(new_n25288));
  xor_4  g22940(.A(new_n25288), .B(new_n25273), .Y(new_n25289));
  or_5   g22941(.A(new_n25289), .B(new_n19843), .Y(new_n25290));
  nand_5 g22942(.A(new_n25289), .B(new_n19843), .Y(new_n25291));
  nand_5 g22943(.A(new_n25257), .B(new_n25256_1), .Y(new_n25292));
  xor_4  g22944(.A(new_n25292), .B(new_n25271), .Y(new_n25293_1));
  or_5   g22945(.A(new_n25293_1), .B(new_n19851), .Y(new_n25294));
  nand_5 g22946(.A(new_n25293_1), .B(new_n19851), .Y(new_n25295));
  nand_5 g22947(.A(new_n25259), .B(new_n25258), .Y(new_n25296_1));
  xor_4  g22948(.A(new_n25296_1), .B(new_n25269), .Y(new_n25297));
  or_5   g22949(.A(new_n25297), .B(new_n19859), .Y(new_n25298));
  nand_5 g22950(.A(new_n25297), .B(new_n19859), .Y(new_n25299));
  nand_5 g22951(.A(new_n25261), .B(new_n25260), .Y(new_n25300));
  xor_4  g22952(.A(new_n25300), .B(new_n25267), .Y(new_n25301));
  or_5   g22953(.A(new_n25301), .B(new_n19867), .Y(new_n25302));
  nand_5 g22954(.A(new_n25301), .B(new_n19867), .Y(new_n25303));
  nand_5 g22955(.A(new_n25263), .B(new_n25262), .Y(new_n25304));
  xor_4  g22956(.A(new_n25304), .B(new_n25265), .Y(new_n25305));
  or_5   g22957(.A(new_n25305), .B(new_n19875), .Y(new_n25306));
  nand_5 g22958(.A(new_n25305), .B(new_n19875), .Y(new_n25307));
  nand_5 g22959(.A(new_n10964), .B(new_n10925), .Y(new_n25308));
  nand_5 g22960(.A(new_n25308), .B(new_n10963), .Y(new_n25309));
  nand_5 g22961(.A(new_n25309), .B(new_n25307), .Y(new_n25310));
  nand_5 g22962(.A(new_n25310), .B(new_n25306), .Y(new_n25311));
  nand_5 g22963(.A(new_n25311), .B(new_n25303), .Y(new_n25312));
  nand_5 g22964(.A(new_n25312), .B(new_n25302), .Y(new_n25313));
  nand_5 g22965(.A(new_n25313), .B(new_n25299), .Y(new_n25314));
  nand_5 g22966(.A(new_n25314), .B(new_n25298), .Y(new_n25315));
  nand_5 g22967(.A(new_n25315), .B(new_n25295), .Y(new_n25316_1));
  nand_5 g22968(.A(new_n25316_1), .B(new_n25294), .Y(new_n25317));
  nand_5 g22969(.A(new_n25317), .B(new_n25291), .Y(new_n25318));
  nand_5 g22970(.A(new_n25318), .B(new_n25290), .Y(new_n25319));
  nand_5 g22971(.A(new_n25319), .B(new_n25287), .Y(new_n25320));
  nand_5 g22972(.A(new_n25320), .B(new_n25286), .Y(new_n25321));
  nand_5 g22973(.A(new_n25321), .B(new_n25283), .Y(new_n25322));
  nand_5 g22974(.A(new_n25322), .B(new_n25282), .Y(new_n25323));
  xnor_4 g22975(.A(new_n25323), .B(new_n25281), .Y(n10165));
  nand_5 g22976(.A(new_n14961), .B(new_n14960), .Y(new_n25325));
  xor_4  g22977(.A(new_n25325), .B(new_n14963), .Y(n10236));
  nand_5 g22978(.A(new_n16585), .B(new_n16584_1), .Y(new_n25327));
  xor_4  g22979(.A(new_n25327), .B(new_n16613), .Y(n10239));
  nor_5  g22980(.A(new_n7233_1), .B(new_n7231), .Y(new_n25329));
  xor_4  g22981(.A(new_n25329), .B(new_n7290), .Y(n10244));
  nand_5 g22982(.A(new_n20801), .B(new_n20800), .Y(new_n25331_1));
  xnor_4 g22983(.A(new_n25331_1), .B(new_n20818), .Y(n10261));
  nand_5 g22984(.A(new_n18080), .B(new_n18079), .Y(new_n25333));
  xnor_4 g22985(.A(new_n25333), .B(new_n18096), .Y(n10262));
  nor_5  g22986(.A(new_n19477_1), .B(new_n19476), .Y(new_n25335));
  nor_5  g22987(.A(new_n25335), .B(new_n19479), .Y(n10287));
  not_8  g22988(.A(new_n24624), .Y(new_n25337_1));
  nand_5 g22989(.A(new_n25337_1), .B(new_n24619), .Y(new_n25338));
  nand_5 g22990(.A(new_n24624), .B(new_n24618_1), .Y(new_n25339));
  nand_5 g22991(.A(new_n25339), .B(new_n25338), .Y(new_n25340));
  nand_5 g22992(.A(new_n24641), .B(new_n24628), .Y(new_n25341));
  nand_5 g22993(.A(new_n25341), .B(new_n24630), .Y(new_n25342));
  xor_4  g22994(.A(new_n25342), .B(new_n25340), .Y(n10295));
  nand_5 g22995(.A(new_n17089), .B(new_n17086), .Y(new_n25344));
  xor_4  g22996(.A(new_n25344), .B(new_n17093), .Y(n10321));
  nand_5 g22997(.A(new_n16581), .B(new_n16580), .Y(new_n25346));
  xor_4  g22998(.A(new_n25346), .B(new_n16615), .Y(n10326));
  nand_5 g22999(.A(new_n2964), .B(new_n2963), .Y(new_n25348));
  xnor_4 g23000(.A(new_n25348), .B(new_n2980), .Y(n10327));
  or_5   g23001(.A(new_n23375), .B(new_n23370), .Y(new_n25350));
  nand_5 g23002(.A(new_n25350), .B(new_n23376), .Y(new_n25351));
  xor_4  g23003(.A(new_n25351), .B(new_n23357), .Y(n10330));
  nand_5 g23004(.A(new_n24060), .B(new_n24061), .Y(new_n25353));
  xor_4  g23005(.A(new_n25353), .B(new_n24100), .Y(n10340));
  nand_5 g23006(.A(new_n19482), .B(new_n19486), .Y(new_n25355));
  xor_4  g23007(.A(new_n25355), .B(new_n19485), .Y(n10345));
  not_8  g23008(.A(new_n5492), .Y(new_n25357));
  nand_5 g23009(.A(new_n21980), .B(new_n25357), .Y(new_n25358));
  nand_5 g23010(.A(new_n21979), .B(new_n5492), .Y(new_n25359));
  or_5   g23011(.A(new_n21982), .B(new_n5495), .Y(new_n25360));
  nand_5 g23012(.A(new_n21982), .B(new_n5495), .Y(new_n25361));
  or_5   g23013(.A(new_n21989), .B(new_n5500), .Y(new_n25362_1));
  nand_5 g23014(.A(new_n21989), .B(new_n5500), .Y(new_n25363));
  or_5   g23015(.A(new_n21994), .B(new_n5506), .Y(new_n25364));
  nand_5 g23016(.A(new_n21994), .B(new_n5506), .Y(new_n25365_1));
  or_5   g23017(.A(new_n22000), .B(new_n5512), .Y(new_n25366));
  nand_5 g23018(.A(new_n22000), .B(new_n5512), .Y(new_n25367));
  nand_5 g23019(.A(new_n10846), .B(new_n5516), .Y(new_n25368));
  nand_5 g23020(.A(new_n10845), .B(new_n5518), .Y(new_n25369));
  or_5   g23021(.A(new_n10775_1), .B(new_n5524_1), .Y(new_n25370_1));
  nand_5 g23022(.A(new_n10775_1), .B(new_n5524_1), .Y(new_n25371));
  or_5   g23023(.A(new_n10779), .B(new_n5530), .Y(new_n25372));
  nand_5 g23024(.A(new_n10779), .B(new_n5530), .Y(new_n25373));
  or_5   g23025(.A(new_n10787), .B(new_n5536), .Y(new_n25374));
  nand_5 g23026(.A(new_n10787), .B(new_n5536), .Y(new_n25375));
  or_5   g23027(.A(new_n10793), .B(new_n5542), .Y(new_n25376));
  nand_5 g23028(.A(new_n10793), .B(new_n5542), .Y(new_n25377));
  nand_5 g23029(.A(new_n20559), .B(new_n5550), .Y(new_n25378));
  or_5   g23030(.A(new_n25378), .B(new_n10797), .Y(new_n25379));
  nand_5 g23031(.A(new_n25378), .B(new_n10797), .Y(new_n25380));
  nand_5 g23032(.A(new_n25380), .B(new_n5546), .Y(new_n25381_1));
  nand_5 g23033(.A(new_n25381_1), .B(new_n25379), .Y(new_n25382));
  nand_5 g23034(.A(new_n25382), .B(new_n25377), .Y(new_n25383));
  nand_5 g23035(.A(new_n25383), .B(new_n25376), .Y(new_n25384));
  nand_5 g23036(.A(new_n25384), .B(new_n25375), .Y(new_n25385));
  nand_5 g23037(.A(new_n25385), .B(new_n25374), .Y(new_n25386));
  nand_5 g23038(.A(new_n25386), .B(new_n25373), .Y(new_n25387));
  nand_5 g23039(.A(new_n25387), .B(new_n25372), .Y(new_n25388));
  nand_5 g23040(.A(new_n25388), .B(new_n25371), .Y(new_n25389));
  nand_5 g23041(.A(new_n25389), .B(new_n25370_1), .Y(new_n25390));
  nand_5 g23042(.A(new_n25390), .B(new_n25369), .Y(new_n25391));
  nand_5 g23043(.A(new_n25391), .B(new_n25368), .Y(new_n25392));
  nand_5 g23044(.A(new_n25392), .B(new_n25367), .Y(new_n25393));
  nand_5 g23045(.A(new_n25393), .B(new_n25366), .Y(new_n25394));
  nand_5 g23046(.A(new_n25394), .B(new_n25365_1), .Y(new_n25395));
  nand_5 g23047(.A(new_n25395), .B(new_n25364), .Y(new_n25396));
  nand_5 g23048(.A(new_n25396), .B(new_n25363), .Y(new_n25397));
  nand_5 g23049(.A(new_n25397), .B(new_n25362_1), .Y(new_n25398));
  nand_5 g23050(.A(new_n25398), .B(new_n25361), .Y(new_n25399));
  nand_5 g23051(.A(new_n25399), .B(new_n25360), .Y(new_n25400));
  nand_5 g23052(.A(new_n25400), .B(new_n25359), .Y(new_n25401));
  nand_5 g23053(.A(new_n25401), .B(new_n25358), .Y(n10356));
  nand_5 g23054(.A(new_n22586), .B(new_n22585), .Y(new_n25403));
  xor_4  g23055(.A(new_n25403), .B(new_n22609), .Y(n10385));
  nand_5 g23056(.A(new_n22871_1), .B(new_n22800), .Y(new_n25405));
  nand_5 g23057(.A(new_n25405), .B(new_n22870_1), .Y(new_n25406));
  nor_5  g23058(.A(new_n25406), .B(new_n22796), .Y(n10387));
  nand_5 g23059(.A(new_n23096), .B(new_n23095), .Y(new_n25408));
  xnor_4 g23060(.A(new_n25408), .B(new_n23112), .Y(n10388));
  nand_5 g23061(.A(new_n17772), .B(new_n17771), .Y(new_n25410));
  xor_4  g23062(.A(new_n25410), .B(new_n17834), .Y(n10390));
  xor_4  g23063(.A(new_n10912), .B(new_n10911), .Y(n10404));
  nand_5 g23064(.A(new_n18297), .B(new_n18296), .Y(new_n25413));
  xnor_4 g23065(.A(new_n25413), .B(new_n18299), .Y(n10409));
  xor_4  g23066(.A(new_n18536), .B(new_n18534), .Y(n10420));
  xor_4  g23067(.A(new_n20811), .B(new_n13537), .Y(n10432));
  nand_5 g23068(.A(new_n24182), .B(new_n23507), .Y(new_n25417));
  nand_5 g23069(.A(new_n24292), .B(new_n23508), .Y(new_n25418));
  nand_5 g23070(.A(new_n25418), .B(new_n25417), .Y(new_n25419));
  nand_5 g23071(.A(new_n23818), .B(new_n23816), .Y(new_n25420));
  nand_5 g23072(.A(new_n25420), .B(new_n23817), .Y(new_n25421));
  xor_4  g23073(.A(new_n25421), .B(new_n25419), .Y(new_n25422));
  or_5   g23074(.A(new_n25422), .B(new_n13244), .Y(new_n25423));
  nand_5 g23075(.A(new_n25422), .B(new_n13244), .Y(new_n25424));
  nand_5 g23076(.A(new_n25424), .B(new_n25423), .Y(new_n25425));
  nand_5 g23077(.A(new_n23822), .B(new_n23814), .Y(new_n25426));
  nand_5 g23078(.A(new_n25426), .B(new_n23821), .Y(new_n25427));
  xor_4  g23079(.A(new_n25427), .B(new_n25425), .Y(n10484));
  nand_5 g23080(.A(new_n13096_1), .B(new_n13097), .Y(new_n25429));
  xnor_4 g23081(.A(new_n25429), .B(new_n13110_1), .Y(n10489));
  xor_4  g23082(.A(new_n15455), .B(new_n3829), .Y(n10525));
  nand_5 g23083(.A(new_n20096_1), .B(new_n20095), .Y(new_n25432));
  xor_4  g23084(.A(new_n25432), .B(new_n20103_1), .Y(n10540));
  nand_5 g23085(.A(new_n18387), .B(new_n18385), .Y(new_n25434));
  xnor_4 g23086(.A(new_n25434), .B(new_n18417), .Y(n10561));
  nand_5 g23087(.A(new_n17758), .B(new_n17757), .Y(new_n25436));
  xor_4  g23088(.A(new_n25436), .B(new_n17838), .Y(n10564));
  xor_4  g23089(.A(new_n11599), .B(new_n11597), .Y(n10588));
  nand_5 g23090(.A(new_n11596), .B(new_n11594), .Y(new_n25439));
  xor_4  g23091(.A(new_n25439), .B(new_n11601), .Y(n10595));
  nand_5 g23092(.A(new_n23920), .B(new_n23918), .Y(new_n25441));
  xnor_4 g23093(.A(new_n25441), .B(new_n23935_1), .Y(n10617));
  nand_5 g23094(.A(new_n14247), .B(new_n14248), .Y(new_n25443));
  xor_4  g23095(.A(new_n25443), .B(new_n14325), .Y(n10628));
  or_5   g23096(.A(new_n12240), .B(new_n6473), .Y(new_n25445));
  nand_5 g23097(.A(new_n12240), .B(new_n6473), .Y(new_n25446));
  or_5   g23098(.A(new_n12245), .B(new_n6479), .Y(new_n25447));
  nand_5 g23099(.A(new_n12245), .B(new_n6479), .Y(new_n25448));
  nand_5 g23100(.A(new_n6541), .B(new_n6484), .Y(new_n25449));
  or_5   g23101(.A(new_n25449), .B(new_n6548), .Y(new_n25450));
  nand_5 g23102(.A(new_n25449), .B(new_n6548), .Y(new_n25451));
  nand_5 g23103(.A(new_n25451), .B(new_n6495), .Y(new_n25452));
  nand_5 g23104(.A(new_n25452), .B(new_n25450), .Y(new_n25453));
  nand_5 g23105(.A(new_n25453), .B(new_n25448), .Y(new_n25454));
  nand_5 g23106(.A(new_n25454), .B(new_n25447), .Y(new_n25455));
  nand_5 g23107(.A(new_n25455), .B(new_n25446), .Y(new_n25456));
  nand_5 g23108(.A(new_n25456), .B(new_n25445), .Y(new_n25457));
  or_5   g23109(.A(new_n12235_1), .B(new_n6467), .Y(new_n25458));
  nand_5 g23110(.A(new_n12235_1), .B(new_n6467), .Y(new_n25459));
  nand_5 g23111(.A(new_n25459), .B(new_n25458), .Y(new_n25460_1));
  xnor_4 g23112(.A(new_n25460_1), .B(new_n25457), .Y(n10647));
  nand_5 g23113(.A(new_n3847), .B(new_n3768), .Y(new_n25462));
  nand_5 g23114(.A(new_n25462), .B(new_n3771), .Y(new_n25463));
  and_5  g23115(.A(new_n25463), .B(new_n3708), .Y(new_n25464_1));
  nand_5 g23116(.A(new_n25464_1), .B(new_n15414), .Y(new_n25465));
  nand_5 g23117(.A(new_n25465), .B(new_n9565), .Y(new_n25466));
  nor_5  g23118(.A(new_n25465), .B(new_n9565), .Y(new_n25467));
  not_8  g23119(.A(new_n25467), .Y(new_n25468_1));
  nand_5 g23120(.A(new_n25468_1), .B(new_n25466), .Y(new_n25469));
  not_8  g23121(.A(new_n9567), .Y(new_n25470));
  xor_4  g23122(.A(new_n25464_1), .B(new_n15414), .Y(new_n25471_1));
  or_5   g23123(.A(new_n25471_1), .B(new_n25470), .Y(new_n25472));
  nand_5 g23124(.A(new_n25471_1), .B(new_n25470), .Y(new_n25473));
  nand_5 g23125(.A(new_n4062), .B(new_n3984_1), .Y(new_n25474));
  nand_5 g23126(.A(new_n25474), .B(new_n3983_1), .Y(new_n25475_1));
  nand_5 g23127(.A(new_n25475_1), .B(new_n25473), .Y(new_n25476));
  nand_5 g23128(.A(new_n25476), .B(new_n25472), .Y(new_n25477));
  xnor_4 g23129(.A(new_n25477), .B(new_n25469), .Y(n10653));
  xor_4  g23130(.A(new_n10424), .B(new_n10423), .Y(n10692));
  xor_4  g23131(.A(new_n16799), .B(new_n4754), .Y(n10694));
  nand_5 g23132(.A(new_n22899), .B(new_n22898), .Y(new_n25481));
  xnor_4 g23133(.A(new_n25481), .B(new_n22925), .Y(n10701));
  nand_5 g23134(.A(new_n6954), .B(new_n6953), .Y(new_n25483));
  xnor_4 g23135(.A(new_n25483), .B(new_n6975_1), .Y(n10756));
  nand_5 g23136(.A(new_n18194), .B(new_n18163), .Y(new_n25485));
  nand_5 g23137(.A(new_n25485), .B(new_n18161), .Y(new_n25486));
  not_8  g23138(.A(new_n25486), .Y(new_n25487));
  nand_5 g23139(.A(new_n18196), .B(new_n18160), .Y(new_n25488));
  nand_5 g23140(.A(new_n21941), .B(new_n18201), .Y(new_n25489));
  or_5   g23141(.A(new_n21941), .B(new_n18201), .Y(new_n25490));
  nand_5 g23142(.A(new_n25490), .B(new_n18205), .Y(new_n25491));
  nand_5 g23143(.A(new_n25491), .B(new_n25489), .Y(new_n25492));
  nand_5 g23144(.A(new_n18197), .B(n13419), .Y(new_n25493));
  nand_5 g23145(.A(new_n25493), .B(new_n25492), .Y(new_n25494_1));
  nand_5 g23146(.A(new_n25494_1), .B(new_n25488), .Y(new_n25495));
  nor_5  g23147(.A(new_n25495), .B(new_n25487), .Y(new_n25496));
  xor_4  g23148(.A(new_n25496), .B(new_n3440), .Y(new_n25497));
  xor_4  g23149(.A(new_n25495), .B(new_n25487), .Y(new_n25498));
  nor_5  g23150(.A(new_n25498), .B(new_n3595), .Y(new_n25499_1));
  xor_4  g23151(.A(new_n25492), .B(new_n18200), .Y(new_n25500));
  nand_5 g23152(.A(new_n25500), .B(new_n3458), .Y(new_n25501));
  or_5   g23153(.A(new_n25500), .B(new_n3458), .Y(new_n25502));
  nand_5 g23154(.A(new_n21945), .B(new_n21937), .Y(new_n25503));
  nand_5 g23155(.A(new_n25503), .B(new_n21943_1), .Y(new_n25504));
  nand_5 g23156(.A(new_n25504), .B(new_n25502), .Y(new_n25505));
  nand_5 g23157(.A(new_n25505), .B(new_n25501), .Y(new_n25506));
  nor_5  g23158(.A(new_n25506), .B(new_n25499_1), .Y(new_n25507));
  and_5  g23159(.A(new_n25498), .B(new_n3595), .Y(new_n25508));
  nor_5  g23160(.A(new_n25508), .B(new_n25507), .Y(new_n25509));
  xor_4  g23161(.A(new_n25509), .B(new_n25497), .Y(n10775));
  nand_5 g23162(.A(new_n23840), .B(new_n23841), .Y(new_n25511));
  xnor_4 g23163(.A(new_n25511), .B(new_n23846), .Y(n10780));
  nand_5 g23164(.A(new_n10998), .B(new_n4559), .Y(new_n25513_1));
  nand_5 g23165(.A(n22591), .B(n22274), .Y(new_n25514));
  nand_5 g23166(.A(new_n25514), .B(new_n25513_1), .Y(new_n25515));
  xor_4  g23167(.A(new_n25515), .B(new_n10259), .Y(new_n25516));
  or_5   g23168(.A(new_n10263), .B(new_n10973), .Y(new_n25517));
  nand_5 g23169(.A(new_n10263), .B(new_n10973), .Y(new_n25518_1));
  nand_5 g23170(.A(new_n25518_1), .B(new_n25517), .Y(new_n25519));
  xor_4  g23171(.A(new_n25519), .B(new_n25516), .Y(new_n25520));
  not_8  g23172(.A(new_n25520), .Y(new_n25521));
  or_5   g23173(.A(new_n25521), .B(new_n21016), .Y(new_n25522));
  nand_5 g23174(.A(new_n25521), .B(new_n21016), .Y(new_n25523_1));
  nand_5 g23175(.A(new_n25523_1), .B(new_n10267), .Y(new_n25524));
  nand_5 g23176(.A(new_n25524), .B(new_n25522), .Y(new_n25525));
  nand_5 g23177(.A(new_n25518_1), .B(new_n25516), .Y(new_n25526));
  nand_5 g23178(.A(new_n25526), .B(new_n25517), .Y(new_n25527));
  nand_5 g23179(.A(new_n25514), .B(new_n10258), .Y(new_n25528));
  nand_5 g23180(.A(new_n25528), .B(new_n25513_1), .Y(new_n25529));
  not_8  g23181(.A(new_n25529), .Y(new_n25530));
  nand_5 g23182(.A(new_n10997), .B(new_n4604), .Y(new_n25531));
  nand_5 g23183(.A(n17095), .B(n1689), .Y(new_n25532_1));
  nand_5 g23184(.A(new_n25532_1), .B(new_n25531), .Y(new_n25533));
  xor_4  g23185(.A(new_n25533), .B(new_n25530), .Y(new_n25534));
  not_8  g23186(.A(new_n25534), .Y(new_n25535));
  nand_5 g23187(.A(new_n25535), .B(new_n10969), .Y(new_n25536));
  nand_5 g23188(.A(new_n25534), .B(n21749), .Y(new_n25537));
  nand_5 g23189(.A(new_n25537), .B(new_n25536), .Y(new_n25538));
  xor_4  g23190(.A(new_n25538), .B(new_n25527), .Y(new_n25539_1));
  nand_5 g23191(.A(new_n25539_1), .B(new_n21009), .Y(new_n25540));
  or_5   g23192(.A(new_n25539_1), .B(new_n21009), .Y(new_n25541));
  nand_5 g23193(.A(new_n25541), .B(new_n25540), .Y(new_n25542));
  xnor_4 g23194(.A(new_n25542), .B(new_n25525), .Y(n10817));
  not_8  g23195(.A(new_n24648), .Y(new_n25544));
  nor_5  g23196(.A(new_n24652), .B(new_n25544), .Y(new_n25545));
  nand_5 g23197(.A(new_n24644), .B(new_n23130), .Y(new_n25546));
  nand_5 g23198(.A(new_n24649), .B(new_n25546), .Y(new_n25547));
  nor_5  g23199(.A(new_n25547), .B(new_n25545), .Y(new_n25548));
  nor_5  g23200(.A(new_n25548), .B(new_n8841), .Y(new_n25549));
  xor_4  g23201(.A(new_n25548), .B(new_n8840), .Y(new_n25550_1));
  nand_5 g23202(.A(new_n24660), .B(new_n24655), .Y(new_n25551));
  nand_5 g23203(.A(new_n25551), .B(new_n24656), .Y(new_n25552));
  nor_5  g23204(.A(new_n25552), .B(new_n25550_1), .Y(new_n25553));
  nor_5  g23205(.A(new_n25553), .B(new_n25549), .Y(n10834));
  xor_4  g23206(.A(new_n24932), .B(new_n24915), .Y(n10851));
  nand_5 g23207(.A(new_n24394), .B(new_n24393), .Y(new_n25556));
  xor_4  g23208(.A(new_n25556), .B(new_n24402), .Y(n10874));
  nor_5  g23209(.A(new_n25123), .B(new_n25116), .Y(new_n25558));
  nor_5  g23210(.A(new_n25558), .B(new_n25126_1), .Y(new_n25559));
  xor_4  g23211(.A(new_n25559), .B(new_n9225), .Y(n10924));
  nor_5  g23212(.A(new_n12817), .B(new_n12822), .Y(new_n25561));
  nor_5  g23213(.A(new_n12891), .B(new_n12818), .Y(new_n25562));
  nor_5  g23214(.A(new_n25562), .B(new_n25561), .Y(n10943));
  nand_5 g23215(.A(new_n13683_1), .B(new_n13682), .Y(new_n25564));
  xor_4  g23216(.A(new_n25564), .B(new_n13732), .Y(n10961));
  nand_5 g23217(.A(new_n12173), .B(new_n12171), .Y(new_n25566));
  xor_4  g23218(.A(new_n25566), .B(new_n12185), .Y(n11005));
  nand_5 g23219(.A(new_n24144), .B(new_n24145_1), .Y(new_n25568));
  xor_4  g23220(.A(new_n25568), .B(new_n24153), .Y(n11023));
  nand_5 g23221(.A(new_n20660), .B(new_n8356), .Y(new_n25570));
  nand_5 g23222(.A(new_n20659), .B(new_n8360), .Y(new_n25571));
  or_5   g23223(.A(new_n20664), .B(new_n17115), .Y(new_n25572));
  nand_5 g23224(.A(new_n20664), .B(new_n17115), .Y(new_n25573));
  nand_5 g23225(.A(new_n19308), .B(new_n8370), .Y(new_n25574));
  nand_5 g23226(.A(new_n19307), .B(new_n17041), .Y(new_n25575));
  nand_5 g23227(.A(new_n13988), .B(new_n13982), .Y(new_n25576));
  nand_5 g23228(.A(new_n25576), .B(new_n13987), .Y(new_n25577));
  nand_5 g23229(.A(new_n25577), .B(new_n25575), .Y(new_n25578));
  nand_5 g23230(.A(new_n25578), .B(new_n25574), .Y(new_n25579));
  nand_5 g23231(.A(new_n25579), .B(new_n25573), .Y(new_n25580));
  nand_5 g23232(.A(new_n25580), .B(new_n25572), .Y(new_n25581));
  nand_5 g23233(.A(new_n25581), .B(new_n25571), .Y(new_n25582));
  nand_5 g23234(.A(new_n25582), .B(new_n25570), .Y(new_n25583));
  nand_5 g23235(.A(new_n25583), .B(new_n8333), .Y(new_n25584));
  nor_5  g23236(.A(new_n25584), .B(new_n20657), .Y(new_n25585));
  xor_4  g23237(.A(new_n25583), .B(new_n8333), .Y(new_n25586_1));
  xor_4  g23238(.A(new_n25586_1), .B(new_n20658_1), .Y(new_n25587));
  nand_5 g23239(.A(new_n25587), .B(new_n25081), .Y(new_n25588));
  or_5   g23240(.A(new_n25587), .B(new_n25081), .Y(new_n25589));
  nand_5 g23241(.A(new_n25571), .B(new_n25570), .Y(new_n25590));
  xor_4  g23242(.A(new_n25590), .B(new_n25581), .Y(new_n25591));
  nand_5 g23243(.A(new_n25591), .B(new_n25087), .Y(new_n25592));
  or_5   g23244(.A(new_n25591), .B(new_n25087), .Y(new_n25593));
  nand_5 g23245(.A(new_n25573), .B(new_n25572), .Y(new_n25594));
  xnor_4 g23246(.A(new_n25594), .B(new_n25579), .Y(new_n25595));
  or_5   g23247(.A(new_n25595), .B(new_n25091), .Y(new_n25596));
  nand_5 g23248(.A(new_n25595), .B(new_n25091), .Y(new_n25597));
  not_8  g23249(.A(new_n20121), .Y(new_n25598));
  nand_5 g23250(.A(new_n25575), .B(new_n25574), .Y(new_n25599));
  xor_4  g23251(.A(new_n25599), .B(new_n25577), .Y(new_n25600));
  nand_5 g23252(.A(new_n25600), .B(new_n25598), .Y(new_n25601));
  not_8  g23253(.A(new_n25601), .Y(new_n25602));
  not_8  g23254(.A(new_n25600), .Y(new_n25603));
  nand_5 g23255(.A(new_n25603), .B(new_n20121), .Y(new_n25604));
  not_8  g23256(.A(new_n25604), .Y(new_n25605));
  nand_5 g23257(.A(new_n13992), .B(new_n13972), .Y(new_n25606));
  nand_5 g23258(.A(new_n25606), .B(new_n13991), .Y(new_n25607));
  nor_5  g23259(.A(new_n25607), .B(new_n25605), .Y(new_n25608));
  nor_5  g23260(.A(new_n25608), .B(new_n25602), .Y(new_n25609));
  not_8  g23261(.A(new_n25609), .Y(new_n25610));
  nand_5 g23262(.A(new_n25610), .B(new_n25597), .Y(new_n25611_1));
  nand_5 g23263(.A(new_n25611_1), .B(new_n25596), .Y(new_n25612));
  nand_5 g23264(.A(new_n25612), .B(new_n25593), .Y(new_n25613));
  nand_5 g23265(.A(new_n25613), .B(new_n25592), .Y(new_n25614_1));
  nand_5 g23266(.A(new_n25614_1), .B(new_n25589), .Y(new_n25615));
  nand_5 g23267(.A(new_n25615), .B(new_n25588), .Y(new_n25616));
  xor_4  g23268(.A(new_n25616), .B(new_n25585), .Y(new_n25617));
  not_8  g23269(.A(new_n25617), .Y(new_n25618));
  nor_5  g23270(.A(new_n25585), .B(new_n25107), .Y(new_n25619_1));
  nor_5  g23271(.A(new_n25619_1), .B(new_n25618), .Y(n11025));
  nand_5 g23272(.A(new_n21772), .B(new_n7178), .Y(new_n25621));
  nand_5 g23273(.A(new_n21773), .B(n4590), .Y(new_n25622));
  and_5  g23274(.A(new_n25622), .B(new_n25621), .Y(new_n25623));
  or_5   g23275(.A(new_n25623), .B(new_n10100), .Y(new_n25624));
  nand_5 g23276(.A(new_n25623), .B(new_n10100), .Y(new_n25625));
  nand_5 g23277(.A(new_n21777), .B(new_n21771), .Y(new_n25626));
  nand_5 g23278(.A(new_n25626), .B(new_n21776), .Y(new_n25627));
  nand_5 g23279(.A(new_n25627), .B(new_n25625), .Y(new_n25628));
  nand_5 g23280(.A(new_n25628), .B(new_n25624), .Y(new_n25629_1));
  nor_5  g23281(.A(new_n25621), .B(n25464), .Y(new_n25630));
  not_8  g23282(.A(new_n25630), .Y(new_n25631));
  nand_5 g23283(.A(new_n25621), .B(n25464), .Y(new_n25632));
  and_5  g23284(.A(new_n25632), .B(new_n25631), .Y(new_n25633));
  or_5   g23285(.A(new_n25633), .B(new_n10092), .Y(new_n25634));
  nand_5 g23286(.A(new_n25633), .B(new_n10092), .Y(new_n25635));
  nand_5 g23287(.A(new_n25635), .B(new_n25634), .Y(new_n25636));
  xor_4  g23288(.A(new_n25636), .B(new_n25629_1), .Y(new_n25637));
  not_8  g23289(.A(new_n25637), .Y(new_n25638));
  nand_5 g23290(.A(new_n18845), .B(n1293), .Y(new_n25639));
  nand_5 g23291(.A(new_n18847), .B(new_n7838), .Y(new_n25640));
  nand_5 g23292(.A(new_n21784_1), .B(new_n21782), .Y(new_n25641));
  nand_5 g23293(.A(new_n25641), .B(new_n21783), .Y(new_n25642));
  nand_5 g23294(.A(new_n25642), .B(new_n25640), .Y(new_n25643_1));
  nand_5 g23295(.A(new_n25643_1), .B(new_n25639), .Y(new_n25644));
  nand_5 g23296(.A(new_n18840), .B(n13775), .Y(new_n25645));
  nand_5 g23297(.A(new_n18842), .B(new_n7882), .Y(new_n25646));
  nand_5 g23298(.A(new_n25646), .B(new_n25645), .Y(new_n25647));
  xor_4  g23299(.A(new_n25647), .B(new_n25644), .Y(new_n25648));
  or_5   g23300(.A(new_n25648), .B(new_n25638), .Y(new_n25649));
  nand_5 g23301(.A(new_n25648), .B(new_n25638), .Y(new_n25650));
  nand_5 g23302(.A(new_n25625), .B(new_n25624), .Y(new_n25651));
  xor_4  g23303(.A(new_n25651), .B(new_n25627), .Y(new_n25652));
  not_8  g23304(.A(new_n25652), .Y(new_n25653));
  nand_5 g23305(.A(new_n25640), .B(new_n25639), .Y(new_n25654));
  xor_4  g23306(.A(new_n25654), .B(new_n25642), .Y(new_n25655));
  or_5   g23307(.A(new_n25655), .B(new_n25653), .Y(new_n25656));
  nand_5 g23308(.A(new_n25655), .B(new_n25653), .Y(new_n25657));
  nand_5 g23309(.A(new_n21788), .B(new_n21769), .Y(new_n25658));
  nand_5 g23310(.A(new_n25658), .B(new_n21787), .Y(new_n25659));
  nand_5 g23311(.A(new_n25659), .B(new_n25657), .Y(new_n25660));
  nand_5 g23312(.A(new_n25660), .B(new_n25656), .Y(new_n25661));
  nand_5 g23313(.A(new_n25661), .B(new_n25650), .Y(new_n25662));
  nand_5 g23314(.A(new_n25662), .B(new_n25649), .Y(new_n25663));
  nand_5 g23315(.A(new_n25635), .B(new_n25629_1), .Y(new_n25664));
  nand_5 g23316(.A(new_n25664), .B(new_n25634), .Y(new_n25665_1));
  nand_5 g23317(.A(new_n25630), .B(new_n7170), .Y(new_n25666));
  nand_5 g23318(.A(new_n25631), .B(n3795), .Y(new_n25667));
  and_5  g23319(.A(new_n25667), .B(new_n25666), .Y(new_n25668));
  or_5   g23320(.A(new_n25668), .B(new_n10087), .Y(new_n25669));
  nand_5 g23321(.A(new_n25668), .B(new_n10087), .Y(new_n25670));
  nand_5 g23322(.A(new_n25670), .B(new_n25669), .Y(new_n25671));
  xor_4  g23323(.A(new_n25671), .B(new_n25665_1), .Y(new_n25672));
  not_8  g23324(.A(new_n25672), .Y(new_n25673));
  nand_5 g23325(.A(new_n25646), .B(new_n25644), .Y(new_n25674));
  nand_5 g23326(.A(new_n25674), .B(new_n25645), .Y(new_n25675));
  nand_5 g23327(.A(new_n18835), .B(n21915), .Y(new_n25676));
  nand_5 g23328(.A(new_n18837), .B(new_n7974), .Y(new_n25677));
  nand_5 g23329(.A(new_n25677), .B(new_n25676), .Y(new_n25678));
  xor_4  g23330(.A(new_n25678), .B(new_n25675), .Y(new_n25679));
  or_5   g23331(.A(new_n25679), .B(new_n25673), .Y(new_n25680));
  nand_5 g23332(.A(new_n25679), .B(new_n25673), .Y(new_n25681));
  nand_5 g23333(.A(new_n25681), .B(new_n25680), .Y(new_n25682));
  xnor_4 g23334(.A(new_n25682), .B(new_n25663), .Y(n11063));
  nand_5 g23335(.A(new_n23101), .B(new_n23100), .Y(new_n25684));
  xnor_4 g23336(.A(new_n25684), .B(new_n23110), .Y(n11078));
  nand_5 g23337(.A(new_n23838), .B(new_n23839), .Y(new_n25686));
  xnor_4 g23338(.A(new_n25686), .B(new_n23848), .Y(n11080));
  nand_5 g23339(.A(new_n15783), .B(new_n15782), .Y(new_n25688));
  xor_4  g23340(.A(new_n25688), .B(new_n15800), .Y(n11094));
  nand_5 g23341(.A(new_n25303), .B(new_n25302), .Y(new_n25690));
  xnor_4 g23342(.A(new_n25690), .B(new_n25311), .Y(n11101));
  xor_4  g23343(.A(new_n23931), .B(new_n16419_1), .Y(new_n25692));
  xor_4  g23344(.A(new_n25692), .B(new_n23927), .Y(n11103));
  nand_5 g23345(.A(new_n7431), .B(new_n7433), .Y(new_n25694_1));
  xor_4  g23346(.A(new_n25694_1), .B(new_n7463), .Y(n11120));
  nand_5 g23347(.A(new_n5640), .B(new_n5638), .Y(new_n25696));
  xnor_4 g23348(.A(new_n25696), .B(new_n5642), .Y(n11127));
  nand_5 g23349(.A(new_n17080), .B(new_n17079), .Y(new_n25698));
  xor_4  g23350(.A(new_n25698), .B(new_n17095_1), .Y(n11132));
  nand_5 g23351(.A(new_n12833), .B(new_n12832), .Y(new_n25700));
  xor_4  g23352(.A(new_n25700), .B(new_n12885), .Y(n11134));
  nand_5 g23353(.A(new_n4041), .B(new_n4040), .Y(new_n25702));
  xnor_4 g23354(.A(new_n25702), .B(new_n4046), .Y(n11138));
  nand_5 g23355(.A(new_n12080), .B(new_n12079), .Y(new_n25704));
  xnor_4 g23356(.A(new_n25704), .B(new_n12091), .Y(n11182));
  nor_5  g23357(.A(new_n15759), .B(new_n15758), .Y(new_n25706_1));
  xor_4  g23358(.A(new_n25706_1), .B(new_n15811), .Y(n11234));
  nand_5 g23359(.A(new_n24627), .B(new_n21207), .Y(new_n25708));
  or_5   g23360(.A(new_n24627), .B(new_n21207), .Y(new_n25709));
  nand_5 g23361(.A(new_n25709), .B(new_n25708), .Y(new_n25710));
  nand_5 g23362(.A(new_n24260_1), .B(new_n24236), .Y(new_n25711));
  nand_5 g23363(.A(new_n25711), .B(new_n24238), .Y(new_n25712));
  xor_4  g23364(.A(new_n25712), .B(new_n25710), .Y(n11245));
  nor_5  g23365(.A(new_n9900), .B(new_n9898), .Y(new_n25714));
  xor_4  g23366(.A(new_n25714), .B(new_n9917_1), .Y(n11261));
  nand_5 g23367(.A(new_n25650), .B(new_n25649), .Y(new_n25716));
  xnor_4 g23368(.A(new_n25716), .B(new_n25661), .Y(n11275));
  nand_5 g23369(.A(new_n15478), .B(new_n15410), .Y(n11290));
  nand_5 g23370(.A(new_n10800), .B(new_n10801), .Y(new_n25719_1));
  xnor_4 g23371(.A(new_n25719_1), .B(new_n10807), .Y(n11313));
  nor_5  g23372(.A(new_n19238), .B(new_n19236), .Y(new_n25721));
  xor_4  g23373(.A(new_n25721), .B(new_n19240), .Y(n11325));
  or_5   g23374(.A(new_n15848), .B(new_n15845), .Y(new_n25723));
  xor_4  g23375(.A(new_n25723), .B(new_n15847), .Y(n11326));
  nand_5 g23376(.A(new_n19451), .B(new_n19449), .Y(new_n25725));
  xnor_4 g23377(.A(new_n25725), .B(new_n19494_1), .Y(n11330));
  nand_5 g23378(.A(new_n12848), .B(new_n12847), .Y(new_n25727));
  xor_4  g23379(.A(new_n25727), .B(new_n12879), .Y(n11347));
  nand_5 g23380(.A(new_n25377), .B(new_n25376), .Y(new_n25729));
  xor_4  g23381(.A(new_n25729), .B(new_n25382), .Y(n11348));
  nand_5 g23382(.A(new_n17261), .B(new_n17260), .Y(new_n25731));
  xnor_4 g23383(.A(new_n25731), .B(new_n17269), .Y(n11352));
  nor_5  g23384(.A(new_n20286), .B(new_n20269), .Y(new_n25733));
  nand_5 g23385(.A(new_n20286), .B(new_n20270), .Y(new_n25734));
  not_8  g23386(.A(new_n25734), .Y(new_n25735));
  nor_5  g23387(.A(new_n25735), .B(new_n25733), .Y(new_n25736));
  nand_5 g23388(.A(n22442), .B(new_n18124), .Y(new_n25737));
  nand_5 g23389(.A(new_n8016), .B(n3324), .Y(new_n25738_1));
  nand_5 g23390(.A(new_n18127), .B(n468), .Y(new_n25739));
  nand_5 g23391(.A(n17911), .B(new_n8019), .Y(new_n25740));
  nand_5 g23392(.A(new_n19721), .B(new_n19719), .Y(new_n25741));
  nand_5 g23393(.A(new_n25741), .B(new_n19720), .Y(new_n25742));
  nand_5 g23394(.A(new_n25742), .B(new_n25740), .Y(new_n25743));
  nand_5 g23395(.A(new_n25743), .B(new_n25739), .Y(new_n25744));
  nand_5 g23396(.A(new_n25744), .B(new_n25738_1), .Y(new_n25745));
  nand_5 g23397(.A(new_n25745), .B(new_n25737), .Y(new_n25746));
  nor_5  g23398(.A(new_n25746), .B(new_n25736), .Y(new_n25747));
  and_5  g23399(.A(new_n25746), .B(new_n25736), .Y(new_n25748));
  nor_5  g23400(.A(new_n25748), .B(new_n25747), .Y(new_n25749_1));
  nand_5 g23401(.A(new_n25746), .B(new_n20288), .Y(new_n25750));
  not_8  g23402(.A(new_n25746), .Y(new_n25751_1));
  nand_5 g23403(.A(new_n25751_1), .B(new_n20287_1), .Y(new_n25752));
  not_8  g23404(.A(new_n25752), .Y(new_n25753));
  nand_5 g23405(.A(new_n25738_1), .B(new_n25737), .Y(new_n25754));
  xor_4  g23406(.A(new_n25754), .B(new_n25744), .Y(new_n25755));
  or_5   g23407(.A(new_n25755), .B(new_n20294), .Y(new_n25756_1));
  nand_5 g23408(.A(new_n25755), .B(new_n20294), .Y(new_n25757));
  not_8  g23409(.A(new_n20298), .Y(new_n25758_1));
  nand_5 g23410(.A(new_n25740), .B(new_n25739), .Y(new_n25759));
  xor_4  g23411(.A(new_n25759), .B(new_n25742), .Y(new_n25760));
  or_5   g23412(.A(new_n25760), .B(new_n25758_1), .Y(new_n25761));
  nand_5 g23413(.A(new_n25760), .B(new_n25758_1), .Y(new_n25762));
  not_8  g23414(.A(new_n19703), .Y(new_n25763));
  nor_5  g23415(.A(new_n19726), .B(new_n25763), .Y(new_n25764));
  nor_5  g23416(.A(new_n25764), .B(new_n19725), .Y(new_n25765));
  not_8  g23417(.A(new_n25765), .Y(new_n25766));
  nand_5 g23418(.A(new_n25766), .B(new_n25762), .Y(new_n25767));
  nand_5 g23419(.A(new_n25767), .B(new_n25761), .Y(new_n25768));
  nand_5 g23420(.A(new_n25768), .B(new_n25757), .Y(new_n25769));
  nand_5 g23421(.A(new_n25769), .B(new_n25756_1), .Y(new_n25770));
  nor_5  g23422(.A(new_n25770), .B(new_n25753), .Y(new_n25771));
  not_8  g23423(.A(new_n25771), .Y(new_n25772));
  nand_5 g23424(.A(new_n25772), .B(new_n25750), .Y(new_n25773_1));
  xor_4  g23425(.A(new_n25773_1), .B(new_n25749_1), .Y(n11375));
  nand_5 g23426(.A(new_n14351), .B(new_n14352), .Y(new_n25775));
  xor_4  g23427(.A(new_n25775), .B(new_n8253), .Y(n11379));
  nand_5 g23428(.A(new_n18827), .B(new_n18797), .Y(new_n25777));
  nand_5 g23429(.A(new_n25777), .B(new_n18796), .Y(new_n25778));
  not_8  g23430(.A(new_n25778), .Y(new_n25779));
  nand_5 g23431(.A(new_n25779), .B(new_n13748), .Y(new_n25780));
  or_5   g23432(.A(new_n25779), .B(new_n13748), .Y(new_n25781));
  nand_5 g23433(.A(new_n25781), .B(new_n25780), .Y(new_n25782));
  nand_5 g23434(.A(new_n18877), .B(new_n18830_1), .Y(new_n25783));
  nand_5 g23435(.A(new_n25783), .B(new_n18832), .Y(new_n25784_1));
  xor_4  g23436(.A(new_n25784_1), .B(new_n25782), .Y(new_n25785));
  nand_5 g23437(.A(new_n25785), .B(new_n7206), .Y(new_n25786));
  or_5   g23438(.A(new_n25785), .B(new_n7206), .Y(new_n25787));
  nand_5 g23439(.A(new_n25787), .B(new_n25786), .Y(new_n25788));
  nand_5 g23440(.A(new_n18919_1), .B(new_n18880_1), .Y(new_n25789));
  nand_5 g23441(.A(new_n25789), .B(new_n18879), .Y(new_n25790));
  xnor_4 g23442(.A(new_n25790), .B(new_n25788), .Y(n11386));
  nand_5 g23443(.A(new_n21915_1), .B(new_n21916), .Y(new_n25792_1));
  xnor_4 g23444(.A(new_n25792_1), .B(new_n21926), .Y(n11391));
  nand_5 g23445(.A(new_n24211), .B(new_n24212), .Y(new_n25794));
  xor_4  g23446(.A(new_n25794), .B(new_n24218), .Y(n11398));
  xor_4  g23447(.A(new_n14693), .B(new_n14691), .Y(n11403));
  nand_5 g23448(.A(new_n14067), .B(new_n14068), .Y(new_n25797_1));
  xnor_4 g23449(.A(new_n25797_1), .B(new_n14074), .Y(n11419));
  nand_5 g23450(.A(new_n21710), .B(new_n21709), .Y(new_n25799));
  xnor_4 g23451(.A(new_n25799), .B(new_n21727), .Y(n11439));
  nand_5 g23452(.A(new_n19592), .B(new_n18795), .Y(new_n25801));
  nand_5 g23453(.A(n7569), .B(n2570), .Y(new_n25802));
  nand_5 g23454(.A(new_n25802), .B(new_n25801), .Y(new_n25803));
  nand_5 g23455(.A(new_n18655), .B(new_n13166), .Y(new_n25804));
  nand_5 g23456(.A(n19033), .B(n17037), .Y(new_n25805));
  nand_5 g23457(.A(new_n13191), .B(new_n18801), .Y(new_n25806));
  nand_5 g23458(.A(n5386), .B(n655), .Y(new_n25807));
  nand_5 g23459(.A(new_n13167), .B(new_n17984), .Y(new_n25808));
  nand_5 g23460(.A(n26191), .B(n18145), .Y(new_n25809));
  or_5   g23461(.A(n26512), .B(n10712), .Y(new_n25810));
  nand_5 g23462(.A(n26512), .B(n10712), .Y(new_n25811));
  or_5   g23463(.A(n25126), .B(n19575), .Y(new_n25812));
  nand_5 g23464(.A(n25126), .B(n19575), .Y(new_n25813));
  nand_5 g23465(.A(new_n18811), .B(new_n11028), .Y(new_n25814));
  nand_5 g23466(.A(n19608), .B(n15378), .Y(new_n25815));
  nand_5 g23467(.A(new_n25532_1), .B(new_n25529), .Y(new_n25816_1));
  nand_5 g23468(.A(new_n25816_1), .B(new_n25531), .Y(new_n25817));
  nand_5 g23469(.A(new_n25817), .B(new_n25815), .Y(new_n25818));
  nand_5 g23470(.A(new_n25818), .B(new_n25814), .Y(new_n25819));
  nand_5 g23471(.A(new_n25819), .B(new_n25813), .Y(new_n25820));
  nand_5 g23472(.A(new_n25820), .B(new_n25812), .Y(new_n25821));
  nand_5 g23473(.A(new_n25821), .B(new_n25811), .Y(new_n25822));
  nand_5 g23474(.A(new_n25822), .B(new_n25810), .Y(new_n25823));
  nand_5 g23475(.A(new_n25823), .B(new_n25809), .Y(new_n25824));
  nand_5 g23476(.A(new_n25824), .B(new_n25808), .Y(new_n25825));
  nand_5 g23477(.A(new_n25825), .B(new_n25807), .Y(new_n25826_1));
  nand_5 g23478(.A(new_n25826_1), .B(new_n25806), .Y(new_n25827));
  nand_5 g23479(.A(new_n25827), .B(new_n25805), .Y(new_n25828));
  nand_5 g23480(.A(new_n25828), .B(new_n25804), .Y(new_n25829));
  xor_4  g23481(.A(new_n25829), .B(new_n25803), .Y(new_n25830));
  nand_5 g23482(.A(new_n25830), .B(new_n13220), .Y(new_n25831));
  or_5   g23483(.A(new_n25830), .B(new_n13220), .Y(new_n25832));
  nand_5 g23484(.A(new_n25805), .B(new_n25804), .Y(new_n25833));
  xor_4  g23485(.A(new_n25833), .B(new_n25827), .Y(new_n25834));
  nand_5 g23486(.A(new_n25834), .B(new_n13224), .Y(new_n25835));
  or_5   g23487(.A(new_n25834), .B(new_n13224), .Y(new_n25836));
  nand_5 g23488(.A(new_n25807), .B(new_n25806), .Y(new_n25837));
  xor_4  g23489(.A(new_n25837), .B(new_n25825), .Y(new_n25838));
  nand_5 g23490(.A(new_n25838), .B(new_n13227), .Y(new_n25839_1));
  or_5   g23491(.A(new_n25838), .B(new_n13227), .Y(new_n25840_1));
  nand_5 g23492(.A(new_n25809), .B(new_n25808), .Y(new_n25841));
  xor_4  g23493(.A(new_n25841), .B(new_n25823), .Y(new_n25842));
  nand_5 g23494(.A(new_n25842), .B(new_n12632), .Y(new_n25843));
  or_5   g23495(.A(new_n25842), .B(new_n12632), .Y(new_n25844));
  nand_5 g23496(.A(new_n25811), .B(new_n25810), .Y(new_n25845));
  xor_4  g23497(.A(new_n25845), .B(new_n25821), .Y(new_n25846));
  nand_5 g23498(.A(new_n25846), .B(new_n12539), .Y(new_n25847));
  or_5   g23499(.A(new_n25846), .B(new_n12539), .Y(new_n25848));
  nand_5 g23500(.A(new_n25813), .B(new_n25812), .Y(new_n25849));
  xor_4  g23501(.A(new_n25849), .B(new_n25819), .Y(new_n25850));
  nand_5 g23502(.A(new_n25850), .B(new_n11063_1), .Y(new_n25851));
  nor_5  g23503(.A(new_n25850), .B(new_n11063_1), .Y(new_n25852));
  not_8  g23504(.A(new_n25852), .Y(new_n25853));
  nand_5 g23505(.A(new_n25815), .B(new_n25814), .Y(new_n25854));
  xor_4  g23506(.A(new_n25854), .B(new_n25817), .Y(new_n25855));
  nand_5 g23507(.A(new_n25855), .B(new_n10982), .Y(new_n25856));
  nor_5  g23508(.A(new_n25855), .B(new_n10982), .Y(new_n25857));
  not_8  g23509(.A(new_n25536), .Y(new_n25858));
  not_8  g23510(.A(new_n25537), .Y(new_n25859));
  nor_5  g23511(.A(new_n25859), .B(new_n25527), .Y(new_n25860));
  nor_5  g23512(.A(new_n25860), .B(new_n25858), .Y(new_n25861));
  or_5   g23513(.A(new_n25861), .B(new_n25857), .Y(new_n25862));
  nand_5 g23514(.A(new_n25862), .B(new_n25856), .Y(new_n25863));
  nand_5 g23515(.A(new_n25863), .B(new_n25853), .Y(new_n25864));
  nand_5 g23516(.A(new_n25864), .B(new_n25851), .Y(new_n25865));
  nand_5 g23517(.A(new_n25865), .B(new_n25848), .Y(new_n25866));
  nand_5 g23518(.A(new_n25866), .B(new_n25847), .Y(new_n25867));
  nand_5 g23519(.A(new_n25867), .B(new_n25844), .Y(new_n25868));
  nand_5 g23520(.A(new_n25868), .B(new_n25843), .Y(new_n25869));
  nand_5 g23521(.A(new_n25869), .B(new_n25840_1), .Y(new_n25870));
  nand_5 g23522(.A(new_n25870), .B(new_n25839_1), .Y(new_n25871));
  nand_5 g23523(.A(new_n25871), .B(new_n25836), .Y(new_n25872_1));
  nand_5 g23524(.A(new_n25872_1), .B(new_n25835), .Y(new_n25873_1));
  nand_5 g23525(.A(new_n25873_1), .B(new_n25832), .Y(new_n25874));
  nand_5 g23526(.A(new_n25874), .B(new_n25831), .Y(new_n25875));
  nand_5 g23527(.A(new_n25829), .B(new_n25802), .Y(new_n25876));
  nand_5 g23528(.A(new_n25876), .B(new_n25801), .Y(new_n25877_1));
  xor_4  g23529(.A(new_n25877_1), .B(new_n25875), .Y(new_n25878));
  nor_5  g23530(.A(new_n25666), .B(n6105), .Y(new_n25879));
  xor_4  g23531(.A(new_n25879), .B(new_n12822), .Y(new_n25880));
  xor_4  g23532(.A(new_n25666), .B(n6105), .Y(new_n25881));
  or_5   g23533(.A(new_n25881), .B(new_n10078), .Y(new_n25882));
  nand_5 g23534(.A(new_n25881), .B(new_n10078), .Y(new_n25883));
  nand_5 g23535(.A(new_n25670), .B(new_n25665_1), .Y(new_n25884));
  nand_5 g23536(.A(new_n25884), .B(new_n25669), .Y(new_n25885));
  nand_5 g23537(.A(new_n25885), .B(new_n25883), .Y(new_n25886));
  nand_5 g23538(.A(new_n25886), .B(new_n25882), .Y(new_n25887));
  xor_4  g23539(.A(new_n25887), .B(new_n25880), .Y(new_n25888));
  and_5  g23540(.A(new_n25888), .B(new_n25878), .Y(new_n25889));
  nor_5  g23541(.A(new_n25888), .B(new_n25878), .Y(new_n25890));
  nor_5  g23542(.A(new_n25890), .B(new_n25889), .Y(new_n25891));
  nand_5 g23543(.A(new_n25832), .B(new_n25831), .Y(new_n25892));
  xor_4  g23544(.A(new_n25892), .B(new_n25873_1), .Y(new_n25893));
  nand_5 g23545(.A(new_n25883), .B(new_n25882), .Y(new_n25894));
  xor_4  g23546(.A(new_n25894), .B(new_n25885), .Y(new_n25895));
  not_8  g23547(.A(new_n25895), .Y(new_n25896));
  or_5   g23548(.A(new_n25896), .B(new_n25893), .Y(new_n25897));
  nand_5 g23549(.A(new_n25896), .B(new_n25893), .Y(new_n25898));
  nand_5 g23550(.A(new_n25836), .B(new_n25835), .Y(new_n25899));
  xor_4  g23551(.A(new_n25899), .B(new_n25871), .Y(new_n25900));
  or_5   g23552(.A(new_n25900), .B(new_n25673), .Y(new_n25901));
  nand_5 g23553(.A(new_n25900), .B(new_n25673), .Y(new_n25902));
  nand_5 g23554(.A(new_n25840_1), .B(new_n25839_1), .Y(new_n25903));
  xor_4  g23555(.A(new_n25903), .B(new_n25869), .Y(new_n25904));
  or_5   g23556(.A(new_n25904), .B(new_n25638), .Y(new_n25905));
  nand_5 g23557(.A(new_n25904), .B(new_n25638), .Y(new_n25906));
  nand_5 g23558(.A(new_n25844), .B(new_n25843), .Y(new_n25907));
  xor_4  g23559(.A(new_n25907), .B(new_n25867), .Y(new_n25908));
  or_5   g23560(.A(new_n25908), .B(new_n25653), .Y(new_n25909));
  nand_5 g23561(.A(new_n25908), .B(new_n25653), .Y(new_n25910));
  nand_5 g23562(.A(new_n25848), .B(new_n25847), .Y(new_n25911));
  xor_4  g23563(.A(new_n25911), .B(new_n25865), .Y(new_n25912));
  or_5   g23564(.A(new_n25912), .B(new_n21780), .Y(new_n25913));
  nand_5 g23565(.A(new_n25912), .B(new_n21780), .Y(new_n25914));
  nand_5 g23566(.A(new_n25853), .B(new_n25851), .Y(new_n25915));
  xor_4  g23567(.A(new_n25915), .B(new_n25863), .Y(new_n25916));
  or_5   g23568(.A(new_n25916), .B(new_n21041), .Y(new_n25917));
  nand_5 g23569(.A(new_n25916), .B(new_n21041), .Y(new_n25918));
  not_8  g23570(.A(new_n25857), .Y(new_n25919));
  nand_5 g23571(.A(new_n25919), .B(new_n25856), .Y(new_n25920));
  xor_4  g23572(.A(new_n25920), .B(new_n25861), .Y(new_n25921));
  nand_5 g23573(.A(new_n25921), .B(new_n20991), .Y(new_n25922));
  or_5   g23574(.A(new_n25921), .B(new_n20991), .Y(new_n25923_1));
  nand_5 g23575(.A(new_n25541), .B(new_n25525), .Y(new_n25924));
  nand_5 g23576(.A(new_n25924), .B(new_n25540), .Y(new_n25925));
  nand_5 g23577(.A(new_n25925), .B(new_n25923_1), .Y(new_n25926_1));
  nand_5 g23578(.A(new_n25926_1), .B(new_n25922), .Y(new_n25927));
  nand_5 g23579(.A(new_n25927), .B(new_n25918), .Y(new_n25928));
  nand_5 g23580(.A(new_n25928), .B(new_n25917), .Y(new_n25929));
  nand_5 g23581(.A(new_n25929), .B(new_n25914), .Y(new_n25930));
  nand_5 g23582(.A(new_n25930), .B(new_n25913), .Y(new_n25931));
  nand_5 g23583(.A(new_n25931), .B(new_n25910), .Y(new_n25932));
  nand_5 g23584(.A(new_n25932), .B(new_n25909), .Y(new_n25933));
  nand_5 g23585(.A(new_n25933), .B(new_n25906), .Y(new_n25934_1));
  nand_5 g23586(.A(new_n25934_1), .B(new_n25905), .Y(new_n25935));
  nand_5 g23587(.A(new_n25935), .B(new_n25902), .Y(new_n25936));
  nand_5 g23588(.A(new_n25936), .B(new_n25901), .Y(new_n25937));
  nand_5 g23589(.A(new_n25937), .B(new_n25898), .Y(new_n25938_1));
  nand_5 g23590(.A(new_n25938_1), .B(new_n25897), .Y(new_n25939));
  xor_4  g23591(.A(new_n25939), .B(new_n25891), .Y(n11462));
  nand_5 g23592(.A(new_n23088), .B(new_n23087), .Y(new_n25941));
  xnor_4 g23593(.A(new_n25941), .B(new_n23116), .Y(n11470));
  nand_5 g23594(.A(new_n17610), .B(new_n17612), .Y(new_n25943));
  xor_4  g23595(.A(new_n25943), .B(new_n17628), .Y(n11472));
  nand_5 g23596(.A(new_n21556), .B(new_n21555), .Y(new_n25945));
  xnor_4 g23597(.A(new_n25945), .B(new_n21572), .Y(n11496));
  nand_5 g23598(.A(new_n22818), .B(new_n22816), .Y(new_n25947));
  xnor_4 g23599(.A(new_n25947), .B(new_n22860), .Y(n11506));
  nand_5 g23600(.A(new_n18043_1), .B(new_n6449), .Y(new_n25949));
  or_5   g23601(.A(new_n18043_1), .B(new_n6449), .Y(new_n25950));
  or_5   g23602(.A(new_n12320), .B(new_n6455), .Y(new_n25951));
  nand_5 g23603(.A(new_n12320), .B(new_n6455), .Y(new_n25952));
  or_5   g23604(.A(new_n12269), .B(new_n6461), .Y(new_n25953));
  nand_5 g23605(.A(new_n12269), .B(new_n6461), .Y(new_n25954));
  nand_5 g23606(.A(new_n25459), .B(new_n25457), .Y(new_n25955));
  nand_5 g23607(.A(new_n25955), .B(new_n25458), .Y(new_n25956));
  nand_5 g23608(.A(new_n25956), .B(new_n25954), .Y(new_n25957));
  nand_5 g23609(.A(new_n25957), .B(new_n25953), .Y(new_n25958));
  nand_5 g23610(.A(new_n25958), .B(new_n25952), .Y(new_n25959));
  and_5  g23611(.A(new_n25959), .B(new_n25951), .Y(new_n25960));
  nand_5 g23612(.A(new_n25960), .B(new_n25950), .Y(new_n25961));
  nand_5 g23613(.A(new_n25961), .B(new_n25949), .Y(new_n25962));
  or_5   g23614(.A(new_n24816), .B(new_n6443), .Y(new_n25963));
  nand_5 g23615(.A(new_n24816), .B(new_n6443), .Y(new_n25964));
  nand_5 g23616(.A(new_n25964), .B(new_n25963), .Y(new_n25965));
  xor_4  g23617(.A(new_n25965), .B(new_n25962), .Y(n11515));
  nand_5 g23618(.A(new_n23828), .B(new_n23829), .Y(new_n25967));
  xnor_4 g23619(.A(new_n25967), .B(new_n23858), .Y(n11538));
  nand_5 g23620(.A(new_n21320), .B(new_n21319), .Y(new_n25969));
  xnor_4 g23621(.A(new_n25969), .B(new_n21322), .Y(n11548));
  nand_5 g23622(.A(new_n21591), .B(new_n21592), .Y(new_n25971));
  xor_4  g23623(.A(new_n25971), .B(new_n21599_1), .Y(n11564));
  not_8  g23624(.A(new_n24687), .Y(new_n25973));
  not_8  g23625(.A(new_n24686), .Y(new_n25974_1));
  nor_5  g23626(.A(new_n25974_1), .B(new_n24685), .Y(new_n25975));
  nor_5  g23627(.A(new_n25975), .B(new_n25973), .Y(new_n25976));
  nand_5 g23628(.A(new_n25976), .B(new_n8593), .Y(new_n25977));
  or_5   g23629(.A(new_n25976), .B(new_n8593), .Y(new_n25978));
  nand_5 g23630(.A(new_n24694), .B(new_n24691), .Y(new_n25979));
  nand_5 g23631(.A(new_n25979), .B(new_n24690), .Y(new_n25980));
  nand_5 g23632(.A(new_n25980), .B(new_n25978), .Y(new_n25981));
  nand_5 g23633(.A(new_n25981), .B(new_n25977), .Y(new_n25982));
  nand_5 g23634(.A(new_n24701), .B(new_n24698), .Y(new_n25983));
  nand_5 g23635(.A(new_n25983), .B(new_n24697), .Y(new_n25984));
  not_8  g23636(.A(new_n25984), .Y(new_n25985_1));
  and_5  g23637(.A(new_n25985_1), .B(new_n25982), .Y(new_n25986));
  nor_5  g23638(.A(new_n25985_1), .B(new_n25982), .Y(new_n25987));
  nor_5  g23639(.A(new_n25987), .B(new_n25986), .Y(new_n25988));
  nand_5 g23640(.A(new_n25978), .B(new_n25977), .Y(new_n25989));
  xor_4  g23641(.A(new_n25989), .B(new_n25980), .Y(new_n25990));
  not_8  g23642(.A(new_n25990), .Y(new_n25991));
  nand_5 g23643(.A(new_n25991), .B(new_n25985_1), .Y(new_n25992));
  nand_5 g23644(.A(new_n25990), .B(new_n25984), .Y(new_n25993));
  nor_5  g23645(.A(new_n24709), .B(new_n24705), .Y(new_n25994_1));
  nor_5  g23646(.A(new_n25994_1), .B(new_n24704), .Y(new_n25995));
  not_8  g23647(.A(new_n25995), .Y(new_n25996));
  nand_5 g23648(.A(new_n25996), .B(new_n25993), .Y(new_n25997));
  nand_5 g23649(.A(new_n25997), .B(new_n25992), .Y(new_n25998));
  not_8  g23650(.A(new_n25998), .Y(new_n25999));
  xor_4  g23651(.A(new_n25999), .B(new_n25988), .Y(n11591));
  nand_5 g23652(.A(new_n9554_1), .B(new_n9547), .Y(new_n26001));
  nand_5 g23653(.A(new_n9629), .B(new_n9569), .Y(new_n26002));
  nand_5 g23654(.A(new_n26002), .B(new_n9568), .Y(new_n26003));
  nand_5 g23655(.A(new_n26003), .B(new_n26001), .Y(new_n26004));
  nor_5  g23656(.A(new_n26004), .B(new_n9566), .Y(n11607));
  nand_5 g23657(.A(new_n21238_1), .B(new_n21237), .Y(new_n26006));
  xnor_4 g23658(.A(new_n26006), .B(new_n21267), .Y(n11647));
  nand_5 g23659(.A(new_n25762), .B(new_n25761), .Y(new_n26008));
  xor_4  g23660(.A(new_n26008), .B(new_n25765), .Y(n11674));
  xor_4  g23661(.A(new_n22289), .B(new_n23480_1), .Y(new_n26010));
  nand_5 g23662(.A(new_n24220), .B(new_n24208), .Y(new_n26011));
  nand_5 g23663(.A(new_n26011), .B(new_n24209), .Y(new_n26012));
  xor_4  g23664(.A(new_n26012), .B(new_n26010), .Y(n11682));
  nand_5 g23665(.A(new_n24920), .B(new_n24918), .Y(new_n26014));
  xor_4  g23666(.A(new_n26014), .B(new_n24930), .Y(n11710));
  nand_5 g23667(.A(new_n15773), .B(new_n15772), .Y(new_n26016));
  xor_4  g23668(.A(new_n26016), .B(new_n15804), .Y(n11712));
  nand_5 g23669(.A(new_n24537), .B(new_n24536), .Y(new_n26018));
  xnor_4 g23670(.A(new_n26018), .B(new_n24552), .Y(n11724));
  nand_5 g23671(.A(new_n20611), .B(new_n20612), .Y(new_n26020));
  xor_4  g23672(.A(new_n26020), .B(new_n20614), .Y(n11741));
  xor_4  g23673(.A(new_n20335), .B(new_n3246), .Y(n11770));
  nand_5 g23674(.A(new_n9594), .B(new_n9593), .Y(new_n26023));
  xor_4  g23675(.A(new_n26023), .B(new_n9617), .Y(n11771));
  nor_5  g23676(.A(new_n21411), .B(new_n21410), .Y(new_n26025));
  xor_4  g23677(.A(new_n26025), .B(new_n21447), .Y(n11818));
  nand_5 g23678(.A(new_n25447), .B(new_n25448), .Y(new_n26027));
  xnor_4 g23679(.A(new_n26027), .B(new_n25453), .Y(n11837));
  nand_5 g23680(.A(new_n18555), .B(n2743), .Y(new_n26029));
  nor_5  g23681(.A(new_n18555), .B(n2743), .Y(new_n26030));
  not_8  g23682(.A(new_n26030), .Y(new_n26031));
  and_5  g23683(.A(new_n26031), .B(new_n26029), .Y(new_n26032));
  or_5   g23684(.A(new_n26032), .B(new_n6709), .Y(new_n26033));
  nand_5 g23685(.A(new_n26032), .B(new_n6709), .Y(new_n26034));
  nand_5 g23686(.A(new_n18559), .B(new_n18553), .Y(new_n26035));
  nand_5 g23687(.A(new_n26035), .B(new_n18558_1), .Y(new_n26036_1));
  nand_5 g23688(.A(new_n26036_1), .B(new_n26034), .Y(new_n26037));
  nand_5 g23689(.A(new_n26037), .B(new_n26033), .Y(new_n26038));
  not_8  g23690(.A(new_n26038), .Y(new_n26039));
  nand_5 g23691(.A(new_n26030), .B(new_n15343), .Y(new_n26040));
  nand_5 g23692(.A(new_n26031), .B(new_n15344), .Y(new_n26041));
  nand_5 g23693(.A(new_n26041), .B(new_n26040), .Y(new_n26042));
  xor_4  g23694(.A(new_n26042), .B(new_n26039), .Y(new_n26043));
  nand_5 g23695(.A(new_n26043), .B(new_n24621), .Y(new_n26044));
  or_5   g23696(.A(new_n26043), .B(new_n24621), .Y(new_n26045));
  nand_5 g23697(.A(new_n26045), .B(new_n26044), .Y(new_n26046));
  nand_5 g23698(.A(new_n26034), .B(new_n26033), .Y(new_n26047));
  xnor_4 g23699(.A(new_n26047), .B(new_n26036_1), .Y(new_n26048));
  nand_5 g23700(.A(new_n26048), .B(new_n24123), .Y(new_n26049));
  or_5   g23701(.A(new_n26048), .B(new_n24123), .Y(new_n26050));
  nor_5  g23702(.A(new_n18572_1), .B(new_n18551), .Y(new_n26051));
  nor_5  g23703(.A(new_n26051), .B(new_n18570), .Y(new_n26052));
  not_8  g23704(.A(new_n26052), .Y(new_n26053_1));
  nand_5 g23705(.A(new_n26053_1), .B(new_n26050), .Y(new_n26054_1));
  nand_5 g23706(.A(new_n26054_1), .B(new_n26049), .Y(new_n26055));
  xor_4  g23707(.A(new_n26055), .B(new_n26046), .Y(n11842));
  nand_5 g23708(.A(new_n17952), .B(new_n17951), .Y(new_n26057));
  xnor_4 g23709(.A(new_n26057), .B(new_n17974), .Y(n11843));
  nand_5 g23710(.A(new_n21007), .B(new_n21006), .Y(new_n26059));
  xnor_4 g23711(.A(new_n26059), .B(new_n21028), .Y(n11905));
  nand_5 g23712(.A(new_n13100), .B(new_n13101), .Y(new_n26061));
  xnor_4 g23713(.A(new_n26061), .B(new_n13106), .Y(n11965));
  nand_5 g23714(.A(new_n20912), .B(new_n20913), .Y(new_n26063));
  xor_4  g23715(.A(new_n26063), .B(new_n20915_1), .Y(n12000));
  nand_5 g23716(.A(new_n18636), .B(new_n18637), .Y(new_n26065));
  xor_4  g23717(.A(new_n26065), .B(new_n18639), .Y(n12003));
  nand_5 g23718(.A(new_n19291), .B(new_n19292), .Y(new_n26067));
  xor_4  g23719(.A(new_n26067), .B(new_n19294), .Y(n12011));
  nand_5 g23720(.A(new_n19876), .B(new_n19877), .Y(new_n26069));
  xor_4  g23721(.A(new_n26069), .B(new_n19891), .Y(n12072));
  nand_5 g23722(.A(new_n12281), .B(new_n12282), .Y(new_n26071));
  xor_4  g23723(.A(new_n26071), .B(new_n12298), .Y(n12131));
  nand_5 g23724(.A(new_n18592), .B(new_n18593), .Y(new_n26073));
  xnor_4 g23725(.A(new_n26073), .B(new_n18623), .Y(n12146));
  nand_5 g23726(.A(new_n18905), .B(new_n18904), .Y(new_n26075));
  xnor_4 g23727(.A(new_n26075), .B(new_n18907_1), .Y(n12157));
  nand_5 g23728(.A(new_n11760), .B(new_n11761), .Y(new_n26077));
  xor_4  g23729(.A(new_n26077), .B(new_n11830), .Y(n12158));
  nand_5 g23730(.A(new_n25008), .B(new_n25007), .Y(new_n26079));
  xnor_4 g23731(.A(new_n26079), .B(new_n25028), .Y(n12179));
  nor_5  g23732(.A(new_n7224), .B(new_n7222), .Y(new_n26081));
  xor_4  g23733(.A(new_n26081), .B(new_n7292), .Y(n12192));
  nand_5 g23734(.A(new_n25375), .B(new_n25374), .Y(new_n26083));
  xor_4  g23735(.A(new_n26083), .B(new_n25384), .Y(n12223));
  nand_5 g23736(.A(new_n11767), .B(new_n11768), .Y(new_n26085));
  xor_4  g23737(.A(new_n26085), .B(new_n11828), .Y(n12225));
  nand_5 g23738(.A(new_n25445), .B(new_n25446), .Y(new_n26087));
  xnor_4 g23739(.A(new_n26087), .B(new_n25455), .Y(n12228));
  xor_4  g23740(.A(new_n15265), .B(new_n8282), .Y(n12235));
  nand_5 g23741(.A(new_n10405_1), .B(new_n10404_1), .Y(new_n26090));
  xor_4  g23742(.A(new_n26090), .B(new_n10440), .Y(n12302));
  nand_5 g23743(.A(new_n19024), .B(new_n19025), .Y(new_n26092));
  xor_4  g23744(.A(new_n26092), .B(new_n19057), .Y(n12304));
  nand_5 g23745(.A(n21226), .B(new_n7360), .Y(new_n26094));
  nand_5 g23746(.A(new_n7009), .B(n8244), .Y(new_n26095));
  nand_5 g23747(.A(new_n7329), .B(n4426), .Y(new_n26096_1));
  nand_5 g23748(.A(n9493), .B(new_n7012), .Y(new_n26097));
  nand_5 g23749(.A(new_n22225), .B(new_n22223), .Y(new_n26098));
  nand_5 g23750(.A(new_n26098), .B(new_n22224), .Y(new_n26099));
  nand_5 g23751(.A(new_n26099), .B(new_n26097), .Y(new_n26100));
  nand_5 g23752(.A(new_n26100), .B(new_n26096_1), .Y(new_n26101));
  nand_5 g23753(.A(new_n26101), .B(new_n26095), .Y(new_n26102));
  nand_5 g23754(.A(new_n26102), .B(new_n26094), .Y(new_n26103));
  nand_5 g23755(.A(n23586), .B(new_n7416), .Y(new_n26104));
  nand_5 g23756(.A(new_n7118), .B(n4858), .Y(new_n26105));
  nand_5 g23757(.A(new_n26105), .B(new_n26104), .Y(new_n26106));
  xor_4  g23758(.A(new_n26106), .B(new_n26103), .Y(new_n26107_1));
  or_5   g23759(.A(new_n26107_1), .B(new_n20635), .Y(new_n26108));
  nand_5 g23760(.A(new_n26107_1), .B(new_n20635), .Y(new_n26109));
  nand_5 g23761(.A(new_n26095), .B(new_n26094), .Y(new_n26110));
  xor_4  g23762(.A(new_n26110), .B(new_n26101), .Y(new_n26111_1));
  or_5   g23763(.A(new_n26111_1), .B(new_n20599), .Y(new_n26112));
  nand_5 g23764(.A(new_n26111_1), .B(new_n20599), .Y(new_n26113_1));
  nand_5 g23765(.A(new_n26097), .B(new_n26096_1), .Y(new_n26114));
  xor_4  g23766(.A(new_n26114), .B(new_n26099), .Y(new_n26115));
  or_5   g23767(.A(new_n26115), .B(new_n20603), .Y(new_n26116));
  nand_5 g23768(.A(new_n26115), .B(new_n20603), .Y(new_n26117));
  nand_5 g23769(.A(new_n22229), .B(new_n22221), .Y(new_n26118));
  nand_5 g23770(.A(new_n26118), .B(new_n22228), .Y(new_n26119));
  nand_5 g23771(.A(new_n26119), .B(new_n26117), .Y(new_n26120));
  nand_5 g23772(.A(new_n26120), .B(new_n26116), .Y(new_n26121));
  nand_5 g23773(.A(new_n26121), .B(new_n26113_1), .Y(new_n26122));
  nand_5 g23774(.A(new_n26122), .B(new_n26112), .Y(new_n26123));
  nand_5 g23775(.A(new_n26123), .B(new_n26109), .Y(new_n26124));
  nand_5 g23776(.A(new_n26124), .B(new_n26108), .Y(new_n26125));
  nand_5 g23777(.A(new_n26105), .B(new_n26103), .Y(new_n26126));
  nand_5 g23778(.A(new_n26126), .B(new_n26104), .Y(new_n26127));
  nand_5 g23779(.A(n19196), .B(new_n7491), .Y(new_n26128));
  nand_5 g23780(.A(new_n7003), .B(n1742), .Y(new_n26129));
  nand_5 g23781(.A(new_n26129), .B(new_n26128), .Y(new_n26130));
  xnor_4 g23782(.A(new_n26130), .B(new_n26127), .Y(new_n26131));
  nand_5 g23783(.A(new_n26131), .B(new_n22147), .Y(new_n26132));
  or_5   g23784(.A(new_n26131), .B(new_n22147), .Y(new_n26133));
  nand_5 g23785(.A(new_n26133), .B(new_n26132), .Y(new_n26134));
  xnor_4 g23786(.A(new_n26134), .B(new_n26125), .Y(n12324));
  nand_5 g23787(.A(new_n24213), .B(new_n24214), .Y(new_n26136));
  xor_4  g23788(.A(new_n26136), .B(new_n24216), .Y(n12325));
  nand_5 g23789(.A(new_n12073), .B(new_n12072_1), .Y(new_n26138));
  xnor_4 g23790(.A(new_n26138), .B(new_n12093), .Y(n12329));
  nor_5  g23791(.A(new_n9912), .B(new_n9911), .Y(new_n26140));
  xor_4  g23792(.A(new_n26140), .B(new_n9915), .Y(n12330));
  nand_5 g23793(.A(new_n6451), .B(new_n6450), .Y(new_n26142));
  xnor_4 g23794(.A(new_n26142), .B(new_n6507), .Y(n12346));
  nand_5 g23795(.A(new_n8724), .B(new_n8723), .Y(new_n26144));
  xor_4  g23796(.A(new_n26144), .B(new_n8744_1), .Y(n12349));
  nand_5 g23797(.A(new_n21921), .B(new_n21922), .Y(new_n26146));
  xor_4  g23798(.A(new_n26146), .B(new_n14930), .Y(n12364));
  nor_5  g23799(.A(new_n24907), .B(new_n6522), .Y(new_n26148));
  xor_4  g23800(.A(new_n24906), .B(new_n6522), .Y(new_n26149));
  nand_5 g23801(.A(new_n24906), .B(new_n6380), .Y(new_n26150));
  nand_5 g23802(.A(new_n24907), .B(new_n6381_1), .Y(new_n26151));
  nand_5 g23803(.A(new_n24812), .B(new_n6437_1), .Y(new_n26152));
  or_5   g23804(.A(new_n24812), .B(new_n6437_1), .Y(new_n26153));
  nand_5 g23805(.A(new_n25963), .B(new_n25962), .Y(new_n26154));
  nand_5 g23806(.A(new_n26154), .B(new_n25964), .Y(new_n26155));
  nand_5 g23807(.A(new_n26155), .B(new_n26153), .Y(new_n26156_1));
  nand_5 g23808(.A(new_n26156_1), .B(new_n26152), .Y(new_n26157));
  nand_5 g23809(.A(new_n26157), .B(new_n26151), .Y(new_n26158));
  nand_5 g23810(.A(new_n26158), .B(new_n26150), .Y(new_n26159_1));
  nor_5  g23811(.A(new_n26159_1), .B(new_n26149), .Y(new_n26160));
  nor_5  g23812(.A(new_n26160), .B(new_n26148), .Y(n12383));
  xor_4  g23813(.A(new_n9813), .B(new_n18534), .Y(n12397));
  nand_5 g23814(.A(new_n19471), .B(new_n19470), .Y(new_n26163));
  xor_4  g23815(.A(new_n26163), .B(new_n19488), .Y(n12408));
  nor_5  g23816(.A(new_n22289), .B(new_n17664_1), .Y(new_n26165));
  nor_5  g23817(.A(new_n26012), .B(new_n26010), .Y(new_n26166));
  nor_5  g23818(.A(new_n26166), .B(new_n26165), .Y(n12449));
  nand_5 g23819(.A(new_n23901), .B(new_n23902), .Y(new_n26168));
  xnor_4 g23820(.A(new_n26168), .B(new_n23943), .Y(n12461));
  nand_5 g23821(.A(new_n23769), .B(new_n13748), .Y(new_n26170));
  or_5   g23822(.A(new_n26170), .B(new_n19631), .Y(new_n26171));
  nand_5 g23823(.A(new_n26170), .B(new_n19631), .Y(new_n26172));
  nand_5 g23824(.A(new_n23781), .B(new_n23772), .Y(new_n26173));
  nand_5 g23825(.A(new_n26173), .B(new_n23771), .Y(new_n26174));
  nand_5 g23826(.A(new_n26174), .B(new_n26172), .Y(new_n26175));
  and_5  g23827(.A(new_n26175), .B(new_n26171), .Y(n12462));
  xor_4  g23828(.A(new_n25034), .B(new_n24996), .Y(n12467));
  nand_5 g23829(.A(new_n18250), .B(new_n18199), .Y(new_n26178));
  nand_5 g23830(.A(new_n26178), .B(new_n18198), .Y(new_n26179_1));
  xor_4  g23831(.A(new_n26179_1), .B(new_n25486), .Y(new_n26180_1));
  nand_5 g23832(.A(new_n18158), .B(new_n18123), .Y(new_n26181));
  nand_5 g23833(.A(new_n26181), .B(new_n18125), .Y(new_n26182));
  not_8  g23834(.A(new_n26182), .Y(new_n26183));
  nand_5 g23835(.A(new_n26183), .B(new_n24647), .Y(new_n26184));
  not_8  g23836(.A(new_n26184), .Y(new_n26185));
  nor_5  g23837(.A(new_n26183), .B(new_n24647), .Y(new_n26186));
  nor_5  g23838(.A(new_n26186), .B(new_n26185), .Y(new_n26187));
  nand_5 g23839(.A(new_n26187), .B(new_n26180_1), .Y(new_n26188));
  or_5   g23840(.A(new_n26187), .B(new_n26180_1), .Y(new_n26189));
  nand_5 g23841(.A(new_n18311_1), .B(new_n18253), .Y(new_n26190));
  nand_5 g23842(.A(new_n26190), .B(new_n18252), .Y(new_n26191_1));
  nand_5 g23843(.A(new_n26191_1), .B(new_n26189), .Y(new_n26192));
  nand_5 g23844(.A(new_n26192), .B(new_n26188), .Y(new_n26193));
  nor_5  g23845(.A(new_n26179_1), .B(new_n25486), .Y(new_n26194));
  xor_4  g23846(.A(new_n26194), .B(new_n26184), .Y(new_n26195));
  xor_4  g23847(.A(new_n26195), .B(new_n26193), .Y(n12469));
  nand_5 g23848(.A(new_n12594), .B(new_n12595), .Y(new_n26197));
  xnor_4 g23849(.A(new_n26197), .B(new_n12625), .Y(n12515));
  nand_5 g23850(.A(n10250), .B(new_n14201), .Y(new_n26199));
  nand_5 g23851(.A(new_n7040), .B(n5140), .Y(new_n26200));
  nand_5 g23852(.A(n7674), .B(new_n14204), .Y(new_n26201));
  nand_5 g23853(.A(new_n6991), .B(n6204), .Y(new_n26202));
  nand_5 g23854(.A(n6397), .B(new_n14207), .Y(new_n26203));
  nand_5 g23855(.A(new_n6997), .B(n3349), .Y(new_n26204));
  nand_5 g23856(.A(new_n26129), .B(new_n26127), .Y(new_n26205));
  nand_5 g23857(.A(new_n26205), .B(new_n26128), .Y(new_n26206));
  nand_5 g23858(.A(new_n26206), .B(new_n26204), .Y(new_n26207));
  nand_5 g23859(.A(new_n26207), .B(new_n26203), .Y(new_n26208));
  nand_5 g23860(.A(new_n26208), .B(new_n26202), .Y(new_n26209));
  nand_5 g23861(.A(new_n26209), .B(new_n26201), .Y(new_n26210));
  nand_5 g23862(.A(new_n26210), .B(new_n26200), .Y(new_n26211));
  nand_5 g23863(.A(new_n26211), .B(new_n26199), .Y(new_n26212));
  not_8  g23864(.A(new_n26212), .Y(new_n26213));
  nand_5 g23865(.A(new_n26212), .B(new_n23487), .Y(new_n26214));
  nand_5 g23866(.A(new_n26200), .B(new_n26199), .Y(new_n26215));
  xor_4  g23867(.A(new_n26215), .B(new_n26210), .Y(new_n26216));
  or_5   g23868(.A(new_n26216), .B(new_n23493_1), .Y(new_n26217));
  nand_5 g23869(.A(new_n26216), .B(new_n23493_1), .Y(new_n26218));
  nand_5 g23870(.A(new_n26202), .B(new_n26201), .Y(new_n26219));
  xor_4  g23871(.A(new_n26219), .B(new_n26208), .Y(new_n26220_1));
  or_5   g23872(.A(new_n26220_1), .B(new_n22168), .Y(new_n26221));
  nand_5 g23873(.A(new_n26220_1), .B(new_n22168), .Y(new_n26222));
  nand_5 g23874(.A(new_n26204), .B(new_n26203), .Y(new_n26223));
  xor_4  g23875(.A(new_n26223), .B(new_n26206), .Y(new_n26224_1));
  or_5   g23876(.A(new_n26224_1), .B(new_n22142), .Y(new_n26225));
  nand_5 g23877(.A(new_n26224_1), .B(new_n22142), .Y(new_n26226));
  nand_5 g23878(.A(new_n26133), .B(new_n26125), .Y(new_n26227));
  nand_5 g23879(.A(new_n26227), .B(new_n26132), .Y(new_n26228));
  nand_5 g23880(.A(new_n26228), .B(new_n26226), .Y(new_n26229_1));
  nand_5 g23881(.A(new_n26229_1), .B(new_n26225), .Y(new_n26230));
  nand_5 g23882(.A(new_n26230), .B(new_n26222), .Y(new_n26231));
  nand_5 g23883(.A(new_n26231), .B(new_n26221), .Y(new_n26232));
  nand_5 g23884(.A(new_n26232), .B(new_n26218), .Y(new_n26233));
  nand_5 g23885(.A(new_n26233), .B(new_n26217), .Y(new_n26234));
  nand_5 g23886(.A(new_n26234), .B(new_n26214), .Y(new_n26235));
  nand_5 g23887(.A(new_n26213), .B(new_n23488), .Y(new_n26236));
  nand_5 g23888(.A(new_n26236), .B(new_n26235), .Y(new_n26237_1));
  xor_4  g23889(.A(new_n26237_1), .B(new_n24740), .Y(new_n26238));
  xor_4  g23890(.A(new_n26238), .B(new_n26213), .Y(n12516));
  nand_5 g23891(.A(new_n8532), .B(new_n8531), .Y(new_n26240));
  xor_4  g23892(.A(new_n26240), .B(new_n8546), .Y(n12540));
  nand_5 g23893(.A(new_n13462), .B(new_n13460_1), .Y(new_n26242));
  xor_4  g23894(.A(new_n26242), .B(new_n13473), .Y(n12545));
  nand_5 g23895(.A(new_n23092), .B(new_n23091), .Y(new_n26244));
  xnor_4 g23896(.A(new_n26244), .B(new_n23114), .Y(n12552));
  nand_5 g23897(.A(new_n9386), .B(new_n9385), .Y(new_n26246));
  xnor_4 g23898(.A(new_n26246), .B(new_n9411), .Y(n12566));
  nand_5 g23899(.A(new_n15181), .B(new_n15180_1), .Y(new_n26248));
  xnor_4 g23900(.A(new_n26248), .B(new_n15200), .Y(n12569));
  nand_5 g23901(.A(new_n7207), .B(new_n7208), .Y(new_n26250_1));
  xor_4  g23902(.A(new_n26250_1), .B(new_n7297), .Y(n12607));
  or_5   g23903(.A(new_n11531), .B(new_n11530), .Y(new_n26252));
  xor_4  g23904(.A(new_n26252), .B(new_n11619), .Y(n12620));
  nand_5 g23905(.A(new_n4006), .B(new_n4005), .Y(new_n26254));
  xnor_4 g23906(.A(new_n26254), .B(new_n4056), .Y(n12621));
  nand_5 g23907(.A(new_n20808), .B(new_n20809), .Y(new_n26256));
  xor_4  g23908(.A(new_n26256), .B(new_n20813), .Y(n12654));
  xor_4  g23909(.A(new_n22210), .B(new_n17155), .Y(n12665));
  nand_5 g23910(.A(new_n19515_1), .B(new_n19516), .Y(new_n26259));
  xor_4  g23911(.A(new_n26259), .B(new_n19525), .Y(n12670));
  xor_4  g23912(.A(new_n8733), .B(new_n2544), .Y(n12707));
  nand_5 g23913(.A(new_n8241), .B(new_n8240), .Y(new_n26262));
  xor_4  g23914(.A(new_n26262), .B(new_n8257), .Y(n12725));
  nand_5 g23915(.A(new_n18261), .B(new_n18260), .Y(new_n26264_1));
  xnor_4 g23916(.A(new_n26264_1), .B(new_n18309), .Y(n12727));
  nand_5 g23917(.A(new_n11187), .B(new_n11188), .Y(new_n26266));
  xor_4  g23918(.A(new_n26266), .B(new_n11216), .Y(n12740));
  nand_5 g23919(.A(new_n23454), .B(new_n23451), .Y(new_n26268));
  xor_4  g23920(.A(new_n26268), .B(new_n23453), .Y(n12742));
  xor_4  g23921(.A(new_n23661), .B(new_n23659), .Y(n12746));
  xor_4  g23922(.A(new_n10625), .B(new_n5105), .Y(new_n26271));
  xor_4  g23923(.A(new_n26271), .B(new_n10631), .Y(n12756));
  nand_5 g23924(.A(new_n8205), .B(new_n8204), .Y(new_n26273));
  xor_4  g23925(.A(new_n26273), .B(new_n8269), .Y(n12783));
  nand_5 g23926(.A(new_n26236), .B(new_n26214), .Y(new_n26275));
  xnor_4 g23927(.A(new_n26275), .B(new_n26234), .Y(n12801));
  nand_5 g23928(.A(new_n20232), .B(new_n20231), .Y(new_n26277));
  xor_4  g23929(.A(new_n26277), .B(new_n20234), .Y(n12812));
  nor_5  g23930(.A(new_n18504), .B(new_n18502), .Y(new_n26279));
  xor_4  g23931(.A(new_n26279), .B(new_n18549), .Y(n12816));
  nand_5 g23932(.A(new_n20893), .B(new_n20873), .Y(new_n26281));
  nand_5 g23933(.A(new_n26281), .B(new_n20874), .Y(new_n26282));
  xor_4  g23934(.A(new_n26282), .B(new_n22484_1), .Y(new_n26283));
  nor_5  g23935(.A(new_n26283), .B(new_n26187), .Y(new_n26284));
  nand_5 g23936(.A(new_n20923_1), .B(new_n20895), .Y(new_n26285));
  nand_5 g23937(.A(new_n26285), .B(new_n20896), .Y(new_n26286));
  nor_5  g23938(.A(new_n26286), .B(new_n26284), .Y(new_n26287_1));
  nor_5  g23939(.A(new_n26282), .B(new_n22484_1), .Y(new_n26288));
  not_8  g23940(.A(new_n26288), .Y(new_n26289));
  nand_5 g23941(.A(new_n26283), .B(new_n26187), .Y(new_n26290));
  nand_5 g23942(.A(new_n26290), .B(new_n26289), .Y(new_n26291));
  nor_5  g23943(.A(new_n26291), .B(new_n26287_1), .Y(new_n26292));
  nor_5  g23944(.A(new_n26292), .B(new_n26185), .Y(n12843));
  nand_5 g23945(.A(new_n23711), .B(new_n23712), .Y(new_n26294));
  xor_4  g23946(.A(new_n26294), .B(new_n23714_1), .Y(n12864));
  not_8  g23947(.A(new_n25137), .Y(new_n26296));
  not_8  g23948(.A(new_n25136), .Y(new_n26297));
  nor_5  g23949(.A(new_n25163), .B(new_n26297), .Y(new_n26298));
  nor_5  g23950(.A(new_n26298), .B(new_n26296), .Y(new_n26299));
  or_5   g23951(.A(new_n26299), .B(new_n5493), .Y(new_n26300));
  nand_5 g23952(.A(new_n26299), .B(new_n5493), .Y(new_n26301));
  nand_5 g23953(.A(new_n26301), .B(new_n26300), .Y(new_n26302));
  nand_5 g23954(.A(new_n25193), .B(new_n25166), .Y(new_n26303));
  nand_5 g23955(.A(new_n26303), .B(new_n25165), .Y(new_n26304));
  xor_4  g23956(.A(new_n26304), .B(new_n26302), .Y(new_n26305));
  or_5   g23957(.A(new_n26305), .B(new_n21310), .Y(new_n26306));
  nand_5 g23958(.A(new_n26305), .B(new_n21310), .Y(new_n26307));
  nand_5 g23959(.A(new_n25223), .B(new_n25196), .Y(new_n26308));
  nand_5 g23960(.A(new_n26308), .B(new_n25195), .Y(new_n26309));
  nand_5 g23961(.A(new_n26309), .B(new_n26307), .Y(new_n26310));
  nand_5 g23962(.A(new_n26310), .B(new_n26306), .Y(new_n26311));
  nand_5 g23963(.A(new_n26304), .B(new_n26300), .Y(new_n26312));
  nand_5 g23964(.A(new_n26312), .B(new_n26301), .Y(new_n26313));
  nor_5  g23965(.A(new_n26313), .B(new_n26311), .Y(n12865));
  nand_5 g23966(.A(new_n14767), .B(new_n14766), .Y(new_n26315));
  xor_4  g23967(.A(new_n26315), .B(new_n14788), .Y(n12870));
  nand_5 g23968(.A(new_n23646), .B(new_n23645), .Y(new_n26317_1));
  xor_4  g23969(.A(new_n26317_1), .B(new_n23668), .Y(n12873));
  nand_5 g23970(.A(new_n25337_1), .B(new_n21115), .Y(new_n26319));
  nand_5 g23971(.A(new_n24624), .B(new_n21116), .Y(new_n26320));
  nand_5 g23972(.A(new_n25712), .B(new_n25708), .Y(new_n26321));
  nand_5 g23973(.A(new_n26321), .B(new_n25709), .Y(new_n26322));
  nand_5 g23974(.A(new_n26322), .B(new_n26320), .Y(new_n26323));
  nand_5 g23975(.A(new_n26323), .B(new_n26319), .Y(n12904));
  nand_5 g23976(.A(new_n12058), .B(new_n12057), .Y(new_n26325));
  xnor_4 g23977(.A(new_n26325), .B(new_n12097), .Y(n12941));
  nand_5 g23978(.A(new_n12929), .B(new_n12928), .Y(new_n26327));
  xnor_4 g23979(.A(new_n26327), .B(new_n12939), .Y(n12942));
  xor_4  g23980(.A(new_n6622), .B(new_n4204_1), .Y(new_n26329));
  xor_4  g23981(.A(new_n26329), .B(new_n6627), .Y(n12978));
  xor_4  g23982(.A(new_n11255), .B(new_n9071), .Y(n12980));
  xor_4  g23983(.A(new_n7449), .B(new_n5193), .Y(n12985));
  nand_5 g23984(.A(new_n16577), .B(new_n16576), .Y(new_n26333));
  xor_4  g23985(.A(new_n26333), .B(new_n16617_1), .Y(n12987));
  nand_5 g23986(.A(new_n19165), .B(new_n19149), .Y(new_n26335));
  nand_5 g23987(.A(new_n26335), .B(new_n19150), .Y(new_n26336));
  nor_5  g23988(.A(new_n26336), .B(new_n16906), .Y(new_n26337));
  not_8  g23989(.A(new_n26336), .Y(new_n26338));
  nor_5  g23990(.A(new_n26338), .B(new_n16907), .Y(new_n26339));
  or_5   g23991(.A(new_n26339), .B(new_n26337), .Y(new_n26340));
  nand_5 g23992(.A(new_n19189), .B(new_n19167), .Y(new_n26341));
  nand_5 g23993(.A(new_n26341), .B(new_n19168), .Y(new_n26342));
  xor_4  g23994(.A(new_n26342), .B(new_n26340), .Y(n12992));
  not_8  g23995(.A(new_n24970), .Y(new_n26344));
  nand_5 g23996(.A(new_n26344), .B(new_n18162), .Y(new_n26345));
  not_8  g23997(.A(new_n26345), .Y(new_n26346));
  nand_5 g23998(.A(new_n23952), .B(new_n23947), .Y(new_n26347));
  nand_5 g23999(.A(new_n26347), .B(new_n23951), .Y(new_n26348));
  nor_5  g24000(.A(new_n26348), .B(new_n26346), .Y(new_n26349));
  nand_5 g24001(.A(new_n24970), .B(n6659), .Y(new_n26350));
  nand_5 g24002(.A(new_n26350), .B(new_n24965), .Y(new_n26351));
  nor_5  g24003(.A(new_n26351), .B(new_n26349), .Y(new_n26352));
  nand_5 g24004(.A(new_n26352), .B(new_n22498), .Y(new_n26353_1));
  not_8  g24005(.A(new_n26352), .Y(new_n26354));
  nand_5 g24006(.A(new_n26354), .B(new_n22508), .Y(new_n26355));
  nand_5 g24007(.A(new_n26355), .B(new_n26353_1), .Y(new_n26356));
  nand_5 g24008(.A(new_n26350), .B(new_n26345), .Y(new_n26357));
  xor_4  g24009(.A(new_n26357), .B(new_n26348), .Y(new_n26358));
  or_5   g24010(.A(new_n26358), .B(new_n22516), .Y(new_n26359));
  not_8  g24011(.A(new_n26359), .Y(new_n26360));
  nand_5 g24012(.A(new_n26358), .B(new_n22516), .Y(new_n26361));
  not_8  g24013(.A(new_n26361), .Y(new_n26362));
  nor_5  g24014(.A(new_n23957), .B(new_n23945), .Y(new_n26363));
  nor_5  g24015(.A(new_n26363), .B(new_n23956), .Y(new_n26364));
  nor_5  g24016(.A(new_n26364), .B(new_n26362), .Y(new_n26365));
  nor_5  g24017(.A(new_n26365), .B(new_n26360), .Y(new_n26366));
  xnor_4 g24018(.A(new_n26366), .B(new_n26356), .Y(n13005));
  nor_5  g24019(.A(new_n22596), .B(new_n18993), .Y(new_n26368));
  nor_5  g24020(.A(new_n26368), .B(new_n22598), .Y(n13043));
  nand_5 g24021(.A(new_n20295), .B(new_n20296), .Y(new_n26370));
  xor_4  g24022(.A(new_n26370), .B(new_n20316), .Y(n13048));
  nand_5 g24023(.A(new_n17584), .B(new_n17583_1), .Y(new_n26372));
  xor_4  g24024(.A(new_n26372), .B(new_n17586), .Y(n13054));
  nand_5 g24025(.A(new_n20477), .B(new_n20476), .Y(new_n26374));
  xnor_4 g24026(.A(new_n26374), .B(new_n20492), .Y(n13082));
  nand_5 g24027(.A(new_n8229), .B(new_n8228), .Y(new_n26376));
  xor_4  g24028(.A(new_n26376), .B(new_n8261), .Y(n13096));
  nand_5 g24029(.A(new_n20471), .B(new_n20470_1), .Y(new_n26378));
  xnor_4 g24030(.A(new_n26378), .B(new_n20494), .Y(n13116));
  nand_5 g24031(.A(new_n22574), .B(new_n22573), .Y(new_n26380));
  xor_4  g24032(.A(new_n26380), .B(new_n22615), .Y(n13122));
  nand_5 g24033(.A(new_n7274), .B(new_n7272), .Y(new_n26382));
  xnor_4 g24034(.A(new_n26382), .B(new_n7278), .Y(n13141));
  nand_5 g24035(.A(new_n22430), .B(new_n22429), .Y(new_n26384));
  xor_4  g24036(.A(new_n26384), .B(new_n22442_1), .Y(n13144));
  nand_5 g24037(.A(new_n23079), .B(new_n23078), .Y(new_n26386));
  xnor_4 g24038(.A(new_n26386), .B(new_n23120_1), .Y(n13168));
  nand_5 g24039(.A(new_n23834), .B(new_n23835), .Y(new_n26388));
  xnor_4 g24040(.A(new_n26388), .B(new_n23852), .Y(n13198));
  nand_5 g24041(.A(new_n16589_1), .B(new_n16588), .Y(new_n26390));
  xnor_4 g24042(.A(new_n26390), .B(new_n16610), .Y(n13199));
  nor_5  g24043(.A(new_n16728), .B(new_n16727), .Y(new_n26392));
  xor_4  g24044(.A(new_n26392), .B(new_n16747), .Y(n13204));
  nand_5 g24045(.A(new_n11788), .B(new_n11789), .Y(new_n26394));
  xor_4  g24046(.A(new_n26394), .B(new_n11822), .Y(n13209));
  nand_5 g24047(.A(new_n22189), .B(new_n22188), .Y(new_n26396_1));
  xor_4  g24048(.A(new_n26396_1), .B(new_n22197), .Y(n13270));
  nand_5 g24049(.A(new_n15074), .B(new_n15073), .Y(new_n26398));
  xor_4  g24050(.A(new_n26398), .B(new_n15098), .Y(n13273));
  nand_5 g24051(.A(new_n25004), .B(new_n25003), .Y(new_n26400));
  xnor_4 g24052(.A(new_n26400), .B(new_n25030), .Y(n13285));
  or_5   g24053(.A(new_n24302), .B(new_n24301), .Y(new_n26402));
  xor_4  g24054(.A(new_n26402), .B(new_n24325), .Y(n13338));
  nand_5 g24055(.A(new_n9057), .B(new_n9056), .Y(new_n26404));
  xor_4  g24056(.A(new_n26404), .B(new_n9090_1), .Y(n13407));
  nand_5 g24057(.A(new_n18606), .B(new_n18607), .Y(new_n26406));
  xnor_4 g24058(.A(new_n26406), .B(new_n18609), .Y(n13409));
  nand_5 g24059(.A(new_n6084_1), .B(new_n6085), .Y(new_n26408_1));
  xor_4  g24060(.A(new_n26408_1), .B(new_n6126), .Y(n13456));
  nor_5  g24061(.A(new_n24163), .B(new_n23504), .Y(new_n26410));
  and_5  g24062(.A(new_n24166), .B(new_n23505), .Y(new_n26411));
  nand_5 g24063(.A(new_n25421), .B(new_n25418), .Y(new_n26412));
  nand_5 g24064(.A(new_n26412), .B(new_n25417), .Y(new_n26413));
  nor_5  g24065(.A(new_n26413), .B(new_n26411), .Y(new_n26414));
  nand_5 g24066(.A(new_n26414), .B(new_n26410), .Y(new_n26415));
  xor_4  g24067(.A(new_n24163), .B(new_n23505), .Y(new_n26416));
  xor_4  g24068(.A(new_n26416), .B(new_n26414), .Y(new_n26417));
  xor_4  g24069(.A(new_n24166), .B(new_n23504), .Y(new_n26418));
  xor_4  g24070(.A(new_n26418), .B(new_n26413), .Y(new_n26419));
  nand_5 g24071(.A(new_n26419), .B(new_n13239), .Y(new_n26420));
  or_5   g24072(.A(new_n26419), .B(new_n13239), .Y(new_n26421));
  nand_5 g24073(.A(new_n25427), .B(new_n25423), .Y(new_n26422));
  nand_5 g24074(.A(new_n26422), .B(new_n25424), .Y(new_n26423));
  nand_5 g24075(.A(new_n26423), .B(new_n26421), .Y(new_n26424));
  nand_5 g24076(.A(new_n26424), .B(new_n26420), .Y(new_n26425));
  nand_5 g24077(.A(new_n26425), .B(new_n26417), .Y(new_n26426));
  nand_5 g24078(.A(new_n26426), .B(new_n26415), .Y(n13457));
  nand_5 g24079(.A(new_n14005), .B(new_n14004_1), .Y(new_n26428));
  xor_4  g24080(.A(new_n26428), .B(new_n14014), .Y(n13477));
  nand_5 g24081(.A(new_n14341), .B(new_n14340), .Y(new_n26430));
  xor_4  g24082(.A(new_n26430), .B(new_n14362), .Y(n13484));
  nand_5 g24083(.A(new_n23298), .B(new_n23299), .Y(new_n26432));
  xor_4  g24084(.A(new_n26432), .B(new_n23333_1), .Y(n13486));
  nand_5 g24085(.A(new_n24917), .B(new_n24355), .Y(new_n26434));
  nand_5 g24086(.A(new_n24919), .B(new_n24337), .Y(new_n26435));
  nand_5 g24087(.A(new_n26435), .B(new_n26434), .Y(new_n26436));
  nand_5 g24088(.A(new_n24853_1), .B(new_n24825), .Y(new_n26437));
  nand_5 g24089(.A(new_n26437), .B(new_n24827), .Y(new_n26438));
  xor_4  g24090(.A(new_n26438), .B(new_n26436), .Y(n13487));
  nand_5 g24091(.A(new_n5832), .B(new_n5831), .Y(new_n26440));
  xnor_4 g24092(.A(new_n26440), .B(new_n5854), .Y(n13500));
  nand_5 g24093(.A(new_n5101_1), .B(new_n5100), .Y(new_n26442));
  xnor_4 g24094(.A(new_n26442), .B(new_n5115_1), .Y(n13501));
  nand_5 g24095(.A(new_n7256_1), .B(new_n7254), .Y(new_n26444));
  xnor_4 g24096(.A(new_n26444), .B(new_n7284), .Y(n13506));
  nand_5 g24097(.A(new_n6960), .B(new_n6959), .Y(new_n26446));
  xor_4  g24098(.A(new_n26446), .B(new_n6973), .Y(n13548));
  nand_5 g24099(.A(new_n25910), .B(new_n25909), .Y(new_n26448));
  xnor_4 g24100(.A(new_n26448), .B(new_n25931), .Y(n13551));
  nand_5 g24101(.A(new_n5623), .B(new_n5622), .Y(new_n26450));
  xor_4  g24102(.A(new_n26450), .B(new_n5647), .Y(n13602));
  nand_5 g24103(.A(new_n19924), .B(new_n19923_1), .Y(new_n26452_1));
  xor_4  g24104(.A(new_n26452_1), .B(new_n19933), .Y(n13626));
  nand_5 g24105(.A(new_n9398), .B(new_n9397), .Y(new_n26454));
  xnor_4 g24106(.A(new_n26454), .B(new_n9407), .Y(n13683));
  nand_5 g24107(.A(new_n22813), .B(new_n22811), .Y(new_n26456));
  xnor_4 g24108(.A(new_n26456), .B(new_n22862), .Y(n13710));
  nand_5 g24109(.A(new_n22421), .B(new_n22422), .Y(new_n26458));
  xnor_4 g24110(.A(new_n26458), .B(new_n22446), .Y(n13722));
  xor_4  g24111(.A(new_n16167_1), .B(new_n16169), .Y(new_n26460));
  xor_4  g24112(.A(new_n26460), .B(new_n16259), .Y(n13754));
  nand_5 g24113(.A(new_n2943), .B(new_n2942), .Y(new_n26462));
  xnor_4 g24114(.A(new_n26462), .B(new_n2986), .Y(n13764));
  xor_4  g24115(.A(new_n16423), .B(new_n16419_1), .Y(new_n26464));
  xor_4  g24116(.A(new_n26464), .B(new_n16415), .Y(n13798));
  nand_5 g24117(.A(new_n19920), .B(new_n19919), .Y(new_n26466));
  xor_4  g24118(.A(new_n26466), .B(new_n19937), .Y(n13835));
  nand_5 g24119(.A(new_n18084), .B(new_n18083), .Y(new_n26468));
  xnor_4 g24120(.A(new_n26468), .B(new_n18094), .Y(n13850));
  xor_4  g24121(.A(new_n20479), .B(new_n8917), .Y(n13922));
  nand_5 g24122(.A(new_n22143), .B(new_n22144_1), .Y(new_n26471));
  xor_4  g24123(.A(new_n26471), .B(new_n22154), .Y(n13923));
  nand_5 g24124(.A(new_n13453_1), .B(new_n13452), .Y(new_n26473));
  xor_4  g24125(.A(new_n26473), .B(new_n13477_1), .Y(n14004));
  nand_5 g24126(.A(new_n13676), .B(new_n13674), .Y(new_n26475));
  xnor_4 g24127(.A(new_n26475), .B(new_n13735), .Y(n14036));
  nand_5 g24128(.A(new_n24390), .B(new_n24389), .Y(new_n26477));
  xor_4  g24129(.A(new_n26477), .B(new_n24404), .Y(n14059));
  nand_5 g24130(.A(new_n19699), .B(new_n19698), .Y(new_n26479));
  xnor_4 g24131(.A(new_n26479), .B(new_n19701_1), .Y(n14081));
  nand_5 g24132(.A(new_n21564), .B(new_n21563), .Y(new_n26481));
  xor_4  g24133(.A(new_n26481), .B(new_n21567), .Y(n14095));
  xor_4  g24134(.A(new_n7693_1), .B(new_n3656), .Y(n14107));
  nor_5  g24135(.A(new_n10198), .B(new_n10197), .Y(new_n26484));
  xor_4  g24136(.A(new_n26484), .B(new_n10242), .Y(n14121));
  xor_4  g24137(.A(new_n13958), .B(new_n13957), .Y(n14126));
  nand_5 g24138(.A(new_n22413), .B(new_n22414), .Y(new_n26487));
  xnor_4 g24139(.A(new_n26487), .B(new_n22450), .Y(n14136));
  nor_5  g24140(.A(new_n26336), .B(new_n25237), .Y(new_n26489));
  and_5  g24141(.A(new_n26336), .B(new_n25237), .Y(new_n26490));
  nor_5  g24142(.A(new_n26490), .B(new_n26489), .Y(new_n26491));
  nor_5  g24143(.A(new_n26342), .B(new_n26339), .Y(new_n26492_1));
  nor_5  g24144(.A(new_n26492_1), .B(new_n26337), .Y(new_n26493));
  xor_4  g24145(.A(new_n26493), .B(new_n26491), .Y(n14147));
  nand_5 g24146(.A(new_n24056), .B(new_n24057), .Y(new_n26495));
  xor_4  g24147(.A(new_n26495), .B(new_n24102), .Y(n14174));
  nand_5 g24148(.A(new_n18889), .B(new_n18888), .Y(new_n26497));
  xnor_4 g24149(.A(new_n26497), .B(new_n18915), .Y(n14190));
  nand_5 g24150(.A(new_n6092), .B(new_n6091), .Y(new_n26499));
  xor_4  g24151(.A(new_n26499), .B(new_n6124), .Y(n14211));
  nand_5 g24152(.A(new_n19128), .B(new_n19127), .Y(new_n26501));
  xnor_4 g24153(.A(new_n26501), .B(new_n19131), .Y(n14222));
  nor_5  g24154(.A(new_n15422), .B(new_n15420), .Y(new_n26503));
  xor_4  g24155(.A(new_n26503), .B(new_n15472), .Y(n14267));
  nand_5 g24156(.A(new_n6481), .B(new_n6480), .Y(new_n26505));
  xnor_4 g24157(.A(new_n26505), .B(new_n6497), .Y(n14271));
  nand_5 g24158(.A(new_n10794), .B(new_n10795), .Y(new_n26507));
  xnor_4 g24159(.A(new_n26507), .B(new_n10809), .Y(n14277));
  nand_5 g24160(.A(new_n9603), .B(new_n9601), .Y(new_n26509));
  xor_4  g24161(.A(new_n26509), .B(new_n9613), .Y(n14294));
  nand_5 g24162(.A(new_n25898), .B(new_n25897), .Y(new_n26511));
  xnor_4 g24163(.A(new_n26511), .B(new_n25937), .Y(n14310));
  nand_5 g24164(.A(new_n25953), .B(new_n25954), .Y(new_n26513));
  xnor_4 g24165(.A(new_n26513), .B(new_n25956), .Y(n14326));
  nand_5 g24166(.A(new_n14261), .B(new_n14262), .Y(new_n26515_1));
  xor_4  g24167(.A(new_n26515_1), .B(new_n14321), .Y(n14342));
  nand_5 g24168(.A(new_n21014), .B(new_n21013), .Y(new_n26517));
  xnor_4 g24169(.A(new_n26517), .B(new_n21026), .Y(n14353));
  nor_5  g24170(.A(new_n24406_1), .B(new_n24385), .Y(new_n26519));
  nor_5  g24171(.A(new_n26519), .B(new_n24383), .Y(new_n26520));
  nor_5  g24172(.A(new_n24384), .B(new_n13503), .Y(new_n26521));
  nor_5  g24173(.A(new_n26521), .B(new_n26520), .Y(new_n26522));
  nor_5  g24174(.A(new_n24382), .B(new_n13506_1), .Y(new_n26523));
  nor_5  g24175(.A(new_n26523), .B(new_n26519), .Y(new_n26524));
  nor_5  g24176(.A(new_n26524), .B(new_n26522), .Y(n14364));
  nand_5 g24177(.A(new_n24923), .B(new_n24924), .Y(new_n26526));
  xor_4  g24178(.A(new_n26526), .B(new_n24926), .Y(n14375));
  nand_5 g24179(.A(new_n25367), .B(new_n25366), .Y(new_n26528));
  xor_4  g24180(.A(new_n26528), .B(new_n25392), .Y(n14412));
  nor_5  g24181(.A(new_n20211), .B(new_n7082), .Y(new_n26530));
  nor_5  g24182(.A(new_n26530), .B(new_n13411), .Y(new_n26531));
  and_5  g24183(.A(new_n26530), .B(new_n13411), .Y(new_n26532));
  nor_5  g24184(.A(new_n26532), .B(new_n26531), .Y(new_n26533));
  nand_5 g24185(.A(new_n20242), .B(new_n20215), .Y(new_n26534));
  nand_5 g24186(.A(new_n26534), .B(new_n20213_1), .Y(new_n26535));
  xor_4  g24187(.A(new_n26535), .B(new_n26533), .Y(n14414));
  xor_4  g24188(.A(new_n17820_1), .B(new_n17819), .Y(n14457));
  nand_5 g24189(.A(new_n5609_1), .B(new_n5608), .Y(new_n26538_1));
  xor_4  g24190(.A(new_n26538_1), .B(new_n5651), .Y(n14464));
  nand_5 g24191(.A(new_n12598), .B(new_n12599), .Y(new_n26540));
  xnor_4 g24192(.A(new_n26540), .B(new_n12623), .Y(n14471));
  nand_5 g24193(.A(new_n22495), .B(new_n22485), .Y(new_n26542));
  not_8  g24194(.A(new_n26542), .Y(new_n26543));
  nor_5  g24195(.A(new_n26543), .B(new_n26354), .Y(new_n26544));
  nor_5  g24196(.A(new_n26542), .B(new_n26352), .Y(new_n26545));
  nor_5  g24197(.A(new_n26545), .B(new_n26544), .Y(new_n26546));
  nand_5 g24198(.A(new_n26366), .B(new_n26355), .Y(new_n26547));
  nand_5 g24199(.A(new_n26547), .B(new_n26353_1), .Y(new_n26548));
  not_8  g24200(.A(new_n26548), .Y(new_n26549));
  xor_4  g24201(.A(new_n26549), .B(new_n26546), .Y(n14475));
  nand_5 g24202(.A(new_n14304), .B(new_n14305), .Y(new_n26551));
  xor_4  g24203(.A(new_n26551), .B(new_n14307), .Y(n14541));
  nand_5 g24204(.A(new_n24674), .B(new_n24666), .Y(new_n26553_1));
  nand_5 g24205(.A(new_n26553_1), .B(new_n24665), .Y(n14546));
  nand_5 g24206(.A(new_n12869), .B(new_n12868), .Y(new_n26555));
  xor_4  g24207(.A(new_n26555), .B(new_n12871_1), .Y(n14547));
  nand_5 g24208(.A(new_n14674), .B(new_n14673), .Y(new_n26557));
  xor_4  g24209(.A(new_n26557), .B(new_n14698), .Y(n14593));
  nand_5 g24210(.A(new_n10782), .B(new_n10783), .Y(new_n26559));
  xnor_4 g24211(.A(new_n26559), .B(new_n10813), .Y(n14636));
  nand_5 g24212(.A(new_n26109), .B(new_n26108), .Y(new_n26561));
  xnor_4 g24213(.A(new_n26561), .B(new_n26123), .Y(n14701));
  nand_5 g24214(.A(new_n14065), .B(new_n14066), .Y(new_n26563));
  xnor_4 g24215(.A(new_n26563), .B(new_n14076), .Y(n14734));
  nand_5 g24216(.A(new_n8211), .B(new_n8210), .Y(new_n26565_1));
  xor_4  g24217(.A(new_n26565_1), .B(new_n8267_1), .Y(n14746));
  xor_4  g24218(.A(new_n11209), .B(new_n11208), .Y(n14763));
  nand_5 g24219(.A(new_n25597), .B(new_n25596), .Y(new_n26568));
  xor_4  g24220(.A(new_n26568), .B(new_n25609), .Y(n14772));
  nand_5 g24221(.A(new_n24922), .B(new_n24921), .Y(new_n26570));
  xor_4  g24222(.A(new_n26570), .B(new_n24928), .Y(n14801));
  or_5   g24223(.A(new_n24433), .B(new_n24432), .Y(new_n26572_1));
  xor_4  g24224(.A(new_n26572_1), .B(new_n24455), .Y(n14819));
  nand_5 g24225(.A(new_n16708), .B(new_n16706), .Y(new_n26574));
  xor_4  g24226(.A(new_n26574), .B(new_n16756), .Y(n14827));
  nand_5 g24227(.A(new_n23777), .B(new_n23776), .Y(new_n26576));
  xnor_4 g24228(.A(new_n26576), .B(new_n23779), .Y(n14839));
  nand_5 g24229(.A(new_n19928), .B(new_n19927), .Y(new_n26578));
  xor_4  g24230(.A(new_n26578), .B(new_n19929), .Y(n14849));
  not_8  g24231(.A(new_n23617), .Y(new_n26580));
  nor_5  g24232(.A(new_n23682), .B(new_n26580), .Y(new_n26581));
  nand_5 g24233(.A(new_n23616), .B(new_n23610), .Y(new_n26582));
  nor_5  g24234(.A(new_n26582), .B(new_n26581), .Y(n14891));
  xor_4  g24235(.A(new_n7390_1), .B(new_n5266), .Y(n14931));
  nor_5  g24236(.A(new_n26535), .B(new_n26531), .Y(new_n26585));
  not_8  g24237(.A(new_n26535), .Y(new_n26586));
  nor_5  g24238(.A(new_n26586), .B(new_n26532), .Y(new_n26587));
  nor_5  g24239(.A(new_n26587), .B(new_n26585), .Y(n14944));
  xor_4  g24240(.A(new_n21022), .B(new_n10256), .Y(n14977));
  nor_5  g24241(.A(new_n14648), .B(new_n14647), .Y(new_n26590_1));
  xor_4  g24242(.A(new_n26590_1), .B(new_n14707), .Y(n14989));
  nand_5 g24243(.A(new_n12498), .B(new_n12496), .Y(new_n26592));
  xor_4  g24244(.A(new_n26592), .B(new_n12509), .Y(n15002));
  nand_5 g24245(.A(new_n25450), .B(new_n25451), .Y(new_n26594));
  xor_4  g24246(.A(new_n26594), .B(new_n6494), .Y(n15004));
  nand_5 g24247(.A(new_n10391), .B(new_n10390_1), .Y(new_n26596));
  xor_4  g24248(.A(new_n26596), .B(new_n10444), .Y(n15011));
  nand_5 g24249(.A(new_n25502), .B(new_n25501), .Y(new_n26598_1));
  xor_4  g24250(.A(new_n26598_1), .B(new_n25504), .Y(n15019));
  nand_5 g24251(.A(new_n17592_1), .B(new_n17570), .Y(new_n26600));
  nand_5 g24252(.A(new_n26600), .B(new_n17569), .Y(n15031));
  xor_4  g24253(.A(new_n20481), .B(new_n20479), .Y(n15033));
  xor_4  g24254(.A(new_n13834), .B(new_n8282), .Y(n15052));
  nand_5 g24255(.A(new_n22350), .B(new_n22348), .Y(new_n26604));
  xnor_4 g24256(.A(new_n26604), .B(new_n22338), .Y(n15082));
  nand_5 g24257(.A(new_n9392), .B(new_n9391), .Y(new_n26606));
  xnor_4 g24258(.A(new_n26606), .B(new_n9409), .Y(n15094));
  nand_5 g24259(.A(new_n13523), .B(new_n13524), .Y(new_n26608));
  xnor_4 g24260(.A(new_n26608), .B(new_n13526), .Y(n15118));
  nand_5 g24261(.A(new_n26320), .B(new_n26319), .Y(new_n26610));
  xor_4  g24262(.A(new_n26610), .B(new_n26322), .Y(n15128));
  nand_5 g24263(.A(new_n21401), .B(new_n21400), .Y(new_n26612));
  xor_4  g24264(.A(new_n26612), .B(new_n21452), .Y(n15139));
  or_5   g24265(.A(new_n19248), .B(new_n19246), .Y(new_n26614));
  xor_4  g24266(.A(new_n26614), .B(new_n19242), .Y(n15145));
  nand_5 g24267(.A(new_n16959), .B(new_n16957), .Y(new_n26616));
  xor_4  g24268(.A(new_n26616), .B(new_n16995), .Y(n15165));
  xor_4  g24269(.A(new_n17482), .B(new_n5698), .Y(n15176));
  nand_5 g24270(.A(new_n23106), .B(new_n23105), .Y(new_n26619));
  xnor_4 g24271(.A(new_n26619), .B(new_n23108), .Y(n15180));
  nand_5 g24272(.A(new_n18590), .B(new_n18591), .Y(new_n26621));
  xnor_4 g24273(.A(new_n26621), .B(new_n18625), .Y(n15205));
  xor_4  g24274(.A(new_n6114), .B(new_n18608), .Y(n15230));
  nand_5 g24275(.A(new_n19519), .B(new_n19520), .Y(new_n26624));
  xor_4  g24276(.A(new_n26624), .B(new_n19521), .Y(n15255));
  nand_5 g24277(.A(new_n11175), .B(new_n11176), .Y(new_n26626));
  xor_4  g24278(.A(new_n26626), .B(new_n11220_1), .Y(n15275));
  nand_5 g24279(.A(new_n15997), .B(new_n15996), .Y(new_n26628));
  xor_4  g24280(.A(new_n26628), .B(new_n16000), .Y(n15300));
  nor_5  g24281(.A(new_n26041), .B(new_n26039), .Y(new_n26630));
  nor_5  g24282(.A(new_n26040), .B(new_n26038), .Y(new_n26631));
  nor_5  g24283(.A(new_n26631), .B(new_n26630), .Y(new_n26632));
  xor_4  g24284(.A(new_n26632), .B(new_n24619), .Y(new_n26633));
  nand_5 g24285(.A(new_n26055), .B(new_n26044), .Y(new_n26634));
  nand_5 g24286(.A(new_n26634), .B(new_n26045), .Y(new_n26635));
  xor_4  g24287(.A(new_n26635), .B(new_n26633), .Y(n15307));
  nand_5 g24288(.A(new_n22808), .B(new_n22806), .Y(new_n26637));
  xnor_4 g24289(.A(new_n26637), .B(new_n22864), .Y(n15327));
  nor_5  g24290(.A(new_n22841), .B(new_n22840), .Y(new_n26639));
  xor_4  g24291(.A(new_n26639), .B(new_n22850), .Y(n15345));
  nand_5 g24292(.A(new_n14682), .B(new_n14681), .Y(new_n26641));
  xor_4  g24293(.A(new_n26641), .B(new_n14696), .Y(n15353));
  xor_4  g24294(.A(new_n26159_1), .B(new_n26149), .Y(n15366));
  xnor_4 g24295(.A(new_n26313), .B(new_n26311), .Y(n15382));
  nand_5 g24296(.A(new_n10613), .B(new_n10611_1), .Y(new_n26645));
  xnor_4 g24297(.A(new_n26645), .B(new_n10637), .Y(n15407));
  xor_4  g24298(.A(new_n17146), .B(new_n15528), .Y(n15428));
  not_8  g24299(.A(new_n25877_1), .Y(new_n26648));
  nor_5  g24300(.A(new_n26648), .B(new_n25875), .Y(new_n26649));
  nor_5  g24301(.A(new_n25939), .B(new_n25889), .Y(new_n26650));
  nor_5  g24302(.A(new_n26650), .B(new_n25890), .Y(new_n26651));
  nor_5  g24303(.A(new_n26651), .B(new_n26649), .Y(new_n26652));
  nor_5  g24304(.A(new_n25879), .B(new_n12822), .Y(new_n26653));
  nand_5 g24305(.A(new_n25887), .B(new_n26653), .Y(new_n26654));
  nor_5  g24306(.A(new_n26654), .B(new_n26649), .Y(new_n26655));
  nor_5  g24307(.A(new_n26655), .B(new_n26650), .Y(new_n26656_1));
  nor_5  g24308(.A(new_n26656_1), .B(new_n26652), .Y(n15435));
  nand_5 g24309(.A(new_n25477), .B(new_n25466), .Y(new_n26658));
  nand_5 g24310(.A(new_n26658), .B(new_n25468_1), .Y(new_n26659));
  xnor_4 g24311(.A(new_n26659), .B(new_n25465), .Y(n15438));
  nand_5 g24312(.A(new_n25906), .B(new_n25905), .Y(new_n26661));
  xnor_4 g24313(.A(new_n26661), .B(new_n25933), .Y(n15465));
  xor_4  g24314(.A(new_n18534), .B(new_n7593_1), .Y(n15467));
  nand_5 g24315(.A(new_n9021), .B(new_n9020), .Y(new_n26664));
  xor_4  g24316(.A(new_n26664), .B(new_n9100), .Y(n15470));
  nand_5 g24317(.A(new_n16698), .B(new_n16697), .Y(new_n26666));
  xnor_4 g24318(.A(new_n26666), .B(new_n16761), .Y(n15477));
  nand_5 g24319(.A(new_n26222), .B(new_n26221), .Y(new_n26668));
  xnor_4 g24320(.A(new_n26668), .B(new_n26230), .Y(n15481));
  nand_5 g24321(.A(new_n17265), .B(new_n17264), .Y(new_n26670));
  xnor_4 g24322(.A(new_n26670), .B(new_n17267), .Y(n15496));
  nor_5  g24323(.A(new_n13926), .B(new_n13925), .Y(new_n26672));
  xor_4  g24324(.A(new_n26672), .B(new_n13969), .Y(n15501));
  nand_5 g24325(.A(new_n21560), .B(new_n21559), .Y(new_n26674_1));
  xnor_4 g24326(.A(new_n26674_1), .B(new_n21570), .Y(n15555));
  nand_5 g24327(.A(new_n24244), .B(new_n24243), .Y(new_n26676));
  xor_4  g24328(.A(new_n26676), .B(new_n24258_1), .Y(n15558));
  nand_5 g24329(.A(new_n25342), .B(new_n25339), .Y(new_n26678));
  nand_5 g24330(.A(new_n26678), .B(new_n25338), .Y(n15559));
  nand_5 g24331(.A(new_n23196), .B(new_n23181), .Y(new_n26680));
  nand_5 g24332(.A(new_n26680), .B(new_n23180), .Y(new_n26681_1));
  nor_5  g24333(.A(new_n26681_1), .B(new_n24653), .Y(new_n26682));
  nand_5 g24334(.A(new_n23229), .B(new_n23199), .Y(new_n26683));
  nand_5 g24335(.A(new_n26683), .B(new_n23198), .Y(new_n26684));
  nor_5  g24336(.A(new_n26684), .B(new_n26682), .Y(new_n26685));
  and_5  g24337(.A(new_n26681_1), .B(new_n25548), .Y(new_n26686));
  nor_5  g24338(.A(new_n26686), .B(new_n26685), .Y(new_n26687));
  and_5  g24339(.A(new_n26681_1), .B(new_n24653), .Y(new_n26688));
  nor_5  g24340(.A(new_n26688), .B(new_n26685), .Y(new_n26689));
  nor_5  g24341(.A(new_n26681_1), .B(new_n25548), .Y(new_n26690));
  nor_5  g24342(.A(new_n26690), .B(new_n26689), .Y(new_n26691));
  nor_5  g24343(.A(new_n26691), .B(new_n26687), .Y(n15570));
  nand_5 g24344(.A(new_n14242), .B(new_n14241), .Y(new_n26693));
  xnor_4 g24345(.A(new_n26693), .B(new_n14327), .Y(n15573));
  nor_5  g24346(.A(new_n13424_1), .B(new_n13423), .Y(new_n26695));
  xor_4  g24347(.A(new_n26695), .B(new_n13488), .Y(n15588));
  nand_5 g24348(.A(new_n24441), .B(new_n24440), .Y(new_n26697));
  xor_4  g24349(.A(new_n26697), .B(new_n24451), .Y(n15590));
  nand_5 g24350(.A(new_n25089), .B(new_n25088), .Y(new_n26699));
  xor_4  g24351(.A(new_n26699), .B(new_n25100), .Y(n15598));
  nand_5 g24352(.A(new_n10776), .B(new_n10777), .Y(new_n26701));
  xnor_4 g24353(.A(new_n26701), .B(new_n10815), .Y(n15614));
  nand_5 g24354(.A(new_n25589), .B(new_n25588), .Y(new_n26703));
  xnor_4 g24355(.A(new_n26703), .B(new_n25614_1), .Y(n15662));
  nand_5 g24356(.A(new_n3631), .B(new_n3632), .Y(new_n26705));
  xnor_4 g24357(.A(new_n26705), .B(new_n3675), .Y(n15716));
  nand_5 g24358(.A(new_n16573), .B(new_n16572), .Y(new_n26707_1));
  xor_4  g24359(.A(new_n26707_1), .B(new_n16619), .Y(n15749));
  nand_5 g24360(.A(new_n21468), .B(new_n21469), .Y(new_n26709));
  xnor_4 g24361(.A(new_n26709), .B(new_n21471_1), .Y(n15762));
  nor_5  g24362(.A(new_n9071), .B(new_n9068), .Y(new_n26711));
  nor_5  g24363(.A(new_n26711), .B(new_n9073), .Y(n15793));
  nand_5 g24364(.A(new_n25373), .B(new_n25372), .Y(new_n26713));
  xor_4  g24365(.A(new_n26713), .B(new_n25386), .Y(n15812));
  nand_5 g24366(.A(new_n14254), .B(new_n14255), .Y(new_n26715));
  xor_4  g24367(.A(new_n26715), .B(new_n14323_1), .Y(n15815));
  or_5   g24368(.A(new_n9609), .B(new_n9607), .Y(new_n26717));
  xor_4  g24369(.A(new_n26717), .B(new_n9611), .Y(n15816));
  nand_5 g24370(.A(new_n13824), .B(new_n13823), .Y(new_n26719_1));
  xor_4  g24371(.A(new_n26719_1), .B(new_n13839), .Y(n15831));
  nor_5  g24372(.A(new_n11052), .B(new_n11050), .Y(new_n26721));
  xor_4  g24373(.A(new_n26721), .B(new_n8288_1), .Y(n15846));
  nand_5 g24374(.A(new_n9645), .B(new_n9644), .Y(new_n26723));
  xor_4  g24375(.A(new_n26723), .B(new_n9660), .Y(n15859));
  nand_5 g24376(.A(new_n22720), .B(new_n22704), .Y(new_n26725_1));
  nand_5 g24377(.A(new_n26725_1), .B(new_n22705), .Y(new_n26726));
  nor_5  g24378(.A(new_n26726), .B(new_n9274), .Y(new_n26727_1));
  not_8  g24379(.A(new_n26727_1), .Y(new_n26728));
  nand_5 g24380(.A(new_n26728), .B(new_n22975), .Y(new_n26729_1));
  nand_5 g24381(.A(new_n26727_1), .B(new_n22976), .Y(new_n26730));
  nand_5 g24382(.A(new_n26730), .B(new_n26729_1), .Y(new_n26731));
  nand_5 g24383(.A(new_n26726), .B(new_n9274), .Y(new_n26732));
  nand_5 g24384(.A(new_n26732), .B(new_n26728), .Y(new_n26733));
  or_5   g24385(.A(new_n26733), .B(new_n22977), .Y(new_n26734));
  nand_5 g24386(.A(new_n26733), .B(new_n22977), .Y(new_n26735));
  nand_5 g24387(.A(new_n22751), .B(new_n22723), .Y(new_n26736));
  nand_5 g24388(.A(new_n26736), .B(new_n22722), .Y(new_n26737));
  nand_5 g24389(.A(new_n26737), .B(new_n26735), .Y(new_n26738));
  nand_5 g24390(.A(new_n26738), .B(new_n26734), .Y(new_n26739));
  xnor_4 g24391(.A(new_n26739), .B(new_n26731), .Y(n15869));
  nand_5 g24392(.A(new_n21581), .B(new_n21582), .Y(new_n26741));
  xor_4  g24393(.A(new_n26741), .B(new_n21609), .Y(n15885));
  nor_5  g24394(.A(new_n24052_1), .B(new_n17843), .Y(new_n26743));
  nor_5  g24395(.A(new_n26743), .B(new_n24104), .Y(new_n26744_1));
  xor_4  g24396(.A(new_n26744_1), .B(new_n24052_1), .Y(n15889));
  nand_5 g24397(.A(new_n21596), .B(new_n21597), .Y(new_n26746));
  xor_4  g24398(.A(new_n26746), .B(new_n15847), .Y(n15917));
  xor_4  g24399(.A(new_n15840), .B(new_n15839), .Y(n15922));
  xor_4  g24400(.A(new_n8245), .B(new_n8243), .Y(n15947));
  nand_5 g24401(.A(new_n23701), .B(new_n23691), .Y(new_n26750));
  xor_4  g24402(.A(new_n26750), .B(new_n22295), .Y(new_n26751));
  nand_5 g24403(.A(new_n23716), .B(new_n23705), .Y(new_n26752_1));
  nand_5 g24404(.A(new_n26752_1), .B(new_n23706), .Y(new_n26753));
  xor_4  g24405(.A(new_n26753), .B(new_n26751), .Y(n15956));
  xor_4  g24406(.A(new_n15581), .B(new_n15579), .Y(n15958));
  xor_4  g24407(.A(new_n19562), .B(new_n19555), .Y(new_n26756));
  and_5  g24408(.A(new_n26756), .B(new_n19556), .Y(n15986));
  nand_5 g24409(.A(new_n26049), .B(new_n26050), .Y(new_n26758));
  xor_4  g24410(.A(new_n26758), .B(new_n26053_1), .Y(n16013));
  nand_5 g24411(.A(new_n24889), .B(new_n24878), .Y(new_n26760));
  nand_5 g24412(.A(new_n26760), .B(new_n24877), .Y(new_n26761));
  or_5   g24413(.A(new_n26750), .B(new_n24876), .Y(new_n26762));
  nand_5 g24414(.A(new_n26750), .B(new_n24876), .Y(new_n26763));
  nand_5 g24415(.A(new_n26763), .B(new_n26762), .Y(new_n26764));
  xnor_4 g24416(.A(new_n26764), .B(new_n26761), .Y(n16060));
  nand_5 g24417(.A(new_n18829), .B(new_n9943), .Y(new_n26766));
  nand_5 g24418(.A(new_n18831_1), .B(n25972), .Y(new_n26767));
  nand_5 g24419(.A(new_n25677), .B(new_n25675), .Y(new_n26768));
  nand_5 g24420(.A(new_n26768), .B(new_n25676), .Y(new_n26769));
  not_8  g24421(.A(new_n26769), .Y(new_n26770));
  nand_5 g24422(.A(new_n26770), .B(new_n26767), .Y(new_n26771));
  nand_5 g24423(.A(new_n26771), .B(new_n26766), .Y(new_n26772));
  not_8  g24424(.A(new_n26772), .Y(new_n26773));
  nand_5 g24425(.A(new_n26773), .B(new_n25778), .Y(new_n26774));
  not_8  g24426(.A(new_n26774), .Y(new_n26775_1));
  nor_5  g24427(.A(new_n26773), .B(new_n25778), .Y(new_n26776));
  nor_5  g24428(.A(new_n26776), .B(new_n26775_1), .Y(new_n26777));
  nand_5 g24429(.A(new_n26777), .B(new_n25888), .Y(new_n26778));
  or_5   g24430(.A(new_n26777), .B(new_n25888), .Y(new_n26779));
  nand_5 g24431(.A(new_n26766), .B(new_n26767), .Y(new_n26780_1));
  xor_4  g24432(.A(new_n26780_1), .B(new_n26770), .Y(new_n26781));
  nand_5 g24433(.A(new_n26781), .B(new_n25895), .Y(new_n26782));
  or_5   g24434(.A(new_n26781), .B(new_n25895), .Y(new_n26783));
  nand_5 g24435(.A(new_n25681), .B(new_n25663), .Y(new_n26784));
  nand_5 g24436(.A(new_n26784), .B(new_n25680), .Y(new_n26785));
  nand_5 g24437(.A(new_n26785), .B(new_n26783), .Y(new_n26786));
  nand_5 g24438(.A(new_n26786), .B(new_n26782), .Y(new_n26787));
  nand_5 g24439(.A(new_n26787), .B(new_n26779), .Y(new_n26788));
  nand_5 g24440(.A(new_n26788), .B(new_n26778), .Y(new_n26789));
  xor_4  g24441(.A(new_n26775_1), .B(new_n26654), .Y(new_n26790));
  xor_4  g24442(.A(new_n26790), .B(new_n26789), .Y(n16062));
  nand_5 g24443(.A(new_n26151), .B(new_n26150), .Y(new_n26792));
  xor_4  g24444(.A(new_n26792), .B(new_n26157), .Y(n16068));
  nand_5 g24445(.A(new_n26421), .B(new_n26420), .Y(new_n26794_1));
  xor_4  g24446(.A(new_n26794_1), .B(new_n26423), .Y(n16080));
  nand_5 g24447(.A(new_n25790), .B(new_n25787), .Y(new_n26796));
  nand_5 g24448(.A(new_n26796), .B(new_n25786), .Y(new_n26797_1));
  nand_5 g24449(.A(new_n25784_1), .B(new_n25780), .Y(new_n26798));
  and_5  g24450(.A(new_n26798), .B(new_n25781), .Y(new_n26799));
  xnor_4 g24451(.A(new_n26799), .B(new_n26797_1), .Y(n16098));
  nand_5 g24452(.A(new_n20167), .B(new_n20166), .Y(new_n26801_1));
  xor_4  g24453(.A(new_n26801_1), .B(new_n20177), .Y(n16110));
  nand_5 g24454(.A(new_n17373), .B(new_n17375), .Y(new_n26803));
  xor_4  g24455(.A(new_n26803), .B(new_n17407), .Y(n16142));
  nand_5 g24456(.A(new_n19036), .B(new_n19037), .Y(new_n26805));
  xor_4  g24457(.A(new_n26805), .B(new_n19051), .Y(n16185));
  nand_5 g24458(.A(new_n14343), .B(new_n14342_1), .Y(new_n26807));
  xor_4  g24459(.A(new_n26807), .B(new_n14360), .Y(n16196));
  nand_5 g24460(.A(new_n23727), .B(new_n23728), .Y(new_n26809));
  xor_4  g24461(.A(new_n26809), .B(new_n23730), .Y(n16206));
  nand_5 g24462(.A(new_n23809), .B(new_n23808), .Y(new_n26811));
  xor_4  g24463(.A(new_n26811), .B(new_n23812), .Y(n16215));
  nand_5 g24464(.A(new_n21714), .B(new_n21713), .Y(new_n26813));
  xor_4  g24465(.A(new_n26813), .B(new_n21724), .Y(n16218));
  nor_5  g24466(.A(new_n4265), .B(new_n4264), .Y(new_n26815_1));
  nor_5  g24467(.A(new_n26815_1), .B(new_n4266_1), .Y(n16219));
  nand_5 g24468(.A(new_n7931), .B(new_n7932), .Y(new_n26817));
  xnor_4 g24469(.A(new_n26817), .B(new_n7938), .Y(n16230));
  nand_5 g24470(.A(new_n9649), .B(new_n9648_1), .Y(new_n26819));
  xor_4  g24471(.A(new_n26819), .B(new_n9658), .Y(n16243));
  nand_5 g24472(.A(new_n19878), .B(new_n19879), .Y(new_n26821));
  xor_4  g24473(.A(new_n26821), .B(new_n19889), .Y(n16275));
  nand_5 g24474(.A(new_n11781), .B(new_n11782), .Y(new_n26823_1));
  xor_4  g24475(.A(new_n26823_1), .B(new_n11824), .Y(n16279));
  nand_5 g24476(.A(new_n23343), .B(new_n23275), .Y(new_n26825));
  nand_5 g24477(.A(new_n26825), .B(new_n23274), .Y(n16322));
  nand_5 g24478(.A(new_n19853), .B(new_n19852), .Y(new_n26827));
  xor_4  g24479(.A(new_n26827), .B(new_n19897), .Y(n16327));
  nand_5 g24480(.A(new_n24248), .B(new_n24247), .Y(new_n26829));
  xor_4  g24481(.A(new_n26829), .B(new_n24254), .Y(n16350));
  xor_4  g24482(.A(new_n7593_1), .B(new_n19083), .Y(n16367));
  nand_5 g24483(.A(new_n21829), .B(new_n21828), .Y(new_n26832));
  xnor_4 g24484(.A(new_n26832), .B(new_n21857), .Y(n16379));
  nand_5 g24485(.A(new_n22833), .B(new_n22831), .Y(new_n26834));
  xnor_4 g24486(.A(new_n26834), .B(new_n22854), .Y(n16398));
  nand_5 g24487(.A(new_n15536), .B(new_n15537), .Y(new_n26836));
  xor_4  g24488(.A(new_n26836), .B(new_n15539_1), .Y(n16406));
  nand_5 g24489(.A(new_n25104), .B(new_n25082), .Y(new_n26838));
  xor_4  g24490(.A(new_n26838), .B(new_n25102), .Y(n16407));
  nand_5 g24491(.A(new_n26779), .B(new_n26778), .Y(new_n26840));
  xnor_4 g24492(.A(new_n26840), .B(new_n26787), .Y(n16419));
  nand_5 g24493(.A(new_n9578), .B(new_n9577), .Y(new_n26842));
  xor_4  g24494(.A(new_n26842), .B(new_n9625), .Y(n16424));
  nand_5 g24495(.A(new_n15965), .B(new_n15964), .Y(new_n26844));
  xor_4  g24496(.A(new_n26844), .B(new_n16014), .Y(n16428));
  nand_5 g24497(.A(new_n13792), .B(new_n13791), .Y(new_n26846));
  xor_4  g24498(.A(new_n26846), .B(new_n13855), .Y(n16433));
  nand_5 g24499(.A(new_n13800), .B(new_n13799), .Y(new_n26848));
  xor_4  g24500(.A(new_n26848), .B(new_n13851_1), .Y(n16440));
  nand_5 g24501(.A(new_n20163), .B(new_n20162), .Y(new_n26850));
  xor_4  g24502(.A(new_n26850), .B(new_n20179_1), .Y(n16445));
  nand_5 g24503(.A(new_n16183), .B(new_n16182), .Y(new_n26852));
  xor_4  g24504(.A(new_n26852), .B(new_n16255), .Y(n16460));
  nand_5 g24505(.A(new_n22736), .B(new_n22735), .Y(new_n26854));
  xnor_4 g24506(.A(new_n26854), .B(new_n22747), .Y(n16481));
  nor_5  g24507(.A(new_n16947), .B(new_n12817), .Y(new_n26856));
  xor_4  g24508(.A(new_n16949), .B(new_n12817), .Y(new_n26857));
  nand_5 g24509(.A(new_n23406), .B(new_n23391), .Y(new_n26858));
  nand_5 g24510(.A(new_n26858), .B(new_n23390), .Y(new_n26859));
  nor_5  g24511(.A(new_n26859), .B(new_n26857), .Y(new_n26860));
  nor_5  g24512(.A(new_n26860), .B(new_n26856), .Y(n16493));
  nand_5 g24513(.A(new_n5251), .B(new_n5250), .Y(new_n26862));
  xnor_4 g24514(.A(new_n26862), .B(new_n5285), .Y(n16506));
  nand_5 g24515(.A(new_n9707), .B(new_n6962), .Y(new_n26864));
  nand_5 g24516(.A(new_n26864), .B(new_n14777), .Y(new_n26865));
  xor_4  g24517(.A(new_n26865), .B(new_n14780), .Y(n16516));
  nand_5 g24518(.A(new_n25213), .B(new_n25212), .Y(new_n26867));
  xnor_4 g24519(.A(new_n26867), .B(new_n25215_1), .Y(n16517));
  xor_4  g24520(.A(new_n17962), .B(new_n6592), .Y(new_n26869));
  xor_4  g24521(.A(new_n26869), .B(new_n17967), .Y(n16527));
  nand_5 g24522(.A(new_n12501), .B(new_n10565), .Y(new_n26871));
  nand_5 g24523(.A(new_n26871), .B(new_n12502), .Y(n16554));
  xor_4  g24524(.A(new_n6969), .B(new_n6568), .Y(n16583));
  nor_5  g24525(.A(new_n24584), .B(new_n24582), .Y(new_n26874));
  xor_4  g24526(.A(new_n26874), .B(new_n24578), .Y(n16584));
  nand_5 g24527(.A(new_n21909), .B(new_n21907), .Y(new_n26876));
  xor_4  g24528(.A(new_n26876), .B(new_n21931), .Y(n16589));
  nand_5 g24529(.A(new_n22307), .B(new_n22310), .Y(new_n26878));
  xor_4  g24530(.A(new_n26878), .B(new_n22319), .Y(n16596));
  nand_5 g24531(.A(new_n25361), .B(new_n25360), .Y(new_n26880));
  xor_4  g24532(.A(new_n26880), .B(new_n25398), .Y(n16617));
  nand_5 g24533(.A(new_n8716_1), .B(new_n8715), .Y(new_n26882_1));
  xor_4  g24534(.A(new_n26882_1), .B(new_n8748), .Y(n16630));
  nand_5 g24535(.A(new_n25380), .B(new_n25379), .Y(new_n26884));
  xor_4  g24536(.A(new_n26884), .B(new_n5546), .Y(n16640));
  xor_4  g24537(.A(new_n2545), .B(new_n2544), .Y(n16656));
  nand_5 g24538(.A(new_n7892), .B(new_n7891), .Y(new_n26887));
  xnor_4 g24539(.A(new_n26887), .B(new_n7950_1), .Y(n16674));
  nand_5 g24540(.A(new_n16189), .B(new_n16188), .Y(new_n26889));
  xor_4  g24541(.A(new_n26889), .B(new_n16253), .Y(n16682));
  nand_5 g24542(.A(new_n25295), .B(new_n25294), .Y(new_n26891));
  xnor_4 g24543(.A(new_n26891), .B(new_n25315), .Y(n16684));
  nand_5 g24544(.A(new_n12181), .B(new_n12179_1), .Y(new_n26893));
  xor_4  g24545(.A(new_n26893), .B(new_n12183), .Y(n16688));
  nand_5 g24546(.A(new_n7269), .B(new_n7267), .Y(new_n26895));
  xnor_4 g24547(.A(new_n26895), .B(new_n7280_1), .Y(n16733));
  nand_5 g24548(.A(new_n9083), .B(new_n9082), .Y(new_n26897));
  xor_4  g24549(.A(new_n26897), .B(new_n9086), .Y(n16798));
  nand_5 g24550(.A(new_n19177), .B(new_n19176_1), .Y(new_n26899));
  xor_4  g24551(.A(new_n26899), .B(new_n19185), .Y(n16834));
  nand_5 g24552(.A(new_n3215), .B(new_n3214), .Y(new_n26901));
  xnor_4 g24553(.A(new_n26901), .B(new_n3268), .Y(n16837));
  nand_5 g24554(.A(new_n24883), .B(new_n24882), .Y(new_n26903));
  xor_4  g24555(.A(new_n26903), .B(new_n24886), .Y(n16841));
  nand_5 g24556(.A(new_n5696_1), .B(new_n5695), .Y(new_n26905_1));
  xor_4  g24557(.A(new_n26905_1), .B(new_n5703), .Y(n16885));
  nand_5 g24558(.A(new_n9425), .B(new_n9350), .Y(new_n26907));
  xnor_4 g24559(.A(new_n26907), .B(new_n9423_1), .Y(n16905));
  xor_4  g24560(.A(new_n24789), .B(new_n20772), .Y(n16951));
  nand_5 g24561(.A(new_n18602), .B(new_n18603), .Y(new_n26910));
  xnor_4 g24562(.A(new_n26910), .B(new_n18613), .Y(n16954));
  xor_4  g24563(.A(new_n9604), .B(new_n4043), .Y(n16989));
  nand_5 g24564(.A(new_n21825), .B(new_n21824), .Y(new_n26913_1));
  xnor_4 g24565(.A(new_n26913_1), .B(new_n21859), .Y(n17006));
  nand_5 g24566(.A(new_n15454), .B(new_n15453), .Y(new_n26915));
  xnor_4 g24567(.A(new_n26915), .B(new_n15456), .Y(n17068));
  nand_5 g24568(.A(new_n17397), .B(new_n17398), .Y(new_n26917));
  xor_4  g24569(.A(new_n26917), .B(new_n17399), .Y(n17070));
  or_5   g24570(.A(new_n23284), .B(new_n23283), .Y(new_n26919));
  xor_4  g24571(.A(new_n26919), .B(new_n23339), .Y(n17075));
  nand_5 g24572(.A(new_n19463), .B(new_n19464), .Y(new_n26921_1));
  xnor_4 g24573(.A(new_n26921_1), .B(new_n19490), .Y(n17084));
  nor_5  g24574(.A(new_n5278), .B(new_n5274_1), .Y(new_n26923_1));
  xor_4  g24575(.A(new_n26923_1), .B(new_n5276), .Y(n17104));
  nand_5 g24576(.A(new_n15174), .B(new_n15173), .Y(new_n26925));
  xnor_4 g24577(.A(new_n26925), .B(new_n15202), .Y(n17106));
  nand_5 g24578(.A(new_n11199), .B(new_n11200), .Y(new_n26927));
  xor_4  g24579(.A(new_n26927), .B(new_n11212), .Y(n17119));
  or_5   g24580(.A(new_n15062), .B(new_n15060), .Y(new_n26929_1));
  xor_4  g24581(.A(new_n26929_1), .B(new_n15102), .Y(n17130));
  nand_5 g24582(.A(new_n25914), .B(new_n25913), .Y(new_n26931));
  xnor_4 g24583(.A(new_n26931), .B(new_n25929), .Y(n17138));
  nand_5 g24584(.A(new_n25209_1), .B(new_n25208), .Y(new_n26933));
  xnor_4 g24585(.A(new_n26933), .B(new_n25217), .Y(n17163));
  nand_5 g24586(.A(new_n22903_1), .B(new_n22902), .Y(new_n26935));
  xnor_4 g24587(.A(new_n26935), .B(new_n22923), .Y(n17168));
  nand_5 g24588(.A(new_n13265), .B(new_n13264), .Y(new_n26937));
  xor_4  g24589(.A(new_n26937), .B(new_n13274), .Y(n17202));
  nand_5 g24590(.A(new_n22085), .B(new_n22084), .Y(new_n26939));
  xor_4  g24591(.A(new_n26939), .B(new_n22088), .Y(n17219));
  nand_5 g24592(.A(new_n21231), .B(new_n21230), .Y(new_n26941));
  xnor_4 g24593(.A(new_n26941), .B(new_n21269), .Y(n17232));
  nand_5 g24594(.A(new_n17529_1), .B(new_n17530), .Y(new_n26943_1));
  xor_4  g24595(.A(new_n26943_1), .B(new_n17532), .Y(n17236));
  nand_5 g24596(.A(new_n12044), .B(new_n12043), .Y(new_n26945));
  xor_4  g24597(.A(new_n26945), .B(new_n12101), .Y(n17243));
  nand_5 g24598(.A(new_n12858), .B(new_n12857), .Y(new_n26947));
  xor_4  g24599(.A(new_n26947), .B(new_n12875_1), .Y(n17263));
  nor_5  g24600(.A(new_n22300), .B(new_n22289), .Y(new_n26949));
  nor_5  g24601(.A(new_n22323), .B(new_n22296), .Y(new_n26950));
  nor_5  g24602(.A(new_n26950), .B(new_n26949), .Y(n17285));
  nand_5 g24603(.A(new_n13445), .B(new_n13444), .Y(new_n26952));
  xor_4  g24604(.A(new_n26952), .B(new_n13481), .Y(n17320));
  nand_5 g24605(.A(new_n2929_1), .B(new_n2928), .Y(new_n26954));
  xnor_4 g24606(.A(new_n26954), .B(new_n2990), .Y(n17337));
  nand_5 g24607(.A(new_n25015), .B(new_n25016), .Y(new_n26956));
  xnor_4 g24608(.A(new_n26956), .B(new_n25024), .Y(n17344));
  nand_5 g24609(.A(new_n25000), .B(new_n24999), .Y(new_n26958));
  xnor_4 g24610(.A(new_n26958), .B(new_n25032_1), .Y(n17359));
  nand_5 g24611(.A(new_n16236), .B(new_n24947), .Y(new_n26960));
  nand_5 g24612(.A(new_n26960), .B(new_n19538), .Y(n17387));
  nor_5  g24613(.A(new_n5702), .B(new_n5698), .Y(new_n26962));
  nor_5  g24614(.A(new_n26962), .B(new_n5704_1), .Y(n17391));
  nand_5 g24615(.A(new_n21833), .B(new_n21832_1), .Y(new_n26964));
  xnor_4 g24616(.A(new_n26964), .B(new_n21855), .Y(n17392));
  nand_5 g24617(.A(new_n25291), .B(new_n25290), .Y(new_n26966));
  xnor_4 g24618(.A(new_n26966), .B(new_n25317), .Y(n17421));
  nor_5  g24619(.A(new_n14012), .B(new_n14011), .Y(new_n26968));
  xor_4  g24620(.A(new_n26968), .B(new_n7454), .Y(n17432));
  nand_5 g24621(.A(new_n24072), .B(new_n24073), .Y(new_n26970_1));
  xor_4  g24622(.A(new_n26970_1), .B(new_n24094), .Y(n17436));
  xor_4  g24623(.A(new_n8243), .B(new_n5192), .Y(n17440));
  xor_4  g24624(.A(new_n9713), .B(new_n6567_1), .Y(n17450));
  not_8  g24625(.A(new_n8563_1), .Y(new_n26974));
  nor_5  g24626(.A(new_n26974), .B(new_n8475), .Y(new_n26975));
  nor_5  g24627(.A(new_n26975), .B(new_n8472), .Y(new_n26976));
  nor_5  g24628(.A(new_n21576), .B(new_n8474), .Y(new_n26977));
  nor_5  g24629(.A(new_n26977), .B(new_n26976), .Y(new_n26978));
  nor_5  g24630(.A(new_n21575), .B(new_n8471), .Y(new_n26979_1));
  nor_5  g24631(.A(new_n26979_1), .B(new_n26975), .Y(new_n26980));
  nor_5  g24632(.A(new_n26980), .B(new_n26978), .Y(n17461));
  nor_5  g24633(.A(new_n26362), .B(new_n26360), .Y(new_n26982));
  xor_4  g24634(.A(new_n26982), .B(new_n26364), .Y(n17466));
  nand_5 g24635(.A(new_n15425), .B(new_n15426), .Y(new_n26984));
  xnor_4 g24636(.A(new_n26984), .B(new_n15470_1), .Y(n17493));
  nand_5 g24637(.A(new_n24635), .B(new_n24634), .Y(new_n26986_1));
  xor_4  g24638(.A(new_n26986_1), .B(new_n24637), .Y(n17500));
  nand_5 g24639(.A(new_n25604), .B(new_n25601), .Y(new_n26988));
  xor_4  g24640(.A(new_n26988), .B(new_n25607), .Y(n17524));
  nand_5 g24641(.A(new_n6457_1), .B(new_n6456_1), .Y(new_n26990));
  xnor_4 g24642(.A(new_n26990), .B(new_n6505), .Y(n17529));
  nand_5 g24643(.A(new_n17182), .B(new_n17183), .Y(new_n26992));
  xor_4  g24644(.A(new_n26992), .B(new_n17185), .Y(n17557));
  nand_5 g24645(.A(new_n19020), .B(new_n19021), .Y(new_n26994));
  xor_4  g24646(.A(new_n26994), .B(new_n19059), .Y(n17583));
  nand_5 g24647(.A(new_n16213), .B(new_n16212), .Y(new_n26996));
  xor_4  g24648(.A(new_n26996), .B(new_n16245), .Y(n17592));
  nand_5 g24649(.A(new_n9598_1), .B(new_n9597), .Y(new_n26998));
  xor_4  g24650(.A(new_n26998), .B(new_n9615), .Y(n17638));
  nand_5 g24651(.A(new_n22730), .B(new_n22729), .Y(new_n27000));
  xnor_4 g24652(.A(new_n27000), .B(new_n22749), .Y(n17687));
  nor_5  g24653(.A(new_n15764), .B(new_n15763), .Y(new_n27002));
  xor_4  g24654(.A(new_n27002), .B(new_n15809), .Y(n17721));
  nand_5 g24655(.A(new_n24833), .B(new_n24832), .Y(new_n27004_1));
  xor_4  g24656(.A(new_n27004_1), .B(new_n24851), .Y(n17735));
  nor_5  g24657(.A(new_n24175), .B(new_n24168), .Y(new_n27006));
  nor_5  g24658(.A(new_n24176), .B(new_n24167_1), .Y(new_n27007));
  nor_5  g24659(.A(new_n27007), .B(new_n27006), .Y(new_n27008));
  nor_5  g24660(.A(new_n27008), .B(new_n24163), .Y(new_n27009));
  nand_5 g24661(.A(new_n24192), .B(new_n24178), .Y(new_n27010));
  nand_5 g24662(.A(new_n27010), .B(new_n24179), .Y(new_n27011_1));
  nor_5  g24663(.A(new_n27011_1), .B(new_n27009), .Y(new_n27012));
  not_8  g24664(.A(new_n27006), .Y(new_n27013));
  nand_5 g24665(.A(new_n27008), .B(new_n24163), .Y(new_n27014));
  nand_5 g24666(.A(new_n27014), .B(new_n27013), .Y(new_n27015));
  nor_5  g24667(.A(new_n27015), .B(new_n27012), .Y(n17738));
  nand_5 g24668(.A(new_n17620), .B(new_n17622), .Y(new_n27017));
  xor_4  g24669(.A(new_n27017), .B(new_n17624), .Y(n17746));
  nand_5 g24670(.A(new_n26117), .B(new_n26116), .Y(new_n27019_1));
  xnor_4 g24671(.A(new_n27019_1), .B(new_n26119), .Y(n17749));
  nor_5  g24672(.A(new_n21421), .B(new_n21420), .Y(new_n27021));
  xor_4  g24673(.A(new_n27021), .B(new_n21443), .Y(n17820));
  nand_5 g24674(.A(new_n16220), .B(new_n16219_1), .Y(new_n27023));
  xor_4  g24675(.A(new_n27023), .B(new_n16243_1), .Y(n17855));
  nor_5  g24676(.A(new_n5570), .B(new_n5494), .Y(new_n27025));
  nand_5 g24677(.A(new_n5570), .B(new_n25357), .Y(new_n27026));
  not_8  g24678(.A(new_n27026), .Y(new_n27027));
  nand_5 g24679(.A(new_n5661), .B(new_n5572), .Y(new_n27028));
  nand_5 g24680(.A(new_n27028), .B(new_n5573), .Y(new_n27029));
  nor_5  g24681(.A(new_n27029), .B(new_n27027), .Y(new_n27030));
  nor_5  g24682(.A(new_n27030), .B(new_n27025), .Y(n17877));
  nand_5 g24683(.A(new_n17750), .B(new_n17751), .Y(new_n27032));
  xor_4  g24684(.A(new_n27032), .B(new_n17840), .Y(n17889));
  nor_5  g24685(.A(new_n25999), .B(new_n25987), .Y(new_n27034));
  not_8  g24686(.A(new_n25997), .Y(new_n27035));
  nor_5  g24687(.A(new_n27035), .B(new_n25986), .Y(new_n27036));
  nor_5  g24688(.A(new_n27036), .B(new_n27034), .Y(n17912));
  nand_5 g24689(.A(new_n25307), .B(new_n25306), .Y(new_n27038));
  xnor_4 g24690(.A(new_n27038), .B(new_n25309), .Y(n17927));
  nand_5 g24691(.A(new_n25369), .B(new_n25368), .Y(new_n27040));
  xor_4  g24692(.A(new_n27040), .B(new_n25390), .Y(n17931));
  nand_5 g24693(.A(new_n9077), .B(new_n9075), .Y(new_n27042));
  xnor_4 g24694(.A(new_n27042), .B(new_n9079), .Y(n17948));
  nand_5 g24695(.A(new_n18088), .B(new_n18087), .Y(new_n27044));
  xor_4  g24696(.A(new_n27044), .B(new_n18091), .Y(n17956));
  nand_5 g24697(.A(new_n14717), .B(new_n14512), .Y(new_n27046));
  nand_5 g24698(.A(new_n27046), .B(new_n14716), .Y(n17963));
  nand_5 g24699(.A(new_n20154), .B(new_n20139), .Y(new_n27048));
  nand_5 g24700(.A(new_n27048), .B(new_n20138_1), .Y(new_n27049));
  nor_5  g24701(.A(new_n27049), .B(new_n15059), .Y(new_n27050));
  not_8  g24702(.A(new_n27049), .Y(new_n27051_1));
  nor_5  g24703(.A(new_n27051_1), .B(new_n15061), .Y(new_n27052));
  nand_5 g24704(.A(new_n20181), .B(new_n20158), .Y(new_n27053));
  nand_5 g24705(.A(new_n27053), .B(new_n20157), .Y(new_n27054));
  nor_5  g24706(.A(new_n27054), .B(new_n27052), .Y(new_n27055));
  nor_5  g24707(.A(new_n27055), .B(new_n27050), .Y(new_n27056));
  nor_5  g24708(.A(new_n27051_1), .B(new_n15054), .Y(new_n27057));
  nor_5  g24709(.A(new_n27057), .B(new_n27056), .Y(new_n27058));
  nor_5  g24710(.A(new_n27049), .B(new_n15030), .Y(new_n27059));
  nor_5  g24711(.A(new_n27059), .B(new_n27055), .Y(new_n27060));
  nor_5  g24712(.A(new_n27060), .B(new_n27058), .Y(n17976));
  nand_5 g24713(.A(new_n8217), .B(new_n8216), .Y(new_n27062));
  xor_4  g24714(.A(new_n27062), .B(new_n8265), .Y(n17998));
  xor_4  g24715(.A(new_n16740), .B(new_n23659), .Y(n18025));
  nand_5 g24716(.A(new_n23630), .B(new_n23629), .Y(new_n27065));
  xor_4  g24717(.A(new_n27065), .B(new_n23676), .Y(n18043));
  nand_5 g24718(.A(new_n25228), .B(new_n25227), .Y(new_n27067));
  xor_4  g24719(.A(new_n27067), .B(new_n25230), .Y(n18045));
  nand_5 g24720(.A(new_n4256_1), .B(new_n4255), .Y(new_n27069));
  xnor_4 g24721(.A(new_n27069), .B(new_n4268), .Y(n18059));
  or_5   g24722(.A(new_n23289_1), .B(new_n23288), .Y(new_n27071));
  xor_4  g24723(.A(new_n27071), .B(new_n23337), .Y(n18061));
  nand_5 g24724(.A(new_n3606), .B(new_n3605), .Y(new_n27073));
  xnor_4 g24725(.A(new_n27073), .B(new_n3683), .Y(n18071));
  or_5   g24726(.A(new_n11537), .B(new_n11536), .Y(new_n27075));
  xor_4  g24727(.A(new_n27075), .B(new_n11617), .Y(n18143));
  nand_5 g24728(.A(new_n24633), .B(new_n24632), .Y(new_n27077));
  xor_4  g24729(.A(new_n27077), .B(new_n24639), .Y(n18152));
  nand_5 g24730(.A(new_n8732), .B(new_n8731), .Y(new_n27079_1));
  xor_4  g24731(.A(new_n27079_1), .B(new_n8740), .Y(n18193));
  nor_5  g24732(.A(new_n13534), .B(new_n13532), .Y(new_n27081));
  xor_4  g24733(.A(new_n27081), .B(new_n13530), .Y(n18232));
  nand_5 g24734(.A(new_n19458_1), .B(new_n19456), .Y(new_n27083));
  xnor_4 g24735(.A(new_n27083), .B(new_n19492), .Y(n18238));
  nand_5 g24736(.A(new_n21257), .B(new_n21256), .Y(new_n27085));
  xnor_4 g24737(.A(new_n27085), .B(new_n21259), .Y(n18241));
  nand_5 g24738(.A(new_n24080), .B(new_n24081), .Y(new_n27087));
  xor_4  g24739(.A(new_n27087), .B(new_n24090), .Y(n18254));
  nand_5 g24740(.A(new_n24835), .B(new_n24834), .Y(new_n27089_1));
  xor_4  g24741(.A(new_n27089_1), .B(new_n24849), .Y(n18288));
  nand_5 g24742(.A(new_n14052), .B(new_n14050), .Y(new_n27091));
  xor_4  g24743(.A(new_n27091), .B(new_n14090_1), .Y(n18301));
  nand_5 g24744(.A(new_n25205), .B(new_n25204), .Y(new_n27093));
  xnor_4 g24745(.A(new_n27093), .B(new_n25219), .Y(n18304));
  nand_5 g24746(.A(new_n15416), .B(new_n15415), .Y(new_n27095));
  xor_4  g24747(.A(new_n27095), .B(new_n15475), .Y(n18310));
  nand_5 g24748(.A(new_n7588_1), .B(new_n7587), .Y(new_n27097));
  xor_4  g24749(.A(new_n27097), .B(new_n7594), .Y(n18311));
  nand_5 g24750(.A(new_n20299), .B(new_n20300), .Y(new_n27099));
  xor_4  g24751(.A(new_n27099), .B(new_n20314), .Y(n18323));
  nand_5 g24752(.A(new_n6078), .B(new_n6079), .Y(new_n27101));
  xor_4  g24753(.A(new_n27101), .B(new_n6128), .Y(n18332));
  nand_5 g24754(.A(new_n25359), .B(new_n25358), .Y(new_n27103));
  xor_4  g24755(.A(new_n27103), .B(new_n25400), .Y(n18343));
  nand_5 g24756(.A(new_n22193), .B(new_n22192), .Y(new_n27105));
  xor_4  g24757(.A(new_n27105), .B(new_n22195), .Y(n18350));
  nand_5 g24758(.A(new_n20805), .B(new_n20804), .Y(new_n27107));
  xor_4  g24759(.A(new_n27107), .B(new_n20815), .Y(n18362));
  nand_5 g24760(.A(new_n5587), .B(new_n5586), .Y(new_n27109));
  xor_4  g24761(.A(new_n27109), .B(new_n5657), .Y(n18377));
  nand_5 g24762(.A(new_n4455), .B(new_n4456), .Y(new_n27111));
  xnor_4 g24763(.A(new_n27111), .B(new_n4483), .Y(n18405));
  nand_5 g24764(.A(new_n19285), .B(new_n19286), .Y(new_n27113));
  xor_4  g24765(.A(new_n27113), .B(new_n19296), .Y(n18414));
  nand_5 g24766(.A(new_n16797), .B(new_n16795), .Y(new_n27115));
  xor_4  g24767(.A(new_n27115), .B(new_n16807), .Y(n18418));
  nand_5 g24768(.A(new_n9368), .B(new_n9367), .Y(new_n27117));
  xnor_4 g24769(.A(new_n27117), .B(new_n9417), .Y(n18437));
  nor_5  g24770(.A(new_n23074), .B(new_n23073), .Y(new_n27119));
  xor_4  g24771(.A(new_n27119), .B(new_n23122), .Y(n18439));
  nand_5 g24772(.A(new_n12933), .B(new_n12932), .Y(new_n27121));
  xor_4  g24773(.A(new_n27121), .B(new_n12936), .Y(n18445));
  nand_5 g24774(.A(new_n7899), .B(new_n7898), .Y(new_n27123));
  xnor_4 g24775(.A(new_n27123), .B(new_n7948), .Y(n18467));
  nand_5 g24776(.A(new_n21210), .B(new_n21209), .Y(new_n27125));
  xnor_4 g24777(.A(new_n27125), .B(new_n21275), .Y(n18482));
  nand_5 g24778(.A(new_n21583), .B(new_n21584), .Y(new_n27127));
  xor_4  g24779(.A(new_n27127), .B(new_n21607), .Y(n18509));
  nor_5  g24780(.A(new_n16034), .B(new_n16033), .Y(new_n27129));
  xor_4  g24781(.A(new_n27129), .B(new_n10431), .Y(n18513));
  nand_5 g24782(.A(new_n17381), .B(new_n17383), .Y(new_n27131));
  xor_4  g24783(.A(new_n27131), .B(new_n17405), .Y(n18515));
  nand_5 g24784(.A(new_n18392), .B(new_n18390), .Y(new_n27133));
  xnor_4 g24785(.A(new_n27133), .B(new_n18415), .Y(n18572));
  xor_4  g24786(.A(new_n26789), .B(new_n26774), .Y(new_n27135));
  and_5  g24787(.A(new_n26790), .B(new_n27135), .Y(n18574));
  nand_5 g24788(.A(new_n24250), .B(new_n24249), .Y(new_n27137));
  xor_4  g24789(.A(new_n27137), .B(new_n24252), .Y(n18576));
  nand_5 g24790(.A(new_n25757), .B(new_n25756_1), .Y(new_n27139));
  xnor_4 g24791(.A(new_n27139), .B(new_n25768), .Y(n18582));
  nand_5 g24792(.A(new_n22837), .B(new_n22836), .Y(new_n27141));
  xnor_4 g24793(.A(new_n27141), .B(new_n22852), .Y(n18583));
  nand_5 g24794(.A(new_n23320), .B(new_n23322), .Y(new_n27143));
  xnor_4 g24795(.A(new_n27143), .B(new_n23321), .Y(n18610));
  xor_4  g24796(.A(new_n25241), .B(new_n25239), .Y(n18635));
  nand_5 g24797(.A(new_n7686_1), .B(new_n7687), .Y(new_n27146));
  xnor_4 g24798(.A(new_n27146), .B(new_n7704), .Y(n18653));
  nand_5 g24799(.A(new_n3992), .B(new_n3991), .Y(new_n27148));
  xnor_4 g24800(.A(new_n27148), .B(new_n4060), .Y(n18679));
  nand_5 g24801(.A(new_n23457), .B(new_n23448), .Y(new_n27150));
  xor_4  g24802(.A(new_n27150), .B(new_n23456), .Y(n18693));
  nand_5 g24803(.A(new_n3222), .B(new_n3221), .Y(new_n27152));
  xnor_4 g24804(.A(new_n27152), .B(new_n3266), .Y(n18708));
  nand_5 g24805(.A(new_n26172), .B(new_n26171), .Y(new_n27154));
  xnor_4 g24806(.A(new_n27154), .B(new_n26174), .Y(n18721));
  nand_5 g24807(.A(new_n21406), .B(new_n21405), .Y(new_n27156));
  xor_4  g24808(.A(new_n27156), .B(new_n21450), .Y(n18725));
  nand_5 g24809(.A(new_n23832), .B(new_n23833), .Y(new_n27158_1));
  xnor_4 g24810(.A(new_n27158_1), .B(new_n23854), .Y(n18751));
  nand_5 g24811(.A(new_n19032), .B(new_n19033_1), .Y(new_n27160));
  xor_4  g24812(.A(new_n27160), .B(new_n19053), .Y(n18780));
  nand_5 g24813(.A(new_n22402), .B(new_n22401), .Y(new_n27162));
  xor_4  g24814(.A(new_n27162), .B(new_n22457), .Y(n18782));
  nor_5  g24815(.A(new_n8758), .B(new_n8688), .Y(new_n27164));
  nor_5  g24816(.A(new_n8757), .B(new_n8685), .Y(new_n27165));
  nor_5  g24817(.A(new_n27165), .B(new_n27164), .Y(n18802));
  nand_5 g24818(.A(new_n12607_1), .B(new_n12606), .Y(new_n27167));
  xor_4  g24819(.A(new_n27167), .B(new_n12619), .Y(n18830));
  nand_5 g24820(.A(new_n14805), .B(new_n14806), .Y(new_n27169));
  xor_4  g24821(.A(new_n27169), .B(new_n14811), .Y(n18831));
  nand_5 g24822(.A(new_n13828), .B(new_n13827), .Y(new_n27171));
  xor_4  g24823(.A(new_n27171), .B(new_n13837), .Y(n18843));
  nand_5 g24824(.A(new_n3236), .B(new_n3235_1), .Y(new_n27173));
  xnor_4 g24825(.A(new_n27173), .B(new_n3262), .Y(n18858));
  nand_5 g24826(.A(new_n11581), .B(new_n11580_1), .Y(new_n27175));
  xor_4  g24827(.A(new_n27175), .B(new_n11605), .Y(n18859));
  nand_5 g24828(.A(new_n19845), .B(new_n19844), .Y(new_n27177));
  xor_4  g24829(.A(new_n27177), .B(new_n19899), .Y(n18864));
  nand_5 g24830(.A(new_n5050), .B(new_n5048), .Y(new_n27179));
  xnor_4 g24831(.A(new_n27179), .B(new_n5131_1), .Y(n18865));
  nand_5 g24832(.A(new_n24542), .B(new_n24540), .Y(new_n27181));
  xnor_4 g24833(.A(new_n27181), .B(new_n24550), .Y(n18886));
  nand_5 g24834(.A(new_n19040), .B(new_n19041), .Y(new_n27183));
  xor_4  g24835(.A(new_n27183), .B(new_n19049), .Y(n18887));
  nor_5  g24836(.A(new_n10191), .B(new_n10190), .Y(new_n27185));
  xor_4  g24837(.A(new_n27185), .B(new_n10244_1), .Y(n18919));
  nor_5  g24838(.A(new_n14296), .B(new_n14295), .Y(new_n27187));
  xor_4  g24839(.A(new_n27187), .B(new_n14310_1), .Y(n18940));
  nand_5 g24840(.A(new_n26307), .B(new_n26306), .Y(new_n27189));
  xnor_4 g24841(.A(new_n27189), .B(new_n26309), .Y(n18945));
  nand_5 g24842(.A(new_n25950), .B(new_n25949), .Y(new_n27191));
  xor_4  g24843(.A(new_n27191), .B(new_n25960), .Y(n18970));
  nand_5 g24844(.A(new_n19558), .B(new_n19557), .Y(new_n27193));
  xor_4  g24845(.A(new_n27193), .B(new_n19560), .Y(n18977));
  nand_5 g24846(.A(new_n17524_1), .B(new_n17525), .Y(new_n27195));
  xor_4  g24847(.A(new_n27195), .B(new_n17534), .Y(n18982));
  nand_5 g24848(.A(new_n23910), .B(new_n23909), .Y(new_n27197));
  xnor_4 g24849(.A(new_n27197), .B(new_n23939), .Y(n18999));
  nand_5 g24850(.A(new_n6438), .B(new_n6439), .Y(new_n27199));
  xor_4  g24851(.A(new_n27199), .B(new_n6512), .Y(n19044));
  nand_5 g24852(.A(new_n17177), .B(new_n17179), .Y(new_n27201));
  xnor_4 g24853(.A(new_n27201), .B(new_n17188), .Y(n19125));
  nand_5 g24854(.A(new_n6445), .B(new_n6444), .Y(new_n27203));
  xnor_4 g24855(.A(new_n27203), .B(new_n6509), .Y(n19141));
  nand_5 g24856(.A(new_n20022), .B(new_n16179), .Y(new_n27205));
  not_8  g24857(.A(new_n16179), .Y(new_n27206));
  nand_5 g24858(.A(new_n20023), .B(new_n27206), .Y(new_n27207));
  nand_5 g24859(.A(new_n27207), .B(new_n27205), .Y(new_n27208));
  nand_5 g24860(.A(new_n20027), .B(new_n16185_1), .Y(new_n27209));
  not_8  g24861(.A(new_n27209), .Y(new_n27210));
  nor_5  g24862(.A(new_n20027), .B(new_n16185_1), .Y(new_n27211));
  not_8  g24863(.A(new_n21477), .Y(new_n27212));
  nor_5  g24864(.A(new_n21480), .B(new_n27212), .Y(new_n27213));
  nor_5  g24865(.A(new_n27213), .B(new_n21479), .Y(new_n27214));
  nor_5  g24866(.A(new_n27214), .B(new_n27211), .Y(new_n27215));
  nor_5  g24867(.A(new_n27215), .B(new_n27210), .Y(new_n27216));
  xor_4  g24868(.A(new_n27216), .B(new_n27208), .Y(n19164));
  nand_5 g24869(.A(new_n9586), .B(new_n9585), .Y(new_n27218));
  xor_4  g24870(.A(new_n27218), .B(new_n9621), .Y(n19174));
  nand_5 g24871(.A(new_n24148), .B(new_n24149), .Y(new_n27220));
  xor_4  g24872(.A(new_n27220), .B(new_n24151), .Y(n19176));
  nand_5 g24873(.A(new_n25201), .B(new_n25200_1), .Y(new_n27222));
  xnor_4 g24874(.A(new_n27222), .B(new_n25221), .Y(n19202));
  nand_5 g24875(.A(new_n23214), .B(new_n23213), .Y(new_n27224));
  xnor_4 g24876(.A(new_n27224), .B(new_n23225), .Y(n19220));
  nand_5 g24877(.A(new_n9027), .B(new_n9026), .Y(new_n27226));
  xor_4  g24878(.A(new_n27226), .B(new_n9098), .Y(n19221));
  nand_5 g24879(.A(new_n13098), .B(new_n13099), .Y(new_n27228));
  xnor_4 g24880(.A(new_n27228), .B(new_n13108), .Y(n19223));
  nand_5 g24881(.A(new_n19883), .B(new_n19884), .Y(new_n27230));
  xor_4  g24882(.A(new_n27230), .B(new_n19885), .Y(n19224));
  nand_5 g24883(.A(new_n18021), .B(new_n18011), .Y(new_n27232));
  xnor_4 g24884(.A(new_n27232), .B(new_n18019), .Y(n19233));
  nand_5 g24885(.A(new_n14759), .B(new_n14758), .Y(new_n27234));
  xor_4  g24886(.A(new_n27234), .B(new_n14794), .Y(n19244));
  nor_5  g24887(.A(new_n10184), .B(new_n10183), .Y(new_n27236));
  xor_4  g24888(.A(new_n27236), .B(new_n10246), .Y(n19314));
  nand_5 g24889(.A(new_n12493), .B(new_n12492), .Y(new_n27238));
  xor_4  g24890(.A(new_n27238), .B(new_n12511), .Y(n19315));
  nand_5 g24891(.A(new_n15433), .B(new_n15434), .Y(new_n27240));
  xnor_4 g24892(.A(new_n27240), .B(new_n15466), .Y(n19323));
  nand_5 g24893(.A(new_n25019), .B(new_n25020), .Y(new_n27242));
  xnor_4 g24894(.A(new_n27242), .B(new_n25022), .Y(n19333));
  not_8  g24895(.A(new_n20014), .Y(new_n27244));
  nand_5 g24896(.A(new_n27244), .B(new_n11521), .Y(new_n27245));
  nand_5 g24897(.A(new_n20014), .B(new_n11522), .Y(new_n27246));
  nand_5 g24898(.A(new_n20041), .B(new_n20018), .Y(new_n27247));
  nand_5 g24899(.A(new_n27247), .B(new_n20019), .Y(new_n27248));
  nand_5 g24900(.A(new_n27248), .B(new_n27246), .Y(new_n27249));
  nand_5 g24901(.A(new_n27249), .B(new_n27245), .Y(n19348));
  not_8  g24902(.A(new_n19416), .Y(new_n27251));
  nor_5  g24903(.A(new_n27251), .B(new_n19415), .Y(new_n27252));
  xor_4  g24904(.A(new_n27252), .B(new_n19504), .Y(n19354));
  nand_5 g24905(.A(new_n12843_1), .B(new_n12842), .Y(new_n27254));
  xor_4  g24906(.A(new_n27254), .B(new_n12881), .Y(n19367));
  nand_5 g24907(.A(new_n21985), .B(new_n21984), .Y(new_n27256));
  xor_4  g24908(.A(new_n27256), .B(new_n22012), .Y(n19385));
  nand_5 g24909(.A(new_n19634), .B(new_n19623_1), .Y(new_n27258));
  xor_4  g24910(.A(new_n27258), .B(new_n19631), .Y(new_n27259));
  xor_4  g24911(.A(new_n27259), .B(new_n19673), .Y(n19389));
  nand_5 g24912(.A(new_n18885), .B(new_n18884), .Y(new_n27261));
  xnor_4 g24913(.A(new_n27261), .B(new_n18917), .Y(n19401));
  or_5   g24914(.A(new_n25508), .B(new_n25499_1), .Y(new_n27263));
  xor_4  g24915(.A(new_n27263), .B(new_n25506), .Y(n19414));
  nand_5 g24916(.A(new_n22219), .B(new_n22218), .Y(new_n27265));
  xor_4  g24917(.A(new_n27265), .B(new_n20614), .Y(n19424));
  nand_5 g24918(.A(new_n24556), .B(new_n24533), .Y(new_n27267));
  xnor_4 g24919(.A(new_n27267), .B(new_n24554), .Y(n19450));
  nand_5 g24920(.A(new_n27244), .B(new_n16169), .Y(new_n27269));
  nand_5 g24921(.A(new_n20014), .B(new_n16109), .Y(new_n27270));
  nand_5 g24922(.A(new_n20017_1), .B(new_n16171), .Y(new_n27271));
  nand_5 g24923(.A(new_n20016), .B(new_n16172), .Y(new_n27272));
  not_8  g24924(.A(new_n27205), .Y(new_n27273));
  not_8  g24925(.A(new_n27207), .Y(new_n27274));
  nor_5  g24926(.A(new_n27216), .B(new_n27274), .Y(new_n27275));
  nor_5  g24927(.A(new_n27275), .B(new_n27273), .Y(new_n27276));
  not_8  g24928(.A(new_n27276), .Y(new_n27277));
  nand_5 g24929(.A(new_n27277), .B(new_n27272), .Y(new_n27278));
  and_5  g24930(.A(new_n27278), .B(new_n27271), .Y(new_n27279));
  nand_5 g24931(.A(new_n27279), .B(new_n27270), .Y(new_n27280));
  nand_5 g24932(.A(new_n27280), .B(new_n27269), .Y(n19458));
  nand_5 g24933(.A(new_n17615), .B(new_n17617), .Y(new_n27282));
  xor_4  g24934(.A(new_n27282), .B(new_n17626), .Y(n19467));
  nand_5 g24935(.A(new_n9362), .B(new_n9361), .Y(new_n27284));
  xnor_4 g24936(.A(new_n27284), .B(new_n9419_1), .Y(n19496));
  nand_5 g24937(.A(new_n17580), .B(new_n17579), .Y(new_n27286));
  xor_4  g24938(.A(new_n27286), .B(new_n17588), .Y(n19523));
  nand_5 g24939(.A(new_n5077_1), .B(new_n5076), .Y(new_n27288));
  xnor_4 g24940(.A(new_n27288), .B(new_n5123), .Y(n19570));
  not_8  g24941(.A(new_n13949), .Y(new_n27290));
  nand_5 g24942(.A(new_n27290), .B(new_n13948), .Y(new_n27291));
  xor_4  g24943(.A(new_n27291), .B(new_n13961), .Y(n19602));
  nand_5 g24944(.A(new_n14349), .B(new_n14348), .Y(new_n27293));
  xor_4  g24945(.A(new_n27293), .B(new_n14354), .Y(n19617));
  nand_5 g24946(.A(new_n15768), .B(new_n15767), .Y(new_n27295));
  xor_4  g24947(.A(new_n27295), .B(new_n15806), .Y(n19623));
  xor_4  g24948(.A(new_n25552), .B(new_n25550_1), .Y(n19641));
  nand_5 g24949(.A(new_n25287), .B(new_n25286), .Y(new_n27298));
  xnor_4 g24950(.A(new_n27298), .B(new_n25319), .Y(n19648));
  nand_5 g24951(.A(new_n18397), .B(new_n18395), .Y(new_n27300));
  xnor_4 g24952(.A(new_n27300), .B(new_n18413), .Y(n19664));
  nand_5 g24953(.A(new_n22907_1), .B(new_n22906), .Y(new_n27302));
  xnor_4 g24954(.A(new_n27302), .B(new_n22921), .Y(n19736));
  nor_5  g24955(.A(new_n25496), .B(new_n3440), .Y(new_n27304));
  nor_5  g24956(.A(new_n25507), .B(new_n27304), .Y(new_n27305));
  nor_5  g24957(.A(new_n25509), .B(new_n25496), .Y(new_n27306));
  nor_5  g24958(.A(new_n27306), .B(new_n27305), .Y(n19749));
  nand_5 g24959(.A(new_n17257), .B(new_n17256), .Y(new_n27308));
  xnor_4 g24960(.A(new_n27308), .B(new_n17271), .Y(n19756));
  or_5   g24961(.A(new_n13956), .B(new_n13955), .Y(new_n27310));
  xor_4  g24962(.A(new_n27310), .B(new_n13959), .Y(n19767));
  nand_5 g24963(.A(new_n3598), .B(new_n3599), .Y(new_n27312));
  xnor_4 g24964(.A(new_n27312), .B(new_n3685), .Y(n19780));
  nand_5 g24965(.A(new_n26189), .B(new_n26188), .Y(new_n27314));
  xnor_4 g24966(.A(new_n27314), .B(new_n26191_1), .Y(n19792));
  nand_5 g24967(.A(new_n23650), .B(new_n23649), .Y(new_n27316));
  xor_4  g24968(.A(new_n27316), .B(new_n23666), .Y(n19798));
  nand_5 g24969(.A(new_n19181), .B(new_n19180), .Y(new_n27318));
  xor_4  g24970(.A(new_n27318), .B(new_n19183), .Y(n19873));
  nor_5  g24971(.A(new_n21292), .B(new_n21294), .Y(new_n27320));
  nor_5  g24972(.A(new_n21304), .B(new_n27320), .Y(new_n27321));
  xor_4  g24973(.A(new_n27321), .B(new_n21294), .Y(n19909));
  nand_5 g24974(.A(new_n22911), .B(new_n22910_1), .Y(new_n27323));
  xnor_4 g24975(.A(new_n27323), .B(new_n22919), .Y(n19916));
  nand_5 g24976(.A(new_n23642), .B(new_n23641), .Y(new_n27325));
  xor_4  g24977(.A(new_n27325), .B(new_n23670), .Y(n19923));
  nand_5 g24978(.A(new_n21821), .B(new_n21820_1), .Y(new_n27327));
  xnor_4 g24979(.A(new_n27327), .B(new_n21861), .Y(n19930));
  nor_5  g24980(.A(new_n7301), .B(new_n7299), .Y(new_n27329));
  or_5   g24981(.A(new_n27329), .B(n588), .Y(n19968));
  nand_5 g24982(.A(new_n22425), .B(new_n22426), .Y(new_n27331));
  xnor_4 g24983(.A(new_n27331), .B(new_n22444_1), .Y(n19988));
  not_8  g24984(.A(new_n23749), .Y(new_n27333));
  nand_5 g24985(.A(new_n27333), .B(new_n23746), .Y(new_n27334));
  nand_5 g24986(.A(new_n27334), .B(new_n23745), .Y(new_n27335));
  nand_5 g24987(.A(new_n24580), .B(new_n23743), .Y(new_n27336));
  nand_5 g24988(.A(new_n27336), .B(new_n27335), .Y(new_n27337));
  nand_5 g24989(.A(new_n24581), .B(new_n23744), .Y(new_n27338));
  nand_5 g24990(.A(new_n27338), .B(new_n27334), .Y(new_n27339));
  and_5  g24991(.A(new_n27339), .B(new_n27337), .Y(n20004));
  nand_5 g24992(.A(new_n23836), .B(new_n23837), .Y(new_n27341));
  xnor_4 g24993(.A(new_n27341), .B(new_n23850), .Y(n20017));
  nand_5 g24994(.A(new_n21224), .B(new_n21223), .Y(new_n27343));
  xnor_4 g24995(.A(new_n27343), .B(new_n21271), .Y(n20033));
  nand_5 g24996(.A(new_n15989), .B(new_n15988), .Y(new_n27345));
  xnor_4 g24997(.A(new_n27345), .B(new_n16005), .Y(n20061));
  nand_5 g24998(.A(new_n20759), .B(new_n20758), .Y(new_n27347));
  xor_4  g24999(.A(new_n27347), .B(new_n20762), .Y(n20069));
  nand_5 g25000(.A(new_n16766), .B(new_n16685), .Y(new_n27349));
  nand_5 g25001(.A(new_n27349), .B(new_n16684_1), .Y(n20086));
  nand_5 g25002(.A(new_n22313), .B(new_n22315), .Y(new_n27351));
  xor_4  g25003(.A(new_n27351), .B(new_n22317_1), .Y(n20096));
  nand_5 g25004(.A(new_n15450), .B(new_n15449), .Y(new_n27353));
  xnor_4 g25005(.A(new_n27353), .B(new_n15458), .Y(n20103));
  nand_5 g25006(.A(new_n13438), .B(new_n13437), .Y(new_n27355));
  xor_4  g25007(.A(new_n27355), .B(new_n13483), .Y(n20126));
  or_5   g25008(.A(new_n24291), .B(new_n24290), .Y(new_n27357));
  xor_4  g25009(.A(new_n27357), .B(new_n24329), .Y(n20149));
  nand_5 g25010(.A(new_n13804), .B(new_n13803), .Y(new_n27359));
  xor_4  g25011(.A(new_n27359), .B(new_n13849), .Y(n20187));
  nand_5 g25012(.A(new_n20080), .B(new_n20079), .Y(new_n27361));
  xor_4  g25013(.A(new_n27361), .B(new_n20111), .Y(n20279));
  not_8  g25014(.A(new_n25773_1), .Y(new_n27363));
  nand_5 g25015(.A(new_n27363), .B(new_n25748), .Y(new_n27364));
  nand_5 g25016(.A(new_n25773_1), .B(new_n25747), .Y(new_n27365));
  nand_5 g25017(.A(new_n27365), .B(new_n27364), .Y(n20287));
  nand_5 g25018(.A(new_n23494), .B(new_n23495), .Y(new_n27367));
  xor_4  g25019(.A(new_n27367), .B(new_n23497), .Y(n20301));
  nor_5  g25020(.A(new_n9426), .B(new_n9427), .Y(new_n27369));
  nor_5  g25021(.A(new_n27369), .B(new_n9224), .Y(n20330));
  nand_5 g25022(.A(new_n13812), .B(new_n13811), .Y(new_n27371));
  xor_4  g25023(.A(new_n27371), .B(new_n13845), .Y(n20333));
  not_8  g25024(.A(new_n12107), .Y(new_n27373));
  nor_5  g25025(.A(new_n27373), .B(new_n11974), .Y(new_n27374));
  nand_5 g25026(.A(new_n27373), .B(new_n12020), .Y(new_n27375));
  nand_5 g25027(.A(new_n27375), .B(new_n12023), .Y(new_n27376));
  nor_5  g25028(.A(new_n27376), .B(new_n27374), .Y(n20355));
  xor_4  g25029(.A(new_n9650), .B(new_n5839), .Y(n20366));
  nand_5 g25030(.A(new_n22057), .B(new_n22051), .Y(new_n27379));
  xnor_4 g25031(.A(new_n27379), .B(new_n22053), .Y(n20388));
  nand_5 g25032(.A(new_n25371), .B(new_n25370_1), .Y(new_n27381));
  xor_4  g25033(.A(new_n27381), .B(new_n25388), .Y(n20402));
  nand_5 g25034(.A(new_n17793), .B(new_n17792), .Y(new_n27383));
  xor_4  g25035(.A(new_n27383), .B(new_n17828), .Y(n20403));
  xor_4  g25036(.A(new_n3250), .B(new_n3247), .Y(n20424));
  nor_5  g25037(.A(new_n23313), .B(new_n23311), .Y(new_n27386));
  xor_4  g25038(.A(new_n27386), .B(new_n23326), .Y(n20436));
  nor_5  g25039(.A(new_n9405), .B(new_n9404), .Y(new_n27388));
  xor_4  g25040(.A(new_n27388), .B(new_n2627), .Y(n20441));
  or_5   g25041(.A(new_n8694_1), .B(new_n8692), .Y(new_n27390));
  xor_4  g25042(.A(new_n27390), .B(new_n8756), .Y(n20445));
  nand_5 g25043(.A(new_n5580), .B(new_n5579_1), .Y(new_n27392));
  xor_4  g25044(.A(new_n27392), .B(new_n5659), .Y(n20450));
  nand_5 g25045(.A(new_n19087), .B(new_n19083), .Y(new_n27394));
  nand_5 g25046(.A(new_n27394), .B(new_n19089), .Y(n20490));
  nand_5 g25047(.A(new_n23221), .B(new_n23220), .Y(new_n27396));
  xnor_4 g25048(.A(new_n27396), .B(new_n23223), .Y(n20495));
  not_8  g25049(.A(new_n17845), .Y(new_n27398));
  xor_4  g25050(.A(new_n17842), .B(new_n17844), .Y(new_n27399));
  nor_5  g25051(.A(new_n27399), .B(new_n27398), .Y(n20515));
  nor_5  g25052(.A(new_n26193), .B(new_n26194), .Y(new_n27401));
  nor_5  g25053(.A(new_n27401), .B(new_n26185), .Y(n20533));
  nand_5 g25054(.A(new_n20609_1), .B(new_n20610), .Y(new_n27403));
  xnor_4 g25055(.A(new_n27403), .B(new_n20617), .Y(n20582));
  nand_5 g25056(.A(new_n22578), .B(new_n22577), .Y(new_n27405));
  xor_4  g25057(.A(new_n27405), .B(new_n22613), .Y(n20590));
  nand_5 g25058(.A(new_n3665_1), .B(new_n3662), .Y(new_n27407));
  xnor_4 g25059(.A(new_n27407), .B(new_n3667), .Y(n20602));
  nand_5 g25060(.A(new_n19045), .B(new_n19044_1), .Y(new_n27409));
  xor_4  g25061(.A(new_n27409), .B(new_n19047), .Y(n20609));
  nand_5 g25062(.A(new_n7447), .B(new_n7448), .Y(new_n27411));
  xor_4  g25063(.A(new_n27411), .B(new_n7457), .Y(n20623));
  nand_5 g25064(.A(new_n23622), .B(new_n23621), .Y(new_n27413));
  xor_4  g25065(.A(new_n27413), .B(new_n23680), .Y(n20629));
  nand_5 g25066(.A(new_n15993), .B(new_n15992), .Y(new_n27415));
  xnor_4 g25067(.A(new_n27415), .B(new_n16003), .Y(n20661));
  nand_5 g25068(.A(new_n9711), .B(new_n9709), .Y(new_n27417));
  xor_4  g25069(.A(new_n27417), .B(new_n9718), .Y(n20673));
  nand_5 g25070(.A(new_n23634), .B(new_n23633), .Y(new_n27419));
  xor_4  g25071(.A(new_n27419), .B(new_n23674), .Y(n20678));
  nand_5 g25072(.A(new_n17277), .B(new_n17244), .Y(new_n27421));
  nand_5 g25073(.A(new_n27421), .B(new_n17243_1), .Y(new_n27422));
  nor_5  g25074(.A(new_n27422), .B(new_n17237), .Y(n20680));
  nand_5 g25075(.A(new_n7277_1), .B(new_n4577), .Y(new_n27424));
  nand_5 g25076(.A(new_n27424), .B(new_n7278), .Y(n20685));
  nor_5  g25077(.A(new_n27059), .B(new_n27057), .Y(new_n27426));
  xor_4  g25078(.A(new_n27426), .B(new_n27056), .Y(n20691));
  nand_5 g25079(.A(new_n18401), .B(new_n18400), .Y(new_n27428));
  xnor_4 g25080(.A(new_n27428), .B(new_n18411), .Y(n20696));
  nand_5 g25081(.A(new_n25918), .B(new_n25917), .Y(new_n27430));
  xnor_4 g25082(.A(new_n27430), .B(new_n25927), .Y(n20704));
  nand_5 g25083(.A(new_n24840_1), .B(new_n24841_1), .Y(new_n27432));
  xnor_4 g25084(.A(new_n27432), .B(new_n24843), .Y(n20705));
  nand_5 g25085(.A(new_n11543), .B(new_n11544), .Y(new_n27434));
  xor_4  g25086(.A(new_n27434), .B(new_n11615_1), .Y(n20709));
  nand_5 g25087(.A(new_n17066), .B(new_n17065), .Y(new_n27436));
  xnor_4 g25088(.A(new_n27436), .B(new_n17100), .Y(n20713));
  nand_5 g25089(.A(new_n9904), .B(new_n9903), .Y(new_n27438));
  xor_4  g25090(.A(new_n27438), .B(new_n9907), .Y(n20722));
  not_8  g25091(.A(new_n22507), .Y(new_n27440));
  not_8  g25092(.A(new_n22510), .Y(new_n27441));
  nor_5  g25093(.A(new_n22523), .B(new_n27441), .Y(new_n27442));
  nor_5  g25094(.A(new_n27442), .B(new_n27440), .Y(new_n27443));
  nor_5  g25095(.A(new_n26542), .B(new_n22506), .Y(new_n27444));
  nor_5  g25096(.A(new_n27444), .B(new_n27443), .Y(new_n27445));
  nor_5  g25097(.A(new_n26543), .B(new_n22509), .Y(new_n27446));
  nor_5  g25098(.A(new_n27446), .B(new_n27442), .Y(new_n27447));
  nor_5  g25099(.A(new_n27447), .B(new_n27445), .Y(n20723));
  nand_5 g25100(.A(new_n25750), .B(new_n25752), .Y(new_n27449));
  xnor_4 g25101(.A(new_n27449), .B(new_n25770), .Y(n20748));
  nand_5 g25102(.A(new_n6106), .B(new_n6105_1), .Y(new_n27451));
  xor_4  g25103(.A(new_n27451), .B(new_n6120), .Y(n20761));
  or_5   g25104(.A(new_n23295), .B(new_n23294), .Y(new_n27453));
  xor_4  g25105(.A(new_n27453), .B(new_n23335), .Y(n20774));
  nand_5 g25106(.A(new_n27270), .B(new_n27269), .Y(new_n27455));
  xor_4  g25107(.A(new_n27455), .B(new_n27279), .Y(n20788));
  nor_5  g25108(.A(new_n26493), .B(new_n26490), .Y(new_n27457));
  nor_5  g25109(.A(new_n26492_1), .B(new_n26489), .Y(new_n27458));
  nor_5  g25110(.A(new_n27458), .B(new_n27457), .Y(n20795));
  nor_5  g25111(.A(new_n23370), .B(new_n23367), .Y(new_n27460));
  or_5   g25112(.A(new_n27460), .B(new_n23371_1), .Y(new_n27461));
  nand_5 g25113(.A(new_n23376), .B(new_n23358), .Y(new_n27462));
  nand_5 g25114(.A(new_n27462), .B(new_n25350), .Y(new_n27463));
  xor_4  g25115(.A(new_n27463), .B(new_n27461), .Y(n20803));
  or_5   g25116(.A(new_n27025), .B(new_n27027), .Y(new_n27465));
  xor_4  g25117(.A(new_n27465), .B(new_n27029), .Y(n20869));
  nand_5 g25118(.A(new_n26113_1), .B(new_n26112), .Y(new_n27467));
  xnor_4 g25119(.A(new_n27467), .B(new_n26121), .Y(n20879));
  nand_5 g25120(.A(new_n7248), .B(new_n7246), .Y(new_n27469));
  xnor_4 g25121(.A(new_n27469), .B(new_n7286), .Y(n20915));
  nand_5 g25122(.A(new_n8335), .B(n2160), .Y(new_n27471));
  nand_5 g25123(.A(n19282), .B(new_n13565), .Y(new_n27472));
  nand_5 g25124(.A(new_n24863), .B(new_n24860), .Y(new_n27473));
  nand_5 g25125(.A(new_n27473), .B(new_n24862), .Y(new_n27474));
  nand_5 g25126(.A(new_n27474), .B(new_n27472), .Y(new_n27475));
  nand_5 g25127(.A(new_n27475), .B(new_n27471), .Y(new_n27476));
  nand_5 g25128(.A(new_n27476), .B(new_n25991), .Y(new_n27477));
  nand_5 g25129(.A(new_n27472), .B(new_n27471), .Y(new_n27478));
  xor_4  g25130(.A(new_n27478), .B(new_n27474), .Y(new_n27479));
  nand_5 g25131(.A(new_n27479), .B(new_n24695), .Y(new_n27480));
  or_5   g25132(.A(new_n27479), .B(new_n24695), .Y(new_n27481));
  nand_5 g25133(.A(new_n24867), .B(new_n24858), .Y(new_n27482));
  nand_5 g25134(.A(new_n27482), .B(new_n24866), .Y(new_n27483));
  nand_5 g25135(.A(new_n27483), .B(new_n27481), .Y(new_n27484));
  nand_5 g25136(.A(new_n27484), .B(new_n27480), .Y(new_n27485));
  not_8  g25137(.A(new_n27485), .Y(new_n27486));
  nand_5 g25138(.A(new_n27486), .B(new_n27477), .Y(new_n27487));
  not_8  g25139(.A(new_n27476), .Y(new_n27488));
  nand_5 g25140(.A(new_n27488), .B(new_n25990), .Y(new_n27489));
  nand_5 g25141(.A(new_n27489), .B(new_n27485), .Y(new_n27490));
  nand_5 g25142(.A(new_n27490), .B(new_n27487), .Y(new_n27491));
  xor_4  g25143(.A(new_n27488), .B(new_n25982), .Y(new_n27492));
  nor_5  g25144(.A(new_n27492), .B(new_n27491), .Y(n20935));
  nand_5 g25145(.A(new_n25299), .B(new_n25298), .Y(new_n27494));
  xnor_4 g25146(.A(new_n27494), .B(new_n25313), .Y(n20936));
  nand_5 g25147(.A(new_n19536), .B(new_n19537), .Y(new_n27496));
  xnor_4 g25148(.A(new_n27496), .B(new_n19538), .Y(n21008));
  nand_5 g25149(.A(new_n22405), .B(new_n22406), .Y(new_n27498));
  xnor_4 g25150(.A(new_n27498), .B(new_n22454), .Y(n21017));
  nand_5 g25151(.A(new_n26632), .B(new_n24618_1), .Y(new_n27500));
  nor_5  g25152(.A(new_n26632), .B(new_n24618_1), .Y(new_n27501));
  or_5   g25153(.A(new_n26635), .B(new_n27501), .Y(new_n27502));
  nand_5 g25154(.A(new_n27502), .B(new_n27500), .Y(new_n27503));
  nor_5  g25155(.A(new_n27503), .B(new_n26631), .Y(n21034));
  nand_5 g25156(.A(new_n25473), .B(new_n25472), .Y(new_n27505));
  xnor_4 g25157(.A(new_n27505), .B(new_n25475_1), .Y(n21046));
  nand_5 g25158(.A(new_n9795), .B(new_n9796), .Y(new_n27507));
  xnor_4 g25159(.A(new_n27507), .B(new_n9818), .Y(n21062));
  not_8  g25160(.A(new_n26292), .Y(new_n27509));
  nand_5 g25161(.A(new_n26287_1), .B(new_n26288), .Y(new_n27510));
  nand_5 g25162(.A(new_n27510), .B(new_n27509), .Y(new_n27511));
  xor_4  g25163(.A(new_n27511), .B(new_n26185), .Y(n21093));
  nand_5 g25164(.A(new_n11274), .B(new_n11273_1), .Y(new_n27513));
  xnor_4 g25165(.A(new_n27513), .B(new_n9079), .Y(n21094));
  nand_5 g25166(.A(new_n16966), .B(new_n16965), .Y(new_n27515));
  xor_4  g25167(.A(new_n27515), .B(new_n16993), .Y(n21123));
  nor_5  g25168(.A(new_n21722), .B(new_n21721), .Y(new_n27517));
  xor_4  g25169(.A(new_n27517), .B(new_n21631), .Y(n21154));
  nand_5 g25170(.A(new_n17947), .B(new_n17946), .Y(new_n27519));
  xnor_4 g25171(.A(new_n27519), .B(new_n17976_1), .Y(n21157));
  nor_5  g25172(.A(new_n24312), .B(new_n24311), .Y(new_n27521));
  xor_4  g25173(.A(new_n27521), .B(new_n24320), .Y(n21168));
  xor_4  g25174(.A(new_n8536), .B(new_n8535_1), .Y(n21173));
  nand_5 g25175(.A(new_n5089), .B(new_n5088), .Y(new_n27524));
  xnor_4 g25176(.A(new_n27524), .B(new_n5119), .Y(n21176));
  nand_5 g25177(.A(new_n16597), .B(new_n16596_1), .Y(new_n27526));
  xnor_4 g25178(.A(new_n27526), .B(new_n16606), .Y(n21182));
  nand_5 g25179(.A(new_n25323), .B(new_n25280), .Y(new_n27528));
  nand_5 g25180(.A(new_n27528), .B(new_n25279), .Y(new_n27529));
  xor_4  g25181(.A(new_n27529), .B(new_n25278), .Y(n21193));
  nand_5 g25182(.A(new_n10921), .B(new_n10916), .Y(new_n27531));
  xor_4  g25183(.A(new_n27531), .B(new_n19882), .Y(n21203));
  xor_4  g25184(.A(new_n19046), .B(new_n2618), .Y(n21225));
  nand_5 g25185(.A(new_n22868), .B(new_n22803), .Y(new_n27534));
  xnor_4 g25186(.A(new_n27534), .B(new_n22866), .Y(n21238));
  nand_5 g25187(.A(new_n15984), .B(new_n15985), .Y(new_n27536));
  xnor_4 g25188(.A(new_n27536), .B(new_n16007), .Y(n21254));
  nand_5 g25189(.A(new_n23084), .B(new_n23083), .Y(new_n27538));
  xnor_4 g25190(.A(new_n27538), .B(new_n23118), .Y(n21298));
  xor_4  g25191(.A(new_n22846), .B(new_n20559), .Y(n21302));
  nand_5 g25192(.A(new_n22915), .B(new_n22914_1), .Y(new_n27541));
  xnor_4 g25193(.A(new_n27541), .B(new_n22917), .Y(n21349));
  nand_5 g25194(.A(new_n18600), .B(new_n18601), .Y(new_n27543));
  xnor_4 g25195(.A(new_n27543), .B(new_n18615), .Y(n21365));
  nand_5 g25196(.A(new_n17576), .B(new_n17575), .Y(new_n27545));
  xor_4  g25197(.A(new_n27545), .B(new_n17590), .Y(n21367));
  nor_5  g25198(.A(new_n13689), .B(new_n13688), .Y(new_n27547));
  xor_4  g25199(.A(new_n27547), .B(new_n13729), .Y(n21396));
  nand_5 g25200(.A(new_n8700), .B(new_n8699), .Y(new_n27549));
  xor_4  g25201(.A(new_n27549), .B(new_n8754), .Y(n21399));
  xor_4  g25202(.A(new_n3691), .B(new_n3687), .Y(n21404));
  nand_5 g25203(.A(new_n9703), .B(new_n9702), .Y(new_n27552));
  xor_4  g25204(.A(new_n27552), .B(new_n9720), .Y(n21446));
  or_5   g25205(.A(new_n13520), .B(new_n13519), .Y(new_n27554));
  xor_4  g25206(.A(new_n27554), .B(new_n13528), .Y(n21472));
  nand_5 g25207(.A(new_n8497), .B(new_n8496), .Y(new_n27556));
  xnor_4 g25208(.A(new_n27556), .B(new_n8557), .Y(n21525));
  nand_5 g25209(.A(new_n19915), .B(new_n19914), .Y(new_n27558));
  xor_4  g25210(.A(new_n27558), .B(new_n19939), .Y(n21549));
  nand_5 g25211(.A(new_n22742), .B(new_n22743), .Y(new_n27560));
  xnor_4 g25212(.A(new_n27560), .B(new_n22745), .Y(n21615));
  nor_5  g25213(.A(new_n25736), .B(new_n9009), .Y(new_n27562));
  xor_4  g25214(.A(new_n25736), .B(new_n9011), .Y(new_n27563));
  nand_5 g25215(.A(new_n20318), .B(new_n20290), .Y(new_n27564));
  nand_5 g25216(.A(new_n27564), .B(new_n20289), .Y(new_n27565));
  nor_5  g25217(.A(new_n27565), .B(new_n27563), .Y(new_n27566));
  nor_5  g25218(.A(new_n27566), .B(new_n27562), .Y(n21628));
  nor_5  g25219(.A(new_n24913), .B(new_n24337), .Y(new_n27568));
  xor_4  g25220(.A(new_n24913), .B(new_n24355), .Y(new_n27569));
  nand_5 g25221(.A(new_n26438), .B(new_n26435), .Y(new_n27570));
  nand_5 g25222(.A(new_n27570), .B(new_n26434), .Y(new_n27571));
  nor_5  g25223(.A(new_n27571), .B(new_n27569), .Y(new_n27572));
  nor_5  g25224(.A(new_n27572), .B(new_n27568), .Y(n21637));
  nand_5 g25225(.A(new_n24839), .B(new_n24838), .Y(new_n27574));
  xor_4  g25226(.A(new_n27574), .B(new_n24845), .Y(n21645));
  xor_4  g25227(.A(new_n14006), .B(new_n7449), .Y(n21665));
  nand_5 g25228(.A(new_n17249), .B(new_n17248), .Y(new_n27577));
  xnor_4 g25229(.A(new_n27577), .B(new_n17275), .Y(n21680));
  nand_5 g25230(.A(new_n25363), .B(new_n25362_1), .Y(new_n27579));
  xor_4  g25231(.A(new_n27579), .B(new_n25396), .Y(n21685));
  nor_5  g25232(.A(new_n21416), .B(new_n21415), .Y(new_n27581));
  xor_4  g25233(.A(new_n27581), .B(new_n21445), .Y(n21717));
  nand_5 g25234(.A(new_n19517), .B(new_n19518), .Y(new_n27583));
  xor_4  g25235(.A(new_n27583), .B(new_n19523_1), .Y(n21719));
  nand_5 g25236(.A(new_n21435), .B(new_n21434), .Y(new_n27585));
  xnor_4 g25237(.A(new_n27585), .B(new_n21437), .Y(n21750));
  nand_5 g25238(.A(new_n25124), .B(new_n25119_1), .Y(new_n27587));
  xor_4  g25239(.A(new_n27587), .B(new_n25121), .Y(n21765));
  nand_5 g25240(.A(new_n27481), .B(new_n27480), .Y(new_n27589));
  xor_4  g25241(.A(new_n27589), .B(new_n27483), .Y(n21800));
  nand_5 g25242(.A(new_n4751), .B(new_n4752), .Y(new_n27591));
  xor_4  g25243(.A(new_n27591), .B(new_n4758), .Y(n21820));
  nand_5 g25244(.A(new_n22417), .B(new_n22418), .Y(new_n27593));
  xnor_4 g25245(.A(new_n27593), .B(new_n22448), .Y(n21874));
  nand_5 g25246(.A(new_n15446), .B(new_n15445), .Y(new_n27595));
  xnor_4 g25247(.A(new_n27595), .B(new_n15460), .Y(n21943));
  nand_5 g25248(.A(new_n18596), .B(new_n18597), .Y(new_n27597));
  xnor_4 g25249(.A(new_n27597), .B(new_n18619), .Y(n21960));
  nand_5 g25250(.A(new_n8251), .B(new_n8250), .Y(new_n27599));
  xor_4  g25251(.A(new_n27599), .B(new_n8253), .Y(n21976));
  nand_5 g25252(.A(new_n13086), .B(new_n13088), .Y(new_n27601));
  xnor_4 g25253(.A(new_n27601), .B(new_n13116_1), .Y(n21986));
  nand_5 g25254(.A(new_n12838), .B(new_n12837), .Y(new_n27603));
  xor_4  g25255(.A(new_n27603), .B(new_n12883), .Y(n22016));
  nor_5  g25256(.A(new_n21431), .B(new_n21430), .Y(new_n27605));
  xor_4  g25257(.A(new_n27605), .B(new_n21439), .Y(n22027));
  nand_5 g25258(.A(new_n15188), .B(new_n15187), .Y(new_n27607));
  xnor_4 g25259(.A(new_n27607), .B(new_n15198), .Y(n22050));
  nand_5 g25260(.A(new_n4580), .B(new_n4577), .Y(new_n27609));
  nand_5 g25261(.A(new_n27609), .B(new_n4581), .Y(n22063));
  nand_5 g25262(.A(new_n24316), .B(new_n24315), .Y(new_n27611));
  xnor_4 g25263(.A(new_n27611), .B(new_n24318), .Y(n22076));
  nor_5  g25264(.A(new_n23361), .B(new_n15930), .Y(new_n27613));
  nor_5  g25265(.A(new_n23738), .B(new_n23720), .Y(new_n27614));
  nor_5  g25266(.A(new_n27614), .B(new_n27613), .Y(n22090));
  nand_5 g25267(.A(new_n25951), .B(new_n25952), .Y(new_n27616));
  xnor_4 g25268(.A(new_n27616), .B(new_n25958), .Y(n22107));
  nand_5 g25269(.A(new_n20464), .B(new_n20463), .Y(new_n27618));
  xnor_4 g25270(.A(new_n27618), .B(new_n20496), .Y(n22113));
  not_8  g25271(.A(new_n16016), .Y(new_n27620));
  nor_5  g25272(.A(new_n27620), .B(new_n15958_1), .Y(new_n27621));
  not_8  g25273(.A(new_n16015), .Y(new_n27622));
  nor_5  g25274(.A(new_n27622), .B(new_n15959), .Y(new_n27623));
  nor_5  g25275(.A(new_n27623), .B(new_n27621), .Y(n22124));
  nor_5  g25276(.A(new_n26750), .B(new_n22300), .Y(new_n27625));
  nor_5  g25277(.A(new_n26753), .B(new_n26751), .Y(new_n27626));
  nor_5  g25278(.A(new_n27626), .B(new_n27625), .Y(n22126));
  xor_4  g25279(.A(new_n27491), .B(new_n25982), .Y(n22130));
  nand_5 g25280(.A(new_n20708), .B(new_n20709_1), .Y(new_n27629));
  xor_4  g25281(.A(new_n27629), .B(new_n20711), .Y(n22144));
  or_5   g25282(.A(new_n26425), .B(new_n26417), .Y(new_n27631));
  nand_5 g25283(.A(new_n27631), .B(new_n26426), .Y(n22150));
  nand_5 g25284(.A(new_n22656), .B(new_n22655), .Y(new_n27633));
  xnor_4 g25285(.A(new_n27633), .B(new_n22663), .Y(n22157));
  or_5   g25286(.A(new_n27211), .B(new_n27210), .Y(new_n27635));
  xor_4  g25287(.A(new_n27635), .B(new_n27214), .Y(n22213));
  nand_5 g25288(.A(new_n12087), .B(new_n12086), .Y(new_n27637));
  xor_4  g25289(.A(new_n27637), .B(new_n12089), .Y(n22283));
  nand_5 g25290(.A(new_n23397), .B(new_n23398), .Y(new_n27639));
  xnor_4 g25291(.A(new_n27639), .B(new_n23400), .Y(n22311));
  nor_5  g25292(.A(new_n10177), .B(new_n10176), .Y(new_n27641));
  xor_4  g25293(.A(new_n27641), .B(new_n10248), .Y(n22317));
  nand_5 g25294(.A(new_n20224), .B(new_n20223), .Y(new_n27643));
  xor_4  g25295(.A(new_n27643), .B(new_n20238), .Y(n22341));
  or_5   g25296(.A(new_n8273), .B(new_n8190), .Y(new_n27645));
  nand_5 g25297(.A(new_n8273), .B(new_n8192), .Y(new_n27646));
  nand_5 g25298(.A(new_n27646), .B(new_n27645), .Y(new_n27647));
  not_8  g25299(.A(new_n27647), .Y(new_n27648));
  xor_4  g25300(.A(new_n27648), .B(new_n21053), .Y(n22353));
  nand_5 g25301(.A(new_n20228), .B(new_n20227), .Y(new_n27650));
  xor_4  g25302(.A(new_n27650), .B(new_n20236), .Y(n22444));
  nand_5 g25303(.A(new_n11813), .B(new_n11812), .Y(new_n27652));
  xnor_4 g25304(.A(new_n27652), .B(new_n11815), .Y(n22467));
  nor_5  g25305(.A(new_n10224), .B(new_n10221), .Y(new_n27654));
  nor_5  g25306(.A(new_n27654), .B(new_n10226), .Y(n22484));
  nand_5 g25307(.A(new_n5057), .B(new_n5055), .Y(new_n27656));
  xnor_4 g25308(.A(new_n27656), .B(new_n5129), .Y(n22489));
  nand_5 g25309(.A(new_n9574), .B(new_n9573), .Y(new_n27658));
  xor_4  g25310(.A(new_n27658), .B(new_n9627), .Y(n22494));
  nand_5 g25311(.A(new_n12066), .B(new_n12064), .Y(new_n27660));
  xnor_4 g25312(.A(new_n27660), .B(new_n12095), .Y(n22533));
  nand_5 g25313(.A(new_n25923_1), .B(new_n25922), .Y(new_n27662));
  xnor_4 g25314(.A(new_n27662), .B(new_n25925), .Y(n22584));
  nor_5  g25315(.A(new_n20722_1), .B(new_n24963), .Y(n22589));
  nand_5 g25316(.A(new_n27272), .B(new_n27271), .Y(new_n27665));
  xor_4  g25317(.A(new_n27665), .B(new_n27276), .Y(n22620));
  xor_4  g25318(.A(new_n9716), .B(new_n14779), .Y(n22623));
  nand_5 g25319(.A(new_n19652_1), .B(new_n19650), .Y(new_n27668));
  xnor_4 g25320(.A(new_n27668), .B(new_n19668), .Y(n22697));
  nand_5 g25321(.A(new_n10212), .B(new_n10213), .Y(new_n27670));
  xnor_4 g25322(.A(new_n27670), .B(new_n10238), .Y(n22714));
  nand_5 g25323(.A(new_n13796), .B(new_n13795), .Y(new_n27672));
  xor_4  g25324(.A(new_n27672), .B(new_n13853), .Y(n22761));
  nor_5  g25325(.A(new_n21913), .B(new_n21912), .Y(new_n27674));
  xor_4  g25326(.A(new_n27674), .B(new_n21928), .Y(n22779));
  nand_5 g25327(.A(new_n25902), .B(new_n25901), .Y(new_n27676));
  xnor_4 g25328(.A(new_n27676), .B(new_n25935), .Y(n22787));
  nor_5  g25329(.A(new_n2524), .B(new_n2523), .Y(new_n27678));
  xor_4  g25330(.A(new_n27678), .B(new_n2563), .Y(n22819));
  xor_4  g25331(.A(new_n10630), .B(new_n5112), .Y(n22858));
  nor_5  g25332(.A(new_n26523), .B(new_n26521), .Y(new_n27681));
  xor_4  g25333(.A(new_n27681), .B(new_n26520), .Y(n22870));
  nand_5 g25334(.A(new_n11193), .B(new_n11194), .Y(new_n27683));
  xor_4  g25335(.A(new_n27683), .B(new_n11214), .Y(n22891));
  nand_5 g25336(.A(new_n22590), .B(new_n22589_1), .Y(new_n27685));
  xor_4  g25337(.A(new_n27685), .B(new_n22607), .Y(n22897));
  nand_5 g25338(.A(new_n11753), .B(new_n11754), .Y(new_n27687));
  xor_4  g25339(.A(new_n27687), .B(new_n11832), .Y(n22903));
  nand_5 g25340(.A(new_n16569), .B(new_n16568), .Y(new_n27689));
  xor_4  g25341(.A(new_n27689), .B(new_n16621), .Y(n22907));
  nand_5 g25342(.A(new_n8235), .B(new_n8234), .Y(new_n27691));
  xor_4  g25343(.A(new_n27691), .B(new_n8259_1), .Y(n22910));
  xnor_4 g25344(.A(new_n14334), .B(new_n14329), .Y(n22914));
  xor_4  g25345(.A(new_n6541), .B(new_n6484), .Y(n22939));
  nor_5  g25346(.A(new_n22056), .B(new_n22048), .Y(new_n27695));
  xor_4  g25347(.A(new_n27695), .B(new_n22059), .Y(n22998));
  nor_5  g25348(.A(new_n10231), .B(new_n10230), .Y(new_n27697));
  xor_4  g25349(.A(new_n27697), .B(new_n14071_1), .Y(n23006));
  nand_5 g25350(.A(new_n14803), .B(new_n14804), .Y(new_n27699));
  xor_4  g25351(.A(new_n27699), .B(new_n14813), .Y(n23007));
  nand_5 g25352(.A(new_n20935_1), .B(new_n20934), .Y(new_n27701));
  xor_4  g25353(.A(new_n27701), .B(new_n20937), .Y(n23009));
  nand_5 g25354(.A(new_n19423), .B(new_n19421), .Y(new_n27703));
  xnor_4 g25355(.A(new_n27703), .B(new_n19502), .Y(n23014));
  xor_4  g25356(.A(new_n27571), .B(new_n27569), .Y(n23047));
  nand_5 g25357(.A(new_n20301_1), .B(new_n20302), .Y(new_n27706));
  xor_4  g25358(.A(new_n27706), .B(new_n20312), .Y(n23058));
  or_5   g25359(.A(new_n21331), .B(new_n12020), .Y(new_n27708));
  nand_5 g25360(.A(new_n27708), .B(new_n21333), .Y(new_n27709));
  xor_4  g25361(.A(new_n27709), .B(new_n21330), .Y(n23067));
  nand_5 g25362(.A(new_n18604), .B(new_n18605), .Y(new_n27711));
  xnor_4 g25363(.A(new_n27711), .B(new_n18611), .Y(n23238));
  nand_5 g25364(.A(new_n20025), .B(new_n20024), .Y(new_n27713));
  xor_4  g25365(.A(new_n27713), .B(new_n20039), .Y(n23247));
  nand_5 g25366(.A(new_n17392_1), .B(new_n17393), .Y(new_n27715));
  xor_4  g25367(.A(new_n27715), .B(new_n17401), .Y(n23248));
  nand_5 g25368(.A(new_n20092), .B(new_n20091), .Y(new_n27717));
  xor_4  g25369(.A(new_n27717), .B(new_n20105), .Y(n23270));
  nand_5 g25370(.A(new_n25993), .B(new_n25992), .Y(new_n27719));
  xor_4  g25371(.A(new_n27719), .B(new_n25995), .Y(n23289));
  nand_5 g25372(.A(new_n6072), .B(new_n6073), .Y(new_n27721));
  xor_4  g25373(.A(new_n27721), .B(new_n6130), .Y(n23305));
  nand_5 g25374(.A(new_n24086), .B(new_n24085_1), .Y(new_n27723));
  xor_4  g25375(.A(new_n27723), .B(new_n24088), .Y(n23341));
  xor_4  g25376(.A(new_n10803), .B(new_n5550), .Y(n23342));
  nor_5  g25377(.A(new_n24457), .B(new_n24430), .Y(new_n27726));
  nor_5  g25378(.A(new_n24456), .B(new_n24428), .Y(new_n27727));
  nor_5  g25379(.A(new_n27727), .B(new_n27726), .Y(n23355));
  nand_5 g25380(.A(new_n22149), .B(new_n22148), .Y(new_n27729));
  xnor_4 g25381(.A(new_n27729), .B(new_n22151), .Y(n23371));
  nand_5 g25382(.A(new_n17779), .B(new_n17778), .Y(new_n27731));
  xor_4  g25383(.A(new_n27731), .B(new_n17832), .Y(n23401));
  nand_5 g25384(.A(new_n15196), .B(new_n15192), .Y(new_n27733));
  xor_4  g25385(.A(new_n27733), .B(new_n15194), .Y(n23414));
  nand_5 g25386(.A(new_n20084), .B(new_n20083), .Y(new_n27735));
  xor_4  g25387(.A(new_n27735), .B(new_n20109), .Y(n23429));
  nand_5 g25388(.A(new_n24728), .B(new_n24725), .Y(new_n27737));
  xor_4  g25389(.A(new_n27737), .B(new_n23065_1), .Y(n23433));
  nand_5 g25390(.A(new_n21249), .B(new_n21248), .Y(new_n27739));
  xnor_4 g25391(.A(new_n27739), .B(new_n21263), .Y(n23434));
  nand_5 g25392(.A(new_n26762), .B(new_n26761), .Y(new_n27741));
  nand_5 g25393(.A(new_n27741), .B(new_n26763), .Y(new_n27742));
  xor_4  g25394(.A(new_n27742), .B(new_n24876), .Y(n23450));
  nand_5 g25395(.A(new_n19430), .B(new_n19428), .Y(new_n27744));
  xnor_4 g25396(.A(new_n27744), .B(new_n19500), .Y(n23471));
  nand_5 g25397(.A(new_n24064), .B(new_n24065), .Y(new_n27746));
  xor_4  g25398(.A(new_n27746), .B(new_n24098), .Y(n23480));
  xor_4  g25399(.A(new_n20549), .B(new_n20543), .Y(n23546));
  nand_5 g25400(.A(new_n23654), .B(new_n23653), .Y(new_n27749));
  xor_4  g25401(.A(new_n27749), .B(new_n23664), .Y(n23550));
  nand_5 g25402(.A(new_n8518), .B(new_n8517), .Y(new_n27751));
  xnor_4 g25403(.A(new_n27751), .B(new_n8551), .Y(n23585));
  nor_5  g25404(.A(new_n22595), .B(new_n22594), .Y(new_n27753));
  xor_4  g25405(.A(new_n27753), .B(new_n22604), .Y(n23588));
  nand_5 g25406(.A(new_n23915), .B(new_n23913_1), .Y(new_n27755));
  xnor_4 g25407(.A(new_n27755), .B(new_n23937), .Y(n23619));
  nand_5 g25408(.A(new_n3243), .B(new_n3242), .Y(new_n27757));
  xnor_4 g25409(.A(new_n27757), .B(new_n3260_1), .Y(n23624));
  nor_5  g25410(.A(new_n13711), .B(new_n13710_1), .Y(new_n27759));
  xor_4  g25411(.A(new_n27759), .B(new_n13720), .Y(n23628));
  nand_5 g25412(.A(new_n25011), .B(new_n25012), .Y(new_n27761));
  xnor_4 g25413(.A(new_n27761), .B(new_n25026), .Y(n23637));
  nand_5 g25414(.A(new_n25657), .B(new_n25656), .Y(new_n27763));
  xnor_4 g25415(.A(new_n27763), .B(new_n25659), .Y(n23663));
  not_8  g25416(.A(new_n13705), .Y(new_n27765));
  nand_5 g25417(.A(new_n27765), .B(new_n13704), .Y(new_n27766));
  xor_4  g25418(.A(new_n27766), .B(new_n13723), .Y(n23669));
  nand_5 g25419(.A(new_n15068), .B(new_n15067), .Y(new_n27768));
  xor_4  g25420(.A(new_n27768), .B(new_n15100), .Y(n23684));
  nand_5 g25421(.A(new_n21841), .B(new_n21840), .Y(new_n27770));
  xnor_4 g25422(.A(new_n27770), .B(new_n21851), .Y(n23690));
  nand_5 g25423(.A(new_n25365_1), .B(new_n25364), .Y(new_n27772));
  xor_4  g25424(.A(new_n27772), .B(new_n25394), .Y(n23714));
  nor_5  g25425(.A(new_n26799), .B(new_n26797_1), .Y(n23719));
  nand_5 g25426(.A(new_n24398), .B(new_n24397), .Y(new_n27775));
  xor_4  g25427(.A(new_n27775), .B(new_n24400), .Y(n23748));
  nand_5 g25428(.A(new_n12611), .B(new_n8279), .Y(new_n27777));
  nand_5 g25429(.A(new_n27777), .B(new_n12613), .Y(n23856));
  nand_5 g25430(.A(new_n8525), .B(new_n8524), .Y(new_n27779));
  xnor_4 g25431(.A(new_n27779), .B(new_n8549), .Y(n23883));
  nand_5 g25432(.A(new_n16602), .B(new_n16600), .Y(new_n27781));
  xnor_4 g25433(.A(new_n27781), .B(new_n16604), .Y(n23888));
  nand_5 g25434(.A(new_n3637), .B(new_n3638), .Y(new_n27783));
  xnor_4 g25435(.A(new_n27783), .B(new_n3673), .Y(n23899));
  xor_4  g25436(.A(new_n17184), .B(new_n10910), .Y(n23903));
  nand_5 g25437(.A(new_n14761), .B(new_n14760), .Y(new_n27786));
  xor_4  g25438(.A(new_n27786), .B(new_n14792), .Y(n23924));
  nand_5 g25439(.A(new_n19124), .B(new_n19123), .Y(new_n27788));
  xnor_4 g25440(.A(new_n27788), .B(new_n19133), .Y(n23935));
  nand_5 g25441(.A(new_n15080), .B(new_n15079), .Y(new_n27790));
  xor_4  g25442(.A(new_n27790), .B(new_n15096), .Y(n23942));
  nor_5  g25443(.A(new_n20334), .B(new_n20332), .Y(new_n27792));
  xor_4  g25444(.A(new_n27792), .B(new_n20342), .Y(n23954));
  nor_5  g25445(.A(new_n21503), .B(new_n21502), .Y(new_n27794));
  xor_4  g25446(.A(new_n27794), .B(new_n21526), .Y(n23958));
  nand_5 g25447(.A(new_n25523_1), .B(new_n25522), .Y(new_n27796));
  xor_4  g25448(.A(new_n27796), .B(new_n10266), .Y(n23986));
  nand_5 g25449(.A(new_n19534), .B(new_n19535), .Y(new_n27798));
  xnor_4 g25450(.A(new_n27798), .B(new_n19540), .Y(n24002));
  nand_5 g25451(.A(new_n14957), .B(new_n14956), .Y(new_n27800));
  xor_4  g25452(.A(new_n27800), .B(new_n14965), .Y(n24039));
  nand_5 g25453(.A(new_n26735), .B(new_n26734), .Y(new_n27802));
  xnor_4 g25454(.A(new_n27802), .B(new_n26737), .Y(n24052));
  nand_5 g25455(.A(new_n23306), .B(new_n23307), .Y(new_n27804));
  xor_4  g25456(.A(new_n27804), .B(new_n23329), .Y(n24092));
  nand_5 g25457(.A(new_n17956_1), .B(new_n17955), .Y(new_n27806));
  xnor_4 g25458(.A(new_n27806), .B(new_n17972), .Y(n24096));
  nand_5 g25459(.A(new_n14057), .B(new_n14058), .Y(new_n27808));
  xnor_4 g25460(.A(new_n27808), .B(new_n14084), .Y(n24097));
  nand_5 g25461(.A(new_n13695), .B(new_n13693), .Y(new_n27810));
  xnor_4 g25462(.A(new_n27810), .B(new_n13727), .Y(n24105));
  nand_5 g25463(.A(new_n20900), .B(new_n20901), .Y(new_n27812));
  xor_4  g25464(.A(new_n27812), .B(new_n20921), .Y(n24119));
  nand_5 g25465(.A(new_n17253), .B(new_n17252), .Y(new_n27814));
  xnor_4 g25466(.A(new_n27814), .B(new_n17273), .Y(n24133));
  nand_5 g25467(.A(new_n22823), .B(new_n22821), .Y(new_n27816));
  xnor_4 g25468(.A(new_n27816), .B(new_n22858_1), .Y(n24141));
  nand_5 g25469(.A(new_n24288), .B(new_n24287), .Y(new_n27818));
  xor_4  g25470(.A(new_n27818), .B(new_n24331), .Y(n24145));
  nand_5 g25471(.A(new_n25096), .B(new_n25095), .Y(new_n27820));
  xor_4  g25472(.A(new_n27820), .B(new_n25098), .Y(n24146));
  nor_5  g25473(.A(new_n14641), .B(new_n14640), .Y(new_n27822));
  xor_4  g25474(.A(new_n27822), .B(new_n14709), .Y(n24155));
  or_5   g25475(.A(new_n27052), .B(new_n27050), .Y(new_n27824));
  xor_4  g25476(.A(new_n27824), .B(new_n27054), .Y(n24160));
  nand_5 g25477(.A(new_n10599), .B(new_n10597), .Y(new_n27826));
  xnor_4 g25478(.A(new_n27826), .B(new_n10643), .Y(n24167));
  nand_5 g25479(.A(new_n16593), .B(new_n16592), .Y(new_n27828));
  xnor_4 g25480(.A(new_n27828), .B(new_n16608_1), .Y(n24177));
  xor_4  g25481(.A(new_n26859), .B(new_n26857), .Y(n24228));
  nand_5 g25482(.A(new_n20220), .B(new_n20219), .Y(new_n27831));
  xor_4  g25483(.A(new_n27831), .B(new_n20240), .Y(n24258));
  xor_4  g25484(.A(new_n21053), .B(new_n8273), .Y(new_n27833));
  nor_5  g25485(.A(new_n27833), .B(new_n27648), .Y(n24260));
  nand_5 g25486(.A(new_n21905_1), .B(new_n21903), .Y(new_n27835));
  xor_4  g25487(.A(new_n27835), .B(new_n21933), .Y(n24289));
  nand_5 g25488(.A(new_n5265_1), .B(new_n5264), .Y(new_n27837));
  xor_4  g25489(.A(new_n27837), .B(new_n5280), .Y(n24297));
  nand_5 g25490(.A(new_n13718), .B(new_n13717), .Y(new_n27839));
  xnor_4 g25491(.A(new_n27839), .B(new_n4258), .Y(n24307));
  nand_5 g25492(.A(new_n2542), .B(new_n2541), .Y(new_n27841));
  xor_4  g25493(.A(new_n27841), .B(new_n2556), .Y(n24342));
  nand_5 g25494(.A(new_n18598), .B(new_n18599), .Y(new_n27843));
  xnor_4 g25495(.A(new_n27843), .B(new_n18617), .Y(n24345));
  nand_5 g25496(.A(new_n10907), .B(new_n10906), .Y(new_n27845));
  xnor_4 g25497(.A(new_n27845), .B(new_n10923), .Y(n24347));
  nand_5 g25498(.A(new_n5595), .B(new_n5594), .Y(new_n27847));
  xor_4  g25499(.A(new_n27847), .B(new_n5655), .Y(n24373));
  nor_5  g25500(.A(new_n20857), .B(new_n20854), .Y(new_n27849));
  nor_5  g25501(.A(new_n27849), .B(new_n20859), .Y(n24406));
  nand_5 g25502(.A(new_n15837), .B(new_n15836), .Y(new_n27851));
  xor_4  g25503(.A(new_n27851), .B(new_n15850), .Y(n24415));
  nand_5 g25504(.A(new_n12503), .B(new_n12504), .Y(new_n27853));
  xor_4  g25505(.A(new_n27853), .B(new_n12507_1), .Y(n24421));
  nand_5 g25506(.A(new_n15633), .B(new_n15632), .Y(new_n27855));
  xnor_4 g25507(.A(new_n27855), .B(new_n15662_1), .Y(n24431));
  nand_5 g25508(.A(new_n13816), .B(new_n13815), .Y(new_n27857));
  xor_4  g25509(.A(new_n27857), .B(new_n13843), .Y(n24472));
  xor_4  g25510(.A(new_n9565), .B(new_n26001), .Y(new_n27859));
  xor_4  g25511(.A(new_n27859), .B(new_n26003), .Y(n24476));
  nand_5 g25512(.A(new_n11774), .B(new_n11775_1), .Y(new_n27861));
  xor_4  g25513(.A(new_n27861), .B(new_n11826), .Y(n24483));
  xor_4  g25514(.A(new_n15532), .B(new_n15529), .Y(n24501));
  nand_5 g25515(.A(new_n20953), .B(new_n20952), .Y(new_n27864));
  xor_4  g25516(.A(new_n27864), .B(new_n20956), .Y(n24512));
  nand_5 g25517(.A(new_n5258), .B(new_n5257), .Y(new_n27866));
  xnor_4 g25518(.A(new_n27866), .B(new_n5283), .Y(n24558));
  xor_4  g25519(.A(new_n2977), .B(new_n2976), .Y(n24576));
  xor_4  g25520(.A(new_n2968), .B(new_n2966), .Y(new_n27869));
  xor_4  g25521(.A(new_n27869), .B(new_n2978_1), .Y(n24579));
  nand_5 g25522(.A(new_n23394), .B(new_n23393), .Y(new_n27871));
  xor_4  g25523(.A(new_n27871), .B(new_n23404), .Y(n24602));
  nand_5 g25524(.A(new_n16386), .B(new_n16385), .Y(new_n27873));
  xnor_4 g25525(.A(new_n27873), .B(new_n16431), .Y(n24604));
  nand_5 g25526(.A(new_n26153), .B(new_n26152), .Y(new_n27875));
  xor_4  g25527(.A(new_n27875), .B(new_n26155), .Y(n24626));
  xor_4  g25528(.A(new_n25107), .B(new_n25057), .Y(new_n27877));
  xor_4  g25529(.A(new_n27877), .B(new_n25105), .Y(n24629));
  nand_5 g25530(.A(new_n24837), .B(new_n24836), .Y(new_n27879));
  xor_4  g25531(.A(new_n27879), .B(new_n24847), .Y(n24636));
  not_8  g25532(.A(new_n24546), .Y(new_n27881));
  nand_5 g25533(.A(new_n27881), .B(new_n24545), .Y(new_n27882));
  xor_4  g25534(.A(new_n27882), .B(new_n24548), .Y(n24715));
  or_5   g25535(.A(new_n23279), .B(new_n23278), .Y(new_n27884));
  xor_4  g25536(.A(new_n27884), .B(new_n23341_1), .Y(n24723));
  nor_5  g25537(.A(new_n19512), .B(new_n19509), .Y(new_n27886));
  xor_4  g25538(.A(new_n27886), .B(new_n19506), .Y(n24749));
  nand_5 g25539(.A(new_n23302), .B(new_n23303), .Y(new_n27888));
  xor_4  g25540(.A(new_n27888), .B(new_n23331), .Y(n24758));
  nand_5 g25541(.A(new_n26226), .B(new_n26225), .Y(new_n27890));
  xnor_4 g25542(.A(new_n27890), .B(new_n26228), .Y(n24784));
  nand_5 g25543(.A(new_n18769), .B(new_n18768), .Y(new_n27892));
  xor_4  g25544(.A(new_n27892), .B(new_n18771), .Y(n24807));
  xor_4  g25545(.A(new_n11266_1), .B(new_n9068), .Y(n24826));
  nand_5 g25546(.A(new_n8712), .B(new_n8711), .Y(new_n27895));
  xor_4  g25547(.A(new_n27895), .B(new_n8750), .Y(n24840));
  nand_5 g25548(.A(new_n11588), .B(new_n11587), .Y(new_n27897));
  xor_4  g25549(.A(new_n27897), .B(new_n11603), .Y(n24841));
  nand_5 g25550(.A(new_n5838), .B(new_n5837), .Y(new_n27899));
  xor_4  g25551(.A(new_n27899), .B(new_n5851), .Y(n24853));
  nand_5 g25552(.A(new_n3229), .B(new_n3228_1), .Y(new_n27901));
  xnor_4 g25553(.A(new_n27901), .B(new_n3264), .Y(n24857));
  nand_5 g25554(.A(new_n7264), .B(new_n7262), .Y(new_n27903));
  xnor_4 g25555(.A(new_n27903), .B(new_n7282), .Y(n24887));
  nand_5 g25556(.A(new_n10623), .B(new_n10621), .Y(new_n27905));
  xnor_4 g25557(.A(new_n27905), .B(new_n10633), .Y(n24934));
  nand_5 g25558(.A(new_n8483), .B(new_n8482), .Y(new_n27907));
  xnor_4 g25559(.A(new_n27907), .B(new_n8561), .Y(n24998));
  nand_5 g25560(.A(new_n13457_1), .B(new_n13456_1), .Y(new_n27909));
  xor_4  g25561(.A(new_n27909), .B(new_n13475), .Y(n25006));
  nand_5 g25562(.A(new_n23724), .B(new_n23723), .Y(new_n27911));
  xor_4  g25563(.A(new_n27911), .B(new_n23734), .Y(n25032));
  nand_5 g25564(.A(new_n18711), .B(new_n18710), .Y(new_n27913));
  xnor_4 g25565(.A(new_n27913), .B(new_n18731), .Y(n25062));
  nor_5  g25566(.A(new_n22464), .B(new_n22462), .Y(new_n27915));
  xor_4  g25567(.A(new_n27915), .B(new_n22461), .Y(n25083));
  nand_5 g25568(.A(new_n15090), .B(new_n15089), .Y(new_n27917));
  xor_4  g25569(.A(new_n27917), .B(new_n15092), .Y(n25097));
  nand_5 g25570(.A(new_n20538), .B(new_n20537), .Y(new_n27919));
  xor_4  g25571(.A(new_n27919), .B(new_n20540), .Y(n25133));
  nand_5 g25572(.A(new_n21245), .B(new_n21244), .Y(new_n27921));
  xnor_4 g25573(.A(new_n27921), .B(new_n21265), .Y(n25155));
  nand_5 g25574(.A(new_n27489), .B(new_n27477), .Y(new_n27923));
  xor_4  g25575(.A(new_n27923), .B(new_n27486), .Y(n25181));
  nand_5 g25576(.A(new_n23722), .B(new_n23721), .Y(new_n27925));
  xor_4  g25577(.A(new_n27925), .B(new_n23736), .Y(n25200));
  nand_5 g25578(.A(new_n24560), .B(new_n24558_1), .Y(new_n27927));
  xnor_4 g25579(.A(new_n27927), .B(new_n24529), .Y(n25209));
  nand_5 g25580(.A(new_n17476), .B(new_n17477), .Y(new_n27929));
  xor_4  g25581(.A(new_n27929), .B(new_n17485), .Y(n25215));
  xor_4  g25582(.A(new_n21057), .B(new_n21055), .Y(n25244));
  nand_5 g25583(.A(new_n20600), .B(new_n20601), .Y(new_n27932));
  xnor_4 g25584(.A(new_n27932), .B(new_n20621), .Y(n25254));
  nand_5 g25585(.A(new_n23905), .B(new_n23906), .Y(new_n27934));
  xnor_4 g25586(.A(new_n27934), .B(new_n23941), .Y(n25256));
  or_5   g25587(.A(new_n26690), .B(new_n26686), .Y(new_n27936));
  xor_4  g25588(.A(new_n27936), .B(new_n26689), .Y(n25293));
  nand_5 g25589(.A(new_n23923_1), .B(new_n23924_1), .Y(new_n27938));
  xnor_4 g25590(.A(new_n27938), .B(new_n23933), .Y(n25328));
  xor_4  g25591(.A(new_n12866), .B(new_n4757), .Y(n25332));
  xor_4  g25592(.A(new_n26237_1), .B(new_n26212), .Y(new_n27941));
  nor_5  g25593(.A(new_n27941), .B(new_n26238), .Y(n25337));
  nand_5 g25594(.A(new_n13270_1), .B(new_n13268), .Y(new_n27943));
  xor_4  g25595(.A(new_n27943), .B(new_n13272), .Y(n25356));
  nand_5 g25596(.A(new_n10419), .B(new_n10418), .Y(new_n27945));
  xor_4  g25597(.A(new_n27945), .B(new_n10435), .Y(n25362));
  nor_5  g25598(.A(new_n16723), .B(new_n16722_1), .Y(new_n27947));
  xor_4  g25599(.A(new_n27947), .B(new_n16749), .Y(n25412));
  nand_5 g25600(.A(new_n17816), .B(new_n17814), .Y(new_n27949));
  xor_4  g25601(.A(new_n27949), .B(new_n17822), .Y(n25460));
  nand_5 g25602(.A(new_n8511), .B(new_n8510_1), .Y(new_n27951));
  xnor_4 g25603(.A(new_n27951), .B(new_n8553), .Y(n25468));
  nand_5 g25604(.A(new_n16718), .B(new_n16716), .Y(new_n27953));
  xor_4  g25605(.A(new_n27953), .B(new_n16752), .Y(n25499));
  nand_5 g25606(.A(new_n22845), .B(new_n22844), .Y(new_n27955));
  xor_4  g25607(.A(new_n27955), .B(new_n22848), .Y(n25513));
  nand_5 g25608(.A(new_n14059_1), .B(new_n14060), .Y(new_n27957));
  xnor_4 g25609(.A(new_n27957), .B(new_n14082), .Y(n25518));
  nand_5 g25610(.A(new_n15430), .B(new_n15429), .Y(new_n27959));
  xnor_4 g25611(.A(new_n27959), .B(new_n15468), .Y(n25532));
  nand_5 g25612(.A(new_n23207), .B(new_n23206), .Y(new_n27961));
  xnor_4 g25613(.A(new_n27961), .B(new_n23227), .Y(n25539));
  nand_5 g25614(.A(new_n19657), .B(new_n19655), .Y(new_n27963));
  xnor_4 g25615(.A(new_n27963), .B(new_n19666), .Y(n25550));
  nand_5 g25616(.A(new_n24076), .B(new_n24077), .Y(new_n27965));
  xor_4  g25617(.A(new_n27965), .B(new_n24092_1), .Y(n25611));
  nand_5 g25618(.A(new_n6113), .B(new_n6111), .Y(new_n27967));
  xor_4  g25619(.A(new_n27967), .B(new_n6118), .Y(n25614));
  nand_5 g25620(.A(new_n14764), .B(new_n14763_1), .Y(new_n27969));
  xor_4  g25621(.A(new_n27969), .B(new_n14790_1), .Y(n25619));
  nor_5  g25622(.A(new_n26549), .B(new_n26545), .Y(new_n27971));
  not_8  g25623(.A(new_n26547), .Y(new_n27972));
  nor_5  g25624(.A(new_n27972), .B(new_n26544), .Y(new_n27973));
  nor_5  g25625(.A(new_n27973), .B(new_n27971), .Y(n25665));
  nand_5 g25626(.A(new_n10608), .B(new_n10606), .Y(new_n27975));
  xnor_4 g25627(.A(new_n27975), .B(new_n10639), .Y(n25706));
  nor_5  g25628(.A(new_n27446), .B(new_n27444), .Y(new_n27977));
  xor_4  g25629(.A(new_n27977), .B(new_n27443), .Y(n25719));
  nand_5 g25630(.A(new_n11169), .B(new_n11170), .Y(new_n27979));
  xor_4  g25631(.A(new_n27979), .B(new_n11222), .Y(n25756));
  nor_5  g25632(.A(new_n15104), .B(new_n15056), .Y(new_n27981));
  nor_5  g25633(.A(new_n15103), .B(new_n15053_1), .Y(new_n27982));
  nor_5  g25634(.A(new_n27982), .B(new_n27981), .Y(n25758));
  nor_5  g25635(.A(new_n17184), .B(new_n6554), .Y(new_n27984));
  nor_5  g25636(.A(new_n27984), .B(new_n17186), .Y(n25773));
  nand_5 g25637(.A(new_n23843), .B(new_n23844), .Y(new_n27986));
  xor_4  g25638(.A(new_n27986), .B(new_n20489_1), .Y(n25784));
  nand_5 g25639(.A(new_n9590), .B(new_n9589), .Y(new_n27988));
  xor_4  g25640(.A(new_n27988), .B(new_n9619), .Y(n25792));
  nand_5 g25641(.A(new_n7906), .B(new_n7905), .Y(new_n27990));
  xnor_4 g25642(.A(new_n27990), .B(new_n7946), .Y(n25816));
  nand_5 g25643(.A(new_n7239), .B(new_n7240), .Y(new_n27992));
  xnor_4 g25644(.A(new_n27992), .B(new_n7288), .Y(n25826));
  xor_4  g25645(.A(new_n14300), .B(new_n14298), .Y(n25839));
  nand_5 g25646(.A(new_n16195), .B(new_n16194), .Y(new_n27995));
  xor_4  g25647(.A(new_n27995), .B(new_n16251), .Y(n25840));
  nand_5 g25648(.A(new_n9380_1), .B(new_n9379), .Y(new_n27997));
  xnor_4 g25649(.A(new_n27997), .B(new_n9413), .Y(n25873));
  xor_4  g25650(.A(new_n27565), .B(new_n27563), .Y(n25934));
  or_5   g25651(.A(new_n24307_1), .B(new_n24306), .Y(new_n28000));
  xor_4  g25652(.A(new_n28000), .B(new_n24323_1), .Y(n25938));
  nand_5 g25653(.A(new_n24669), .B(new_n24670), .Y(new_n28002));
  xor_4  g25654(.A(new_n28002), .B(new_n24672), .Y(n25985));
  xor_4  g25655(.A(new_n16029_1), .B(new_n10423), .Y(n25994));
  nand_5 g25656(.A(new_n21278), .B(new_n21203_1), .Y(new_n28005));
  nand_5 g25657(.A(new_n28005), .B(new_n21204), .Y(n26084));
  nand_5 g25658(.A(new_n26218), .B(new_n26217), .Y(new_n28007));
  xnor_4 g25659(.A(new_n28007), .B(new_n26232), .Y(n26096));
  nor_5  g25660(.A(new_n13494_1), .B(new_n13409_1), .Y(n26111));
  nand_5 g25661(.A(new_n13449), .B(new_n13448), .Y(new_n28010));
  xor_4  g25662(.A(new_n28010), .B(new_n13479), .Y(n26113));
  nand_5 g25663(.A(new_n23345), .B(new_n23346), .Y(new_n28012));
  xnor_4 g25664(.A(new_n28012), .B(new_n23348), .Y(n26156));
  nand_5 g25665(.A(new_n19869), .B(new_n19868), .Y(new_n28014));
  xor_4  g25666(.A(new_n28014), .B(new_n19893), .Y(n26159));
  nand_5 g25667(.A(new_n3999), .B(new_n3998), .Y(new_n28016));
  xnor_4 g25668(.A(new_n28016), .B(new_n4058), .Y(n26179));
  xor_4  g25669(.A(new_n16238), .B(new_n16237), .Y(n26220));
  not_8  g25670(.A(new_n26284), .Y(new_n28019));
  nand_5 g25671(.A(new_n26290), .B(new_n28019), .Y(new_n28020));
  xor_4  g25672(.A(new_n28020), .B(new_n26286), .Y(n26229));
  nor_5  g25673(.A(new_n14662), .B(new_n14661), .Y(new_n28022));
  xor_4  g25674(.A(new_n28022), .B(new_n14703), .Y(n26237));
  nand_5 g25675(.A(new_n18286), .B(new_n18285), .Y(new_n28024));
  xnor_4 g25676(.A(new_n28024), .B(new_n18303), .Y(n26250));
  nand_5 g25677(.A(new_n24360), .B(new_n24359), .Y(new_n28026));
  xor_4  g25678(.A(new_n28026), .B(new_n24362), .Y(n26274));
  nand_5 g25679(.A(new_n18268), .B(new_n18267), .Y(new_n28028));
  xnor_4 g25680(.A(new_n28028), .B(new_n18307), .Y(n26287));
  nand_5 g25681(.A(new_n27338), .B(new_n27336), .Y(new_n28030));
  xor_4  g25682(.A(new_n28030), .B(new_n27335), .Y(n26317));
  nand_5 g25683(.A(new_n21577), .B(new_n21574), .Y(new_n28032));
  nand_5 g25684(.A(new_n28032), .B(new_n21578), .Y(new_n28033));
  xor_4  g25685(.A(new_n28033), .B(new_n21554), .Y(n26353));
  nand_5 g25686(.A(new_n23396), .B(new_n23395), .Y(new_n28035));
  xor_4  g25687(.A(new_n28035), .B(new_n23402), .Y(n26375));
  nand_5 g25688(.A(new_n26739), .B(new_n26729_1), .Y(new_n28037));
  nand_5 g25689(.A(new_n28037), .B(new_n26730), .Y(n26396));
  xor_4  g25690(.A(new_n6116), .B(new_n6114), .Y(n26429));
  nand_5 g25691(.A(new_n16792), .B(new_n16790), .Y(new_n28040));
  xor_4  g25692(.A(new_n28040), .B(new_n16809), .Y(n26431));
  nand_5 g25693(.A(new_n8199), .B(new_n8198), .Y(new_n28042));
  xor_4  g25694(.A(new_n28042), .B(new_n8271), .Y(n26439));
  nand_5 g25695(.A(new_n23658), .B(new_n23657_1), .Y(new_n28044));
  xor_4  g25696(.A(new_n28044), .B(new_n23662), .Y(n26492));
  nand_5 g25697(.A(new_n11797), .B(new_n11795), .Y(new_n28046));
  xor_4  g25698(.A(new_n28046), .B(new_n11820), .Y(n26515));
  nand_5 g25699(.A(new_n2530), .B(new_n2529), .Y(new_n28048));
  xnor_4 g25700(.A(new_n28048), .B(new_n2561_1), .Y(n26538));
  nand_5 g25701(.A(new_n17387_1), .B(new_n17388), .Y(new_n28050));
  xor_4  g25702(.A(new_n28050), .B(new_n17403), .Y(n26590));
  nor_5  g25703(.A(new_n22434), .B(new_n19476), .Y(new_n28052));
  nor_5  g25704(.A(new_n28052), .B(new_n22436), .Y(n26598));
  nor_5  g25705(.A(new_n26688), .B(new_n26682), .Y(new_n28054));
  xor_4  g25706(.A(new_n28054), .B(new_n26684), .Y(n26605));
  xor_4  g25707(.A(new_n26654), .B(new_n26649), .Y(new_n28056));
  xnor_4 g25708(.A(new_n28056), .B(new_n26651), .Y(n26656));
  nand_5 g25709(.A(new_n13468), .B(new_n13466), .Y(new_n28058));
  xor_4  g25710(.A(new_n28058), .B(new_n13471), .Y(n26674));
  nand_5 g25711(.A(new_n11037), .B(new_n11036), .Y(new_n28060));
  xor_4  g25712(.A(new_n28060), .B(new_n11057), .Y(n26675));
  nand_5 g25713(.A(new_n23638), .B(new_n23637_1), .Y(new_n28062));
  xor_4  g25714(.A(new_n28062), .B(new_n23672), .Y(n26681));
  nand_5 g25715(.A(new_n6522), .B(new_n6515), .Y(new_n28064));
  nand_5 g25716(.A(new_n6523), .B(new_n6518), .Y(new_n28065));
  nand_5 g25717(.A(new_n28065), .B(new_n28064), .Y(n26696));
  nand_5 g25718(.A(new_n17073), .B(new_n17072), .Y(new_n28067));
  xnor_4 g25719(.A(new_n28067), .B(new_n17098), .Y(n26698));
  nor_5  g25720(.A(new_n17966), .B(new_n6579), .Y(new_n28069));
  nor_5  g25721(.A(new_n28069), .B(new_n17968_1), .Y(n26707));
  nand_5 g25722(.A(new_n27246), .B(new_n27245), .Y(new_n28071));
  xor_4  g25723(.A(new_n28071), .B(new_n27248), .Y(n26719));
  nand_5 g25724(.A(new_n10618), .B(new_n10616), .Y(new_n28073));
  xnor_4 g25725(.A(new_n28073), .B(new_n10635), .Y(n26727));
  nor_5  g25726(.A(new_n24740), .B(new_n22260), .Y(new_n28075));
  nor_5  g25727(.A(new_n24743), .B(new_n24741), .Y(new_n28076));
  nor_5  g25728(.A(new_n28076), .B(new_n28075), .Y(n26729));
  nor_5  g25729(.A(new_n24774), .B(new_n24772), .Y(new_n28078));
  xor_4  g25730(.A(new_n28078), .B(new_n24776), .Y(n26745));
  nand_5 g25731(.A(new_n9049), .B(new_n9048), .Y(new_n28080));
  xor_4  g25732(.A(new_n28080), .B(new_n9092), .Y(n26775));
  nand_5 g25733(.A(new_n12165), .B(new_n12163), .Y(new_n28082));
  xor_4  g25734(.A(new_n28082), .B(new_n12187), .Y(n26780));
  xor_4  g25735(.A(new_n25232), .B(new_n25226), .Y(n26794));
  nand_5 g25736(.A(new_n3612), .B(new_n3611), .Y(new_n28085));
  xnor_4 g25737(.A(new_n28085), .B(new_n3681), .Y(n26795));
  nand_5 g25738(.A(new_n12473), .B(new_n12472), .Y(new_n28087));
  xor_4  g25739(.A(new_n28087), .B(new_n12521), .Y(n26801));
  nand_5 g25740(.A(new_n12921), .B(new_n12920), .Y(new_n28089));
  xnor_4 g25741(.A(new_n28089), .B(new_n12943), .Y(n26815));
  nand_5 g25742(.A(new_n26783), .B(new_n26782), .Y(new_n28091));
  xnor_4 g25743(.A(new_n28091), .B(new_n26785), .Y(n26847));
  nor_5  g25744(.A(new_n26979_1), .B(new_n26977), .Y(new_n28093));
  xor_4  g25745(.A(new_n28093), .B(new_n26976), .Y(n26900));
  nor_5  g25746(.A(new_n21703), .B(new_n21702), .Y(new_n28095));
  xor_4  g25747(.A(new_n28095), .B(new_n21729), .Y(n26902));
  nor_5  g25748(.A(new_n20172), .B(new_n20171), .Y(new_n28097));
  xor_4  g25749(.A(new_n28097), .B(new_n20174), .Y(n26905));
  nand_5 g25750(.A(new_n9374), .B(new_n9373), .Y(new_n28099));
  xnor_4 g25751(.A(new_n28099), .B(new_n9415), .Y(n26921));
  nand_5 g25752(.A(new_n25593), .B(new_n25592), .Y(new_n28101));
  xnor_4 g25753(.A(new_n28101), .B(new_n25612), .Y(n26923));
  nand_5 g25754(.A(new_n12615), .B(new_n12614), .Y(new_n28103));
  xor_4  g25755(.A(new_n28103), .B(new_n12617), .Y(n26929));
  xor_4  g25756(.A(new_n14625), .B(new_n14624), .Y(new_n28105));
  xor_4  g25757(.A(new_n28105), .B(new_n14713), .Y(n26930));
  nand_5 g25758(.A(new_n18277), .B(new_n18276), .Y(new_n28107));
  xnor_4 g25759(.A(new_n28107), .B(new_n18305), .Y(n26943));
  nand_5 g25760(.A(new_n16712), .B(new_n16713), .Y(new_n28109));
  xor_4  g25761(.A(new_n28109), .B(new_n16754), .Y(n26970));
  nand_5 g25762(.A(new_n24246), .B(new_n24245), .Y(new_n28111));
  xor_4  g25763(.A(new_n28111), .B(new_n24256), .Y(n27004));
  nand_5 g25764(.A(new_n12031), .B(new_n12029), .Y(new_n28113));
  xor_4  g25765(.A(new_n28113), .B(new_n12105), .Y(n27011));
  or_5   g25766(.A(new_n22398), .B(new_n22397), .Y(new_n28115));
  xor_4  g25767(.A(new_n28115), .B(new_n22459), .Y(n27019));
  nand_5 g25768(.A(new_n5629), .B(new_n5628), .Y(new_n28117));
  xor_4  g25769(.A(new_n28117), .B(new_n5645), .Y(n27031));
  nand_5 g25770(.A(new_n25283), .B(new_n25282), .Y(new_n28119));
  xnor_4 g25771(.A(new_n28119), .B(new_n25321), .Y(n27051));
  nand_5 g25772(.A(new_n20032), .B(new_n20033_1), .Y(new_n28121));
  xor_4  g25773(.A(new_n28121), .B(new_n20035), .Y(n27072));
  nand_5 g25774(.A(new_n17765), .B(new_n17764), .Y(new_n28123));
  xor_4  g25775(.A(new_n28123), .B(new_n17836), .Y(n27079));
  xor_4  g25776(.A(new_n4757), .B(new_n4754), .Y(n27096));
  nand_5 g25777(.A(new_n16408), .B(new_n16409), .Y(new_n28126));
  xnor_4 g25778(.A(new_n28126), .B(new_n16425), .Y(n27110));
  nand_5 g25779(.A(new_n15793_1), .B(new_n15792), .Y(new_n28128));
  xor_4  g25780(.A(new_n28128), .B(new_n15796), .Y(n27112));
  xor_4  g25781(.A(new_n25617), .B(new_n25107), .Y(n27130));
  nand_5 g25782(.A(new_n18719), .B(new_n18718), .Y(new_n28131));
  xnor_4 g25783(.A(new_n28131), .B(new_n18727), .Y(n27145));
  nor_5  g25784(.A(new_n19245), .B(new_n16868), .Y(new_n28133));
  nor_5  g25785(.A(new_n24945), .B(new_n24943), .Y(new_n28134));
  nor_5  g25786(.A(new_n28134), .B(new_n28133), .Y(n27158));
  nand_5 g25787(.A(new_n24471), .B(new_n24472_1), .Y(new_n28136));
  xor_4  g25788(.A(new_n28136), .B(new_n24475), .Y(n27163));
  xor_4  g25789(.A(new_n27008), .B(new_n24164), .Y(new_n28138));
  xor_4  g25790(.A(new_n28138), .B(new_n27011_1), .Y(n27194));
endmodule


