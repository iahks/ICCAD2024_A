// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Wed Aug 14 23:35:30 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519,
    pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549,
    pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559,
    pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569,
    pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579,
    pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589,
    pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599,
    pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609,
    pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639,
    pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649,
    pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659,
    pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669,
    pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679,
    pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689,
    pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699,
    pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729,
    pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739,
    pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749,
    pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759,
    pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768, pi769,
    pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778, pi779,
    pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789,
    pi790, pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818, pi819,
    pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827, pi828, pi829,
    pi830, pi831, pi832, pi833, pi834, pi835, pi836, pi837, pi838, pi839,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232,
    po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241,
    po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250,
    po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259,
    po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268,
    po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277,
    po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286,
    po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295,
    po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304,
    po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313,
    po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322,
    po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331,
    po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340,
    po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349,
    po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358,
    po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367,
    po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376,
    po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385,
    po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394,
    po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403,
    po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412,
    po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421,
    po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430,
    po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439,
    po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448,
    po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457,
    po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466,
    po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475,
    po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484,
    po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493,
    po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502,
    po1503, po1504, po1505, po1506, po1507  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518,
    pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528,
    pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558,
    pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568,
    pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578,
    pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588,
    pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598,
    pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608,
    pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618,
    pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648,
    pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658,
    pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668,
    pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678,
    pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688,
    pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698,
    pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708,
    pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738,
    pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748,
    pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758,
    pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768,
    pi769, pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778,
    pi779, pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788,
    pi789, pi790, pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798,
    pi799, pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827, pi828,
    pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836, pi837, pi838,
    pi839;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231,
    po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240,
    po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249,
    po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258,
    po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267,
    po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276,
    po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285,
    po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294,
    po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303,
    po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312,
    po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321,
    po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330,
    po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339,
    po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348,
    po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357,
    po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366,
    po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375,
    po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384,
    po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393,
    po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402,
    po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411,
    po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420,
    po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429,
    po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438,
    po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447,
    po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456,
    po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465,
    po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474,
    po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483,
    po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492,
    po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501,
    po1502, po1503, po1504, po1505, po1506, po1507;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2564, new_n2565, new_n2566,
    new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2572,
    new_n2573, new_n2575, new_n2576, new_n2577, new_n2578, new_n2579,
    new_n2580, new_n2581, new_n2582, new_n2583, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659, new_n2660, new_n2661, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703, new_n2704, new_n2705,
    new_n2706, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125, new_n3126, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161, new_n3162, new_n3163,
    new_n3164, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319,
    new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340, new_n3341, new_n3342, new_n3343,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617, new_n3618, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4024, new_n4025,
    new_n4026, new_n4027, new_n4028, new_n4029, new_n4030, new_n4031,
    new_n4032, new_n4033, new_n4034, new_n4035, new_n4036, new_n4037,
    new_n4038, new_n4039, new_n4040, new_n4041, new_n4042, new_n4043,
    new_n4044, new_n4045, new_n4046, new_n4047, new_n4048, new_n4049,
    new_n4050, new_n4051, new_n4052, new_n4053, new_n4054, new_n4055,
    new_n4056, new_n4057, new_n4058, new_n4059, new_n4060, new_n4061,
    new_n4062, new_n4063, new_n4064, new_n4065, new_n4066, new_n4067,
    new_n4068, new_n4069, new_n4070, new_n4071, new_n4072, new_n4073,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4130, new_n4131, new_n4132, new_n4133, new_n4134, new_n4135,
    new_n4136, new_n4137, new_n4138, new_n4139, new_n4140, new_n4141,
    new_n4142, new_n4143, new_n4144, new_n4145, new_n4146, new_n4147,
    new_n4148, new_n4149, new_n4150, new_n4151, new_n4152, new_n4153,
    new_n4154, new_n4155, new_n4156, new_n4157, new_n4158, new_n4159,
    new_n4160, new_n4161, new_n4162, new_n4163, new_n4164, new_n4165,
    new_n4166, new_n4167, new_n4168, new_n4169, new_n4170, new_n4171,
    new_n4172, new_n4173, new_n4174, new_n4175, new_n4176, new_n4177,
    new_n4178, new_n4179, new_n4180, new_n4181, new_n4182, new_n4183,
    new_n4184, new_n4185, new_n4186, new_n4187, new_n4188, new_n4189,
    new_n4190, new_n4191, new_n4192, new_n4193, new_n4194, new_n4195,
    new_n4196, new_n4197, new_n4198, new_n4199, new_n4200, new_n4201,
    new_n4202, new_n4203, new_n4204, new_n4205, new_n4206, new_n4207,
    new_n4208, new_n4209, new_n4210, new_n4211, new_n4212, new_n4213,
    new_n4214, new_n4215, new_n4216, new_n4217, new_n4218, new_n4219,
    new_n4220, new_n4221, new_n4222, new_n4223, new_n4224, new_n4225,
    new_n4226, new_n4227, new_n4228, new_n4229, new_n4230, new_n4231,
    new_n4232, new_n4233, new_n4234, new_n4235, new_n4236, new_n4237,
    new_n4238, new_n4239, new_n4240, new_n4241, new_n4242, new_n4243,
    new_n4244, new_n4245, new_n4246, new_n4247, new_n4248, new_n4249,
    new_n4250, new_n4251, new_n4253, new_n4254, new_n4255, new_n4256,
    new_n4257, new_n4258, new_n4259, new_n4260, new_n4261, new_n4262,
    new_n4263, new_n4264, new_n4265, new_n4266, new_n4267, new_n4268,
    new_n4269, new_n4270, new_n4271, new_n4272, new_n4273, new_n4274,
    new_n4275, new_n4276, new_n4277, new_n4278, new_n4279, new_n4280,
    new_n4281, new_n4282, new_n4283, new_n4284, new_n4285, new_n4286,
    new_n4287, new_n4288, new_n4289, new_n4290, new_n4291, new_n4292,
    new_n4293, new_n4294, new_n4295, new_n4296, new_n4297, new_n4298,
    new_n4299, new_n4300, new_n4301, new_n4302, new_n4303, new_n4304,
    new_n4305, new_n4306, new_n4307, new_n4308, new_n4309, new_n4310,
    new_n4311, new_n4312, new_n4313, new_n4314, new_n4315, new_n4316,
    new_n4317, new_n4318, new_n4319, new_n4320, new_n4321, new_n4322,
    new_n4323, new_n4324, new_n4325, new_n4326, new_n4327, new_n4328,
    new_n4329, new_n4330, new_n4331, new_n4332, new_n4333, new_n4334,
    new_n4335, new_n4336, new_n4337, new_n4338, new_n4339, new_n4340,
    new_n4341, new_n4342, new_n4343, new_n4344, new_n4345, new_n4346,
    new_n4347, new_n4348, new_n4349, new_n4350, new_n4351, new_n4352,
    new_n4353, new_n4354, new_n4355, new_n4356, new_n4357, new_n4358,
    new_n4359, new_n4360, new_n4361, new_n4362, new_n4363, new_n4364,
    new_n4365, new_n4366, new_n4367, new_n4368, new_n4369, new_n4370,
    new_n4371, new_n4372, new_n4373, new_n4374, new_n4375, new_n4376,
    new_n4377, new_n4378, new_n4379, new_n4380, new_n4381, new_n4382,
    new_n4383, new_n4384, new_n4385, new_n4386, new_n4387, new_n4388,
    new_n4389, new_n4390, new_n4391, new_n4392, new_n4393, new_n4394,
    new_n4395, new_n4396, new_n4397, new_n4398, new_n4399, new_n4400,
    new_n4401, new_n4402, new_n4403, new_n4404, new_n4405, new_n4406,
    new_n4407, new_n4408, new_n4409, new_n4410, new_n4411, new_n4412,
    new_n4413, new_n4414, new_n4415, new_n4416, new_n4417, new_n4418,
    new_n4419, new_n4420, new_n4421, new_n4422, new_n4423, new_n4424,
    new_n4425, new_n4426, new_n4427, new_n4428, new_n4429, new_n4430,
    new_n4431, new_n4432, new_n4433, new_n4434, new_n4435, new_n4436,
    new_n4437, new_n4438, new_n4439, new_n4440, new_n4441, new_n4442,
    new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448,
    new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454,
    new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496,
    new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502,
    new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508,
    new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514,
    new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520,
    new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526,
    new_n4527, new_n4528, new_n4529, new_n4530, new_n4531, new_n4533,
    new_n4534, new_n4535, new_n4536, new_n4537, new_n4538, new_n4539,
    new_n4540, new_n4541, new_n4542, new_n4543, new_n4544, new_n4545,
    new_n4546, new_n4547, new_n4548, new_n4549, new_n4550, new_n4551,
    new_n4552, new_n4553, new_n4554, new_n4555, new_n4556, new_n4557,
    new_n4558, new_n4559, new_n4560, new_n4561, new_n4562, new_n4563,
    new_n4564, new_n4565, new_n4566, new_n4567, new_n4568, new_n4569,
    new_n4570, new_n4571, new_n4572, new_n4573, new_n4574, new_n4575,
    new_n4576, new_n4577, new_n4578, new_n4579, new_n4580, new_n4581,
    new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587,
    new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593,
    new_n4594, new_n4595, new_n4596, new_n4597, new_n4598, new_n4599,
    new_n4600, new_n4601, new_n4602, new_n4603, new_n4604, new_n4605,
    new_n4606, new_n4607, new_n4608, new_n4609, new_n4610, new_n4611,
    new_n4612, new_n4613, new_n4614, new_n4615, new_n4616, new_n4617,
    new_n4618, new_n4619, new_n4620, new_n4621, new_n4622, new_n4623,
    new_n4624, new_n4625, new_n4626, new_n4627, new_n4628, new_n4629,
    new_n4630, new_n4631, new_n4632, new_n4633, new_n4634, new_n4635,
    new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641,
    new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686, new_n4687, new_n4688, new_n4689,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4716, new_n4717, new_n4718, new_n4719, new_n4720,
    new_n4721, new_n4722, new_n4723, new_n4724, new_n4725, new_n4726,
    new_n4727, new_n4728, new_n4729, new_n4730, new_n4731, new_n4732,
    new_n4733, new_n4734, new_n4735, new_n4736, new_n4737, new_n4738,
    new_n4739, new_n4740, new_n4741, new_n4742, new_n4743, new_n4744,
    new_n4745, new_n4746, new_n4747, new_n4748, new_n4749, new_n4750,
    new_n4751, new_n4752, new_n4753, new_n4754, new_n4755, new_n4756,
    new_n4757, new_n4758, new_n4759, new_n4760, new_n4761, new_n4762,
    new_n4763, new_n4764, new_n4765, new_n4766, new_n4767, new_n4768,
    new_n4769, new_n4770, new_n4771, new_n4772, new_n4773, new_n4774,
    new_n4775, new_n4776, new_n4777, new_n4778, new_n4779, new_n4780,
    new_n4781, new_n4782, new_n4783, new_n4784, new_n4785, new_n4786,
    new_n4787, new_n4788, new_n4789, new_n4790, new_n4791, new_n4792,
    new_n4793, new_n4794, new_n4795, new_n4796, new_n4797, new_n4798,
    new_n4799, new_n4800, new_n4801, new_n4802, new_n4803, new_n4804,
    new_n4805, new_n4806, new_n4807, new_n4808, new_n4809, new_n4810,
    new_n4811, new_n4812, new_n4813, new_n4814, new_n4815, new_n4816,
    new_n4817, new_n4818, new_n4819, new_n4820, new_n4821, new_n4822,
    new_n4823, new_n4824, new_n4825, new_n4826, new_n4827, new_n4828,
    new_n4829, new_n4830, new_n4831, new_n4832, new_n4833, new_n4834,
    new_n4835, new_n4836, new_n4837, new_n4838, new_n4839, new_n4840,
    new_n4841, new_n4842, new_n4843, new_n4844, new_n4845, new_n4846,
    new_n4847, new_n4848, new_n4849, new_n4850, new_n4851, new_n4852,
    new_n4853, new_n4854, new_n4855, new_n4856, new_n4857, new_n4858,
    new_n4859, new_n4860, new_n4861, new_n4862, new_n4863, new_n4864,
    new_n4865, new_n4866, new_n4867, new_n4868, new_n4869, new_n4870,
    new_n4871, new_n4872, new_n4873, new_n4874, new_n4875, new_n4876,
    new_n4877, new_n4878, new_n4879, new_n4880, new_n4881, new_n4882,
    new_n4883, new_n4884, new_n4885, new_n4886, new_n4887, new_n4888,
    new_n4889, new_n4890, new_n4891, new_n4892, new_n4893, new_n4894,
    new_n4895, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900,
    new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906,
    new_n4907, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912,
    new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918,
    new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936,
    new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942,
    new_n4943, new_n4944, new_n4945, new_n4946, new_n4947, new_n4948,
    new_n4949, new_n4950, new_n4951, new_n4952, new_n4953, new_n4954,
    new_n4955, new_n4956, new_n4957, new_n4958, new_n4959, new_n4960,
    new_n4961, new_n4962, new_n4963, new_n4964, new_n4965, new_n4966,
    new_n4967, new_n4968, new_n4969, new_n4970, new_n4971, new_n4972,
    new_n4973, new_n4974, new_n4975, new_n4976, new_n4977, new_n4978,
    new_n4979, new_n4980, new_n4981, new_n4982, new_n4983, new_n4984,
    new_n4985, new_n4986, new_n4987, new_n4988, new_n4989, new_n4990,
    new_n4991, new_n4992, new_n4993, new_n4994, new_n4995, new_n4996,
    new_n4997, new_n4998, new_n4999, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5021,
    new_n5022, new_n5023, new_n5024, new_n5025, new_n5026, new_n5027,
    new_n5028, new_n5029, new_n5030, new_n5031, new_n5032, new_n5033,
    new_n5034, new_n5035, new_n5036, new_n5037, new_n5038, new_n5039,
    new_n5040, new_n5041, new_n5042, new_n5043, new_n5044, new_n5045,
    new_n5046, new_n5047, new_n5048, new_n5049, new_n5050, new_n5051,
    new_n5052, new_n5053, new_n5054, new_n5055, new_n5056, new_n5057,
    new_n5058, new_n5059, new_n5060, new_n5061, new_n5062, new_n5063,
    new_n5064, new_n5065, new_n5066, new_n5067, new_n5068, new_n5069,
    new_n5070, new_n5071, new_n5072, new_n5073, new_n5074, new_n5075,
    new_n5076, new_n5077, new_n5078, new_n5079, new_n5080, new_n5082,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100,
    new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128, new_n5129, new_n5130,
    new_n5131, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167, new_n5168, new_n5169, new_n5170, new_n5171, new_n5172,
    new_n5173, new_n5174, new_n5175, new_n5176, new_n5177, new_n5178,
    new_n5179, new_n5180, new_n5181, new_n5182, new_n5183, new_n5184,
    new_n5185, new_n5186, new_n5187, new_n5188, new_n5189, new_n5190,
    new_n5191, new_n5192, new_n5193, new_n5194, new_n5195, new_n5196,
    new_n5197, new_n5198, new_n5199, new_n5200, new_n5201, new_n5203,
    new_n5204, new_n5205, new_n5206, new_n5207, new_n5208, new_n5209,
    new_n5210, new_n5211, new_n5212, new_n5213, new_n5214, new_n5215,
    new_n5216, new_n5217, new_n5218, new_n5219, new_n5220, new_n5221,
    new_n5222, new_n5223, new_n5224, new_n5225, new_n5226, new_n5227,
    new_n5228, new_n5229, new_n5230, new_n5231, new_n5232, new_n5233,
    new_n5234, new_n5235, new_n5236, new_n5237, new_n5238, new_n5239,
    new_n5240, new_n5241, new_n5242, new_n5243, new_n5244, new_n5245,
    new_n5246, new_n5247, new_n5248, new_n5249, new_n5250, new_n5251,
    new_n5252, new_n5253, new_n5254, new_n5255, new_n5256, new_n5257,
    new_n5258, new_n5259, new_n5260, new_n5261, new_n5262, new_n5263,
    new_n5264, new_n5265, new_n5266, new_n5267, new_n5268, new_n5269,
    new_n5270, new_n5271, new_n5272, new_n5273, new_n5274, new_n5275,
    new_n5276, new_n5277, new_n5278, new_n5279, new_n5280, new_n5281,
    new_n5282, new_n5283, new_n5284, new_n5285, new_n5286, new_n5287,
    new_n5288, new_n5289, new_n5290, new_n5291, new_n5292, new_n5293,
    new_n5294, new_n5295, new_n5296, new_n5297, new_n5298, new_n5299,
    new_n5300, new_n5301, new_n5302, new_n5303, new_n5304, new_n5305,
    new_n5306, new_n5307, new_n5308, new_n5309, new_n5310, new_n5311,
    new_n5312, new_n5313, new_n5314, new_n5315, new_n5316, new_n5317,
    new_n5318, new_n5319, new_n5320, new_n5321, new_n5322, new_n5323,
    new_n5324, new_n5325, new_n5326, new_n5327, new_n5328, new_n5329,
    new_n5330, new_n5331, new_n5332, new_n5333, new_n5334, new_n5335,
    new_n5336, new_n5337, new_n5338, new_n5339, new_n5340, new_n5341,
    new_n5342, new_n5343, new_n5344, new_n5345, new_n5346, new_n5347,
    new_n5348, new_n5349, new_n5350, new_n5351, new_n5352, new_n5353,
    new_n5354, new_n5355, new_n5356, new_n5357, new_n5358, new_n5359,
    new_n5360, new_n5361, new_n5362, new_n5363, new_n5364, new_n5365,
    new_n5366, new_n5367, new_n5368, new_n5369, new_n5370, new_n5371,
    new_n5372, new_n5373, new_n5374, new_n5375, new_n5376, new_n5377,
    new_n5378, new_n5379, new_n5380, new_n5381, new_n5382, new_n5383,
    new_n5384, new_n5385, new_n5386, new_n5387, new_n5388, new_n5389,
    new_n5390, new_n5391, new_n5392, new_n5393, new_n5394, new_n5395,
    new_n5396, new_n5397, new_n5398, new_n5399, new_n5400, new_n5401,
    new_n5402, new_n5403, new_n5404, new_n5405, new_n5406, new_n5407,
    new_n5408, new_n5409, new_n5410, new_n5411, new_n5412, new_n5413,
    new_n5414, new_n5415, new_n5416, new_n5417, new_n5418, new_n5419,
    new_n5420, new_n5421, new_n5422, new_n5423, new_n5424, new_n5425,
    new_n5426, new_n5427, new_n5428, new_n5429, new_n5430, new_n5431,
    new_n5432, new_n5433, new_n5434, new_n5435, new_n5436, new_n5437,
    new_n5438, new_n5439, new_n5440, new_n5441, new_n5442, new_n5443,
    new_n5444, new_n5445, new_n5446, new_n5447, new_n5448, new_n5449,
    new_n5451, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456,
    new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462,
    new_n5463, new_n5464, new_n5465, new_n5466, new_n5467, new_n5468,
    new_n5469, new_n5470, new_n5471, new_n5472, new_n5473, new_n5474,
    new_n5475, new_n5476, new_n5477, new_n5478, new_n5479, new_n5480,
    new_n5481, new_n5482, new_n5483, new_n5484, new_n5485, new_n5486,
    new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492,
    new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498,
    new_n5499, new_n5500, new_n5501, new_n5502, new_n5503, new_n5504,
    new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510,
    new_n5511, new_n5512, new_n5513, new_n5514, new_n5515, new_n5516,
    new_n5517, new_n5518, new_n5519, new_n5520, new_n5521, new_n5522,
    new_n5523, new_n5524, new_n5525, new_n5526, new_n5527, new_n5528,
    new_n5529, new_n5530, new_n5531, new_n5532, new_n5533, new_n5534,
    new_n5535, new_n5536, new_n5537, new_n5538, new_n5539, new_n5540,
    new_n5541, new_n5542, new_n5543, new_n5544, new_n5545, new_n5546,
    new_n5547, new_n5548, new_n5549, new_n5550, new_n5551, new_n5552,
    new_n5553, new_n5554, new_n5555, new_n5556, new_n5557, new_n5558,
    new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564,
    new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570,
    new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576,
    new_n5577, new_n5578, new_n5579, new_n5580, new_n5581, new_n5582,
    new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588,
    new_n5589, new_n5590, new_n5591, new_n5592, new_n5593, new_n5594,
    new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600,
    new_n5601, new_n5602, new_n5603, new_n5604, new_n5605, new_n5606,
    new_n5607, new_n5608, new_n5609, new_n5610, new_n5611, new_n5612,
    new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618,
    new_n5619, new_n5620, new_n5621, new_n5622, new_n5623, new_n5624,
    new_n5625, new_n5626, new_n5627, new_n5628, new_n5629, new_n5630,
    new_n5631, new_n5632, new_n5633, new_n5634, new_n5635, new_n5636,
    new_n5637, new_n5638, new_n5639, new_n5640, new_n5641, new_n5642,
    new_n5643, new_n5644, new_n5645, new_n5646, new_n5647, new_n5648,
    new_n5649, new_n5650, new_n5651, new_n5652, new_n5653, new_n5654,
    new_n5655, new_n5656, new_n5657, new_n5658, new_n5659, new_n5660,
    new_n5661, new_n5662, new_n5663, new_n5664, new_n5665, new_n5666,
    new_n5667, new_n5668, new_n5669, new_n5670, new_n5671, new_n5672,
    new_n5673, new_n5674, new_n5675, new_n5676, new_n5677, new_n5678,
    new_n5679, new_n5680, new_n5681, new_n5682, new_n5683, new_n5684,
    new_n5685, new_n5686, new_n5687, new_n5688, new_n5689, new_n5690,
    new_n5691, new_n5692, new_n5693, new_n5694, new_n5695, new_n5696,
    new_n5697, new_n5698, new_n5699, new_n5700, new_n5701, new_n5702,
    new_n5703, new_n5704, new_n5705, new_n5706, new_n5707, new_n5708,
    new_n5709, new_n5710, new_n5711, new_n5712, new_n5713, new_n5714,
    new_n5715, new_n5716, new_n5717, new_n5718, new_n5719, new_n5720,
    new_n5721, new_n5722, new_n5723, new_n5724, new_n5725, new_n5726,
    new_n5727, new_n5728, new_n5729, new_n5730, new_n5731, new_n5732,
    new_n5733, new_n5734, new_n5735, new_n5736, new_n5737, new_n5738,
    new_n5739, new_n5740, new_n5741, new_n5742, new_n5743, new_n5744,
    new_n5745, new_n5746, new_n5747, new_n5748, new_n5749, new_n5750,
    new_n5751, new_n5752, new_n5753, new_n5754, new_n5755, new_n5757,
    new_n5758, new_n5759, new_n5760, new_n5761, new_n5762, new_n5763,
    new_n5764, new_n5765, new_n5766, new_n5767, new_n5768, new_n5769,
    new_n5770, new_n5771, new_n5772, new_n5773, new_n5774, new_n5775,
    new_n5776, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5807, new_n5808, new_n5809,
    new_n5810, new_n5811, new_n5812, new_n5813, new_n5814, new_n5815,
    new_n5816, new_n5817, new_n5818, new_n5819, new_n5820, new_n5821,
    new_n5822, new_n5823, new_n5824, new_n5825, new_n5826, new_n5827,
    new_n5828, new_n5829, new_n5830, new_n5831, new_n5832, new_n5833,
    new_n5834, new_n5835, new_n5836, new_n5838, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857, new_n5858, new_n5859, new_n5860,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980,
    new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986,
    new_n5987, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992,
    new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998,
    new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004,
    new_n6005, new_n6006, new_n6007, new_n6008, new_n6009, new_n6010,
    new_n6011, new_n6012, new_n6013, new_n6014, new_n6015, new_n6016,
    new_n6017, new_n6018, new_n6019, new_n6020, new_n6021, new_n6022,
    new_n6023, new_n6024, new_n6025, new_n6026, new_n6027, new_n6028,
    new_n6029, new_n6030, new_n6031, new_n6032, new_n6033, new_n6034,
    new_n6035, new_n6036, new_n6037, new_n6038, new_n6039, new_n6040,
    new_n6041, new_n6042, new_n6043, new_n6044, new_n6045, new_n6046,
    new_n6047, new_n6048, new_n6049, new_n6050, new_n6051, new_n6052,
    new_n6053, new_n6054, new_n6055, new_n6056, new_n6057, new_n6058,
    new_n6059, new_n6060, new_n6061, new_n6062, new_n6063, new_n6064,
    new_n6065, new_n6066, new_n6067, new_n6068, new_n6069, new_n6070,
    new_n6071, new_n6072, new_n6073, new_n6074, new_n6075, new_n6076,
    new_n6077, new_n6078, new_n6079, new_n6080, new_n6081, new_n6082,
    new_n6083, new_n6084, new_n6085, new_n6086, new_n6087, new_n6088,
    new_n6089, new_n6090, new_n6091, new_n6092, new_n6093, new_n6094,
    new_n6095, new_n6096, new_n6097, new_n6098, new_n6099, new_n6100,
    new_n6101, new_n6102, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254, new_n6255, new_n6256, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271, new_n6272, new_n6273, new_n6274, new_n6275,
    new_n6276, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281,
    new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287,
    new_n6288, new_n6289, new_n6290, new_n6291, new_n6292, new_n6293,
    new_n6294, new_n6295, new_n6296, new_n6297, new_n6298, new_n6299,
    new_n6300, new_n6301, new_n6302, new_n6303, new_n6304, new_n6305,
    new_n6306, new_n6307, new_n6308, new_n6309, new_n6310, new_n6311,
    new_n6312, new_n6313, new_n6314, new_n6315, new_n6316, new_n6317,
    new_n6318, new_n6319, new_n6320, new_n6321, new_n6322, new_n6323,
    new_n6324, new_n6325, new_n6326, new_n6327, new_n6328, new_n6329,
    new_n6330, new_n6331, new_n6332, new_n6333, new_n6334, new_n6335,
    new_n6336, new_n6337, new_n6338, new_n6339, new_n6340, new_n6341,
    new_n6342, new_n6343, new_n6344, new_n6345, new_n6346, new_n6347,
    new_n6348, new_n6349, new_n6350, new_n6351, new_n6352, new_n6353,
    new_n6354, new_n6355, new_n6356, new_n6357, new_n6358, new_n6359,
    new_n6360, new_n6361, new_n6362, new_n6363, new_n6364, new_n6365,
    new_n6366, new_n6367, new_n6368, new_n6369, new_n6370, new_n6371,
    new_n6372, new_n6373, new_n6374, new_n6375, new_n6376, new_n6377,
    new_n6378, new_n6379, new_n6380, new_n6381, new_n6382, new_n6383,
    new_n6384, new_n6385, new_n6386, new_n6387, new_n6388, new_n6389,
    new_n6390, new_n6391, new_n6392, new_n6393, new_n6394, new_n6395,
    new_n6396, new_n6397, new_n6398, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504,
    new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6527, new_n6528,
    new_n6529, new_n6530, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558,
    new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6568, new_n6569, new_n6570, new_n6572,
    new_n6573, new_n6574, new_n6575, new_n6576, new_n6577, new_n6578,
    new_n6579, new_n6580, new_n6581, new_n6582, new_n6583, new_n6584,
    new_n6585, new_n6586, new_n6587, new_n6588, new_n6589, new_n6590,
    new_n6591, new_n6592, new_n6593, new_n6594, new_n6595, new_n6596,
    new_n6597, new_n6598, new_n6599, new_n6600, new_n6601, new_n6602,
    new_n6603, new_n6604, new_n6605, new_n6606, new_n6607, new_n6608,
    new_n6609, new_n6610, new_n6611, new_n6612, new_n6613, new_n6614,
    new_n6615, new_n6616, new_n6617, new_n6618, new_n6619, new_n6620,
    new_n6621, new_n6622, new_n6623, new_n6624, new_n6625, new_n6626,
    new_n6627, new_n6628, new_n6629, new_n6630, new_n6631, new_n6632,
    new_n6633, new_n6634, new_n6635, new_n6636, new_n6637, new_n6638,
    new_n6639, new_n6640, new_n6641, new_n6642, new_n6643, new_n6644,
    new_n6645, new_n6646, new_n6647, new_n6648, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687,
    new_n6688, new_n6689, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6714, new_n6715, new_n6716, new_n6717, new_n6718,
    new_n6719, new_n6720, new_n6721, new_n6722, new_n6723, new_n6724,
    new_n6725, new_n6726, new_n6727, new_n6728, new_n6729, new_n6730,
    new_n6731, new_n6732, new_n6733, new_n6734, new_n6735, new_n6736,
    new_n6737, new_n6738, new_n6739, new_n6740, new_n6741, new_n6742,
    new_n6743, new_n6744, new_n6745, new_n6746, new_n6747, new_n6748,
    new_n6749, new_n6750, new_n6751, new_n6752, new_n6753, new_n6754,
    new_n6755, new_n6756, new_n6757, new_n6758, new_n6759, new_n6760,
    new_n6761, new_n6762, new_n6763, new_n6764, new_n6765, new_n6766,
    new_n6767, new_n6768, new_n6769, new_n6770, new_n6771, new_n6772,
    new_n6773, new_n6774, new_n6775, new_n6776, new_n6777, new_n6778,
    new_n6779, new_n6780, new_n6781, new_n6782, new_n6783, new_n6784,
    new_n6785, new_n6786, new_n6787, new_n6788, new_n6789, new_n6790,
    new_n6791, new_n6792, new_n6793, new_n6794, new_n6795, new_n6796,
    new_n6797, new_n6798, new_n6799, new_n6800, new_n6801, new_n6802,
    new_n6803, new_n6804, new_n6805, new_n6806, new_n6807, new_n6808,
    new_n6809, new_n6810, new_n6811, new_n6812, new_n6813, new_n6814,
    new_n6815, new_n6816, new_n6817, new_n6818, new_n6819, new_n6820,
    new_n6821, new_n6822, new_n6823, new_n6824, new_n6825, new_n6826,
    new_n6827, new_n6828, new_n6829, new_n6830, new_n6831, new_n6832,
    new_n6833, new_n6834, new_n6835, new_n6836, new_n6837, new_n6838,
    new_n6839, new_n6840, new_n6841, new_n6842, new_n6843, new_n6844,
    new_n6845, new_n6846, new_n6847, new_n6848, new_n6849, new_n6850,
    new_n6851, new_n6852, new_n6853, new_n6854, new_n6855, new_n6856,
    new_n6857, new_n6858, new_n6859, new_n6860, new_n6861, new_n6862,
    new_n6863, new_n6864, new_n6865, new_n6866, new_n6867, new_n6868,
    new_n6869, new_n6870, new_n6871, new_n6872, new_n6873, new_n6874,
    new_n6875, new_n6876, new_n6877, new_n6878, new_n6879, new_n6880,
    new_n6881, new_n6882, new_n6883, new_n6884, new_n6885, new_n6886,
    new_n6887, new_n6888, new_n6889, new_n6890, new_n6891, new_n6892,
    new_n6893, new_n6894, new_n6895, new_n6896, new_n6897, new_n6898,
    new_n6899, new_n6900, new_n6901, new_n6902, new_n6903, new_n6904,
    new_n6905, new_n6906, new_n6907, new_n6908, new_n6909, new_n6910,
    new_n6911, new_n6912, new_n6913, new_n6914, new_n6915, new_n6916,
    new_n6917, new_n6918, new_n6919, new_n6920, new_n6921, new_n6922,
    new_n6923, new_n6924, new_n6925, new_n6926, new_n6927, new_n6928,
    new_n6929, new_n6930, new_n6931, new_n6932, new_n6933, new_n6934,
    new_n6935, new_n6936, new_n6937, new_n6938, new_n6939, new_n6940,
    new_n6941, new_n6942, new_n6943, new_n6944, new_n6945, new_n6946,
    new_n6947, new_n6948, new_n6949, new_n6951, new_n6952, new_n6953,
    new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959,
    new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965,
    new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971,
    new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977,
    new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983,
    new_n6984, new_n6985, new_n6986, new_n6987, new_n6988, new_n6989,
    new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995,
    new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001,
    new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007,
    new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7013,
    new_n7014, new_n7015, new_n7016, new_n7017, new_n7018, new_n7019,
    new_n7020, new_n7021, new_n7022, new_n7023, new_n7024, new_n7025,
    new_n7026, new_n7027, new_n7028, new_n7029, new_n7030, new_n7031,
    new_n7032, new_n7033, new_n7034, new_n7035, new_n7036, new_n7037,
    new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159, new_n7160, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7254, new_n7255,
    new_n7256, new_n7257, new_n7258, new_n7259, new_n7260, new_n7261,
    new_n7262, new_n7263, new_n7264, new_n7265, new_n7266, new_n7267,
    new_n7268, new_n7269, new_n7270, new_n7271, new_n7272, new_n7273,
    new_n7274, new_n7275, new_n7276, new_n7277, new_n7278, new_n7279,
    new_n7280, new_n7281, new_n7282, new_n7283, new_n7284, new_n7285,
    new_n7286, new_n7287, new_n7288, new_n7289, new_n7290, new_n7291,
    new_n7292, new_n7293, new_n7294, new_n7295, new_n7296, new_n7297,
    new_n7298, new_n7299, new_n7300, new_n7301, new_n7302, new_n7303,
    new_n7304, new_n7305, new_n7306, new_n7307, new_n7308, new_n7309,
    new_n7310, new_n7311, new_n7312, new_n7313, new_n7314, new_n7315,
    new_n7316, new_n7317, new_n7318, new_n7319, new_n7320, new_n7321,
    new_n7322, new_n7323, new_n7324, new_n7325, new_n7326, new_n7327,
    new_n7328, new_n7329, new_n7330, new_n7331, new_n7332, new_n7333,
    new_n7334, new_n7335, new_n7336, new_n7337, new_n7338, new_n7339,
    new_n7340, new_n7341, new_n7342, new_n7343, new_n7344, new_n7345,
    new_n7346, new_n7347, new_n7348, new_n7349, new_n7350, new_n7351,
    new_n7352, new_n7353, new_n7354, new_n7355, new_n7356, new_n7357,
    new_n7358, new_n7359, new_n7360, new_n7361, new_n7362, new_n7363,
    new_n7364, new_n7365, new_n7366, new_n7367, new_n7368, new_n7369,
    new_n7370, new_n7371, new_n7372, new_n7373, new_n7374, new_n7375,
    new_n7376, new_n7377, new_n7378, new_n7379, new_n7380, new_n7381,
    new_n7382, new_n7383, new_n7384, new_n7385, new_n7386, new_n7387,
    new_n7388, new_n7389, new_n7390, new_n7391, new_n7392, new_n7393,
    new_n7394, new_n7395, new_n7396, new_n7397, new_n7398, new_n7399,
    new_n7400, new_n7401, new_n7402, new_n7403, new_n7404, new_n7405,
    new_n7406, new_n7407, new_n7408, new_n7409, new_n7410, new_n7411,
    new_n7412, new_n7413, new_n7414, new_n7415, new_n7416, new_n7417,
    new_n7418, new_n7419, new_n7420, new_n7421, new_n7422, new_n7423,
    new_n7424, new_n7425, new_n7426, new_n7427, new_n7428, new_n7429,
    new_n7430, new_n7431, new_n7432, new_n7433, new_n7434, new_n7435,
    new_n7436, new_n7437, new_n7438, new_n7439, new_n7440, new_n7441,
    new_n7442, new_n7443, new_n7444, new_n7445, new_n7446, new_n7447,
    new_n7448, new_n7449, new_n7450, new_n7451, new_n7452, new_n7453,
    new_n7454, new_n7455, new_n7456, new_n7457, new_n7458, new_n7459,
    new_n7460, new_n7461, new_n7462, new_n7463, new_n7464, new_n7465,
    new_n7466, new_n7467, new_n7468, new_n7469, new_n7470, new_n7471,
    new_n7472, new_n7473, new_n7474, new_n7475, new_n7476, new_n7477,
    new_n7478, new_n7479, new_n7480, new_n7481, new_n7482, new_n7483,
    new_n7484, new_n7485, new_n7486, new_n7487, new_n7488, new_n7489,
    new_n7490, new_n7491, new_n7492, new_n7493, new_n7494, new_n7495,
    new_n7496, new_n7497, new_n7498, new_n7499, new_n7500, new_n7501,
    new_n7502, new_n7503, new_n7504, new_n7505, new_n7506, new_n7507,
    new_n7508, new_n7509, new_n7510, new_n7511, new_n7512, new_n7514,
    new_n7515, new_n7516, new_n7517, new_n7518, new_n7519, new_n7520,
    new_n7521, new_n7522, new_n7523, new_n7524, new_n7525, new_n7526,
    new_n7527, new_n7528, new_n7529, new_n7530, new_n7531, new_n7532,
    new_n7533, new_n7534, new_n7535, new_n7536, new_n7537, new_n7538,
    new_n7539, new_n7540, new_n7541, new_n7542, new_n7543, new_n7544,
    new_n7545, new_n7546, new_n7547, new_n7548, new_n7549, new_n7550,
    new_n7551, new_n7552, new_n7553, new_n7554, new_n7555, new_n7556,
    new_n7557, new_n7558, new_n7559, new_n7560, new_n7561, new_n7562,
    new_n7563, new_n7564, new_n7565, new_n7566, new_n7567, new_n7568,
    new_n7569, new_n7570, new_n7571, new_n7572, new_n7573, new_n7574,
    new_n7575, new_n7576, new_n7577, new_n7578, new_n7579, new_n7580,
    new_n7581, new_n7582, new_n7583, new_n7584, new_n7585, new_n7586,
    new_n7587, new_n7588, new_n7589, new_n7590, new_n7591, new_n7592,
    new_n7593, new_n7594, new_n7595, new_n7596, new_n7597, new_n7598,
    new_n7599, new_n7600, new_n7601, new_n7602, new_n7603, new_n7604,
    new_n7605, new_n7606, new_n7607, new_n7608, new_n7609, new_n7610,
    new_n7611, new_n7612, new_n7613, new_n7614, new_n7615, new_n7616,
    new_n7617, new_n7618, new_n7619, new_n7620, new_n7621, new_n7622,
    new_n7623, new_n7624, new_n7625, new_n7626, new_n7627, new_n7628,
    new_n7629, new_n7630, new_n7631, new_n7632, new_n7633, new_n7634,
    new_n7635, new_n7636, new_n7637, new_n7638, new_n7639, new_n7640,
    new_n7641, new_n7642, new_n7643, new_n7644, new_n7645, new_n7646,
    new_n7647, new_n7648, new_n7649, new_n7650, new_n7651, new_n7652,
    new_n7653, new_n7654, new_n7655, new_n7656, new_n7657, new_n7658,
    new_n7659, new_n7660, new_n7661, new_n7662, new_n7663, new_n7664,
    new_n7665, new_n7666, new_n7667, new_n7668, new_n7669, new_n7670,
    new_n7671, new_n7672, new_n7673, new_n7674, new_n7675, new_n7676,
    new_n7677, new_n7678, new_n7679, new_n7680, new_n7681, new_n7682,
    new_n7683, new_n7684, new_n7685, new_n7686, new_n7687, new_n7688,
    new_n7689, new_n7690, new_n7691, new_n7692, new_n7693, new_n7694,
    new_n7695, new_n7696, new_n7697, new_n7698, new_n7700, new_n7701,
    new_n7702, new_n7703, new_n7704, new_n7705, new_n7706, new_n7707,
    new_n7708, new_n7709, new_n7710, new_n7711, new_n7712, new_n7713,
    new_n7714, new_n7715, new_n7716, new_n7717, new_n7718, new_n7719,
    new_n7720, new_n7721, new_n7722, new_n7723, new_n7724, new_n7725,
    new_n7726, new_n7727, new_n7728, new_n7729, new_n7730, new_n7731,
    new_n7732, new_n7733, new_n7734, new_n7735, new_n7736, new_n7737,
    new_n7738, new_n7739, new_n7740, new_n7741, new_n7742, new_n7743,
    new_n7744, new_n7745, new_n7746, new_n7747, new_n7748, new_n7749,
    new_n7750, new_n7751, new_n7752, new_n7753, new_n7754, new_n7755,
    new_n7756, new_n7757, new_n7758, new_n7759, new_n7760, new_n7761,
    new_n7762, new_n7763, new_n7764, new_n7765, new_n7766, new_n7767,
    new_n7768, new_n7769, new_n7770, new_n7771, new_n7772, new_n7773,
    new_n7774, new_n7775, new_n7776, new_n7777, new_n7778, new_n7779,
    new_n7780, new_n7781, new_n7782, new_n7783, new_n7784, new_n7785,
    new_n7786, new_n7787, new_n7788, new_n7789, new_n7790, new_n7791,
    new_n7792, new_n7793, new_n7794, new_n7795, new_n7796, new_n7797,
    new_n7798, new_n7799, new_n7800, new_n7801, new_n7802, new_n7803,
    new_n7804, new_n7805, new_n7806, new_n7807, new_n7808, new_n7809,
    new_n7810, new_n7811, new_n7812, new_n7813, new_n7814, new_n7815,
    new_n7816, new_n7817, new_n7818, new_n7819, new_n7820, new_n7821,
    new_n7822, new_n7823, new_n7824, new_n7825, new_n7826, new_n7827,
    new_n7828, new_n7829, new_n7830, new_n7831, new_n7832, new_n7833,
    new_n7834, new_n7835, new_n7836, new_n7837, new_n7838, new_n7839,
    new_n7840, new_n7841, new_n7842, new_n7843, new_n7844, new_n7845,
    new_n7846, new_n7847, new_n7848, new_n7849, new_n7850, new_n7851,
    new_n7852, new_n7853, new_n7854, new_n7855, new_n7856, new_n7857,
    new_n7858, new_n7859, new_n7860, new_n7861, new_n7862, new_n7863,
    new_n7864, new_n7865, new_n7866, new_n7867, new_n7868, new_n7869,
    new_n7870, new_n7871, new_n7872, new_n7873, new_n7874, new_n7875,
    new_n7876, new_n7877, new_n7878, new_n7879, new_n7880, new_n7881,
    new_n7882, new_n7883, new_n7884, new_n7885, new_n7886, new_n7887,
    new_n7888, new_n7889, new_n7890, new_n7891, new_n7892, new_n7893,
    new_n7894, new_n7895, new_n7896, new_n7897, new_n7898, new_n7899,
    new_n7900, new_n7901, new_n7902, new_n7903, new_n7904, new_n7905,
    new_n7906, new_n7907, new_n7908, new_n7909, new_n7910, new_n7911,
    new_n7912, new_n7913, new_n7914, new_n7915, new_n7916, new_n7917,
    new_n7918, new_n7919, new_n7920, new_n7921, new_n7922, new_n7923,
    new_n7924, new_n7925, new_n7926, new_n7927, new_n7928, new_n7929,
    new_n7930, new_n7931, new_n7932, new_n7933, new_n7934, new_n7935,
    new_n7936, new_n7937, new_n7938, new_n7939, new_n7940, new_n7941,
    new_n7942, new_n7943, new_n7944, new_n7945, new_n7946, new_n7947,
    new_n7948, new_n7949, new_n7950, new_n7951, new_n7952, new_n7953,
    new_n7954, new_n7955, new_n7956, new_n7957, new_n7958, new_n7959,
    new_n7960, new_n7961, new_n7962, new_n7963, new_n7964, new_n7965,
    new_n7966, new_n7967, new_n7968, new_n7969, new_n7970, new_n7971,
    new_n7972, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977,
    new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983,
    new_n7984, new_n7985, new_n7986, new_n7987, new_n7988, new_n7989,
    new_n7990, new_n7991, new_n7992, new_n7993, new_n7994, new_n7995,
    new_n7996, new_n7997, new_n7999, new_n8000, new_n8001, new_n8002,
    new_n8003, new_n8004, new_n8005, new_n8006, new_n8007, new_n8008,
    new_n8009, new_n8010, new_n8011, new_n8012, new_n8013, new_n8014,
    new_n8015, new_n8016, new_n8017, new_n8018, new_n8019, new_n8020,
    new_n8021, new_n8022, new_n8023, new_n8024, new_n8025, new_n8026,
    new_n8027, new_n8028, new_n8029, new_n8030, new_n8031, new_n8032,
    new_n8033, new_n8034, new_n8035, new_n8036, new_n8037, new_n8038,
    new_n8039, new_n8040, new_n8041, new_n8042, new_n8043, new_n8044,
    new_n8045, new_n8046, new_n8047, new_n8048, new_n8049, new_n8050,
    new_n8051, new_n8052, new_n8053, new_n8054, new_n8055, new_n8056,
    new_n8057, new_n8058, new_n8059, new_n8060, new_n8061, new_n8062,
    new_n8063, new_n8064, new_n8065, new_n8066, new_n8067, new_n8068,
    new_n8069, new_n8070, new_n8071, new_n8072, new_n8073, new_n8074,
    new_n8075, new_n8076, new_n8077, new_n8078, new_n8079, new_n8080,
    new_n8081, new_n8082, new_n8083, new_n8084, new_n8085, new_n8086,
    new_n8087, new_n8088, new_n8089, new_n8090, new_n8091, new_n8092,
    new_n8093, new_n8094, new_n8095, new_n8096, new_n8097, new_n8098,
    new_n8099, new_n8100, new_n8101, new_n8102, new_n8103, new_n8104,
    new_n8105, new_n8106, new_n8107, new_n8108, new_n8109, new_n8110,
    new_n8111, new_n8112, new_n8113, new_n8114, new_n8115, new_n8116,
    new_n8117, new_n8118, new_n8119, new_n8120, new_n8121, new_n8122,
    new_n8123, new_n8124, new_n8125, new_n8126, new_n8127, new_n8128,
    new_n8129, new_n8130, new_n8131, new_n8132, new_n8133, new_n8134,
    new_n8135, new_n8136, new_n8137, new_n8138, new_n8139, new_n8140,
    new_n8141, new_n8142, new_n8143, new_n8144, new_n8145, new_n8146,
    new_n8147, new_n8148, new_n8149, new_n8150, new_n8151, new_n8152,
    new_n8153, new_n8154, new_n8155, new_n8156, new_n8157, new_n8158,
    new_n8159, new_n8160, new_n8161, new_n8162, new_n8163, new_n8164,
    new_n8165, new_n8166, new_n8167, new_n8168, new_n8169, new_n8170,
    new_n8171, new_n8172, new_n8173, new_n8174, new_n8175, new_n8176,
    new_n8177, new_n8178, new_n8179, new_n8180, new_n8181, new_n8182,
    new_n8183, new_n8184, new_n8185, new_n8186, new_n8187, new_n8188,
    new_n8189, new_n8190, new_n8191, new_n8192, new_n8193, new_n8194,
    new_n8195, new_n8196, new_n8197, new_n8198, new_n8199, new_n8200,
    new_n8201, new_n8202, new_n8203, new_n8204, new_n8205, new_n8206,
    new_n8207, new_n8208, new_n8209, new_n8210, new_n8211, new_n8212,
    new_n8213, new_n8214, new_n8215, new_n8216, new_n8217, new_n8218,
    new_n8219, new_n8220, new_n8221, new_n8222, new_n8223, new_n8224,
    new_n8225, new_n8226, new_n8227, new_n8228, new_n8229, new_n8230,
    new_n8231, new_n8232, new_n8233, new_n8234, new_n8235, new_n8236,
    new_n8237, new_n8238, new_n8239, new_n8240, new_n8241, new_n8242,
    new_n8243, new_n8244, new_n8245, new_n8246, new_n8247, new_n8248,
    new_n8249, new_n8250, new_n8251, new_n8252, new_n8253, new_n8254,
    new_n8255, new_n8256, new_n8257, new_n8258, new_n8259, new_n8260,
    new_n8261, new_n8262, new_n8263, new_n8264, new_n8265, new_n8266,
    new_n8267, new_n8268, new_n8269, new_n8270, new_n8271, new_n8272,
    new_n8273, new_n8274, new_n8275, new_n8276, new_n8277, new_n8278,
    new_n8279, new_n8280, new_n8281, new_n8282, new_n8283, new_n8284,
    new_n8285, new_n8286, new_n8287, new_n8288, new_n8289, new_n8290,
    new_n8291, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8431, new_n8432, new_n8433, new_n8434, new_n8435, new_n8436,
    new_n8437, new_n8438, new_n8439, new_n8440, new_n8441, new_n8442,
    new_n8443, new_n8444, new_n8445, new_n8446, new_n8447, new_n8448,
    new_n8449, new_n8450, new_n8451, new_n8452, new_n8453, new_n8454,
    new_n8455, new_n8456, new_n8457, new_n8458, new_n8459, new_n8461,
    new_n8462, new_n8463, new_n8464, new_n8465, new_n8466, new_n8467,
    new_n8468, new_n8469, new_n8470, new_n8471, new_n8472, new_n8473,
    new_n8474, new_n8475, new_n8476, new_n8477, new_n8478, new_n8479,
    new_n8480, new_n8481, new_n8482, new_n8483, new_n8484, new_n8485,
    new_n8486, new_n8487, new_n8488, new_n8489, new_n8490, new_n8491,
    new_n8492, new_n8493, new_n8494, new_n8495, new_n8496, new_n8497,
    new_n8498, new_n8499, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8548, new_n8549, new_n8550, new_n8551, new_n8552, new_n8553,
    new_n8554, new_n8555, new_n8556, new_n8557, new_n8558, new_n8559,
    new_n8560, new_n8561, new_n8562, new_n8563, new_n8564, new_n8565,
    new_n8566, new_n8567, new_n8568, new_n8569, new_n8570, new_n8571,
    new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577,
    new_n8578, new_n8579, new_n8580, new_n8581, new_n8582, new_n8583,
    new_n8584, new_n8585, new_n8586, new_n8587, new_n8588, new_n8589,
    new_n8590, new_n8591, new_n8592, new_n8593, new_n8594, new_n8595,
    new_n8596, new_n8597, new_n8598, new_n8599, new_n8600, new_n8601,
    new_n8602, new_n8603, new_n8604, new_n8605, new_n8606, new_n8607,
    new_n8608, new_n8609, new_n8610, new_n8611, new_n8612, new_n8613,
    new_n8614, new_n8615, new_n8616, new_n8617, new_n8618, new_n8619,
    new_n8620, new_n8621, new_n8622, new_n8623, new_n8624, new_n8625,
    new_n8626, new_n8627, new_n8628, new_n8629, new_n8630, new_n8631,
    new_n8632, new_n8633, new_n8634, new_n8635, new_n8636, new_n8637,
    new_n8638, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8644, new_n8645, new_n8646, new_n8648, new_n8649, new_n8650,
    new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656,
    new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662,
    new_n8663, new_n8664, new_n8665, new_n8666, new_n8667, new_n8668,
    new_n8669, new_n8670, new_n8671, new_n8672, new_n8673, new_n8674,
    new_n8675, new_n8676, new_n8677, new_n8678, new_n8679, new_n8680,
    new_n8681, new_n8682, new_n8683, new_n8684, new_n8685, new_n8686,
    new_n8687, new_n8688, new_n8689, new_n8690, new_n8691, new_n8692,
    new_n8693, new_n8694, new_n8695, new_n8696, new_n8697, new_n8698,
    new_n8699, new_n8700, new_n8701, new_n8702, new_n8703, new_n8704,
    new_n8705, new_n8706, new_n8707, new_n8708, new_n8709, new_n8710,
    new_n8711, new_n8712, new_n8713, new_n8714, new_n8715, new_n8716,
    new_n8717, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744, new_n8745, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819,
    new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825,
    new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861,
    new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909,
    new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921,
    new_n8922, new_n8923, new_n8924, new_n8925, new_n8926, new_n8927,
    new_n8928, new_n8929, new_n8930, new_n8931, new_n8932, new_n8933,
    new_n8934, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8996, new_n8997, new_n8998, new_n8999, new_n9000, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9207,
    new_n9208, new_n9209, new_n9210, new_n9211, new_n9212, new_n9213,
    new_n9214, new_n9215, new_n9216, new_n9217, new_n9218, new_n9219,
    new_n9220, new_n9221, new_n9222, new_n9223, new_n9224, new_n9225,
    new_n9226, new_n9227, new_n9228, new_n9229, new_n9230, new_n9231,
    new_n9232, new_n9233, new_n9234, new_n9235, new_n9236, new_n9237,
    new_n9238, new_n9239, new_n9240, new_n9241, new_n9242, new_n9243,
    new_n9244, new_n9245, new_n9246, new_n9247, new_n9248, new_n9249,
    new_n9250, new_n9251, new_n9252, new_n9253, new_n9254, new_n9255,
    new_n9256, new_n9257, new_n9258, new_n9259, new_n9260, new_n9261,
    new_n9262, new_n9263, new_n9264, new_n9265, new_n9266, new_n9267,
    new_n9268, new_n9269, new_n9270, new_n9271, new_n9272, new_n9273,
    new_n9274, new_n9275, new_n9276, new_n9277, new_n9278, new_n9279,
    new_n9280, new_n9281, new_n9282, new_n9283, new_n9284, new_n9285,
    new_n9286, new_n9287, new_n9288, new_n9289, new_n9290, new_n9291,
    new_n9292, new_n9293, new_n9294, new_n9295, new_n9296, new_n9297,
    new_n9298, new_n9299, new_n9300, new_n9301, new_n9302, new_n9303,
    new_n9304, new_n9305, new_n9306, new_n9307, new_n9308, new_n9309,
    new_n9310, new_n9311, new_n9312, new_n9313, new_n9314, new_n9315,
    new_n9316, new_n9317, new_n9318, new_n9319, new_n9320, new_n9321,
    new_n9322, new_n9323, new_n9324, new_n9325, new_n9326, new_n9327,
    new_n9328, new_n9329, new_n9330, new_n9331, new_n9332, new_n9333,
    new_n9334, new_n9335, new_n9336, new_n9337, new_n9338, new_n9339,
    new_n9340, new_n9341, new_n9342, new_n9343, new_n9344, new_n9345,
    new_n9346, new_n9347, new_n9348, new_n9349, new_n9350, new_n9351,
    new_n9353, new_n9354, new_n9355, new_n9356, new_n9357, new_n9358,
    new_n9359, new_n9360, new_n9361, new_n9362, new_n9363, new_n9364,
    new_n9365, new_n9366, new_n9367, new_n9368, new_n9369, new_n9370,
    new_n9371, new_n9372, new_n9373, new_n9378, new_n9379, new_n9380,
    new_n9381, new_n9382, new_n9383, new_n9384, new_n9385, new_n9386,
    new_n9387, new_n9388, new_n9389, new_n9390, new_n9391, new_n9392,
    new_n9393, new_n9394, new_n9395, new_n9396, new_n9397, new_n9398,
    new_n9399, new_n9400, new_n9401, new_n9402, new_n9403, new_n9404,
    new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410,
    new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416,
    new_n9417, new_n9418, new_n9419, new_n9420, new_n9421, new_n9422,
    new_n9423, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428,
    new_n9429, new_n9430, new_n9431, new_n9432, new_n9433, new_n9434,
    new_n9435, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440,
    new_n9441, new_n9442, new_n9443, new_n9444, new_n9445, new_n9446,
    new_n9447, new_n9448, new_n9449, new_n9450, new_n9451, new_n9452,
    new_n9453, new_n9454, new_n9455, new_n9456, new_n9457, new_n9458,
    new_n9459, new_n9460, new_n9461, new_n9462, new_n9463, new_n9464,
    new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507, new_n9508, new_n9509, new_n9510, new_n9511, new_n9512,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554,
    new_n9555, new_n9556, new_n9557, new_n9558, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9567,
    new_n9568, new_n9569, new_n9570, new_n9571, new_n9572, new_n9573,
    new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579,
    new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585,
    new_n9586, new_n9587, new_n9588, new_n9589, new_n9590, new_n9591,
    new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597,
    new_n9598, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603,
    new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609,
    new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615,
    new_n9616, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621,
    new_n9622, new_n9623, new_n9624, new_n9625, new_n9626, new_n9627,
    new_n9628, new_n9629, new_n9630, new_n9631, new_n9632, new_n9633,
    new_n9634, new_n9635, new_n9636, new_n9637, new_n9638, new_n9639,
    new_n9640, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9726,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762,
    new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768,
    new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832, new_n9833, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840,
    new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846,
    new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9854,
    new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860,
    new_n9861, new_n9863, new_n9864, new_n9865, new_n9866, new_n9867,
    new_n9868, new_n9869, new_n9870, new_n9871, new_n9872, new_n9873,
    new_n9874, new_n9875, new_n9876, new_n9877, new_n9878, new_n9879,
    new_n9880, new_n9881, new_n9882, new_n9883, new_n9884, new_n9886,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022, new_n10023, new_n10024, new_n10025,
    new_n10026, new_n10027, new_n10028, new_n10029, new_n10030, new_n10031,
    new_n10032, new_n10033, new_n10034, new_n10035, new_n10036, new_n10037,
    new_n10038, new_n10039, new_n10040, new_n10041, new_n10042, new_n10043,
    new_n10044, new_n10045, new_n10046, new_n10047, new_n10048, new_n10049,
    new_n10050, new_n10051, new_n10052, new_n10053, new_n10054, new_n10055,
    new_n10056, new_n10057, new_n10058, new_n10059, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096, new_n10097,
    new_n10098, new_n10099, new_n10100, new_n10101, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111, new_n10112, new_n10113, new_n10114, new_n10115,
    new_n10116, new_n10117, new_n10118, new_n10119, new_n10120, new_n10121,
    new_n10122, new_n10123, new_n10124, new_n10125, new_n10126, new_n10127,
    new_n10128, new_n10129, new_n10130, new_n10131, new_n10132, new_n10133,
    new_n10134, new_n10135, new_n10136, new_n10137, new_n10138, new_n10139,
    new_n10140, new_n10141, new_n10142, new_n10143, new_n10144, new_n10145,
    new_n10146, new_n10147, new_n10148, new_n10149, new_n10150, new_n10151,
    new_n10152, new_n10153, new_n10154, new_n10155, new_n10156, new_n10157,
    new_n10158, new_n10159, new_n10160, new_n10161, new_n10162, new_n10163,
    new_n10164, new_n10165, new_n10166, new_n10167, new_n10168, new_n10169,
    new_n10170, new_n10171, new_n10172, new_n10173, new_n10174, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10427, new_n10428, new_n10429,
    new_n10430, new_n10431, new_n10432, new_n10433, new_n10434, new_n10435,
    new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476, new_n10477,
    new_n10478, new_n10479, new_n10480, new_n10481, new_n10482, new_n10483,
    new_n10484, new_n10485, new_n10486, new_n10487, new_n10488, new_n10489,
    new_n10490, new_n10491, new_n10492, new_n10493, new_n10494, new_n10495,
    new_n10496, new_n10497, new_n10498, new_n10499, new_n10500, new_n10501,
    new_n10502, new_n10503, new_n10504, new_n10505, new_n10506, new_n10507,
    new_n10508, new_n10509, new_n10510, new_n10511, new_n10512, new_n10513,
    new_n10514, new_n10515, new_n10516, new_n10517, new_n10518, new_n10519,
    new_n10520, new_n10521, new_n10522, new_n10523, new_n10524, new_n10525,
    new_n10526, new_n10527, new_n10528, new_n10529, new_n10530, new_n10531,
    new_n10532, new_n10533, new_n10534, new_n10535, new_n10536, new_n10537,
    new_n10538, new_n10539, new_n10540, new_n10541, new_n10542, new_n10543,
    new_n10544, new_n10545, new_n10546, new_n10547, new_n10548, new_n10549,
    new_n10550, new_n10551, new_n10552, new_n10553, new_n10554, new_n10555,
    new_n10556, new_n10557, new_n10558, new_n10559, new_n10560, new_n10561,
    new_n10562, new_n10563, new_n10564, new_n10565, new_n10566, new_n10567,
    new_n10568, new_n10569, new_n10570, new_n10571, new_n10572, new_n10573,
    new_n10574, new_n10575, new_n10576, new_n10577, new_n10578, new_n10579,
    new_n10580, new_n10581, new_n10582, new_n10583, new_n10584, new_n10585,
    new_n10586, new_n10587, new_n10588, new_n10589, new_n10590, new_n10591,
    new_n10592, new_n10593, new_n10594, new_n10595, new_n10596, new_n10597,
    new_n10598, new_n10599, new_n10600, new_n10601, new_n10602, new_n10603,
    new_n10604, new_n10605, new_n10606, new_n10607, new_n10608, new_n10609,
    new_n10610, new_n10611, new_n10612, new_n10613, new_n10614, new_n10615,
    new_n10616, new_n10617, new_n10618, new_n10619, new_n10620, new_n10621,
    new_n10622, new_n10623, new_n10624, new_n10625, new_n10626, new_n10627,
    new_n10628, new_n10629, new_n10630, new_n10631, new_n10632, new_n10633,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644, new_n10645, new_n10646,
    new_n10647, new_n10648, new_n10649, new_n10650, new_n10651, new_n10652,
    new_n10653, new_n10654, new_n10655, new_n10656, new_n10657, new_n10658,
    new_n10659, new_n10660, new_n10661, new_n10662, new_n10663, new_n10664,
    new_n10665, new_n10666, new_n10667, new_n10668, new_n10669, new_n10670,
    new_n10671, new_n10672, new_n10673, new_n10674, new_n10675, new_n10676,
    new_n10677, new_n10678, new_n10679, new_n10680, new_n10681, new_n10682,
    new_n10683, new_n10684, new_n10685, new_n10686, new_n10687, new_n10688,
    new_n10689, new_n10690, new_n10691, new_n10692, new_n10693, new_n10694,
    new_n10695, new_n10696, new_n10697, new_n10698, new_n10699, new_n10700,
    new_n10701, new_n10702, new_n10703, new_n10704, new_n10705, new_n10706,
    new_n10707, new_n10708, new_n10709, new_n10710, new_n10711, new_n10712,
    new_n10713, new_n10714, new_n10715, new_n10716, new_n10717, new_n10718,
    new_n10719, new_n10720, new_n10721, new_n10722, new_n10724, new_n10725,
    new_n10726, new_n10727, new_n10728, new_n10729, new_n10730, new_n10731,
    new_n10732, new_n10733, new_n10734, new_n10735, new_n10736, new_n10737,
    new_n10738, new_n10739, new_n10740, new_n10741, new_n10742, new_n10743,
    new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749,
    new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755,
    new_n10756, new_n10757, new_n10758, new_n10759, new_n10760, new_n10761,
    new_n10762, new_n10763, new_n10764, new_n10765, new_n10766, new_n10767,
    new_n10768, new_n10769, new_n10770, new_n10771, new_n10772, new_n10773,
    new_n10774, new_n10775, new_n10776, new_n10777, new_n10778, new_n10779,
    new_n10780, new_n10781, new_n10782, new_n10783, new_n10784, new_n10785,
    new_n10786, new_n10787, new_n10788, new_n10789, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923, new_n10924,
    new_n10925, new_n10926, new_n10927, new_n10928, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954,
    new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961, new_n10962, new_n10963, new_n10964, new_n10965, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10978, new_n10979,
    new_n10980, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023, new_n11024, new_n11025, new_n11026, new_n11027, new_n11028,
    new_n11029, new_n11030, new_n11031, new_n11032, new_n11033, new_n11034,
    new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040,
    new_n11041, new_n11042, new_n11043, new_n11044, new_n11045, new_n11046,
    new_n11048, new_n11049, new_n11050, new_n11051, new_n11052, new_n11053,
    new_n11055, new_n11056, new_n11057, new_n11058, new_n11059, new_n11060,
    new_n11061, new_n11062, new_n11063, new_n11064, new_n11065, new_n11066,
    new_n11067, new_n11068, new_n11069, new_n11070, new_n11071, new_n11072,
    new_n11073, new_n11074, new_n11075, new_n11076, new_n11077, new_n11078,
    new_n11079, new_n11080, new_n11081, new_n11082, new_n11083, new_n11084,
    new_n11085, new_n11087, new_n11088, new_n11089, new_n11090, new_n11091,
    new_n11092, new_n11093, new_n11094, new_n11095, new_n11096, new_n11097,
    new_n11098, new_n11099, new_n11100, new_n11101, new_n11102, new_n11103,
    new_n11104, new_n11105, new_n11106, new_n11107, new_n11108, new_n11109,
    new_n11110, new_n11111, new_n11112, new_n11113, new_n11114, new_n11115,
    new_n11116, new_n11117, new_n11118, new_n11119, new_n11120, new_n11121,
    new_n11122, new_n11123, new_n11124, new_n11125, new_n11126, new_n11127,
    new_n11128, new_n11129, new_n11130, new_n11131, new_n11132, new_n11133,
    new_n11134, new_n11135, new_n11136, new_n11137, new_n11138, new_n11139,
    new_n11140, new_n11141, new_n11142, new_n11143, new_n11144, new_n11145,
    new_n11146, new_n11147, new_n11148, new_n11149, new_n11150, new_n11151,
    new_n11152, new_n11153, new_n11154, new_n11155, new_n11156, new_n11157,
    new_n11158, new_n11159, new_n11160, new_n11161, new_n11162, new_n11163,
    new_n11164, new_n11165, new_n11166, new_n11167, new_n11168, new_n11169,
    new_n11170, new_n11171, new_n11172, new_n11173, new_n11174, new_n11175,
    new_n11176, new_n11177, new_n11178, new_n11179, new_n11180, new_n11181,
    new_n11182, new_n11183, new_n11184, new_n11185, new_n11186, new_n11187,
    new_n11188, new_n11189, new_n11190, new_n11191, new_n11192, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201, new_n11202, new_n11203, new_n11204, new_n11205,
    new_n11206, new_n11207, new_n11208, new_n11209, new_n11210, new_n11211,
    new_n11212, new_n11213, new_n11214, new_n11215, new_n11216, new_n11217,
    new_n11218, new_n11219, new_n11220, new_n11221, new_n11222, new_n11223,
    new_n11224, new_n11225, new_n11226, new_n11227, new_n11228, new_n11229,
    new_n11230, new_n11231, new_n11232, new_n11233, new_n11234, new_n11235,
    new_n11236, new_n11237, new_n11238, new_n11239, new_n11240, new_n11241,
    new_n11242, new_n11243, new_n11244, new_n11245, new_n11246, new_n11247,
    new_n11248, new_n11249, new_n11250, new_n11251, new_n11252, new_n11253,
    new_n11254, new_n11255, new_n11256, new_n11257, new_n11258, new_n11259,
    new_n11260, new_n11261, new_n11262, new_n11263, new_n11264, new_n11265,
    new_n11266, new_n11267, new_n11268, new_n11269, new_n11270, new_n11271,
    new_n11272, new_n11273, new_n11274, new_n11275, new_n11276, new_n11277,
    new_n11278, new_n11279, new_n11280, new_n11281, new_n11282, new_n11283,
    new_n11284, new_n11285, new_n11286, new_n11287, new_n11288, new_n11289,
    new_n11290, new_n11291, new_n11293, new_n11294, new_n11295, new_n11296,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311, new_n11312, new_n11313, new_n11314,
    new_n11315, new_n11316, new_n11317, new_n11318, new_n11319, new_n11320,
    new_n11321, new_n11322, new_n11323, new_n11324, new_n11325, new_n11326,
    new_n11327, new_n11328, new_n11329, new_n11330, new_n11331, new_n11332,
    new_n11333, new_n11334, new_n11335, new_n11336, new_n11337, new_n11338,
    new_n11339, new_n11340, new_n11341, new_n11342, new_n11343, new_n11344,
    new_n11345, new_n11346, new_n11347, new_n11348, new_n11349, new_n11350,
    new_n11351, new_n11352, new_n11353, new_n11354, new_n11356, new_n11357,
    new_n11358, new_n11359, new_n11360, new_n11361, new_n11362, new_n11363,
    new_n11364, new_n11365, new_n11366, new_n11367, new_n11368, new_n11369,
    new_n11370, new_n11371, new_n11372, new_n11374, new_n11375, new_n11376,
    new_n11377, new_n11378, new_n11379, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386, new_n11387, new_n11388,
    new_n11389, new_n11390, new_n11391, new_n11392, new_n11393, new_n11394,
    new_n11395, new_n11396, new_n11397, new_n11398, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403, new_n11404, new_n11405, new_n11406,
    new_n11407, new_n11408, new_n11409, new_n11410, new_n11411, new_n11412,
    new_n11413, new_n11414, new_n11415, new_n11416, new_n11417, new_n11418,
    new_n11419, new_n11420, new_n11421, new_n11422, new_n11423, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477, new_n11478,
    new_n11479, new_n11480, new_n11481, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486, new_n11487, new_n11488, new_n11489, new_n11490,
    new_n11491, new_n11492, new_n11493, new_n11494, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535, new_n11536,
    new_n11537, new_n11538, new_n11539, new_n11540, new_n11541, new_n11542,
    new_n11543, new_n11544, new_n11545, new_n11546, new_n11547, new_n11548,
    new_n11549, new_n11550, new_n11551, new_n11552, new_n11553, new_n11554,
    new_n11555, new_n11556, new_n11557, new_n11558, new_n11559, new_n11560,
    new_n11561, new_n11562, new_n11563, new_n11564, new_n11565, new_n11566,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579, new_n11580, new_n11581, new_n11582, new_n11583, new_n11584,
    new_n11585, new_n11586, new_n11587, new_n11588, new_n11589, new_n11590,
    new_n11591, new_n11592, new_n11593, new_n11594, new_n11595, new_n11596,
    new_n11597, new_n11598, new_n11599, new_n11600, new_n11601, new_n11602,
    new_n11603, new_n11604, new_n11605, new_n11606, new_n11607, new_n11608,
    new_n11609, new_n11610, new_n11611, new_n11612, new_n11613, new_n11614,
    new_n11615, new_n11616, new_n11617, new_n11618, new_n11619, new_n11620,
    new_n11621, new_n11622, new_n11623, new_n11624, new_n11625, new_n11626,
    new_n11627, new_n11628, new_n11629, new_n11630, new_n11631, new_n11632,
    new_n11633, new_n11634, new_n11635, new_n11636, new_n11637, new_n11638,
    new_n11640, new_n11641, new_n11642, new_n11643, new_n11644, new_n11645,
    new_n11646, new_n11647, new_n11648, new_n11649, new_n11650, new_n11651,
    new_n11652, new_n11653, new_n11654, new_n11655, new_n11656, new_n11657,
    new_n11658, new_n11659, new_n11660, new_n11661, new_n11662, new_n11663,
    new_n11664, new_n11665, new_n11666, new_n11667, new_n11668, new_n11669,
    new_n11670, new_n11671, new_n11672, new_n11673, new_n11674, new_n11675,
    new_n11676, new_n11677, new_n11678, new_n11679, new_n11680, new_n11681,
    new_n11682, new_n11683, new_n11684, new_n11685, new_n11686, new_n11687,
    new_n11688, new_n11689, new_n11690, new_n11691, new_n11692, new_n11693,
    new_n11694, new_n11695, new_n11696, new_n11697, new_n11698, new_n11699,
    new_n11700, new_n11701, new_n11702, new_n11703, new_n11704, new_n11705,
    new_n11706, new_n11707, new_n11708, new_n11709, new_n11710, new_n11711,
    new_n11712, new_n11713, new_n11714, new_n11715, new_n11716, new_n11717,
    new_n11718, new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724, new_n11725, new_n11726, new_n11727, new_n11728, new_n11729,
    new_n11730, new_n11731, new_n11732, new_n11733, new_n11734, new_n11735,
    new_n11736, new_n11737, new_n11738, new_n11739, new_n11740, new_n11741,
    new_n11742, new_n11743, new_n11744, new_n11745, new_n11746, new_n11747,
    new_n11748, new_n11749, new_n11750, new_n11751, new_n11752, new_n11753,
    new_n11754, new_n11755, new_n11756, new_n11757, new_n11758, new_n11759,
    new_n11760, new_n11761, new_n11762, new_n11763, new_n11764, new_n11765,
    new_n11766, new_n11767, new_n11768, new_n11769, new_n11770, new_n11771,
    new_n11772, new_n11773, new_n11774, new_n11775, new_n11776, new_n11777,
    new_n11778, new_n11779, new_n11780, new_n11781, new_n11782, new_n11783,
    new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789,
    new_n11790, new_n11791, new_n11792, new_n11793, new_n11794, new_n11795,
    new_n11796, new_n11797, new_n11798, new_n11799, new_n11800, new_n11801,
    new_n11802, new_n11803, new_n11804, new_n11805, new_n11806, new_n11807,
    new_n11808, new_n11809, new_n11810, new_n11811, new_n11812, new_n11813,
    new_n11814, new_n11815, new_n11816, new_n11817, new_n11818, new_n11819,
    new_n11820, new_n11821, new_n11822, new_n11823, new_n11824, new_n11825,
    new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831,
    new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837,
    new_n11838, new_n11839, new_n11840, new_n11841, new_n11842, new_n11843,
    new_n11844, new_n11845, new_n11846, new_n11847, new_n11848, new_n11849,
    new_n11850, new_n11851, new_n11852, new_n11853, new_n11854, new_n11855,
    new_n11857, new_n11860, new_n11861, new_n11862, new_n11863, new_n11864,
    new_n11868, new_n11869, new_n11870, new_n11871, new_n11872, new_n11873,
    new_n11874, new_n11875, new_n11876, new_n11877, new_n11878, new_n11879,
    new_n11880, new_n11881, new_n11882, new_n11883, new_n11884, new_n11885,
    new_n11886, new_n11887, new_n11888, new_n11889, new_n11890, new_n11891,
    new_n11892, new_n11893, new_n11894, new_n11897, new_n11898, new_n11899,
    new_n11900, new_n11901, new_n11902, new_n11903, new_n11904, new_n11905,
    new_n11906, new_n11907, new_n11908, new_n11909, new_n11910, new_n11911,
    new_n11912, new_n11913, new_n11914, new_n11915, new_n11916, new_n11917,
    new_n11918, new_n11919, new_n11920, new_n11921, new_n11922, new_n11923,
    new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965,
    new_n11966, new_n11967, new_n11968, new_n11969, new_n11970, new_n11971,
    new_n11972, new_n11973, new_n11974, new_n11975, new_n11976, new_n11977,
    new_n11978, new_n11979, new_n11980, new_n11981, new_n11982, new_n11983,
    new_n11984, new_n11985, new_n11986, new_n11987, new_n11988, new_n11989,
    new_n11990, new_n11991, new_n11992, new_n11993, new_n11994, new_n11995,
    new_n11996, new_n11997, new_n11998, new_n11999, new_n12000, new_n12001,
    new_n12002, new_n12003, new_n12004, new_n12005, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014, new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020, new_n12021, new_n12022, new_n12023, new_n12024, new_n12025,
    new_n12026, new_n12027, new_n12028, new_n12029, new_n12030, new_n12031,
    new_n12032, new_n12033, new_n12034, new_n12035, new_n12036, new_n12037,
    new_n12038, new_n12039, new_n12040, new_n12041, new_n12042, new_n12043,
    new_n12044, new_n12045, new_n12046, new_n12047, new_n12048, new_n12049,
    new_n12050, new_n12051, new_n12052, new_n12053, new_n12054, new_n12055,
    new_n12056, new_n12057, new_n12058, new_n12059, new_n12060, new_n12061,
    new_n12062, new_n12063, new_n12064, new_n12065, new_n12066, new_n12067,
    new_n12068, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075,
    new_n12076, new_n12077, new_n12078, new_n12079, new_n12080, new_n12081,
    new_n12082, new_n12083, new_n12084, new_n12085, new_n12086, new_n12087,
    new_n12088, new_n12089, new_n12090, new_n12091, new_n12092, new_n12093,
    new_n12094, new_n12095, new_n12096, new_n12097, new_n12098, new_n12099,
    new_n12100, new_n12101, new_n12102, new_n12103, new_n12104, new_n12105,
    new_n12106, new_n12107, new_n12108, new_n12109, new_n12110, new_n12111,
    new_n12112, new_n12113, new_n12114, new_n12115, new_n12116, new_n12117,
    new_n12118, new_n12119, new_n12120, new_n12121, new_n12122, new_n12123,
    new_n12124, new_n12125, new_n12126, new_n12127, new_n12128, new_n12129,
    new_n12130, new_n12131, new_n12132, new_n12133, new_n12134, new_n12135,
    new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141,
    new_n12142, new_n12143, new_n12144, new_n12145, new_n12146, new_n12147,
    new_n12148, new_n12149, new_n12150, new_n12151, new_n12152, new_n12153,
    new_n12154, new_n12155, new_n12156, new_n12157, new_n12158, new_n12159,
    new_n12160, new_n12161, new_n12162, new_n12163, new_n12164, new_n12165,
    new_n12166, new_n12167, new_n12168, new_n12169, new_n12170, new_n12171,
    new_n12172, new_n12173, new_n12174, new_n12175, new_n12176, new_n12177,
    new_n12178, new_n12179, new_n12180, new_n12181, new_n12182, new_n12183,
    new_n12184, new_n12185, new_n12186, new_n12187, new_n12188, new_n12189,
    new_n12190, new_n12191, new_n12192, new_n12193, new_n12194, new_n12195,
    new_n12196, new_n12197, new_n12198, new_n12199, new_n12200, new_n12201,
    new_n12203, new_n12205, new_n12206, new_n12207, new_n12208, new_n12209,
    new_n12210, new_n12211, new_n12212, new_n12213, new_n12214, new_n12215,
    new_n12216, new_n12217, new_n12218, new_n12219, new_n12220, new_n12221,
    new_n12222, new_n12223, new_n12224, new_n12225, new_n12226, new_n12227,
    new_n12228, new_n12229, new_n12230, new_n12231, new_n12232, new_n12233,
    new_n12234, new_n12235, new_n12236, new_n12237, new_n12238, new_n12239,
    new_n12240, new_n12241, new_n12242, new_n12243, new_n12244, new_n12245,
    new_n12246, new_n12247, new_n12248, new_n12249, new_n12250, new_n12251,
    new_n12252, new_n12253, new_n12254, new_n12255, new_n12256, new_n12257,
    new_n12258, new_n12259, new_n12260, new_n12261, new_n12262, new_n12263,
    new_n12264, new_n12265, new_n12266, new_n12267, new_n12268, new_n12269,
    new_n12270, new_n12271, new_n12272, new_n12273, new_n12274, new_n12275,
    new_n12276, new_n12277, new_n12278, new_n12279, new_n12280, new_n12281,
    new_n12282, new_n12283, new_n12284, new_n12285, new_n12286, new_n12287,
    new_n12288, new_n12289, new_n12290, new_n12291, new_n12292, new_n12293,
    new_n12294, new_n12295, new_n12296, new_n12297, new_n12298, new_n12299,
    new_n12300, new_n12301, new_n12302, new_n12303, new_n12305, new_n12306,
    new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312,
    new_n12313, new_n12314, new_n12315, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12322, new_n12323, new_n12324,
    new_n12325, new_n12326, new_n12327, new_n12328, new_n12329, new_n12330,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12339,
    new_n12340, new_n12341, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346, new_n12347, new_n12348, new_n12349, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12354, new_n12355, new_n12356, new_n12357,
    new_n12358, new_n12359, new_n12360, new_n12361, new_n12362, new_n12363,
    new_n12364, new_n12365, new_n12366, new_n12367, new_n12368, new_n12369,
    new_n12370, new_n12371, new_n12372, new_n12373, new_n12374, new_n12375,
    new_n12376, new_n12377, new_n12378, new_n12379, new_n12380, new_n12381,
    new_n12382, new_n12383, new_n12384, new_n12385, new_n12386, new_n12387,
    new_n12388, new_n12389, new_n12390, new_n12391, new_n12392, new_n12393,
    new_n12394, new_n12395, new_n12396, new_n12397, new_n12398, new_n12399,
    new_n12400, new_n12401, new_n12402, new_n12403, new_n12404, new_n12405,
    new_n12406, new_n12407, new_n12408, new_n12409, new_n12410, new_n12411,
    new_n12413, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419,
    new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425,
    new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444, new_n12445, new_n12446, new_n12447, new_n12448, new_n12449,
    new_n12450, new_n12451, new_n12452, new_n12453, new_n12454, new_n12455,
    new_n12456, new_n12457, new_n12458, new_n12459, new_n12460, new_n12461,
    new_n12462, new_n12463, new_n12464, new_n12465, new_n12466, new_n12467,
    new_n12468, new_n12469, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495, new_n12496, new_n12497,
    new_n12498, new_n12499, new_n12500, new_n12501, new_n12502, new_n12503,
    new_n12504, new_n12505, new_n12506, new_n12507, new_n12508, new_n12509,
    new_n12510, new_n12511, new_n12512, new_n12513, new_n12514, new_n12515,
    new_n12516, new_n12517, new_n12518, new_n12519, new_n12520, new_n12521,
    new_n12522, new_n12523, new_n12524, new_n12525, new_n12526, new_n12527,
    new_n12528, new_n12529, new_n12530, new_n12531, new_n12532, new_n12533,
    new_n12534, new_n12535, new_n12536, new_n12537, new_n12538, new_n12539,
    new_n12540, new_n12541, new_n12542, new_n12543, new_n12544, new_n12545,
    new_n12546, new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557,
    new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563,
    new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587,
    new_n12588, new_n12589, new_n12590, new_n12591, new_n12592, new_n12593,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607, new_n12608, new_n12609, new_n12610, new_n12611,
    new_n12612, new_n12613, new_n12614, new_n12615, new_n12616, new_n12617,
    new_n12618, new_n12619, new_n12620, new_n12621, new_n12622, new_n12623,
    new_n12624, new_n12625, new_n12626, new_n12627, new_n12628, new_n12629,
    new_n12630, new_n12631, new_n12632, new_n12633, new_n12634, new_n12635,
    new_n12636, new_n12637, new_n12638, new_n12639, new_n12640, new_n12641,
    new_n12642, new_n12643, new_n12644, new_n12645, new_n12646, new_n12647,
    new_n12648, new_n12649, new_n12650, new_n12651, new_n12652, new_n12653,
    new_n12654, new_n12655, new_n12656, new_n12657, new_n12658, new_n12659,
    new_n12660, new_n12661, new_n12662, new_n12663, new_n12664, new_n12665,
    new_n12666, new_n12667, new_n12668, new_n12669, new_n12670, new_n12671,
    new_n12672, new_n12673, new_n12674, new_n12675, new_n12676, new_n12679,
    new_n12680, new_n12681, new_n12682, new_n12683, new_n12684, new_n12685,
    new_n12686, new_n12687, new_n12688, new_n12689, new_n12690, new_n12691,
    new_n12692, new_n12693, new_n12694, new_n12695, new_n12696, new_n12697,
    new_n12698, new_n12699, new_n12700, new_n12701, new_n12702, new_n12703,
    new_n12704, new_n12705, new_n12706, new_n12707, new_n12708, new_n12709,
    new_n12710, new_n12711, new_n12712, new_n12713, new_n12714, new_n12715,
    new_n12716, new_n12718, new_n12719, new_n12720, new_n12721, new_n12722,
    new_n12723, new_n12724, new_n12725, new_n12726, new_n12727, new_n12728,
    new_n12729, new_n12730, new_n12731, new_n12732, new_n12733, new_n12734,
    new_n12735, new_n12736, new_n12737, new_n12738, new_n12739, new_n12740,
    new_n12741, new_n12742, new_n12743, new_n12744, new_n12745, new_n12746,
    new_n12747, new_n12748, new_n12749, new_n12750, new_n12751, new_n12752,
    new_n12753, new_n12754, new_n12755, new_n12756, new_n12757, new_n12758,
    new_n12759, new_n12760, new_n12761, new_n12762, new_n12763, new_n12764,
    new_n12765, new_n12766, new_n12767, new_n12768, new_n12769, new_n12770,
    new_n12771, new_n12772, new_n12773, new_n12774, new_n12775, new_n12776,
    new_n12777, new_n12778, new_n12779, new_n12780, new_n12781, new_n12782,
    new_n12783, new_n12784, new_n12785, new_n12786, new_n12787, new_n12788,
    new_n12789, new_n12790, new_n12791, new_n12792, new_n12793, new_n12794,
    new_n12795, new_n12796, new_n12797, new_n12798, new_n12799, new_n12800,
    new_n12801, new_n12802, new_n12803, new_n12804, new_n12805, new_n12806,
    new_n12807, new_n12808, new_n12809, new_n12810, new_n12811, new_n12812,
    new_n12813, new_n12814, new_n12815, new_n12816, new_n12817, new_n12818,
    new_n12819, new_n12820, new_n12821, new_n12822, new_n12823, new_n12824,
    new_n12825, new_n12826, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925, new_n12926,
    new_n12927, new_n12928, new_n12929, new_n12930, new_n12931, new_n12932,
    new_n12933, new_n12934, new_n12935, new_n12936, new_n12937, new_n12938,
    new_n12939, new_n12940, new_n12941, new_n12942, new_n12943, new_n12944,
    new_n12945, new_n12946, new_n12947, new_n12948, new_n12949, new_n12950,
    new_n12951, new_n12952, new_n12953, new_n12954, new_n12955, new_n12956,
    new_n12957, new_n12958, new_n12959, new_n12960, new_n12961, new_n12962,
    new_n12963, new_n12964, new_n12965, new_n12966, new_n12967, new_n12968,
    new_n12969, new_n12970, new_n12971, new_n12972, new_n12973, new_n12974,
    new_n12975, new_n12976, new_n12977, new_n12978, new_n12979, new_n12980,
    new_n12981, new_n12982, new_n12983, new_n12984, new_n12985, new_n12986,
    new_n12987, new_n12988, new_n12989, new_n12990, new_n12991, new_n12992,
    new_n12993, new_n12994, new_n12995, new_n12996, new_n12997, new_n12998,
    new_n12999, new_n13000, new_n13001, new_n13002, new_n13003, new_n13004,
    new_n13005, new_n13006, new_n13007, new_n13008, new_n13009, new_n13010,
    new_n13011, new_n13012, new_n13013, new_n13014, new_n13015, new_n13016,
    new_n13017, new_n13018, new_n13019, new_n13020, new_n13021, new_n13022,
    new_n13023, new_n13024, new_n13025, new_n13026, new_n13027, new_n13028,
    new_n13029, new_n13030, new_n13031, new_n13032, new_n13033, new_n13034,
    new_n13035, new_n13036, new_n13037, new_n13038, new_n13039, new_n13040,
    new_n13041, new_n13042, new_n13043, new_n13044, new_n13045, new_n13046,
    new_n13047, new_n13048, new_n13049, new_n13050, new_n13053, new_n13054,
    new_n13055, new_n13056, new_n13057, new_n13058, new_n13059, new_n13060,
    new_n13061, new_n13062, new_n13063, new_n13064, new_n13065, new_n13066,
    new_n13067, new_n13068, new_n13069, new_n13070, new_n13071, new_n13072,
    new_n13073, new_n13074, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082, new_n13083, new_n13084,
    new_n13085, new_n13086, new_n13087, new_n13088, new_n13089, new_n13090,
    new_n13091, new_n13092, new_n13093, new_n13094, new_n13095, new_n13096,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116, new_n13117, new_n13118, new_n13119, new_n13120,
    new_n13121, new_n13122, new_n13123, new_n13128, new_n13129, new_n13130,
    new_n13131, new_n13132, new_n13133, new_n13134, new_n13135, new_n13136,
    new_n13137, new_n13138, new_n13139, new_n13140, new_n13141, new_n13142,
    new_n13146, new_n13147, new_n13148, new_n13149, new_n13150, new_n13151,
    new_n13152, new_n13153, new_n13154, new_n13155, new_n13156, new_n13157,
    new_n13158, new_n13159, new_n13160, new_n13161, new_n13162, new_n13163,
    new_n13164, new_n13165, new_n13166, new_n13167, new_n13168, new_n13169,
    new_n13171, new_n13174, new_n13175, new_n13176, new_n13177, new_n13178,
    new_n13179, new_n13180, new_n13181, new_n13182, new_n13183, new_n13184,
    new_n13185, new_n13186, new_n13187, new_n13188, new_n13189, new_n13190,
    new_n13191, new_n13192, new_n13193, new_n13194, new_n13195, new_n13196,
    new_n13197, new_n13198, new_n13199, new_n13200, new_n13201, new_n13202,
    new_n13203, new_n13205, new_n13206, new_n13207, new_n13208, new_n13209,
    new_n13210, new_n13211, new_n13212, new_n13213, new_n13214, new_n13215,
    new_n13216, new_n13217, new_n13218, new_n13219, new_n13220, new_n13221,
    new_n13222, new_n13223, new_n13224, new_n13225, new_n13226, new_n13227,
    new_n13228, new_n13229, new_n13230, new_n13231, new_n13232, new_n13233,
    new_n13234, new_n13235, new_n13236, new_n13237, new_n13238, new_n13241,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263, new_n13264, new_n13265, new_n13266,
    new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272,
    new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13283, new_n13284, new_n13285, new_n13286,
    new_n13287, new_n13288, new_n13289, new_n13290, new_n13291, new_n13292,
    new_n13293, new_n13294, new_n13295, new_n13296, new_n13297, new_n13298,
    new_n13299, new_n13300, new_n13301, new_n13302, new_n13303, new_n13304,
    new_n13305, new_n13306, new_n13307, new_n13308, new_n13309, new_n13310,
    new_n13311, new_n13312, new_n13313, new_n13314, new_n13315, new_n13316,
    new_n13317, new_n13318, new_n13319, new_n13320, new_n13321, new_n13322,
    new_n13323, new_n13324, new_n13325, new_n13326, new_n13327, new_n13328,
    new_n13329, new_n13330, new_n13331, new_n13332, new_n13333, new_n13334,
    new_n13335, new_n13336, new_n13337, new_n13338, new_n13339, new_n13340,
    new_n13341, new_n13342, new_n13343, new_n13344, new_n13345, new_n13346,
    new_n13347, new_n13348, new_n13349, new_n13350, new_n13351, new_n13352,
    new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358,
    new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364,
    new_n13365, new_n13366, new_n13367, new_n13368, new_n13369, new_n13370,
    new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13377,
    new_n13378, new_n13379, new_n13380, new_n13381, new_n13382, new_n13383,
    new_n13384, new_n13385, new_n13386, new_n13387, new_n13388, new_n13389,
    new_n13390, new_n13391, new_n13392, new_n13393, new_n13394, new_n13395,
    new_n13396, new_n13397, new_n13398, new_n13399, new_n13400, new_n13401,
    new_n13402, new_n13403, new_n13404, new_n13405, new_n13406, new_n13407,
    new_n13408, new_n13409, new_n13410, new_n13411, new_n13412, new_n13413,
    new_n13414, new_n13415, new_n13416, new_n13417, new_n13418, new_n13419,
    new_n13420, new_n13421, new_n13422, new_n13423, new_n13424, new_n13425,
    new_n13426, new_n13427, new_n13428, new_n13429, new_n13430, new_n13431,
    new_n13432, new_n13433, new_n13434, new_n13435, new_n13436, new_n13437,
    new_n13438, new_n13439, new_n13440, new_n13441, new_n13442, new_n13443,
    new_n13444, new_n13445, new_n13446, new_n13447, new_n13448, new_n13449,
    new_n13450, new_n13451, new_n13452, new_n13453, new_n13454, new_n13455,
    new_n13456, new_n13457, new_n13458, new_n13459, new_n13460, new_n13461,
    new_n13462, new_n13463, new_n13464, new_n13465, new_n13466, new_n13467,
    new_n13468, new_n13469, new_n13470, new_n13471, new_n13472, new_n13473,
    new_n13474, new_n13475, new_n13476, new_n13477, new_n13478, new_n13479,
    new_n13480, new_n13481, new_n13482, new_n13483, new_n13484, new_n13485,
    new_n13486, new_n13487, new_n13488, new_n13489, new_n13491, new_n13492,
    new_n13493, new_n13494, new_n13495, new_n13496, new_n13497, new_n13498,
    new_n13499, new_n13500, new_n13501, new_n13502, new_n13503, new_n13504,
    new_n13505, new_n13506, new_n13507, new_n13508, new_n13509, new_n13510,
    new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13532, new_n13535, new_n13536,
    new_n13537, new_n13538, new_n13539, new_n13540, new_n13541, new_n13542,
    new_n13543, new_n13544, new_n13545, new_n13546, new_n13547, new_n13549,
    new_n13550, new_n13551, new_n13552, new_n13553, new_n13554, new_n13555,
    new_n13556, new_n13557, new_n13558, new_n13559, new_n13560, new_n13561,
    new_n13562, new_n13563, new_n13564, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591,
    new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597,
    new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603,
    new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609,
    new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615,
    new_n13616, new_n13617, new_n13618, new_n13619, new_n13620, new_n13621,
    new_n13622, new_n13623, new_n13624, new_n13625, new_n13626, new_n13627,
    new_n13628, new_n13629, new_n13630, new_n13631, new_n13632, new_n13633,
    new_n13634, new_n13635, new_n13636, new_n13637, new_n13638, new_n13639,
    new_n13640, new_n13641, new_n13642, new_n13643, new_n13644, new_n13645,
    new_n13646, new_n13647, new_n13648, new_n13649, new_n13650, new_n13651,
    new_n13652, new_n13653, new_n13654, new_n13655, new_n13656, new_n13657,
    new_n13658, new_n13659, new_n13660, new_n13661, new_n13662, new_n13663,
    new_n13664, new_n13665, new_n13666, new_n13667, new_n13668, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677, new_n13678, new_n13679, new_n13680, new_n13681,
    new_n13682, new_n13683, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708, new_n13709, new_n13710, new_n13711,
    new_n13712, new_n13713, new_n13714, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719, new_n13720, new_n13721, new_n13722, new_n13723,
    new_n13724, new_n13725, new_n13726, new_n13729, new_n13730, new_n13731,
    new_n13732, new_n13733, new_n13734, new_n13735, new_n13736, new_n13737,
    new_n13738, new_n13739, new_n13740, new_n13741, new_n13742, new_n13743,
    new_n13744, new_n13745, new_n13746, new_n13747, new_n13748, new_n13749,
    new_n13750, new_n13751, new_n13752, new_n13753, new_n13754, new_n13755,
    new_n13756, new_n13757, new_n13758, new_n13759, new_n13760, new_n13761,
    new_n13762, new_n13763, new_n13764, new_n13765, new_n13766, new_n13767,
    new_n13768, new_n13769, new_n13770, new_n13771, new_n13772, new_n13773,
    new_n13774, new_n13775, new_n13776, new_n13777, new_n13778, new_n13779,
    new_n13780, new_n13781, new_n13782, new_n13783, new_n13784, new_n13785,
    new_n13786, new_n13787, new_n13788, new_n13789, new_n13790, new_n13791,
    new_n13792, new_n13793, new_n13794, new_n13795, new_n13796, new_n13797,
    new_n13798, new_n13799, new_n13800, new_n13801, new_n13802, new_n13803,
    new_n13804, new_n13805, new_n13806, new_n13807, new_n13808, new_n13809,
    new_n13810, new_n13811, new_n13812, new_n13813, new_n13814, new_n13816,
    new_n13817, new_n13818, new_n13819, new_n13820, new_n13821, new_n13822,
    new_n13823, new_n13824, new_n13825, new_n13826, new_n13827, new_n13828,
    new_n13829, new_n13830, new_n13833, new_n13834, new_n13835, new_n13836,
    new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842,
    new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848,
    new_n13849, new_n13850, new_n13851, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860,
    new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866,
    new_n13867, new_n13868, new_n13869, new_n13870, new_n13871, new_n13872,
    new_n13873, new_n13874, new_n13875, new_n13876, new_n13877, new_n13878,
    new_n13879, new_n13880, new_n13881, new_n13882, new_n13883, new_n13884,
    new_n13885, new_n13886, new_n13887, new_n13888, new_n13889, new_n13890,
    new_n13891, new_n13892, new_n13893, new_n13894, new_n13895, new_n13896,
    new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902,
    new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908,
    new_n13909, new_n13910, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14030, new_n14031,
    new_n14032, new_n14033, new_n14034, new_n14035, new_n14036, new_n14037,
    new_n14038, new_n14039, new_n14040, new_n14041, new_n14042, new_n14043,
    new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049,
    new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055,
    new_n14056, new_n14057, new_n14058, new_n14059, new_n14060, new_n14061,
    new_n14062, new_n14063, new_n14064, new_n14065, new_n14066, new_n14067,
    new_n14068, new_n14069, new_n14070, new_n14071, new_n14072, new_n14073,
    new_n14074, new_n14077, new_n14078, new_n14079, new_n14080, new_n14081,
    new_n14082, new_n14083, new_n14084, new_n14085, new_n14086, new_n14087,
    new_n14088, new_n14089, new_n14090, new_n14091, new_n14092, new_n14093,
    new_n14094, new_n14095, new_n14096, new_n14097, new_n14098, new_n14099,
    new_n14100, new_n14101, new_n14102, new_n14103, new_n14104, new_n14105,
    new_n14106, new_n14107, new_n14108, new_n14109, new_n14110, new_n14111,
    new_n14112, new_n14113, new_n14114, new_n14115, new_n14116, new_n14117,
    new_n14118, new_n14119, new_n14120, new_n14121, new_n14122, new_n14123,
    new_n14124, new_n14125, new_n14126, new_n14127, new_n14128, new_n14129,
    new_n14130, new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136, new_n14137, new_n14138, new_n14139, new_n14140, new_n14141,
    new_n14142, new_n14143, new_n14144, new_n14145, new_n14146, new_n14147,
    new_n14148, new_n14149, new_n14150, new_n14151, new_n14152, new_n14153,
    new_n14154, new_n14155, new_n14156, new_n14157, new_n14158, new_n14159,
    new_n14160, new_n14161, new_n14162, new_n14163, new_n14164, new_n14165,
    new_n14166, new_n14167, new_n14168, new_n14169, new_n14170, new_n14171,
    new_n14172, new_n14173, new_n14174, new_n14175, new_n14176, new_n14177,
    new_n14178, new_n14179, new_n14180, new_n14181, new_n14182, new_n14183,
    new_n14184, new_n14185, new_n14186, new_n14187, new_n14188, new_n14189,
    new_n14190, new_n14191, new_n14192, new_n14193, new_n14194, new_n14195,
    new_n14196, new_n14197, new_n14198, new_n14199, new_n14200, new_n14201,
    new_n14202, new_n14203, new_n14204, new_n14205, new_n14206, new_n14207,
    new_n14208, new_n14209, new_n14210, new_n14211, new_n14212, new_n14213,
    new_n14215, new_n14216, new_n14217, new_n14218, new_n14219, new_n14221,
    new_n14222, new_n14223, new_n14224, new_n14225, new_n14226, new_n14227,
    new_n14228, new_n14229, new_n14230, new_n14231, new_n14232, new_n14233,
    new_n14234, new_n14235, new_n14236, new_n14237, new_n14238, new_n14239,
    new_n14240, new_n14241, new_n14242, new_n14243, new_n14244, new_n14245,
    new_n14246, new_n14247, new_n14248, new_n14249, new_n14250, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258,
    new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264,
    new_n14265, new_n14266, new_n14267, new_n14268, new_n14269, new_n14270,
    new_n14271, new_n14272, new_n14273, new_n14274, new_n14275, new_n14276,
    new_n14277, new_n14278, new_n14279, new_n14280, new_n14281, new_n14282,
    new_n14283, new_n14284, new_n14285, new_n14286, new_n14287, new_n14288,
    new_n14289, new_n14290, new_n14291, new_n14292, new_n14293, new_n14294,
    new_n14295, new_n14296, new_n14297, new_n14298, new_n14299, new_n14300,
    new_n14301, new_n14302, new_n14303, new_n14304, new_n14305, new_n14306,
    new_n14307, new_n14308, new_n14309, new_n14310, new_n14311, new_n14312,
    new_n14313, new_n14314, new_n14315, new_n14316, new_n14317, new_n14318,
    new_n14319, new_n14320, new_n14321, new_n14322, new_n14323, new_n14324,
    new_n14325, new_n14326, new_n14327, new_n14328, new_n14329, new_n14330,
    new_n14331, new_n14332, new_n14333, new_n14334, new_n14335, new_n14336,
    new_n14337, new_n14338, new_n14339, new_n14340, new_n14341, new_n14342,
    new_n14343, new_n14344, new_n14345, new_n14346, new_n14347, new_n14348,
    new_n14349, new_n14350, new_n14351, new_n14352, new_n14353, new_n14354,
    new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360,
    new_n14361, new_n14362, new_n14363, new_n14364, new_n14365, new_n14366,
    new_n14367, new_n14368, new_n14369, new_n14370, new_n14371, new_n14372,
    new_n14373, new_n14374, new_n14375, new_n14376, new_n14377, new_n14378,
    new_n14379, new_n14380, new_n14381, new_n14382, new_n14383, new_n14384,
    new_n14385, new_n14386, new_n14387, new_n14388, new_n14389, new_n14390,
    new_n14391, new_n14392, new_n14393, new_n14394, new_n14395, new_n14396,
    new_n14397, new_n14398, new_n14399, new_n14400, new_n14401, new_n14402,
    new_n14403, new_n14404, new_n14405, new_n14406, new_n14407, new_n14408,
    new_n14409, new_n14410, new_n14411, new_n14412, new_n14413, new_n14414,
    new_n14415, new_n14416, new_n14417, new_n14418, new_n14419, new_n14420,
    new_n14421, new_n14422, new_n14423, new_n14424, new_n14425, new_n14426,
    new_n14427, new_n14428, new_n14429, new_n14430, new_n14431, new_n14432,
    new_n14434, new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440, new_n14441, new_n14442, new_n14443, new_n14444, new_n14445,
    new_n14446, new_n14447, new_n14448, new_n14449, new_n14450, new_n14451,
    new_n14452, new_n14453, new_n14454, new_n14455, new_n14456, new_n14457,
    new_n14458, new_n14459, new_n14460, new_n14461, new_n14462, new_n14463,
    new_n14464, new_n14465, new_n14466, new_n14467, new_n14468, new_n14469,
    new_n14470, new_n14471, new_n14472, new_n14473, new_n14474, new_n14475,
    new_n14477, new_n14478, new_n14480, new_n14481, new_n14482, new_n14483,
    new_n14484, new_n14485, new_n14486, new_n14487, new_n14488, new_n14489,
    new_n14490, new_n14491, new_n14492, new_n14493, new_n14494, new_n14495,
    new_n14496, new_n14497, new_n14498, new_n14499, new_n14500, new_n14501,
    new_n14502, new_n14503, new_n14504, new_n14505, new_n14506, new_n14507,
    new_n14508, new_n14509, new_n14510, new_n14511, new_n14512, new_n14513,
    new_n14514, new_n14515, new_n14516, new_n14517, new_n14518, new_n14519,
    new_n14520, new_n14521, new_n14522, new_n14523, new_n14524, new_n14525,
    new_n14526, new_n14527, new_n14528, new_n14529, new_n14530, new_n14531,
    new_n14532, new_n14533, new_n14534, new_n14535, new_n14536, new_n14537,
    new_n14538, new_n14539, new_n14540, new_n14541, new_n14542, new_n14543,
    new_n14544, new_n14545, new_n14546, new_n14547, new_n14548, new_n14549,
    new_n14550, new_n14551, new_n14552, new_n14553, new_n14554, new_n14555,
    new_n14556, new_n14557, new_n14558, new_n14559, new_n14560, new_n14561,
    new_n14562, new_n14563, new_n14564, new_n14565, new_n14566, new_n14567,
    new_n14568, new_n14569, new_n14570, new_n14571, new_n14572, new_n14573,
    new_n14574, new_n14575, new_n14576, new_n14577, new_n14578, new_n14579,
    new_n14580, new_n14581, new_n14582, new_n14583, new_n14584, new_n14585,
    new_n14586, new_n14587, new_n14588, new_n14589, new_n14590, new_n14591,
    new_n14592, new_n14593, new_n14594, new_n14595, new_n14596, new_n14597,
    new_n14598, new_n14599, new_n14600, new_n14601, new_n14602, new_n14603,
    new_n14604, new_n14605, new_n14606, new_n14607, new_n14608, new_n14609,
    new_n14610, new_n14611, new_n14612, new_n14613, new_n14614, new_n14615,
    new_n14616, new_n14617, new_n14618, new_n14619, new_n14620, new_n14621,
    new_n14622, new_n14623, new_n14624, new_n14625, new_n14626, new_n14627,
    new_n14628, new_n14629, new_n14630, new_n14631, new_n14632, new_n14634,
    new_n14635, new_n14636, new_n14637, new_n14638, new_n14639, new_n14640,
    new_n14641, new_n14642, new_n14643, new_n14644, new_n14645, new_n14646,
    new_n14647, new_n14648, new_n14649, new_n14650, new_n14651, new_n14652,
    new_n14653, new_n14654, new_n14655, new_n14656, new_n14657, new_n14658,
    new_n14659, new_n14660, new_n14661, new_n14662, new_n14663, new_n14664,
    new_n14665, new_n14666, new_n14667, new_n14668, new_n14669, new_n14670,
    new_n14671, new_n14672, new_n14673, new_n14674, new_n14675, new_n14676,
    new_n14677, new_n14678, new_n14679, new_n14680, new_n14681, new_n14682,
    new_n14683, new_n14684, new_n14685, new_n14686, new_n14687, new_n14688,
    new_n14689, new_n14690, new_n14691, new_n14692, new_n14693, new_n14694,
    new_n14695, new_n14696, new_n14697, new_n14698, new_n14699, new_n14700,
    new_n14701, new_n14702, new_n14703, new_n14704, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724,
    new_n14725, new_n14726, new_n14727, new_n14728, new_n14729, new_n14730,
    new_n14731, new_n14732, new_n14733, new_n14734, new_n14735, new_n14736,
    new_n14737, new_n14738, new_n14739, new_n14740, new_n14741, new_n14742,
    new_n14743, new_n14744, new_n14745, new_n14746, new_n14747, new_n14748,
    new_n14749, new_n14750, new_n14751, new_n14752, new_n14753, new_n14754,
    new_n14755, new_n14756, new_n14757, new_n14758, new_n14759, new_n14760,
    new_n14762, new_n14763, new_n14764, new_n14765, new_n14766, new_n14767,
    new_n14768, new_n14769, new_n14770, new_n14771, new_n14772, new_n14773,
    new_n14774, new_n14775, new_n14776, new_n14777, new_n14778, new_n14779,
    new_n14780, new_n14781, new_n14782, new_n14783, new_n14784, new_n14785,
    new_n14786, new_n14787, new_n14788, new_n14789, new_n14790, new_n14791,
    new_n14792, new_n14793, new_n14794, new_n14795, new_n14796, new_n14797,
    new_n14798, new_n14799, new_n14800, new_n14801, new_n14802, new_n14803,
    new_n14804, new_n14805, new_n14806, new_n14807, new_n14808, new_n14809,
    new_n14810, new_n14812, new_n14813, new_n14814, new_n14815, new_n14816,
    new_n14817, new_n14818, new_n14819, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826, new_n14827, new_n14828,
    new_n14829, new_n14830, new_n14831, new_n14832, new_n14833, new_n14834,
    new_n14835, new_n14836, new_n14837, new_n14838, new_n14839, new_n14840,
    new_n14841, new_n14842, new_n14843, new_n14844, new_n14845, new_n14846,
    new_n14847, new_n14848, new_n14849, new_n14850, new_n14851, new_n14852,
    new_n14853, new_n14854, new_n14855, new_n14856, new_n14857, new_n14858,
    new_n14859, new_n14860, new_n14861, new_n14862, new_n14863, new_n14864,
    new_n14865, new_n14866, new_n14867, new_n14868, new_n14869, new_n14870,
    new_n14871, new_n14872, new_n14873, new_n14874, new_n14875, new_n14876,
    new_n14877, new_n14878, new_n14879, new_n14880, new_n14881, new_n14882,
    new_n14883, new_n14884, new_n14885, new_n14886, new_n14887, new_n14888,
    new_n14889, new_n14890, new_n14891, new_n14892, new_n14893, new_n14894,
    new_n14895, new_n14896, new_n14897, new_n14898, new_n14899, new_n14900,
    new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906,
    new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912,
    new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918,
    new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924,
    new_n14925, new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931, new_n14932, new_n14934, new_n14935, new_n14936, new_n14937,
    new_n14938, new_n14939, new_n14940, new_n14941, new_n14942, new_n14943,
    new_n14944, new_n14945, new_n14946, new_n14947, new_n14948, new_n14949,
    new_n14950, new_n14951, new_n14952, new_n14953, new_n14954, new_n14955,
    new_n14956, new_n14957, new_n14958, new_n14959, new_n14960, new_n14961,
    new_n14962, new_n14963, new_n14964, new_n14965, new_n14966, new_n14967,
    new_n14968, new_n14969, new_n14970, new_n14971, new_n14972, new_n14973,
    new_n14974, new_n14975, new_n14976, new_n14977, new_n14978, new_n14979,
    new_n14980, new_n14981, new_n14982, new_n14983, new_n14984, new_n14985,
    new_n14986, new_n14987, new_n14988, new_n14989, new_n14990, new_n14991,
    new_n14994, new_n14995, new_n14996, new_n14997, new_n14998, new_n14999,
    new_n15000, new_n15001, new_n15002, new_n15003, new_n15004, new_n15005,
    new_n15006, new_n15007, new_n15008, new_n15009, new_n15010, new_n15011,
    new_n15012, new_n15013, new_n15014, new_n15015, new_n15016, new_n15017,
    new_n15018, new_n15019, new_n15020, new_n15021, new_n15022, new_n15023,
    new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029,
    new_n15030, new_n15031, new_n15032, new_n15033, new_n15034, new_n15035,
    new_n15036, new_n15037, new_n15038, new_n15039, new_n15040, new_n15041,
    new_n15042, new_n15043, new_n15044, new_n15045, new_n15046, new_n15047,
    new_n15048, new_n15049, new_n15050, new_n15051, new_n15052, new_n15053,
    new_n15054, new_n15055, new_n15056, new_n15057, new_n15058, new_n15059,
    new_n15060, new_n15061, new_n15062, new_n15063, new_n15064, new_n15065,
    new_n15066, new_n15067, new_n15068, new_n15069, new_n15070, new_n15071,
    new_n15072, new_n15073, new_n15074, new_n15075, new_n15076, new_n15077,
    new_n15078, new_n15079, new_n15080, new_n15081, new_n15082, new_n15083,
    new_n15084, new_n15085, new_n15086, new_n15087, new_n15088, new_n15089,
    new_n15090, new_n15091, new_n15092, new_n15093, new_n15094, new_n15095,
    new_n15096, new_n15097, new_n15098, new_n15099, new_n15100, new_n15101,
    new_n15102, new_n15103, new_n15104, new_n15105, new_n15106, new_n15107,
    new_n15109, new_n15110, new_n15111, new_n15112, new_n15113, new_n15114,
    new_n15115, new_n15116, new_n15117, new_n15118, new_n15119, new_n15120,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128, new_n15129, new_n15130, new_n15131, new_n15132,
    new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138,
    new_n15139, new_n15140, new_n15141, new_n15142, new_n15143, new_n15144,
    new_n15145, new_n15146, new_n15147, new_n15148, new_n15149, new_n15150,
    new_n15151, new_n15152, new_n15153, new_n15154, new_n15155, new_n15156,
    new_n15157, new_n15158, new_n15159, new_n15160, new_n15161, new_n15162,
    new_n15163, new_n15164, new_n15165, new_n15166, new_n15167, new_n15168,
    new_n15169, new_n15170, new_n15171, new_n15172, new_n15173, new_n15174,
    new_n15175, new_n15176, new_n15177, new_n15178, new_n15179, new_n15180,
    new_n15181, new_n15182, new_n15183, new_n15184, new_n15185, new_n15186,
    new_n15187, new_n15188, new_n15189, new_n15190, new_n15191, new_n15192,
    new_n15193, new_n15194, new_n15195, new_n15196, new_n15197, new_n15198,
    new_n15199, new_n15200, new_n15201, new_n15202, new_n15203, new_n15204,
    new_n15205, new_n15206, new_n15207, new_n15208, new_n15209, new_n15210,
    new_n15211, new_n15212, new_n15213, new_n15214, new_n15215, new_n15216,
    new_n15217, new_n15220, new_n15226, new_n15228, new_n15229, new_n15230,
    new_n15231, new_n15232, new_n15233, new_n15234, new_n15235, new_n15236,
    new_n15237, new_n15238, new_n15239, new_n15240, new_n15241, new_n15242,
    new_n15243, new_n15244, new_n15245, new_n15246, new_n15247, new_n15248,
    new_n15249, new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15256, new_n15258, new_n15259, new_n15260, new_n15261, new_n15262,
    new_n15263, new_n15264, new_n15265, new_n15266, new_n15267, new_n15268,
    new_n15269, new_n15270, new_n15271, new_n15272, new_n15273, new_n15274,
    new_n15275, new_n15276, new_n15277, new_n15278, new_n15279, new_n15280,
    new_n15281, new_n15282, new_n15283, new_n15284, new_n15285, new_n15286,
    new_n15287, new_n15288, new_n15289, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300, new_n15301, new_n15302, new_n15303, new_n15304,
    new_n15305, new_n15306, new_n15307, new_n15308, new_n15309, new_n15310,
    new_n15311, new_n15312, new_n15313, new_n15314, new_n15315, new_n15316,
    new_n15317, new_n15318, new_n15319, new_n15320, new_n15325, new_n15326,
    new_n15327, new_n15328, new_n15329, new_n15330, new_n15331, new_n15332,
    new_n15333, new_n15334, new_n15335, new_n15336, new_n15337, new_n15338,
    new_n15339, new_n15340, new_n15341, new_n15342, new_n15343, new_n15344,
    new_n15345, new_n15346, new_n15347, new_n15348, new_n15349, new_n15350,
    new_n15351, new_n15352, new_n15353, new_n15354, new_n15355, new_n15356,
    new_n15357, new_n15358, new_n15359, new_n15360, new_n15361, new_n15362,
    new_n15363, new_n15364, new_n15365, new_n15366, new_n15367, new_n15368,
    new_n15369, new_n15370, new_n15371, new_n15372, new_n15373, new_n15374,
    new_n15375, new_n15376, new_n15377, new_n15378, new_n15379, new_n15380,
    new_n15381, new_n15382, new_n15383, new_n15384, new_n15385, new_n15386,
    new_n15387, new_n15388, new_n15389, new_n15390, new_n15391, new_n15392,
    new_n15393, new_n15394, new_n15395, new_n15396, new_n15397, new_n15398,
    new_n15399, new_n15400, new_n15401, new_n15402, new_n15403, new_n15404,
    new_n15405, new_n15406, new_n15407, new_n15408, new_n15409, new_n15410,
    new_n15411, new_n15412, new_n15413, new_n15414, new_n15415, new_n15416,
    new_n15417, new_n15418, new_n15419, new_n15420, new_n15421, new_n15422,
    new_n15423, new_n15424, new_n15425, new_n15426, new_n15427, new_n15428,
    new_n15429, new_n15430, new_n15433, new_n15434, new_n15435, new_n15436,
    new_n15437, new_n15438, new_n15439, new_n15440, new_n15441, new_n15442,
    new_n15443, new_n15444, new_n15445, new_n15446, new_n15447, new_n15448,
    new_n15449, new_n15450, new_n15451, new_n15452, new_n15453, new_n15454,
    new_n15455, new_n15456, new_n15457, new_n15458, new_n15459, new_n15460,
    new_n15461, new_n15462, new_n15463, new_n15464, new_n15465, new_n15466,
    new_n15467, new_n15468, new_n15469, new_n15470, new_n15471, new_n15472,
    new_n15473, new_n15474, new_n15475, new_n15476, new_n15477, new_n15478,
    new_n15479, new_n15480, new_n15481, new_n15482, new_n15483, new_n15484,
    new_n15485, new_n15486, new_n15487, new_n15488, new_n15489, new_n15491,
    new_n15492, new_n15493, new_n15494, new_n15495, new_n15496, new_n15497,
    new_n15498, new_n15499, new_n15500, new_n15501, new_n15502, new_n15503,
    new_n15504, new_n15505, new_n15506, new_n15507, new_n15508, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15527, new_n15528, new_n15529,
    new_n15530, new_n15531, new_n15532, new_n15533, new_n15534, new_n15535,
    new_n15536, new_n15537, new_n15538, new_n15539, new_n15540, new_n15541,
    new_n15542, new_n15543, new_n15544, new_n15545, new_n15546, new_n15547,
    new_n15548, new_n15549, new_n15550, new_n15551, new_n15552, new_n15553,
    new_n15554, new_n15555, new_n15556, new_n15557, new_n15558, new_n15559,
    new_n15560, new_n15561, new_n15562, new_n15563, new_n15564, new_n15565,
    new_n15566, new_n15567, new_n15568, new_n15569, new_n15570, new_n15571,
    new_n15572, new_n15573, new_n15574, new_n15575, new_n15576, new_n15577,
    new_n15578, new_n15579, new_n15581, new_n15582, new_n15583, new_n15584,
    new_n15585, new_n15586, new_n15587, new_n15588, new_n15589, new_n15590,
    new_n15591, new_n15592, new_n15593, new_n15594, new_n15595, new_n15596,
    new_n15597, new_n15598, new_n15599, new_n15600, new_n15601, new_n15602,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613, new_n15614,
    new_n15615, new_n15616, new_n15617, new_n15618, new_n15620, new_n15621,
    new_n15622, new_n15623, new_n15624, new_n15625, new_n15626, new_n15627,
    new_n15628, new_n15629, new_n15630, new_n15631, new_n15632, new_n15633,
    new_n15634, new_n15635, new_n15636, new_n15637, new_n15638, new_n15639,
    new_n15640, new_n15641, new_n15642, new_n15643, new_n15644, new_n15645,
    new_n15646, new_n15647, new_n15648, new_n15649, new_n15650, new_n15651,
    new_n15652, new_n15653, new_n15654, new_n15655, new_n15656, new_n15657,
    new_n15658, new_n15659, new_n15660, new_n15661, new_n15662, new_n15663,
    new_n15664, new_n15665, new_n15666, new_n15667, new_n15668, new_n15669,
    new_n15670, new_n15671, new_n15672, new_n15673, new_n15674, new_n15675,
    new_n15676, new_n15677, new_n15678, new_n15679, new_n15680, new_n15681,
    new_n15682, new_n15683, new_n15684, new_n15685, new_n15686, new_n15687,
    new_n15688, new_n15689, new_n15690, new_n15691, new_n15692, new_n15693,
    new_n15694, new_n15695, new_n15696, new_n15697, new_n15698, new_n15699,
    new_n15700, new_n15701, new_n15702, new_n15703, new_n15704, new_n15705,
    new_n15706, new_n15707, new_n15708, new_n15709, new_n15710, new_n15711,
    new_n15712, new_n15713, new_n15714, new_n15715, new_n15716, new_n15717,
    new_n15718, new_n15719, new_n15720, new_n15721, new_n15722, new_n15723,
    new_n15724, new_n15725, new_n15726, new_n15727, new_n15728, new_n15729,
    new_n15730, new_n15731, new_n15732, new_n15733, new_n15734, new_n15735,
    new_n15736, new_n15737, new_n15738, new_n15739, new_n15740, new_n15741,
    new_n15742, new_n15743, new_n15744, new_n15745, new_n15746, new_n15747,
    new_n15748, new_n15749, new_n15750, new_n15751, new_n15752, new_n15753,
    new_n15754, new_n15755, new_n15756, new_n15757, new_n15758, new_n15759,
    new_n15760, new_n15761, new_n15762, new_n15763, new_n15764, new_n15765,
    new_n15766, new_n15767, new_n15768, new_n15769, new_n15770, new_n15771,
    new_n15772, new_n15773, new_n15774, new_n15775, new_n15776, new_n15777,
    new_n15778, new_n15779, new_n15780, new_n15781, new_n15782, new_n15783,
    new_n15784, new_n15785, new_n15786, new_n15787, new_n15788, new_n15789,
    new_n15790, new_n15791, new_n15792, new_n15793, new_n15794, new_n15795,
    new_n15796, new_n15797, new_n15798, new_n15799, new_n15800, new_n15801,
    new_n15802, new_n15803, new_n15804, new_n15805, new_n15806, new_n15807,
    new_n15808, new_n15809, new_n15810, new_n15811, new_n15812, new_n15813,
    new_n15814, new_n15815, new_n15816, new_n15817, new_n15818, new_n15819,
    new_n15820, new_n15821, new_n15822, new_n15823, new_n15828, new_n15829,
    new_n15830, new_n15831, new_n15832, new_n15833, new_n15834, new_n15835,
    new_n15836, new_n15837, new_n15838, new_n15839, new_n15840, new_n15841,
    new_n15844, new_n15845, new_n15846, new_n15847, new_n15848, new_n15849,
    new_n15850, new_n15851, new_n15852, new_n15853, new_n15854, new_n15855,
    new_n15856, new_n15857, new_n15858, new_n15859, new_n15860, new_n15861,
    new_n15862, new_n15863, new_n15864, new_n15865, new_n15866, new_n15867,
    new_n15868, new_n15869, new_n15870, new_n15871, new_n15872, new_n15873,
    new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879,
    new_n15880, new_n15881, new_n15882, new_n15883, new_n15884, new_n15885,
    new_n15886, new_n15887, new_n15888, new_n15889, new_n15890, new_n15891,
    new_n15892, new_n15893, new_n15894, new_n15895, new_n15896, new_n15897,
    new_n15898, new_n15899, new_n15900, new_n15901, new_n15902, new_n15903,
    new_n15904, new_n15905, new_n15906, new_n15907, new_n15908, new_n15909,
    new_n15910, new_n15911, new_n15912, new_n15913, new_n15914, new_n15915,
    new_n15916, new_n15917, new_n15918, new_n15919, new_n15920, new_n15921,
    new_n15922, new_n15923, new_n15924, new_n15925, new_n15926, new_n15927,
    new_n15928, new_n15929, new_n15930, new_n15931, new_n15932, new_n15933,
    new_n15934, new_n15936, new_n15937, new_n15939, new_n15940, new_n15941,
    new_n15942, new_n15943, new_n15944, new_n15945, new_n15946, new_n15947,
    new_n15948, new_n15949, new_n15950, new_n15951, new_n15952, new_n15953,
    new_n15954, new_n15955, new_n15956, new_n15957, new_n15958, new_n15959,
    new_n15960, new_n15961, new_n15962, new_n15963, new_n15964, new_n15965,
    new_n15966, new_n15967, new_n15968, new_n15969, new_n15970, new_n15971,
    new_n15972, new_n15973, new_n15974, new_n15975, new_n15976, new_n15978,
    new_n15979, new_n15980, new_n15981, new_n15982, new_n15983, new_n15984,
    new_n15985, new_n15986, new_n15987, new_n15988, new_n15989, new_n15990,
    new_n15991, new_n15992, new_n15993, new_n15994, new_n15995, new_n15996,
    new_n15997, new_n15998, new_n15999, new_n16000, new_n16001, new_n16003,
    new_n16005, new_n16006, new_n16007, new_n16008, new_n16009, new_n16010,
    new_n16011, new_n16012, new_n16013, new_n16014, new_n16015, new_n16016,
    new_n16017, new_n16018, new_n16019, new_n16020, new_n16021, new_n16022,
    new_n16023, new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029, new_n16030, new_n16031, new_n16032, new_n16033, new_n16034,
    new_n16035, new_n16036, new_n16037, new_n16038, new_n16039, new_n16040,
    new_n16041, new_n16042, new_n16044, new_n16045, new_n16046, new_n16047,
    new_n16048, new_n16049, new_n16050, new_n16051, new_n16052, new_n16053,
    new_n16054, new_n16055, new_n16056, new_n16057, new_n16058, new_n16059,
    new_n16060, new_n16061, new_n16062, new_n16063, new_n16064, new_n16065,
    new_n16066, new_n16067, new_n16068, new_n16069, new_n16070, new_n16071,
    new_n16072, new_n16073, new_n16074, new_n16075, new_n16076, new_n16077,
    new_n16078, new_n16079, new_n16080, new_n16081, new_n16082, new_n16083,
    new_n16084, new_n16085, new_n16086, new_n16087, new_n16088, new_n16089,
    new_n16090, new_n16091, new_n16092, new_n16093, new_n16094, new_n16095,
    new_n16096, new_n16097, new_n16098, new_n16099, new_n16100, new_n16101,
    new_n16102, new_n16103, new_n16104, new_n16105, new_n16106, new_n16107,
    new_n16108, new_n16109, new_n16110, new_n16111, new_n16112, new_n16113,
    new_n16114, new_n16115, new_n16116, new_n16117, new_n16118, new_n16119,
    new_n16120, new_n16121, new_n16122, new_n16123, new_n16124, new_n16125,
    new_n16126, new_n16127, new_n16128, new_n16129, new_n16130, new_n16131,
    new_n16132, new_n16133, new_n16134, new_n16135, new_n16136, new_n16137,
    new_n16138, new_n16139, new_n16140, new_n16141, new_n16142, new_n16143,
    new_n16144, new_n16145, new_n16146, new_n16147, new_n16148, new_n16149,
    new_n16150, new_n16151, new_n16152, new_n16153, new_n16154, new_n16155,
    new_n16156, new_n16157, new_n16158, new_n16159, new_n16160, new_n16161,
    new_n16162, new_n16163, new_n16164, new_n16165, new_n16166, new_n16167,
    new_n16168, new_n16169, new_n16170, new_n16171, new_n16172, new_n16173,
    new_n16174, new_n16175, new_n16176, new_n16177, new_n16178, new_n16179,
    new_n16180, new_n16181, new_n16182, new_n16183, new_n16184, new_n16185,
    new_n16186, new_n16187, new_n16188, new_n16189, new_n16190, new_n16191,
    new_n16192, new_n16193, new_n16194, new_n16195, new_n16196, new_n16197,
    new_n16198, new_n16199, new_n16200, new_n16201, new_n16202, new_n16203,
    new_n16204, new_n16205, new_n16206, new_n16207, new_n16208, new_n16209,
    new_n16210, new_n16211, new_n16212, new_n16213, new_n16214, new_n16215,
    new_n16216, new_n16217, new_n16218, new_n16219, new_n16220, new_n16221,
    new_n16222, new_n16223, new_n16224, new_n16225, new_n16226, new_n16227,
    new_n16228, new_n16229, new_n16230, new_n16231, new_n16233, new_n16234,
    new_n16235, new_n16236, new_n16237, new_n16238, new_n16239, new_n16240,
    new_n16241, new_n16242, new_n16243, new_n16244, new_n16245, new_n16246,
    new_n16247, new_n16248, new_n16249, new_n16250, new_n16251, new_n16252,
    new_n16253, new_n16254, new_n16255, new_n16256, new_n16257, new_n16258,
    new_n16259, new_n16260, new_n16261, new_n16262, new_n16263, new_n16264,
    new_n16265, new_n16266, new_n16267, new_n16268, new_n16269, new_n16270,
    new_n16271, new_n16272, new_n16273, new_n16274, new_n16275, new_n16276,
    new_n16277, new_n16278, new_n16279, new_n16280, new_n16281, new_n16282,
    new_n16283, new_n16284, new_n16285, new_n16286, new_n16287, new_n16288,
    new_n16289, new_n16290, new_n16291, new_n16292, new_n16293, new_n16294,
    new_n16295, new_n16296, new_n16297, new_n16298, new_n16299, new_n16300,
    new_n16302, new_n16303, new_n16304, new_n16305, new_n16306, new_n16307,
    new_n16308, new_n16309, new_n16310, new_n16311, new_n16312, new_n16313,
    new_n16314, new_n16315, new_n16316, new_n16317, new_n16318, new_n16319,
    new_n16320, new_n16321, new_n16322, new_n16323, new_n16324, new_n16325,
    new_n16326, new_n16327, new_n16328, new_n16329, new_n16330, new_n16331,
    new_n16332, new_n16333, new_n16334, new_n16335, new_n16336, new_n16337,
    new_n16338, new_n16339, new_n16340, new_n16341, new_n16342, new_n16343,
    new_n16344, new_n16345, new_n16346, new_n16347, new_n16348, new_n16349,
    new_n16350, new_n16351, new_n16353, new_n16355, new_n16356, new_n16357,
    new_n16358, new_n16359, new_n16360, new_n16361, new_n16362, new_n16363,
    new_n16364, new_n16365, new_n16366, new_n16367, new_n16368, new_n16369,
    new_n16370, new_n16371, new_n16372, new_n16373, new_n16374, new_n16375,
    new_n16376, new_n16377, new_n16378, new_n16379, new_n16380, new_n16381,
    new_n16382, new_n16383, new_n16384, new_n16385, new_n16386, new_n16387,
    new_n16388, new_n16389, new_n16390, new_n16391, new_n16392, new_n16393,
    new_n16394, new_n16395, new_n16396, new_n16397, new_n16398, new_n16399,
    new_n16400, new_n16401, new_n16402, new_n16403, new_n16404, new_n16405,
    new_n16406, new_n16407, new_n16408, new_n16409, new_n16410, new_n16411,
    new_n16412, new_n16413, new_n16414, new_n16415, new_n16416, new_n16417,
    new_n16418, new_n16419, new_n16420, new_n16421, new_n16422, new_n16423,
    new_n16424, new_n16425, new_n16426, new_n16427, new_n16428, new_n16429,
    new_n16430, new_n16431, new_n16432, new_n16433, new_n16434, new_n16435,
    new_n16436, new_n16437, new_n16438, new_n16439, new_n16440, new_n16441,
    new_n16442, new_n16443, new_n16445, new_n16446, new_n16447, new_n16448,
    new_n16449, new_n16450, new_n16451, new_n16452, new_n16453, new_n16454,
    new_n16455, new_n16456, new_n16457, new_n16458, new_n16459, new_n16460,
    new_n16461, new_n16462, new_n16463, new_n16464, new_n16465, new_n16466,
    new_n16467, new_n16468, new_n16469, new_n16470, new_n16471, new_n16472,
    new_n16473, new_n16474, new_n16475, new_n16476, new_n16477, new_n16478,
    new_n16479, new_n16480, new_n16481, new_n16482, new_n16483, new_n16484,
    new_n16485, new_n16486, new_n16487, new_n16488, new_n16489, new_n16490,
    new_n16491, new_n16492, new_n16493, new_n16494, new_n16495, new_n16496,
    new_n16497, new_n16499, new_n16500, new_n16501, new_n16502, new_n16503,
    new_n16504, new_n16505, new_n16506, new_n16507, new_n16508, new_n16509,
    new_n16510, new_n16511, new_n16512, new_n16513, new_n16514, new_n16515,
    new_n16516, new_n16517, new_n16518, new_n16519, new_n16522, new_n16523,
    new_n16524, new_n16525, new_n16526, new_n16527, new_n16528, new_n16529,
    new_n16530, new_n16531, new_n16532, new_n16533, new_n16534, new_n16535,
    new_n16536, new_n16537, new_n16538, new_n16539, new_n16540, new_n16541,
    new_n16542, new_n16543, new_n16544, new_n16545, new_n16546, new_n16547,
    new_n16548, new_n16549, new_n16550, new_n16551, new_n16552, new_n16553,
    new_n16554, new_n16555, new_n16556, new_n16557, new_n16558, new_n16559,
    new_n16560, new_n16561, new_n16562, new_n16563, new_n16564, new_n16565,
    new_n16566, new_n16567, new_n16568, new_n16569, new_n16570, new_n16571,
    new_n16572, new_n16573, new_n16574, new_n16575, new_n16576, new_n16577,
    new_n16578, new_n16579, new_n16580, new_n16581, new_n16582, new_n16583,
    new_n16584, new_n16585, new_n16586, new_n16587, new_n16588, new_n16589,
    new_n16591, new_n16592, new_n16593, new_n16594, new_n16598, new_n16599,
    new_n16600, new_n16601, new_n16602, new_n16603, new_n16604, new_n16605,
    new_n16606, new_n16607, new_n16611, new_n16612, new_n16613, new_n16614,
    new_n16615, new_n16616, new_n16617, new_n16618, new_n16619, new_n16620,
    new_n16621, new_n16622, new_n16623, new_n16624, new_n16625, new_n16626,
    new_n16627, new_n16628, new_n16629, new_n16630, new_n16631, new_n16632,
    new_n16633, new_n16634, new_n16635, new_n16636, new_n16637, new_n16638,
    new_n16639, new_n16640, new_n16641, new_n16642, new_n16643, new_n16644,
    new_n16645, new_n16646, new_n16649, new_n16650, new_n16651, new_n16652,
    new_n16653, new_n16654, new_n16655, new_n16656, new_n16657, new_n16658,
    new_n16659, new_n16660, new_n16661, new_n16662, new_n16663, new_n16664,
    new_n16665, new_n16666, new_n16667, new_n16668, new_n16669, new_n16670,
    new_n16671, new_n16672, new_n16673, new_n16674, new_n16675, new_n16676,
    new_n16677, new_n16678, new_n16679, new_n16680, new_n16681, new_n16682,
    new_n16683, new_n16684, new_n16685, new_n16686, new_n16687, new_n16688,
    new_n16689, new_n16690, new_n16691, new_n16692, new_n16693, new_n16694,
    new_n16695, new_n16696, new_n16697, new_n16698, new_n16699, new_n16700,
    new_n16701, new_n16702, new_n16703, new_n16704, new_n16705, new_n16706,
    new_n16707, new_n16708, new_n16709, new_n16710, new_n16711, new_n16712,
    new_n16713, new_n16714, new_n16715, new_n16716, new_n16717, new_n16718,
    new_n16719, new_n16720, new_n16721, new_n16722, new_n16723, new_n16724,
    new_n16725, new_n16726, new_n16727, new_n16728, new_n16729, new_n16730,
    new_n16731, new_n16732, new_n16733, new_n16734, new_n16735, new_n16736,
    new_n16737, new_n16738, new_n16739, new_n16740, new_n16741, new_n16742,
    new_n16743, new_n16744, new_n16745, new_n16746, new_n16747, new_n16748,
    new_n16749, new_n16750, new_n16751, new_n16752, new_n16753, new_n16754,
    new_n16755, new_n16756, new_n16757, new_n16758, new_n16759, new_n16762,
    new_n16763, new_n16764, new_n16765, new_n16766, new_n16767, new_n16768,
    new_n16769, new_n16770, new_n16771, new_n16772, new_n16773, new_n16774,
    new_n16775, new_n16776, new_n16777, new_n16778, new_n16779, new_n16780,
    new_n16781, new_n16782, new_n16783, new_n16784, new_n16785, new_n16786,
    new_n16787, new_n16788, new_n16789, new_n16790, new_n16791, new_n16792,
    new_n16793, new_n16794, new_n16795, new_n16796, new_n16797, new_n16798,
    new_n16799, new_n16800, new_n16801, new_n16802, new_n16803, new_n16804,
    new_n16805, new_n16806, new_n16807, new_n16808, new_n16809, new_n16810,
    new_n16811, new_n16812, new_n16813, new_n16814, new_n16815, new_n16816,
    new_n16817, new_n16818, new_n16819, new_n16820, new_n16821, new_n16822,
    new_n16823, new_n16824, new_n16825, new_n16826, new_n16827, new_n16828,
    new_n16829, new_n16830, new_n16831, new_n16832, new_n16833, new_n16834,
    new_n16835, new_n16836, new_n16837, new_n16838, new_n16839, new_n16840,
    new_n16841, new_n16842, new_n16843, new_n16844, new_n16845, new_n16846,
    new_n16847, new_n16848, new_n16849, new_n16850, new_n16851, new_n16852,
    new_n16853, new_n16854, new_n16855, new_n16856, new_n16857, new_n16858,
    new_n16859, new_n16860, new_n16861, new_n16862, new_n16863, new_n16864,
    new_n16865, new_n16866, new_n16867, new_n16868, new_n16869, new_n16870,
    new_n16871, new_n16872, new_n16873, new_n16874, new_n16875, new_n16876,
    new_n16877, new_n16878, new_n16879, new_n16880, new_n16881, new_n16882,
    new_n16883, new_n16884, new_n16886, new_n16887, new_n16888, new_n16889,
    new_n16890, new_n16891, new_n16892, new_n16893, new_n16895, new_n16897,
    new_n16898, new_n16899, new_n16900, new_n16901, new_n16902, new_n16903,
    new_n16904, new_n16905, new_n16906, new_n16907, new_n16908, new_n16909,
    new_n16910, new_n16911, new_n16912, new_n16913, new_n16914, new_n16915,
    new_n16916, new_n16917, new_n16918, new_n16919, new_n16920, new_n16921,
    new_n16922, new_n16923, new_n16924, new_n16925, new_n16926, new_n16927,
    new_n16928, new_n16929, new_n16930, new_n16931, new_n16932, new_n16933,
    new_n16934, new_n16935, new_n16936, new_n16937, new_n16938, new_n16939,
    new_n16941, new_n16942, new_n16943, new_n16944, new_n16945, new_n16946,
    new_n16947, new_n16948, new_n16949, new_n16950, new_n16951, new_n16952,
    new_n16953, new_n16954, new_n16955, new_n16956, new_n16957, new_n16958,
    new_n16959, new_n16960, new_n16961, new_n16962, new_n16963, new_n16964,
    new_n16965, new_n16966, new_n16967, new_n16968, new_n16969, new_n16970,
    new_n16971, new_n16972, new_n16973, new_n16974, new_n16975, new_n16976,
    new_n16977, new_n16978, new_n16979, new_n16980, new_n16981, new_n16982,
    new_n16984, new_n16985, new_n16986, new_n16987, new_n16988, new_n16989,
    new_n16990, new_n16991, new_n16992, new_n16993, new_n16994, new_n16995,
    new_n16996, new_n16997, new_n16998, new_n16999, new_n17000, new_n17001,
    new_n17002, new_n17003, new_n17004, new_n17005, new_n17006, new_n17007,
    new_n17008, new_n17009, new_n17010, new_n17011, new_n17012, new_n17013,
    new_n17014, new_n17015, new_n17016, new_n17017, new_n17020, new_n17021,
    new_n17022, new_n17023, new_n17024, new_n17025, new_n17026, new_n17027,
    new_n17028, new_n17029, new_n17030, new_n17031, new_n17032, new_n17033,
    new_n17034, new_n17036, new_n17037, new_n17038, new_n17039, new_n17040,
    new_n17041, new_n17042, new_n17043, new_n17044, new_n17045, new_n17046,
    new_n17047, new_n17048, new_n17049, new_n17050, new_n17051, new_n17052,
    new_n17053, new_n17054, new_n17055, new_n17056, new_n17057, new_n17058,
    new_n17059, new_n17060, new_n17061, new_n17062, new_n17063, new_n17064,
    new_n17065, new_n17066, new_n17067, new_n17068, new_n17069, new_n17070,
    new_n17071, new_n17072, new_n17073, new_n17074, new_n17075, new_n17076,
    new_n17077, new_n17078, new_n17079, new_n17080, new_n17081, new_n17082,
    new_n17083, new_n17084, new_n17085, new_n17086, new_n17087, new_n17088,
    new_n17089, new_n17090, new_n17091, new_n17092, new_n17093, new_n17094,
    new_n17095, new_n17096, new_n17097, new_n17098, new_n17099, new_n17100,
    new_n17101, new_n17102, new_n17103, new_n17105, new_n17106, new_n17107,
    new_n17108, new_n17109, new_n17110, new_n17111, new_n17112, new_n17113,
    new_n17114, new_n17115, new_n17116, new_n17117, new_n17118, new_n17119,
    new_n17120, new_n17121, new_n17122, new_n17123, new_n17124, new_n17125,
    new_n17126, new_n17127, new_n17128, new_n17129, new_n17130, new_n17131,
    new_n17132, new_n17133, new_n17134, new_n17135, new_n17136, new_n17137,
    new_n17138, new_n17139, new_n17140, new_n17141, new_n17142, new_n17143,
    new_n17144, new_n17145, new_n17146, new_n17147, new_n17148, new_n17149,
    new_n17150, new_n17151, new_n17152, new_n17153, new_n17154, new_n17155,
    new_n17156, new_n17157, new_n17158, new_n17159, new_n17160, new_n17161,
    new_n17162, new_n17163, new_n17164, new_n17165, new_n17166, new_n17167,
    new_n17168, new_n17169, new_n17170, new_n17171, new_n17172, new_n17173,
    new_n17174, new_n17175, new_n17176, new_n17177, new_n17178, new_n17179,
    new_n17180, new_n17181, new_n17182, new_n17183, new_n17184, new_n17185,
    new_n17186, new_n17187, new_n17188, new_n17189, new_n17190, new_n17191,
    new_n17192, new_n17193, new_n17194, new_n17195, new_n17196, new_n17197,
    new_n17198, new_n17199, new_n17200, new_n17201, new_n17202, new_n17203,
    new_n17204, new_n17205, new_n17206, new_n17207, new_n17208, new_n17209,
    new_n17210, new_n17211, new_n17212, new_n17213, new_n17214, new_n17215,
    new_n17216, new_n17217, new_n17218, new_n17219, new_n17220, new_n17221,
    new_n17222, new_n17223, new_n17224, new_n17225, new_n17226, new_n17227,
    new_n17228, new_n17229, new_n17230, new_n17231, new_n17232, new_n17233,
    new_n17234, new_n17235, new_n17236, new_n17237, new_n17238, new_n17239,
    new_n17240, new_n17241, new_n17242, new_n17243, new_n17244, new_n17245,
    new_n17246, new_n17247, new_n17248, new_n17249, new_n17250, new_n17251,
    new_n17252, new_n17253, new_n17254, new_n17255, new_n17256, new_n17257,
    new_n17258, new_n17259, new_n17260, new_n17261, new_n17262, new_n17263,
    new_n17264, new_n17265, new_n17266, new_n17267, new_n17268, new_n17269,
    new_n17270, new_n17271, new_n17272, new_n17273, new_n17274, new_n17275,
    new_n17276, new_n17277, new_n17278, new_n17279, new_n17280, new_n17281,
    new_n17282, new_n17283, new_n17284, new_n17285, new_n17286, new_n17287,
    new_n17288, new_n17289, new_n17290, new_n17292, new_n17293, new_n17294,
    new_n17295, new_n17296, new_n17297, new_n17298, new_n17299, new_n17300,
    new_n17301, new_n17302, new_n17303, new_n17304, new_n17305, new_n17306,
    new_n17308, new_n17310, new_n17311, new_n17312, new_n17313, new_n17314,
    new_n17315, new_n17316, new_n17317, new_n17318, new_n17319, new_n17320,
    new_n17321, new_n17326, new_n17327, new_n17328, new_n17329, new_n17330,
    new_n17331, new_n17332, new_n17333, new_n17334, new_n17341, new_n17342,
    new_n17343, new_n17344, new_n17345, new_n17346, new_n17347, new_n17348,
    new_n17349, new_n17350, new_n17351, new_n17352, new_n17353, new_n17354,
    new_n17355, new_n17356, new_n17357, new_n17358, new_n17359, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366,
    new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372,
    new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378,
    new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384,
    new_n17385, new_n17386, new_n17387, new_n17388, new_n17389, new_n17390,
    new_n17391, new_n17392, new_n17393, new_n17394, new_n17395, new_n17396,
    new_n17397, new_n17398, new_n17399, new_n17400, new_n17401, new_n17402,
    new_n17403, new_n17404, new_n17405, new_n17406, new_n17407, new_n17408,
    new_n17409, new_n17410, new_n17411, new_n17412, new_n17413, new_n17414,
    new_n17415, new_n17416, new_n17417, new_n17418, new_n17419, new_n17420,
    new_n17421, new_n17422, new_n17423, new_n17424, new_n17425, new_n17426,
    new_n17427, new_n17428, new_n17429, new_n17430, new_n17431, new_n17432,
    new_n17433, new_n17434, new_n17435, new_n17436, new_n17437, new_n17438,
    new_n17439, new_n17440, new_n17442, new_n17443, new_n17444, new_n17445,
    new_n17446, new_n17447, new_n17448, new_n17449, new_n17450, new_n17451,
    new_n17452, new_n17453, new_n17454, new_n17455, new_n17456, new_n17457,
    new_n17458, new_n17459, new_n17460, new_n17461, new_n17462, new_n17463,
    new_n17464, new_n17465, new_n17466, new_n17467, new_n17468, new_n17469,
    new_n17470, new_n17471, new_n17472, new_n17473, new_n17474, new_n17475,
    new_n17476, new_n17477, new_n17478, new_n17479, new_n17480, new_n17481,
    new_n17482, new_n17484, new_n17485, new_n17486, new_n17487, new_n17488,
    new_n17489, new_n17490, new_n17491, new_n17492, new_n17493, new_n17494,
    new_n17495, new_n17496, new_n17497, new_n17498, new_n17499, new_n17500,
    new_n17501, new_n17502, new_n17503, new_n17504, new_n17505, new_n17506,
    new_n17507, new_n17508, new_n17509, new_n17510, new_n17511, new_n17512,
    new_n17513, new_n17514, new_n17515, new_n17516, new_n17517, new_n17518,
    new_n17519, new_n17520, new_n17521, new_n17522, new_n17523, new_n17524,
    new_n17525, new_n17526, new_n17527, new_n17528, new_n17529, new_n17530,
    new_n17531, new_n17532, new_n17533, new_n17534, new_n17535, new_n17536,
    new_n17537, new_n17538, new_n17539, new_n17540, new_n17541, new_n17542,
    new_n17543, new_n17544, new_n17545, new_n17546, new_n17547, new_n17548,
    new_n17549, new_n17550, new_n17551, new_n17552, new_n17553, new_n17554,
    new_n17555, new_n17556, new_n17557, new_n17558, new_n17559, new_n17560,
    new_n17561, new_n17562, new_n17563, new_n17564, new_n17565, new_n17566,
    new_n17567, new_n17568, new_n17569, new_n17570, new_n17571, new_n17572,
    new_n17573, new_n17574, new_n17575, new_n17576, new_n17577, new_n17578,
    new_n17579, new_n17580, new_n17581, new_n17582, new_n17583, new_n17584,
    new_n17585, new_n17586, new_n17587, new_n17588, new_n17589, new_n17590,
    new_n17591, new_n17592, new_n17593, new_n17594, new_n17595, new_n17596,
    new_n17597, new_n17598, new_n17599, new_n17600, new_n17601, new_n17602,
    new_n17603, new_n17604, new_n17605, new_n17606, new_n17607, new_n17608,
    new_n17610, new_n17611, new_n17612, new_n17613, new_n17614, new_n17615,
    new_n17616, new_n17617, new_n17618, new_n17619, new_n17620, new_n17621,
    new_n17622, new_n17623, new_n17624, new_n17625, new_n17626, new_n17627,
    new_n17628, new_n17629, new_n17630, new_n17631, new_n17632, new_n17633,
    new_n17634, new_n17635, new_n17636, new_n17637, new_n17638, new_n17639,
    new_n17640, new_n17641, new_n17642, new_n17643, new_n17644, new_n17645,
    new_n17646, new_n17647, new_n17648, new_n17649, new_n17650, new_n17651,
    new_n17652, new_n17653, new_n17654, new_n17657, new_n17658, new_n17659,
    new_n17660, new_n17661, new_n17662, new_n17663, new_n17664, new_n17665,
    new_n17666, new_n17667, new_n17668, new_n17669, new_n17670, new_n17671,
    new_n17672, new_n17673, new_n17676, new_n17677, new_n17678, new_n17679,
    new_n17680, new_n17681, new_n17682, new_n17683, new_n17684, new_n17685,
    new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694,
    new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700,
    new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706,
    new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712,
    new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718,
    new_n17719, new_n17720, new_n17721, new_n17722, new_n17723, new_n17724,
    new_n17725, new_n17726, new_n17727, new_n17728, new_n17729, new_n17730,
    new_n17731, new_n17732, new_n17733, new_n17734, new_n17735, new_n17736,
    new_n17737, new_n17740, new_n17741, new_n17742, new_n17743, new_n17744,
    new_n17745, new_n17746, new_n17747, new_n17748, new_n17749, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780,
    new_n17781, new_n17782, new_n17783, new_n17784, new_n17785, new_n17786,
    new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792,
    new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798,
    new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17806, new_n17807, new_n17809, new_n17810, new_n17811,
    new_n17812, new_n17813, new_n17814, new_n17815, new_n17816, new_n17817,
    new_n17818, new_n17819, new_n17820, new_n17821, new_n17822, new_n17823,
    new_n17824, new_n17825, new_n17826, new_n17827, new_n17828, new_n17829,
    new_n17830, new_n17831, new_n17832, new_n17833, new_n17834, new_n17835,
    new_n17836, new_n17837, new_n17838, new_n17839, new_n17840, new_n17841,
    new_n17842, new_n17843, new_n17844, new_n17845, new_n17846, new_n17847,
    new_n17849, new_n17850, new_n17851, new_n17852, new_n17853, new_n17854,
    new_n17855, new_n17856, new_n17857, new_n17858, new_n17859, new_n17860,
    new_n17861, new_n17862, new_n17863, new_n17864, new_n17865, new_n17866,
    new_n17867, new_n17868, new_n17869, new_n17870, new_n17871, new_n17872,
    new_n17873, new_n17874, new_n17875, new_n17876, new_n17877, new_n17878,
    new_n17879, new_n17880, new_n17881, new_n17882, new_n17883, new_n17884,
    new_n17885, new_n17886, new_n17887, new_n17888, new_n17889, new_n17890,
    new_n17891, new_n17892, new_n17893, new_n17894, new_n17895, new_n17896,
    new_n17897, new_n17898, new_n17899, new_n17900, new_n17901, new_n17902,
    new_n17903, new_n17904, new_n17906, new_n17911, new_n17912, new_n17913,
    new_n17914, new_n17915, new_n17916, new_n17917, new_n17918, new_n17919,
    new_n17920, new_n17921, new_n17922, new_n17923, new_n17924, new_n17925,
    new_n17926, new_n17927, new_n17928, new_n17929, new_n17930, new_n17931,
    new_n17932, new_n17933, new_n17934, new_n17935, new_n17936, new_n17937,
    new_n17938, new_n17939, new_n17940, new_n17941, new_n17942, new_n17943,
    new_n17944, new_n17945, new_n17946, new_n17947, new_n17948, new_n17949,
    new_n17950, new_n17951, new_n17952, new_n17953, new_n17954, new_n17955,
    new_n17956, new_n17957, new_n17958, new_n17959, new_n17960, new_n17961,
    new_n17962, new_n17963, new_n17964, new_n17965, new_n17966, new_n17967,
    new_n17968, new_n17969, new_n17970, new_n17971, new_n17972, new_n17973,
    new_n17974, new_n17975, new_n17976, new_n17977, new_n17978, new_n17979,
    new_n17980, new_n17981, new_n17982, new_n17983, new_n17984, new_n17985,
    new_n17986, new_n17987, new_n17988, new_n17989, new_n17990, new_n17993,
    new_n17994, new_n17995, new_n17996, new_n17997, new_n17998, new_n17999,
    new_n18000, new_n18001, new_n18002, new_n18003, new_n18004, new_n18005,
    new_n18006, new_n18007, new_n18008, new_n18009, new_n18010, new_n18011,
    new_n18012, new_n18013, new_n18014, new_n18015, new_n18016, new_n18017,
    new_n18018, new_n18019, new_n18020, new_n18021, new_n18024, new_n18025,
    new_n18026, new_n18027, new_n18028, new_n18029, new_n18030, new_n18031,
    new_n18032, new_n18033, new_n18034, new_n18035, new_n18036, new_n18037,
    new_n18038, new_n18039, new_n18040, new_n18041, new_n18042, new_n18043,
    new_n18044, new_n18045, new_n18046, new_n18047, new_n18048, new_n18049,
    new_n18050, new_n18051, new_n18052, new_n18057, new_n18058, new_n18059,
    new_n18061, new_n18062, new_n18063, new_n18064, new_n18065, new_n18066,
    new_n18067, new_n18068, new_n18069, new_n18070, new_n18071, new_n18072,
    new_n18073, new_n18074, new_n18075, new_n18076, new_n18077, new_n18078,
    new_n18079, new_n18080, new_n18081, new_n18082, new_n18083, new_n18084,
    new_n18085, new_n18086, new_n18087, new_n18088, new_n18089, new_n18090,
    new_n18091, new_n18092, new_n18093, new_n18094, new_n18095, new_n18096,
    new_n18097, new_n18098, new_n18099, new_n18100, new_n18101, new_n18102,
    new_n18103, new_n18104, new_n18105, new_n18106, new_n18107, new_n18108,
    new_n18109, new_n18110, new_n18111, new_n18112, new_n18113, new_n18114,
    new_n18115, new_n18116, new_n18117, new_n18118, new_n18119, new_n18120,
    new_n18121, new_n18122, new_n18123, new_n18124, new_n18125, new_n18126,
    new_n18127, new_n18128, new_n18129, new_n18130, new_n18131, new_n18132,
    new_n18133, new_n18134, new_n18135, new_n18136, new_n18137, new_n18138,
    new_n18139, new_n18140, new_n18141, new_n18142, new_n18143, new_n18144,
    new_n18145, new_n18146, new_n18147, new_n18148, new_n18149, new_n18150,
    new_n18151, new_n18152, new_n18153, new_n18154, new_n18155, new_n18156,
    new_n18157, new_n18158, new_n18159, new_n18160, new_n18161, new_n18162,
    new_n18163, new_n18164, new_n18165, new_n18166, new_n18170, new_n18171,
    new_n18172, new_n18173, new_n18174, new_n18175, new_n18176, new_n18177,
    new_n18178, new_n18179, new_n18180, new_n18181, new_n18182, new_n18183,
    new_n18184, new_n18185, new_n18186, new_n18187, new_n18188, new_n18189,
    new_n18190, new_n18191, new_n18192, new_n18193, new_n18194, new_n18201,
    new_n18202, new_n18203, new_n18204, new_n18205, new_n18206, new_n18207,
    new_n18208, new_n18209, new_n18210, new_n18211, new_n18212, new_n18213,
    new_n18214, new_n18215, new_n18216, new_n18217, new_n18218, new_n18219,
    new_n18220, new_n18221, new_n18222, new_n18223, new_n18224, new_n18225,
    new_n18226, new_n18227, new_n18228, new_n18229, new_n18230, new_n18231,
    new_n18232, new_n18233, new_n18234, new_n18235, new_n18236, new_n18237,
    new_n18238, new_n18239, new_n18240, new_n18241, new_n18242, new_n18243,
    new_n18244, new_n18245, new_n18246, new_n18247, new_n18248, new_n18249,
    new_n18250, new_n18251, new_n18252, new_n18253, new_n18254, new_n18255,
    new_n18256, new_n18257, new_n18258, new_n18259, new_n18260, new_n18261,
    new_n18262, new_n18263, new_n18264, new_n18265, new_n18266, new_n18267,
    new_n18268, new_n18269, new_n18270, new_n18271, new_n18272, new_n18273,
    new_n18274, new_n18275, new_n18276, new_n18277, new_n18278, new_n18279,
    new_n18280, new_n18281, new_n18282, new_n18283, new_n18284, new_n18285,
    new_n18286, new_n18288, new_n18290, new_n18291, new_n18292, new_n18293,
    new_n18294, new_n18295, new_n18296, new_n18297, new_n18298, new_n18299,
    new_n18300, new_n18301, new_n18302, new_n18303, new_n18304, new_n18305,
    new_n18306, new_n18307, new_n18308, new_n18309, new_n18310, new_n18311,
    new_n18312, new_n18313, new_n18314, new_n18315, new_n18316, new_n18317,
    new_n18318, new_n18319, new_n18320, new_n18321, new_n18322, new_n18323,
    new_n18324, new_n18325, new_n18326, new_n18327, new_n18328, new_n18329,
    new_n18330, new_n18331, new_n18332, new_n18333, new_n18334, new_n18335,
    new_n18336, new_n18337, new_n18338, new_n18339, new_n18340, new_n18341,
    new_n18342, new_n18343, new_n18344, new_n18345, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18350, new_n18351, new_n18352, new_n18353,
    new_n18354, new_n18355, new_n18356, new_n18357, new_n18358, new_n18359,
    new_n18360, new_n18361, new_n18362, new_n18363, new_n18364, new_n18365,
    new_n18366, new_n18367, new_n18368, new_n18369, new_n18370, new_n18371,
    new_n18372, new_n18373, new_n18374, new_n18375, new_n18376, new_n18378,
    new_n18379, new_n18380, new_n18381, new_n18382, new_n18383, new_n18384,
    new_n18385, new_n18386, new_n18387, new_n18388, new_n18389, new_n18390,
    new_n18391, new_n18392, new_n18393, new_n18394, new_n18395, new_n18396,
    new_n18397, new_n18398, new_n18399, new_n18400, new_n18401, new_n18402,
    new_n18403, new_n18404, new_n18405, new_n18406, new_n18407, new_n18408,
    new_n18409, new_n18410, new_n18411, new_n18412, new_n18413, new_n18414,
    new_n18415, new_n18416, new_n18417, new_n18418, new_n18419, new_n18420,
    new_n18421, new_n18422, new_n18423, new_n18424, new_n18425, new_n18426,
    new_n18427, new_n18428, new_n18429, new_n18430, new_n18431, new_n18432,
    new_n18433, new_n18434, new_n18435, new_n18436, new_n18437, new_n18439,
    new_n18440, new_n18441, new_n18443, new_n18444, new_n18445, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451, new_n18452,
    new_n18453, new_n18454, new_n18455, new_n18456, new_n18457, new_n18458,
    new_n18459, new_n18460, new_n18461, new_n18462, new_n18463, new_n18464,
    new_n18465, new_n18466, new_n18467, new_n18468, new_n18469, new_n18470,
    new_n18471, new_n18472, new_n18473, new_n18474, new_n18475, new_n18476,
    new_n18481, new_n18482, new_n18483, new_n18484, new_n18485, new_n18486,
    new_n18487, new_n18488, new_n18489, new_n18490, new_n18491, new_n18492,
    new_n18493, new_n18494, new_n18495, new_n18496, new_n18497, new_n18498,
    new_n18499, new_n18500, new_n18501, new_n18506, new_n18507, new_n18508,
    new_n18509, new_n18510, new_n18511, new_n18512, new_n18513, new_n18514,
    new_n18515, new_n18516, new_n18517, new_n18518, new_n18519, new_n18520,
    new_n18521, new_n18522, new_n18523, new_n18524, new_n18525, new_n18526,
    new_n18527, new_n18528, new_n18529, new_n18530, new_n18531, new_n18532,
    new_n18533, new_n18534, new_n18535, new_n18536, new_n18537, new_n18538,
    new_n18539, new_n18540, new_n18541, new_n18542, new_n18543, new_n18544,
    new_n18545, new_n18546, new_n18547, new_n18548, new_n18549, new_n18550,
    new_n18551, new_n18553, new_n18554, new_n18555, new_n18557, new_n18558,
    new_n18559, new_n18560, new_n18561, new_n18562, new_n18563, new_n18564,
    new_n18565, new_n18566, new_n18567, new_n18568, new_n18569, new_n18573,
    new_n18574, new_n18575, new_n18576, new_n18577, new_n18578, new_n18579,
    new_n18580, new_n18581, new_n18582, new_n18583, new_n18584, new_n18585,
    new_n18586, new_n18587, new_n18588, new_n18589, new_n18590, new_n18591,
    new_n18592, new_n18594, new_n18595, new_n18596, new_n18597, new_n18598,
    new_n18599, new_n18600, new_n18601, new_n18602, new_n18603, new_n18604,
    new_n18605, new_n18606, new_n18607, new_n18608, new_n18609, new_n18610,
    new_n18611, new_n18612, new_n18613, new_n18614, new_n18615, new_n18616,
    new_n18617, new_n18618, new_n18619, new_n18620, new_n18621, new_n18622,
    new_n18623, new_n18624, new_n18625, new_n18626, new_n18627, new_n18628,
    new_n18629, new_n18630, new_n18631, new_n18632, new_n18633, new_n18634,
    new_n18635, new_n18636, new_n18637, new_n18638, new_n18639, new_n18640,
    new_n18641, new_n18642, new_n18643, new_n18644, new_n18645, new_n18646,
    new_n18647, new_n18648, new_n18649, new_n18650, new_n18651, new_n18652,
    new_n18653, new_n18654, new_n18655, new_n18656, new_n18657, new_n18658,
    new_n18659, new_n18660, new_n18662, new_n18663, new_n18664, new_n18665,
    new_n18666, new_n18667, new_n18668, new_n18669, new_n18671, new_n18672,
    new_n18673, new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679, new_n18680, new_n18681, new_n18682, new_n18683, new_n18684,
    new_n18685, new_n18686, new_n18687, new_n18688, new_n18689, new_n18690,
    new_n18691, new_n18692, new_n18693, new_n18694, new_n18695, new_n18696,
    new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702,
    new_n18703, new_n18704, new_n18705, new_n18706, new_n18707, new_n18708,
    new_n18709, new_n18710, new_n18711, new_n18712, new_n18713, new_n18714,
    new_n18715, new_n18716, new_n18717, new_n18718, new_n18719, new_n18720,
    new_n18721, new_n18722, new_n18723, new_n18724, new_n18725, new_n18726,
    new_n18727, new_n18728, new_n18729, new_n18730, new_n18731, new_n18732,
    new_n18733, new_n18734, new_n18735, new_n18736, new_n18737, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745, new_n18746, new_n18747, new_n18748, new_n18749, new_n18750,
    new_n18751, new_n18752, new_n18753, new_n18754, new_n18755, new_n18756,
    new_n18757, new_n18758, new_n18759, new_n18760, new_n18761, new_n18762,
    new_n18763, new_n18764, new_n18765, new_n18766, new_n18767, new_n18768,
    new_n18769, new_n18770, new_n18771, new_n18772, new_n18773, new_n18774,
    new_n18775, new_n18776, new_n18777, new_n18778, new_n18779, new_n18780,
    new_n18781, new_n18782, new_n18783, new_n18784, new_n18785, new_n18786,
    new_n18787, new_n18788, new_n18789, new_n18790, new_n18791, new_n18792,
    new_n18793, new_n18794, new_n18795, new_n18796, new_n18797, new_n18798,
    new_n18799, new_n18800, new_n18801, new_n18802, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822,
    new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828,
    new_n18829, new_n18830, new_n18831, new_n18832, new_n18833, new_n18834,
    new_n18835, new_n18836, new_n18837, new_n18838, new_n18839, new_n18840,
    new_n18841, new_n18842, new_n18843, new_n18844, new_n18845, new_n18846,
    new_n18847, new_n18848, new_n18849, new_n18850, new_n18851, new_n18852,
    new_n18853, new_n18854, new_n18855, new_n18856, new_n18857, new_n18858,
    new_n18859, new_n18860, new_n18861, new_n18862, new_n18863, new_n18864,
    new_n18865, new_n18866, new_n18867, new_n18868, new_n18869, new_n18870,
    new_n18871, new_n18872, new_n18873, new_n18874, new_n18875, new_n18876,
    new_n18877, new_n18878, new_n18879, new_n18880, new_n18881, new_n18882,
    new_n18883, new_n18884, new_n18885, new_n18886, new_n18887, new_n18888,
    new_n18889, new_n18890, new_n18891, new_n18892, new_n18893, new_n18894,
    new_n18895, new_n18896, new_n18897, new_n18898, new_n18899, new_n18900,
    new_n18901, new_n18902, new_n18903, new_n18904, new_n18905, new_n18907,
    new_n18908, new_n18909, new_n18910, new_n18911, new_n18912, new_n18913,
    new_n18914, new_n18915, new_n18916, new_n18917, new_n18918, new_n18919,
    new_n18920, new_n18921, new_n18922, new_n18923, new_n18924, new_n18925,
    new_n18926, new_n18927, new_n18928, new_n18929, new_n18930, new_n18931,
    new_n18932, new_n18933, new_n18934, new_n18935, new_n18936, new_n18937,
    new_n18938, new_n18939, new_n18940, new_n18941, new_n18942, new_n18943,
    new_n18944, new_n18946, new_n18947, new_n18948, new_n18949, new_n18950,
    new_n18951, new_n18952, new_n18953, new_n18954, new_n18955, new_n18956,
    new_n18957, new_n18958, new_n18959, new_n18960, new_n18961, new_n18964,
    new_n18965, new_n18966, new_n18967, new_n18968, new_n18973, new_n18974,
    new_n18975, new_n18976, new_n18977, new_n18978, new_n18979, new_n18980,
    new_n18981, new_n18982, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999, new_n19000, new_n19001, new_n19002, new_n19003, new_n19004,
    new_n19005, new_n19006, new_n19007, new_n19008, new_n19009, new_n19010,
    new_n19011, new_n19012, new_n19013, new_n19014, new_n19015, new_n19016,
    new_n19017, new_n19018, new_n19019, new_n19020, new_n19021, new_n19022,
    new_n19023, new_n19024, new_n19025, new_n19026, new_n19027, new_n19028,
    new_n19029, new_n19030, new_n19031, new_n19032, new_n19033, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042, new_n19043, new_n19044, new_n19045, new_n19046,
    new_n19047, new_n19048, new_n19049, new_n19050, new_n19051, new_n19052,
    new_n19053, new_n19054, new_n19055, new_n19056, new_n19057, new_n19058,
    new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19067,
    new_n19068, new_n19069, new_n19070, new_n19071, new_n19072, new_n19073,
    new_n19074, new_n19075, new_n19076, new_n19077, new_n19078, new_n19079,
    new_n19080, new_n19081, new_n19082, new_n19083, new_n19084, new_n19086,
    new_n19087, new_n19088, new_n19089, new_n19090, new_n19091, new_n19092,
    new_n19093, new_n19094, new_n19095, new_n19096, new_n19097, new_n19098,
    new_n19099, new_n19100, new_n19101, new_n19102, new_n19103, new_n19104,
    new_n19105, new_n19106, new_n19107, new_n19108, new_n19109, new_n19110,
    new_n19111, new_n19112, new_n19113, new_n19114, new_n19115, new_n19116,
    new_n19117, new_n19118, new_n19119, new_n19120, new_n19121, new_n19122,
    new_n19123, new_n19124, new_n19125, new_n19126, new_n19127, new_n19128,
    new_n19129, new_n19130, new_n19131, new_n19132, new_n19133, new_n19134,
    new_n19135, new_n19138, new_n19139, new_n19140, new_n19141, new_n19142,
    new_n19143, new_n19144, new_n19145, new_n19146, new_n19147, new_n19148,
    new_n19149, new_n19150, new_n19151, new_n19152, new_n19153, new_n19154,
    new_n19155, new_n19156, new_n19157, new_n19158, new_n19159, new_n19160,
    new_n19161, new_n19162, new_n19163, new_n19164, new_n19165, new_n19166,
    new_n19167, new_n19168, new_n19169, new_n19170, new_n19171, new_n19172,
    new_n19173, new_n19174, new_n19175, new_n19176, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19185,
    new_n19186, new_n19187, new_n19188, new_n19189, new_n19190, new_n19191,
    new_n19192, new_n19193, new_n19194, new_n19195, new_n19196, new_n19197,
    new_n19198, new_n19199, new_n19200, new_n19201, new_n19202, new_n19203,
    new_n19204, new_n19205, new_n19206, new_n19207, new_n19208, new_n19209,
    new_n19210, new_n19211, new_n19212, new_n19213, new_n19214, new_n19215,
    new_n19216, new_n19217, new_n19218, new_n19219, new_n19220, new_n19225,
    new_n19226, new_n19227, new_n19228, new_n19229, new_n19230, new_n19231,
    new_n19232, new_n19233, new_n19234, new_n19235, new_n19236, new_n19237,
    new_n19238, new_n19239, new_n19240, new_n19241, new_n19242, new_n19243,
    new_n19244, new_n19245, new_n19246, new_n19247, new_n19248, new_n19249,
    new_n19250, new_n19251, new_n19252, new_n19253, new_n19254, new_n19255,
    new_n19256, new_n19261, new_n19262, new_n19263, new_n19264, new_n19265,
    new_n19266, new_n19267, new_n19268, new_n19269, new_n19270, new_n19271,
    new_n19272, new_n19273, new_n19274, new_n19275, new_n19276, new_n19277,
    new_n19278, new_n19279, new_n19280, new_n19281, new_n19282, new_n19283,
    new_n19284, new_n19285, new_n19286, new_n19287, new_n19288, new_n19289,
    new_n19290, new_n19291, new_n19292, new_n19293, new_n19294, new_n19295,
    new_n19296, new_n19297, new_n19298, new_n19299, new_n19300, new_n19301,
    new_n19302, new_n19303, new_n19304, new_n19305, new_n19306, new_n19307,
    new_n19308, new_n19309, new_n19310, new_n19311, new_n19312, new_n19313,
    new_n19314, new_n19315, new_n19316, new_n19317, new_n19318, new_n19319,
    new_n19320, new_n19321, new_n19322, new_n19323, new_n19324, new_n19325,
    new_n19326, new_n19327, new_n19328, new_n19329, new_n19330, new_n19331,
    new_n19332, new_n19333, new_n19334, new_n19335, new_n19336, new_n19337,
    new_n19338, new_n19339, new_n19340, new_n19341, new_n19342, new_n19343,
    new_n19344, new_n19345, new_n19346, new_n19352, new_n19353, new_n19354,
    new_n19355, new_n19356, new_n19357, new_n19358, new_n19359, new_n19360,
    new_n19361, new_n19362, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367, new_n19368, new_n19370, new_n19371, new_n19372, new_n19373,
    new_n19374, new_n19375, new_n19376, new_n19377, new_n19378, new_n19379,
    new_n19380, new_n19381, new_n19382, new_n19383, new_n19384, new_n19385,
    new_n19386, new_n19387, new_n19388, new_n19389, new_n19390, new_n19391,
    new_n19392, new_n19393, new_n19394, new_n19395, new_n19396, new_n19397,
    new_n19398, new_n19399, new_n19400, new_n19401, new_n19402, new_n19403,
    new_n19404, new_n19405, new_n19406, new_n19407, new_n19408, new_n19409,
    new_n19410, new_n19411, new_n19412, new_n19413, new_n19414, new_n19415,
    new_n19416, new_n19417, new_n19418, new_n19419, new_n19420, new_n19421,
    new_n19422, new_n19423, new_n19424, new_n19425, new_n19426, new_n19427,
    new_n19428, new_n19429, new_n19430, new_n19431, new_n19432, new_n19433,
    new_n19434, new_n19435, new_n19436, new_n19437, new_n19438, new_n19439,
    new_n19440, new_n19441, new_n19442, new_n19443, new_n19444, new_n19445,
    new_n19446, new_n19447, new_n19448, new_n19449, new_n19450, new_n19455,
    new_n19456, new_n19457, new_n19458, new_n19459, new_n19460, new_n19461,
    new_n19462, new_n19463, new_n19464, new_n19465, new_n19466, new_n19467,
    new_n19468, new_n19469, new_n19470, new_n19471, new_n19472, new_n19473,
    new_n19474, new_n19475, new_n19476, new_n19477, new_n19478, new_n19479,
    new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485,
    new_n19486, new_n19487, new_n19488, new_n19489, new_n19490, new_n19491,
    new_n19493, new_n19494, new_n19495, new_n19496, new_n19497, new_n19498,
    new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504,
    new_n19505, new_n19506, new_n19507, new_n19508, new_n19509, new_n19510,
    new_n19511, new_n19512, new_n19513, new_n19514, new_n19515, new_n19516,
    new_n19517, new_n19518, new_n19519, new_n19520, new_n19523, new_n19524,
    new_n19525, new_n19526, new_n19527, new_n19528, new_n19529, new_n19530,
    new_n19531, new_n19532, new_n19533, new_n19534, new_n19535, new_n19536,
    new_n19537, new_n19538, new_n19539, new_n19540, new_n19541, new_n19542,
    new_n19543, new_n19544, new_n19545, new_n19546, new_n19547, new_n19548,
    new_n19549, new_n19550, new_n19551, new_n19552, new_n19553, new_n19554,
    new_n19555, new_n19556, new_n19557, new_n19558, new_n19559, new_n19560,
    new_n19561, new_n19562, new_n19563, new_n19564, new_n19565, new_n19566,
    new_n19567, new_n19568, new_n19569, new_n19570, new_n19571, new_n19572,
    new_n19573, new_n19574, new_n19575, new_n19576, new_n19577, new_n19578,
    new_n19579, new_n19580, new_n19581, new_n19582, new_n19583, new_n19584,
    new_n19585, new_n19586, new_n19587, new_n19588, new_n19591, new_n19592,
    new_n19593, new_n19594, new_n19595, new_n19596, new_n19597, new_n19598,
    new_n19599, new_n19600, new_n19601, new_n19602, new_n19603, new_n19604,
    new_n19605, new_n19606, new_n19607, new_n19608, new_n19609, new_n19611,
    new_n19612, new_n19613, new_n19614, new_n19615, new_n19616, new_n19617,
    new_n19618, new_n19619, new_n19620, new_n19621, new_n19622, new_n19623,
    new_n19624, new_n19625, new_n19626, new_n19627, new_n19628, new_n19629,
    new_n19630, new_n19631, new_n19632, new_n19633, new_n19634, new_n19636,
    new_n19637, new_n19638, new_n19639, new_n19640, new_n19641, new_n19642,
    new_n19643, new_n19644, new_n19645, new_n19646, new_n19647, new_n19648,
    new_n19649, new_n19650, new_n19651, new_n19652, new_n19653, new_n19654,
    new_n19655, new_n19656, new_n19657, new_n19658, new_n19659, new_n19660,
    new_n19661, new_n19662, new_n19663, new_n19664, new_n19665, new_n19666,
    new_n19667, new_n19668, new_n19669, new_n19670, new_n19671, new_n19672,
    new_n19673, new_n19674, new_n19675, new_n19676, new_n19680, new_n19681,
    new_n19682, new_n19683, new_n19684, new_n19685, new_n19686, new_n19687,
    new_n19688, new_n19689, new_n19690, new_n19691, new_n19692, new_n19693,
    new_n19694, new_n19695, new_n19696, new_n19697, new_n19698, new_n19699,
    new_n19700, new_n19701, new_n19702, new_n19703, new_n19704, new_n19705,
    new_n19706, new_n19707, new_n19708, new_n19709, new_n19710, new_n19711,
    new_n19712, new_n19713, new_n19714, new_n19715, new_n19716, new_n19717,
    new_n19718, new_n19719, new_n19720, new_n19721, new_n19722, new_n19723,
    new_n19724, new_n19725, new_n19727, new_n19728, new_n19729, new_n19730,
    new_n19731, new_n19732, new_n19733, new_n19734, new_n19735, new_n19736,
    new_n19737, new_n19738, new_n19739, new_n19740, new_n19741, new_n19742,
    new_n19743, new_n19744, new_n19745, new_n19746, new_n19747, new_n19748,
    new_n19749, new_n19750, new_n19751, new_n19752, new_n19753, new_n19754,
    new_n19755, new_n19756, new_n19757, new_n19759, new_n19760, new_n19761,
    new_n19762, new_n19763, new_n19764, new_n19765, new_n19766, new_n19767,
    new_n19768, new_n19769, new_n19770, new_n19771, new_n19772, new_n19773,
    new_n19774, new_n19775, new_n19776, new_n19777, new_n19781, new_n19783,
    new_n19784, new_n19785, new_n19786, new_n19787, new_n19788, new_n19789,
    new_n19790, new_n19791, new_n19792, new_n19793, new_n19794, new_n19797,
    new_n19798, new_n19799, new_n19800, new_n19801, new_n19802, new_n19803,
    new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809,
    new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815,
    new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821,
    new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827,
    new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833,
    new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839,
    new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845,
    new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851,
    new_n19852, new_n19853, new_n19854, new_n19855, new_n19856, new_n19857,
    new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863,
    new_n19864, new_n19865, new_n19866, new_n19867, new_n19872, new_n19873,
    new_n19874, new_n19875, new_n19876, new_n19877, new_n19878, new_n19879,
    new_n19880, new_n19881, new_n19882, new_n19883, new_n19884, new_n19885,
    new_n19886, new_n19890, new_n19891, new_n19892, new_n19893, new_n19894,
    new_n19895, new_n19896, new_n19897, new_n19898, new_n19899, new_n19900,
    new_n19901, new_n19902, new_n19903, new_n19904, new_n19905, new_n19906,
    new_n19907, new_n19908, new_n19909, new_n19910, new_n19911, new_n19912,
    new_n19913, new_n19914, new_n19915, new_n19916, new_n19917, new_n19918,
    new_n19919, new_n19920, new_n19921, new_n19922, new_n19923, new_n19924,
    new_n19925, new_n19926, new_n19927, new_n19928, new_n19929, new_n19930,
    new_n19931, new_n19932, new_n19933, new_n19934, new_n19935, new_n19936,
    new_n19937, new_n19938, new_n19939, new_n19940, new_n19941, new_n19942,
    new_n19943, new_n19944, new_n19945, new_n19946, new_n19947, new_n19948,
    new_n19949, new_n19950, new_n19951, new_n19952, new_n19953, new_n19954,
    new_n19955, new_n19956, new_n19957, new_n19958, new_n19959, new_n19960,
    new_n19961, new_n19962, new_n19963, new_n19964, new_n19965, new_n19966,
    new_n19967, new_n19968, new_n19969, new_n19970, new_n19971, new_n19972,
    new_n19973, new_n19974, new_n19975, new_n19976, new_n19977, new_n19978,
    new_n19979, new_n19980, new_n19981, new_n19982, new_n19983, new_n19984,
    new_n19985, new_n19986, new_n19987, new_n19988, new_n19989, new_n19990,
    new_n19991, new_n19992, new_n19993, new_n19994, new_n19995, new_n19996,
    new_n19997, new_n19998, new_n19999, new_n20000, new_n20002, new_n20009,
    new_n20010, new_n20011, new_n20012, new_n20013, new_n20014, new_n20015,
    new_n20016, new_n20017, new_n20018, new_n20019, new_n20020, new_n20021,
    new_n20022, new_n20023, new_n20024, new_n20025, new_n20026, new_n20027,
    new_n20028, new_n20029, new_n20030, new_n20031, new_n20032, new_n20033,
    new_n20034, new_n20035, new_n20036, new_n20037, new_n20038, new_n20039,
    new_n20040, new_n20041, new_n20042, new_n20043, new_n20044, new_n20045,
    new_n20046, new_n20047, new_n20048, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061, new_n20062, new_n20063, new_n20064, new_n20065, new_n20066,
    new_n20067, new_n20068, new_n20069, new_n20070, new_n20071, new_n20072,
    new_n20073, new_n20074, new_n20075, new_n20076, new_n20077, new_n20078,
    new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084,
    new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096,
    new_n20097, new_n20098, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108,
    new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114,
    new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126,
    new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20133,
    new_n20134, new_n20135, new_n20136, new_n20137, new_n20138, new_n20139,
    new_n20140, new_n20144, new_n20145, new_n20146, new_n20147, new_n20148,
    new_n20149, new_n20150, new_n20151, new_n20152, new_n20153, new_n20154,
    new_n20155, new_n20156, new_n20157, new_n20158, new_n20159, new_n20160,
    new_n20161, new_n20162, new_n20163, new_n20164, new_n20165, new_n20166,
    new_n20167, new_n20168, new_n20169, new_n20170, new_n20171, new_n20173,
    new_n20174, new_n20175, new_n20176, new_n20177, new_n20178, new_n20179,
    new_n20180, new_n20181, new_n20182, new_n20183, new_n20184, new_n20185,
    new_n20186, new_n20187, new_n20188, new_n20189, new_n20190, new_n20191,
    new_n20192, new_n20193, new_n20194, new_n20195, new_n20196, new_n20197,
    new_n20198, new_n20199, new_n20200, new_n20201, new_n20202, new_n20203,
    new_n20204, new_n20205, new_n20206, new_n20207, new_n20208, new_n20209,
    new_n20210, new_n20211, new_n20212, new_n20213, new_n20214, new_n20215,
    new_n20216, new_n20217, new_n20218, new_n20219, new_n20220, new_n20221,
    new_n20222, new_n20223, new_n20224, new_n20225, new_n20226, new_n20227,
    new_n20228, new_n20229, new_n20230, new_n20231, new_n20232, new_n20233,
    new_n20234, new_n20235, new_n20236, new_n20239, new_n20241, new_n20242,
    new_n20243, new_n20244, new_n20245, new_n20246, new_n20247, new_n20248,
    new_n20249, new_n20250, new_n20251, new_n20252, new_n20253, new_n20254,
    new_n20255, new_n20256, new_n20257, new_n20258, new_n20259, new_n20260,
    new_n20261, new_n20262, new_n20263, new_n20264, new_n20265, new_n20266,
    new_n20267, new_n20268, new_n20269, new_n20270, new_n20271, new_n20272,
    new_n20273, new_n20274, new_n20275, new_n20276, new_n20277, new_n20278,
    new_n20279, new_n20280, new_n20281, new_n20282, new_n20283, new_n20284,
    new_n20285, new_n20286, new_n20287, new_n20288, new_n20289, new_n20290,
    new_n20291, new_n20292, new_n20293, new_n20294, new_n20295, new_n20296,
    new_n20297, new_n20298, new_n20299, new_n20300, new_n20301, new_n20302,
    new_n20303, new_n20304, new_n20305, new_n20306, new_n20307, new_n20308,
    new_n20309, new_n20310, new_n20311, new_n20312, new_n20313, new_n20314,
    new_n20315, new_n20316, new_n20317, new_n20318, new_n20319, new_n20320,
    new_n20321, new_n20322, new_n20323, new_n20324, new_n20325, new_n20326,
    new_n20327, new_n20328, new_n20329, new_n20330, new_n20331, new_n20332,
    new_n20333, new_n20334, new_n20335, new_n20336, new_n20337, new_n20338,
    new_n20339, new_n20340, new_n20341, new_n20342, new_n20343, new_n20344,
    new_n20345, new_n20346, new_n20347, new_n20348, new_n20349, new_n20350,
    new_n20351, new_n20352, new_n20353, new_n20354, new_n20355, new_n20356,
    new_n20357, new_n20358, new_n20359, new_n20360, new_n20361, new_n20362,
    new_n20363, new_n20364, new_n20365, new_n20366, new_n20367, new_n20368,
    new_n20369, new_n20370, new_n20371, new_n20372, new_n20373, new_n20374,
    new_n20375, new_n20376, new_n20377, new_n20378, new_n20379, new_n20380,
    new_n20381, new_n20382, new_n20383, new_n20384, new_n20385, new_n20386,
    new_n20387, new_n20388, new_n20389, new_n20390, new_n20391, new_n20394,
    new_n20395, new_n20396, new_n20397, new_n20398, new_n20399, new_n20400,
    new_n20401, new_n20402, new_n20403, new_n20404, new_n20405, new_n20406,
    new_n20407, new_n20408, new_n20409, new_n20410, new_n20411, new_n20412,
    new_n20413, new_n20414, new_n20415, new_n20416, new_n20417, new_n20418,
    new_n20419, new_n20420, new_n20421, new_n20422, new_n20423, new_n20424,
    new_n20425, new_n20426, new_n20427, new_n20428, new_n20429, new_n20430,
    new_n20431, new_n20432, new_n20433, new_n20434, new_n20435, new_n20436,
    new_n20437, new_n20438, new_n20439, new_n20440, new_n20441, new_n20442,
    new_n20443, new_n20444, new_n20445, new_n20446, new_n20447, new_n20448,
    new_n20449, new_n20450, new_n20451, new_n20452, new_n20453, new_n20454,
    new_n20455, new_n20456, new_n20457, new_n20458, new_n20459, new_n20460,
    new_n20461, new_n20462, new_n20463, new_n20464, new_n20465, new_n20466,
    new_n20467, new_n20473, new_n20475, new_n20479, new_n20480, new_n20481,
    new_n20482, new_n20483, new_n20484, new_n20485, new_n20486, new_n20487,
    new_n20488, new_n20489, new_n20490, new_n20491, new_n20492, new_n20493,
    new_n20494, new_n20495, new_n20496, new_n20497, new_n20498, new_n20499,
    new_n20500, new_n20501, new_n20502, new_n20503, new_n20504, new_n20505,
    new_n20506, new_n20507, new_n20508, new_n20509, new_n20510, new_n20511,
    new_n20512, new_n20513, new_n20514, new_n20515, new_n20516, new_n20517,
    new_n20518, new_n20519, new_n20520, new_n20521, new_n20522, new_n20523,
    new_n20524, new_n20525, new_n20526, new_n20527, new_n20528, new_n20529,
    new_n20530, new_n20531, new_n20532, new_n20533, new_n20534, new_n20535,
    new_n20536, new_n20537, new_n20538, new_n20539, new_n20540, new_n20541,
    new_n20542, new_n20543, new_n20544, new_n20545, new_n20546, new_n20547,
    new_n20548, new_n20549, new_n20550, new_n20551, new_n20552, new_n20553,
    new_n20554, new_n20555, new_n20556, new_n20557, new_n20558, new_n20559,
    new_n20560, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565,
    new_n20566, new_n20567, new_n20568, new_n20569, new_n20570, new_n20571,
    new_n20572, new_n20573, new_n20574, new_n20575, new_n20576, new_n20577,
    new_n20578, new_n20579, new_n20580, new_n20581, new_n20582, new_n20583,
    new_n20584, new_n20585, new_n20586, new_n20587, new_n20588, new_n20589,
    new_n20590, new_n20591, new_n20592, new_n20593, new_n20594, new_n20595,
    new_n20596, new_n20597, new_n20598, new_n20599, new_n20600, new_n20601,
    new_n20602, new_n20603, new_n20604, new_n20605, new_n20606, new_n20607,
    new_n20608, new_n20609, new_n20610, new_n20611, new_n20612, new_n20613,
    new_n20614, new_n20615, new_n20616, new_n20617, new_n20618, new_n20619,
    new_n20620, new_n20621, new_n20622, new_n20623, new_n20624, new_n20625,
    new_n20626, new_n20627, new_n20628, new_n20629, new_n20630, new_n20631,
    new_n20632, new_n20633, new_n20634, new_n20635, new_n20636, new_n20637,
    new_n20638, new_n20639, new_n20640, new_n20641, new_n20642, new_n20643,
    new_n20644, new_n20645, new_n20646, new_n20647, new_n20648, new_n20651,
    new_n20652, new_n20653, new_n20654, new_n20655, new_n20656, new_n20657,
    new_n20658, new_n20659, new_n20660, new_n20661, new_n20662, new_n20663,
    new_n20664, new_n20665, new_n20666, new_n20667, new_n20668, new_n20669,
    new_n20670, new_n20671, new_n20672, new_n20673, new_n20674, new_n20675,
    new_n20676, new_n20677, new_n20678, new_n20679, new_n20680, new_n20681,
    new_n20682, new_n20683, new_n20684, new_n20685, new_n20686, new_n20687,
    new_n20688, new_n20689, new_n20690, new_n20691, new_n20692, new_n20693,
    new_n20694, new_n20695, new_n20696, new_n20697, new_n20698, new_n20699,
    new_n20700, new_n20701, new_n20702, new_n20703, new_n20704, new_n20705,
    new_n20706, new_n20707, new_n20708, new_n20709, new_n20710, new_n20711,
    new_n20712, new_n20713, new_n20714, new_n20715, new_n20716, new_n20717,
    new_n20718, new_n20719, new_n20720, new_n20721, new_n20722, new_n20723,
    new_n20724, new_n20725, new_n20726, new_n20727, new_n20728, new_n20729,
    new_n20730, new_n20731, new_n20732, new_n20733, new_n20734, new_n20735,
    new_n20736, new_n20737, new_n20738, new_n20739, new_n20740, new_n20741,
    new_n20746, new_n20747, new_n20748, new_n20749, new_n20750, new_n20751,
    new_n20752, new_n20753, new_n20754, new_n20755, new_n20756, new_n20757,
    new_n20758, new_n20759, new_n20760, new_n20761, new_n20762, new_n20763,
    new_n20764, new_n20765, new_n20766, new_n20767, new_n20768, new_n20769,
    new_n20770, new_n20771, new_n20772, new_n20773, new_n20774, new_n20775,
    new_n20776, new_n20777, new_n20778, new_n20779, new_n20780, new_n20781,
    new_n20782, new_n20783, new_n20784, new_n20785, new_n20786, new_n20787,
    new_n20788, new_n20789, new_n20790, new_n20791, new_n20792, new_n20793,
    new_n20794, new_n20795, new_n20796, new_n20797, new_n20798, new_n20799,
    new_n20800, new_n20801, new_n20802, new_n20803, new_n20804, new_n20805,
    new_n20806, new_n20807, new_n20808, new_n20809, new_n20810, new_n20811,
    new_n20812, new_n20813, new_n20814, new_n20815, new_n20816, new_n20817,
    new_n20818, new_n20819, new_n20820, new_n20821, new_n20822, new_n20823,
    new_n20824, new_n20825, new_n20826, new_n20827, new_n20828, new_n20829,
    new_n20830, new_n20831, new_n20832, new_n20833, new_n20834, new_n20835,
    new_n20836, new_n20837, new_n20838, new_n20839, new_n20840, new_n20841,
    new_n20842, new_n20843, new_n20844, new_n20845, new_n20846, new_n20848,
    new_n20849, new_n20850, new_n20851, new_n20852, new_n20853, new_n20854,
    new_n20855, new_n20857, new_n20858, new_n20859, new_n20860, new_n20861,
    new_n20862, new_n20863, new_n20864, new_n20865, new_n20866, new_n20867,
    new_n20868, new_n20869, new_n20870, new_n20871, new_n20872, new_n20873,
    new_n20874, new_n20875, new_n20876, new_n20877, new_n20878, new_n20879,
    new_n20880, new_n20881, new_n20883, new_n20885, new_n20890, new_n20891,
    new_n20892, new_n20893, new_n20894, new_n20895, new_n20896, new_n20897,
    new_n20898, new_n20899, new_n20900, new_n20901, new_n20902, new_n20903,
    new_n20904, new_n20905, new_n20906, new_n20907, new_n20908, new_n20918,
    new_n20921, new_n20922, new_n20923, new_n20924, new_n20925, new_n20926,
    new_n20927, new_n20928, new_n20929, new_n20930, new_n20931, new_n20932,
    new_n20933, new_n20934, new_n20935, new_n20936, new_n20937, new_n20938,
    new_n20939, new_n20940, new_n20941, new_n20942, new_n20943, new_n20944,
    new_n20945, new_n20946, new_n20947, new_n20948, new_n20949, new_n20950,
    new_n20951, new_n20953, new_n20954, new_n20955, new_n20956, new_n20957,
    new_n20958, new_n20959, new_n20960, new_n20961, new_n20962, new_n20963,
    new_n20964, new_n20965, new_n20966, new_n20967, new_n20968, new_n20969,
    new_n20970, new_n20971, new_n20972, new_n20973, new_n20974, new_n20975,
    new_n20976, new_n20977, new_n20978, new_n20979, new_n20980, new_n20981,
    new_n20982, new_n20983, new_n20984, new_n20985, new_n20986, new_n20987,
    new_n20988, new_n20989, new_n20990, new_n20991, new_n20992, new_n20993,
    new_n20994, new_n20995, new_n20997, new_n20998, new_n20999, new_n21000,
    new_n21001, new_n21002, new_n21003, new_n21004, new_n21005, new_n21006,
    new_n21007, new_n21008, new_n21009, new_n21010, new_n21011, new_n21012,
    new_n21013, new_n21014, new_n21015, new_n21016, new_n21017, new_n21018,
    new_n21019, new_n21020, new_n21021, new_n21022, new_n21023, new_n21024,
    new_n21025, new_n21026, new_n21027, new_n21028, new_n21029, new_n21030,
    new_n21031, new_n21032, new_n21033, new_n21034, new_n21035, new_n21036,
    new_n21037, new_n21038, new_n21039, new_n21040, new_n21041, new_n21042,
    new_n21043, new_n21044, new_n21045, new_n21046, new_n21047, new_n21048,
    new_n21049, new_n21050, new_n21051, new_n21052, new_n21053, new_n21054,
    new_n21055, new_n21056, new_n21057, new_n21058, new_n21059, new_n21060,
    new_n21061, new_n21062, new_n21063, new_n21064, new_n21065, new_n21066,
    new_n21067, new_n21068, new_n21069, new_n21070, new_n21071, new_n21072,
    new_n21073, new_n21074, new_n21075, new_n21076, new_n21077, new_n21078,
    new_n21079, new_n21080, new_n21081, new_n21082, new_n21083, new_n21084,
    new_n21085, new_n21086, new_n21087, new_n21088, new_n21089, new_n21090,
    new_n21091, new_n21092, new_n21093, new_n21094, new_n21095, new_n21096,
    new_n21097, new_n21098, new_n21099, new_n21100, new_n21101, new_n21102,
    new_n21103, new_n21104, new_n21105, new_n21106, new_n21107, new_n21108,
    new_n21109, new_n21110, new_n21111, new_n21112, new_n21113, new_n21114,
    new_n21115, new_n21116, new_n21117, new_n21118, new_n21119, new_n21120,
    new_n21121, new_n21122, new_n21123, new_n21124, new_n21125, new_n21126,
    new_n21127, new_n21128, new_n21129, new_n21130, new_n21131, new_n21132,
    new_n21133, new_n21134, new_n21135, new_n21136, new_n21137, new_n21138,
    new_n21139, new_n21140, new_n21141, new_n21142, new_n21143, new_n21144,
    new_n21145, new_n21146, new_n21147, new_n21148, new_n21149, new_n21150,
    new_n21151, new_n21152, new_n21153, new_n21154, new_n21155, new_n21156,
    new_n21157, new_n21158, new_n21159, new_n21160, new_n21161, new_n21162,
    new_n21163, new_n21164, new_n21165, new_n21166, new_n21167, new_n21168,
    new_n21169, new_n21170, new_n21171, new_n21172, new_n21173, new_n21174,
    new_n21175, new_n21176, new_n21177, new_n21178, new_n21179, new_n21180,
    new_n21181, new_n21182, new_n21183, new_n21184, new_n21185, new_n21186,
    new_n21187, new_n21188, new_n21189, new_n21190, new_n21191, new_n21192,
    new_n21193, new_n21194, new_n21195, new_n21196, new_n21197, new_n21198,
    new_n21199, new_n21200, new_n21201, new_n21202, new_n21203, new_n21204,
    new_n21205, new_n21206, new_n21207, new_n21212, new_n21213, new_n21214,
    new_n21215, new_n21216, new_n21217, new_n21218, new_n21219, new_n21220,
    new_n21221, new_n21222, new_n21223, new_n21224, new_n21225, new_n21226,
    new_n21227, new_n21228, new_n21229, new_n21230, new_n21231, new_n21232,
    new_n21233, new_n21234, new_n21235, new_n21236, new_n21237, new_n21238,
    new_n21241, new_n21242, new_n21243, new_n21244, new_n21245, new_n21246,
    new_n21247, new_n21248, new_n21249, new_n21250, new_n21251, new_n21252,
    new_n21253, new_n21254, new_n21255, new_n21256, new_n21257, new_n21258,
    new_n21259, new_n21260, new_n21261, new_n21262, new_n21263, new_n21264,
    new_n21265, new_n21266, new_n21269, new_n21270, new_n21271, new_n21272,
    new_n21273, new_n21274, new_n21275, new_n21276, new_n21277, new_n21282,
    new_n21283, new_n21284, new_n21288, new_n21289, new_n21290, new_n21291,
    new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297,
    new_n21298, new_n21299, new_n21300, new_n21301, new_n21302, new_n21303,
    new_n21304, new_n21305, new_n21309, new_n21310, new_n21311, new_n21312,
    new_n21313, new_n21314, new_n21315, new_n21316, new_n21317, new_n21318,
    new_n21319, new_n21321, new_n21322, new_n21323, new_n21324, new_n21325,
    new_n21326, new_n21327, new_n21328, new_n21329, new_n21330, new_n21331,
    new_n21332, new_n21333, new_n21334, new_n21335, new_n21336, new_n21337,
    new_n21338, new_n21339, new_n21340, new_n21341, new_n21342, new_n21344,
    new_n21345, new_n21346, new_n21347, new_n21348, new_n21349, new_n21350,
    new_n21351, new_n21352, new_n21353, new_n21354, new_n21355, new_n21356,
    new_n21357, new_n21358, new_n21359, new_n21360, new_n21361, new_n21362,
    new_n21363, new_n21364, new_n21365, new_n21366, new_n21367, new_n21368,
    new_n21369, new_n21370, new_n21371, new_n21372, new_n21373, new_n21374,
    new_n21375, new_n21376, new_n21377, new_n21378, new_n21379, new_n21380,
    new_n21381, new_n21382, new_n21383, new_n21385, new_n21386, new_n21387,
    new_n21388, new_n21389, new_n21390, new_n21391, new_n21392, new_n21393,
    new_n21394, new_n21395, new_n21396, new_n21397, new_n21398, new_n21399,
    new_n21400, new_n21401, new_n21402, new_n21403, new_n21404, new_n21405,
    new_n21406, new_n21407, new_n21408, new_n21409, new_n21410, new_n21411,
    new_n21412, new_n21413, new_n21414, new_n21415, new_n21416, new_n21417,
    new_n21418, new_n21419, new_n21420, new_n21421, new_n21422, new_n21423,
    new_n21424, new_n21425, new_n21426, new_n21427, new_n21428, new_n21429,
    new_n21430, new_n21431, new_n21432, new_n21433, new_n21434, new_n21435,
    new_n21436, new_n21437, new_n21438, new_n21439, new_n21440, new_n21441,
    new_n21442, new_n21443, new_n21444, new_n21445, new_n21446, new_n21447,
    new_n21448, new_n21449, new_n21450, new_n21451, new_n21452, new_n21453,
    new_n21454, new_n21455, new_n21456, new_n21457, new_n21458, new_n21459,
    new_n21460, new_n21461, new_n21462, new_n21463, new_n21464, new_n21469,
    new_n21470, new_n21471, new_n21472, new_n21473, new_n21474, new_n21475,
    new_n21476, new_n21477, new_n21478, new_n21479, new_n21480, new_n21481,
    new_n21482, new_n21483, new_n21484, new_n21485, new_n21486, new_n21487,
    new_n21488, new_n21489, new_n21490, new_n21491, new_n21492, new_n21493,
    new_n21494, new_n21495, new_n21496, new_n21497, new_n21498, new_n21499,
    new_n21500, new_n21501, new_n21502, new_n21503, new_n21504, new_n21505,
    new_n21506, new_n21507, new_n21508, new_n21509, new_n21510, new_n21511,
    new_n21512, new_n21513, new_n21514, new_n21515, new_n21516, new_n21517,
    new_n21518, new_n21519, new_n21520, new_n21521, new_n21522, new_n21523,
    new_n21524, new_n21525, new_n21526, new_n21527, new_n21528, new_n21529,
    new_n21530, new_n21531, new_n21532, new_n21533, new_n21534, new_n21535,
    new_n21536, new_n21537, new_n21538, new_n21539, new_n21540, new_n21541,
    new_n21542, new_n21543, new_n21544, new_n21545, new_n21546, new_n21547,
    new_n21548, new_n21549, new_n21550, new_n21551, new_n21552, new_n21553,
    new_n21554, new_n21555, new_n21556, new_n21557, new_n21558, new_n21559,
    new_n21560, new_n21561, new_n21562, new_n21563, new_n21564, new_n21565,
    new_n21566, new_n21567, new_n21568, new_n21569, new_n21570, new_n21571,
    new_n21572, new_n21573, new_n21574, new_n21575, new_n21576, new_n21577,
    new_n21578, new_n21579, new_n21580, new_n21581, new_n21582, new_n21583,
    new_n21584, new_n21585, new_n21586, new_n21587, new_n21588, new_n21589,
    new_n21590, new_n21591, new_n21592, new_n21593, new_n21594, new_n21595,
    new_n21596, new_n21597, new_n21598, new_n21600, new_n21601, new_n21607,
    new_n21608, new_n21609, new_n21610, new_n21611, new_n21612, new_n21613,
    new_n21614, new_n21615, new_n21616, new_n21617, new_n21618, new_n21619,
    new_n21620, new_n21621, new_n21622, new_n21623, new_n21624, new_n21625,
    new_n21626, new_n21627, new_n21628, new_n21629, new_n21630, new_n21631,
    new_n21632, new_n21633, new_n21634, new_n21635, new_n21636, new_n21637,
    new_n21638, new_n21639, new_n21640, new_n21641, new_n21642, new_n21643,
    new_n21644, new_n21645, new_n21646, new_n21647, new_n21649, new_n21650,
    new_n21651, new_n21652, new_n21653, new_n21654, new_n21655, new_n21656,
    new_n21657, new_n21658, new_n21659, new_n21660, new_n21661, new_n21662,
    new_n21663, new_n21664, new_n21665, new_n21666, new_n21667, new_n21668,
    new_n21669, new_n21670, new_n21671, new_n21672, new_n21673, new_n21674,
    new_n21675, new_n21676, new_n21677, new_n21678, new_n21679, new_n21680,
    new_n21681, new_n21682, new_n21683, new_n21684, new_n21685, new_n21686,
    new_n21695, new_n21696, new_n21697, new_n21698, new_n21699, new_n21700,
    new_n21701, new_n21702, new_n21703, new_n21704, new_n21705, new_n21706,
    new_n21707, new_n21708, new_n21709, new_n21713, new_n21714, new_n21715,
    new_n21716, new_n21717, new_n21718, new_n21719, new_n21720, new_n21721,
    new_n21722, new_n21723, new_n21724, new_n21725, new_n21726, new_n21727,
    new_n21728, new_n21729, new_n21730, new_n21731, new_n21732, new_n21733,
    new_n21734, new_n21735, new_n21736, new_n21737, new_n21738, new_n21739,
    new_n21740, new_n21741, new_n21742, new_n21743, new_n21744, new_n21745,
    new_n21746, new_n21747, new_n21750, new_n21751, new_n21752, new_n21753,
    new_n21754, new_n21755, new_n21756, new_n21757, new_n21758, new_n21759,
    new_n21760, new_n21761, new_n21762, new_n21763, new_n21764, new_n21765,
    new_n21766, new_n21767, new_n21768, new_n21769, new_n21770, new_n21771,
    new_n21772, new_n21773, new_n21774, new_n21775, new_n21776, new_n21777,
    new_n21778, new_n21779, new_n21780, new_n21781, new_n21782, new_n21783,
    new_n21784, new_n21785, new_n21786, new_n21787, new_n21788, new_n21789,
    new_n21790, new_n21791, new_n21792, new_n21793, new_n21794, new_n21795,
    new_n21796, new_n21797, new_n21798, new_n21799, new_n21800, new_n21801,
    new_n21802, new_n21803, new_n21804, new_n21805, new_n21806, new_n21807,
    new_n21808, new_n21809, new_n21810, new_n21811, new_n21812, new_n21813,
    new_n21814, new_n21815, new_n21816, new_n21817, new_n21818, new_n21820,
    new_n21821, new_n21822, new_n21823, new_n21824, new_n21825, new_n21826,
    new_n21827, new_n21828, new_n21829, new_n21830, new_n21831, new_n21832,
    new_n21833, new_n21834, new_n21835, new_n21836, new_n21837, new_n21838,
    new_n21839, new_n21840, new_n21841, new_n21842, new_n21843, new_n21844,
    new_n21845, new_n21846, new_n21847, new_n21848, new_n21850, new_n21851,
    new_n21853, new_n21854, new_n21855, new_n21856, new_n21857, new_n21858,
    new_n21859, new_n21860, new_n21861, new_n21862, new_n21863, new_n21864,
    new_n21865, new_n21866, new_n21867, new_n21868, new_n21869, new_n21870,
    new_n21871, new_n21872, new_n21873, new_n21874, new_n21875, new_n21876,
    new_n21877, new_n21878, new_n21879, new_n21880, new_n21881, new_n21882,
    new_n21883, new_n21884, new_n21885, new_n21886, new_n21887, new_n21888,
    new_n21891, new_n21892, new_n21895, new_n21896, new_n21897, new_n21898,
    new_n21899, new_n21900, new_n21901, new_n21902, new_n21903, new_n21904,
    new_n21905, new_n21906, new_n21907, new_n21908, new_n21909, new_n21910,
    new_n21911, new_n21912, new_n21913, new_n21914, new_n21915, new_n21916,
    new_n21917, new_n21918, new_n21919, new_n21920, new_n21921, new_n21922,
    new_n21923, new_n21924, new_n21925, new_n21926, new_n21927, new_n21928,
    new_n21929, new_n21930, new_n21931, new_n21932, new_n21933, new_n21934,
    new_n21935, new_n21936, new_n21937, new_n21938, new_n21939, new_n21940,
    new_n21941, new_n21944, new_n21945, new_n21946, new_n21947, new_n21948,
    new_n21949, new_n21950, new_n21951, new_n21952, new_n21953, new_n21954,
    new_n21955, new_n21956, new_n21957, new_n21958, new_n21959, new_n21960,
    new_n21961, new_n21962, new_n21963, new_n21964, new_n21972, new_n21973,
    new_n21974, new_n21975, new_n21976, new_n21977, new_n21978, new_n21979,
    new_n21980, new_n21981, new_n21982, new_n21983, new_n21984, new_n21985,
    new_n21986, new_n21987, new_n21988, new_n21989, new_n21990, new_n21991,
    new_n21992, new_n21993, new_n21994, new_n21995, new_n21996, new_n21997,
    new_n21998, new_n21999, new_n22000, new_n22001, new_n22002, new_n22003,
    new_n22004, new_n22005, new_n22006, new_n22007, new_n22008, new_n22009,
    new_n22010, new_n22011, new_n22012, new_n22013, new_n22014, new_n22015,
    new_n22016, new_n22017, new_n22018, new_n22019, new_n22020, new_n22021,
    new_n22022, new_n22023, new_n22024, new_n22025, new_n22027, new_n22029,
    new_n22038, new_n22039, new_n22040, new_n22041, new_n22042, new_n22047,
    new_n22048, new_n22049, new_n22050, new_n22051, new_n22052, new_n22053,
    new_n22054, new_n22055, new_n22056, new_n22057, new_n22058, new_n22061,
    new_n22067, new_n22073, new_n22074, new_n22075, new_n22076, new_n22077,
    new_n22078, new_n22079, new_n22080, new_n22081, new_n22082, new_n22083,
    new_n22084, new_n22085, new_n22086, new_n22087, new_n22088, new_n22089,
    new_n22090, new_n22091, new_n22092, new_n22093, new_n22094, new_n22095,
    new_n22096, new_n22097, new_n22098, new_n22099, new_n22100, new_n22101,
    new_n22102, new_n22103, new_n22104, new_n22105, new_n22106, new_n22107,
    new_n22109, new_n22110, new_n22111, new_n22112, new_n22113, new_n22114,
    new_n22115, new_n22116, new_n22117, new_n22118, new_n22119, new_n22120,
    new_n22121, new_n22122, new_n22123, new_n22124, new_n22125, new_n22127,
    new_n22128, new_n22129, new_n22130, new_n22131, new_n22132, new_n22133,
    new_n22134, new_n22135, new_n22136, new_n22137, new_n22138, new_n22139,
    new_n22140, new_n22145, new_n22146, new_n22147, new_n22148, new_n22149,
    new_n22150, new_n22151, new_n22152, new_n22153, new_n22154, new_n22155,
    new_n22156, new_n22157, new_n22158, new_n22159, new_n22160, new_n22161,
    new_n22162, new_n22163, new_n22166, new_n22173, new_n22174, new_n22175,
    new_n22176, new_n22177, new_n22178, new_n22179, new_n22180, new_n22185,
    new_n22186, new_n22187, new_n22188, new_n22189, new_n22190, new_n22194,
    new_n22201, new_n22202, new_n22203, new_n22204, new_n22205, new_n22206,
    new_n22207, new_n22208, new_n22209, new_n22210, new_n22211, new_n22212,
    new_n22213, new_n22214, new_n22215, new_n22216, new_n22217, new_n22218,
    new_n22219, new_n22220, new_n22221, new_n22222, new_n22225, new_n22228,
    new_n22229, new_n22230, new_n22231, new_n22233, new_n22239, new_n22240,
    new_n22241, new_n22242, new_n22243, new_n22244, new_n22245, new_n22246,
    new_n22247, new_n22248, new_n22249, new_n22250, new_n22251, new_n22252,
    new_n22253, new_n22254, new_n22255, new_n22256, new_n22257, new_n22258,
    new_n22259, new_n22260, new_n22261, new_n22262, new_n22263, new_n22264,
    new_n22265, new_n22266, new_n22267, new_n22268, new_n22269, new_n22270,
    new_n22271, new_n22272, new_n22273, new_n22274, new_n22275, new_n22276,
    new_n22277, new_n22278, new_n22279, new_n22280, new_n22281, new_n22282,
    new_n22283, new_n22284, new_n22285, new_n22286, new_n22289, new_n22290,
    new_n22291, new_n22292, new_n22293, new_n22294, new_n22295, new_n22296,
    new_n22297, new_n22298, new_n22299, new_n22300, new_n22301, new_n22303,
    new_n22304, new_n22305, new_n22306, new_n22307, new_n22308, new_n22309,
    new_n22310, new_n22311, new_n22312, new_n22313, new_n22314, new_n22315,
    new_n22316, new_n22317, new_n22318, new_n22319, new_n22320, new_n22321,
    new_n22322, new_n22323, new_n22326, new_n22328, new_n22331, new_n22336,
    new_n22337, new_n22338, new_n22339, new_n22340, new_n22341, new_n22342,
    new_n22343, new_n22344, new_n22345, new_n22346, new_n22347, new_n22348,
    new_n22349, new_n22350, new_n22351, new_n22352, new_n22353, new_n22354,
    new_n22355, new_n22356, new_n22357, new_n22358, new_n22359, new_n22360,
    new_n22361, new_n22362, new_n22363, new_n22364, new_n22365, new_n22366,
    new_n22367, new_n22368, new_n22369, new_n22375, new_n22376, new_n22377,
    new_n22378, new_n22388, new_n22389, new_n22390, new_n22391, new_n22392,
    new_n22393, new_n22394, new_n22395, new_n22396, new_n22397, new_n22398,
    new_n22399, new_n22400, new_n22401, new_n22402, new_n22403, new_n22404,
    new_n22405, new_n22406, new_n22407, new_n22408, new_n22409, new_n22410,
    new_n22411, new_n22412, new_n22413, new_n22414, new_n22415, new_n22416,
    new_n22417, new_n22418, new_n22419, new_n22420, new_n22421, new_n22422,
    new_n22423, new_n22424, new_n22425, new_n22426, new_n22427, new_n22428,
    new_n22429, new_n22430, new_n22431, new_n22432, new_n22433, new_n22434,
    new_n22435, new_n22436, new_n22437, new_n22438, new_n22439, new_n22440,
    new_n22441, new_n22442, new_n22443, new_n22444, new_n22445, new_n22446,
    new_n22447, new_n22448, new_n22449, new_n22450, new_n22451, new_n22452,
    new_n22453, new_n22454, new_n22455, new_n22456, new_n22457, new_n22458,
    new_n22459, new_n22460, new_n22461, new_n22462, new_n22464, new_n22465,
    new_n22466, new_n22467, new_n22468, new_n22469, new_n22470, new_n22471,
    new_n22472, new_n22473, new_n22474, new_n22475, new_n22476, new_n22477,
    new_n22478, new_n22479, new_n22480, new_n22481, new_n22482, new_n22483,
    new_n22484, new_n22485, new_n22486, new_n22487, new_n22488, new_n22489,
    new_n22490, new_n22491, new_n22492, new_n22493, new_n22494, new_n22495,
    new_n22496, new_n22497, new_n22498, new_n22499, new_n22500, new_n22501,
    new_n22502, new_n22503, new_n22504, new_n22505, new_n22506, new_n22507,
    new_n22508, new_n22509, new_n22510, new_n22511, new_n22512, new_n22513,
    new_n22514, new_n22515, new_n22516, new_n22517, new_n22518, new_n22519,
    new_n22520, new_n22521, new_n22522, new_n22523, new_n22524, new_n22525,
    new_n22526, new_n22527, new_n22528, new_n22529, new_n22530, new_n22531,
    new_n22532, new_n22533, new_n22534, new_n22535, new_n22536, new_n22539,
    new_n22540, new_n22541, new_n22542, new_n22543, new_n22544, new_n22545,
    new_n22546, new_n22547, new_n22548, new_n22549, new_n22550, new_n22551,
    new_n22552, new_n22553, new_n22556, new_n22560, new_n22561, new_n22562,
    new_n22563, new_n22564, new_n22565, new_n22566, new_n22567, new_n22568,
    new_n22569, new_n22570, new_n22571, new_n22572, new_n22573, new_n22574,
    new_n22575, new_n22576, new_n22577, new_n22578, new_n22579, new_n22580,
    new_n22581, new_n22582, new_n22583, new_n22584, new_n22585, new_n22586,
    new_n22587, new_n22588, new_n22589, new_n22590, new_n22591, new_n22592,
    new_n22593, new_n22594, new_n22595, new_n22596, new_n22597, new_n22598,
    new_n22599, new_n22600, new_n22601, new_n22602, new_n22603, new_n22604,
    new_n22605, new_n22606, new_n22607, new_n22608, new_n22609, new_n22610,
    new_n22611, new_n22612, new_n22613, new_n22614, new_n22615, new_n22616,
    new_n22617, new_n22618, new_n22619, new_n22620, new_n22621, new_n22622,
    new_n22623, new_n22624, new_n22625, new_n22626, new_n22627, new_n22628,
    new_n22629, new_n22630, new_n22631, new_n22632, new_n22633, new_n22634,
    new_n22635, new_n22636, new_n22638, new_n22639, new_n22640, new_n22641,
    new_n22642, new_n22643, new_n22644, new_n22645, new_n22646, new_n22647,
    new_n22650, new_n22651, new_n22652, new_n22653, new_n22654, new_n22655,
    new_n22656, new_n22657, new_n22658, new_n22660, new_n22661, new_n22666,
    new_n22667, new_n22668, new_n22669, new_n22670, new_n22671, new_n22672,
    new_n22673, new_n22674, new_n22675, new_n22676, new_n22677, new_n22678,
    new_n22679, new_n22680, new_n22681, new_n22682, new_n22683, new_n22684,
    new_n22685, new_n22686, new_n22687, new_n22688, new_n22689, new_n22690,
    new_n22691, new_n22692, new_n22693, new_n22694, new_n22695, new_n22696,
    new_n22697, new_n22698, new_n22699, new_n22700, new_n22701, new_n22702,
    new_n22703, new_n22704, new_n22705, new_n22706, new_n22707, new_n22708,
    new_n22709, new_n22710, new_n22711, new_n22712, new_n22713, new_n22714,
    new_n22715, new_n22716, new_n22717, new_n22718, new_n22719, new_n22720,
    new_n22721, new_n22722, new_n22723, new_n22724, new_n22725, new_n22726,
    new_n22727, new_n22728, new_n22729, new_n22730, new_n22731, new_n22732,
    new_n22733, new_n22734, new_n22735, new_n22736, new_n22737, new_n22738,
    new_n22739, new_n22740, new_n22748, new_n22749, new_n22750, new_n22751,
    new_n22752, new_n22753, new_n22754, new_n22759, new_n22763, new_n22764,
    new_n22765, new_n22766, new_n22767, new_n22768, new_n22769, new_n22770,
    new_n22771, new_n22772, new_n22773, new_n22774, new_n22775, new_n22776,
    new_n22777, new_n22778, new_n22779, new_n22780, new_n22781, new_n22782,
    new_n22783, new_n22784, new_n22785, new_n22786, new_n22787, new_n22788,
    new_n22789, new_n22790, new_n22791, new_n22792, new_n22793, new_n22794,
    new_n22795, new_n22796, new_n22797, new_n22798, new_n22799, new_n22800,
    new_n22801, new_n22802, new_n22803, new_n22804, new_n22805, new_n22806,
    new_n22807, new_n22808, new_n22811, new_n22812, new_n22813, new_n22819,
    new_n22821, new_n22823, new_n22824, new_n22825, new_n22826, new_n22827,
    new_n22828, new_n22829, new_n22830, new_n22831, new_n22832, new_n22836,
    new_n22844, new_n22845, new_n22846, new_n22847, new_n22848, new_n22849,
    new_n22850, new_n22851, new_n22852, new_n22853, new_n22854, new_n22855,
    new_n22856, new_n22857, new_n22858, new_n22859, new_n22860, new_n22861,
    new_n22862, new_n22863, new_n22864, new_n22865, new_n22866, new_n22867,
    new_n22868, new_n22869, new_n22870, new_n22871, new_n22873, new_n22874,
    new_n22875, new_n22876, new_n22877, new_n22878, new_n22879, new_n22880,
    new_n22881, new_n22882, new_n22883, new_n22884, new_n22885, new_n22886,
    new_n22887, new_n22888, new_n22889, new_n22890, new_n22896, new_n22897,
    new_n22898, new_n22899, new_n22900, new_n22901, new_n22902, new_n22903,
    new_n22904, new_n22905, new_n22906, new_n22907, new_n22908, new_n22909,
    new_n22910, new_n22911, new_n22912, new_n22913, new_n22914, new_n22915,
    new_n22916, new_n22917, new_n22918, new_n22919, new_n22920, new_n22921,
    new_n22922, new_n22923, new_n22924, new_n22925, new_n22928, new_n22929,
    new_n22930, new_n22931, new_n22932, new_n22933, new_n22934, new_n22935,
    new_n22936, new_n22937, new_n22938, new_n22939, new_n22940, new_n22941,
    new_n22942, new_n22943, new_n22944, new_n22945, new_n22946, new_n22947,
    new_n22948, new_n22949, new_n22950, new_n22951, new_n22952, new_n22953,
    new_n22954, new_n22955, new_n22957, new_n22958, new_n22959, new_n22960,
    new_n22961, new_n22962, new_n22963, new_n22964, new_n22965, new_n22966,
    new_n22967, new_n22971, new_n22972, new_n22974, new_n22975, new_n22976,
    new_n22981, new_n22982, new_n22983, new_n22984, new_n22985, new_n22986,
    new_n22987, new_n22988, new_n22989, new_n22990, new_n22991, new_n22992,
    new_n22993, new_n22994, new_n22995, new_n22996, new_n22997, new_n22998,
    new_n22999, new_n23000, new_n23001, new_n23002, new_n23003, new_n23004,
    new_n23005, new_n23006, new_n23007, new_n23008, new_n23009, new_n23010,
    new_n23011, new_n23012, new_n23013, new_n23014, new_n23015, new_n23016,
    new_n23017, new_n23018, new_n23019, new_n23020, new_n23021, new_n23022,
    new_n23023, new_n23024, new_n23026, new_n23027, new_n23028, new_n23029,
    new_n23030, new_n23031, new_n23032, new_n23033, new_n23034, new_n23035,
    new_n23036, new_n23037, new_n23038, new_n23039, new_n23040, new_n23041,
    new_n23042, new_n23043, new_n23044, new_n23045, new_n23046, new_n23047,
    new_n23048, new_n23049, new_n23050, new_n23051, new_n23052, new_n23053,
    new_n23054, new_n23055, new_n23056, new_n23057, new_n23058, new_n23059,
    new_n23060, new_n23061, new_n23062, new_n23063, new_n23064, new_n23065,
    new_n23066, new_n23067, new_n23068, new_n23069, new_n23070, new_n23071,
    new_n23075, new_n23080, new_n23087, new_n23088, new_n23089, new_n23090,
    new_n23095, new_n23097, new_n23104, new_n23105, new_n23106, new_n23107,
    new_n23108, new_n23109, new_n23110, new_n23111, new_n23112, new_n23113,
    new_n23114, new_n23115, new_n23116, new_n23117, new_n23118, new_n23119,
    new_n23120, new_n23121, new_n23122, new_n23123, new_n23124, new_n23125,
    new_n23126, new_n23127, new_n23128, new_n23129, new_n23130, new_n23131,
    new_n23132, new_n23133, new_n23134, new_n23135, new_n23136, new_n23137,
    new_n23138, new_n23139, new_n23140, new_n23141, new_n23142, new_n23143,
    new_n23144, new_n23145, new_n23148, new_n23149, new_n23150, new_n23151,
    new_n23152, new_n23153, new_n23154, new_n23155, new_n23156, new_n23157,
    new_n23158, new_n23159, new_n23160, new_n23164, new_n23168, new_n23169,
    new_n23170, new_n23171, new_n23172, new_n23173, new_n23174, new_n23175,
    new_n23176, new_n23177, new_n23178, new_n23179, new_n23180, new_n23181,
    new_n23182, new_n23183, new_n23184, new_n23185, new_n23186, new_n23187,
    new_n23188, new_n23189, new_n23190, new_n23191, new_n23192, new_n23193,
    new_n23194, new_n23195, new_n23196, new_n23197, new_n23198, new_n23199,
    new_n23200, new_n23201, new_n23202, new_n23203, new_n23204, new_n23205,
    new_n23206, new_n23207, new_n23208, new_n23209, new_n23210, new_n23211,
    new_n23212, new_n23213, new_n23214, new_n23215, new_n23216, new_n23217,
    new_n23218, new_n23219, new_n23220, new_n23221, new_n23222, new_n23223,
    new_n23224, new_n23225, new_n23226, new_n23227, new_n23228, new_n23229,
    new_n23230, new_n23231, new_n23232, new_n23233, new_n23234, new_n23235,
    new_n23236, new_n23237, new_n23238, new_n23239, new_n23240, new_n23241,
    new_n23242, new_n23243, new_n23244, new_n23245, new_n23246, new_n23247,
    new_n23248, new_n23249, new_n23250, new_n23251, new_n23252, new_n23253,
    new_n23254, new_n23255, new_n23256, new_n23257, new_n23258, new_n23259,
    new_n23260, new_n23261, new_n23262, new_n23263, new_n23264, new_n23265,
    new_n23266, new_n23267, new_n23268, new_n23269, new_n23270, new_n23271,
    new_n23272, new_n23273, new_n23274, new_n23275, new_n23276, new_n23277,
    new_n23278, new_n23279, new_n23280, new_n23281, new_n23282, new_n23283,
    new_n23284, new_n23285, new_n23286, new_n23287, new_n23288, new_n23289,
    new_n23290, new_n23291, new_n23292, new_n23293, new_n23294, new_n23295,
    new_n23296, new_n23297, new_n23298, new_n23299, new_n23300, new_n23301,
    new_n23302, new_n23303, new_n23304, new_n23305, new_n23306, new_n23307,
    new_n23308, new_n23309, new_n23310, new_n23311, new_n23312, new_n23316,
    new_n23319, new_n23320, new_n23321, new_n23322, new_n23323, new_n23324,
    new_n23325, new_n23326, new_n23327, new_n23328, new_n23329, new_n23330,
    new_n23331, new_n23332, new_n23333, new_n23334, new_n23338, new_n23340,
    new_n23341, new_n23342, new_n23343, new_n23344, new_n23345, new_n23346,
    new_n23347, new_n23348, new_n23349, new_n23350, new_n23351, new_n23352,
    new_n23353, new_n23354, new_n23355, new_n23356, new_n23357, new_n23358,
    new_n23359, new_n23360, new_n23361, new_n23362, new_n23363, new_n23365,
    new_n23366, new_n23367, new_n23368, new_n23372, new_n23373, new_n23374,
    new_n23375, new_n23376, new_n23386, new_n23387, new_n23388, new_n23389,
    new_n23390, new_n23391, new_n23392, new_n23393, new_n23394, new_n23395,
    new_n23396, new_n23397, new_n23398, new_n23399, new_n23400, new_n23401,
    new_n23402, new_n23403, new_n23404, new_n23405, new_n23418, new_n23422,
    new_n23428, new_n23429, new_n23430, new_n23431, new_n23432, new_n23433,
    new_n23434, new_n23435, new_n23436, new_n23437, new_n23438, new_n23439,
    new_n23440, new_n23441, new_n23442, new_n23443, new_n23444, new_n23445,
    new_n23446, new_n23447, new_n23448, new_n23449, new_n23450, new_n23451,
    new_n23452, new_n23453, new_n23454, new_n23455, new_n23456, new_n23457,
    new_n23458, new_n23459, new_n23460, new_n23461, new_n23462, new_n23463,
    new_n23464, new_n23465, new_n23466, new_n23467, new_n23471, new_n23473,
    new_n23476, new_n23477, new_n23478, new_n23479, new_n23480, new_n23481,
    new_n23482, new_n23483, new_n23484, new_n23485, new_n23486, new_n23487,
    new_n23488, new_n23489, new_n23490, new_n23491, new_n23492, new_n23493,
    new_n23494, new_n23495, new_n23496, new_n23497, new_n23501, new_n23502,
    new_n23505, new_n23506, new_n23507, new_n23508, new_n23509, new_n23510,
    new_n23511, new_n23514, new_n23515, new_n23516, new_n23517, new_n23518,
    new_n23519, new_n23520, new_n23521, new_n23522, new_n23523, new_n23524,
    new_n23525, new_n23526, new_n23527, new_n23528, new_n23529, new_n23530,
    new_n23531, new_n23532, new_n23533, new_n23534, new_n23535, new_n23536,
    new_n23537, new_n23538, new_n23539, new_n23540, new_n23541, new_n23542,
    new_n23543, new_n23544, new_n23545, new_n23546, new_n23547, new_n23548,
    new_n23549, new_n23552, new_n23553, new_n23554, new_n23555, new_n23556,
    new_n23557, new_n23558, new_n23559, new_n23560, new_n23561, new_n23562,
    new_n23563, new_n23564, new_n23565, new_n23566, new_n23567, new_n23568,
    new_n23569, new_n23570, new_n23571, new_n23572, new_n23573, new_n23574,
    new_n23575, new_n23576, new_n23577, new_n23578, new_n23579, new_n23580,
    new_n23581, new_n23582, new_n23583, new_n23584, new_n23585, new_n23586,
    new_n23587, new_n23588, new_n23589, new_n23590, new_n23591, new_n23592,
    new_n23605, new_n23610, new_n23612, new_n23616, new_n23620, new_n23621,
    new_n23622, new_n23623, new_n23624, new_n23625, new_n23626, new_n23627,
    new_n23628, new_n23629, new_n23630, new_n23631, new_n23632, new_n23633,
    new_n23634, new_n23635, new_n23638, new_n23639, new_n23640, new_n23641,
    new_n23642, new_n23643, new_n23644, new_n23645, new_n23646, new_n23647,
    new_n23648, new_n23649, new_n23650, new_n23651, new_n23652, new_n23653,
    new_n23654, new_n23655, new_n23656, new_n23657, new_n23661, new_n23662,
    new_n23663, new_n23664, new_n23665, new_n23666, new_n23667, new_n23668,
    new_n23669, new_n23677, new_n23678, new_n23679, new_n23680, new_n23681,
    new_n23682, new_n23683, new_n23685, new_n23686, new_n23687, new_n23688,
    new_n23689, new_n23690, new_n23691, new_n23692, new_n23693, new_n23694,
    new_n23695, new_n23696, new_n23697, new_n23698, new_n23699, new_n23700,
    new_n23701, new_n23702, new_n23703, new_n23704, new_n23722, new_n23728,
    new_n23729, new_n23730, new_n23731, new_n23732, new_n23733, new_n23734,
    new_n23735, new_n23736, new_n23737, new_n23738, new_n23739, new_n23740,
    new_n23741, new_n23742, new_n23743, new_n23744, new_n23745, new_n23746,
    new_n23751, new_n23752, new_n23753, new_n23754, new_n23762, new_n23772,
    new_n23783, new_n23784, new_n23785, new_n23786, new_n23787, new_n23788,
    new_n23789, new_n23792, new_n23804, new_n23805, new_n23806, new_n23810,
    new_n23811, new_n23812, new_n23813, new_n23814, new_n23815, new_n23816,
    new_n23817, new_n23822, new_n23823, new_n23824, new_n23825, new_n23826,
    new_n23827, new_n23829, new_n23830, new_n23831, new_n23833, new_n23834,
    new_n23838, new_n23850, new_n23851, new_n23852, new_n23855, new_n23856,
    new_n23864, new_n23865, new_n23868, new_n23871, new_n23876, new_n23877,
    new_n23887, new_n23888, new_n23889, new_n23890, new_n23891, new_n23892,
    new_n23893, new_n23895, new_n23897, new_n23899, new_n23902, new_n23903,
    new_n23904, new_n23905, new_n23906, new_n23907, new_n23908, new_n23909,
    new_n23913, new_n23914, new_n23915, new_n23916, new_n23917, new_n23918,
    new_n23920, new_n23921, new_n23927, new_n23931, new_n23932, new_n23933,
    new_n23936, new_n23937, new_n23939, new_n23940, new_n23941, new_n23942,
    new_n23943, new_n23944, new_n23945, new_n23946, new_n23947, new_n23948,
    new_n23949, new_n23950, new_n23951, new_n23952, new_n23953, new_n23954,
    new_n23955, new_n23960, new_n23974, new_n23975, new_n23976, new_n23977,
    new_n23978, new_n23979, new_n23980, new_n23981, new_n23982, new_n23983,
    new_n23984, new_n23985, new_n23986, new_n23989, new_n23990, new_n23991,
    new_n23996, new_n23997, new_n23998, new_n23999, new_n24000, new_n24002,
    new_n24006, new_n24007, new_n24008, new_n24009, new_n24010, new_n24011,
    new_n24012, new_n24013, new_n24014, new_n24015, new_n24016, new_n24018,
    new_n24019, new_n24020, new_n24021, new_n24022, new_n24023, new_n24024,
    new_n24025, new_n24026, new_n24027, new_n24028, new_n24029, new_n24030,
    new_n24031, new_n24032, new_n24033, new_n24034, new_n24035, new_n24036,
    new_n24037, new_n24038, new_n24039, new_n24040, new_n24041, new_n24042,
    new_n24043, new_n24044, new_n24045, new_n24046, new_n24047, new_n24048,
    new_n24050, new_n24051, new_n24052, new_n24053, new_n24054, new_n24055,
    new_n24056, new_n24057, new_n24058, new_n24059, new_n24060, new_n24061,
    new_n24062, new_n24063, new_n24064, new_n24065, new_n24066, new_n24068,
    new_n24070, new_n24071, new_n24072, new_n24073, new_n24074, new_n24075,
    new_n24076, new_n24087, new_n24091, new_n24092, new_n24093, new_n24107,
    new_n24110, new_n24111, new_n24112, new_n24113, new_n24114, new_n24115,
    new_n24122, new_n24124, new_n24125, new_n24126, new_n24127, new_n24128,
    new_n24129, new_n24130, new_n24137, new_n24150, new_n24151, new_n24152,
    new_n24154, new_n24165, new_n24168, new_n24174, new_n24178, new_n24179,
    new_n24183, new_n24185, new_n24186, new_n24187, new_n24188, new_n24189,
    new_n24190, new_n24191, new_n24192, new_n24202, new_n24203, new_n24204,
    new_n24218, new_n24219, new_n24220, new_n24221, new_n24222, new_n24223,
    new_n24229, new_n24230, new_n24231, new_n24232, new_n24233, new_n24234,
    new_n24235, new_n24236, new_n24237, new_n24240, new_n24241, new_n24242,
    new_n24243, new_n24249, new_n24250, new_n24251, new_n24253, new_n24254,
    new_n24255, new_n24256, new_n24257, new_n24258, new_n24259, new_n24260,
    new_n24261, new_n24262, new_n24263, new_n24264, new_n24265, new_n24266,
    new_n24269, new_n24274, new_n24279, new_n24281, new_n24291, new_n24301,
    new_n24305, new_n24309, new_n24310, new_n24314, new_n24315, new_n24318,
    new_n24323, new_n24326, new_n24329, new_n24335, new_n24336, new_n24349,
    new_n24358, new_n24359, new_n24360, new_n24361, new_n24362, new_n24363,
    new_n24364, new_n24365, new_n24366, new_n24367, new_n24368, new_n24383,
    new_n24384, new_n24385, new_n24386, new_n24387, new_n24388, new_n24389,
    new_n24390, new_n24391, new_n24400, new_n24402, new_n24403, new_n24404,
    new_n24405, new_n24406, new_n24407, new_n24408, new_n24409, new_n24410,
    new_n24411, new_n24417, new_n24419, new_n24421, new_n24424, new_n24427,
    new_n24429, new_n24430, new_n24431, new_n24439, new_n24440, new_n24441,
    new_n24445, new_n24449, new_n24450, new_n24456, new_n24463, new_n24465,
    new_n24466, new_n24467, new_n24470, new_n24473, new_n24474, new_n24475,
    new_n24486, new_n24488, new_n24489, new_n24490, new_n24492, new_n24499,
    new_n24503, new_n24505, new_n24506, new_n24508, new_n24514, new_n24518,
    new_n24519, new_n24520, new_n24521, new_n24522, new_n24523, new_n24524,
    new_n24526, new_n24531, new_n24532, new_n24534, new_n24535, new_n24540,
    new_n24541, new_n24542, new_n24543, new_n24544, new_n24545, new_n24546,
    new_n24547, new_n24548, new_n24549, new_n24550, new_n24551, new_n24552,
    new_n24553, new_n24554, new_n24555, new_n24556, new_n24557, new_n24558,
    new_n24559, new_n24560, new_n24561, new_n24562, new_n24563, new_n24564,
    new_n24565, new_n24566, new_n24567, new_n24568, new_n24569, new_n24570,
    new_n24571, new_n24572, new_n24577, new_n24581, new_n24582, new_n24583,
    new_n24584, new_n24585, new_n24595, new_n24596, new_n24605, new_n24611,
    new_n24613, new_n24618, new_n24619, new_n24620, new_n24621, new_n24622,
    new_n24624, new_n24625, new_n24626, new_n24627, new_n24628, new_n24629,
    new_n24630, new_n24652, new_n24653, new_n24656, new_n24658, new_n24659,
    new_n24661, new_n24662, new_n24663, new_n24664, new_n24665, new_n24667,
    new_n24676, new_n24677, new_n24678, new_n24679, new_n24680, new_n24681,
    new_n24682, new_n24683, new_n24684, new_n24685, new_n24686, new_n24687,
    new_n24688, new_n24689, new_n24690, new_n24691, new_n24695, new_n24701,
    new_n24716, new_n24720, new_n24727, new_n24730, new_n24734, new_n24739,
    new_n24740, new_n24746, new_n24747, new_n24748, new_n24751, new_n24752,
    new_n24756, new_n24757, new_n24758, new_n24759, new_n24760, new_n24762,
    new_n24776, new_n24784, new_n24789, new_n24795, new_n24797, new_n24801,
    new_n24805, new_n24812, new_n24817, new_n24823, new_n24828, new_n24834,
    new_n24840, new_n24841, new_n24842, new_n24843, new_n24844, new_n24849,
    new_n24853, new_n24858, new_n24863, new_n24864, new_n24865, new_n24869,
    new_n24870, new_n24874, new_n24875, new_n24884, new_n24903, new_n24904,
    new_n24907, new_n24908, new_n24909, new_n24910, new_n24911, new_n24926,
    new_n24928, new_n24929, new_n24932, new_n24939, new_n24940, new_n24945,
    new_n24947, new_n24948, new_n24949, new_n24950, new_n24951, new_n24952,
    new_n24954, new_n24957, new_n24958, new_n24960, new_n24969, new_n24971,
    new_n24972, new_n24973, new_n24974, new_n24979, new_n24980, new_n24981,
    new_n24982, new_n24988, new_n24989, new_n24999, new_n25000, new_n25001,
    new_n25002, new_n25003, new_n25015, new_n25016, new_n25017, new_n25018,
    new_n25019, new_n25020, new_n25021, new_n25022, new_n25023, new_n25025,
    new_n25032, new_n25035, new_n25036, new_n25039, new_n25040;
  xor_4  g00000(.A(pi683), .B(pi439), .Y(new_n2349));
  nand_5 g00001(.A(pi822), .B(pi567), .Y(new_n2350));
  xor_4  g00002(.A(pi822), .B(pi567), .Y(new_n2351));
  nand_5 g00003(.A(pi100), .B(pi088), .Y(new_n2352));
  nand_5 g00004(.A(pi605), .B(pi117), .Y(new_n2353));
  not_8  g00005(.A(new_n2353), .Y(new_n2354));
  xor_4  g00006(.A(pi605), .B(pi117), .Y(new_n2355));
  not_8  g00007(.A(new_n2355), .Y(new_n2356));
  not_8  g00008(.A(pi434), .Y(new_n2357));
  not_8  g00009(.A(pi514), .Y(new_n2358));
  nor_5  g00010(.A(new_n2358), .B(new_n2357), .Y(new_n2359));
  not_8  g00011(.A(pi369), .Y(new_n2360));
  not_8  g00012(.A(pi552), .Y(new_n2361));
  nor_5  g00013(.A(new_n2361), .B(new_n2360), .Y(new_n2362));
  xor_4  g00014(.A(pi552), .B(pi369), .Y(new_n2363));
  not_8  g00015(.A(new_n2363), .Y(new_n2364));
  nand_5 g00016(.A(pi438), .B(pi190), .Y(new_n2365));
  nor_5  g00017(.A(new_n2365), .B(new_n2364), .Y(new_n2366));
  nor_5  g00018(.A(new_n2366), .B(new_n2362), .Y(new_n2367));
  xor_4  g00019(.A(pi514), .B(new_n2357), .Y(new_n2368));
  nor_5  g00020(.A(new_n2368), .B(new_n2367), .Y(new_n2369));
  nor_5  g00021(.A(new_n2369), .B(new_n2359), .Y(new_n2370));
  nor_5  g00022(.A(new_n2370), .B(new_n2356), .Y(new_n2371));
  nor_5  g00023(.A(new_n2371), .B(new_n2354), .Y(new_n2372));
  not_8  g00024(.A(pi088), .Y(new_n2373));
  xor_4  g00025(.A(pi100), .B(new_n2373), .Y(new_n2374));
  or_6   g00026(.A(new_n2374), .B(new_n2372), .Y(new_n2375));
  nand_5 g00027(.A(new_n2375), .B(new_n2352), .Y(new_n2376));
  nand_5 g00028(.A(new_n2376), .B(new_n2351), .Y(new_n2377));
  nand_5 g00029(.A(new_n2377), .B(new_n2350), .Y(new_n2378));
  xor_4  g00030(.A(new_n2378), .B(new_n2349), .Y(new_n2379));
  not_8  g00031(.A(new_n2379), .Y(new_n2380));
  xor_4  g00032(.A(pi429), .B(pi253), .Y(new_n2381));
  nand_5 g00033(.A(pi829), .B(pi699), .Y(new_n2382));
  xor_4  g00034(.A(pi829), .B(pi699), .Y(new_n2383));
  nand_5 g00035(.A(pi153), .B(pi055), .Y(new_n2384));
  not_8  g00036(.A(pi289), .Y(new_n2385));
  not_8  g00037(.A(pi749), .Y(new_n2386));
  nor_5  g00038(.A(new_n2386), .B(new_n2385), .Y(new_n2387));
  not_8  g00039(.A(pi486), .Y(new_n2388));
  not_8  g00040(.A(pi755), .Y(new_n2389));
  nor_5  g00041(.A(new_n2389), .B(new_n2388), .Y(new_n2390));
  not_8  g00042(.A(pi132), .Y(new_n2391));
  not_8  g00043(.A(pi611), .Y(new_n2392));
  nor_5  g00044(.A(new_n2392), .B(new_n2391), .Y(new_n2393));
  xor_4  g00045(.A(pi611), .B(pi132), .Y(new_n2394));
  not_8  g00046(.A(new_n2394), .Y(new_n2395));
  nand_5 g00047(.A(pi390), .B(pi223), .Y(new_n2396));
  nor_5  g00048(.A(new_n2396), .B(new_n2395), .Y(new_n2397));
  nor_5  g00049(.A(new_n2397), .B(new_n2393), .Y(new_n2398));
  xor_4  g00050(.A(pi755), .B(new_n2388), .Y(new_n2399));
  nor_5  g00051(.A(new_n2399), .B(new_n2398), .Y(new_n2400));
  nor_5  g00052(.A(new_n2400), .B(new_n2390), .Y(new_n2401));
  xor_4  g00053(.A(pi749), .B(new_n2385), .Y(new_n2402));
  nor_5  g00054(.A(new_n2402), .B(new_n2401), .Y(new_n2403));
  nor_5  g00055(.A(new_n2403), .B(new_n2387), .Y(new_n2404));
  not_8  g00056(.A(pi055), .Y(new_n2405));
  xor_4  g00057(.A(pi153), .B(new_n2405), .Y(new_n2406));
  or_6   g00058(.A(new_n2406), .B(new_n2404), .Y(new_n2407));
  nand_5 g00059(.A(new_n2407), .B(new_n2384), .Y(new_n2408));
  nand_5 g00060(.A(new_n2408), .B(new_n2383), .Y(new_n2409));
  nand_5 g00061(.A(new_n2409), .B(new_n2382), .Y(new_n2410));
  xor_4  g00062(.A(new_n2410), .B(new_n2381), .Y(new_n2411));
  not_8  g00063(.A(new_n2411), .Y(new_n2412));
  xor_4  g00064(.A(new_n2408), .B(new_n2383), .Y(new_n2413));
  xor_4  g00065(.A(new_n2368), .B(new_n2367), .Y(new_n2414));
  xor_4  g00066(.A(new_n2399), .B(new_n2398), .Y(new_n2415));
  not_8  g00067(.A(new_n2415), .Y(new_n2416));
  or_6   g00068(.A(new_n2416), .B(new_n2414), .Y(new_n2417));
  xor_4  g00069(.A(new_n2416), .B(new_n2414), .Y(new_n2418));
  not_8  g00070(.A(pi190), .Y(new_n2419));
  not_8  g00071(.A(pi438), .Y(new_n2420));
  nand_5 g00072(.A(new_n2420), .B(new_n2419), .Y(new_n2421));
  nor_5  g00073(.A(new_n2421), .B(new_n2363), .Y(new_n2422));
  nor_5  g00074(.A(new_n2422), .B(new_n2366), .Y(new_n2423));
  not_8  g00075(.A(new_n2396), .Y(new_n2424));
  or_6   g00076(.A(new_n2424), .B(new_n2365), .Y(new_n2425));
  not_8  g00077(.A(new_n2425), .Y(new_n2426));
  not_8  g00078(.A(new_n2421), .Y(new_n2427));
  not_8  g00079(.A(pi223), .Y(new_n2428));
  not_8  g00080(.A(pi390), .Y(new_n2429));
  nand_5 g00081(.A(new_n2429), .B(new_n2428), .Y(new_n2430));
  nor_5  g00082(.A(new_n2430), .B(new_n2427), .Y(new_n2431));
  not_8  g00083(.A(new_n2431), .Y(new_n2432));
  nand_5 g00084(.A(new_n2427), .B(new_n2424), .Y(new_n2433));
  nand_5 g00085(.A(new_n2433), .B(new_n2432), .Y(new_n2434));
  nor_5  g00086(.A(new_n2434), .B(new_n2426), .Y(new_n2435));
  and_6  g00087(.A(new_n2430), .B(new_n2364), .Y(new_n2436));
  nand_5 g00088(.A(new_n2436), .B(new_n2435), .Y(new_n2437));
  and_6  g00089(.A(new_n2433), .B(new_n2395), .Y(new_n2438));
  nand_5 g00090(.A(new_n2438), .B(new_n2437), .Y(new_n2439));
  nor_5  g00091(.A(new_n2432), .B(new_n2364), .Y(new_n2440));
  nor_5  g00092(.A(new_n2440), .B(new_n2397), .Y(new_n2441));
  nand_5 g00093(.A(new_n2441), .B(new_n2439), .Y(new_n2442));
  nand_5 g00094(.A(new_n2442), .B(new_n2423), .Y(new_n2443));
  nand_5 g00095(.A(new_n2443), .B(new_n2418), .Y(new_n2444));
  nand_5 g00096(.A(new_n2444), .B(new_n2417), .Y(new_n2445));
  xor_4  g00097(.A(new_n2370), .B(new_n2355), .Y(new_n2446));
  nor_5  g00098(.A(new_n2446), .B(new_n2445), .Y(new_n2447));
  not_8  g00099(.A(new_n2446), .Y(new_n2448));
  xor_4  g00100(.A(new_n2448), .B(new_n2445), .Y(new_n2449));
  xor_4  g00101(.A(new_n2402), .B(new_n2401), .Y(new_n2450));
  nor_5  g00102(.A(new_n2450), .B(new_n2449), .Y(new_n2451));
  or_6   g00103(.A(new_n2451), .B(new_n2447), .Y(new_n2452));
  xor_4  g00104(.A(new_n2406), .B(new_n2404), .Y(new_n2453));
  not_8  g00105(.A(new_n2453), .Y(new_n2454));
  nor_5  g00106(.A(new_n2454), .B(new_n2452), .Y(new_n2455));
  xor_4  g00107(.A(new_n2374), .B(new_n2372), .Y(new_n2456));
  xor_4  g00108(.A(new_n2453), .B(new_n2452), .Y(new_n2457));
  nor_5  g00109(.A(new_n2457), .B(new_n2456), .Y(new_n2458));
  or_6   g00110(.A(new_n2458), .B(new_n2455), .Y(new_n2459));
  nor_5  g00111(.A(new_n2459), .B(new_n2413), .Y(new_n2460));
  xor_4  g00112(.A(new_n2376), .B(new_n2351), .Y(new_n2461));
  not_8  g00113(.A(new_n2461), .Y(new_n2462));
  xnor_4 g00114(.A(new_n2459), .B(new_n2413), .Y(new_n2463));
  nor_5  g00115(.A(new_n2463), .B(new_n2462), .Y(new_n2464));
  nor_5  g00116(.A(new_n2464), .B(new_n2460), .Y(new_n2465));
  xor_4  g00117(.A(new_n2465), .B(new_n2412), .Y(new_n2466));
  xor_4  g00118(.A(new_n2466), .B(new_n2380), .Y(new_n2467));
  not_8  g00119(.A(pi324), .Y(new_n2468));
  xor_4  g00120(.A(pi348), .B(new_n2468), .Y(new_n2469));
  not_8  g00121(.A(pi659), .Y(new_n2470));
  nand_5 g00122(.A(pi790), .B(new_n2470), .Y(new_n2471));
  not_8  g00123(.A(pi662), .Y(new_n2472));
  nand_5 g00124(.A(new_n2472), .B(pi316), .Y(new_n2473));
  not_8  g00125(.A(pi316), .Y(new_n2474));
  xor_4  g00126(.A(pi662), .B(new_n2474), .Y(new_n2475));
  not_8  g00127(.A(pi831), .Y(new_n2476));
  nand_5 g00128(.A(new_n2476), .B(pi102), .Y(new_n2477));
  not_8  g00129(.A(pi102), .Y(new_n2478));
  xor_4  g00130(.A(pi831), .B(new_n2478), .Y(new_n2479));
  not_8  g00131(.A(pi501), .Y(new_n2480));
  nand_5 g00132(.A(new_n2480), .B(pi204), .Y(new_n2481));
  not_8  g00133(.A(pi204), .Y(new_n2482));
  xor_4  g00134(.A(pi501), .B(new_n2482), .Y(new_n2483));
  not_8  g00135(.A(pi589), .Y(new_n2484));
  nand_5 g00136(.A(pi612), .B(new_n2484), .Y(new_n2485));
  xor_4  g00137(.A(pi612), .B(new_n2484), .Y(new_n2486));
  not_8  g00138(.A(pi077), .Y(new_n2487));
  nand_5 g00139(.A(pi302), .B(new_n2487), .Y(new_n2488));
  not_8  g00140(.A(new_n2488), .Y(new_n2489));
  nand_5 g00141(.A(new_n2489), .B(new_n2486), .Y(new_n2490));
  nand_5 g00142(.A(new_n2490), .B(new_n2485), .Y(new_n2491));
  nand_5 g00143(.A(new_n2491), .B(new_n2483), .Y(new_n2492));
  nand_5 g00144(.A(new_n2492), .B(new_n2481), .Y(new_n2493));
  nand_5 g00145(.A(new_n2493), .B(new_n2479), .Y(new_n2494));
  nand_5 g00146(.A(new_n2494), .B(new_n2477), .Y(new_n2495));
  nand_5 g00147(.A(new_n2495), .B(new_n2475), .Y(new_n2496));
  nand_5 g00148(.A(new_n2496), .B(new_n2473), .Y(new_n2497));
  xor_4  g00149(.A(pi790), .B(new_n2470), .Y(new_n2498));
  nand_5 g00150(.A(new_n2498), .B(new_n2497), .Y(new_n2499));
  nand_5 g00151(.A(new_n2499), .B(new_n2471), .Y(new_n2500));
  xor_4  g00152(.A(new_n2500), .B(new_n2469), .Y(new_n2501));
  xor_4  g00153(.A(new_n2501), .B(new_n2467), .Y(new_n2502));
  xor_4  g00154(.A(new_n2463), .B(new_n2462), .Y(new_n2503));
  xor_4  g00155(.A(new_n2498), .B(new_n2497), .Y(new_n2504));
  or_6   g00156(.A(new_n2504), .B(new_n2503), .Y(new_n2505));
  not_8  g00157(.A(new_n2456), .Y(new_n2506));
  xor_4  g00158(.A(new_n2457), .B(new_n2506), .Y(new_n2507));
  xor_4  g00159(.A(new_n2495), .B(new_n2475), .Y(new_n2508));
  nor_5  g00160(.A(new_n2508), .B(new_n2507), .Y(new_n2509));
  xnor_4 g00161(.A(new_n2450), .B(new_n2449), .Y(new_n2510));
  xor_4  g00162(.A(new_n2493), .B(new_n2479), .Y(new_n2511));
  not_8  g00163(.A(new_n2511), .Y(new_n2512));
  nor_5  g00164(.A(new_n2512), .B(new_n2510), .Y(new_n2513));
  xor_4  g00165(.A(new_n2511), .B(new_n2510), .Y(new_n2514));
  xor_4  g00166(.A(new_n2443), .B(new_n2418), .Y(new_n2515));
  not_8  g00167(.A(new_n2515), .Y(new_n2516));
  xor_4  g00168(.A(new_n2491), .B(new_n2483), .Y(new_n2517));
  or_6   g00169(.A(new_n2517), .B(new_n2516), .Y(new_n2518));
  nand_5 g00170(.A(new_n2517), .B(new_n2516), .Y(new_n2519));
  nand_5 g00171(.A(new_n2430), .B(new_n2396), .Y(new_n2520));
  nand_5 g00172(.A(new_n2421), .B(new_n2365), .Y(new_n2521));
  xor_4  g00173(.A(new_n2521), .B(new_n2520), .Y(new_n2522));
  not_8  g00174(.A(new_n2522), .Y(new_n2523));
  or_6   g00175(.A(new_n2523), .B(new_n2490), .Y(new_n2524));
  not_8  g00176(.A(new_n2486), .Y(new_n2525));
  xor_4  g00177(.A(new_n2435), .B(new_n2364), .Y(new_n2526));
  xor_4  g00178(.A(new_n2526), .B(new_n2395), .Y(new_n2527));
  nand_5 g00179(.A(new_n2523), .B(new_n2489), .Y(new_n2528));
  nor_5  g00180(.A(pi302), .B(new_n2487), .Y(new_n2529));
  nand_5 g00181(.A(new_n2529), .B(new_n2522), .Y(new_n2530));
  nand_5 g00182(.A(new_n2530), .B(new_n2528), .Y(new_n2531));
  xor_4  g00183(.A(new_n2531), .B(new_n2527), .Y(new_n2532));
  or_6   g00184(.A(new_n2532), .B(new_n2525), .Y(new_n2533));
  not_8  g00185(.A(new_n2527), .Y(new_n2534));
  nor_5  g00186(.A(new_n2531), .B(new_n2534), .Y(new_n2535));
  nor_5  g00187(.A(new_n2528), .B(new_n2486), .Y(new_n2536));
  nor_5  g00188(.A(new_n2536), .B(new_n2535), .Y(new_n2537));
  nand_5 g00189(.A(new_n2537), .B(new_n2533), .Y(new_n2538));
  nand_5 g00190(.A(new_n2538), .B(new_n2524), .Y(new_n2539));
  nand_5 g00191(.A(new_n2539), .B(new_n2519), .Y(new_n2540));
  nand_5 g00192(.A(new_n2540), .B(new_n2518), .Y(new_n2541));
  nor_5  g00193(.A(new_n2541), .B(new_n2514), .Y(new_n2542));
  or_6   g00194(.A(new_n2542), .B(new_n2513), .Y(new_n2543));
  not_8  g00195(.A(new_n2507), .Y(new_n2544));
  xor_4  g00196(.A(new_n2508), .B(new_n2544), .Y(new_n2545));
  nor_5  g00197(.A(new_n2545), .B(new_n2543), .Y(new_n2546));
  or_6   g00198(.A(new_n2546), .B(new_n2509), .Y(new_n2547));
  xor_4  g00199(.A(new_n2504), .B(new_n2503), .Y(new_n2548));
  nand_5 g00200(.A(new_n2548), .B(new_n2547), .Y(new_n2549));
  nand_5 g00201(.A(new_n2549), .B(new_n2505), .Y(new_n2550));
  xor_4  g00202(.A(new_n2550), .B(new_n2502), .Y(po0000));
  not_8  g00203(.A(pi149), .Y(new_n2552));
  xor_4  g00204(.A(pi122), .B(pi049), .Y(new_n2553));
  xor_4  g00205(.A(new_n2553), .B(new_n2552), .Y(new_n2554));
  not_8  g00206(.A(pi010), .Y(new_n2555));
  nand_5 g00207(.A(pi702), .B(new_n2555), .Y(new_n2556));
  not_8  g00208(.A(new_n2556), .Y(new_n2557));
  not_8  g00209(.A(pi702), .Y(new_n2558));
  nand_5 g00210(.A(new_n2558), .B(pi010), .Y(new_n2559));
  not_8  g00211(.A(new_n2559), .Y(new_n2560));
  nor_5  g00212(.A(new_n2560), .B(new_n2557), .Y(new_n2561));
  xor_4  g00213(.A(new_n2561), .B(pi677), .Y(new_n2562));
  xor_4  g00214(.A(new_n2562), .B(new_n2554), .Y(po0001));
  not_8  g00215(.A(pi799), .Y(new_n2564));
  not_8  g00216(.A(pi445), .Y(new_n2565));
  xor_4  g00217(.A(pi648), .B(new_n2565), .Y(new_n2566));
  xor_4  g00218(.A(new_n2566), .B(new_n2564), .Y(new_n2567));
  not_8  g00219(.A(pi219), .Y(new_n2568));
  nand_5 g00220(.A(pi606), .B(new_n2568), .Y(new_n2569));
  not_8  g00221(.A(pi606), .Y(new_n2570));
  nand_5 g00222(.A(new_n2570), .B(pi219), .Y(new_n2571));
  nand_5 g00223(.A(new_n2571), .B(new_n2569), .Y(new_n2572));
  xor_4  g00224(.A(new_n2572), .B(pi656), .Y(new_n2573));
  xor_4  g00225(.A(new_n2573), .B(new_n2567), .Y(po0002));
  nand_5 g00226(.A(pi592), .B(pi059), .Y(new_n2575));
  xor_4  g00227(.A(pi592), .B(pi059), .Y(new_n2576));
  nand_5 g00228(.A(pi771), .B(pi551), .Y(new_n2577));
  xor_4  g00229(.A(pi771), .B(pi551), .Y(new_n2578));
  nand_5 g00230(.A(pi420), .B(pi304), .Y(new_n2579));
  xor_4  g00231(.A(pi420), .B(pi304), .Y(new_n2580));
  nand_5 g00232(.A(pi588), .B(pi115), .Y(new_n2581));
  xor_4  g00233(.A(pi588), .B(pi115), .Y(new_n2582));
  nand_5 g00234(.A(pi359), .B(pi173), .Y(new_n2583));
  xor_4  g00235(.A(pi359), .B(pi173), .Y(new_n2584));
  nand_5 g00236(.A(pi535), .B(pi167), .Y(new_n2585));
  xor_4  g00237(.A(pi535), .B(pi167), .Y(new_n2586));
  nor_5  g00238(.A(pi820), .B(pi719), .Y(new_n2587));
  nand_5 g00239(.A(pi376), .B(pi024), .Y(new_n2588));
  not_8  g00240(.A(new_n2588), .Y(new_n2589));
  not_8  g00241(.A(pi719), .Y(new_n2590));
  xor_4  g00242(.A(pi820), .B(new_n2590), .Y(new_n2591));
  nor_5  g00243(.A(new_n2591), .B(new_n2589), .Y(new_n2592));
  nor_5  g00244(.A(new_n2592), .B(new_n2587), .Y(new_n2593));
  nand_5 g00245(.A(new_n2593), .B(new_n2586), .Y(new_n2594));
  nand_5 g00246(.A(new_n2594), .B(new_n2585), .Y(new_n2595));
  nand_5 g00247(.A(new_n2595), .B(new_n2584), .Y(new_n2596));
  nand_5 g00248(.A(new_n2596), .B(new_n2583), .Y(new_n2597));
  nand_5 g00249(.A(new_n2597), .B(new_n2582), .Y(new_n2598));
  nand_5 g00250(.A(new_n2598), .B(new_n2581), .Y(new_n2599));
  nand_5 g00251(.A(new_n2599), .B(new_n2580), .Y(new_n2600));
  nand_5 g00252(.A(new_n2600), .B(new_n2579), .Y(new_n2601));
  nand_5 g00253(.A(new_n2601), .B(new_n2578), .Y(new_n2602));
  nand_5 g00254(.A(new_n2602), .B(new_n2577), .Y(new_n2603));
  nand_5 g00255(.A(new_n2603), .B(new_n2576), .Y(new_n2604));
  nand_5 g00256(.A(new_n2604), .B(new_n2575), .Y(new_n2605));
  nand_5 g00257(.A(pi610), .B(pi308), .Y(new_n2606));
  not_8  g00258(.A(pi308), .Y(new_n2607));
  not_8  g00259(.A(pi610), .Y(new_n2608));
  nand_5 g00260(.A(new_n2608), .B(new_n2607), .Y(new_n2609));
  nand_5 g00261(.A(new_n2609), .B(new_n2606), .Y(new_n2610));
  not_8  g00262(.A(new_n2610), .Y(new_n2611));
  xor_4  g00263(.A(new_n2611), .B(new_n2605), .Y(new_n2612));
  not_8  g00264(.A(pi778), .Y(new_n2613));
  not_8  g00265(.A(pi463), .Y(new_n2614));
  xor_4  g00266(.A(new_n2603), .B(new_n2576), .Y(new_n2615));
  not_8  g00267(.A(new_n2615), .Y(new_n2616));
  nand_5 g00268(.A(new_n2616), .B(new_n2614), .Y(new_n2617));
  xor_4  g00269(.A(new_n2615), .B(pi463), .Y(new_n2618));
  not_8  g00270(.A(new_n2618), .Y(new_n2619));
  xor_4  g00271(.A(new_n2601), .B(new_n2578), .Y(new_n2620));
  nand_5 g00272(.A(new_n2620), .B(pi581), .Y(new_n2621));
  or_6   g00273(.A(new_n2620), .B(pi581), .Y(new_n2622));
  xor_4  g00274(.A(new_n2599), .B(new_n2580), .Y(new_n2623));
  nand_5 g00275(.A(new_n2623), .B(pi286), .Y(new_n2624));
  or_6   g00276(.A(new_n2623), .B(pi286), .Y(new_n2625));
  xor_4  g00277(.A(new_n2597), .B(new_n2582), .Y(new_n2626));
  nand_5 g00278(.A(new_n2626), .B(pi759), .Y(new_n2627));
  or_6   g00279(.A(new_n2626), .B(pi759), .Y(new_n2628));
  xor_4  g00280(.A(new_n2595), .B(new_n2584), .Y(new_n2629));
  nand_5 g00281(.A(new_n2629), .B(pi815), .Y(new_n2630));
  or_6   g00282(.A(new_n2629), .B(pi815), .Y(new_n2631));
  xor_4  g00283(.A(new_n2593), .B(new_n2586), .Y(new_n2632));
  nand_5 g00284(.A(new_n2632), .B(pi496), .Y(new_n2633));
  xor_4  g00285(.A(new_n2591), .B(new_n2588), .Y(new_n2634));
  or_6   g00286(.A(new_n2634), .B(pi283), .Y(new_n2635));
  xor_4  g00287(.A(new_n2634), .B(pi283), .Y(new_n2636));
  not_8  g00288(.A(pi502), .Y(new_n2637));
  not_8  g00289(.A(pi024), .Y(new_n2638));
  xor_4  g00290(.A(pi376), .B(new_n2638), .Y(new_n2639));
  nor_5  g00291(.A(new_n2639), .B(new_n2637), .Y(new_n2640));
  xor_4  g00292(.A(new_n2639), .B(new_n2637), .Y(new_n2641));
  not_8  g00293(.A(new_n2641), .Y(new_n2642));
  nand_5 g00294(.A(pi648), .B(pi580), .Y(new_n2643));
  or_6   g00295(.A(pi648), .B(pi580), .Y(new_n2644));
  nand_5 g00296(.A(new_n2644), .B(pi725), .Y(new_n2645));
  and_6  g00297(.A(new_n2645), .B(new_n2643), .Y(new_n2646));
  nor_5  g00298(.A(new_n2646), .B(new_n2642), .Y(new_n2647));
  nor_5  g00299(.A(new_n2647), .B(new_n2640), .Y(new_n2648));
  nand_5 g00300(.A(new_n2648), .B(new_n2636), .Y(new_n2649));
  nand_5 g00301(.A(new_n2649), .B(new_n2635), .Y(new_n2650));
  not_8  g00302(.A(pi496), .Y(new_n2651));
  xor_4  g00303(.A(new_n2632), .B(new_n2651), .Y(new_n2652));
  or_6   g00304(.A(new_n2652), .B(new_n2650), .Y(new_n2653));
  nand_5 g00305(.A(new_n2653), .B(new_n2633), .Y(new_n2654));
  nand_5 g00306(.A(new_n2654), .B(new_n2631), .Y(new_n2655));
  nand_5 g00307(.A(new_n2655), .B(new_n2630), .Y(new_n2656));
  nand_5 g00308(.A(new_n2656), .B(new_n2628), .Y(new_n2657));
  nand_5 g00309(.A(new_n2657), .B(new_n2627), .Y(new_n2658));
  nand_5 g00310(.A(new_n2658), .B(new_n2625), .Y(new_n2659));
  nand_5 g00311(.A(new_n2659), .B(new_n2624), .Y(new_n2660));
  nand_5 g00312(.A(new_n2660), .B(new_n2622), .Y(new_n2661));
  nand_5 g00313(.A(new_n2661), .B(new_n2621), .Y(new_n2662));
  or_6   g00314(.A(new_n2662), .B(new_n2619), .Y(new_n2663));
  nand_5 g00315(.A(new_n2663), .B(new_n2617), .Y(new_n2664));
  nand_5 g00316(.A(new_n2664), .B(new_n2613), .Y(new_n2665));
  nor_5  g00317(.A(new_n2664), .B(new_n2613), .Y(new_n2666));
  not_8  g00318(.A(new_n2666), .Y(new_n2667));
  nand_5 g00319(.A(new_n2667), .B(new_n2665), .Y(new_n2668));
  xor_4  g00320(.A(new_n2668), .B(new_n2612), .Y(new_n2669));
  xor_4  g00321(.A(new_n2662), .B(new_n2619), .Y(new_n2670));
  not_8  g00322(.A(pi306), .Y(new_n2671));
  xor_4  g00323(.A(pi691), .B(new_n2671), .Y(new_n2672));
  nand_5 g00324(.A(pi407), .B(pi213), .Y(new_n2673));
  not_8  g00325(.A(pi213), .Y(new_n2674));
  not_8  g00326(.A(pi407), .Y(new_n2675));
  nand_5 g00327(.A(new_n2675), .B(new_n2674), .Y(new_n2676));
  nand_5 g00328(.A(pi476), .B(pi116), .Y(new_n2677));
  or_6   g00329(.A(pi476), .B(pi116), .Y(new_n2678));
  nand_5 g00330(.A(pi558), .B(pi211), .Y(new_n2679));
  or_6   g00331(.A(pi558), .B(pi211), .Y(new_n2680));
  nand_5 g00332(.A(pi703), .B(pi231), .Y(new_n2681));
  xor_4  g00333(.A(pi703), .B(pi231), .Y(new_n2682));
  nor_5  g00334(.A(pi449), .B(pi447), .Y(new_n2683));
  xor_4  g00335(.A(pi449), .B(pi447), .Y(new_n2684));
  nand_5 g00336(.A(pi763), .B(pi025), .Y(new_n2685));
  and_6  g00337(.A(new_n2685), .B(new_n2684), .Y(new_n2686));
  nor_5  g00338(.A(new_n2686), .B(new_n2683), .Y(new_n2687));
  nand_5 g00339(.A(new_n2687), .B(new_n2682), .Y(new_n2688));
  nand_5 g00340(.A(new_n2688), .B(new_n2681), .Y(new_n2689));
  nand_5 g00341(.A(new_n2689), .B(new_n2680), .Y(new_n2690));
  nand_5 g00342(.A(new_n2690), .B(new_n2679), .Y(new_n2691));
  nand_5 g00343(.A(new_n2691), .B(new_n2678), .Y(new_n2692));
  nand_5 g00344(.A(new_n2692), .B(new_n2677), .Y(new_n2693));
  nand_5 g00345(.A(new_n2693), .B(new_n2676), .Y(new_n2694));
  nand_5 g00346(.A(new_n2694), .B(new_n2673), .Y(new_n2695));
  xor_4  g00347(.A(new_n2695), .B(new_n2672), .Y(new_n2696));
  not_8  g00348(.A(new_n2696), .Y(new_n2697));
  nand_5 g00349(.A(new_n2673), .B(new_n2676), .Y(new_n2698));
  xor_4  g00350(.A(new_n2698), .B(new_n2693), .Y(new_n2699));
  nand_5 g00351(.A(new_n2678), .B(new_n2677), .Y(new_n2700));
  xor_4  g00352(.A(new_n2700), .B(new_n2691), .Y(new_n2701));
  not_8  g00353(.A(new_n2701), .Y(new_n2702));
  or_6   g00354(.A(new_n2702), .B(pi720), .Y(new_n2703));
  nand_5 g00355(.A(new_n2702), .B(pi720), .Y(new_n2704));
  not_8  g00356(.A(pi521), .Y(new_n2705));
  xor_4  g00357(.A(new_n2685), .B(new_n2684), .Y(new_n2706));
  not_8  g00358(.A(new_n2706), .Y(new_n2707));
  nand_5 g00359(.A(new_n2707), .B(pi370), .Y(new_n2708));
  nand_5 g00360(.A(new_n2708), .B(new_n2705), .Y(new_n2709));
  xor_4  g00361(.A(new_n2708), .B(new_n2705), .Y(new_n2710));
  xor_4  g00362(.A(new_n2687), .B(new_n2682), .Y(new_n2711));
  not_8  g00363(.A(new_n2711), .Y(new_n2712));
  nand_5 g00364(.A(new_n2712), .B(new_n2710), .Y(new_n2713));
  nand_5 g00365(.A(new_n2713), .B(new_n2709), .Y(new_n2714));
  nand_5 g00366(.A(new_n2680), .B(new_n2679), .Y(new_n2715));
  xor_4  g00367(.A(new_n2715), .B(new_n2689), .Y(new_n2716));
  nand_5 g00368(.A(new_n2716), .B(new_n2714), .Y(new_n2717));
  not_8  g00369(.A(pi339), .Y(new_n2718));
  or_6   g00370(.A(new_n2716), .B(new_n2714), .Y(new_n2719));
  nand_5 g00371(.A(new_n2719), .B(new_n2718), .Y(new_n2720));
  nand_5 g00372(.A(new_n2720), .B(new_n2717), .Y(new_n2721));
  nand_5 g00373(.A(new_n2721), .B(new_n2704), .Y(new_n2722));
  nand_5 g00374(.A(new_n2722), .B(new_n2703), .Y(new_n2723));
  or_6   g00375(.A(new_n2723), .B(new_n2699), .Y(new_n2724));
  nand_5 g00376(.A(new_n2723), .B(new_n2699), .Y(new_n2725));
  nand_5 g00377(.A(new_n2725), .B(pi187), .Y(new_n2726));
  nand_5 g00378(.A(new_n2726), .B(new_n2724), .Y(new_n2727));
  nand_5 g00379(.A(new_n2727), .B(new_n2697), .Y(new_n2728));
  or_6   g00380(.A(new_n2727), .B(new_n2697), .Y(new_n2729));
  nand_5 g00381(.A(new_n2729), .B(pi786), .Y(new_n2730));
  nand_5 g00382(.A(new_n2730), .B(new_n2728), .Y(new_n2731));
  xor_4  g00383(.A(new_n2731), .B(pi279), .Y(new_n2732));
  xor_4  g00384(.A(pi233), .B(pi082), .Y(new_n2733));
  nor_5  g00385(.A(pi691), .B(pi306), .Y(new_n2734));
  nor_5  g00386(.A(new_n2695), .B(new_n2672), .Y(new_n2735));
  nor_5  g00387(.A(new_n2735), .B(new_n2734), .Y(new_n2736));
  xor_4  g00388(.A(new_n2736), .B(new_n2733), .Y(new_n2737));
  not_8  g00389(.A(new_n2737), .Y(new_n2738));
  xor_4  g00390(.A(new_n2738), .B(new_n2732), .Y(new_n2739));
  nand_5 g00391(.A(new_n2622), .B(new_n2621), .Y(new_n2740));
  xor_4  g00392(.A(new_n2740), .B(new_n2660), .Y(new_n2741));
  not_8  g00393(.A(new_n2741), .Y(new_n2742));
  or_6   g00394(.A(new_n2742), .B(new_n2739), .Y(new_n2743));
  xor_4  g00395(.A(new_n2646), .B(new_n2641), .Y(new_n2744));
  not_8  g00396(.A(new_n2744), .Y(new_n2745));
  not_8  g00397(.A(pi544), .Y(new_n2746));
  not_8  g00398(.A(pi025), .Y(new_n2747));
  xor_4  g00399(.A(pi763), .B(new_n2747), .Y(new_n2748));
  nand_5 g00400(.A(new_n2748), .B(new_n2746), .Y(new_n2749));
  not_8  g00401(.A(new_n2748), .Y(new_n2750));
  nand_5 g00402(.A(new_n2750), .B(pi544), .Y(new_n2751));
  not_8  g00403(.A(pi580), .Y(new_n2752));
  xor_4  g00404(.A(pi725), .B(new_n2752), .Y(new_n2753));
  xor_4  g00405(.A(new_n2753), .B(pi648), .Y(new_n2754));
  not_8  g00406(.A(new_n2754), .Y(new_n2755));
  nand_5 g00407(.A(new_n2755), .B(new_n2751), .Y(new_n2756));
  nand_5 g00408(.A(new_n2756), .B(new_n2749), .Y(new_n2757));
  nor_5  g00409(.A(new_n2757), .B(new_n2745), .Y(new_n2758));
  xor_4  g00410(.A(new_n2706), .B(pi370), .Y(new_n2759));
  xor_4  g00411(.A(new_n2757), .B(new_n2744), .Y(new_n2760));
  nor_5  g00412(.A(new_n2760), .B(new_n2759), .Y(new_n2761));
  or_6   g00413(.A(new_n2761), .B(new_n2758), .Y(new_n2762));
  xor_4  g00414(.A(new_n2648), .B(new_n2636), .Y(new_n2763));
  nand_5 g00415(.A(new_n2763), .B(new_n2762), .Y(new_n2764));
  not_8  g00416(.A(new_n2763), .Y(new_n2765));
  xor_4  g00417(.A(new_n2765), .B(new_n2762), .Y(new_n2766));
  xor_4  g00418(.A(new_n2712), .B(new_n2710), .Y(new_n2767));
  or_6   g00419(.A(new_n2767), .B(new_n2766), .Y(new_n2768));
  nand_5 g00420(.A(new_n2768), .B(new_n2764), .Y(new_n2769));
  xor_4  g00421(.A(new_n2652), .B(new_n2650), .Y(new_n2770));
  not_8  g00422(.A(new_n2770), .Y(new_n2771));
  nand_5 g00423(.A(new_n2771), .B(new_n2769), .Y(new_n2772));
  nand_5 g00424(.A(new_n2719), .B(new_n2717), .Y(new_n2773));
  xor_4  g00425(.A(new_n2773), .B(pi339), .Y(new_n2774));
  xor_4  g00426(.A(new_n2770), .B(new_n2769), .Y(new_n2775));
  or_6   g00427(.A(new_n2775), .B(new_n2774), .Y(new_n2776));
  nand_5 g00428(.A(new_n2776), .B(new_n2772), .Y(new_n2777));
  nand_5 g00429(.A(new_n2631), .B(new_n2630), .Y(new_n2778));
  xor_4  g00430(.A(new_n2778), .B(new_n2654), .Y(new_n2779));
  or_6   g00431(.A(new_n2779), .B(new_n2777), .Y(new_n2780));
  nand_5 g00432(.A(new_n2704), .B(new_n2703), .Y(new_n2781));
  xor_4  g00433(.A(new_n2781), .B(new_n2721), .Y(new_n2782));
  not_8  g00434(.A(new_n2782), .Y(new_n2783));
  xor_4  g00435(.A(new_n2779), .B(new_n2777), .Y(new_n2784));
  nand_5 g00436(.A(new_n2784), .B(new_n2783), .Y(new_n2785));
  nand_5 g00437(.A(new_n2785), .B(new_n2780), .Y(new_n2786));
  nand_5 g00438(.A(new_n2628), .B(new_n2627), .Y(new_n2787));
  xor_4  g00439(.A(new_n2787), .B(new_n2656), .Y(new_n2788));
  not_8  g00440(.A(new_n2788), .Y(new_n2789));
  nor_5  g00441(.A(new_n2789), .B(new_n2786), .Y(new_n2790));
  nand_5 g00442(.A(new_n2725), .B(new_n2724), .Y(new_n2791));
  xor_4  g00443(.A(new_n2791), .B(pi187), .Y(new_n2792));
  xor_4  g00444(.A(new_n2788), .B(new_n2786), .Y(new_n2793));
  nor_5  g00445(.A(new_n2793), .B(new_n2792), .Y(new_n2794));
  or_6   g00446(.A(new_n2794), .B(new_n2790), .Y(new_n2795));
  nand_5 g00447(.A(new_n2625), .B(new_n2624), .Y(new_n2796));
  xor_4  g00448(.A(new_n2796), .B(new_n2658), .Y(new_n2797));
  nand_5 g00449(.A(new_n2797), .B(new_n2795), .Y(new_n2798));
  nand_5 g00450(.A(new_n2729), .B(new_n2728), .Y(new_n2799));
  xor_4  g00451(.A(new_n2799), .B(pi786), .Y(new_n2800));
  not_8  g00452(.A(new_n2797), .Y(new_n2801));
  xor_4  g00453(.A(new_n2801), .B(new_n2795), .Y(new_n2802));
  or_6   g00454(.A(new_n2802), .B(new_n2800), .Y(new_n2803));
  nand_5 g00455(.A(new_n2803), .B(new_n2798), .Y(new_n2804));
  xor_4  g00456(.A(new_n2742), .B(new_n2739), .Y(new_n2805));
  nand_5 g00457(.A(new_n2805), .B(new_n2804), .Y(new_n2806));
  nand_5 g00458(.A(new_n2806), .B(new_n2743), .Y(new_n2807));
  nand_5 g00459(.A(new_n2807), .B(new_n2670), .Y(new_n2808));
  nand_5 g00460(.A(new_n2731), .B(pi279), .Y(new_n2809));
  nand_5 g00461(.A(new_n2737), .B(new_n2732), .Y(new_n2810));
  nand_5 g00462(.A(new_n2810), .B(new_n2809), .Y(new_n2811));
  xor_4  g00463(.A(pi291), .B(pi016), .Y(new_n2812));
  not_8  g00464(.A(pi082), .Y(new_n2813));
  not_8  g00465(.A(pi233), .Y(new_n2814));
  nand_5 g00466(.A(new_n2814), .B(new_n2813), .Y(new_n2815));
  not_8  g00467(.A(new_n2815), .Y(new_n2816));
  not_8  g00468(.A(new_n2733), .Y(new_n2817));
  nor_5  g00469(.A(new_n2736), .B(new_n2817), .Y(new_n2818));
  nor_5  g00470(.A(new_n2818), .B(new_n2816), .Y(new_n2819));
  xor_4  g00471(.A(new_n2819), .B(new_n2812), .Y(new_n2820));
  nand_5 g00472(.A(new_n2820), .B(new_n2811), .Y(new_n2821));
  nor_5  g00473(.A(new_n2820), .B(new_n2811), .Y(new_n2822));
  not_8  g00474(.A(new_n2822), .Y(new_n2823));
  nand_5 g00475(.A(new_n2823), .B(new_n2821), .Y(new_n2824));
  xor_4  g00476(.A(new_n2824), .B(pi701), .Y(new_n2825));
  not_8  g00477(.A(new_n2670), .Y(new_n2826));
  xor_4  g00478(.A(new_n2807), .B(new_n2826), .Y(new_n2827));
  or_6   g00479(.A(new_n2827), .B(new_n2825), .Y(new_n2828));
  nand_5 g00480(.A(new_n2828), .B(new_n2808), .Y(new_n2829));
  nand_5 g00481(.A(new_n2829), .B(new_n2669), .Y(new_n2830));
  nor_5  g00482(.A(new_n2829), .B(new_n2669), .Y(new_n2831));
  not_8  g00483(.A(new_n2831), .Y(new_n2832));
  nand_5 g00484(.A(new_n2832), .B(new_n2830), .Y(new_n2833));
  nand_5 g00485(.A(new_n2823), .B(pi701), .Y(new_n2834));
  nand_5 g00486(.A(new_n2834), .B(new_n2821), .Y(new_n2835));
  xor_4  g00487(.A(pi679), .B(pi095), .Y(new_n2836));
  not_8  g00488(.A(pi016), .Y(new_n2837));
  not_8  g00489(.A(pi291), .Y(new_n2838));
  nand_5 g00490(.A(new_n2838), .B(new_n2837), .Y(new_n2839));
  not_8  g00491(.A(new_n2839), .Y(new_n2840));
  not_8  g00492(.A(new_n2812), .Y(new_n2841));
  nor_5  g00493(.A(new_n2819), .B(new_n2841), .Y(new_n2842));
  nor_5  g00494(.A(new_n2842), .B(new_n2840), .Y(new_n2843));
  xor_4  g00495(.A(new_n2843), .B(new_n2836), .Y(new_n2844));
  nand_5 g00496(.A(new_n2844), .B(pi443), .Y(new_n2845));
  not_8  g00497(.A(pi443), .Y(new_n2846));
  not_8  g00498(.A(new_n2844), .Y(new_n2847));
  nand_5 g00499(.A(new_n2847), .B(new_n2846), .Y(new_n2848));
  nand_5 g00500(.A(new_n2848), .B(new_n2845), .Y(new_n2849));
  not_8  g00501(.A(new_n2849), .Y(new_n2850));
  xor_4  g00502(.A(new_n2850), .B(new_n2835), .Y(new_n2851));
  xor_4  g00503(.A(new_n2851), .B(new_n2833), .Y(po0003));
  xor_4  g00504(.A(pi687), .B(new_n2837), .Y(new_n2853));
  nand_5 g00505(.A(new_n2814), .B(pi047), .Y(new_n2854));
  not_8  g00506(.A(pi047), .Y(new_n2855));
  xor_4  g00507(.A(pi233), .B(new_n2855), .Y(new_n2856));
  not_8  g00508(.A(pi691), .Y(new_n2857));
  nand_5 g00509(.A(new_n2857), .B(pi410), .Y(new_n2858));
  not_8  g00510(.A(pi410), .Y(new_n2859));
  xor_4  g00511(.A(pi691), .B(new_n2859), .Y(new_n2860));
  nand_5 g00512(.A(new_n2675), .B(pi061), .Y(new_n2861));
  not_8  g00513(.A(pi061), .Y(new_n2862));
  xor_4  g00514(.A(pi407), .B(new_n2862), .Y(new_n2863));
  not_8  g00515(.A(pi116), .Y(new_n2864));
  nand_5 g00516(.A(pi172), .B(new_n2864), .Y(new_n2865));
  xor_4  g00517(.A(pi172), .B(new_n2864), .Y(new_n2866));
  not_8  g00518(.A(pi558), .Y(new_n2867));
  nand_5 g00519(.A(new_n2867), .B(pi151), .Y(new_n2868));
  not_8  g00520(.A(pi231), .Y(new_n2869));
  nand_5 g00521(.A(pi570), .B(new_n2869), .Y(new_n2870));
  not_8  g00522(.A(new_n2870), .Y(new_n2871));
  not_8  g00523(.A(pi144), .Y(new_n2872));
  nand_5 g00524(.A(pi447), .B(new_n2872), .Y(new_n2873));
  not_8  g00525(.A(pi181), .Y(new_n2874));
  not_8  g00526(.A(pi447), .Y(new_n2875));
  nand_5 g00527(.A(new_n2875), .B(pi144), .Y(new_n2876));
  nand_5 g00528(.A(new_n2876), .B(new_n2874), .Y(new_n2877));
  nand_5 g00529(.A(new_n2877), .B(new_n2873), .Y(new_n2878));
  xor_4  g00530(.A(pi570), .B(pi231), .Y(new_n2879));
  nor_5  g00531(.A(new_n2879), .B(new_n2878), .Y(new_n2880));
  nor_5  g00532(.A(new_n2880), .B(new_n2871), .Y(new_n2881));
  not_8  g00533(.A(new_n2881), .Y(new_n2882));
  not_8  g00534(.A(pi151), .Y(new_n2883));
  xor_4  g00535(.A(pi558), .B(new_n2883), .Y(new_n2884));
  nand_5 g00536(.A(new_n2884), .B(new_n2882), .Y(new_n2885));
  nand_5 g00537(.A(new_n2885), .B(new_n2868), .Y(new_n2886));
  nand_5 g00538(.A(new_n2886), .B(new_n2866), .Y(new_n2887));
  nand_5 g00539(.A(new_n2887), .B(new_n2865), .Y(new_n2888));
  nand_5 g00540(.A(new_n2888), .B(new_n2863), .Y(new_n2889));
  nand_5 g00541(.A(new_n2889), .B(new_n2861), .Y(new_n2890));
  nand_5 g00542(.A(new_n2890), .B(new_n2860), .Y(new_n2891));
  nand_5 g00543(.A(new_n2891), .B(new_n2858), .Y(new_n2892));
  nand_5 g00544(.A(new_n2892), .B(new_n2856), .Y(new_n2893));
  nand_5 g00545(.A(new_n2893), .B(new_n2854), .Y(new_n2894));
  xor_4  g00546(.A(new_n2894), .B(new_n2853), .Y(new_n2895));
  xor_4  g00547(.A(pi349), .B(pi224), .Y(new_n2896));
  not_8  g00548(.A(pi239), .Y(new_n2897));
  not_8  g00549(.A(pi600), .Y(new_n2898));
  nand_5 g00550(.A(new_n2898), .B(new_n2897), .Y(new_n2899));
  not_8  g00551(.A(new_n2899), .Y(new_n2900));
  xor_4  g00552(.A(pi600), .B(pi239), .Y(new_n2901));
  not_8  g00553(.A(new_n2901), .Y(new_n2902));
  nor_5  g00554(.A(pi724), .B(pi632), .Y(new_n2903));
  nor_5  g00555(.A(pi756), .B(pi229), .Y(new_n2904));
  xor_4  g00556(.A(pi756), .B(pi229), .Y(new_n2905));
  not_8  g00557(.A(new_n2905), .Y(new_n2906));
  nand_5 g00558(.A(pi406), .B(pi171), .Y(new_n2907));
  not_8  g00559(.A(pi171), .Y(new_n2908));
  not_8  g00560(.A(pi406), .Y(new_n2909));
  nand_5 g00561(.A(new_n2909), .B(new_n2908), .Y(new_n2910));
  nand_5 g00562(.A(pi414), .B(pi023), .Y(new_n2911));
  not_8  g00563(.A(pi023), .Y(new_n2912));
  not_8  g00564(.A(pi414), .Y(new_n2913));
  nand_5 g00565(.A(new_n2913), .B(new_n2912), .Y(new_n2914));
  nand_5 g00566(.A(pi801), .B(pi550), .Y(new_n2915));
  xor_4  g00567(.A(pi801), .B(pi550), .Y(new_n2916));
  nor_5  g00568(.A(pi209), .B(pi044), .Y(new_n2917));
  nand_5 g00569(.A(pi491), .B(pi038), .Y(new_n2918));
  not_8  g00570(.A(new_n2918), .Y(new_n2919));
  not_8  g00571(.A(pi044), .Y(new_n2920));
  xor_4  g00572(.A(pi209), .B(new_n2920), .Y(new_n2921));
  nor_5  g00573(.A(new_n2921), .B(new_n2919), .Y(new_n2922));
  nor_5  g00574(.A(new_n2922), .B(new_n2917), .Y(new_n2923));
  nand_5 g00575(.A(new_n2923), .B(new_n2916), .Y(new_n2924));
  nand_5 g00576(.A(new_n2924), .B(new_n2915), .Y(new_n2925));
  nand_5 g00577(.A(new_n2925), .B(new_n2914), .Y(new_n2926));
  nand_5 g00578(.A(new_n2926), .B(new_n2911), .Y(new_n2927));
  nand_5 g00579(.A(new_n2927), .B(new_n2910), .Y(new_n2928));
  nand_5 g00580(.A(new_n2928), .B(new_n2907), .Y(new_n2929));
  nor_5  g00581(.A(new_n2929), .B(new_n2906), .Y(new_n2930));
  nor_5  g00582(.A(new_n2930), .B(new_n2904), .Y(new_n2931));
  not_8  g00583(.A(pi632), .Y(new_n2932));
  xor_4  g00584(.A(pi724), .B(new_n2932), .Y(new_n2933));
  nor_5  g00585(.A(new_n2933), .B(new_n2931), .Y(new_n2934));
  nor_5  g00586(.A(new_n2934), .B(new_n2903), .Y(new_n2935));
  nor_5  g00587(.A(new_n2935), .B(new_n2902), .Y(new_n2936));
  nor_5  g00588(.A(new_n2936), .B(new_n2900), .Y(new_n2937));
  xor_4  g00589(.A(new_n2937), .B(new_n2896), .Y(new_n2938));
  not_8  g00590(.A(pi380), .Y(new_n2939));
  not_8  g00591(.A(pi527), .Y(new_n2940));
  nand_5 g00592(.A(new_n2940), .B(new_n2939), .Y(new_n2941));
  nand_5 g00593(.A(pi816), .B(pi346), .Y(new_n2942));
  not_8  g00594(.A(pi346), .Y(new_n2943));
  not_8  g00595(.A(pi816), .Y(new_n2944));
  nand_5 g00596(.A(new_n2944), .B(new_n2943), .Y(new_n2945));
  nand_5 g00597(.A(pi709), .B(pi636), .Y(new_n2946));
  nand_5 g00598(.A(pi590), .B(pi263), .Y(new_n2947));
  not_8  g00599(.A(pi328), .Y(new_n2948));
  not_8  g00600(.A(pi766), .Y(new_n2949));
  nand_5 g00601(.A(new_n2949), .B(new_n2948), .Y(new_n2950));
  xor_4  g00602(.A(pi766), .B(pi328), .Y(new_n2951));
  nor_5  g00603(.A(pi504), .B(pi277), .Y(new_n2952));
  nor_5  g00604(.A(pi313), .B(pi309), .Y(new_n2953));
  nand_5 g00605(.A(pi832), .B(pi062), .Y(new_n2954));
  not_8  g00606(.A(new_n2954), .Y(new_n2955));
  not_8  g00607(.A(pi309), .Y(new_n2956));
  xor_4  g00608(.A(pi313), .B(new_n2956), .Y(new_n2957));
  nor_5  g00609(.A(new_n2957), .B(new_n2955), .Y(new_n2958));
  nor_5  g00610(.A(new_n2958), .B(new_n2953), .Y(new_n2959));
  not_8  g00611(.A(pi277), .Y(new_n2960));
  xor_4  g00612(.A(pi504), .B(new_n2960), .Y(new_n2961));
  nor_5  g00613(.A(new_n2961), .B(new_n2959), .Y(new_n2962));
  or_6   g00614(.A(new_n2962), .B(new_n2952), .Y(new_n2963));
  nand_5 g00615(.A(new_n2963), .B(new_n2951), .Y(new_n2964));
  nand_5 g00616(.A(new_n2964), .B(new_n2950), .Y(new_n2965));
  not_8  g00617(.A(pi263), .Y(new_n2966));
  xor_4  g00618(.A(pi590), .B(new_n2966), .Y(new_n2967));
  or_6   g00619(.A(new_n2967), .B(new_n2965), .Y(new_n2968));
  nand_5 g00620(.A(new_n2968), .B(new_n2947), .Y(new_n2969));
  xor_4  g00621(.A(pi709), .B(pi636), .Y(new_n2970));
  nand_5 g00622(.A(new_n2970), .B(new_n2969), .Y(new_n2971));
  nand_5 g00623(.A(new_n2971), .B(new_n2946), .Y(new_n2972));
  nand_5 g00624(.A(new_n2972), .B(new_n2945), .Y(new_n2973));
  nand_5 g00625(.A(new_n2973), .B(new_n2942), .Y(new_n2974));
  nand_5 g00626(.A(new_n2974), .B(new_n2941), .Y(new_n2975));
  nand_5 g00627(.A(pi527), .B(pi380), .Y(new_n2976));
  nand_5 g00628(.A(new_n2976), .B(new_n2975), .Y(new_n2977));
  not_8  g00629(.A(pi404), .Y(new_n2978));
  xor_4  g00630(.A(pi835), .B(new_n2978), .Y(new_n2979));
  xor_4  g00631(.A(new_n2979), .B(new_n2977), .Y(new_n2980));
  xor_4  g00632(.A(new_n2980), .B(new_n2938), .Y(new_n2981));
  xor_4  g00633(.A(new_n2935), .B(new_n2901), .Y(new_n2982));
  nand_5 g00634(.A(new_n2976), .B(new_n2941), .Y(new_n2983));
  xor_4  g00635(.A(new_n2983), .B(new_n2974), .Y(new_n2984));
  nand_5 g00636(.A(new_n2984), .B(new_n2982), .Y(new_n2985));
  xor_4  g00637(.A(new_n2984), .B(new_n2982), .Y(new_n2986));
  xor_4  g00638(.A(new_n2933), .B(new_n2931), .Y(new_n2987));
  not_8  g00639(.A(new_n2987), .Y(new_n2988));
  nand_5 g00640(.A(new_n2945), .B(new_n2942), .Y(new_n2989));
  xor_4  g00641(.A(new_n2989), .B(new_n2972), .Y(new_n2990));
  nand_5 g00642(.A(new_n2990), .B(new_n2988), .Y(new_n2991));
  xor_4  g00643(.A(new_n2990), .B(new_n2988), .Y(new_n2992));
  xor_4  g00644(.A(new_n2929), .B(new_n2905), .Y(new_n2993));
  xor_4  g00645(.A(new_n2970), .B(new_n2969), .Y(new_n2994));
  not_8  g00646(.A(new_n2994), .Y(new_n2995));
  nand_5 g00647(.A(new_n2995), .B(new_n2993), .Y(new_n2996));
  xor_4  g00648(.A(new_n2994), .B(new_n2993), .Y(new_n2997));
  and_6  g00649(.A(new_n2907), .B(new_n2910), .Y(new_n2998));
  xor_4  g00650(.A(new_n2998), .B(new_n2927), .Y(new_n2999));
  xor_4  g00651(.A(new_n2967), .B(new_n2965), .Y(new_n3000));
  not_8  g00652(.A(new_n3000), .Y(new_n3001));
  nand_5 g00653(.A(new_n3001), .B(new_n2999), .Y(new_n3002));
  not_8  g00654(.A(new_n3002), .Y(new_n3003));
  nand_5 g00655(.A(new_n2914), .B(new_n2911), .Y(new_n3004));
  xor_4  g00656(.A(new_n3004), .B(new_n2925), .Y(new_n3005));
  xnor_4 g00657(.A(new_n2963), .B(new_n2951), .Y(new_n3006));
  nand_5 g00658(.A(new_n3006), .B(new_n3005), .Y(new_n3007));
  not_8  g00659(.A(new_n3005), .Y(new_n3008));
  xor_4  g00660(.A(new_n3006), .B(new_n3008), .Y(new_n3009));
  xor_4  g00661(.A(new_n2923), .B(new_n2916), .Y(new_n3010));
  xor_4  g00662(.A(new_n2961), .B(new_n2959), .Y(new_n3011));
  nand_5 g00663(.A(new_n3011), .B(new_n3010), .Y(new_n3012));
  not_8  g00664(.A(new_n3010), .Y(new_n3013));
  not_8  g00665(.A(new_n3011), .Y(new_n3014));
  nand_5 g00666(.A(new_n3014), .B(new_n3013), .Y(new_n3015));
  xor_4  g00667(.A(new_n2921), .B(new_n2919), .Y(new_n3016));
  not_8  g00668(.A(new_n3016), .Y(new_n3017));
  xor_4  g00669(.A(pi491), .B(pi038), .Y(new_n3018));
  not_8  g00670(.A(new_n3018), .Y(new_n3019));
  not_8  g00671(.A(pi062), .Y(new_n3020));
  xor_4  g00672(.A(pi832), .B(new_n3020), .Y(new_n3021));
  not_8  g00673(.A(new_n3021), .Y(new_n3022));
  nand_5 g00674(.A(new_n3022), .B(new_n3019), .Y(new_n3023));
  nand_5 g00675(.A(new_n3023), .B(new_n3017), .Y(new_n3024));
  xor_4  g00676(.A(new_n2957), .B(new_n2955), .Y(new_n3025));
  not_8  g00677(.A(new_n3025), .Y(new_n3026));
  xor_4  g00678(.A(new_n3023), .B(new_n3016), .Y(new_n3027));
  or_6   g00679(.A(new_n3027), .B(new_n3026), .Y(new_n3028));
  nand_5 g00680(.A(new_n3028), .B(new_n3024), .Y(new_n3029));
  nand_5 g00681(.A(new_n3029), .B(new_n3015), .Y(new_n3030));
  nand_5 g00682(.A(new_n3030), .B(new_n3012), .Y(new_n3031));
  or_6   g00683(.A(new_n3031), .B(new_n3009), .Y(new_n3032));
  nand_5 g00684(.A(new_n3032), .B(new_n3007), .Y(new_n3033));
  not_8  g00685(.A(new_n2999), .Y(new_n3034));
  xor_4  g00686(.A(new_n3000), .B(new_n3034), .Y(new_n3035));
  not_8  g00687(.A(new_n3035), .Y(new_n3036));
  nor_5  g00688(.A(new_n3036), .B(new_n3033), .Y(new_n3037));
  nor_5  g00689(.A(new_n3037), .B(new_n3003), .Y(new_n3038));
  or_6   g00690(.A(new_n3038), .B(new_n2997), .Y(new_n3039));
  nand_5 g00691(.A(new_n3039), .B(new_n2996), .Y(new_n3040));
  nand_5 g00692(.A(new_n3040), .B(new_n2992), .Y(new_n3041));
  nand_5 g00693(.A(new_n3041), .B(new_n2991), .Y(new_n3042));
  nand_5 g00694(.A(new_n3042), .B(new_n2986), .Y(new_n3043));
  nand_5 g00695(.A(new_n3043), .B(new_n2985), .Y(new_n3044));
  xor_4  g00696(.A(new_n3044), .B(new_n2981), .Y(new_n3045));
  xor_4  g00697(.A(new_n3045), .B(new_n2895), .Y(new_n3046));
  xor_4  g00698(.A(new_n3042), .B(new_n2986), .Y(new_n3047));
  not_8  g00699(.A(new_n3047), .Y(new_n3048));
  xnor_4 g00700(.A(new_n2892), .B(new_n2856), .Y(new_n3049));
  or_6   g00701(.A(new_n3049), .B(new_n3048), .Y(new_n3050));
  xor_4  g00702(.A(new_n3049), .B(new_n3048), .Y(new_n3051));
  xnor_4 g00703(.A(new_n2890), .B(new_n2860), .Y(new_n3052));
  xor_4  g00704(.A(new_n3040), .B(new_n2992), .Y(new_n3053));
  not_8  g00705(.A(new_n3053), .Y(new_n3054));
  or_6   g00706(.A(new_n3054), .B(new_n3052), .Y(new_n3055));
  xor_4  g00707(.A(new_n3054), .B(new_n3052), .Y(new_n3056));
  xnor_4 g00708(.A(new_n2888), .B(new_n2863), .Y(new_n3057));
  xnor_4 g00709(.A(new_n3038), .B(new_n2997), .Y(new_n3058));
  or_6   g00710(.A(new_n3058), .B(new_n3057), .Y(new_n3059));
  xor_4  g00711(.A(new_n3058), .B(new_n3057), .Y(new_n3060));
  xor_4  g00712(.A(new_n2886), .B(new_n2866), .Y(new_n3061));
  not_8  g00713(.A(new_n3061), .Y(new_n3062));
  xor_4  g00714(.A(new_n3035), .B(new_n3033), .Y(new_n3063));
  nand_5 g00715(.A(new_n3063), .B(new_n3062), .Y(new_n3064));
  xor_4  g00716(.A(new_n3063), .B(new_n3061), .Y(new_n3065));
  xor_4  g00717(.A(new_n3031), .B(new_n3009), .Y(new_n3066));
  xor_4  g00718(.A(new_n2884), .B(new_n2881), .Y(new_n3067));
  nand_5 g00719(.A(new_n3067), .B(new_n3066), .Y(new_n3068));
  xor_4  g00720(.A(new_n2879), .B(new_n2878), .Y(new_n3069));
  nand_5 g00721(.A(new_n3012), .B(new_n3015), .Y(new_n3070));
  xor_4  g00722(.A(new_n3070), .B(new_n3029), .Y(new_n3071));
  not_8  g00723(.A(new_n3071), .Y(new_n3072));
  nor_5  g00724(.A(new_n3072), .B(new_n3069), .Y(new_n3073));
  xor_4  g00725(.A(new_n3071), .B(new_n3069), .Y(new_n3074));
  and_6  g00726(.A(new_n2876), .B(new_n2873), .Y(new_n3075));
  xor_4  g00727(.A(new_n3021), .B(new_n3018), .Y(new_n3076));
  nand_5 g00728(.A(pi181), .B(new_n2747), .Y(new_n3077));
  or_6   g00729(.A(new_n3077), .B(new_n3076), .Y(new_n3078));
  nor_5  g00730(.A(pi181), .B(new_n2747), .Y(new_n3079));
  nand_5 g00731(.A(new_n3079), .B(new_n3076), .Y(new_n3080));
  nand_5 g00732(.A(new_n3080), .B(new_n3078), .Y(new_n3081));
  nand_5 g00733(.A(new_n3081), .B(new_n3075), .Y(new_n3082));
  nand_5 g00734(.A(new_n3075), .B(new_n2874), .Y(new_n3083));
  nand_5 g00735(.A(new_n3083), .B(new_n3078), .Y(new_n3084));
  nand_5 g00736(.A(new_n3084), .B(new_n3082), .Y(new_n3085));
  xor_4  g00737(.A(new_n3027), .B(new_n3026), .Y(new_n3086));
  not_8  g00738(.A(new_n3086), .Y(new_n3087));
  xor_4  g00739(.A(new_n3081), .B(new_n3075), .Y(new_n3088));
  or_6   g00740(.A(new_n3088), .B(new_n3087), .Y(new_n3089));
  nand_5 g00741(.A(new_n3089), .B(new_n3085), .Y(new_n3090));
  nor_5  g00742(.A(new_n3090), .B(new_n3074), .Y(new_n3091));
  or_6   g00743(.A(new_n3091), .B(new_n3073), .Y(new_n3092));
  xor_4  g00744(.A(new_n3067), .B(new_n3066), .Y(new_n3093));
  nand_5 g00745(.A(new_n3093), .B(new_n3092), .Y(new_n3094));
  and_6  g00746(.A(new_n3094), .B(new_n3068), .Y(new_n3095));
  or_6   g00747(.A(new_n3095), .B(new_n3065), .Y(new_n3096));
  nand_5 g00748(.A(new_n3096), .B(new_n3064), .Y(new_n3097));
  not_8  g00749(.A(new_n3097), .Y(new_n3098));
  nand_5 g00750(.A(new_n3098), .B(new_n3060), .Y(new_n3099));
  nand_5 g00751(.A(new_n3099), .B(new_n3059), .Y(new_n3100));
  nand_5 g00752(.A(new_n3100), .B(new_n3056), .Y(new_n3101));
  nand_5 g00753(.A(new_n3101), .B(new_n3055), .Y(new_n3102));
  nand_5 g00754(.A(new_n3102), .B(new_n3051), .Y(new_n3103));
  nand_5 g00755(.A(new_n3103), .B(new_n3050), .Y(new_n3104));
  xor_4  g00756(.A(new_n3104), .B(new_n3046), .Y(po0004));
  nand_5 g00757(.A(pi234), .B(pi142), .Y(new_n3106));
  nand_5 g00758(.A(pi721), .B(pi189), .Y(new_n3107));
  xor_4  g00759(.A(pi721), .B(pi189), .Y(new_n3108));
  nand_5 g00760(.A(pi424), .B(pi417), .Y(new_n3109));
  xor_4  g00761(.A(pi424), .B(pi417), .Y(new_n3110));
  nand_5 g00762(.A(pi348), .B(pi018), .Y(new_n3111));
  xor_4  g00763(.A(pi348), .B(pi018), .Y(new_n3112));
  nand_5 g00764(.A(pi659), .B(pi217), .Y(new_n3113));
  xor_4  g00765(.A(pi659), .B(pi217), .Y(new_n3114));
  nand_5 g00766(.A(pi662), .B(pi107), .Y(new_n3115));
  xor_4  g00767(.A(pi662), .B(pi107), .Y(new_n3116));
  nand_5 g00768(.A(pi831), .B(pi629), .Y(new_n3117));
  xor_4  g00769(.A(pi831), .B(pi629), .Y(new_n3118));
  nand_5 g00770(.A(pi501), .B(pi076), .Y(new_n3119));
  xor_4  g00771(.A(pi501), .B(pi076), .Y(new_n3120));
  nor_5  g00772(.A(pi589), .B(pi354), .Y(new_n3121));
  nand_5 g00773(.A(pi500), .B(pi077), .Y(new_n3122));
  not_8  g00774(.A(new_n3122), .Y(new_n3123));
  not_8  g00775(.A(pi354), .Y(new_n3124));
  xor_4  g00776(.A(pi589), .B(new_n3124), .Y(new_n3125));
  nor_5  g00777(.A(new_n3125), .B(new_n3123), .Y(new_n3126));
  nor_5  g00778(.A(new_n3126), .B(new_n3121), .Y(new_n3127));
  nand_5 g00779(.A(new_n3127), .B(new_n3120), .Y(new_n3128));
  nand_5 g00780(.A(new_n3128), .B(new_n3119), .Y(new_n3129));
  nand_5 g00781(.A(new_n3129), .B(new_n3118), .Y(new_n3130));
  nand_5 g00782(.A(new_n3130), .B(new_n3117), .Y(new_n3131));
  nand_5 g00783(.A(new_n3131), .B(new_n3116), .Y(new_n3132));
  nand_5 g00784(.A(new_n3132), .B(new_n3115), .Y(new_n3133));
  nand_5 g00785(.A(new_n3133), .B(new_n3114), .Y(new_n3134));
  nand_5 g00786(.A(new_n3134), .B(new_n3113), .Y(new_n3135));
  nand_5 g00787(.A(new_n3135), .B(new_n3112), .Y(new_n3136));
  nand_5 g00788(.A(new_n3136), .B(new_n3111), .Y(new_n3137));
  nand_5 g00789(.A(new_n3137), .B(new_n3110), .Y(new_n3138));
  nand_5 g00790(.A(new_n3138), .B(new_n3109), .Y(new_n3139));
  nand_5 g00791(.A(new_n3139), .B(new_n3108), .Y(new_n3140));
  nand_5 g00792(.A(new_n3140), .B(new_n3107), .Y(new_n3141));
  xor_4  g00793(.A(pi234), .B(pi142), .Y(new_n3142));
  nand_5 g00794(.A(new_n3142), .B(new_n3141), .Y(new_n3143));
  nand_5 g00795(.A(new_n3143), .B(new_n3106), .Y(new_n3144));
  not_8  g00796(.A(new_n3144), .Y(new_n3145));
  not_8  g00797(.A(pi160), .Y(new_n3146));
  not_8  g00798(.A(pi208), .Y(new_n3147));
  xor_4  g00799(.A(new_n3139), .B(new_n3108), .Y(new_n3148));
  nand_5 g00800(.A(new_n3148), .B(new_n3147), .Y(new_n3149));
  xor_4  g00801(.A(new_n3148), .B(new_n3147), .Y(new_n3150));
  not_8  g00802(.A(new_n3150), .Y(new_n3151));
  xor_4  g00803(.A(new_n3137), .B(new_n3110), .Y(new_n3152));
  not_8  g00804(.A(new_n3152), .Y(new_n3153));
  nand_5 g00805(.A(new_n3153), .B(pi802), .Y(new_n3154));
  not_8  g00806(.A(pi802), .Y(new_n3155));
  xor_4  g00807(.A(new_n3152), .B(new_n3155), .Y(new_n3156));
  not_8  g00808(.A(pi601), .Y(new_n3157));
  xor_4  g00809(.A(new_n3135), .B(new_n3112), .Y(new_n3158));
  nor_5  g00810(.A(new_n3158), .B(new_n3157), .Y(new_n3159));
  xor_4  g00811(.A(new_n3158), .B(new_n3157), .Y(new_n3160));
  not_8  g00812(.A(new_n3160), .Y(new_n3161));
  xor_4  g00813(.A(new_n3133), .B(new_n3114), .Y(new_n3162));
  xor_4  g00814(.A(new_n3129), .B(new_n3118), .Y(new_n3163));
  not_8  g00815(.A(new_n3163), .Y(new_n3164));
  xor_4  g00816(.A(new_n3127), .B(new_n3120), .Y(new_n3165));
  not_8  g00817(.A(new_n3165), .Y(new_n3166));
  nand_5 g00818(.A(new_n3166), .B(pi652), .Y(new_n3167));
  not_8  g00819(.A(pi776), .Y(new_n3168));
  xor_4  g00820(.A(pi500), .B(pi077), .Y(new_n3169));
  not_8  g00821(.A(new_n3169), .Y(new_n3170));
  nor_5  g00822(.A(new_n3170), .B(pi364), .Y(new_n3171));
  nand_5 g00823(.A(new_n3171), .B(new_n3168), .Y(new_n3172));
  xor_4  g00824(.A(new_n3171), .B(new_n3168), .Y(new_n3173));
  xor_4  g00825(.A(new_n3125), .B(new_n3122), .Y(new_n3174));
  nand_5 g00826(.A(new_n3174), .B(new_n3173), .Y(new_n3175));
  nand_5 g00827(.A(new_n3175), .B(new_n3172), .Y(new_n3176));
  xor_4  g00828(.A(new_n3165), .B(pi652), .Y(new_n3177));
  or_6   g00829(.A(new_n3177), .B(new_n3176), .Y(new_n3178));
  nand_5 g00830(.A(new_n3178), .B(new_n3167), .Y(new_n3179));
  or_6   g00831(.A(new_n3179), .B(new_n3164), .Y(new_n3180));
  nand_5 g00832(.A(new_n3180), .B(pi036), .Y(new_n3181));
  nand_5 g00833(.A(new_n3179), .B(new_n3164), .Y(new_n3182));
  nand_5 g00834(.A(new_n3182), .B(new_n3181), .Y(new_n3183));
  xnor_4 g00835(.A(new_n3131), .B(new_n3116), .Y(new_n3184));
  or_6   g00836(.A(new_n3184), .B(new_n3183), .Y(new_n3185));
  not_8  g00837(.A(pi285), .Y(new_n3186));
  nand_5 g00838(.A(new_n3184), .B(new_n3183), .Y(new_n3187));
  nand_5 g00839(.A(new_n3187), .B(new_n3186), .Y(new_n3188));
  nand_5 g00840(.A(new_n3188), .B(new_n3185), .Y(new_n3189));
  nand_5 g00841(.A(new_n3189), .B(new_n3162), .Y(new_n3190));
  not_8  g00842(.A(pi290), .Y(new_n3191));
  xor_4  g00843(.A(new_n3189), .B(new_n3162), .Y(new_n3192));
  nand_5 g00844(.A(new_n3192), .B(new_n3191), .Y(new_n3193));
  nand_5 g00845(.A(new_n3193), .B(new_n3190), .Y(new_n3194));
  nor_5  g00846(.A(new_n3194), .B(new_n3161), .Y(new_n3195));
  or_6   g00847(.A(new_n3195), .B(new_n3159), .Y(new_n3196));
  nand_5 g00848(.A(new_n3196), .B(new_n3156), .Y(new_n3197));
  nand_5 g00849(.A(new_n3197), .B(new_n3154), .Y(new_n3198));
  or_6   g00850(.A(new_n3198), .B(new_n3151), .Y(new_n3199));
  nand_5 g00851(.A(new_n3199), .B(new_n3149), .Y(new_n3200));
  or_6   g00852(.A(new_n3200), .B(new_n3146), .Y(new_n3201));
  xor_4  g00853(.A(new_n3142), .B(new_n3141), .Y(new_n3202));
  nand_5 g00854(.A(new_n3200), .B(new_n3146), .Y(new_n3203));
  nand_5 g00855(.A(new_n3203), .B(new_n3201), .Y(new_n3204));
  or_6   g00856(.A(new_n3204), .B(new_n3202), .Y(new_n3205));
  nand_5 g00857(.A(new_n3205), .B(new_n3201), .Y(new_n3206));
  nand_5 g00858(.A(new_n3206), .B(new_n3145), .Y(new_n3207));
  not_8  g00859(.A(pi166), .Y(new_n3208));
  not_8  g00860(.A(pi244), .Y(new_n3209));
  nand_5 g00861(.A(new_n3209), .B(new_n3208), .Y(new_n3210));
  nand_5 g00862(.A(pi244), .B(pi166), .Y(new_n3211));
  not_8  g00863(.A(pi005), .Y(new_n3212));
  not_8  g00864(.A(pi509), .Y(new_n3213));
  nand_5 g00865(.A(new_n3213), .B(new_n3212), .Y(new_n3214));
  nand_5 g00866(.A(pi509), .B(pi005), .Y(new_n3215));
  or_6   g00867(.A(pi690), .B(pi105), .Y(new_n3216));
  nand_5 g00868(.A(pi690), .B(pi105), .Y(new_n3217));
  not_8  g00869(.A(pi175), .Y(new_n3218));
  not_8  g00870(.A(pi575), .Y(new_n3219));
  nand_5 g00871(.A(new_n3219), .B(new_n3218), .Y(new_n3220));
  nand_5 g00872(.A(pi575), .B(pi175), .Y(new_n3221));
  not_8  g00873(.A(pi225), .Y(new_n3222));
  not_8  g00874(.A(pi792), .Y(new_n3223));
  nand_5 g00875(.A(new_n3223), .B(new_n3222), .Y(new_n3224));
  xor_4  g00876(.A(pi792), .B(pi225), .Y(new_n3225));
  not_8  g00877(.A(pi584), .Y(new_n3226));
  not_8  g00878(.A(pi649), .Y(new_n3227));
  nand_5 g00879(.A(new_n3227), .B(new_n3226), .Y(new_n3228));
  xor_4  g00880(.A(pi649), .B(pi584), .Y(new_n3229));
  not_8  g00881(.A(pi074), .Y(new_n3230));
  not_8  g00882(.A(pi563), .Y(new_n3231));
  nand_5 g00883(.A(new_n3231), .B(new_n3230), .Y(new_n3232));
  nand_5 g00884(.A(pi563), .B(pi074), .Y(new_n3233));
  not_8  g00885(.A(pi457), .Y(new_n3234));
  not_8  g00886(.A(pi468), .Y(new_n3235));
  nand_5 g00887(.A(new_n3235), .B(new_n3234), .Y(new_n3236));
  nand_5 g00888(.A(pi468), .B(pi457), .Y(new_n3237));
  not_8  g00889(.A(pi633), .Y(new_n3238));
  not_8  g00890(.A(pi783), .Y(new_n3239));
  nand_5 g00891(.A(new_n3239), .B(new_n3238), .Y(new_n3240));
  nand_5 g00892(.A(pi783), .B(pi633), .Y(new_n3241));
  nand_5 g00893(.A(pi718), .B(pi508), .Y(new_n3242));
  nand_5 g00894(.A(new_n3242), .B(new_n3241), .Y(new_n3243));
  nand_5 g00895(.A(new_n3243), .B(new_n3240), .Y(new_n3244));
  nand_5 g00896(.A(new_n3244), .B(new_n3237), .Y(new_n3245));
  nand_5 g00897(.A(new_n3245), .B(new_n3236), .Y(new_n3246));
  nand_5 g00898(.A(new_n3246), .B(new_n3233), .Y(new_n3247));
  nand_5 g00899(.A(new_n3247), .B(new_n3232), .Y(new_n3248));
  nand_5 g00900(.A(new_n3248), .B(new_n3229), .Y(new_n3249));
  nand_5 g00901(.A(new_n3249), .B(new_n3228), .Y(new_n3250));
  nand_5 g00902(.A(new_n3250), .B(new_n3225), .Y(new_n3251));
  nand_5 g00903(.A(new_n3251), .B(new_n3224), .Y(new_n3252));
  nand_5 g00904(.A(new_n3252), .B(new_n3221), .Y(new_n3253));
  nand_5 g00905(.A(new_n3253), .B(new_n3220), .Y(new_n3254));
  nand_5 g00906(.A(new_n3254), .B(new_n3217), .Y(new_n3255));
  nand_5 g00907(.A(new_n3255), .B(new_n3216), .Y(new_n3256));
  nand_5 g00908(.A(new_n3256), .B(new_n3215), .Y(new_n3257));
  nand_5 g00909(.A(new_n3257), .B(new_n3214), .Y(new_n3258));
  nand_5 g00910(.A(new_n3258), .B(new_n3211), .Y(new_n3259));
  nand_5 g00911(.A(new_n3259), .B(new_n3210), .Y(new_n3260));
  xor_4  g00912(.A(new_n3204), .B(new_n3202), .Y(new_n3261));
  not_8  g00913(.A(pi325), .Y(new_n3262));
  xnor_4 g00914(.A(new_n3196), .B(new_n3156), .Y(new_n3263));
  not_8  g00915(.A(pi829), .Y(new_n3264));
  xor_4  g00916(.A(new_n3192), .B(pi290), .Y(new_n3265));
  nor_5  g00917(.A(new_n3265), .B(new_n3264), .Y(new_n3266));
  xor_4  g00918(.A(new_n3265), .B(new_n3264), .Y(new_n3267));
  not_8  g00919(.A(new_n3267), .Y(new_n3268));
  xor_4  g00920(.A(new_n3170), .B(pi364), .Y(new_n3269));
  nand_5 g00921(.A(new_n3269), .B(pi390), .Y(new_n3270));
  nand_5 g00922(.A(new_n3270), .B(new_n2391), .Y(new_n3271));
  xor_4  g00923(.A(new_n3270), .B(pi132), .Y(new_n3272));
  xor_4  g00924(.A(new_n3174), .B(new_n3173), .Y(new_n3273));
  or_6   g00925(.A(new_n3273), .B(new_n3272), .Y(new_n3274));
  nand_5 g00926(.A(new_n3274), .B(new_n3271), .Y(new_n3275));
  xor_4  g00927(.A(new_n3177), .B(new_n3176), .Y(new_n3276));
  nand_5 g00928(.A(new_n3276), .B(new_n3275), .Y(new_n3277));
  or_6   g00929(.A(new_n3276), .B(new_n3275), .Y(new_n3278));
  nand_5 g00930(.A(new_n3278), .B(new_n2389), .Y(new_n3279));
  nand_5 g00931(.A(new_n3279), .B(new_n3277), .Y(new_n3280));
  nor_5  g00932(.A(new_n3280), .B(new_n2386), .Y(new_n3281));
  not_8  g00933(.A(pi036), .Y(new_n3282));
  and_6  g00934(.A(new_n3182), .B(new_n3180), .Y(new_n3283));
  xor_4  g00935(.A(new_n3283), .B(new_n3282), .Y(new_n3284));
  not_8  g00936(.A(new_n3284), .Y(new_n3285));
  xor_4  g00937(.A(new_n3280), .B(pi749), .Y(new_n3286));
  nor_5  g00938(.A(new_n3286), .B(new_n3285), .Y(new_n3287));
  or_6   g00939(.A(new_n3287), .B(new_n3281), .Y(new_n3288));
  nand_5 g00940(.A(new_n3187), .B(new_n3185), .Y(new_n3289));
  xor_4  g00941(.A(new_n3289), .B(pi285), .Y(new_n3290));
  nand_5 g00942(.A(new_n3290), .B(new_n3288), .Y(new_n3291));
  or_6   g00943(.A(new_n3290), .B(new_n3288), .Y(new_n3292));
  nand_5 g00944(.A(new_n3292), .B(pi153), .Y(new_n3293));
  and_6  g00945(.A(new_n3293), .B(new_n3291), .Y(new_n3294));
  nor_5  g00946(.A(new_n3294), .B(new_n3268), .Y(new_n3295));
  or_6   g00947(.A(new_n3295), .B(new_n3266), .Y(new_n3296));
  xor_4  g00948(.A(new_n3194), .B(new_n3160), .Y(new_n3297));
  nand_5 g00949(.A(new_n3297), .B(new_n3296), .Y(new_n3298));
  or_6   g00950(.A(new_n3297), .B(new_n3296), .Y(new_n3299));
  nand_5 g00951(.A(new_n3299), .B(pi253), .Y(new_n3300));
  nand_5 g00952(.A(new_n3300), .B(new_n3298), .Y(new_n3301));
  or_6   g00953(.A(new_n3301), .B(new_n3263), .Y(new_n3302));
  not_8  g00954(.A(pi637), .Y(new_n3303));
  nand_5 g00955(.A(new_n3301), .B(new_n3263), .Y(new_n3304));
  nand_5 g00956(.A(new_n3304), .B(new_n3303), .Y(new_n3305));
  nand_5 g00957(.A(new_n3305), .B(new_n3302), .Y(new_n3306));
  nand_5 g00958(.A(new_n3306), .B(new_n3262), .Y(new_n3307));
  xor_4  g00959(.A(new_n3306), .B(pi325), .Y(new_n3308));
  xor_4  g00960(.A(new_n3198), .B(new_n3150), .Y(new_n3309));
  not_8  g00961(.A(new_n3309), .Y(new_n3310));
  or_6   g00962(.A(new_n3310), .B(new_n3308), .Y(new_n3311));
  nand_5 g00963(.A(new_n3311), .B(new_n3307), .Y(new_n3312));
  nand_5 g00964(.A(new_n3312), .B(new_n3261), .Y(new_n3313));
  not_8  g00965(.A(new_n3313), .Y(new_n3314));
  not_8  g00966(.A(new_n3261), .Y(new_n3315));
  xor_4  g00967(.A(new_n3312), .B(new_n3315), .Y(new_n3316));
  nor_5  g00968(.A(new_n3316), .B(pi114), .Y(new_n3317));
  nor_5  g00969(.A(new_n3317), .B(new_n3314), .Y(new_n3318));
  nor_5  g00970(.A(new_n3203), .B(new_n3145), .Y(new_n3319));
  not_8  g00971(.A(new_n3106), .Y(new_n3320));
  nand_5 g00972(.A(new_n3141), .B(new_n3320), .Y(new_n3321));
  nor_5  g00973(.A(new_n3321), .B(new_n3315), .Y(new_n3322));
  nor_5  g00974(.A(new_n3322), .B(new_n3319), .Y(new_n3323));
  nand_5 g00975(.A(new_n3323), .B(new_n3207), .Y(new_n3324));
  xor_4  g00976(.A(new_n3324), .B(new_n3318), .Y(new_n3325));
  nand_5 g00977(.A(new_n3325), .B(new_n3260), .Y(new_n3326));
  not_8  g00978(.A(pi114), .Y(new_n3327));
  xor_4  g00979(.A(new_n3316), .B(new_n3327), .Y(new_n3328));
  not_8  g00980(.A(new_n3258), .Y(new_n3329));
  nand_5 g00981(.A(new_n3210), .B(new_n3211), .Y(new_n3330));
  xor_4  g00982(.A(new_n3330), .B(new_n3329), .Y(new_n3331));
  nand_5 g00983(.A(new_n3331), .B(new_n3328), .Y(new_n3332));
  not_8  g00984(.A(pi253), .Y(new_n3333));
  nand_5 g00985(.A(new_n3299), .B(new_n3298), .Y(new_n3334));
  xor_4  g00986(.A(new_n3334), .B(new_n3333), .Y(new_n3335));
  xor_4  g00987(.A(new_n3250), .B(new_n3225), .Y(new_n3336));
  xor_4  g00988(.A(new_n3248), .B(new_n3229), .Y(new_n3337));
  not_8  g00989(.A(new_n3337), .Y(new_n3338));
  not_8  g00990(.A(pi508), .Y(new_n3339));
  not_8  g00991(.A(pi718), .Y(new_n3340));
  nand_5 g00992(.A(new_n3340), .B(new_n3339), .Y(new_n3341));
  nand_5 g00993(.A(new_n3341), .B(new_n3242), .Y(new_n3342));
  not_8  g00994(.A(new_n3342), .Y(new_n3343));
  xor_4  g00995(.A(new_n3269), .B(new_n2429), .Y(new_n3344));
  and_6  g00996(.A(new_n3344), .B(new_n3343), .Y(new_n3345));
  nand_5 g00997(.A(new_n3241), .B(new_n3240), .Y(new_n3346));
  xor_4  g00998(.A(new_n3346), .B(new_n3242), .Y(new_n3347));
  or_6   g00999(.A(new_n3347), .B(new_n3345), .Y(new_n3348));
  not_8  g01000(.A(new_n3341), .Y(new_n3349));
  nor_5  g01001(.A(new_n3346), .B(new_n3349), .Y(new_n3350));
  nand_5 g01002(.A(new_n3350), .B(new_n3344), .Y(new_n3351));
  nand_5 g01003(.A(new_n3351), .B(new_n3348), .Y(new_n3352));
  xor_4  g01004(.A(new_n3273), .B(new_n3272), .Y(new_n3353));
  or_6   g01005(.A(new_n3353), .B(new_n3352), .Y(new_n3354));
  nand_5 g01006(.A(new_n3354), .B(new_n3348), .Y(new_n3355));
  nand_5 g01007(.A(new_n3237), .B(new_n3236), .Y(new_n3356));
  xor_4  g01008(.A(new_n3356), .B(new_n3244), .Y(new_n3357));
  not_8  g01009(.A(new_n3357), .Y(new_n3358));
  or_6   g01010(.A(new_n3358), .B(new_n3355), .Y(new_n3359));
  xor_4  g01011(.A(new_n3358), .B(new_n3355), .Y(new_n3360));
  nand_5 g01012(.A(new_n3278), .B(new_n3277), .Y(new_n3361));
  xor_4  g01013(.A(new_n3361), .B(pi755), .Y(new_n3362));
  nand_5 g01014(.A(new_n3362), .B(new_n3360), .Y(new_n3363));
  nand_5 g01015(.A(new_n3363), .B(new_n3359), .Y(new_n3364));
  and_6  g01016(.A(new_n3232), .B(new_n3233), .Y(new_n3365));
  xor_4  g01017(.A(new_n3365), .B(new_n3246), .Y(new_n3366));
  not_8  g01018(.A(new_n3366), .Y(new_n3367));
  nand_5 g01019(.A(new_n3367), .B(new_n3364), .Y(new_n3368));
  xor_4  g01020(.A(new_n3366), .B(new_n3364), .Y(new_n3369));
  xor_4  g01021(.A(new_n3286), .B(new_n3284), .Y(new_n3370));
  not_8  g01022(.A(new_n3370), .Y(new_n3371));
  or_6   g01023(.A(new_n3371), .B(new_n3369), .Y(new_n3372));
  nand_5 g01024(.A(new_n3372), .B(new_n3368), .Y(new_n3373));
  nor_5  g01025(.A(new_n3373), .B(new_n3338), .Y(new_n3374));
  nand_5 g01026(.A(new_n3292), .B(new_n3291), .Y(new_n3375));
  xor_4  g01027(.A(new_n3375), .B(pi153), .Y(new_n3376));
  xor_4  g01028(.A(new_n3373), .B(new_n3337), .Y(new_n3377));
  nor_5  g01029(.A(new_n3377), .B(new_n3376), .Y(new_n3378));
  or_6   g01030(.A(new_n3378), .B(new_n3374), .Y(new_n3379));
  nor_5  g01031(.A(new_n3379), .B(new_n3336), .Y(new_n3380));
  xor_4  g01032(.A(new_n3379), .B(new_n3336), .Y(new_n3381));
  xor_4  g01033(.A(new_n3294), .B(new_n3267), .Y(new_n3382));
  nand_5 g01034(.A(new_n3382), .B(new_n3381), .Y(new_n3383));
  not_8  g01035(.A(new_n3383), .Y(new_n3384));
  nor_5  g01036(.A(new_n3384), .B(new_n3380), .Y(new_n3385));
  nand_5 g01037(.A(new_n3385), .B(new_n3335), .Y(new_n3386));
  xnor_4 g01038(.A(new_n3385), .B(new_n3335), .Y(new_n3387));
  nand_5 g01039(.A(new_n3221), .B(new_n3220), .Y(new_n3388));
  xor_4  g01040(.A(new_n3388), .B(new_n3252), .Y(new_n3389));
  or_6   g01041(.A(new_n3389), .B(new_n3387), .Y(new_n3390));
  nand_5 g01042(.A(new_n3390), .B(new_n3386), .Y(new_n3391));
  nand_5 g01043(.A(new_n3217), .B(new_n3216), .Y(new_n3392));
  xor_4  g01044(.A(new_n3392), .B(new_n3254), .Y(new_n3393));
  not_8  g01045(.A(new_n3393), .Y(new_n3394));
  nand_5 g01046(.A(new_n3394), .B(new_n3391), .Y(new_n3395));
  nand_5 g01047(.A(new_n3304), .B(new_n3302), .Y(new_n3396));
  xor_4  g01048(.A(new_n3396), .B(new_n3303), .Y(new_n3397));
  xor_4  g01049(.A(new_n3393), .B(new_n3391), .Y(new_n3398));
  not_8  g01050(.A(new_n3398), .Y(new_n3399));
  nand_5 g01051(.A(new_n3399), .B(new_n3397), .Y(new_n3400));
  nand_5 g01052(.A(new_n3400), .B(new_n3395), .Y(new_n3401));
  xor_4  g01053(.A(new_n3309), .B(new_n3308), .Y(new_n3402));
  nand_5 g01054(.A(new_n3402), .B(new_n3401), .Y(new_n3403));
  xor_4  g01055(.A(new_n3402), .B(new_n3401), .Y(new_n3404));
  nand_5 g01056(.A(new_n3214), .B(new_n3215), .Y(new_n3405));
  xnor_4 g01057(.A(new_n3405), .B(new_n3256), .Y(new_n3406));
  nand_5 g01058(.A(new_n3406), .B(new_n3404), .Y(new_n3407));
  nand_5 g01059(.A(new_n3407), .B(new_n3403), .Y(new_n3408));
  xor_4  g01060(.A(new_n3331), .B(new_n3328), .Y(new_n3409));
  nand_5 g01061(.A(new_n3409), .B(new_n3408), .Y(new_n3410));
  nand_5 g01062(.A(new_n3410), .B(new_n3332), .Y(new_n3411));
  xor_4  g01063(.A(new_n3325), .B(new_n3260), .Y(new_n3412));
  nand_5 g01064(.A(new_n3412), .B(new_n3411), .Y(new_n3413));
  nand_5 g01065(.A(new_n3413), .B(new_n3326), .Y(new_n3414));
  nor_5  g01066(.A(new_n3414), .B(new_n3207), .Y(new_n3415));
  not_8  g01067(.A(new_n3207), .Y(new_n3416));
  or_6   g01068(.A(new_n3318), .B(new_n3416), .Y(new_n3417));
  nand_5 g01069(.A(new_n3323), .B(new_n3318), .Y(new_n3418));
  nand_5 g01070(.A(new_n3418), .B(new_n3417), .Y(new_n3419));
  nand_5 g01071(.A(new_n3414), .B(new_n3207), .Y(new_n3420));
  nand_5 g01072(.A(new_n3420), .B(new_n3419), .Y(new_n3421));
  nor_5  g01073(.A(new_n3421), .B(new_n3415), .Y(po0005));
  not_8  g01074(.A(pi303), .Y(new_n3423));
  not_8  g01075(.A(pi089), .Y(new_n3424));
  xor_4  g01076(.A(pi118), .B(new_n3424), .Y(new_n3425));
  not_8  g01077(.A(pi227), .Y(new_n3426));
  nand_5 g01078(.A(pi466), .B(new_n3426), .Y(new_n3427));
  xor_4  g01079(.A(pi466), .B(new_n3426), .Y(new_n3428));
  not_8  g01080(.A(pi436), .Y(new_n3429));
  nand_5 g01081(.A(pi553), .B(new_n3429), .Y(new_n3430));
  xor_4  g01082(.A(pi553), .B(new_n3429), .Y(new_n3431));
  not_8  g01083(.A(pi008), .Y(new_n3432));
  nand_5 g01084(.A(pi757), .B(new_n3432), .Y(new_n3433));
  xor_4  g01085(.A(pi757), .B(new_n3432), .Y(new_n3434));
  not_8  g01086(.A(pi155), .Y(new_n3435));
  nand_5 g01087(.A(pi531), .B(new_n3435), .Y(new_n3436));
  xor_4  g01088(.A(pi531), .B(new_n3435), .Y(new_n3437));
  not_8  g01089(.A(pi011), .Y(new_n3438));
  nand_5 g01090(.A(pi464), .B(new_n3438), .Y(new_n3439));
  xor_4  g01091(.A(pi464), .B(new_n3438), .Y(new_n3440));
  not_8  g01092(.A(pi518), .Y(new_n3441));
  nand_5 g01093(.A(new_n3441), .B(pi330), .Y(new_n3442));
  not_8  g01094(.A(pi330), .Y(new_n3443));
  xor_4  g01095(.A(pi518), .B(new_n3443), .Y(new_n3444));
  not_8  g01096(.A(pi510), .Y(new_n3445));
  nand_5 g01097(.A(pi523), .B(new_n3445), .Y(new_n3446));
  xor_4  g01098(.A(pi523), .B(new_n3445), .Y(new_n3447));
  not_8  g01099(.A(pi230), .Y(new_n3448));
  nand_5 g01100(.A(pi301), .B(new_n3448), .Y(new_n3449));
  not_8  g01101(.A(new_n3449), .Y(new_n3450));
  nand_5 g01102(.A(new_n3450), .B(new_n3447), .Y(new_n3451));
  nand_5 g01103(.A(new_n3451), .B(new_n3446), .Y(new_n3452));
  nand_5 g01104(.A(new_n3452), .B(new_n3444), .Y(new_n3453));
  nand_5 g01105(.A(new_n3453), .B(new_n3442), .Y(new_n3454));
  nand_5 g01106(.A(new_n3454), .B(new_n3440), .Y(new_n3455));
  nand_5 g01107(.A(new_n3455), .B(new_n3439), .Y(new_n3456));
  nand_5 g01108(.A(new_n3456), .B(new_n3437), .Y(new_n3457));
  nand_5 g01109(.A(new_n3457), .B(new_n3436), .Y(new_n3458));
  nand_5 g01110(.A(new_n3458), .B(pi655), .Y(new_n3459));
  not_8  g01111(.A(pi655), .Y(new_n3460));
  xor_4  g01112(.A(new_n3458), .B(new_n3460), .Y(new_n3461));
  or_6   g01113(.A(new_n3461), .B(pi300), .Y(new_n3462));
  nand_5 g01114(.A(new_n3462), .B(new_n3459), .Y(new_n3463));
  nand_5 g01115(.A(new_n3463), .B(new_n3434), .Y(new_n3464));
  nand_5 g01116(.A(new_n3464), .B(new_n3433), .Y(new_n3465));
  nand_5 g01117(.A(new_n3465), .B(new_n3431), .Y(new_n3466));
  nand_5 g01118(.A(new_n3466), .B(new_n3430), .Y(new_n3467));
  nand_5 g01119(.A(new_n3467), .B(new_n3428), .Y(new_n3468));
  nand_5 g01120(.A(new_n3468), .B(new_n3427), .Y(new_n3469));
  xnor_4 g01121(.A(new_n3469), .B(new_n3425), .Y(new_n3470));
  xor_4  g01122(.A(new_n3470), .B(new_n3423), .Y(new_n3471));
  not_8  g01123(.A(new_n3471), .Y(new_n3472));
  not_8  g01124(.A(pi650), .Y(new_n3473));
  xor_4  g01125(.A(new_n3467), .B(new_n3428), .Y(new_n3474));
  not_8  g01126(.A(new_n3474), .Y(new_n3475));
  nand_5 g01127(.A(new_n3475), .B(new_n3473), .Y(new_n3476));
  xor_4  g01128(.A(new_n3465), .B(new_n3431), .Y(new_n3477));
  nand_5 g01129(.A(new_n3477), .B(pi616), .Y(new_n3478));
  xor_4  g01130(.A(new_n3477), .B(pi616), .Y(new_n3479));
  xor_4  g01131(.A(new_n3463), .B(new_n3434), .Y(new_n3480));
  nor_5  g01132(.A(new_n3480), .B(pi441), .Y(new_n3481));
  xor_4  g01133(.A(new_n3461), .B(pi300), .Y(new_n3482));
  nor_5  g01134(.A(new_n3482), .B(pi246), .Y(new_n3483));
  not_8  g01135(.A(pi246), .Y(new_n3484));
  xor_4  g01136(.A(pi300), .B(new_n3484), .Y(new_n3485));
  xor_4  g01137(.A(new_n3485), .B(new_n3461), .Y(new_n3486));
  xor_4  g01138(.A(new_n3456), .B(new_n3437), .Y(new_n3487));
  xor_4  g01139(.A(new_n3454), .B(new_n3440), .Y(new_n3488));
  not_8  g01140(.A(pi361), .Y(new_n3489));
  xor_4  g01141(.A(new_n3449), .B(new_n3447), .Y(new_n3490));
  not_8  g01142(.A(pi301), .Y(new_n3491));
  nand_5 g01143(.A(new_n3491), .B(pi230), .Y(new_n3492));
  not_8  g01144(.A(pi670), .Y(new_n3493));
  nand_5 g01145(.A(new_n3449), .B(new_n3493), .Y(new_n3494));
  nand_5 g01146(.A(new_n3494), .B(new_n3492), .Y(new_n3495));
  xor_4  g01147(.A(new_n3495), .B(new_n3447), .Y(new_n3496));
  nand_5 g01148(.A(new_n3496), .B(new_n3490), .Y(new_n3497));
  or_6   g01149(.A(new_n3496), .B(pi787), .Y(new_n3498));
  nand_5 g01150(.A(new_n3498), .B(new_n3497), .Y(new_n3499));
  or_6   g01151(.A(new_n3499), .B(new_n3489), .Y(new_n3500));
  xor_4  g01152(.A(new_n3452), .B(new_n3444), .Y(new_n3501));
  xor_4  g01153(.A(new_n3499), .B(new_n3489), .Y(new_n3502));
  nand_5 g01154(.A(new_n3502), .B(new_n3501), .Y(new_n3503));
  nand_5 g01155(.A(new_n3503), .B(new_n3500), .Y(new_n3504));
  nand_5 g01156(.A(new_n3504), .B(new_n3488), .Y(new_n3505));
  or_6   g01157(.A(new_n3504), .B(new_n3488), .Y(new_n3506));
  nand_5 g01158(.A(new_n3506), .B(pi681), .Y(new_n3507));
  nand_5 g01159(.A(new_n3507), .B(new_n3505), .Y(new_n3508));
  nand_5 g01160(.A(new_n3508), .B(new_n3487), .Y(new_n3509));
  or_6   g01161(.A(new_n3508), .B(new_n3487), .Y(new_n3510));
  nand_5 g01162(.A(new_n3510), .B(pi317), .Y(new_n3511));
  nand_5 g01163(.A(new_n3511), .B(new_n3509), .Y(new_n3512));
  nor_5  g01164(.A(new_n3512), .B(new_n3486), .Y(new_n3513));
  nor_5  g01165(.A(new_n3513), .B(new_n3483), .Y(new_n3514));
  and_6  g01166(.A(new_n3480), .B(pi441), .Y(new_n3515));
  nor_5  g01167(.A(new_n3515), .B(new_n3514), .Y(new_n3516));
  nor_5  g01168(.A(new_n3516), .B(new_n3481), .Y(new_n3517));
  nand_5 g01169(.A(new_n3517), .B(new_n3479), .Y(new_n3518));
  nand_5 g01170(.A(new_n3518), .B(new_n3478), .Y(new_n3519));
  xor_4  g01171(.A(new_n3474), .B(new_n3473), .Y(new_n3520));
  or_6   g01172(.A(new_n3520), .B(new_n3519), .Y(new_n3521));
  nand_5 g01173(.A(new_n3521), .B(new_n3476), .Y(new_n3522));
  xor_4  g01174(.A(new_n3522), .B(new_n3472), .Y(new_n3523));
  not_8  g01175(.A(pi740), .Y(new_n3524));
  not_8  g01176(.A(pi446), .Y(new_n3525));
  nand_5 g01177(.A(new_n3525), .B(pi331), .Y(new_n3526));
  not_8  g01178(.A(pi331), .Y(new_n3527));
  nand_5 g01179(.A(pi446), .B(new_n3527), .Y(new_n3528));
  nand_5 g01180(.A(new_n3528), .B(new_n3526), .Y(new_n3529));
  not_8  g01181(.A(pi507), .Y(new_n3530));
  nand_5 g01182(.A(new_n3530), .B(pi428), .Y(new_n3531));
  not_8  g01183(.A(new_n3531), .Y(new_n3532));
  not_8  g01184(.A(pi428), .Y(new_n3533));
  xor_4  g01185(.A(pi507), .B(new_n3533), .Y(new_n3534));
  not_8  g01186(.A(new_n3534), .Y(new_n3535));
  not_8  g01187(.A(pi196), .Y(new_n3536));
  nand_5 g01188(.A(pi324), .B(new_n3536), .Y(new_n3537));
  nand_5 g01189(.A(new_n2468), .B(pi196), .Y(new_n3538));
  not_8  g01190(.A(pi138), .Y(new_n3539));
  nand_5 g01191(.A(pi790), .B(new_n3539), .Y(new_n3540));
  not_8  g01192(.A(new_n3540), .Y(new_n3541));
  not_8  g01193(.A(pi453), .Y(new_n3542));
  nand_5 g01194(.A(new_n3542), .B(pi316), .Y(new_n3543));
  not_8  g01195(.A(new_n3543), .Y(new_n3544));
  not_8  g01196(.A(pi421), .Y(new_n3545));
  nand_5 g01197(.A(new_n3545), .B(pi102), .Y(new_n3546));
  not_8  g01198(.A(new_n3546), .Y(new_n3547));
  xor_4  g01199(.A(pi421), .B(new_n2478), .Y(new_n3548));
  not_8  g01200(.A(new_n3548), .Y(new_n3549));
  nand_5 g01201(.A(pi626), .B(new_n2482), .Y(new_n3550));
  or_6   g01202(.A(pi626), .B(new_n2482), .Y(new_n3551));
  not_8  g01203(.A(pi612), .Y(new_n3552));
  nand_5 g01204(.A(new_n3552), .B(pi045), .Y(new_n3553));
  not_8  g01205(.A(pi045), .Y(new_n3554));
  nand_5 g01206(.A(pi612), .B(new_n3554), .Y(new_n3555));
  not_8  g01207(.A(pi520), .Y(new_n3556));
  nand_5 g01208(.A(new_n3556), .B(pi302), .Y(new_n3557));
  nand_5 g01209(.A(new_n3557), .B(new_n3555), .Y(new_n3558));
  nand_5 g01210(.A(new_n3558), .B(new_n3553), .Y(new_n3559));
  nand_5 g01211(.A(new_n3559), .B(new_n3551), .Y(new_n3560));
  nand_5 g01212(.A(new_n3560), .B(new_n3550), .Y(new_n3561));
  nor_5  g01213(.A(new_n3561), .B(new_n3549), .Y(new_n3562));
  nor_5  g01214(.A(new_n3562), .B(new_n3547), .Y(new_n3563));
  xor_4  g01215(.A(pi453), .B(pi316), .Y(new_n3564));
  nor_5  g01216(.A(new_n3564), .B(new_n3563), .Y(new_n3565));
  nor_5  g01217(.A(new_n3565), .B(new_n3544), .Y(new_n3566));
  xor_4  g01218(.A(pi790), .B(pi138), .Y(new_n3567));
  nor_5  g01219(.A(new_n3567), .B(new_n3566), .Y(new_n3568));
  nor_5  g01220(.A(new_n3568), .B(new_n3541), .Y(new_n3569));
  not_8  g01221(.A(new_n3569), .Y(new_n3570));
  nand_5 g01222(.A(new_n3570), .B(new_n3538), .Y(new_n3571));
  nand_5 g01223(.A(new_n3571), .B(new_n3537), .Y(new_n3572));
  nor_5  g01224(.A(new_n3572), .B(new_n3535), .Y(new_n3573));
  nor_5  g01225(.A(new_n3573), .B(new_n3532), .Y(new_n3574));
  not_8  g01226(.A(new_n3574), .Y(new_n3575));
  xor_4  g01227(.A(new_n3575), .B(new_n3529), .Y(new_n3576));
  xor_4  g01228(.A(new_n3576), .B(new_n3524), .Y(new_n3577));
  xor_4  g01229(.A(new_n3572), .B(new_n3534), .Y(new_n3578));
  xor_4  g01230(.A(new_n3564), .B(new_n3563), .Y(new_n3579));
  xor_4  g01231(.A(new_n3561), .B(new_n3549), .Y(new_n3580));
  not_8  g01232(.A(pi458), .Y(new_n3581));
  and_6  g01233(.A(new_n3555), .B(new_n3553), .Y(new_n3582));
  xor_4  g01234(.A(new_n3582), .B(new_n3557), .Y(new_n3583));
  nand_5 g01235(.A(new_n3583), .B(pi288), .Y(new_n3584));
  nand_5 g01236(.A(new_n3584), .B(new_n3581), .Y(new_n3585));
  xor_4  g01237(.A(new_n3584), .B(pi458), .Y(new_n3586));
  nand_5 g01238(.A(new_n3551), .B(new_n3550), .Y(new_n3587));
  xor_4  g01239(.A(new_n3587), .B(new_n3559), .Y(new_n3588));
  not_8  g01240(.A(new_n3588), .Y(new_n3589));
  or_6   g01241(.A(new_n3589), .B(new_n3586), .Y(new_n3590));
  nand_5 g01242(.A(new_n3590), .B(new_n3585), .Y(new_n3591));
  nor_5  g01243(.A(new_n3591), .B(new_n3580), .Y(new_n3592));
  nand_5 g01244(.A(new_n3591), .B(new_n3580), .Y(new_n3593));
  nand_5 g01245(.A(new_n3593), .B(pi152), .Y(new_n3594));
  not_8  g01246(.A(new_n3594), .Y(new_n3595));
  nor_5  g01247(.A(new_n3595), .B(new_n3592), .Y(new_n3596));
  nand_5 g01248(.A(new_n3596), .B(new_n3579), .Y(new_n3597));
  not_8  g01249(.A(pi037), .Y(new_n3598));
  xor_4  g01250(.A(new_n3596), .B(new_n3579), .Y(new_n3599));
  nand_5 g01251(.A(new_n3599), .B(new_n3598), .Y(new_n3600));
  nand_5 g01252(.A(new_n3600), .B(new_n3597), .Y(new_n3601));
  xor_4  g01253(.A(new_n3567), .B(new_n3566), .Y(new_n3602));
  nand_5 g01254(.A(new_n3602), .B(new_n3601), .Y(new_n3603));
  not_8  g01255(.A(pi585), .Y(new_n3604));
  or_6   g01256(.A(new_n3602), .B(new_n3601), .Y(new_n3605));
  nand_5 g01257(.A(new_n3605), .B(new_n3604), .Y(new_n3606));
  nand_5 g01258(.A(new_n3606), .B(new_n3603), .Y(new_n3607));
  and_6  g01259(.A(new_n3538), .B(new_n3537), .Y(new_n3608));
  xor_4  g01260(.A(new_n3608), .B(new_n3570), .Y(new_n3609));
  nor_5  g01261(.A(new_n3609), .B(new_n3607), .Y(new_n3610));
  not_8  g01262(.A(pi717), .Y(new_n3611));
  not_8  g01263(.A(new_n3609), .Y(new_n3612));
  xor_4  g01264(.A(new_n3612), .B(new_n3607), .Y(new_n3613));
  nor_5  g01265(.A(new_n3613), .B(new_n3611), .Y(new_n3614));
  nor_5  g01266(.A(new_n3614), .B(new_n3610), .Y(new_n3615));
  or_6   g01267(.A(new_n3615), .B(new_n3578), .Y(new_n3616));
  xor_4  g01268(.A(new_n3615), .B(new_n3578), .Y(new_n3617));
  nand_5 g01269(.A(new_n3617), .B(pi409), .Y(new_n3618));
  nand_5 g01270(.A(new_n3618), .B(new_n3616), .Y(new_n3619));
  xor_4  g01271(.A(new_n3619), .B(new_n3577), .Y(new_n3620));
  not_8  g01272(.A(new_n3620), .Y(new_n3621));
  not_8  g01273(.A(pi409), .Y(new_n3622));
  xor_4  g01274(.A(new_n3617), .B(new_n3622), .Y(new_n3623));
  xor_4  g01275(.A(new_n3599), .B(pi037), .Y(new_n3624));
  xor_4  g01276(.A(new_n3502), .B(new_n3501), .Y(new_n3625));
  not_8  g01277(.A(new_n3625), .Y(new_n3626));
  xor_4  g01278(.A(new_n3583), .B(pi288), .Y(new_n3627));
  not_8  g01279(.A(new_n3627), .Y(new_n3628));
  not_8  g01280(.A(pi787), .Y(new_n3629));
  xor_4  g01281(.A(new_n3496), .B(new_n3629), .Y(new_n3630));
  nor_5  g01282(.A(new_n3630), .B(new_n3628), .Y(new_n3631));
  xor_4  g01283(.A(new_n3630), .B(new_n3628), .Y(new_n3632));
  not_8  g01284(.A(new_n3632), .Y(new_n3633));
  nand_5 g01285(.A(new_n3493), .B(pi230), .Y(new_n3634));
  nand_5 g01286(.A(pi670), .B(new_n3448), .Y(new_n3635));
  nand_5 g01287(.A(new_n3635), .B(new_n3634), .Y(new_n3636));
  not_8  g01288(.A(new_n3636), .Y(new_n3637));
  xor_4  g01289(.A(pi559), .B(new_n3491), .Y(new_n3638));
  xor_4  g01290(.A(new_n3638), .B(new_n3637), .Y(new_n3639));
  or_6   g01291(.A(new_n3639), .B(pi559), .Y(new_n3640));
  not_8  g01292(.A(pi302), .Y(new_n3641));
  xor_4  g01293(.A(pi520), .B(new_n3641), .Y(new_n3642));
  nand_5 g01294(.A(new_n3642), .B(new_n3639), .Y(new_n3643));
  nand_5 g01295(.A(new_n3643), .B(new_n3640), .Y(new_n3644));
  nor_5  g01296(.A(new_n3644), .B(new_n3633), .Y(new_n3645));
  or_6   g01297(.A(new_n3645), .B(new_n3631), .Y(new_n3646));
  nand_5 g01298(.A(new_n3646), .B(new_n3626), .Y(new_n3647));
  xor_4  g01299(.A(new_n3588), .B(new_n3586), .Y(new_n3648));
  xor_4  g01300(.A(new_n3646), .B(new_n3626), .Y(new_n3649));
  nand_5 g01301(.A(new_n3649), .B(new_n3648), .Y(new_n3650));
  nand_5 g01302(.A(new_n3650), .B(new_n3647), .Y(new_n3651));
  nand_5 g01303(.A(new_n3506), .B(new_n3505), .Y(new_n3652));
  xor_4  g01304(.A(new_n3652), .B(pi681), .Y(new_n3653));
  nand_5 g01305(.A(new_n3653), .B(new_n3651), .Y(new_n3654));
  xor_4  g01306(.A(new_n3653), .B(new_n3651), .Y(new_n3655));
  not_8  g01307(.A(pi152), .Y(new_n3656));
  xor_4  g01308(.A(new_n3591), .B(new_n3580), .Y(new_n3657));
  xor_4  g01309(.A(new_n3657), .B(new_n3656), .Y(new_n3658));
  not_8  g01310(.A(new_n3658), .Y(new_n3659));
  nand_5 g01311(.A(new_n3659), .B(new_n3655), .Y(new_n3660));
  nand_5 g01312(.A(new_n3660), .B(new_n3654), .Y(new_n3661));
  nor_5  g01313(.A(new_n3661), .B(new_n3624), .Y(new_n3662));
  nand_5 g01314(.A(new_n3510), .B(new_n3509), .Y(new_n3663));
  xor_4  g01315(.A(new_n3663), .B(pi317), .Y(new_n3664));
  xnor_4 g01316(.A(new_n3661), .B(new_n3624), .Y(new_n3665));
  nor_5  g01317(.A(new_n3665), .B(new_n3664), .Y(new_n3666));
  or_6   g01318(.A(new_n3666), .B(new_n3662), .Y(new_n3667));
  nand_5 g01319(.A(new_n3605), .B(new_n3603), .Y(new_n3668));
  xor_4  g01320(.A(new_n3668), .B(pi585), .Y(new_n3669));
  nand_5 g01321(.A(new_n3669), .B(new_n3667), .Y(new_n3670));
  xnor_4 g01322(.A(new_n3669), .B(new_n3667), .Y(new_n3671));
  xor_4  g01323(.A(new_n3512), .B(new_n3486), .Y(new_n3672));
  or_6   g01324(.A(new_n3672), .B(new_n3671), .Y(new_n3673));
  nand_5 g01325(.A(new_n3673), .B(new_n3670), .Y(new_n3674));
  xor_4  g01326(.A(new_n3613), .B(pi717), .Y(new_n3675));
  nand_5 g01327(.A(new_n3675), .B(new_n3674), .Y(new_n3676));
  xnor_4 g01328(.A(new_n3675), .B(new_n3674), .Y(new_n3677));
  or_6   g01329(.A(new_n3515), .B(new_n3481), .Y(new_n3678));
  xor_4  g01330(.A(new_n3678), .B(new_n3514), .Y(new_n3679));
  or_6   g01331(.A(new_n3679), .B(new_n3677), .Y(new_n3680));
  nand_5 g01332(.A(new_n3680), .B(new_n3676), .Y(new_n3681));
  nand_5 g01333(.A(new_n3681), .B(new_n3623), .Y(new_n3682));
  xnor_4 g01334(.A(new_n3517), .B(new_n3479), .Y(new_n3683));
  xnor_4 g01335(.A(new_n3681), .B(new_n3623), .Y(new_n3684));
  or_6   g01336(.A(new_n3684), .B(new_n3683), .Y(new_n3685));
  nand_5 g01337(.A(new_n3685), .B(new_n3682), .Y(new_n3686));
  nand_5 g01338(.A(new_n3686), .B(new_n3621), .Y(new_n3687));
  xor_4  g01339(.A(new_n3686), .B(new_n3620), .Y(new_n3688));
  xor_4  g01340(.A(new_n3520), .B(new_n3519), .Y(new_n3689));
  or_6   g01341(.A(new_n3689), .B(new_n3688), .Y(new_n3690));
  nand_5 g01342(.A(new_n3690), .B(new_n3687), .Y(new_n3691));
  or_6   g01343(.A(new_n3576), .B(new_n3524), .Y(new_n3692));
  nand_5 g01344(.A(new_n3619), .B(new_n3577), .Y(new_n3693));
  nand_5 g01345(.A(new_n3693), .B(new_n3692), .Y(new_n3694));
  not_8  g01346(.A(pi785), .Y(new_n3695));
  nand_5 g01347(.A(new_n3695), .B(pi293), .Y(new_n3696));
  not_8  g01348(.A(pi293), .Y(new_n3697));
  nand_5 g01349(.A(pi785), .B(new_n3697), .Y(new_n3698));
  nand_5 g01350(.A(new_n3698), .B(new_n3696), .Y(new_n3699));
  nand_5 g01351(.A(new_n3575), .B(new_n3528), .Y(new_n3700));
  nand_5 g01352(.A(new_n3700), .B(new_n3526), .Y(new_n3701));
  xnor_4 g01353(.A(new_n3701), .B(new_n3699), .Y(new_n3702));
  and_6  g01354(.A(new_n3702), .B(new_n3694), .Y(new_n3703));
  nor_5  g01355(.A(new_n3702), .B(new_n3694), .Y(new_n3704));
  or_6   g01356(.A(new_n3704), .B(new_n3703), .Y(new_n3705));
  xor_4  g01357(.A(new_n3705), .B(pi807), .Y(new_n3706));
  xnor_4 g01358(.A(new_n3706), .B(new_n3691), .Y(new_n3707));
  xor_4  g01359(.A(new_n3707), .B(new_n3523), .Y(po0006));
  not_8  g01360(.A(pi793), .Y(new_n3709));
  not_8  g01361(.A(pi064), .Y(new_n3710));
  xor_4  g01362(.A(pi583), .B(new_n3710), .Y(new_n3711));
  not_8  g01363(.A(pi695), .Y(new_n3712));
  nand_5 g01364(.A(new_n3712), .B(pi641), .Y(new_n3713));
  not_8  g01365(.A(pi641), .Y(new_n3714));
  xor_4  g01366(.A(pi695), .B(new_n3714), .Y(new_n3715));
  not_8  g01367(.A(pi805), .Y(new_n3716));
  nand_5 g01368(.A(new_n3716), .B(pi201), .Y(new_n3717));
  not_8  g01369(.A(pi201), .Y(new_n3718));
  xor_4  g01370(.A(pi805), .B(new_n3718), .Y(new_n3719));
  not_8  g01371(.A(pi006), .Y(new_n3720));
  nand_5 g01372(.A(pi795), .B(new_n3720), .Y(new_n3721));
  xor_4  g01373(.A(pi795), .B(new_n3720), .Y(new_n3722));
  not_8  g01374(.A(pi495), .Y(new_n3723));
  nor_5  g01375(.A(pi818), .B(new_n3723), .Y(new_n3724));
  xor_4  g01376(.A(pi818), .B(pi495), .Y(new_n3725));
  not_8  g01377(.A(pi422), .Y(new_n3726));
  nand_5 g01378(.A(new_n3726), .B(pi158), .Y(new_n3727));
  not_8  g01379(.A(pi158), .Y(new_n3728));
  nand_5 g01380(.A(pi422), .B(new_n3728), .Y(new_n3729));
  not_8  g01381(.A(pi259), .Y(new_n3730));
  nand_5 g01382(.A(pi781), .B(new_n3730), .Y(new_n3731));
  nand_5 g01383(.A(new_n3731), .B(new_n3729), .Y(new_n3732));
  nand_5 g01384(.A(new_n3732), .B(new_n3727), .Y(new_n3733));
  nor_5  g01385(.A(new_n3733), .B(new_n3725), .Y(new_n3734));
  nor_5  g01386(.A(new_n3734), .B(new_n3724), .Y(new_n3735));
  not_8  g01387(.A(new_n3735), .Y(new_n3736));
  nand_5 g01388(.A(new_n3736), .B(new_n3722), .Y(new_n3737));
  nand_5 g01389(.A(new_n3737), .B(new_n3721), .Y(new_n3738));
  nand_5 g01390(.A(new_n3738), .B(new_n3719), .Y(new_n3739));
  nand_5 g01391(.A(new_n3739), .B(new_n3717), .Y(new_n3740));
  nand_5 g01392(.A(new_n3740), .B(new_n3715), .Y(new_n3741));
  nand_5 g01393(.A(new_n3741), .B(new_n3713), .Y(new_n3742));
  xor_4  g01394(.A(new_n3742), .B(new_n3711), .Y(new_n3743));
  xor_4  g01395(.A(new_n3738), .B(new_n3719), .Y(new_n3744));
  not_8  g01396(.A(new_n3744), .Y(new_n3745));
  not_8  g01397(.A(pi241), .Y(new_n3746));
  nand_5 g01398(.A(new_n3729), .B(new_n3727), .Y(new_n3747));
  xnor_4 g01399(.A(new_n3747), .B(new_n3731), .Y(new_n3748));
  nand_5 g01400(.A(new_n3748), .B(pi488), .Y(new_n3749));
  nor_5  g01401(.A(new_n3749), .B(new_n3746), .Y(new_n3750));
  xor_4  g01402(.A(new_n3749), .B(new_n3746), .Y(new_n3751));
  not_8  g01403(.A(new_n3751), .Y(new_n3752));
  xor_4  g01404(.A(new_n3733), .B(new_n3725), .Y(new_n3753));
  nor_5  g01405(.A(new_n3753), .B(new_n3752), .Y(new_n3754));
  or_6   g01406(.A(new_n3754), .B(new_n3750), .Y(new_n3755));
  xor_4  g01407(.A(new_n3735), .B(new_n3722), .Y(new_n3756));
  nand_5 g01408(.A(new_n3756), .B(new_n3755), .Y(new_n3757));
  not_8  g01409(.A(pi157), .Y(new_n3758));
  xnor_4 g01410(.A(new_n3756), .B(new_n3755), .Y(new_n3759));
  or_6   g01411(.A(new_n3759), .B(new_n3758), .Y(new_n3760));
  nand_5 g01412(.A(new_n3760), .B(new_n3757), .Y(new_n3761));
  nand_5 g01413(.A(new_n3761), .B(new_n3745), .Y(new_n3762));
  not_8  g01414(.A(pi298), .Y(new_n3763));
  xor_4  g01415(.A(new_n3761), .B(new_n3744), .Y(new_n3764));
  or_6   g01416(.A(new_n3764), .B(new_n3763), .Y(new_n3765));
  nand_5 g01417(.A(new_n3765), .B(new_n3762), .Y(new_n3766));
  xnor_4 g01418(.A(new_n3740), .B(new_n3715), .Y(new_n3767));
  or_6   g01419(.A(new_n3767), .B(new_n3766), .Y(new_n3768));
  nand_5 g01420(.A(new_n3768), .B(pi103), .Y(new_n3769));
  nand_5 g01421(.A(new_n3767), .B(new_n3766), .Y(new_n3770));
  nand_5 g01422(.A(new_n3770), .B(new_n3769), .Y(new_n3771));
  xor_4  g01423(.A(new_n3771), .B(new_n3743), .Y(new_n3772));
  xor_4  g01424(.A(new_n3772), .B(new_n3709), .Y(new_n3773));
  not_8  g01425(.A(pi567), .Y(new_n3774));
  nand_5 g01426(.A(pi709), .B(new_n3774), .Y(new_n3775));
  xor_4  g01427(.A(pi709), .B(new_n3774), .Y(new_n3776));
  nand_5 g01428(.A(pi590), .B(new_n2373), .Y(new_n3777));
  xor_4  g01429(.A(pi590), .B(new_n2373), .Y(new_n3778));
  not_8  g01430(.A(pi605), .Y(new_n3779));
  nand_5 g01431(.A(new_n3779), .B(pi328), .Y(new_n3780));
  xor_4  g01432(.A(pi605), .B(new_n2948), .Y(new_n3781));
  nand_5 g01433(.A(new_n2357), .B(pi277), .Y(new_n3782));
  xor_4  g01434(.A(pi434), .B(new_n2960), .Y(new_n3783));
  nand_5 g01435(.A(new_n2361), .B(pi313), .Y(new_n3784));
  not_8  g01436(.A(pi313), .Y(new_n3785));
  xor_4  g01437(.A(pi552), .B(new_n3785), .Y(new_n3786));
  nand_5 g01438(.A(pi832), .B(new_n2419), .Y(new_n3787));
  not_8  g01439(.A(new_n3787), .Y(new_n3788));
  nand_5 g01440(.A(new_n3788), .B(new_n3786), .Y(new_n3789));
  nand_5 g01441(.A(new_n3789), .B(new_n3784), .Y(new_n3790));
  nand_5 g01442(.A(new_n3790), .B(new_n3783), .Y(new_n3791));
  nand_5 g01443(.A(new_n3791), .B(new_n3782), .Y(new_n3792));
  nand_5 g01444(.A(new_n3792), .B(new_n3781), .Y(new_n3793));
  nand_5 g01445(.A(new_n3793), .B(new_n3780), .Y(new_n3794));
  nand_5 g01446(.A(new_n3794), .B(new_n3778), .Y(new_n3795));
  nand_5 g01447(.A(new_n3795), .B(new_n3777), .Y(new_n3796));
  nand_5 g01448(.A(new_n3796), .B(new_n3776), .Y(new_n3797));
  nand_5 g01449(.A(new_n3797), .B(new_n3775), .Y(new_n3798));
  not_8  g01450(.A(pi683), .Y(new_n3799));
  nand_5 g01451(.A(pi816), .B(new_n3799), .Y(new_n3800));
  nand_5 g01452(.A(new_n2944), .B(pi683), .Y(new_n3801));
  and_6  g01453(.A(new_n3801), .B(new_n3800), .Y(new_n3802));
  xor_4  g01454(.A(new_n3802), .B(new_n3798), .Y(new_n3803));
  not_8  g01455(.A(new_n3803), .Y(new_n3804));
  not_8  g01456(.A(pi177), .Y(new_n3805));
  xnor_4 g01457(.A(new_n3796), .B(new_n3776), .Y(new_n3806));
  nor_5  g01458(.A(new_n3806), .B(new_n3805), .Y(new_n3807));
  xor_4  g01459(.A(new_n3806), .B(new_n3805), .Y(new_n3808));
  not_8  g01460(.A(new_n3808), .Y(new_n3809));
  xnor_4 g01461(.A(new_n3794), .B(new_n3778), .Y(new_n3810));
  not_8  g01462(.A(pi027), .Y(new_n3811));
  xor_4  g01463(.A(new_n3792), .B(new_n3781), .Y(new_n3812));
  not_8  g01464(.A(new_n3812), .Y(new_n3813));
  not_8  g01465(.A(pi672), .Y(new_n3814));
  not_8  g01466(.A(pi832), .Y(new_n3815));
  nand_5 g01467(.A(new_n3815), .B(pi190), .Y(new_n3816));
  nand_5 g01468(.A(new_n3816), .B(new_n3787), .Y(new_n3817));
  not_8  g01469(.A(new_n3817), .Y(new_n3818));
  nand_5 g01470(.A(new_n3818), .B(pi385), .Y(new_n3819));
  not_8  g01471(.A(new_n3819), .Y(new_n3820));
  nor_5  g01472(.A(new_n3820), .B(new_n3788), .Y(new_n3821));
  xor_4  g01473(.A(new_n3821), .B(new_n3786), .Y(new_n3822));
  or_6   g01474(.A(new_n3822), .B(new_n3814), .Y(new_n3823));
  nand_5 g01475(.A(new_n3820), .B(new_n3786), .Y(new_n3824));
  nand_5 g01476(.A(new_n3824), .B(new_n3823), .Y(new_n3825));
  nor_5  g01477(.A(new_n3825), .B(pi597), .Y(new_n3826));
  xor_4  g01478(.A(new_n3790), .B(new_n3783), .Y(new_n3827));
  not_8  g01479(.A(pi597), .Y(new_n3828));
  xor_4  g01480(.A(new_n3825), .B(new_n3828), .Y(new_n3829));
  nor_5  g01481(.A(new_n3829), .B(new_n3827), .Y(new_n3830));
  or_6   g01482(.A(new_n3830), .B(new_n3826), .Y(new_n3831));
  or_6   g01483(.A(new_n3831), .B(new_n3813), .Y(new_n3832));
  nand_5 g01484(.A(new_n3832), .B(new_n3811), .Y(new_n3833));
  nand_5 g01485(.A(new_n3831), .B(new_n3813), .Y(new_n3834));
  nand_5 g01486(.A(new_n3834), .B(new_n3833), .Y(new_n3835));
  nand_5 g01487(.A(new_n3835), .B(new_n3810), .Y(new_n3836));
  xnor_4 g01488(.A(new_n3835), .B(new_n3810), .Y(new_n3837));
  or_6   g01489(.A(new_n3837), .B(pi012), .Y(new_n3838));
  nand_5 g01490(.A(new_n3838), .B(new_n3836), .Y(new_n3839));
  nor_5  g01491(.A(new_n3839), .B(new_n3809), .Y(new_n3840));
  nor_5  g01492(.A(new_n3840), .B(new_n3807), .Y(new_n3841));
  or_6   g01493(.A(new_n3841), .B(new_n3804), .Y(new_n3842));
  nand_5 g01494(.A(new_n3841), .B(new_n3804), .Y(new_n3843));
  nand_5 g01495(.A(new_n3843), .B(new_n3842), .Y(new_n3844));
  xor_4  g01496(.A(new_n3844), .B(pi143), .Y(new_n3845));
  not_8  g01497(.A(pi012), .Y(new_n3846));
  xor_4  g01498(.A(new_n3837), .B(new_n3846), .Y(new_n3847));
  xor_4  g01499(.A(new_n3764), .B(new_n3763), .Y(new_n3848));
  not_8  g01500(.A(new_n3848), .Y(new_n3849));
  nand_5 g01501(.A(new_n3849), .B(new_n3847), .Y(new_n3850));
  xor_4  g01502(.A(new_n3848), .B(new_n3847), .Y(new_n3851));
  xor_4  g01503(.A(new_n3759), .B(new_n3758), .Y(new_n3852));
  not_8  g01504(.A(new_n3852), .Y(new_n3853));
  xor_4  g01505(.A(new_n3753), .B(new_n3752), .Y(new_n3854));
  not_8  g01506(.A(new_n3854), .Y(new_n3855));
  xor_4  g01507(.A(new_n3822), .B(new_n3814), .Y(new_n3856));
  not_8  g01508(.A(new_n3856), .Y(new_n3857));
  xor_4  g01509(.A(new_n3748), .B(pi488), .Y(new_n3858));
  nor_5  g01510(.A(new_n3858), .B(new_n3857), .Y(new_n3859));
  not_8  g01511(.A(pi631), .Y(new_n3860));
  xor_4  g01512(.A(pi781), .B(new_n3730), .Y(new_n3861));
  or_6   g01513(.A(new_n3861), .B(new_n3860), .Y(new_n3862));
  not_8  g01514(.A(pi385), .Y(new_n3863));
  xor_4  g01515(.A(new_n3817), .B(new_n3863), .Y(new_n3864));
  not_8  g01516(.A(new_n3864), .Y(new_n3865));
  xor_4  g01517(.A(new_n3861), .B(new_n3860), .Y(new_n3866));
  nand_5 g01518(.A(new_n3866), .B(new_n3865), .Y(new_n3867));
  nand_5 g01519(.A(new_n3867), .B(new_n3862), .Y(new_n3868));
  xor_4  g01520(.A(new_n3858), .B(new_n3856), .Y(new_n3869));
  nor_5  g01521(.A(new_n3869), .B(new_n3868), .Y(new_n3870));
  or_6   g01522(.A(new_n3870), .B(new_n3859), .Y(new_n3871));
  nand_5 g01523(.A(new_n3871), .B(new_n3855), .Y(new_n3872));
  xor_4  g01524(.A(new_n3829), .B(new_n3827), .Y(new_n3873));
  xor_4  g01525(.A(new_n3871), .B(new_n3854), .Y(new_n3874));
  or_6   g01526(.A(new_n3874), .B(new_n3873), .Y(new_n3875));
  nand_5 g01527(.A(new_n3875), .B(new_n3872), .Y(new_n3876));
  and_6  g01528(.A(new_n3876), .B(new_n3853), .Y(new_n3877));
  nand_5 g01529(.A(new_n3834), .B(new_n3832), .Y(new_n3878));
  xor_4  g01530(.A(new_n3878), .B(pi027), .Y(new_n3879));
  xor_4  g01531(.A(new_n3876), .B(new_n3852), .Y(new_n3880));
  nor_5  g01532(.A(new_n3880), .B(new_n3879), .Y(new_n3881));
  nor_5  g01533(.A(new_n3881), .B(new_n3877), .Y(new_n3882));
  or_6   g01534(.A(new_n3882), .B(new_n3851), .Y(new_n3883));
  nand_5 g01535(.A(new_n3883), .B(new_n3850), .Y(new_n3884));
  nand_5 g01536(.A(new_n3770), .B(new_n3768), .Y(new_n3885));
  xor_4  g01537(.A(new_n3885), .B(pi103), .Y(new_n3886));
  nand_5 g01538(.A(new_n3886), .B(new_n3884), .Y(new_n3887));
  xor_4  g01539(.A(new_n3839), .B(new_n3808), .Y(new_n3888));
  xnor_4 g01540(.A(new_n3886), .B(new_n3884), .Y(new_n3889));
  or_6   g01541(.A(new_n3889), .B(new_n3888), .Y(new_n3890));
  nand_5 g01542(.A(new_n3890), .B(new_n3887), .Y(new_n3891));
  xor_4  g01543(.A(new_n3891), .B(new_n3845), .Y(new_n3892));
  xnor_4 g01544(.A(new_n3892), .B(new_n3773), .Y(po0007));
  not_8  g01545(.A(pi568), .Y(new_n3894));
  not_8  g01546(.A(pi497), .Y(new_n3895));
  xor_4  g01547(.A(new_n3895), .B(pi359), .Y(new_n3896));
  not_8  g01548(.A(pi506), .Y(new_n3897));
  nand_5 g01549(.A(new_n3897), .B(pi167), .Y(new_n3898));
  xor_4  g01550(.A(new_n3897), .B(pi167), .Y(new_n3899));
  not_8  g01551(.A(pi374), .Y(new_n3900));
  nand_5 g01552(.A(pi820), .B(new_n3900), .Y(new_n3901));
  not_8  g01553(.A(new_n3901), .Y(new_n3902));
  xor_4  g01554(.A(pi820), .B(new_n3900), .Y(new_n3903));
  not_8  g01555(.A(new_n3903), .Y(new_n3904));
  not_8  g01556(.A(pi688), .Y(new_n3905));
  or_6   g01557(.A(new_n3905), .B(pi376), .Y(new_n3906));
  nand_5 g01558(.A(pi648), .B(new_n2565), .Y(new_n3907));
  nand_5 g01559(.A(new_n3905), .B(pi376), .Y(new_n3908));
  nand_5 g01560(.A(new_n3908), .B(new_n3907), .Y(new_n3909));
  nand_5 g01561(.A(new_n3909), .B(new_n3906), .Y(new_n3910));
  nor_5  g01562(.A(new_n3910), .B(new_n3904), .Y(new_n3911));
  nor_5  g01563(.A(new_n3911), .B(new_n3902), .Y(new_n3912));
  not_8  g01564(.A(new_n3912), .Y(new_n3913));
  nand_5 g01565(.A(new_n3913), .B(new_n3899), .Y(new_n3914));
  nand_5 g01566(.A(new_n3914), .B(new_n3898), .Y(new_n3915));
  xor_4  g01567(.A(new_n3915), .B(new_n3896), .Y(new_n3916));
  xor_4  g01568(.A(new_n3916), .B(new_n3894), .Y(new_n3917));
  xor_4  g01569(.A(new_n3912), .B(new_n3899), .Y(new_n3918));
  not_8  g01570(.A(new_n3918), .Y(new_n3919));
  xor_4  g01571(.A(new_n3910), .B(new_n3903), .Y(new_n3920));
  not_8  g01572(.A(new_n3920), .Y(new_n3921));
  not_8  g01573(.A(pi245), .Y(new_n3922));
  not_8  g01574(.A(new_n2566), .Y(new_n3923));
  nand_5 g01575(.A(new_n3923), .B(pi799), .Y(new_n3924));
  nand_5 g01576(.A(new_n3924), .B(new_n3922), .Y(new_n3925));
  nand_5 g01577(.A(new_n3908), .B(new_n3906), .Y(new_n3926));
  xnor_4 g01578(.A(new_n3926), .B(new_n3907), .Y(new_n3927));
  xor_4  g01579(.A(new_n3924), .B(new_n3922), .Y(new_n3928));
  not_8  g01580(.A(new_n3928), .Y(new_n3929));
  or_6   g01581(.A(new_n3929), .B(new_n3927), .Y(new_n3930));
  nand_5 g01582(.A(new_n3930), .B(new_n3925), .Y(new_n3931));
  nand_5 g01583(.A(new_n3931), .B(new_n3921), .Y(new_n3932));
  not_8  g01584(.A(pi176), .Y(new_n3933));
  or_6   g01585(.A(new_n3931), .B(new_n3921), .Y(new_n3934));
  nand_5 g01586(.A(new_n3934), .B(new_n3933), .Y(new_n3935));
  nand_5 g01587(.A(new_n3935), .B(new_n3932), .Y(new_n3936));
  nand_5 g01588(.A(new_n3936), .B(new_n3919), .Y(new_n3937));
  not_8  g01589(.A(new_n3937), .Y(new_n3938));
  xor_4  g01590(.A(new_n3936), .B(new_n3918), .Y(new_n3939));
  nor_5  g01591(.A(new_n3939), .B(pi183), .Y(new_n3940));
  nor_5  g01592(.A(new_n3940), .B(new_n3938), .Y(new_n3941));
  xor_4  g01593(.A(new_n3941), .B(new_n3917), .Y(new_n3942));
  not_8  g01594(.A(new_n3942), .Y(new_n3943));
  not_8  g01595(.A(pi058), .Y(new_n3944));
  xor_4  g01596(.A(pi338), .B(new_n3944), .Y(new_n3945));
  not_8  g01597(.A(pi362), .Y(new_n3946));
  nand_5 g01598(.A(new_n3946), .B(pi305), .Y(new_n3947));
  not_8  g01599(.A(new_n3947), .Y(new_n3948));
  not_8  g01600(.A(pi305), .Y(new_n3949));
  xor_4  g01601(.A(pi362), .B(new_n3949), .Y(new_n3950));
  not_8  g01602(.A(new_n3950), .Y(new_n3951));
  not_8  g01603(.A(pi350), .Y(new_n3952));
  nand_5 g01604(.A(pi528), .B(new_n3952), .Y(new_n3953));
  not_8  g01605(.A(pi528), .Y(new_n3954));
  nand_5 g01606(.A(new_n3954), .B(pi350), .Y(new_n3955));
  nand_5 g01607(.A(new_n3955), .B(new_n2569), .Y(new_n3956));
  nand_5 g01608(.A(new_n3956), .B(new_n3953), .Y(new_n3957));
  nor_5  g01609(.A(new_n3957), .B(new_n3951), .Y(new_n3958));
  nor_5  g01610(.A(new_n3958), .B(new_n3948), .Y(new_n3959));
  xor_4  g01611(.A(new_n3959), .B(new_n3945), .Y(new_n3960));
  not_8  g01612(.A(new_n3960), .Y(new_n3961));
  not_8  g01613(.A(pi614), .Y(new_n3962));
  not_8  g01614(.A(pi271), .Y(new_n3963));
  nor_5  g01615(.A(pi656), .B(pi218), .Y(new_n3964));
  nand_5 g01616(.A(new_n3964), .B(new_n3963), .Y(new_n3965));
  xor_4  g01617(.A(new_n3965), .B(new_n3962), .Y(new_n3966));
  nand_5 g01618(.A(new_n3966), .B(new_n3961), .Y(new_n3967));
  xor_4  g01619(.A(new_n3957), .B(new_n3951), .Y(new_n3968));
  xor_4  g01620(.A(new_n3964), .B(pi271), .Y(new_n3969));
  and_6  g01621(.A(new_n3969), .B(new_n3968), .Y(new_n3970));
  nand_5 g01622(.A(new_n3955), .B(new_n3953), .Y(new_n3971));
  not_8  g01623(.A(new_n2569), .Y(new_n3972));
  nor_5  g01624(.A(new_n2571), .B(pi218), .Y(new_n3973));
  nor_5  g01625(.A(new_n3973), .B(new_n3972), .Y(new_n3974));
  nor_5  g01626(.A(new_n3974), .B(new_n3971), .Y(new_n3975));
  not_8  g01627(.A(pi218), .Y(new_n3976));
  nand_5 g01628(.A(new_n2571), .B(pi656), .Y(new_n3977));
  nor_5  g01629(.A(new_n3977), .B(new_n3976), .Y(new_n3978));
  not_8  g01630(.A(pi656), .Y(new_n3979));
  nand_5 g01631(.A(new_n3972), .B(new_n3979), .Y(new_n3980));
  nand_5 g01632(.A(new_n3980), .B(new_n3971), .Y(new_n3981));
  nor_5  g01633(.A(new_n3981), .B(new_n3978), .Y(new_n3982));
  nor_5  g01634(.A(new_n3982), .B(new_n3975), .Y(new_n3983));
  nor_5  g01635(.A(new_n3983), .B(new_n3964), .Y(new_n3984));
  xnor_4 g01636(.A(new_n3969), .B(new_n3968), .Y(new_n3985));
  nor_5  g01637(.A(new_n3985), .B(new_n3984), .Y(new_n3986));
  nor_5  g01638(.A(new_n3986), .B(new_n3970), .Y(new_n3987));
  xor_4  g01639(.A(new_n3966), .B(new_n3960), .Y(new_n3988));
  or_6   g01640(.A(new_n3988), .B(new_n3987), .Y(new_n3989));
  nand_5 g01641(.A(new_n3989), .B(new_n3967), .Y(new_n3990));
  not_8  g01642(.A(pi250), .Y(new_n3991));
  xor_4  g01643(.A(pi479), .B(new_n3991), .Y(new_n3992));
  not_8  g01644(.A(pi338), .Y(new_n3993));
  nand_5 g01645(.A(new_n3993), .B(pi058), .Y(new_n3994));
  not_8  g01646(.A(new_n3959), .Y(new_n3995));
  nand_5 g01647(.A(new_n3995), .B(new_n3945), .Y(new_n3996));
  nand_5 g01648(.A(new_n3996), .B(new_n3994), .Y(new_n3997));
  xnor_4 g01649(.A(new_n3997), .B(new_n3992), .Y(new_n3998));
  not_8  g01650(.A(pi602), .Y(new_n3999));
  nor_5  g01651(.A(new_n3965), .B(pi614), .Y(new_n4000));
  xor_4  g01652(.A(new_n4000), .B(new_n3999), .Y(new_n4001));
  xor_4  g01653(.A(new_n4001), .B(new_n3998), .Y(new_n4002));
  xor_4  g01654(.A(new_n4002), .B(new_n3990), .Y(new_n4003));
  nor_5  g01655(.A(new_n4003), .B(new_n3943), .Y(new_n4004));
  not_8  g01656(.A(pi183), .Y(new_n4005));
  xor_4  g01657(.A(new_n3939), .B(new_n4005), .Y(new_n4006));
  xor_4  g01658(.A(new_n3988), .B(new_n3987), .Y(new_n4007));
  not_8  g01659(.A(new_n4007), .Y(new_n4008));
  nor_5  g01660(.A(new_n4008), .B(new_n4006), .Y(new_n4009));
  and_6  g01661(.A(new_n3934), .B(new_n3932), .Y(new_n4010));
  xor_4  g01662(.A(new_n4010), .B(new_n3933), .Y(new_n4011));
  xor_4  g01663(.A(new_n3985), .B(new_n3984), .Y(new_n4012));
  nor_5  g01664(.A(new_n4012), .B(new_n4011), .Y(new_n4013));
  xor_4  g01665(.A(new_n4012), .B(new_n4011), .Y(new_n4014));
  not_8  g01666(.A(new_n4014), .Y(new_n4015));
  xor_4  g01667(.A(new_n3929), .B(new_n3927), .Y(new_n4016));
  xor_4  g01668(.A(new_n3971), .B(new_n3976), .Y(new_n4017));
  nand_5 g01669(.A(new_n2573), .B(new_n2567), .Y(new_n4018));
  nand_5 g01670(.A(new_n3977), .B(new_n2569), .Y(new_n4019));
  not_8  g01671(.A(new_n4019), .Y(new_n4020));
  xor_4  g01672(.A(new_n4020), .B(new_n4018), .Y(new_n4021));
  xor_4  g01673(.A(new_n4021), .B(new_n4016), .Y(new_n4022));
  xor_4  g01674(.A(new_n4022), .B(new_n4017), .Y(po0189));
  nand_5 g01675(.A(po0189), .B(new_n4016), .Y(new_n4024));
  not_8  g01676(.A(new_n4017), .Y(new_n4025));
  nand_5 g01677(.A(new_n4020), .B(new_n4018), .Y(new_n4026));
  nor_5  g01678(.A(new_n4026), .B(new_n4025), .Y(new_n4027));
  nor_5  g01679(.A(new_n4021), .B(new_n4016), .Y(new_n4028));
  or_6   g01680(.A(new_n2571), .B(pi656), .Y(new_n4029));
  nand_5 g01681(.A(new_n4029), .B(new_n4025), .Y(new_n4030));
  nor_5  g01682(.A(new_n4030), .B(new_n4028), .Y(new_n4031));
  nor_5  g01683(.A(new_n4031), .B(new_n4027), .Y(new_n4032));
  nand_5 g01684(.A(new_n4032), .B(new_n4024), .Y(new_n4033));
  nor_5  g01685(.A(new_n4033), .B(new_n4015), .Y(new_n4034));
  or_6   g01686(.A(new_n4034), .B(new_n4013), .Y(new_n4035));
  xor_4  g01687(.A(new_n4007), .B(new_n4006), .Y(new_n4036));
  nor_5  g01688(.A(new_n4036), .B(new_n4035), .Y(new_n4037));
  or_6   g01689(.A(new_n4037), .B(new_n4009), .Y(new_n4038));
  xor_4  g01690(.A(new_n4003), .B(new_n3942), .Y(new_n4039));
  nor_5  g01691(.A(new_n4039), .B(new_n4038), .Y(new_n4040));
  nor_5  g01692(.A(new_n4040), .B(new_n4004), .Y(new_n4041));
  nand_5 g01693(.A(new_n3895), .B(pi359), .Y(new_n4042));
  nand_5 g01694(.A(new_n3915), .B(new_n3896), .Y(new_n4043));
  nand_5 g01695(.A(new_n4043), .B(new_n4042), .Y(new_n4044));
  not_8  g01696(.A(pi351), .Y(new_n4045));
  nand_5 g01697(.A(pi588), .B(new_n4045), .Y(new_n4046));
  or_6   g01698(.A(pi588), .B(new_n4045), .Y(new_n4047));
  and_6  g01699(.A(new_n4047), .B(new_n4046), .Y(new_n4048));
  xor_4  g01700(.A(new_n4048), .B(new_n4044), .Y(new_n4049));
  not_8  g01701(.A(new_n4049), .Y(new_n4050));
  not_8  g01702(.A(new_n3916), .Y(new_n4051));
  nand_5 g01703(.A(new_n4051), .B(pi568), .Y(new_n4052));
  nand_5 g01704(.A(new_n3941), .B(new_n3917), .Y(new_n4053));
  nand_5 g01705(.A(new_n4053), .B(new_n4052), .Y(new_n4054));
  or_6   g01706(.A(new_n4054), .B(new_n4050), .Y(new_n4055));
  nand_5 g01707(.A(new_n4054), .B(new_n4050), .Y(new_n4056));
  nand_5 g01708(.A(new_n4056), .B(new_n4055), .Y(new_n4057));
  xor_4  g01709(.A(new_n4057), .B(pi433), .Y(new_n4058));
  not_8  g01710(.A(new_n4058), .Y(new_n4059));
  not_8  g01711(.A(pi394), .Y(new_n4060));
  nand_5 g01712(.A(pi479), .B(new_n3991), .Y(new_n4061));
  nand_5 g01713(.A(new_n3997), .B(new_n3992), .Y(new_n4062));
  nand_5 g01714(.A(new_n4062), .B(new_n4061), .Y(new_n4063));
  xor_4  g01715(.A(pi791), .B(pi613), .Y(new_n4064));
  xor_4  g01716(.A(new_n4064), .B(new_n4063), .Y(new_n4065));
  xor_4  g01717(.A(new_n4065), .B(new_n4060), .Y(new_n4066));
  nand_5 g01718(.A(new_n4000), .B(new_n3999), .Y(new_n4067));
  or_6   g01719(.A(new_n4001), .B(new_n3998), .Y(new_n4068));
  nand_5 g01720(.A(new_n4002), .B(new_n3990), .Y(new_n4069));
  nand_5 g01721(.A(new_n4069), .B(new_n4068), .Y(new_n4070));
  nand_5 g01722(.A(new_n4070), .B(new_n4067), .Y(new_n4071));
  xnor_4 g01723(.A(new_n4071), .B(new_n4066), .Y(new_n4072));
  xor_4  g01724(.A(new_n4072), .B(new_n4059), .Y(new_n4073));
  xor_4  g01725(.A(new_n4073), .B(new_n4041), .Y(po0008));
  not_8  g01726(.A(pi837), .Y(new_n4075));
  nor_5  g01727(.A(new_n4075), .B(new_n3954), .Y(new_n4076));
  xor_4  g01728(.A(pi837), .B(pi528), .Y(new_n4077));
  nand_5 g01729(.A(pi708), .B(pi219), .Y(new_n4078));
  not_8  g01730(.A(new_n4078), .Y(new_n4079));
  and_6  g01731(.A(new_n4079), .B(new_n4077), .Y(new_n4080));
  nor_5  g01732(.A(new_n4080), .B(new_n4076), .Y(new_n4081));
  xor_4  g01733(.A(pi760), .B(new_n3946), .Y(new_n4082));
  xor_4  g01734(.A(new_n4082), .B(new_n4081), .Y(new_n4083));
  not_8  g01735(.A(pi051), .Y(new_n4084));
  xor_4  g01736(.A(pi609), .B(new_n4084), .Y(new_n4085));
  not_8  g01737(.A(pi356), .Y(new_n4086));
  nand_5 g01738(.A(pi680), .B(new_n4086), .Y(new_n4087));
  not_8  g01739(.A(pi307), .Y(new_n4088));
  nand_5 g01740(.A(pi745), .B(new_n4088), .Y(new_n4089));
  not_8  g01741(.A(new_n4089), .Y(new_n4090));
  xor_4  g01742(.A(pi680), .B(new_n4086), .Y(new_n4091));
  nand_5 g01743(.A(new_n4091), .B(new_n4090), .Y(new_n4092));
  nand_5 g01744(.A(new_n4092), .B(new_n4087), .Y(new_n4093));
  xor_4  g01745(.A(new_n4093), .B(new_n4085), .Y(new_n4094));
  not_8  g01746(.A(new_n4094), .Y(new_n4095));
  xor_4  g01747(.A(new_n4091), .B(new_n4090), .Y(new_n4096));
  xor_4  g01748(.A(new_n4096), .B(new_n4077), .Y(new_n4097));
  nor_5  g01749(.A(pi708), .B(pi219), .Y(new_n4098));
  xor_4  g01750(.A(pi745), .B(new_n4088), .Y(new_n4099));
  nor_5  g01751(.A(new_n4099), .B(new_n4098), .Y(new_n4100));
  nor_5  g01752(.A(new_n4100), .B(new_n4079), .Y(new_n4101));
  not_8  g01753(.A(new_n4101), .Y(new_n4102));
  or_6   g01754(.A(new_n4102), .B(new_n4097), .Y(new_n4103));
  not_8  g01755(.A(new_n4096), .Y(new_n4104));
  nor_5  g01756(.A(new_n4104), .B(new_n4077), .Y(new_n4105));
  nor_5  g01757(.A(new_n4105), .B(new_n4080), .Y(new_n4106));
  nand_5 g01758(.A(new_n4106), .B(new_n4103), .Y(new_n4107));
  xor_4  g01759(.A(new_n4107), .B(new_n4095), .Y(new_n4108));
  xor_4  g01760(.A(new_n4108), .B(new_n4083), .Y(new_n4109));
  nand_5 g01761(.A(pi774), .B(pi245), .Y(new_n4110));
  not_8  g01762(.A(new_n4110), .Y(new_n4111));
  not_8  g01763(.A(pi017), .Y(new_n4112));
  xor_4  g01764(.A(pi176), .B(new_n4112), .Y(new_n4113));
  xor_4  g01765(.A(new_n4113), .B(new_n4111), .Y(new_n4114));
  xor_4  g01766(.A(pi774), .B(pi245), .Y(new_n4115));
  nand_5 g01767(.A(pi799), .B(pi622), .Y(new_n4116));
  xor_4  g01768(.A(pi799), .B(pi622), .Y(new_n4117));
  nor_5  g01769(.A(new_n4098), .B(new_n4079), .Y(new_n4118));
  xor_4  g01770(.A(new_n4118), .B(new_n4099), .Y(new_n4119));
  nand_5 g01771(.A(new_n4119), .B(new_n4117), .Y(new_n4120));
  nand_5 g01772(.A(new_n4120), .B(new_n4116), .Y(new_n4121));
  or_6   g01773(.A(new_n4121), .B(new_n4115), .Y(new_n4122));
  xor_4  g01774(.A(new_n4101), .B(new_n4097), .Y(new_n4123));
  xor_4  g01775(.A(new_n4121), .B(new_n4115), .Y(new_n4124));
  nand_5 g01776(.A(new_n4124), .B(new_n4123), .Y(new_n4125));
  nand_5 g01777(.A(new_n4125), .B(new_n4122), .Y(new_n4126));
  xor_4  g01778(.A(new_n4126), .B(new_n4114), .Y(new_n4127));
  not_8  g01779(.A(new_n4127), .Y(new_n4128));
  xor_4  g01780(.A(new_n4128), .B(new_n4109), .Y(po0009));
  not_8  g01781(.A(pi524), .Y(new_n4130));
  xor_4  g01782(.A(pi795), .B(new_n4130), .Y(new_n4131));
  nand_5 g01783(.A(new_n3723), .B(pi460), .Y(new_n4132));
  not_8  g01784(.A(pi460), .Y(new_n4133));
  xor_4  g01785(.A(pi495), .B(new_n4133), .Y(new_n4134));
  nand_5 g01786(.A(new_n3726), .B(pi215), .Y(new_n4135));
  not_8  g01787(.A(pi781), .Y(new_n4136));
  nand_5 g01788(.A(new_n4136), .B(pi758), .Y(new_n4137));
  not_8  g01789(.A(new_n4137), .Y(new_n4138));
  not_8  g01790(.A(pi215), .Y(new_n4139));
  xor_4  g01791(.A(pi422), .B(new_n4139), .Y(new_n4140));
  nand_5 g01792(.A(new_n4140), .B(new_n4138), .Y(new_n4141));
  nand_5 g01793(.A(new_n4141), .B(new_n4135), .Y(new_n4142));
  nand_5 g01794(.A(new_n4142), .B(new_n4134), .Y(new_n4143));
  nand_5 g01795(.A(new_n4143), .B(new_n4132), .Y(new_n4144));
  xor_4  g01796(.A(new_n4144), .B(new_n4131), .Y(new_n4145));
  not_8  g01797(.A(new_n4145), .Y(new_n4146));
  xor_4  g01798(.A(pi645), .B(new_n3811), .Y(new_n4147));
  not_8  g01799(.A(new_n4147), .Y(new_n4148));
  not_8  g01800(.A(pi825), .Y(new_n4149));
  nand_5 g01801(.A(new_n4149), .B(pi597), .Y(new_n4150));
  nand_5 g01802(.A(pi825), .B(new_n3828), .Y(new_n4151));
  not_8  g01803(.A(pi329), .Y(new_n4152));
  nand_5 g01804(.A(pi672), .B(new_n4152), .Y(new_n4153));
  nand_5 g01805(.A(new_n3863), .B(pi295), .Y(new_n4154));
  nand_5 g01806(.A(new_n3814), .B(pi329), .Y(new_n4155));
  nand_5 g01807(.A(new_n4155), .B(new_n4154), .Y(new_n4156));
  nand_5 g01808(.A(new_n4156), .B(new_n4153), .Y(new_n4157));
  nand_5 g01809(.A(new_n4157), .B(new_n4151), .Y(new_n4158));
  nand_5 g01810(.A(new_n4158), .B(new_n4150), .Y(new_n4159));
  xor_4  g01811(.A(new_n4159), .B(new_n4148), .Y(new_n4160));
  xor_4  g01812(.A(pi558), .B(new_n2948), .Y(new_n4161));
  nand_5 g01813(.A(new_n2960), .B(pi231), .Y(new_n4162));
  not_8  g01814(.A(new_n4162), .Y(new_n4163));
  xor_4  g01815(.A(pi277), .B(new_n2869), .Y(new_n4164));
  not_8  g01816(.A(new_n4164), .Y(new_n4165));
  nand_5 g01817(.A(new_n2875), .B(pi313), .Y(new_n4166));
  nand_5 g01818(.A(pi447), .B(new_n3785), .Y(new_n4167));
  nand_5 g01819(.A(new_n3815), .B(pi025), .Y(new_n4168));
  nand_5 g01820(.A(new_n4168), .B(new_n4167), .Y(new_n4169));
  nand_5 g01821(.A(new_n4169), .B(new_n4166), .Y(new_n4170));
  nor_5  g01822(.A(new_n4170), .B(new_n4165), .Y(new_n4171));
  nor_5  g01823(.A(new_n4171), .B(new_n4163), .Y(new_n4172));
  xor_4  g01824(.A(new_n4172), .B(new_n4161), .Y(new_n4173));
  and_6  g01825(.A(new_n4151), .B(new_n4150), .Y(new_n4174));
  xor_4  g01826(.A(new_n4174), .B(new_n4157), .Y(new_n4175));
  not_8  g01827(.A(new_n4175), .Y(new_n4176));
  xor_4  g01828(.A(new_n4170), .B(new_n4164), .Y(new_n4177));
  not_8  g01829(.A(new_n4177), .Y(new_n4178));
  nand_5 g01830(.A(new_n4178), .B(new_n4176), .Y(new_n4179));
  xor_4  g01831(.A(new_n4177), .B(new_n4175), .Y(new_n4180));
  nand_5 g01832(.A(new_n4155), .B(new_n4153), .Y(new_n4181));
  not_8  g01833(.A(new_n4181), .Y(new_n4182));
  xor_4  g01834(.A(new_n4182), .B(new_n4154), .Y(new_n4183));
  not_8  g01835(.A(pi295), .Y(new_n4184));
  nand_5 g01836(.A(pi385), .B(new_n4184), .Y(new_n4185));
  nand_5 g01837(.A(new_n4185), .B(new_n4154), .Y(new_n4186));
  not_8  g01838(.A(new_n4186), .Y(new_n4187));
  xor_4  g01839(.A(pi832), .B(new_n2747), .Y(new_n4188));
  nor_5  g01840(.A(new_n4188), .B(new_n4187), .Y(new_n4189));
  or_6   g01841(.A(new_n4189), .B(new_n4183), .Y(new_n4190));
  nand_5 g01842(.A(new_n4189), .B(new_n4183), .Y(new_n4191));
  nand_5 g01843(.A(new_n4167), .B(new_n4166), .Y(new_n4192));
  xnor_4 g01844(.A(new_n4192), .B(new_n4168), .Y(new_n4193));
  not_8  g01845(.A(new_n4193), .Y(new_n4194));
  nand_5 g01846(.A(new_n4194), .B(new_n4191), .Y(new_n4195));
  nand_5 g01847(.A(new_n4195), .B(new_n4190), .Y(new_n4196));
  nand_5 g01848(.A(new_n4196), .B(new_n4180), .Y(new_n4197));
  nand_5 g01849(.A(new_n4197), .B(new_n4179), .Y(new_n4198));
  xor_4  g01850(.A(new_n4198), .B(new_n4173), .Y(new_n4199));
  xor_4  g01851(.A(new_n4199), .B(new_n4160), .Y(new_n4200));
  nand_5 g01852(.A(new_n4200), .B(new_n4146), .Y(new_n4201));
  xor_4  g01853(.A(new_n4200), .B(new_n4146), .Y(new_n4202));
  xor_4  g01854(.A(new_n4142), .B(new_n4134), .Y(new_n4203));
  not_8  g01855(.A(pi758), .Y(new_n4204));
  xor_4  g01856(.A(pi781), .B(new_n4204), .Y(new_n4205));
  not_8  g01857(.A(new_n4205), .Y(new_n4206));
  xor_4  g01858(.A(new_n4188), .B(new_n4187), .Y(new_n4207));
  nand_5 g01859(.A(new_n4207), .B(new_n4206), .Y(new_n4208));
  xor_4  g01860(.A(new_n4140), .B(new_n4137), .Y(new_n4209));
  not_8  g01861(.A(new_n4209), .Y(new_n4210));
  nand_5 g01862(.A(new_n4210), .B(new_n4208), .Y(new_n4211));
  xor_4  g01863(.A(new_n4210), .B(new_n4208), .Y(new_n4212));
  nand_5 g01864(.A(new_n4190), .B(new_n4191), .Y(new_n4213));
  xor_4  g01865(.A(new_n4213), .B(new_n4194), .Y(new_n4214));
  not_8  g01866(.A(new_n4214), .Y(new_n4215));
  nand_5 g01867(.A(new_n4215), .B(new_n4212), .Y(new_n4216));
  nand_5 g01868(.A(new_n4216), .B(new_n4211), .Y(new_n4217));
  or_6   g01869(.A(new_n4217), .B(new_n4203), .Y(new_n4218));
  xor_4  g01870(.A(new_n4217), .B(new_n4203), .Y(new_n4219));
  xor_4  g01871(.A(new_n4196), .B(new_n4180), .Y(new_n4220));
  not_8  g01872(.A(new_n4220), .Y(new_n4221));
  nand_5 g01873(.A(new_n4221), .B(new_n4219), .Y(new_n4222));
  nand_5 g01874(.A(new_n4222), .B(new_n4218), .Y(new_n4223));
  nand_5 g01875(.A(new_n4223), .B(new_n4202), .Y(new_n4224));
  nand_5 g01876(.A(new_n4224), .B(new_n4201), .Y(new_n4225));
  xor_4  g01877(.A(pi604), .B(new_n3718), .Y(new_n4226));
  not_8  g01878(.A(pi795), .Y(new_n4227));
  nand_5 g01879(.A(new_n4227), .B(pi524), .Y(new_n4228));
  nand_5 g01880(.A(new_n4144), .B(new_n4131), .Y(new_n4229));
  nand_5 g01881(.A(new_n4229), .B(new_n4228), .Y(new_n4230));
  xor_4  g01882(.A(new_n4230), .B(new_n4226), .Y(new_n4231));
  not_8  g01883(.A(new_n4231), .Y(new_n4232));
  xor_4  g01884(.A(pi590), .B(new_n2864), .Y(new_n4233));
  nand_5 g01885(.A(pi558), .B(new_n2948), .Y(new_n4234));
  not_8  g01886(.A(new_n4172), .Y(new_n4235));
  nand_5 g01887(.A(new_n4235), .B(new_n4161), .Y(new_n4236));
  nand_5 g01888(.A(new_n4236), .B(new_n4234), .Y(new_n4237));
  xor_4  g01889(.A(new_n4237), .B(new_n4233), .Y(new_n4238));
  xor_4  g01890(.A(pi432), .B(new_n3846), .Y(new_n4239));
  nand_5 g01891(.A(pi645), .B(new_n3811), .Y(new_n4240));
  not_8  g01892(.A(new_n4240), .Y(new_n4241));
  nor_5  g01893(.A(new_n4159), .B(new_n4148), .Y(new_n4242));
  nor_5  g01894(.A(new_n4242), .B(new_n4241), .Y(new_n4243));
  xor_4  g01895(.A(new_n4243), .B(new_n4239), .Y(new_n4244));
  not_8  g01896(.A(new_n4173), .Y(new_n4245));
  nor_5  g01897(.A(new_n4198), .B(new_n4245), .Y(new_n4246));
  nor_5  g01898(.A(new_n4199), .B(new_n4160), .Y(new_n4247));
  or_6   g01899(.A(new_n4247), .B(new_n4246), .Y(new_n4248));
  xnor_4 g01900(.A(new_n4248), .B(new_n4244), .Y(new_n4249));
  xor_4  g01901(.A(new_n4249), .B(new_n4238), .Y(new_n4250));
  xor_4  g01902(.A(new_n4250), .B(new_n4232), .Y(new_n4251));
  xor_4  g01903(.A(new_n4251), .B(new_n4225), .Y(po0010));
  nand_5 g01904(.A(pi565), .B(new_n2607), .Y(new_n4253));
  not_8  g01905(.A(new_n4253), .Y(new_n4254));
  xor_4  g01906(.A(pi565), .B(new_n2607), .Y(new_n4255));
  not_8  g01907(.A(new_n4255), .Y(new_n4256));
  not_8  g01908(.A(pi059), .Y(new_n4257));
  nand_5 g01909(.A(pi784), .B(new_n4257), .Y(new_n4258));
  not_8  g01910(.A(new_n4258), .Y(new_n4259));
  xor_4  g01911(.A(pi784), .B(new_n4257), .Y(new_n4260));
  not_8  g01912(.A(new_n4260), .Y(new_n4261));
  not_8  g01913(.A(pi734), .Y(new_n4262));
  nor_5  g01914(.A(pi771), .B(new_n4262), .Y(new_n4263));
  xor_4  g01915(.A(pi771), .B(new_n4262), .Y(new_n4264));
  not_8  g01916(.A(new_n4264), .Y(new_n4265));
  not_8  g01917(.A(pi395), .Y(new_n4266));
  nand_5 g01918(.A(new_n4266), .B(pi304), .Y(new_n4267));
  xor_4  g01919(.A(new_n4266), .B(pi304), .Y(new_n4268));
  nand_5 g01920(.A(new_n4047), .B(new_n4044), .Y(new_n4269));
  nand_5 g01921(.A(new_n4269), .B(new_n4046), .Y(new_n4270));
  nand_5 g01922(.A(new_n4270), .B(new_n4268), .Y(new_n4271));
  nand_5 g01923(.A(new_n4271), .B(new_n4267), .Y(new_n4272));
  nor_5  g01924(.A(new_n4272), .B(new_n4265), .Y(new_n4273));
  nor_5  g01925(.A(new_n4273), .B(new_n4263), .Y(new_n4274));
  nor_5  g01926(.A(new_n4274), .B(new_n4261), .Y(new_n4275));
  nor_5  g01927(.A(new_n4275), .B(new_n4259), .Y(new_n4276));
  nor_5  g01928(.A(new_n4276), .B(new_n4256), .Y(new_n4277));
  nor_5  g01929(.A(new_n4277), .B(new_n4254), .Y(new_n4278));
  not_8  g01930(.A(new_n4278), .Y(new_n4279));
  not_8  g01931(.A(pi503), .Y(new_n4280));
  not_8  g01932(.A(pi761), .Y(new_n4281));
  not_8  g01933(.A(pi741), .Y(new_n4282));
  or_6   g01934(.A(new_n3927), .B(new_n4282), .Y(new_n4283));
  nand_5 g01935(.A(new_n3927), .B(new_n4282), .Y(new_n4284));
  nand_5 g01936(.A(new_n4284), .B(pi702), .Y(new_n4285));
  nand_5 g01937(.A(new_n4285), .B(new_n4283), .Y(new_n4286));
  or_6   g01938(.A(new_n4286), .B(new_n3921), .Y(new_n4287));
  not_8  g01939(.A(pi221), .Y(new_n4288));
  nand_5 g01940(.A(new_n4286), .B(new_n3921), .Y(new_n4289));
  nand_5 g01941(.A(new_n4289), .B(new_n4288), .Y(new_n4290));
  nand_5 g01942(.A(new_n4290), .B(new_n4287), .Y(new_n4291));
  nor_5  g01943(.A(new_n4291), .B(new_n4281), .Y(new_n4292));
  xor_4  g01944(.A(new_n4291), .B(pi761), .Y(new_n4293));
  nor_5  g01945(.A(new_n4293), .B(new_n3918), .Y(new_n4294));
  or_6   g01946(.A(new_n4294), .B(new_n4292), .Y(new_n4295));
  nand_5 g01947(.A(new_n4295), .B(new_n3916), .Y(new_n4296));
  or_6   g01948(.A(new_n4295), .B(new_n3916), .Y(new_n4297));
  nand_5 g01949(.A(new_n4297), .B(pi003), .Y(new_n4298));
  nand_5 g01950(.A(new_n4298), .B(new_n4296), .Y(new_n4299));
  nand_5 g01951(.A(new_n4299), .B(pi400), .Y(new_n4300));
  xor_4  g01952(.A(new_n4299), .B(pi400), .Y(new_n4301));
  nand_5 g01953(.A(new_n4301), .B(new_n4049), .Y(new_n4302));
  nand_5 g01954(.A(new_n4302), .B(new_n4300), .Y(new_n4303));
  xor_4  g01955(.A(new_n4270), .B(new_n4268), .Y(new_n4304));
  or_6   g01956(.A(new_n4304), .B(new_n4303), .Y(new_n4305));
  not_8  g01957(.A(pi780), .Y(new_n4306));
  xor_4  g01958(.A(new_n4304), .B(new_n4303), .Y(new_n4307));
  nand_5 g01959(.A(new_n4307), .B(new_n4306), .Y(new_n4308));
  nand_5 g01960(.A(new_n4308), .B(new_n4305), .Y(new_n4309));
  or_6   g01961(.A(new_n4309), .B(new_n4280), .Y(new_n4310));
  xor_4  g01962(.A(new_n4309), .B(new_n4280), .Y(new_n4311));
  xor_4  g01963(.A(new_n4272), .B(new_n4264), .Y(new_n4312));
  nand_5 g01964(.A(new_n4312), .B(new_n4311), .Y(new_n4313));
  nand_5 g01965(.A(new_n4313), .B(new_n4310), .Y(new_n4314));
  nand_5 g01966(.A(new_n4314), .B(pi748), .Y(new_n4315));
  xor_4  g01967(.A(new_n4314), .B(pi748), .Y(new_n4316));
  xor_4  g01968(.A(new_n4274), .B(new_n4260), .Y(new_n4317));
  nand_5 g01969(.A(new_n4317), .B(new_n4316), .Y(new_n4318));
  nand_5 g01970(.A(new_n4318), .B(new_n4315), .Y(new_n4319));
  xor_4  g01971(.A(new_n4276), .B(new_n4255), .Y(new_n4320));
  nand_5 g01972(.A(new_n4320), .B(new_n4319), .Y(new_n4321));
  xor_4  g01973(.A(new_n4320), .B(new_n4319), .Y(new_n4322));
  nand_5 g01974(.A(new_n4322), .B(pi542), .Y(new_n4323));
  nand_5 g01975(.A(new_n4323), .B(new_n4321), .Y(new_n4324));
  nand_5 g01976(.A(new_n4324), .B(new_n4279), .Y(new_n4325));
  xor_4  g01977(.A(new_n4324), .B(new_n4279), .Y(new_n4326));
  not_8  g01978(.A(pi542), .Y(new_n4327));
  xor_4  g01979(.A(new_n4322), .B(new_n4327), .Y(new_n4328));
  not_8  g01980(.A(pi679), .Y(new_n4329));
  nand_5 g01981(.A(new_n4329), .B(pi663), .Y(new_n4330));
  not_8  g01982(.A(new_n4330), .Y(new_n4331));
  nor_5  g01983(.A(new_n4329), .B(pi663), .Y(new_n4332));
  nor_5  g01984(.A(new_n4332), .B(new_n4331), .Y(new_n4333));
  not_8  g01985(.A(new_n4333), .Y(new_n4334));
  not_8  g01986(.A(pi835), .Y(new_n4335));
  nand_5 g01987(.A(new_n4335), .B(pi291), .Y(new_n4336));
  nand_5 g01988(.A(new_n2939), .B(pi082), .Y(new_n4337));
  xor_4  g01989(.A(pi380), .B(new_n2813), .Y(new_n4338));
  nand_5 g01990(.A(new_n2943), .B(pi306), .Y(new_n4339));
  xor_4  g01991(.A(pi346), .B(new_n2671), .Y(new_n4340));
  not_8  g01992(.A(pi636), .Y(new_n4341));
  nand_5 g01993(.A(new_n4341), .B(pi213), .Y(new_n4342));
  xor_4  g01994(.A(pi636), .B(new_n2674), .Y(new_n4343));
  nand_5 g01995(.A(pi476), .B(new_n2966), .Y(new_n4344));
  xor_4  g01996(.A(pi476), .B(new_n2966), .Y(new_n4345));
  nand_5 g01997(.A(new_n2949), .B(pi211), .Y(new_n4346));
  not_8  g01998(.A(pi504), .Y(new_n4347));
  nand_5 g01999(.A(pi703), .B(new_n4347), .Y(new_n4348));
  xor_4  g02000(.A(pi703), .B(new_n4347), .Y(new_n4349));
  nand_5 g02001(.A(pi763), .B(new_n3020), .Y(new_n4350));
  nand_5 g02002(.A(pi449), .B(new_n2956), .Y(new_n4351));
  nand_5 g02003(.A(new_n4351), .B(new_n4350), .Y(new_n4352));
  not_8  g02004(.A(new_n4352), .Y(new_n4353));
  nor_5  g02005(.A(pi449), .B(new_n2956), .Y(new_n4354));
  nor_5  g02006(.A(new_n4354), .B(new_n4353), .Y(new_n4355));
  nand_5 g02007(.A(new_n4355), .B(new_n4349), .Y(new_n4356));
  nand_5 g02008(.A(new_n4356), .B(new_n4348), .Y(new_n4357));
  xor_4  g02009(.A(pi766), .B(pi211), .Y(new_n4358));
  not_8  g02010(.A(new_n4358), .Y(new_n4359));
  nand_5 g02011(.A(new_n4359), .B(new_n4357), .Y(new_n4360));
  nand_5 g02012(.A(new_n4360), .B(new_n4346), .Y(new_n4361));
  nand_5 g02013(.A(new_n4361), .B(new_n4345), .Y(new_n4362));
  nand_5 g02014(.A(new_n4362), .B(new_n4344), .Y(new_n4363));
  nand_5 g02015(.A(new_n4363), .B(new_n4343), .Y(new_n4364));
  nand_5 g02016(.A(new_n4364), .B(new_n4342), .Y(new_n4365));
  nand_5 g02017(.A(new_n4365), .B(new_n4340), .Y(new_n4366));
  nand_5 g02018(.A(new_n4366), .B(new_n4339), .Y(new_n4367));
  nand_5 g02019(.A(new_n4367), .B(new_n4338), .Y(new_n4368));
  nand_5 g02020(.A(new_n4368), .B(new_n4337), .Y(new_n4369));
  nand_5 g02021(.A(pi835), .B(new_n2838), .Y(new_n4370));
  nand_5 g02022(.A(new_n4370), .B(new_n4369), .Y(new_n4371));
  nand_5 g02023(.A(new_n4371), .B(new_n4336), .Y(new_n4372));
  xor_4  g02024(.A(new_n4372), .B(new_n4334), .Y(new_n4373));
  not_8  g02025(.A(pi368), .Y(new_n4374));
  nand_5 g02026(.A(new_n4370), .B(new_n4336), .Y(new_n4375));
  xnor_4 g02027(.A(new_n4375), .B(new_n4369), .Y(new_n4376));
  nand_5 g02028(.A(new_n4376), .B(new_n4374), .Y(new_n4377));
  or_6   g02029(.A(new_n4376), .B(new_n4374), .Y(new_n4378));
  xnor_4 g02030(.A(new_n4367), .B(new_n4338), .Y(new_n4379));
  or_6   g02031(.A(new_n4379), .B(pi505), .Y(new_n4380));
  xor_4  g02032(.A(new_n4379), .B(pi505), .Y(new_n4381));
  not_8  g02033(.A(pi473), .Y(new_n4382));
  xor_4  g02034(.A(new_n4365), .B(new_n4340), .Y(new_n4383));
  or_6   g02035(.A(new_n4383), .B(new_n4382), .Y(new_n4384));
  not_8  g02036(.A(new_n4384), .Y(new_n4385));
  xnor_4 g02037(.A(new_n4363), .B(new_n4343), .Y(new_n4386));
  nor_5  g02038(.A(new_n4386), .B(pi248), .Y(new_n4387));
  xor_4  g02039(.A(new_n4386), .B(pi248), .Y(new_n4388));
  not_8  g02040(.A(new_n4388), .Y(new_n4389));
  xnor_4 g02041(.A(new_n4361), .B(new_n4345), .Y(new_n4390));
  nand_5 g02042(.A(new_n4390), .B(pi125), .Y(new_n4391));
  xor_4  g02043(.A(new_n4390), .B(pi125), .Y(new_n4392));
  xor_4  g02044(.A(new_n4358), .B(new_n4357), .Y(new_n4393));
  nand_5 g02045(.A(new_n4393), .B(pi618), .Y(new_n4394));
  not_8  g02046(.A(pi618), .Y(new_n4395));
  not_8  g02047(.A(new_n4393), .Y(new_n4396));
  nand_5 g02048(.A(new_n4396), .B(new_n4395), .Y(new_n4397));
  xnor_4 g02049(.A(new_n4355), .B(new_n4349), .Y(new_n4398));
  nor_5  g02050(.A(new_n4398), .B(pi192), .Y(new_n4399));
  xor_4  g02051(.A(new_n4398), .B(pi192), .Y(new_n4400));
  xor_4  g02052(.A(pi449), .B(new_n2956), .Y(new_n4401));
  nor_5  g02053(.A(pi763), .B(new_n3020), .Y(new_n4402));
  not_8  g02054(.A(new_n4402), .Y(new_n4403));
  nand_5 g02055(.A(new_n4403), .B(pi049), .Y(new_n4404));
  not_8  g02056(.A(pi049), .Y(new_n4405));
  nand_5 g02057(.A(new_n4350), .B(new_n4405), .Y(new_n4406));
  nand_5 g02058(.A(new_n4406), .B(new_n4404), .Y(new_n4407));
  xor_4  g02059(.A(new_n4407), .B(new_n4401), .Y(new_n4408));
  nand_5 g02060(.A(new_n4408), .B(pi813), .Y(new_n4409));
  not_8  g02061(.A(new_n4409), .Y(new_n4410));
  nand_5 g02062(.A(new_n4403), .B(new_n4350), .Y(new_n4411));
  nand_5 g02063(.A(new_n4411), .B(pi049), .Y(new_n4412));
  nor_5  g02064(.A(new_n4412), .B(new_n4408), .Y(new_n4413));
  nor_5  g02065(.A(new_n4413), .B(new_n4410), .Y(new_n4414));
  nand_5 g02066(.A(new_n4414), .B(new_n4400), .Y(new_n4415));
  not_8  g02067(.A(new_n4415), .Y(new_n4416));
  nor_5  g02068(.A(new_n4416), .B(new_n4399), .Y(new_n4417));
  nand_5 g02069(.A(new_n4417), .B(new_n4397), .Y(new_n4418));
  nand_5 g02070(.A(new_n4418), .B(new_n4394), .Y(new_n4419));
  nand_5 g02071(.A(new_n4419), .B(new_n4392), .Y(new_n4420));
  nand_5 g02072(.A(new_n4420), .B(new_n4391), .Y(new_n4421));
  nor_5  g02073(.A(new_n4421), .B(new_n4389), .Y(new_n4422));
  or_6   g02074(.A(new_n4422), .B(new_n4387), .Y(new_n4423));
  xor_4  g02075(.A(new_n4383), .B(pi473), .Y(new_n4424));
  nor_5  g02076(.A(new_n4424), .B(new_n4423), .Y(new_n4425));
  nor_5  g02077(.A(new_n4425), .B(new_n4385), .Y(new_n4426));
  nand_5 g02078(.A(new_n4426), .B(new_n4381), .Y(new_n4427));
  nand_5 g02079(.A(new_n4427), .B(new_n4380), .Y(new_n4428));
  nand_5 g02080(.A(new_n4428), .B(new_n4378), .Y(new_n4429));
  nand_5 g02081(.A(new_n4429), .B(new_n4377), .Y(new_n4430));
  xor_4  g02082(.A(new_n4430), .B(pi716), .Y(new_n4431));
  xor_4  g02083(.A(new_n4431), .B(new_n4373), .Y(new_n4432));
  not_8  g02084(.A(new_n4432), .Y(new_n4433));
  nor_5  g02085(.A(new_n4433), .B(new_n4328), .Y(new_n4434));
  xor_4  g02086(.A(new_n4432), .B(new_n4328), .Y(new_n4435));
  not_8  g02087(.A(new_n4317), .Y(new_n4436));
  xor_4  g02088(.A(new_n4436), .B(new_n4316), .Y(new_n4437));
  nand_5 g02089(.A(new_n4377), .B(new_n4378), .Y(new_n4438));
  xor_4  g02090(.A(new_n4438), .B(new_n4428), .Y(new_n4439));
  nand_5 g02091(.A(new_n4439), .B(new_n4437), .Y(new_n4440));
  not_8  g02092(.A(new_n4312), .Y(new_n4441));
  xor_4  g02093(.A(new_n4441), .B(new_n4311), .Y(new_n4442));
  xor_4  g02094(.A(new_n4426), .B(new_n4381), .Y(new_n4443));
  not_8  g02095(.A(new_n4443), .Y(new_n4444));
  and_6  g02096(.A(new_n4444), .B(new_n4442), .Y(new_n4445));
  xor_4  g02097(.A(new_n4443), .B(new_n4442), .Y(new_n4446));
  xor_4  g02098(.A(new_n4307), .B(pi780), .Y(new_n4447));
  xor_4  g02099(.A(new_n4424), .B(new_n4423), .Y(new_n4448));
  not_8  g02100(.A(new_n4448), .Y(new_n4449));
  nand_5 g02101(.A(new_n4449), .B(new_n4447), .Y(new_n4450));
  xor_4  g02102(.A(new_n4293), .B(new_n3919), .Y(new_n4451));
  nand_5 g02103(.A(new_n4394), .B(new_n4397), .Y(new_n4452));
  xor_4  g02104(.A(new_n4452), .B(new_n4417), .Y(new_n4453));
  not_8  g02105(.A(new_n4453), .Y(new_n4454));
  nand_5 g02106(.A(new_n4454), .B(new_n4451), .Y(new_n4455));
  xor_4  g02107(.A(new_n4453), .B(new_n4451), .Y(new_n4456));
  nand_5 g02108(.A(new_n4289), .B(new_n4287), .Y(new_n4457));
  xor_4  g02109(.A(new_n4457), .B(pi221), .Y(new_n4458));
  xor_4  g02110(.A(new_n4414), .B(new_n4400), .Y(new_n4459));
  not_8  g02111(.A(new_n4459), .Y(new_n4460));
  nor_5  g02112(.A(new_n4460), .B(new_n4458), .Y(new_n4461));
  xor_4  g02113(.A(new_n4459), .B(new_n4458), .Y(new_n4462));
  xor_4  g02114(.A(new_n4408), .B(pi813), .Y(new_n4463));
  nand_5 g02115(.A(new_n4284), .B(new_n4283), .Y(new_n4464));
  xor_4  g02116(.A(new_n4411), .B(pi049), .Y(new_n4465));
  nand_5 g02117(.A(new_n2566), .B(pi702), .Y(new_n4466));
  nor_5  g02118(.A(new_n4466), .B(new_n4465), .Y(new_n4467));
  not_8  g02119(.A(new_n4465), .Y(new_n4468));
  nand_5 g02120(.A(new_n3923), .B(new_n2558), .Y(new_n4469));
  nor_5  g02121(.A(new_n4469), .B(new_n4468), .Y(new_n4470));
  or_6   g02122(.A(new_n4470), .B(new_n4467), .Y(new_n4471));
  xnor_4 g02123(.A(new_n4471), .B(new_n4464), .Y(new_n4472));
  nor_5  g02124(.A(new_n4472), .B(new_n4463), .Y(new_n4473));
  nand_5 g02125(.A(new_n4467), .B(new_n4464), .Y(new_n4474));
  nor_5  g02126(.A(new_n4471), .B(new_n4464), .Y(new_n4475));
  nand_5 g02127(.A(new_n4475), .B(new_n2558), .Y(new_n4476));
  nand_5 g02128(.A(new_n4476), .B(new_n4474), .Y(new_n4477));
  nor_5  g02129(.A(new_n4477), .B(new_n4473), .Y(new_n4478));
  nor_5  g02130(.A(new_n4478), .B(new_n4462), .Y(new_n4479));
  or_6   g02131(.A(new_n4479), .B(new_n4461), .Y(new_n4480));
  or_6   g02132(.A(new_n4480), .B(new_n4456), .Y(new_n4481));
  nand_5 g02133(.A(new_n4481), .B(new_n4455), .Y(new_n4482));
  nand_5 g02134(.A(new_n4297), .B(new_n4296), .Y(new_n4483));
  xor_4  g02135(.A(new_n4483), .B(pi003), .Y(new_n4484));
  nand_5 g02136(.A(new_n4484), .B(new_n4482), .Y(new_n4485));
  xor_4  g02137(.A(new_n4484), .B(new_n4482), .Y(new_n4486));
  xor_4  g02138(.A(new_n4419), .B(new_n4392), .Y(new_n4487));
  nand_5 g02139(.A(new_n4487), .B(new_n4486), .Y(new_n4488));
  nand_5 g02140(.A(new_n4488), .B(new_n4485), .Y(new_n4489));
  xor_4  g02141(.A(new_n4421), .B(new_n4388), .Y(new_n4490));
  nand_5 g02142(.A(new_n4490), .B(new_n4489), .Y(new_n4491));
  xor_4  g02143(.A(new_n4490), .B(new_n4489), .Y(new_n4492));
  not_8  g02144(.A(new_n4492), .Y(new_n4493));
  xor_4  g02145(.A(new_n4301), .B(new_n4049), .Y(new_n4494));
  or_6   g02146(.A(new_n4494), .B(new_n4493), .Y(new_n4495));
  nand_5 g02147(.A(new_n4495), .B(new_n4491), .Y(new_n4496));
  xor_4  g02148(.A(new_n4448), .B(new_n4447), .Y(new_n4497));
  or_6   g02149(.A(new_n4497), .B(new_n4496), .Y(new_n4498));
  nand_5 g02150(.A(new_n4498), .B(new_n4450), .Y(new_n4499));
  nor_5  g02151(.A(new_n4499), .B(new_n4446), .Y(new_n4500));
  nor_5  g02152(.A(new_n4500), .B(new_n4445), .Y(new_n4501));
  not_8  g02153(.A(new_n4439), .Y(new_n4502));
  xor_4  g02154(.A(new_n4502), .B(new_n4437), .Y(new_n4503));
  or_6   g02155(.A(new_n4503), .B(new_n4501), .Y(new_n4504));
  nand_5 g02156(.A(new_n4504), .B(new_n4440), .Y(new_n4505));
  nor_5  g02157(.A(new_n4505), .B(new_n4435), .Y(new_n4506));
  or_6   g02158(.A(new_n4506), .B(new_n4434), .Y(new_n4507));
  nor_5  g02159(.A(new_n4507), .B(new_n4326), .Y(new_n4508));
  nor_5  g02160(.A(new_n4372), .B(new_n4334), .Y(new_n4509));
  nor_5  g02161(.A(new_n4509), .B(new_n4331), .Y(new_n4510));
  not_8  g02162(.A(pi716), .Y(new_n4511));
  nor_5  g02163(.A(new_n4430), .B(new_n4511), .Y(new_n4512));
  nand_5 g02164(.A(new_n4372), .B(new_n4332), .Y(new_n4513));
  nor_5  g02165(.A(new_n4513), .B(new_n4512), .Y(new_n4514));
  nand_5 g02166(.A(new_n4430), .B(new_n4511), .Y(new_n4515));
  not_8  g02167(.A(new_n4510), .Y(new_n4516));
  or_6   g02168(.A(new_n4516), .B(new_n4515), .Y(new_n4517));
  nor_5  g02169(.A(new_n4372), .B(new_n4330), .Y(new_n4518));
  nand_5 g02170(.A(new_n4518), .B(new_n4515), .Y(new_n4519));
  nand_5 g02171(.A(new_n4519), .B(new_n4517), .Y(new_n4520));
  nor_5  g02172(.A(new_n4520), .B(new_n4514), .Y(new_n4521));
  nand_5 g02173(.A(new_n4521), .B(new_n4510), .Y(new_n4522));
  not_8  g02174(.A(new_n4522), .Y(new_n4523));
  nand_5 g02175(.A(new_n4523), .B(new_n4508), .Y(new_n4524));
  xor_4  g02176(.A(new_n4507), .B(new_n4326), .Y(new_n4525));
  nand_5 g02177(.A(new_n4516), .B(new_n4512), .Y(new_n4526));
  nand_5 g02178(.A(new_n4526), .B(new_n4521), .Y(new_n4527));
  nand_5 g02179(.A(new_n4527), .B(new_n4525), .Y(new_n4528));
  nor_5  g02180(.A(new_n4523), .B(new_n4508), .Y(new_n4529));
  nand_5 g02181(.A(new_n4529), .B(new_n4528), .Y(new_n4530));
  nand_5 g02182(.A(new_n4530), .B(new_n4524), .Y(new_n4531));
  xor_4  g02183(.A(new_n4531), .B(new_n4325), .Y(po0011));
  xor_4  g02184(.A(pi522), .B(new_n3542), .Y(new_n4533));
  not_8  g02185(.A(pi660), .Y(new_n4534));
  nand_5 g02186(.A(new_n4534), .B(pi421), .Y(new_n4535));
  xor_4  g02187(.A(pi660), .B(new_n3545), .Y(new_n4536));
  not_8  g02188(.A(pi178), .Y(new_n4537));
  nand_5 g02189(.A(pi626), .B(new_n4537), .Y(new_n4538));
  xor_4  g02190(.A(pi626), .B(new_n4537), .Y(new_n4539));
  not_8  g02191(.A(pi168), .Y(new_n4540));
  nand_5 g02192(.A(new_n4540), .B(pi045), .Y(new_n4541));
  xor_4  g02193(.A(pi168), .B(new_n3554), .Y(new_n4542));
  not_8  g02194(.A(pi710), .Y(new_n4543));
  nand_5 g02195(.A(new_n4543), .B(pi520), .Y(new_n4544));
  not_8  g02196(.A(new_n4544), .Y(new_n4545));
  nand_5 g02197(.A(new_n4545), .B(new_n4542), .Y(new_n4546));
  nand_5 g02198(.A(new_n4546), .B(new_n4541), .Y(new_n4547));
  nand_5 g02199(.A(new_n4547), .B(new_n4539), .Y(new_n4548));
  nand_5 g02200(.A(new_n4548), .B(new_n4538), .Y(new_n4549));
  nand_5 g02201(.A(new_n4549), .B(new_n4536), .Y(new_n4550));
  nand_5 g02202(.A(new_n4550), .B(new_n4535), .Y(new_n4551));
  xor_4  g02203(.A(new_n4551), .B(new_n4533), .Y(new_n4552));
  not_8  g02204(.A(pi226), .Y(new_n4553));
  xor_4  g02205(.A(pi750), .B(new_n4553), .Y(new_n4554));
  not_8  g02206(.A(pi240), .Y(new_n4555));
  nand_5 g02207(.A(pi673), .B(new_n4555), .Y(new_n4556));
  xor_4  g02208(.A(pi673), .B(new_n4555), .Y(new_n4557));
  not_8  g02209(.A(pi002), .Y(new_n4558));
  nand_5 g02210(.A(pi311), .B(new_n4558), .Y(new_n4559));
  not_8  g02211(.A(new_n4559), .Y(new_n4560));
  xor_4  g02212(.A(pi311), .B(new_n4558), .Y(new_n4561));
  not_8  g02213(.A(new_n4561), .Y(new_n4562));
  not_8  g02214(.A(pi378), .Y(new_n4563));
  or_6   g02215(.A(pi467), .B(new_n4563), .Y(new_n4564));
  nand_5 g02216(.A(pi467), .B(new_n4563), .Y(new_n4565));
  not_8  g02217(.A(pi426), .Y(new_n4566));
  nand_5 g02218(.A(pi732), .B(new_n4566), .Y(new_n4567));
  nand_5 g02219(.A(new_n4567), .B(new_n4565), .Y(new_n4568));
  nand_5 g02220(.A(new_n4568), .B(new_n4564), .Y(new_n4569));
  nor_5  g02221(.A(new_n4569), .B(new_n4562), .Y(new_n4570));
  nor_5  g02222(.A(new_n4570), .B(new_n4560), .Y(new_n4571));
  not_8  g02223(.A(new_n4571), .Y(new_n4572));
  nand_5 g02224(.A(new_n4572), .B(new_n4557), .Y(new_n4573));
  nand_5 g02225(.A(new_n4573), .B(new_n4556), .Y(new_n4574));
  xor_4  g02226(.A(new_n4574), .B(new_n4554), .Y(new_n4575));
  xor_4  g02227(.A(new_n4575), .B(new_n4552), .Y(new_n4576));
  xor_4  g02228(.A(new_n4549), .B(new_n4536), .Y(new_n4577));
  not_8  g02229(.A(new_n4577), .Y(new_n4578));
  xor_4  g02230(.A(new_n4571), .B(new_n4557), .Y(new_n4579));
  nand_5 g02231(.A(new_n4579), .B(new_n4578), .Y(new_n4580));
  not_8  g02232(.A(new_n4580), .Y(new_n4581));
  xor_4  g02233(.A(new_n4579), .B(new_n4578), .Y(new_n4582));
  not_8  g02234(.A(new_n4582), .Y(new_n4583));
  xor_4  g02235(.A(new_n4547), .B(new_n4539), .Y(new_n4584));
  xor_4  g02236(.A(new_n4569), .B(new_n4561), .Y(new_n4585));
  not_8  g02237(.A(new_n4585), .Y(new_n4586));
  nand_5 g02238(.A(new_n4586), .B(new_n4584), .Y(new_n4587));
  not_8  g02239(.A(new_n4584), .Y(new_n4588));
  xor_4  g02240(.A(new_n4585), .B(new_n4588), .Y(new_n4589));
  nand_5 g02241(.A(pi710), .B(new_n3556), .Y(new_n4590));
  not_8  g02242(.A(new_n4542), .Y(new_n4591));
  and_6  g02243(.A(new_n4565), .B(new_n4564), .Y(new_n4592));
  xor_4  g02244(.A(new_n4592), .B(new_n4591), .Y(new_n4593));
  nor_5  g02245(.A(pi732), .B(new_n4566), .Y(new_n4594));
  not_8  g02246(.A(new_n4594), .Y(new_n4595));
  nor_5  g02247(.A(new_n4595), .B(new_n4590), .Y(new_n4596));
  nand_5 g02248(.A(new_n4590), .B(new_n4544), .Y(new_n4597));
  nand_5 g02249(.A(new_n4595), .B(new_n4567), .Y(new_n4598));
  nor_5  g02250(.A(new_n4598), .B(new_n4597), .Y(new_n4599));
  nand_5 g02251(.A(new_n4595), .B(new_n4590), .Y(new_n4600));
  nor_5  g02252(.A(new_n4600), .B(new_n4599), .Y(new_n4601));
  nor_5  g02253(.A(new_n4601), .B(new_n4596), .Y(new_n4602));
  xor_4  g02254(.A(new_n4602), .B(new_n4593), .Y(new_n4603));
  nor_5  g02255(.A(new_n4603), .B(new_n4590), .Y(new_n4604));
  nand_5 g02256(.A(new_n4544), .B(new_n4542), .Y(new_n4605));
  nor_5  g02257(.A(new_n4605), .B(new_n4604), .Y(new_n4606));
  nor_5  g02258(.A(new_n4592), .B(new_n4542), .Y(new_n4607));
  nand_5 g02259(.A(new_n4601), .B(new_n4607), .Y(new_n4608));
  not_8  g02260(.A(new_n4590), .Y(new_n4609));
  nor_5  g02261(.A(new_n4609), .B(pi732), .Y(new_n4610));
  nand_5 g02262(.A(new_n4610), .B(new_n4591), .Y(new_n4611));
  nand_5 g02263(.A(new_n4611), .B(new_n4598), .Y(new_n4612));
  nand_5 g02264(.A(new_n4612), .B(new_n4592), .Y(new_n4613));
  nand_5 g02265(.A(new_n4613), .B(new_n4608), .Y(new_n4614));
  or_6   g02266(.A(new_n4614), .B(new_n4606), .Y(new_n4615));
  nand_5 g02267(.A(new_n4615), .B(new_n4589), .Y(new_n4616));
  nand_5 g02268(.A(new_n4616), .B(new_n4587), .Y(new_n4617));
  nor_5  g02269(.A(new_n4617), .B(new_n4583), .Y(new_n4618));
  nor_5  g02270(.A(new_n4618), .B(new_n4581), .Y(new_n4619));
  xor_4  g02271(.A(new_n4619), .B(new_n4576), .Y(new_n4620));
  not_8  g02272(.A(pi765), .Y(new_n4621));
  nand_5 g02273(.A(new_n4621), .B(pi386), .Y(new_n4622));
  not_8  g02274(.A(pi386), .Y(new_n4623));
  nand_5 g02275(.A(pi765), .B(new_n4623), .Y(new_n4624));
  nand_5 g02276(.A(new_n4624), .B(new_n4622), .Y(new_n4625));
  not_8  g02277(.A(pi682), .Y(new_n4626));
  nand_5 g02278(.A(new_n4626), .B(pi574), .Y(new_n4627));
  xor_4  g02279(.A(new_n4598), .B(new_n4597), .Y(new_n4628));
  nand_5 g02280(.A(new_n4628), .B(new_n4627), .Y(new_n4629));
  not_8  g02281(.A(new_n4628), .Y(new_n4630));
  not_8  g02282(.A(pi574), .Y(new_n4631));
  nand_5 g02283(.A(pi682), .B(new_n4631), .Y(new_n4632));
  nand_5 g02284(.A(new_n4632), .B(new_n4630), .Y(new_n4633));
  nand_5 g02285(.A(new_n4633), .B(new_n4629), .Y(new_n4634));
  xor_4  g02286(.A(new_n4634), .B(new_n4625), .Y(new_n4635));
  or_6   g02287(.A(new_n4635), .B(new_n4603), .Y(new_n4636));
  nand_5 g02288(.A(new_n4632), .B(new_n4627), .Y(new_n4637));
  nand_5 g02289(.A(new_n4637), .B(new_n4628), .Y(new_n4638));
  nand_5 g02290(.A(new_n4638), .B(new_n4635), .Y(new_n4639));
  nand_5 g02291(.A(new_n4639), .B(new_n4636), .Y(new_n4640));
  not_8  g02292(.A(pi052), .Y(new_n4641));
  xor_4  g02293(.A(pi546), .B(new_n4641), .Y(new_n4642));
  nand_5 g02294(.A(new_n4632), .B(new_n4624), .Y(new_n4643));
  nand_5 g02295(.A(new_n4643), .B(new_n4622), .Y(new_n4644));
  xor_4  g02296(.A(new_n4644), .B(new_n4642), .Y(new_n4645));
  not_8  g02297(.A(new_n4645), .Y(new_n4646));
  nand_5 g02298(.A(new_n4646), .B(new_n4640), .Y(new_n4647));
  xnor_4 g02299(.A(new_n4615), .B(new_n4589), .Y(new_n4648));
  xor_4  g02300(.A(new_n4645), .B(new_n4640), .Y(new_n4649));
  or_6   g02301(.A(new_n4649), .B(new_n4648), .Y(new_n4650));
  nand_5 g02302(.A(new_n4650), .B(new_n4647), .Y(new_n4651));
  not_8  g02303(.A(pi191), .Y(new_n4652));
  xor_4  g02304(.A(pi444), .B(new_n4652), .Y(new_n4653));
  nand_5 g02305(.A(pi546), .B(new_n4641), .Y(new_n4654));
  not_8  g02306(.A(new_n4654), .Y(new_n4655));
  not_8  g02307(.A(new_n4642), .Y(new_n4656));
  nor_5  g02308(.A(new_n4644), .B(new_n4656), .Y(new_n4657));
  nor_5  g02309(.A(new_n4657), .B(new_n4655), .Y(new_n4658));
  xor_4  g02310(.A(new_n4658), .B(new_n4653), .Y(new_n4659));
  not_8  g02311(.A(new_n4659), .Y(new_n4660));
  nand_5 g02312(.A(new_n4660), .B(new_n4651), .Y(new_n4661));
  xor_4  g02313(.A(new_n4617), .B(new_n4583), .Y(new_n4662));
  xor_4  g02314(.A(new_n4659), .B(new_n4651), .Y(new_n4663));
  or_6   g02315(.A(new_n4663), .B(new_n4662), .Y(new_n4664));
  nand_5 g02316(.A(new_n4664), .B(new_n4661), .Y(new_n4665));
  nand_5 g02317(.A(new_n4665), .B(new_n4620), .Y(new_n4666));
  not_8  g02318(.A(pi498), .Y(new_n4667));
  xor_4  g02319(.A(pi743), .B(new_n4667), .Y(new_n4668));
  not_8  g02320(.A(pi444), .Y(new_n4669));
  nand_5 g02321(.A(new_n4669), .B(pi191), .Y(new_n4670));
  not_8  g02322(.A(new_n4658), .Y(new_n4671));
  nand_5 g02323(.A(new_n4671), .B(new_n4653), .Y(new_n4672));
  nand_5 g02324(.A(new_n4672), .B(new_n4670), .Y(new_n4673));
  xnor_4 g02325(.A(new_n4673), .B(new_n4668), .Y(new_n4674));
  not_8  g02326(.A(new_n4620), .Y(new_n4675));
  xor_4  g02327(.A(new_n4665), .B(new_n4675), .Y(new_n4676));
  or_6   g02328(.A(new_n4676), .B(new_n4674), .Y(new_n4677));
  nand_5 g02329(.A(new_n4677), .B(new_n4666), .Y(new_n4678));
  not_8  g02330(.A(pi522), .Y(new_n4679));
  nand_5 g02331(.A(new_n4679), .B(pi453), .Y(new_n4680));
  nand_5 g02332(.A(new_n4551), .B(new_n4533), .Y(new_n4681));
  nand_5 g02333(.A(new_n4681), .B(new_n4680), .Y(new_n4682));
  not_8  g02334(.A(pi040), .Y(new_n4683));
  nand_5 g02335(.A(pi138), .B(new_n4683), .Y(new_n4684));
  nand_5 g02336(.A(new_n3539), .B(pi040), .Y(new_n4685));
  nand_5 g02337(.A(new_n4685), .B(new_n4684), .Y(new_n4686));
  xor_4  g02338(.A(new_n4686), .B(new_n4682), .Y(new_n4687));
  or_6   g02339(.A(pi750), .B(new_n4553), .Y(new_n4688));
  nand_5 g02340(.A(new_n4574), .B(new_n4554), .Y(new_n4689));
  nand_5 g02341(.A(new_n4689), .B(new_n4688), .Y(new_n4690));
  not_8  g02342(.A(pi140), .Y(new_n4691));
  or_6   g02343(.A(pi402), .B(new_n4691), .Y(new_n4692));
  nand_5 g02344(.A(pi402), .B(new_n4691), .Y(new_n4693));
  and_6  g02345(.A(new_n4693), .B(new_n4692), .Y(new_n4694));
  xor_4  g02346(.A(new_n4694), .B(new_n4690), .Y(new_n4695));
  not_8  g02347(.A(new_n4695), .Y(new_n4696));
  xor_4  g02348(.A(new_n4696), .B(new_n4687), .Y(new_n4697));
  not_8  g02349(.A(new_n4552), .Y(new_n4698));
  not_8  g02350(.A(new_n4575), .Y(new_n4699));
  nand_5 g02351(.A(new_n4699), .B(new_n4698), .Y(new_n4700));
  not_8  g02352(.A(new_n4619), .Y(new_n4701));
  nand_5 g02353(.A(new_n4701), .B(new_n4576), .Y(new_n4702));
  and_6  g02354(.A(new_n4702), .B(new_n4700), .Y(new_n4703));
  xnor_4 g02355(.A(new_n4703), .B(new_n4697), .Y(new_n4704));
  not_8  g02356(.A(pi743), .Y(new_n4705));
  nand_5 g02357(.A(new_n4705), .B(pi498), .Y(new_n4706));
  nand_5 g02358(.A(new_n4673), .B(new_n4668), .Y(new_n4707));
  nand_5 g02359(.A(new_n4707), .B(new_n4706), .Y(new_n4708));
  not_8  g02360(.A(pi630), .Y(new_n4709));
  or_6   g02361(.A(pi657), .B(new_n4709), .Y(new_n4710));
  nand_5 g02362(.A(pi657), .B(new_n4709), .Y(new_n4711));
  nand_5 g02363(.A(new_n4711), .B(new_n4710), .Y(new_n4712));
  xor_4  g02364(.A(new_n4712), .B(new_n4708), .Y(new_n4713));
  xor_4  g02365(.A(new_n4713), .B(new_n4704), .Y(new_n4714));
  xnor_4 g02366(.A(new_n4714), .B(new_n4678), .Y(po0012));
  nand_5 g02367(.A(pi323), .B(pi118), .Y(new_n4716));
  xor_4  g02368(.A(pi323), .B(pi118), .Y(new_n4717));
  nand_5 g02369(.A(pi556), .B(pi466), .Y(new_n4718));
  xor_4  g02370(.A(pi556), .B(pi466), .Y(new_n4719));
  nor_5  g02371(.A(pi809), .B(pi553), .Y(new_n4720));
  not_8  g02372(.A(pi553), .Y(new_n4721));
  xor_4  g02373(.A(pi809), .B(new_n4721), .Y(new_n4722));
  nand_5 g02374(.A(pi757), .B(pi583), .Y(new_n4723));
  not_8  g02375(.A(pi583), .Y(new_n4724));
  not_8  g02376(.A(pi757), .Y(new_n4725));
  nand_5 g02377(.A(new_n4725), .B(new_n4724), .Y(new_n4726));
  nand_5 g02378(.A(pi695), .B(pi655), .Y(new_n4727));
  nand_5 g02379(.A(new_n3712), .B(new_n3460), .Y(new_n4728));
  nand_5 g02380(.A(pi805), .B(pi531), .Y(new_n4729));
  xor_4  g02381(.A(pi805), .B(pi531), .Y(new_n4730));
  nor_5  g02382(.A(pi464), .B(pi006), .Y(new_n4731));
  nor_5  g02383(.A(pi818), .B(pi330), .Y(new_n4732));
  xor_4  g02384(.A(pi818), .B(pi330), .Y(new_n4733));
  nand_5 g02385(.A(pi523), .B(pi158), .Y(new_n4734));
  and_6  g02386(.A(new_n4734), .B(new_n4733), .Y(new_n4735));
  nor_5  g02387(.A(new_n4735), .B(new_n4732), .Y(new_n4736));
  xor_4  g02388(.A(pi464), .B(new_n3720), .Y(new_n4737));
  nor_5  g02389(.A(new_n4737), .B(new_n4736), .Y(new_n4738));
  nor_5  g02390(.A(new_n4738), .B(new_n4731), .Y(new_n4739));
  nand_5 g02391(.A(new_n4739), .B(new_n4730), .Y(new_n4740));
  nand_5 g02392(.A(new_n4740), .B(new_n4729), .Y(new_n4741));
  nand_5 g02393(.A(new_n4741), .B(new_n4728), .Y(new_n4742));
  nand_5 g02394(.A(new_n4742), .B(new_n4727), .Y(new_n4743));
  nand_5 g02395(.A(new_n4743), .B(new_n4726), .Y(new_n4744));
  nand_5 g02396(.A(new_n4744), .B(new_n4723), .Y(new_n4745));
  nor_5  g02397(.A(new_n4745), .B(new_n4722), .Y(new_n4746));
  nor_5  g02398(.A(new_n4746), .B(new_n4720), .Y(new_n4747));
  nand_5 g02399(.A(new_n4747), .B(new_n4719), .Y(new_n4748));
  nand_5 g02400(.A(new_n4748), .B(new_n4718), .Y(new_n4749));
  nand_5 g02401(.A(new_n4749), .B(new_n4717), .Y(new_n4750));
  nand_5 g02402(.A(new_n4750), .B(new_n4716), .Y(new_n4751));
  not_8  g02403(.A(new_n4751), .Y(new_n4752));
  xor_4  g02404(.A(pi623), .B(pi547), .Y(new_n4753));
  not_8  g02405(.A(pi236), .Y(new_n4754));
  nand_5 g02406(.A(new_n3709), .B(new_n4754), .Y(new_n4755));
  not_8  g02407(.A(pi103), .Y(new_n4756));
  not_8  g02408(.A(pi375), .Y(new_n4757));
  nand_5 g02409(.A(new_n4757), .B(new_n4756), .Y(new_n4758));
  xor_4  g02410(.A(pi375), .B(pi103), .Y(new_n4759));
  not_8  g02411(.A(pi427), .Y(new_n4760));
  nand_5 g02412(.A(new_n4760), .B(new_n3763), .Y(new_n4761));
  nand_5 g02413(.A(pi427), .B(pi298), .Y(new_n4762));
  not_8  g02414(.A(pi237), .Y(new_n4763));
  nand_5 g02415(.A(new_n4763), .B(new_n3758), .Y(new_n4764));
  not_8  g02416(.A(new_n4764), .Y(new_n4765));
  nor_5  g02417(.A(pi599), .B(pi241), .Y(new_n4766));
  xor_4  g02418(.A(pi599), .B(pi241), .Y(new_n4767));
  not_8  g02419(.A(new_n4767), .Y(new_n4768));
  nor_5  g02420(.A(pi488), .B(pi091), .Y(new_n4769));
  not_8  g02421(.A(pi091), .Y(new_n4770));
  xor_4  g02422(.A(pi488), .B(new_n4770), .Y(new_n4771));
  nand_5 g02423(.A(pi631), .B(pi482), .Y(new_n4772));
  not_8  g02424(.A(new_n4772), .Y(new_n4773));
  nor_5  g02425(.A(new_n4773), .B(new_n4771), .Y(new_n4774));
  nor_5  g02426(.A(new_n4774), .B(new_n4769), .Y(new_n4775));
  nor_5  g02427(.A(new_n4775), .B(new_n4768), .Y(new_n4776));
  nor_5  g02428(.A(new_n4776), .B(new_n4766), .Y(new_n4777));
  xor_4  g02429(.A(pi237), .B(new_n3758), .Y(new_n4778));
  nor_5  g02430(.A(new_n4778), .B(new_n4777), .Y(new_n4779));
  nor_5  g02431(.A(new_n4779), .B(new_n4765), .Y(new_n4780));
  not_8  g02432(.A(new_n4780), .Y(new_n4781));
  nand_5 g02433(.A(new_n4781), .B(new_n4762), .Y(new_n4782));
  nand_5 g02434(.A(new_n4782), .B(new_n4761), .Y(new_n4783));
  nand_5 g02435(.A(new_n4783), .B(new_n4759), .Y(new_n4784));
  nand_5 g02436(.A(new_n4784), .B(new_n4758), .Y(new_n4785));
  xor_4  g02437(.A(pi793), .B(new_n4754), .Y(new_n4786));
  not_8  g02438(.A(new_n4786), .Y(new_n4787));
  nand_5 g02439(.A(new_n4787), .B(new_n4785), .Y(new_n4788));
  nand_5 g02440(.A(new_n4788), .B(new_n4755), .Y(new_n4789));
  xor_4  g02441(.A(new_n4789), .B(new_n4753), .Y(new_n4790));
  not_8  g02442(.A(new_n4790), .Y(new_n4791));
  xor_4  g02443(.A(new_n4786), .B(new_n4785), .Y(new_n4792));
  xor_4  g02444(.A(new_n4783), .B(new_n4759), .Y(new_n4793));
  not_8  g02445(.A(new_n4793), .Y(new_n4794));
  not_8  g02446(.A(pi681), .Y(new_n4795));
  xor_4  g02447(.A(pi631), .B(pi482), .Y(new_n4796));
  not_8  g02448(.A(new_n4796), .Y(new_n4797));
  nor_5  g02449(.A(new_n4797), .B(new_n3493), .Y(new_n4798));
  nand_5 g02450(.A(new_n4798), .B(pi787), .Y(new_n4799));
  xor_4  g02451(.A(new_n4798), .B(pi787), .Y(new_n4800));
  xor_4  g02452(.A(new_n4773), .B(new_n4771), .Y(new_n4801));
  not_8  g02453(.A(new_n4801), .Y(new_n4802));
  nand_5 g02454(.A(new_n4802), .B(new_n4800), .Y(new_n4803));
  nand_5 g02455(.A(new_n4803), .B(new_n4799), .Y(new_n4804));
  xor_4  g02456(.A(new_n4775), .B(new_n4767), .Y(new_n4805));
  nor_5  g02457(.A(new_n4805), .B(new_n4804), .Y(new_n4806));
  nor_5  g02458(.A(new_n4806), .B(new_n3489), .Y(new_n4807));
  nand_5 g02459(.A(new_n4805), .B(new_n4804), .Y(new_n4808));
  not_8  g02460(.A(new_n4808), .Y(new_n4809));
  nor_5  g02461(.A(new_n4809), .B(new_n4807), .Y(new_n4810));
  nand_5 g02462(.A(new_n4810), .B(new_n4795), .Y(new_n4811));
  xor_4  g02463(.A(new_n4778), .B(new_n4777), .Y(new_n4812));
  not_8  g02464(.A(new_n4812), .Y(new_n4813));
  xor_4  g02465(.A(new_n4810), .B(pi681), .Y(new_n4814));
  or_6   g02466(.A(new_n4814), .B(new_n4813), .Y(new_n4815));
  nand_5 g02467(.A(new_n4815), .B(new_n4811), .Y(new_n4816));
  nand_5 g02468(.A(new_n4762), .B(new_n4761), .Y(new_n4817));
  xor_4  g02469(.A(new_n4817), .B(new_n4780), .Y(new_n4818));
  or_6   g02470(.A(new_n4818), .B(new_n4816), .Y(new_n4819));
  nand_5 g02471(.A(new_n4818), .B(new_n4816), .Y(new_n4820));
  nand_5 g02472(.A(new_n4820), .B(pi317), .Y(new_n4821));
  nand_5 g02473(.A(new_n4821), .B(new_n4819), .Y(new_n4822));
  nand_5 g02474(.A(new_n4822), .B(new_n4794), .Y(new_n4823));
  or_6   g02475(.A(new_n4822), .B(new_n4794), .Y(new_n4824));
  nand_5 g02476(.A(new_n4824), .B(pi246), .Y(new_n4825));
  nand_5 g02477(.A(new_n4825), .B(new_n4823), .Y(new_n4826));
  nand_5 g02478(.A(new_n4826), .B(new_n4792), .Y(new_n4827));
  not_8  g02479(.A(pi441), .Y(new_n4828));
  not_8  g02480(.A(new_n4792), .Y(new_n4829));
  xor_4  g02481(.A(new_n4826), .B(new_n4829), .Y(new_n4830));
  or_6   g02482(.A(new_n4830), .B(new_n4828), .Y(new_n4831));
  nand_5 g02483(.A(new_n4831), .B(new_n4827), .Y(new_n4832));
  or_6   g02484(.A(new_n4832), .B(new_n4791), .Y(new_n4833));
  nand_5 g02485(.A(new_n4833), .B(pi616), .Y(new_n4834));
  nand_5 g02486(.A(new_n4832), .B(new_n4791), .Y(new_n4835));
  nand_5 g02487(.A(new_n4835), .B(new_n4834), .Y(new_n4836));
  nand_5 g02488(.A(pi812), .B(pi013), .Y(new_n4837));
  not_8  g02489(.A(pi013), .Y(new_n4838));
  not_8  g02490(.A(pi812), .Y(new_n4839));
  nand_5 g02491(.A(new_n4839), .B(new_n4838), .Y(new_n4840));
  nand_5 g02492(.A(new_n4840), .B(new_n4837), .Y(new_n4841));
  not_8  g02493(.A(pi547), .Y(new_n4842));
  not_8  g02494(.A(pi623), .Y(new_n4843));
  nand_5 g02495(.A(new_n4843), .B(new_n4842), .Y(new_n4844));
  nand_5 g02496(.A(new_n4789), .B(new_n4753), .Y(new_n4845));
  nand_5 g02497(.A(new_n4845), .B(new_n4844), .Y(new_n4846));
  not_8  g02498(.A(new_n4846), .Y(new_n4847));
  xor_4  g02499(.A(new_n4847), .B(new_n4841), .Y(new_n4848));
  not_8  g02500(.A(new_n4848), .Y(new_n4849));
  or_6   g02501(.A(new_n4849), .B(new_n4836), .Y(new_n4850));
  nand_5 g02502(.A(new_n4850), .B(pi650), .Y(new_n4851));
  nand_5 g02503(.A(new_n4849), .B(new_n4836), .Y(new_n4852));
  nand_5 g02504(.A(new_n4852), .B(new_n4851), .Y(new_n4853));
  nor_5  g02505(.A(new_n4853), .B(pi303), .Y(new_n4854));
  xor_4  g02506(.A(new_n4853), .B(new_n3423), .Y(new_n4855));
  nand_5 g02507(.A(pi315), .B(pi097), .Y(new_n4856));
  not_8  g02508(.A(pi097), .Y(new_n4857));
  not_8  g02509(.A(pi315), .Y(new_n4858));
  nand_5 g02510(.A(new_n4858), .B(new_n4857), .Y(new_n4859));
  and_6  g02511(.A(new_n4859), .B(new_n4856), .Y(new_n4860));
  nand_5 g02512(.A(new_n4846), .B(new_n4837), .Y(new_n4861));
  nand_5 g02513(.A(new_n4861), .B(new_n4840), .Y(new_n4862));
  xor_4  g02514(.A(new_n4862), .B(new_n4860), .Y(new_n4863));
  not_8  g02515(.A(new_n4863), .Y(new_n4864));
  nor_5  g02516(.A(new_n4864), .B(new_n4855), .Y(new_n4865));
  or_6   g02517(.A(new_n4865), .B(new_n4854), .Y(new_n4866));
  nand_5 g02518(.A(new_n4862), .B(new_n4856), .Y(new_n4867));
  nand_5 g02519(.A(new_n4867), .B(new_n4859), .Y(new_n4868));
  nand_5 g02520(.A(new_n4868), .B(new_n4866), .Y(new_n4869));
  not_8  g02521(.A(new_n4869), .Y(new_n4870));
  nor_5  g02522(.A(new_n4868), .B(new_n4866), .Y(new_n4871));
  nor_5  g02523(.A(new_n4871), .B(new_n4870), .Y(new_n4872));
  not_8  g02524(.A(pi124), .Y(new_n4873));
  nand_5 g02525(.A(new_n4835), .B(new_n4833), .Y(new_n4874));
  xor_4  g02526(.A(new_n4874), .B(pi616), .Y(new_n4875));
  nor_5  g02527(.A(new_n4875), .B(pi086), .Y(new_n4876));
  xor_4  g02528(.A(new_n4830), .B(pi441), .Y(new_n4877));
  nor_5  g02529(.A(new_n4877), .B(pi752), .Y(new_n4878));
  not_8  g02530(.A(pi752), .Y(new_n4879));
  xor_4  g02531(.A(new_n4877), .B(new_n4879), .Y(new_n4880));
  not_8  g02532(.A(pi676), .Y(new_n4881));
  xor_4  g02533(.A(new_n4801), .B(new_n4800), .Y(new_n4882));
  nand_5 g02534(.A(new_n4882), .B(pi619), .Y(new_n4883));
  not_8  g02535(.A(pi619), .Y(new_n4884));
  xor_4  g02536(.A(new_n4882), .B(new_n4884), .Y(new_n4885));
  not_8  g02537(.A(pi130), .Y(new_n4886));
  xor_4  g02538(.A(new_n4796), .B(pi670), .Y(new_n4887));
  nand_5 g02539(.A(new_n4887), .B(new_n4886), .Y(new_n4888));
  not_8  g02540(.A(new_n4888), .Y(new_n4889));
  or_6   g02541(.A(new_n4889), .B(new_n4885), .Y(new_n4890));
  nand_5 g02542(.A(new_n4890), .B(new_n4883), .Y(new_n4891));
  nor_5  g02543(.A(new_n4809), .B(new_n4806), .Y(new_n4892));
  xor_4  g02544(.A(new_n4892), .B(new_n3489), .Y(new_n4893));
  nand_5 g02545(.A(new_n4893), .B(new_n4891), .Y(new_n4894));
  or_6   g02546(.A(new_n4893), .B(new_n4891), .Y(new_n4895));
  nand_5 g02547(.A(new_n4895), .B(pi796), .Y(new_n4896));
  nand_5 g02548(.A(new_n4896), .B(new_n4894), .Y(new_n4897));
  nor_5  g02549(.A(new_n4897), .B(pi232), .Y(new_n4898));
  xor_4  g02550(.A(new_n4814), .B(new_n4813), .Y(new_n4899));
  not_8  g02551(.A(pi232), .Y(new_n4900));
  xor_4  g02552(.A(new_n4897), .B(new_n4900), .Y(new_n4901));
  nor_5  g02553(.A(new_n4901), .B(new_n4899), .Y(new_n4902));
  or_6   g02554(.A(new_n4902), .B(new_n4898), .Y(new_n4903));
  not_8  g02555(.A(pi317), .Y(new_n4904));
  nand_5 g02556(.A(new_n4820), .B(new_n4819), .Y(new_n4905));
  xor_4  g02557(.A(new_n4905), .B(new_n4904), .Y(new_n4906));
  nand_5 g02558(.A(new_n4906), .B(new_n4903), .Y(new_n4907));
  not_8  g02559(.A(pi634), .Y(new_n4908));
  or_6   g02560(.A(new_n4906), .B(new_n4903), .Y(new_n4909));
  nand_5 g02561(.A(new_n4909), .B(new_n4908), .Y(new_n4910));
  nand_5 g02562(.A(new_n4910), .B(new_n4907), .Y(new_n4911));
  nand_5 g02563(.A(new_n4911), .B(new_n4881), .Y(new_n4912));
  xor_4  g02564(.A(new_n4911), .B(new_n4881), .Y(new_n4913));
  not_8  g02565(.A(new_n4913), .Y(new_n4914));
  nand_5 g02566(.A(new_n4823), .B(new_n4824), .Y(new_n4915));
  xor_4  g02567(.A(new_n4915), .B(pi246), .Y(new_n4916));
  or_6   g02568(.A(new_n4916), .B(new_n4914), .Y(new_n4917));
  nand_5 g02569(.A(new_n4917), .B(new_n4912), .Y(new_n4918));
  not_8  g02570(.A(new_n4918), .Y(new_n4919));
  nor_5  g02571(.A(new_n4919), .B(new_n4880), .Y(new_n4920));
  nor_5  g02572(.A(new_n4920), .B(new_n4878), .Y(new_n4921));
  not_8  g02573(.A(pi086), .Y(new_n4922));
  xor_4  g02574(.A(new_n4875), .B(new_n4922), .Y(new_n4923));
  nor_5  g02575(.A(new_n4923), .B(new_n4921), .Y(new_n4924));
  or_6   g02576(.A(new_n4924), .B(new_n4876), .Y(new_n4925));
  nand_5 g02577(.A(new_n4852), .B(new_n4850), .Y(new_n4926));
  xor_4  g02578(.A(new_n4926), .B(pi650), .Y(new_n4927));
  not_8  g02579(.A(new_n4927), .Y(new_n4928));
  nand_5 g02580(.A(new_n4928), .B(new_n4925), .Y(new_n4929));
  not_8  g02581(.A(pi093), .Y(new_n4930));
  or_6   g02582(.A(new_n4928), .B(new_n4925), .Y(new_n4931));
  nand_5 g02583(.A(new_n4931), .B(new_n4930), .Y(new_n4932));
  nand_5 g02584(.A(new_n4932), .B(new_n4929), .Y(new_n4933));
  or_6   g02585(.A(new_n4933), .B(new_n4873), .Y(new_n4934));
  xor_4  g02586(.A(new_n4864), .B(new_n4855), .Y(new_n4935));
  not_8  g02587(.A(new_n4935), .Y(new_n4936));
  xor_4  g02588(.A(new_n4933), .B(pi124), .Y(new_n4937));
  or_6   g02589(.A(new_n4937), .B(new_n4936), .Y(new_n4938));
  nand_5 g02590(.A(new_n4938), .B(new_n4934), .Y(new_n4939));
  xor_4  g02591(.A(new_n4939), .B(new_n4872), .Y(new_n4940));
  xor_4  g02592(.A(new_n4940), .B(new_n4752), .Y(new_n4941));
  not_8  g02593(.A(new_n4941), .Y(new_n4942));
  xor_4  g02594(.A(new_n4937), .B(new_n4935), .Y(new_n4943));
  xor_4  g02595(.A(new_n4749), .B(new_n4717), .Y(new_n4944));
  not_8  g02596(.A(new_n4944), .Y(new_n4945));
  nand_5 g02597(.A(new_n4945), .B(new_n4943), .Y(new_n4946));
  xor_4  g02598(.A(new_n4747), .B(new_n4719), .Y(new_n4947));
  not_8  g02599(.A(new_n4947), .Y(new_n4948));
  nand_5 g02600(.A(new_n4931), .B(new_n4929), .Y(new_n4949));
  xor_4  g02601(.A(new_n4949), .B(pi093), .Y(new_n4950));
  and_6  g02602(.A(new_n4950), .B(new_n4948), .Y(new_n4951));
  xor_4  g02603(.A(new_n4950), .B(new_n4947), .Y(new_n4952));
  xor_4  g02604(.A(new_n4745), .B(new_n4722), .Y(new_n4953));
  not_8  g02605(.A(new_n4953), .Y(new_n4954));
  xnor_4 g02606(.A(new_n4923), .B(new_n4921), .Y(new_n4955));
  nor_5  g02607(.A(new_n4955), .B(new_n4954), .Y(new_n4956));
  xor_4  g02608(.A(new_n4955), .B(new_n4953), .Y(new_n4957));
  xor_4  g02609(.A(new_n4918), .B(new_n4880), .Y(new_n4958));
  and_6  g02610(.A(new_n4723), .B(new_n4726), .Y(new_n4959));
  xor_4  g02611(.A(new_n4959), .B(new_n4743), .Y(new_n4960));
  nor_5  g02612(.A(new_n4960), .B(new_n4958), .Y(new_n4961));
  nand_5 g02613(.A(new_n4960), .B(new_n4958), .Y(new_n4962));
  xor_4  g02614(.A(new_n4916), .B(new_n4913), .Y(new_n4963));
  nand_5 g02615(.A(new_n4728), .B(new_n4727), .Y(new_n4964));
  xor_4  g02616(.A(new_n4964), .B(new_n4741), .Y(new_n4965));
  not_8  g02617(.A(new_n4965), .Y(new_n4966));
  nor_5  g02618(.A(new_n4966), .B(new_n4963), .Y(new_n4967));
  xor_4  g02619(.A(new_n4965), .B(new_n4963), .Y(new_n4968));
  xor_4  g02620(.A(new_n4739), .B(new_n4730), .Y(new_n4969));
  not_8  g02621(.A(new_n4969), .Y(new_n4970));
  nand_5 g02622(.A(new_n4909), .B(new_n4907), .Y(new_n4971));
  xor_4  g02623(.A(new_n4971), .B(pi634), .Y(new_n4972));
  and_6  g02624(.A(new_n4972), .B(new_n4970), .Y(new_n4973));
  xor_4  g02625(.A(new_n4972), .B(new_n4969), .Y(new_n4974));
  xor_4  g02626(.A(new_n4737), .B(new_n4736), .Y(new_n4975));
  not_8  g02627(.A(new_n4975), .Y(new_n4976));
  xnor_4 g02628(.A(new_n4901), .B(new_n4899), .Y(new_n4977));
  nand_5 g02629(.A(new_n4977), .B(new_n4976), .Y(new_n4978));
  nand_5 g02630(.A(new_n4895), .B(new_n4894), .Y(new_n4979));
  xor_4  g02631(.A(new_n4979), .B(pi796), .Y(new_n4980));
  nor_5  g02632(.A(new_n4980), .B(new_n4733), .Y(new_n4981));
  nor_5  g02633(.A(new_n4981), .B(new_n4735), .Y(new_n4982));
  not_8  g02634(.A(pi523), .Y(new_n4983));
  nand_5 g02635(.A(new_n4983), .B(new_n3728), .Y(new_n4984));
  nand_5 g02636(.A(pi301), .B(pi259), .Y(new_n4985));
  xor_4  g02637(.A(new_n4887), .B(new_n4886), .Y(new_n4986));
  nand_5 g02638(.A(new_n3491), .B(new_n3730), .Y(new_n4987));
  nand_5 g02639(.A(new_n4987), .B(new_n4985), .Y(new_n4988));
  or_6   g02640(.A(new_n4988), .B(new_n4986), .Y(new_n4989));
  nand_5 g02641(.A(new_n4989), .B(new_n4985), .Y(new_n4990));
  not_8  g02642(.A(new_n4990), .Y(new_n4991));
  xor_4  g02643(.A(new_n4888), .B(new_n4885), .Y(new_n4992));
  nand_5 g02644(.A(new_n4992), .B(new_n4991), .Y(new_n4993));
  nand_5 g02645(.A(new_n4993), .B(new_n4984), .Y(new_n4994));
  nor_5  g02646(.A(new_n4994), .B(new_n4982), .Y(new_n4995));
  xor_4  g02647(.A(new_n4734), .B(new_n4733), .Y(new_n4996));
  or_6   g02648(.A(new_n4996), .B(new_n4980), .Y(new_n4997));
  xnor_4 g02649(.A(new_n4996), .B(new_n4980), .Y(new_n4998));
  or_6   g02650(.A(new_n4992), .B(new_n4991), .Y(new_n4999));
  or_6   g02651(.A(new_n4999), .B(new_n4998), .Y(new_n5000));
  nand_5 g02652(.A(new_n5000), .B(new_n4997), .Y(new_n5001));
  nor_5  g02653(.A(new_n5001), .B(new_n4995), .Y(new_n5002));
  xor_4  g02654(.A(new_n4977), .B(new_n4976), .Y(new_n5003));
  not_8  g02655(.A(new_n5003), .Y(new_n5004));
  or_6   g02656(.A(new_n5004), .B(new_n5002), .Y(new_n5005));
  nand_5 g02657(.A(new_n5005), .B(new_n4978), .Y(new_n5006));
  nor_5  g02658(.A(new_n5006), .B(new_n4974), .Y(new_n5007));
  nor_5  g02659(.A(new_n5007), .B(new_n4973), .Y(new_n5008));
  nor_5  g02660(.A(new_n5008), .B(new_n4968), .Y(new_n5009));
  or_6   g02661(.A(new_n5009), .B(new_n4967), .Y(new_n5010));
  and_6  g02662(.A(new_n5010), .B(new_n4962), .Y(new_n5011));
  nor_5  g02663(.A(new_n5011), .B(new_n4961), .Y(new_n5012));
  nor_5  g02664(.A(new_n5012), .B(new_n4957), .Y(new_n5013));
  nor_5  g02665(.A(new_n5013), .B(new_n4956), .Y(new_n5014));
  nor_5  g02666(.A(new_n5014), .B(new_n4952), .Y(new_n5015));
  nor_5  g02667(.A(new_n5015), .B(new_n4951), .Y(new_n5016));
  xor_4  g02668(.A(new_n4944), .B(new_n4943), .Y(new_n5017));
  or_6   g02669(.A(new_n5017), .B(new_n5016), .Y(new_n5018));
  nand_5 g02670(.A(new_n5018), .B(new_n4946), .Y(new_n5019));
  xor_4  g02671(.A(new_n5019), .B(new_n4942), .Y(po0013));
  not_8  g02672(.A(pi276), .Y(new_n5021));
  xor_4  g02673(.A(pi550), .B(pi501), .Y(new_n5022));
  nor_5  g02674(.A(pi589), .B(pi209), .Y(new_n5023));
  nand_5 g02675(.A(pi491), .B(pi077), .Y(new_n5024));
  not_8  g02676(.A(new_n5024), .Y(new_n5025));
  not_8  g02677(.A(pi209), .Y(new_n5026));
  xor_4  g02678(.A(pi589), .B(new_n5026), .Y(new_n5027));
  nor_5  g02679(.A(new_n5027), .B(new_n5025), .Y(new_n5028));
  nor_5  g02680(.A(new_n5028), .B(new_n5023), .Y(new_n5029));
  xor_4  g02681(.A(new_n5029), .B(new_n5022), .Y(new_n5030));
  not_8  g02682(.A(pi617), .Y(new_n5031));
  xor_4  g02683(.A(pi491), .B(pi077), .Y(new_n5032));
  not_8  g02684(.A(new_n5032), .Y(new_n5033));
  nor_5  g02685(.A(new_n5033), .B(pi396), .Y(new_n5034));
  nand_5 g02686(.A(new_n5034), .B(new_n5031), .Y(new_n5035));
  xor_4  g02687(.A(new_n5027), .B(new_n5025), .Y(new_n5036));
  not_8  g02688(.A(new_n5036), .Y(new_n5037));
  xor_4  g02689(.A(new_n5034), .B(new_n5031), .Y(new_n5038));
  nand_5 g02690(.A(new_n5038), .B(new_n5037), .Y(new_n5039));
  nand_5 g02691(.A(new_n5039), .B(new_n5035), .Y(new_n5040));
  xor_4  g02692(.A(new_n5040), .B(new_n5030), .Y(new_n5041));
  xor_4  g02693(.A(new_n5041), .B(new_n5021), .Y(new_n5042));
  not_8  g02694(.A(pi654), .Y(new_n5043));
  nand_5 g02695(.A(new_n5043), .B(pi508), .Y(new_n5044));
  nand_5 g02696(.A(new_n3239), .B(pi733), .Y(new_n5045));
  not_8  g02697(.A(pi733), .Y(new_n5046));
  nand_5 g02698(.A(pi783), .B(new_n5046), .Y(new_n5047));
  and_6  g02699(.A(new_n5047), .B(new_n5045), .Y(new_n5048));
  xor_4  g02700(.A(new_n5048), .B(new_n5044), .Y(new_n5049));
  not_8  g02701(.A(new_n5049), .Y(new_n5050));
  or_6   g02702(.A(new_n5050), .B(pi711), .Y(new_n5051));
  nand_5 g02703(.A(new_n5050), .B(pi711), .Y(new_n5052));
  nand_5 g02704(.A(new_n5052), .B(new_n5051), .Y(new_n5053));
  not_8  g02705(.A(new_n5053), .Y(new_n5054));
  not_8  g02706(.A(pi540), .Y(new_n5055));
  xor_4  g02707(.A(pi654), .B(new_n3339), .Y(new_n5056));
  nand_5 g02708(.A(new_n5056), .B(new_n5055), .Y(new_n5057));
  not_8  g02709(.A(pi396), .Y(new_n5058));
  xor_4  g02710(.A(new_n5032), .B(new_n5058), .Y(new_n5059));
  nor_5  g02711(.A(new_n5056), .B(pi540), .Y(new_n5060));
  not_8  g02712(.A(new_n5060), .Y(new_n5061));
  nand_5 g02713(.A(new_n5056), .B(pi540), .Y(new_n5062));
  nand_5 g02714(.A(new_n5062), .B(new_n5061), .Y(new_n5063));
  nand_5 g02715(.A(new_n5063), .B(new_n5059), .Y(new_n5064));
  nand_5 g02716(.A(new_n5064), .B(new_n5057), .Y(new_n5065));
  or_6   g02717(.A(new_n5065), .B(new_n5054), .Y(new_n5066));
  xor_4  g02718(.A(new_n5038), .B(new_n5037), .Y(new_n5067));
  not_8  g02719(.A(new_n5067), .Y(new_n5068));
  xor_4  g02720(.A(new_n5065), .B(new_n5054), .Y(new_n5069));
  nand_5 g02721(.A(new_n5069), .B(new_n5068), .Y(new_n5070));
  nand_5 g02722(.A(new_n5070), .B(new_n5066), .Y(new_n5071));
  nand_5 g02723(.A(new_n5049), .B(pi711), .Y(new_n5072));
  not_8  g02724(.A(pi355), .Y(new_n5073));
  xor_4  g02725(.A(pi468), .B(pi127), .Y(new_n5074));
  nand_5 g02726(.A(new_n5047), .B(new_n5044), .Y(new_n5075));
  nand_5 g02727(.A(new_n5075), .B(new_n5045), .Y(new_n5076));
  xor_4  g02728(.A(new_n5076), .B(new_n5074), .Y(new_n5077));
  xor_4  g02729(.A(new_n5077), .B(new_n5073), .Y(new_n5078));
  xor_4  g02730(.A(new_n5078), .B(new_n5072), .Y(new_n5079));
  xor_4  g02731(.A(new_n5079), .B(new_n5071), .Y(new_n5080));
  xor_4  g02732(.A(new_n5080), .B(new_n5042), .Y(po0014));
  xor_4  g02733(.A(pi191), .B(pi102), .Y(new_n5082));
  not_8  g02734(.A(pi546), .Y(new_n5083));
  nor_5  g02735(.A(new_n5083), .B(new_n2482), .Y(new_n5084));
  nand_5 g02736(.A(pi765), .B(pi612), .Y(new_n5085));
  xor_4  g02737(.A(pi765), .B(pi612), .Y(new_n5086));
  nand_5 g02738(.A(pi682), .B(pi302), .Y(new_n5087));
  not_8  g02739(.A(new_n5087), .Y(new_n5088));
  nand_5 g02740(.A(new_n5088), .B(new_n5086), .Y(new_n5089));
  and_6  g02741(.A(new_n5089), .B(new_n5085), .Y(new_n5090));
  xor_4  g02742(.A(pi546), .B(new_n2482), .Y(new_n5091));
  nor_5  g02743(.A(new_n5091), .B(new_n5090), .Y(new_n5092));
  nor_5  g02744(.A(new_n5092), .B(new_n5084), .Y(new_n5093));
  xor_4  g02745(.A(new_n5093), .B(new_n5082), .Y(new_n5094));
  xor_4  g02746(.A(new_n5091), .B(new_n5090), .Y(new_n5095));
  or_6   g02747(.A(new_n5095), .B(new_n3166), .Y(new_n5096));
  nand_5 g02748(.A(new_n5095), .B(new_n3166), .Y(new_n5097));
  nor_5  g02749(.A(pi682), .B(pi302), .Y(new_n5098));
  or_6   g02750(.A(new_n5098), .B(new_n5088), .Y(new_n5099));
  nor_5  g02751(.A(new_n5099), .B(new_n3169), .Y(new_n5100));
  nor_5  g02752(.A(new_n5100), .B(new_n5088), .Y(new_n5101));
  not_8  g02753(.A(new_n5101), .Y(new_n5102));
  xor_4  g02754(.A(new_n5086), .B(new_n3174), .Y(new_n5103));
  nor_5  g02755(.A(new_n5103), .B(new_n5102), .Y(new_n5104));
  not_8  g02756(.A(new_n5086), .Y(new_n5105));
  nand_5 g02757(.A(new_n5105), .B(new_n3174), .Y(new_n5106));
  nand_5 g02758(.A(new_n5106), .B(new_n5089), .Y(new_n5107));
  or_6   g02759(.A(new_n5107), .B(new_n5104), .Y(new_n5108));
  nand_5 g02760(.A(new_n5108), .B(new_n5097), .Y(new_n5109));
  nand_5 g02761(.A(new_n5109), .B(new_n5096), .Y(new_n5110));
  nand_5 g02762(.A(new_n5110), .B(new_n5094), .Y(new_n5111));
  xnor_4 g02763(.A(new_n5110), .B(new_n5094), .Y(new_n5112));
  or_6   g02764(.A(new_n5112), .B(new_n3164), .Y(new_n5113));
  nand_5 g02765(.A(new_n5113), .B(new_n5111), .Y(new_n5114));
  nand_5 g02766(.A(pi191), .B(pi102), .Y(new_n5115));
  not_8  g02767(.A(new_n5115), .Y(new_n5116));
  not_8  g02768(.A(new_n5082), .Y(new_n5117));
  nor_5  g02769(.A(new_n5093), .B(new_n5117), .Y(new_n5118));
  nor_5  g02770(.A(new_n5118), .B(new_n5116), .Y(new_n5119));
  not_8  g02771(.A(new_n5119), .Y(new_n5120));
  nand_5 g02772(.A(pi498), .B(pi316), .Y(new_n5121));
  nand_5 g02773(.A(new_n4667), .B(new_n2474), .Y(new_n5122));
  nand_5 g02774(.A(new_n5122), .B(new_n5121), .Y(new_n5123));
  xor_4  g02775(.A(new_n5123), .B(new_n5120), .Y(new_n5124));
  xor_4  g02776(.A(new_n5124), .B(new_n5114), .Y(new_n5125));
  xor_4  g02777(.A(new_n5125), .B(new_n3184), .Y(new_n5126));
  xor_4  g02778(.A(pi653), .B(new_n3542), .Y(new_n5127));
  not_8  g02779(.A(pi548), .Y(new_n5128));
  nand_5 g02780(.A(new_n5128), .B(pi421), .Y(new_n5129));
  xor_4  g02781(.A(pi548), .B(new_n3545), .Y(new_n5130));
  not_8  g02782(.A(pi127), .Y(new_n5131));
  nand_5 g02783(.A(pi626), .B(new_n5131), .Y(new_n5132));
  xor_4  g02784(.A(pi626), .B(new_n5131), .Y(new_n5133));
  nand_5 g02785(.A(new_n5046), .B(pi045), .Y(new_n5134));
  xor_4  g02786(.A(pi733), .B(new_n3554), .Y(new_n5135));
  nand_5 g02787(.A(new_n5043), .B(pi520), .Y(new_n5136));
  not_8  g02788(.A(new_n5136), .Y(new_n5137));
  nand_5 g02789(.A(new_n5137), .B(new_n5135), .Y(new_n5138));
  nand_5 g02790(.A(new_n5138), .B(new_n5134), .Y(new_n5139));
  nand_5 g02791(.A(new_n5139), .B(new_n5133), .Y(new_n5140));
  nand_5 g02792(.A(new_n5140), .B(new_n5132), .Y(new_n5141));
  nand_5 g02793(.A(new_n5141), .B(new_n5130), .Y(new_n5142));
  nand_5 g02794(.A(new_n5142), .B(new_n5129), .Y(new_n5143));
  xor_4  g02795(.A(new_n5143), .B(new_n5127), .Y(new_n5144));
  nand_5 g02796(.A(new_n5144), .B(new_n5126), .Y(new_n5145));
  xnor_4 g02797(.A(new_n5144), .B(new_n5126), .Y(new_n5146));
  xor_4  g02798(.A(new_n5112), .B(new_n3163), .Y(new_n5147));
  xor_4  g02799(.A(new_n5141), .B(new_n5130), .Y(new_n5148));
  or_6   g02800(.A(new_n5148), .B(new_n5147), .Y(new_n5149));
  xor_4  g02801(.A(new_n5148), .B(new_n5147), .Y(new_n5150));
  nand_5 g02802(.A(new_n5097), .B(new_n5096), .Y(new_n5151));
  xor_4  g02803(.A(new_n5151), .B(new_n5108), .Y(new_n5152));
  xor_4  g02804(.A(new_n5139), .B(new_n5133), .Y(new_n5153));
  and_6  g02805(.A(new_n5153), .B(new_n5152), .Y(new_n5154));
  nor_5  g02806(.A(new_n5153), .B(new_n5152), .Y(new_n5155));
  not_8  g02807(.A(new_n5138), .Y(new_n5156));
  xor_4  g02808(.A(new_n5099), .B(new_n3169), .Y(new_n5157));
  xor_4  g02809(.A(new_n5103), .B(new_n5101), .Y(new_n5158));
  nand_5 g02810(.A(new_n5158), .B(new_n5157), .Y(new_n5159));
  nand_5 g02811(.A(new_n5159), .B(new_n5156), .Y(new_n5160));
  not_8  g02812(.A(new_n5157), .Y(new_n5161));
  nor_5  g02813(.A(new_n5043), .B(pi520), .Y(new_n5162));
  nand_5 g02814(.A(new_n5162), .B(new_n5161), .Y(new_n5163));
  nor_5  g02815(.A(new_n5163), .B(new_n5135), .Y(new_n5164));
  nand_5 g02816(.A(new_n5157), .B(new_n5137), .Y(new_n5165));
  nand_5 g02817(.A(new_n5165), .B(new_n5163), .Y(new_n5166));
  xor_4  g02818(.A(new_n5166), .B(new_n5135), .Y(new_n5167));
  nor_5  g02819(.A(new_n5167), .B(new_n5158), .Y(new_n5168));
  nor_5  g02820(.A(new_n5168), .B(new_n5164), .Y(new_n5169));
  nand_5 g02821(.A(new_n5169), .B(new_n5160), .Y(new_n5170));
  nor_5  g02822(.A(new_n5170), .B(new_n5155), .Y(new_n5171));
  nor_5  g02823(.A(new_n5171), .B(new_n5154), .Y(new_n5172));
  nand_5 g02824(.A(new_n5172), .B(new_n5150), .Y(new_n5173));
  nand_5 g02825(.A(new_n5173), .B(new_n5149), .Y(new_n5174));
  or_6   g02826(.A(new_n5174), .B(new_n5146), .Y(new_n5175));
  nand_5 g02827(.A(new_n5175), .B(new_n5145), .Y(new_n5176));
  nand_5 g02828(.A(new_n5122), .B(new_n5120), .Y(new_n5177));
  nand_5 g02829(.A(new_n5177), .B(new_n5121), .Y(new_n5178));
  not_8  g02830(.A(new_n5178), .Y(new_n5179));
  nand_5 g02831(.A(pi790), .B(pi630), .Y(new_n5180));
  not_8  g02832(.A(pi790), .Y(new_n5181));
  nand_5 g02833(.A(new_n5181), .B(new_n4709), .Y(new_n5182));
  and_6  g02834(.A(new_n5182), .B(new_n5180), .Y(new_n5183));
  xor_4  g02835(.A(new_n5183), .B(new_n5179), .Y(new_n5184));
  xor_4  g02836(.A(new_n5184), .B(new_n3162), .Y(new_n5185));
  nand_5 g02837(.A(new_n5124), .B(new_n5114), .Y(new_n5186));
  not_8  g02838(.A(new_n5125), .Y(new_n5187));
  or_6   g02839(.A(new_n5187), .B(new_n3184), .Y(new_n5188));
  nand_5 g02840(.A(new_n5188), .B(new_n5186), .Y(new_n5189));
  xor_4  g02841(.A(new_n5189), .B(new_n5185), .Y(new_n5190));
  not_8  g02842(.A(new_n5190), .Y(new_n5191));
  not_8  g02843(.A(pi653), .Y(new_n5192));
  nand_5 g02844(.A(new_n5192), .B(pi453), .Y(new_n5193));
  nand_5 g02845(.A(new_n5143), .B(new_n5127), .Y(new_n5194));
  nand_5 g02846(.A(new_n5194), .B(new_n5193), .Y(new_n5195));
  not_8  g02847(.A(pi174), .Y(new_n5196));
  nand_5 g02848(.A(new_n5196), .B(pi138), .Y(new_n5197));
  nand_5 g02849(.A(pi174), .B(new_n3539), .Y(new_n5198));
  nand_5 g02850(.A(new_n5198), .B(new_n5197), .Y(new_n5199));
  xnor_4 g02851(.A(new_n5199), .B(new_n5195), .Y(new_n5200));
  xor_4  g02852(.A(new_n5200), .B(new_n5191), .Y(new_n5201));
  xnor_4 g02853(.A(new_n5201), .B(new_n5176), .Y(po0015));
  xor_4  g02854(.A(pi208), .B(new_n3212), .Y(new_n5203));
  nand_5 g02855(.A(new_n3155), .B(pi105), .Y(new_n5204));
  not_8  g02856(.A(pi105), .Y(new_n5205));
  xor_4  g02857(.A(pi802), .B(new_n5205), .Y(new_n5206));
  nand_5 g02858(.A(new_n3157), .B(pi175), .Y(new_n5207));
  xor_4  g02859(.A(pi601), .B(new_n3218), .Y(new_n5208));
  nand_5 g02860(.A(pi792), .B(new_n3191), .Y(new_n5209));
  xor_4  g02861(.A(pi792), .B(new_n3191), .Y(new_n5210));
  nand_5 g02862(.A(pi649), .B(new_n3186), .Y(new_n5211));
  xor_4  g02863(.A(pi649), .B(new_n3186), .Y(new_n5212));
  nand_5 g02864(.A(pi563), .B(new_n3282), .Y(new_n5213));
  xor_4  g02865(.A(pi563), .B(new_n3282), .Y(new_n5214));
  or_6   g02866(.A(pi652), .B(new_n3234), .Y(new_n5215));
  xor_4  g02867(.A(pi652), .B(new_n3234), .Y(new_n5216));
  nand_5 g02868(.A(new_n3168), .B(pi633), .Y(new_n5217));
  nand_5 g02869(.A(pi776), .B(new_n3238), .Y(new_n5218));
  nand_5 g02870(.A(new_n5218), .B(pi718), .Y(new_n5219));
  nand_5 g02871(.A(new_n5219), .B(new_n5217), .Y(new_n5220));
  nand_5 g02872(.A(new_n5220), .B(new_n5216), .Y(new_n5221));
  nand_5 g02873(.A(new_n5221), .B(new_n5215), .Y(new_n5222));
  nand_5 g02874(.A(new_n5222), .B(new_n5214), .Y(new_n5223));
  nand_5 g02875(.A(new_n5223), .B(new_n5213), .Y(new_n5224));
  nand_5 g02876(.A(new_n5224), .B(new_n5212), .Y(new_n5225));
  nand_5 g02877(.A(new_n5225), .B(new_n5211), .Y(new_n5226));
  nand_5 g02878(.A(new_n5226), .B(new_n5210), .Y(new_n5227));
  nand_5 g02879(.A(new_n5227), .B(new_n5209), .Y(new_n5228));
  nand_5 g02880(.A(new_n5228), .B(new_n5208), .Y(new_n5229));
  nand_5 g02881(.A(new_n5229), .B(new_n5207), .Y(new_n5230));
  nand_5 g02882(.A(new_n5230), .B(new_n5206), .Y(new_n5231));
  nand_5 g02883(.A(new_n5231), .B(new_n5204), .Y(new_n5232));
  xnor_4 g02884(.A(new_n5232), .B(new_n5203), .Y(new_n5233));
  xor_4  g02885(.A(pi687), .B(pi325), .Y(new_n5234));
  nand_5 g02886(.A(pi637), .B(pi047), .Y(new_n5235));
  xor_4  g02887(.A(pi637), .B(pi047), .Y(new_n5236));
  nand_5 g02888(.A(pi410), .B(pi253), .Y(new_n5237));
  xor_4  g02889(.A(pi410), .B(pi253), .Y(new_n5238));
  nand_5 g02890(.A(pi829), .B(pi061), .Y(new_n5239));
  xor_4  g02891(.A(pi829), .B(pi061), .Y(new_n5240));
  nand_5 g02892(.A(pi172), .B(pi153), .Y(new_n5241));
  nand_5 g02893(.A(pi749), .B(pi151), .Y(new_n5242));
  not_8  g02894(.A(new_n5242), .Y(new_n5243));
  xor_4  g02895(.A(pi749), .B(pi151), .Y(new_n5244));
  not_8  g02896(.A(new_n5244), .Y(new_n5245));
  not_8  g02897(.A(pi570), .Y(new_n5246));
  nor_5  g02898(.A(new_n2389), .B(new_n5246), .Y(new_n5247));
  nor_5  g02899(.A(new_n2872), .B(new_n2391), .Y(new_n5248));
  xor_4  g02900(.A(pi144), .B(pi132), .Y(new_n5249));
  not_8  g02901(.A(new_n5249), .Y(new_n5250));
  nand_5 g02902(.A(pi390), .B(pi181), .Y(new_n5251));
  nor_5  g02903(.A(new_n5251), .B(new_n5250), .Y(new_n5252));
  nor_5  g02904(.A(new_n5252), .B(new_n5248), .Y(new_n5253));
  xor_4  g02905(.A(pi755), .B(new_n5246), .Y(new_n5254));
  nor_5  g02906(.A(new_n5254), .B(new_n5253), .Y(new_n5255));
  nor_5  g02907(.A(new_n5255), .B(new_n5247), .Y(new_n5256));
  nor_5  g02908(.A(new_n5256), .B(new_n5245), .Y(new_n5257));
  nor_5  g02909(.A(new_n5257), .B(new_n5243), .Y(new_n5258));
  not_8  g02910(.A(pi153), .Y(new_n5259));
  xor_4  g02911(.A(pi172), .B(new_n5259), .Y(new_n5260));
  or_6   g02912(.A(new_n5260), .B(new_n5258), .Y(new_n5261));
  nand_5 g02913(.A(new_n5261), .B(new_n5241), .Y(new_n5262));
  nand_5 g02914(.A(new_n5262), .B(new_n5240), .Y(new_n5263));
  nand_5 g02915(.A(new_n5263), .B(new_n5239), .Y(new_n5264));
  nand_5 g02916(.A(new_n5264), .B(new_n5238), .Y(new_n5265));
  nand_5 g02917(.A(new_n5265), .B(new_n5237), .Y(new_n5266));
  nand_5 g02918(.A(new_n5266), .B(new_n5236), .Y(new_n5267));
  nand_5 g02919(.A(new_n5267), .B(new_n5235), .Y(new_n5268));
  xor_4  g02920(.A(new_n5268), .B(new_n5234), .Y(new_n5269));
  not_8  g02921(.A(new_n5269), .Y(new_n5270));
  xor_4  g02922(.A(pi349), .B(pi189), .Y(new_n5271));
  not_8  g02923(.A(pi424), .Y(new_n5272));
  nand_5 g02924(.A(new_n5272), .B(new_n2897), .Y(new_n5273));
  xor_4  g02925(.A(pi424), .B(pi239), .Y(new_n5274));
  not_8  g02926(.A(pi018), .Y(new_n5275));
  nand_5 g02927(.A(new_n2932), .B(new_n5275), .Y(new_n5276));
  nand_5 g02928(.A(pi229), .B(pi217), .Y(new_n5277));
  not_8  g02929(.A(new_n5277), .Y(new_n5278));
  nand_5 g02930(.A(pi406), .B(pi107), .Y(new_n5279));
  not_8  g02931(.A(new_n5279), .Y(new_n5280));
  xor_4  g02932(.A(pi406), .B(pi107), .Y(new_n5281));
  not_8  g02933(.A(new_n5281), .Y(new_n5282));
  not_8  g02934(.A(pi629), .Y(new_n5283));
  nand_5 g02935(.A(new_n5283), .B(new_n2912), .Y(new_n5284));
  xor_4  g02936(.A(pi629), .B(pi023), .Y(new_n5285));
  not_8  g02937(.A(pi076), .Y(new_n5286));
  not_8  g02938(.A(pi801), .Y(new_n5287));
  nor_5  g02939(.A(new_n5287), .B(new_n5286), .Y(new_n5288));
  xor_4  g02940(.A(pi801), .B(pi076), .Y(new_n5289));
  not_8  g02941(.A(new_n5289), .Y(new_n5290));
  nand_5 g02942(.A(pi500), .B(pi038), .Y(new_n5291));
  nand_5 g02943(.A(pi354), .B(pi044), .Y(new_n5292));
  nand_5 g02944(.A(new_n5292), .B(new_n5291), .Y(new_n5293));
  nand_5 g02945(.A(new_n3124), .B(new_n2920), .Y(new_n5294));
  nand_5 g02946(.A(new_n5294), .B(new_n5293), .Y(new_n5295));
  nor_5  g02947(.A(new_n5295), .B(new_n5290), .Y(new_n5296));
  nor_5  g02948(.A(new_n5296), .B(new_n5288), .Y(new_n5297));
  nand_5 g02949(.A(new_n5297), .B(new_n5285), .Y(new_n5298));
  nand_5 g02950(.A(new_n5298), .B(new_n5284), .Y(new_n5299));
  nor_5  g02951(.A(new_n5299), .B(new_n5282), .Y(new_n5300));
  nor_5  g02952(.A(new_n5300), .B(new_n5280), .Y(new_n5301));
  xor_4  g02953(.A(pi229), .B(pi217), .Y(new_n5302));
  not_8  g02954(.A(new_n5302), .Y(new_n5303));
  nor_5  g02955(.A(new_n5303), .B(new_n5301), .Y(new_n5304));
  nor_5  g02956(.A(new_n5304), .B(new_n5278), .Y(new_n5305));
  xor_4  g02957(.A(pi632), .B(new_n5275), .Y(new_n5306));
  not_8  g02958(.A(new_n5306), .Y(new_n5307));
  nand_5 g02959(.A(new_n5307), .B(new_n5305), .Y(new_n5308));
  nand_5 g02960(.A(new_n5308), .B(new_n5276), .Y(new_n5309));
  nand_5 g02961(.A(new_n5309), .B(new_n5274), .Y(new_n5310));
  nand_5 g02962(.A(new_n5310), .B(new_n5273), .Y(new_n5311));
  xnor_4 g02963(.A(new_n5311), .B(new_n5271), .Y(new_n5312));
  or_6   g02964(.A(new_n5312), .B(new_n5270), .Y(new_n5313));
  nand_5 g02965(.A(new_n5312), .B(new_n5270), .Y(new_n5314));
  nand_5 g02966(.A(new_n5314), .B(new_n5313), .Y(new_n5315));
  xor_4  g02967(.A(new_n5309), .B(new_n5274), .Y(new_n5316));
  not_8  g02968(.A(new_n5316), .Y(new_n5317));
  xnor_4 g02969(.A(new_n5266), .B(new_n5236), .Y(new_n5318));
  nor_5  g02970(.A(new_n5318), .B(new_n5317), .Y(new_n5319));
  xor_4  g02971(.A(new_n5262), .B(new_n5240), .Y(new_n5320));
  xor_4  g02972(.A(new_n5302), .B(new_n5301), .Y(new_n5321));
  nand_5 g02973(.A(new_n5321), .B(new_n5320), .Y(new_n5322));
  xor_4  g02974(.A(new_n5321), .B(new_n5320), .Y(new_n5323));
  not_8  g02975(.A(new_n5323), .Y(new_n5324));
  xor_4  g02976(.A(new_n5260), .B(new_n5258), .Y(new_n5325));
  xor_4  g02977(.A(new_n5299), .B(new_n5281), .Y(new_n5326));
  or_6   g02978(.A(new_n5326), .B(new_n5325), .Y(new_n5327));
  nand_5 g02979(.A(new_n5326), .B(new_n5325), .Y(new_n5328));
  xor_4  g02980(.A(new_n5297), .B(new_n5285), .Y(new_n5329));
  not_8  g02981(.A(new_n5329), .Y(new_n5330));
  xor_4  g02982(.A(new_n5256), .B(new_n5244), .Y(new_n5331));
  nor_5  g02983(.A(new_n5331), .B(new_n5330), .Y(new_n5332));
  xor_4  g02984(.A(new_n5331), .B(new_n5330), .Y(new_n5333));
  not_8  g02985(.A(new_n5333), .Y(new_n5334));
  xor_4  g02986(.A(new_n5254), .B(new_n5253), .Y(new_n5335));
  xor_4  g02987(.A(new_n5295), .B(new_n5289), .Y(new_n5336));
  or_6   g02988(.A(new_n5336), .B(new_n5335), .Y(new_n5337));
  xor_4  g02989(.A(new_n5336), .B(new_n5335), .Y(new_n5338));
  nor_5  g02990(.A(new_n2874), .B(pi038), .Y(new_n5339));
  not_8  g02991(.A(pi038), .Y(new_n5340));
  nor_5  g02992(.A(pi181), .B(new_n5340), .Y(new_n5341));
  nor_5  g02993(.A(new_n5341), .B(new_n5339), .Y(new_n5342));
  or_6   g02994(.A(pi500), .B(new_n2429), .Y(new_n5343));
  nand_5 g02995(.A(pi500), .B(new_n2429), .Y(new_n5344));
  nand_5 g02996(.A(new_n5344), .B(new_n5343), .Y(new_n5345));
  not_8  g02997(.A(new_n5345), .Y(new_n5346));
  xor_4  g02998(.A(new_n5346), .B(new_n5342), .Y(new_n5347));
  not_8  g02999(.A(new_n5347), .Y(new_n5348));
  nand_5 g03000(.A(new_n5348), .B(new_n5251), .Y(new_n5349));
  nand_5 g03001(.A(pi354), .B(new_n2391), .Y(new_n5350));
  nand_5 g03002(.A(new_n3124), .B(pi132), .Y(new_n5351));
  nand_5 g03003(.A(new_n5351), .B(new_n5350), .Y(new_n5352));
  not_8  g03004(.A(new_n5352), .Y(new_n5353));
  xor_4  g03005(.A(pi144), .B(new_n2920), .Y(new_n5354));
  not_8  g03006(.A(new_n5354), .Y(new_n5355));
  nand_5 g03007(.A(new_n2429), .B(new_n2874), .Y(new_n5356));
  nand_5 g03008(.A(new_n5356), .B(new_n5349), .Y(new_n5357));
  and_6  g03009(.A(new_n5357), .B(new_n5291), .Y(new_n5358));
  not_8  g03010(.A(new_n5356), .Y(new_n5359));
  nor_5  g03011(.A(new_n5359), .B(new_n5291), .Y(new_n5360));
  nor_5  g03012(.A(new_n5360), .B(new_n5358), .Y(new_n5361));
  xor_4  g03013(.A(new_n5361), .B(new_n5355), .Y(new_n5362));
  xor_4  g03014(.A(new_n5362), .B(new_n5353), .Y(new_n5363));
  not_8  g03015(.A(new_n5363), .Y(new_n5364));
  nand_5 g03016(.A(new_n5364), .B(new_n5349), .Y(new_n5365));
  nand_5 g03017(.A(new_n5365), .B(new_n5250), .Y(new_n5366));
  nor_5  g03018(.A(new_n5359), .B(new_n5348), .Y(new_n5367));
  nor_5  g03019(.A(new_n5367), .B(new_n5364), .Y(new_n5368));
  nand_5 g03020(.A(new_n5359), .B(new_n5250), .Y(new_n5369));
  not_8  g03021(.A(new_n5369), .Y(new_n5370));
  nor_5  g03022(.A(new_n5370), .B(new_n5252), .Y(new_n5371));
  not_8  g03023(.A(new_n5371), .Y(new_n5372));
  nor_5  g03024(.A(new_n5372), .B(new_n5368), .Y(new_n5373));
  nand_5 g03025(.A(new_n5373), .B(new_n5366), .Y(new_n5374));
  nand_5 g03026(.A(new_n5374), .B(new_n5338), .Y(new_n5375));
  nand_5 g03027(.A(new_n5375), .B(new_n5337), .Y(new_n5376));
  nor_5  g03028(.A(new_n5376), .B(new_n5334), .Y(new_n5377));
  nor_5  g03029(.A(new_n5377), .B(new_n5332), .Y(new_n5378));
  nand_5 g03030(.A(new_n5378), .B(new_n5328), .Y(new_n5379));
  nand_5 g03031(.A(new_n5379), .B(new_n5327), .Y(new_n5380));
  or_6   g03032(.A(new_n5380), .B(new_n5324), .Y(new_n5381));
  nand_5 g03033(.A(new_n5381), .B(new_n5322), .Y(new_n5382));
  xor_4  g03034(.A(new_n5264), .B(new_n5238), .Y(new_n5383));
  xor_4  g03035(.A(new_n5307), .B(new_n5305), .Y(new_n5384));
  and_6  g03036(.A(new_n5384), .B(new_n5383), .Y(new_n5385));
  nor_5  g03037(.A(new_n5385), .B(new_n5382), .Y(new_n5386));
  nor_5  g03038(.A(new_n5384), .B(new_n5383), .Y(new_n5387));
  or_6   g03039(.A(new_n5387), .B(new_n5386), .Y(new_n5388));
  xor_4  g03040(.A(new_n5318), .B(new_n5317), .Y(new_n5389));
  not_8  g03041(.A(new_n5389), .Y(new_n5390));
  nor_5  g03042(.A(new_n5390), .B(new_n5388), .Y(new_n5391));
  nor_5  g03043(.A(new_n5391), .B(new_n5319), .Y(new_n5392));
  xor_4  g03044(.A(new_n5392), .B(new_n5315), .Y(new_n5393));
  xor_4  g03045(.A(new_n5393), .B(new_n5233), .Y(new_n5394));
  xnor_4 g03046(.A(new_n5230), .B(new_n5206), .Y(new_n5395));
  xor_4  g03047(.A(new_n5389), .B(new_n5388), .Y(new_n5396));
  nor_5  g03048(.A(new_n5396), .B(new_n5395), .Y(new_n5397));
  xnor_4 g03049(.A(new_n5228), .B(new_n5208), .Y(new_n5398));
  xnor_4 g03050(.A(new_n5226), .B(new_n5210), .Y(new_n5399));
  xnor_4 g03051(.A(new_n5224), .B(new_n5212), .Y(new_n5400));
  xnor_4 g03052(.A(new_n5222), .B(new_n5214), .Y(new_n5401));
  xor_4  g03053(.A(new_n5376), .B(new_n5333), .Y(new_n5402));
  or_6   g03054(.A(new_n5402), .B(new_n5401), .Y(new_n5403));
  not_8  g03055(.A(new_n5402), .Y(new_n5404));
  xor_4  g03056(.A(new_n5404), .B(new_n5401), .Y(new_n5405));
  and_6  g03057(.A(new_n5217), .B(new_n5218), .Y(new_n5406));
  nand_5 g03058(.A(new_n3340), .B(pi364), .Y(new_n5407));
  or_6   g03059(.A(new_n5407), .B(new_n5348), .Y(new_n5408));
  or_6   g03060(.A(new_n5408), .B(new_n5406), .Y(new_n5409));
  nor_5  g03061(.A(new_n3340), .B(pi364), .Y(new_n5410));
  nand_5 g03062(.A(new_n5410), .B(new_n5348), .Y(new_n5411));
  nand_5 g03063(.A(new_n5411), .B(new_n5408), .Y(new_n5412));
  xor_4  g03064(.A(new_n5412), .B(new_n5406), .Y(new_n5413));
  or_6   g03065(.A(new_n5413), .B(new_n5364), .Y(new_n5414));
  nand_5 g03066(.A(new_n5411), .B(pi718), .Y(new_n5415));
  nand_5 g03067(.A(new_n5415), .B(new_n5413), .Y(new_n5416));
  nand_5 g03068(.A(new_n5416), .B(new_n5414), .Y(new_n5417));
  nand_5 g03069(.A(new_n5417), .B(new_n5409), .Y(new_n5418));
  xnor_4 g03070(.A(new_n5220), .B(new_n5216), .Y(new_n5419));
  nand_5 g03071(.A(new_n5419), .B(new_n5418), .Y(new_n5420));
  xor_4  g03072(.A(new_n5374), .B(new_n5338), .Y(new_n5421));
  xor_4  g03073(.A(new_n5419), .B(new_n5418), .Y(new_n5422));
  nand_5 g03074(.A(new_n5422), .B(new_n5421), .Y(new_n5423));
  nand_5 g03075(.A(new_n5423), .B(new_n5420), .Y(new_n5424));
  or_6   g03076(.A(new_n5424), .B(new_n5405), .Y(new_n5425));
  nand_5 g03077(.A(new_n5425), .B(new_n5403), .Y(new_n5426));
  not_8  g03078(.A(new_n5426), .Y(new_n5427));
  nand_5 g03079(.A(new_n5427), .B(new_n5400), .Y(new_n5428));
  xor_4  g03080(.A(new_n5426), .B(new_n5400), .Y(new_n5429));
  nand_5 g03081(.A(new_n5328), .B(new_n5327), .Y(new_n5430));
  xor_4  g03082(.A(new_n5430), .B(new_n5378), .Y(new_n5431));
  or_6   g03083(.A(new_n5431), .B(new_n5429), .Y(new_n5432));
  nand_5 g03084(.A(new_n5432), .B(new_n5428), .Y(new_n5433));
  nand_5 g03085(.A(new_n5433), .B(new_n5399), .Y(new_n5434));
  xor_4  g03086(.A(new_n5380), .B(new_n5324), .Y(new_n5435));
  not_8  g03087(.A(new_n5435), .Y(new_n5436));
  xor_4  g03088(.A(new_n5433), .B(new_n5399), .Y(new_n5437));
  nand_5 g03089(.A(new_n5437), .B(new_n5436), .Y(new_n5438));
  nand_5 g03090(.A(new_n5438), .B(new_n5434), .Y(new_n5439));
  nand_5 g03091(.A(new_n5439), .B(new_n5398), .Y(new_n5440));
  xor_4  g03092(.A(new_n5439), .B(new_n5398), .Y(new_n5441));
  nor_5  g03093(.A(new_n5387), .B(new_n5385), .Y(new_n5442));
  xor_4  g03094(.A(new_n5442), .B(new_n5382), .Y(new_n5443));
  not_8  g03095(.A(new_n5443), .Y(new_n5444));
  nand_5 g03096(.A(new_n5444), .B(new_n5441), .Y(new_n5445));
  nand_5 g03097(.A(new_n5445), .B(new_n5440), .Y(new_n5446));
  xnor_4 g03098(.A(new_n5396), .B(new_n5395), .Y(new_n5447));
  nor_5  g03099(.A(new_n5447), .B(new_n5446), .Y(new_n5448));
  nor_5  g03100(.A(new_n5448), .B(new_n5397), .Y(new_n5449));
  xnor_4 g03101(.A(new_n5449), .B(new_n5394), .Y(po0016));
  not_8  g03102(.A(pi430), .Y(new_n5451));
  nand_5 g03103(.A(pi565), .B(new_n5451), .Y(new_n5452));
  xor_4  g03104(.A(pi565), .B(new_n5451), .Y(new_n5453));
  not_8  g03105(.A(pi777), .Y(new_n5454));
  nand_5 g03106(.A(pi784), .B(new_n5454), .Y(new_n5455));
  xor_4  g03107(.A(pi784), .B(new_n5454), .Y(new_n5456));
  not_8  g03108(.A(pi319), .Y(new_n5457));
  nand_5 g03109(.A(pi734), .B(new_n5457), .Y(new_n5458));
  nand_5 g03110(.A(new_n4262), .B(pi319), .Y(new_n5459));
  not_8  g03111(.A(pi429), .Y(new_n5460));
  nand_5 g03112(.A(new_n5460), .B(pi395), .Y(new_n5461));
  xor_4  g03113(.A(pi429), .B(new_n4266), .Y(new_n5462));
  not_8  g03114(.A(pi699), .Y(new_n5463));
  nand_5 g03115(.A(new_n5463), .B(pi351), .Y(new_n5464));
  xor_4  g03116(.A(pi699), .B(new_n4045), .Y(new_n5465));
  nand_5 g03117(.A(pi497), .B(new_n2405), .Y(new_n5466));
  xor_4  g03118(.A(pi497), .B(new_n2405), .Y(new_n5467));
  nand_5 g03119(.A(pi506), .B(new_n2385), .Y(new_n5468));
  xor_4  g03120(.A(pi506), .B(new_n2385), .Y(new_n5469));
  nand_5 g03121(.A(new_n2388), .B(pi374), .Y(new_n5470));
  not_8  g03122(.A(new_n5470), .Y(new_n5471));
  xor_4  g03123(.A(pi486), .B(new_n3900), .Y(new_n5472));
  not_8  g03124(.A(new_n5472), .Y(new_n5473));
  nand_5 g03125(.A(new_n3905), .B(pi611), .Y(new_n5474));
  nand_5 g03126(.A(pi688), .B(new_n2392), .Y(new_n5475));
  nand_5 g03127(.A(pi445), .B(new_n2428), .Y(new_n5476));
  nand_5 g03128(.A(new_n5476), .B(new_n5475), .Y(new_n5477));
  nand_5 g03129(.A(new_n5477), .B(new_n5474), .Y(new_n5478));
  nor_5  g03130(.A(new_n5478), .B(new_n5473), .Y(new_n5479));
  nor_5  g03131(.A(new_n5479), .B(new_n5471), .Y(new_n5480));
  not_8  g03132(.A(new_n5480), .Y(new_n5481));
  nand_5 g03133(.A(new_n5481), .B(new_n5469), .Y(new_n5482));
  nand_5 g03134(.A(new_n5482), .B(new_n5468), .Y(new_n5483));
  nand_5 g03135(.A(new_n5483), .B(new_n5467), .Y(new_n5484));
  nand_5 g03136(.A(new_n5484), .B(new_n5466), .Y(new_n5485));
  nand_5 g03137(.A(new_n5485), .B(new_n5465), .Y(new_n5486));
  nand_5 g03138(.A(new_n5486), .B(new_n5464), .Y(new_n5487));
  nand_5 g03139(.A(new_n5487), .B(new_n5462), .Y(new_n5488));
  nand_5 g03140(.A(new_n5488), .B(new_n5461), .Y(new_n5489));
  nand_5 g03141(.A(new_n5489), .B(new_n5459), .Y(new_n5490));
  nand_5 g03142(.A(new_n5490), .B(new_n5458), .Y(new_n5491));
  nand_5 g03143(.A(new_n5491), .B(new_n5456), .Y(new_n5492));
  nand_5 g03144(.A(new_n5492), .B(new_n5455), .Y(new_n5493));
  nand_5 g03145(.A(new_n5493), .B(new_n5453), .Y(new_n5494));
  nand_5 g03146(.A(new_n5494), .B(new_n5452), .Y(new_n5495));
  not_8  g03147(.A(new_n5495), .Y(new_n5496));
  not_8  g03148(.A(pi827), .Y(new_n5497));
  nand_5 g03149(.A(new_n5497), .B(pi334), .Y(new_n5498));
  not_8  g03150(.A(pi737), .Y(new_n5499));
  nand_5 g03151(.A(new_n5499), .B(pi342), .Y(new_n5500));
  not_8  g03152(.A(pi342), .Y(new_n5501));
  xor_4  g03153(.A(pi737), .B(new_n5501), .Y(new_n5502));
  not_8  g03154(.A(pi692), .Y(new_n5503));
  nand_5 g03155(.A(new_n5503), .B(pi549), .Y(new_n5504));
  not_8  g03156(.A(pi549), .Y(new_n5505));
  xor_4  g03157(.A(pi692), .B(new_n5505), .Y(new_n5506));
  not_8  g03158(.A(pi625), .Y(new_n5507));
  nand_5 g03159(.A(new_n5507), .B(pi373), .Y(new_n5508));
  not_8  g03160(.A(pi373), .Y(new_n5509));
  xor_4  g03161(.A(pi625), .B(new_n5509), .Y(new_n5510));
  not_8  g03162(.A(pi128), .Y(new_n5511));
  nand_5 g03163(.A(pi492), .B(new_n5511), .Y(new_n5512));
  not_8  g03164(.A(pi739), .Y(new_n5513));
  nand_5 g03165(.A(new_n5513), .B(pi200), .Y(new_n5514));
  not_8  g03166(.A(pi200), .Y(new_n5515));
  xor_4  g03167(.A(pi739), .B(new_n5515), .Y(new_n5516));
  not_8  g03168(.A(pi067), .Y(new_n5517));
  nand_5 g03169(.A(pi836), .B(new_n5517), .Y(new_n5518));
  xor_4  g03170(.A(pi836), .B(new_n5517), .Y(new_n5519));
  not_8  g03171(.A(pi675), .Y(new_n5520));
  nand_5 g03172(.A(pi839), .B(new_n5520), .Y(new_n5521));
  not_8  g03173(.A(pi839), .Y(new_n5522));
  nand_5 g03174(.A(new_n5522), .B(pi675), .Y(new_n5523));
  nand_5 g03175(.A(new_n5523), .B(pi214), .Y(new_n5524));
  nand_5 g03176(.A(new_n5524), .B(new_n5521), .Y(new_n5525));
  nand_5 g03177(.A(new_n5525), .B(new_n5519), .Y(new_n5526));
  nand_5 g03178(.A(new_n5526), .B(new_n5518), .Y(new_n5527));
  nand_5 g03179(.A(new_n5527), .B(new_n5516), .Y(new_n5528));
  nand_5 g03180(.A(new_n5528), .B(new_n5514), .Y(new_n5529));
  xor_4  g03181(.A(pi492), .B(pi128), .Y(new_n5530));
  not_8  g03182(.A(new_n5530), .Y(new_n5531));
  nand_5 g03183(.A(new_n5531), .B(new_n5529), .Y(new_n5532));
  nand_5 g03184(.A(new_n5532), .B(new_n5512), .Y(new_n5533));
  nand_5 g03185(.A(new_n5533), .B(new_n5510), .Y(new_n5534));
  nand_5 g03186(.A(new_n5534), .B(new_n5508), .Y(new_n5535));
  nand_5 g03187(.A(new_n5535), .B(new_n5506), .Y(new_n5536));
  nand_5 g03188(.A(new_n5536), .B(new_n5504), .Y(new_n5537));
  nand_5 g03189(.A(new_n5537), .B(new_n5502), .Y(new_n5538));
  nand_5 g03190(.A(new_n5538), .B(new_n5500), .Y(new_n5539));
  xor_4  g03191(.A(pi827), .B(pi334), .Y(new_n5540));
  not_8  g03192(.A(new_n5540), .Y(new_n5541));
  nand_5 g03193(.A(new_n5541), .B(new_n5539), .Y(new_n5542));
  nand_5 g03194(.A(new_n5542), .B(new_n5498), .Y(new_n5543));
  nand_5 g03195(.A(pi405), .B(pi403), .Y(new_n5544));
  not_8  g03196(.A(pi403), .Y(new_n5545));
  not_8  g03197(.A(pi405), .Y(new_n5546));
  nand_5 g03198(.A(new_n5546), .B(new_n5545), .Y(new_n5547));
  nand_5 g03199(.A(new_n5547), .B(new_n5544), .Y(new_n5548));
  not_8  g03200(.A(new_n5548), .Y(new_n5549));
  or_6   g03201(.A(new_n5549), .B(new_n5543), .Y(new_n5550));
  nand_5 g03202(.A(new_n5543), .B(new_n5546), .Y(new_n5551));
  nand_5 g03203(.A(new_n5551), .B(new_n5545), .Y(new_n5552));
  nand_5 g03204(.A(new_n5552), .B(new_n5550), .Y(new_n5553));
  nand_5 g03205(.A(new_n5553), .B(new_n5496), .Y(new_n5554));
  xor_4  g03206(.A(new_n5493), .B(new_n5453), .Y(new_n5555));
  xor_4  g03207(.A(new_n5549), .B(new_n5543), .Y(new_n5556));
  or_6   g03208(.A(new_n5556), .B(new_n5555), .Y(new_n5557));
  xor_4  g03209(.A(new_n5556), .B(new_n5555), .Y(new_n5558));
  xor_4  g03210(.A(new_n5540), .B(new_n5539), .Y(new_n5559));
  xor_4  g03211(.A(new_n5491), .B(new_n5456), .Y(new_n5560));
  or_6   g03212(.A(new_n5560), .B(new_n5559), .Y(new_n5561));
  xor_4  g03213(.A(new_n5560), .B(new_n5559), .Y(new_n5562));
  xnor_4 g03214(.A(new_n5537), .B(new_n5502), .Y(new_n5563));
  and_6  g03215(.A(new_n5459), .B(new_n5458), .Y(new_n5564));
  xor_4  g03216(.A(new_n5564), .B(new_n5489), .Y(new_n5565));
  nor_5  g03217(.A(new_n5565), .B(new_n5563), .Y(new_n5566));
  xor_4  g03218(.A(new_n5565), .B(new_n5563), .Y(new_n5567));
  not_8  g03219(.A(new_n5567), .Y(new_n5568));
  xor_4  g03220(.A(new_n5487), .B(new_n5462), .Y(new_n5569));
  xnor_4 g03221(.A(new_n5535), .B(new_n5506), .Y(new_n5570));
  nor_5  g03222(.A(new_n5570), .B(new_n5569), .Y(new_n5571));
  xor_4  g03223(.A(new_n5570), .B(new_n5569), .Y(new_n5572));
  xor_4  g03224(.A(new_n5485), .B(new_n5465), .Y(new_n5573));
  xnor_4 g03225(.A(new_n5533), .B(new_n5510), .Y(new_n5574));
  or_6   g03226(.A(new_n5574), .B(new_n5573), .Y(new_n5575));
  xor_4  g03227(.A(new_n5574), .B(new_n5573), .Y(new_n5576));
  xor_4  g03228(.A(new_n5483), .B(new_n5467), .Y(new_n5577));
  xor_4  g03229(.A(new_n5530), .B(new_n5529), .Y(new_n5578));
  nand_5 g03230(.A(new_n5578), .B(new_n5577), .Y(new_n5579));
  xor_4  g03231(.A(new_n5578), .B(new_n5577), .Y(new_n5580));
  xnor_4 g03232(.A(new_n5527), .B(new_n5516), .Y(new_n5581));
  xor_4  g03233(.A(new_n5480), .B(new_n5469), .Y(new_n5582));
  not_8  g03234(.A(new_n5582), .Y(new_n5583));
  or_6   g03235(.A(new_n5583), .B(new_n5581), .Y(new_n5584));
  xor_4  g03236(.A(new_n5583), .B(new_n5581), .Y(new_n5585));
  not_8  g03237(.A(new_n5585), .Y(new_n5586));
  xor_4  g03238(.A(new_n5478), .B(new_n5472), .Y(new_n5587));
  not_8  g03239(.A(new_n5587), .Y(new_n5588));
  xnor_4 g03240(.A(new_n5525), .B(new_n5519), .Y(new_n5589));
  nand_5 g03241(.A(new_n5589), .B(new_n5588), .Y(new_n5590));
  or_6   g03242(.A(new_n5589), .B(new_n5588), .Y(new_n5591));
  nand_5 g03243(.A(new_n5521), .B(new_n5523), .Y(new_n5592));
  xor_4  g03244(.A(pi445), .B(new_n2428), .Y(new_n5593));
  not_8  g03245(.A(new_n5593), .Y(new_n5594));
  nand_5 g03246(.A(pi214), .B(pi010), .Y(new_n5595));
  not_8  g03247(.A(pi214), .Y(new_n5596));
  nand_5 g03248(.A(new_n5596), .B(new_n2555), .Y(new_n5597));
  nand_5 g03249(.A(new_n5597), .B(new_n5595), .Y(new_n5598));
  nor_5  g03250(.A(new_n5598), .B(new_n5594), .Y(new_n5599));
  nand_5 g03251(.A(new_n5599), .B(pi010), .Y(new_n5600));
  nor_5  g03252(.A(new_n5596), .B(pi010), .Y(new_n5601));
  nand_5 g03253(.A(new_n5601), .B(new_n5594), .Y(new_n5602));
  nand_5 g03254(.A(new_n5602), .B(new_n5600), .Y(new_n5603));
  xor_4  g03255(.A(new_n5603), .B(new_n5592), .Y(new_n5604));
  and_6  g03256(.A(new_n5475), .B(new_n5474), .Y(new_n5605));
  xor_4  g03257(.A(new_n5605), .B(new_n5476), .Y(new_n5606));
  not_8  g03258(.A(new_n5606), .Y(new_n5607));
  nand_5 g03259(.A(new_n5607), .B(new_n5604), .Y(new_n5608));
  nand_5 g03260(.A(new_n5595), .B(new_n5594), .Y(new_n5609));
  nand_5 g03261(.A(new_n5609), .B(new_n5597), .Y(new_n5610));
  or_6   g03262(.A(new_n5610), .B(new_n5604), .Y(new_n5611));
  nand_5 g03263(.A(new_n5611), .B(new_n5608), .Y(new_n5612));
  nand_5 g03264(.A(new_n5612), .B(new_n5591), .Y(new_n5613));
  nand_5 g03265(.A(new_n5613), .B(new_n5590), .Y(new_n5614));
  or_6   g03266(.A(new_n5614), .B(new_n5586), .Y(new_n5615));
  nand_5 g03267(.A(new_n5615), .B(new_n5584), .Y(new_n5616));
  not_8  g03268(.A(new_n5616), .Y(new_n5617));
  nand_5 g03269(.A(new_n5617), .B(new_n5580), .Y(new_n5618));
  nand_5 g03270(.A(new_n5618), .B(new_n5579), .Y(new_n5619));
  not_8  g03271(.A(new_n5619), .Y(new_n5620));
  nand_5 g03272(.A(new_n5620), .B(new_n5576), .Y(new_n5621));
  nand_5 g03273(.A(new_n5621), .B(new_n5575), .Y(new_n5622));
  and_6  g03274(.A(new_n5622), .B(new_n5572), .Y(new_n5623));
  nor_5  g03275(.A(new_n5623), .B(new_n5571), .Y(new_n5624));
  nor_5  g03276(.A(new_n5624), .B(new_n5568), .Y(new_n5625));
  or_6   g03277(.A(new_n5625), .B(new_n5566), .Y(new_n5626));
  nand_5 g03278(.A(new_n5626), .B(new_n5562), .Y(new_n5627));
  nand_5 g03279(.A(new_n5627), .B(new_n5561), .Y(new_n5628));
  nand_5 g03280(.A(new_n5628), .B(new_n5558), .Y(new_n5629));
  nand_5 g03281(.A(new_n5629), .B(new_n5557), .Y(new_n5630));
  xor_4  g03282(.A(new_n5553), .B(new_n5495), .Y(new_n5631));
  or_6   g03283(.A(new_n5631), .B(new_n5630), .Y(new_n5632));
  nand_5 g03284(.A(new_n5632), .B(new_n5554), .Y(new_n5633));
  not_8  g03285(.A(pi282), .Y(new_n5634));
  xor_4  g03286(.A(pi735), .B(new_n5634), .Y(new_n5635));
  not_8  g03287(.A(pi472), .Y(new_n5636));
  nand_5 g03288(.A(pi533), .B(new_n5636), .Y(new_n5637));
  xor_4  g03289(.A(pi533), .B(pi472), .Y(new_n5638));
  not_8  g03290(.A(new_n5638), .Y(new_n5639));
  not_8  g03291(.A(pi834), .Y(new_n5640));
  nand_5 g03292(.A(new_n5640), .B(pi377), .Y(new_n5641));
  not_8  g03293(.A(pi377), .Y(new_n5642));
  nand_5 g03294(.A(pi834), .B(new_n5642), .Y(new_n5643));
  not_8  g03295(.A(pi297), .Y(new_n5644));
  nand_5 g03296(.A(pi714), .B(new_n5644), .Y(new_n5645));
  not_8  g03297(.A(pi613), .Y(new_n5646));
  nand_5 g03298(.A(new_n5646), .B(pi539), .Y(new_n5647));
  not_8  g03299(.A(pi539), .Y(new_n5648));
  xor_4  g03300(.A(pi613), .B(new_n5648), .Y(new_n5649));
  nand_5 g03301(.A(new_n3991), .B(pi242), .Y(new_n5650));
  not_8  g03302(.A(pi242), .Y(new_n5651));
  xor_4  g03303(.A(pi250), .B(new_n5651), .Y(new_n5652));
  nand_5 g03304(.A(new_n3993), .B(pi252), .Y(new_n5653));
  not_8  g03305(.A(pi252), .Y(new_n5654));
  xor_4  g03306(.A(pi338), .B(new_n5654), .Y(new_n5655));
  nand_5 g03307(.A(pi391), .B(new_n3946), .Y(new_n5656));
  xor_4  g03308(.A(pi391), .B(new_n3946), .Y(new_n5657));
  nand_5 g03309(.A(pi638), .B(new_n3954), .Y(new_n5658));
  xor_4  g03310(.A(pi638), .B(new_n3954), .Y(new_n5659));
  nand_5 g03311(.A(new_n5659), .B(pi393), .Y(new_n5660));
  nand_5 g03312(.A(new_n5660), .B(new_n5658), .Y(new_n5661));
  nand_5 g03313(.A(new_n5661), .B(new_n5657), .Y(new_n5662));
  nand_5 g03314(.A(new_n5662), .B(new_n5656), .Y(new_n5663));
  nand_5 g03315(.A(new_n5663), .B(new_n5655), .Y(new_n5664));
  nand_5 g03316(.A(new_n5664), .B(new_n5653), .Y(new_n5665));
  nand_5 g03317(.A(new_n5665), .B(new_n5652), .Y(new_n5666));
  nand_5 g03318(.A(new_n5666), .B(new_n5650), .Y(new_n5667));
  nand_5 g03319(.A(new_n5667), .B(new_n5649), .Y(new_n5668));
  nand_5 g03320(.A(new_n5668), .B(new_n5647), .Y(new_n5669));
  xor_4  g03321(.A(pi714), .B(new_n5644), .Y(new_n5670));
  nand_5 g03322(.A(new_n5670), .B(new_n5669), .Y(new_n5671));
  nand_5 g03323(.A(new_n5671), .B(new_n5645), .Y(new_n5672));
  nand_5 g03324(.A(new_n5672), .B(new_n5643), .Y(new_n5673));
  nand_5 g03325(.A(new_n5673), .B(new_n5641), .Y(new_n5674));
  nand_5 g03326(.A(new_n5674), .B(new_n5639), .Y(new_n5675));
  nand_5 g03327(.A(new_n5675), .B(new_n5637), .Y(new_n5676));
  xor_4  g03328(.A(new_n5676), .B(new_n5635), .Y(new_n5677));
  xor_4  g03329(.A(new_n5674), .B(new_n5638), .Y(new_n5678));
  xnor_4 g03330(.A(new_n5626), .B(new_n5562), .Y(new_n5679));
  or_6   g03331(.A(new_n5679), .B(new_n5678), .Y(new_n5680));
  xor_4  g03332(.A(new_n5679), .B(new_n5678), .Y(new_n5681));
  xor_4  g03333(.A(new_n5624), .B(new_n5567), .Y(new_n5682));
  xor_4  g03334(.A(new_n5667), .B(new_n5649), .Y(new_n5683));
  xor_4  g03335(.A(new_n5665), .B(new_n5652), .Y(new_n5684));
  not_8  g03336(.A(new_n5684), .Y(new_n5685));
  xor_4  g03337(.A(new_n5663), .B(new_n5655), .Y(new_n5686));
  not_8  g03338(.A(new_n5686), .Y(new_n5687));
  xor_4  g03339(.A(new_n5661), .B(new_n5657), .Y(new_n5688));
  xor_4  g03340(.A(new_n5598), .B(new_n5594), .Y(new_n5689));
  nor_5  g03341(.A(pi393), .B(new_n2568), .Y(new_n5690));
  nand_5 g03342(.A(new_n5690), .B(new_n5689), .Y(new_n5691));
  not_8  g03343(.A(new_n5689), .Y(new_n5692));
  not_8  g03344(.A(pi393), .Y(new_n5693));
  nor_5  g03345(.A(new_n5693), .B(pi219), .Y(new_n5694));
  nand_5 g03346(.A(new_n5694), .B(new_n5692), .Y(new_n5695));
  nand_5 g03347(.A(new_n5695), .B(new_n5691), .Y(new_n5696));
  xor_4  g03348(.A(new_n5696), .B(new_n5659), .Y(new_n5697));
  xor_4  g03349(.A(new_n5607), .B(new_n5604), .Y(new_n5698));
  nor_5  g03350(.A(new_n5698), .B(new_n5697), .Y(new_n5699));
  nor_5  g03351(.A(new_n5696), .B(new_n5659), .Y(new_n5700));
  nand_5 g03352(.A(new_n5691), .B(new_n5660), .Y(new_n5701));
  nor_5  g03353(.A(new_n5701), .B(new_n5700), .Y(new_n5702));
  or_6   g03354(.A(new_n5702), .B(new_n5699), .Y(new_n5703));
  nor_5  g03355(.A(new_n5703), .B(new_n5688), .Y(new_n5704));
  xnor_4 g03356(.A(new_n5703), .B(new_n5688), .Y(new_n5705));
  nand_5 g03357(.A(new_n5591), .B(new_n5590), .Y(new_n5706));
  xor_4  g03358(.A(new_n5706), .B(new_n5612), .Y(new_n5707));
  nor_5  g03359(.A(new_n5707), .B(new_n5705), .Y(new_n5708));
  or_6   g03360(.A(new_n5708), .B(new_n5704), .Y(new_n5709));
  nand_5 g03361(.A(new_n5709), .B(new_n5687), .Y(new_n5710));
  xor_4  g03362(.A(new_n5709), .B(new_n5686), .Y(new_n5711));
  xor_4  g03363(.A(new_n5614), .B(new_n5585), .Y(new_n5712));
  not_8  g03364(.A(new_n5712), .Y(new_n5713));
  or_6   g03365(.A(new_n5713), .B(new_n5711), .Y(new_n5714));
  nand_5 g03366(.A(new_n5714), .B(new_n5710), .Y(new_n5715));
  or_6   g03367(.A(new_n5715), .B(new_n5685), .Y(new_n5716));
  xor_4  g03368(.A(new_n5715), .B(new_n5685), .Y(new_n5717));
  xor_4  g03369(.A(new_n5616), .B(new_n5580), .Y(new_n5718));
  nand_5 g03370(.A(new_n5718), .B(new_n5717), .Y(new_n5719));
  nand_5 g03371(.A(new_n5719), .B(new_n5716), .Y(new_n5720));
  nor_5  g03372(.A(new_n5720), .B(new_n5683), .Y(new_n5721));
  xnor_4 g03373(.A(new_n5720), .B(new_n5683), .Y(new_n5722));
  xor_4  g03374(.A(new_n5619), .B(new_n5576), .Y(new_n5723));
  not_8  g03375(.A(new_n5723), .Y(new_n5724));
  nor_5  g03376(.A(new_n5724), .B(new_n5722), .Y(new_n5725));
  or_6   g03377(.A(new_n5725), .B(new_n5721), .Y(new_n5726));
  not_8  g03378(.A(new_n5572), .Y(new_n5727));
  xor_4  g03379(.A(new_n5622), .B(new_n5727), .Y(new_n5728));
  nand_5 g03380(.A(new_n5728), .B(new_n5726), .Y(new_n5729));
  xnor_4 g03381(.A(new_n5728), .B(new_n5726), .Y(new_n5730));
  xor_4  g03382(.A(new_n5670), .B(new_n5669), .Y(new_n5731));
  or_6   g03383(.A(new_n5731), .B(new_n5730), .Y(new_n5732));
  nand_5 g03384(.A(new_n5732), .B(new_n5729), .Y(new_n5733));
  or_6   g03385(.A(new_n5733), .B(new_n5682), .Y(new_n5734));
  nand_5 g03386(.A(new_n5733), .B(new_n5682), .Y(new_n5735));
  nand_5 g03387(.A(new_n5643), .B(new_n5641), .Y(new_n5736));
  xnor_4 g03388(.A(new_n5736), .B(new_n5672), .Y(new_n5737));
  nand_5 g03389(.A(new_n5737), .B(new_n5735), .Y(new_n5738));
  nand_5 g03390(.A(new_n5738), .B(new_n5734), .Y(new_n5739));
  nand_5 g03391(.A(new_n5739), .B(new_n5681), .Y(new_n5740));
  nand_5 g03392(.A(new_n5740), .B(new_n5680), .Y(new_n5741));
  nor_5  g03393(.A(new_n5741), .B(new_n5677), .Y(new_n5742));
  xor_4  g03394(.A(new_n5628), .B(new_n5558), .Y(new_n5743));
  xnor_4 g03395(.A(new_n5741), .B(new_n5677), .Y(new_n5744));
  nor_5  g03396(.A(new_n5744), .B(new_n5743), .Y(new_n5745));
  or_6   g03397(.A(new_n5745), .B(new_n5742), .Y(new_n5746));
  nand_5 g03398(.A(pi735), .B(new_n5634), .Y(new_n5747));
  nand_5 g03399(.A(new_n5676), .B(new_n5635), .Y(new_n5748));
  nand_5 g03400(.A(new_n5748), .B(new_n5747), .Y(new_n5749));
  not_8  g03401(.A(new_n5749), .Y(new_n5750));
  nand_5 g03402(.A(new_n5750), .B(new_n5746), .Y(new_n5751));
  xor_4  g03403(.A(new_n5750), .B(new_n5746), .Y(new_n5752));
  xor_4  g03404(.A(new_n5631), .B(new_n5630), .Y(new_n5753));
  nand_5 g03405(.A(new_n5753), .B(new_n5752), .Y(new_n5754));
  nand_5 g03406(.A(new_n5754), .B(new_n5751), .Y(new_n5755));
  xnor_4 g03407(.A(new_n5755), .B(new_n5633), .Y(po0017));
  nand_5 g03408(.A(new_n2420), .B(pi062), .Y(new_n5757));
  not_8  g03409(.A(new_n5757), .Y(new_n5758));
  xor_4  g03410(.A(pi369), .B(new_n2956), .Y(new_n5759));
  xor_4  g03411(.A(new_n5759), .B(new_n5758), .Y(new_n5760));
  not_8  g03412(.A(new_n5760), .Y(new_n5761));
  xor_4  g03413(.A(pi438), .B(new_n3020), .Y(new_n5762));
  xor_4  g03414(.A(pi751), .B(new_n4405), .Y(new_n5763));
  nor_5  g03415(.A(new_n5763), .B(new_n5762), .Y(new_n5764));
  not_8  g03416(.A(pi751), .Y(new_n5765));
  nand_5 g03417(.A(new_n5765), .B(pi049), .Y(new_n5766));
  not_8  g03418(.A(new_n5766), .Y(new_n5767));
  not_8  g03419(.A(pi797), .Y(new_n5768));
  xor_4  g03420(.A(pi813), .B(new_n5768), .Y(new_n5769));
  xor_4  g03421(.A(new_n5769), .B(new_n5767), .Y(new_n5770));
  xor_4  g03422(.A(new_n5770), .B(new_n5764), .Y(new_n5771));
  xor_4  g03423(.A(new_n5771), .B(new_n5761), .Y(new_n5772));
  xor_4  g03424(.A(new_n5763), .B(new_n5762), .Y(new_n5773));
  and_6  g03425(.A(new_n5773), .B(new_n5594), .Y(new_n5774));
  xor_4  g03426(.A(new_n5774), .B(new_n5606), .Y(new_n5775));
  not_8  g03427(.A(new_n5775), .Y(new_n5776));
  xor_4  g03428(.A(new_n5776), .B(new_n5772), .Y(po0018));
  not_8  g03429(.A(pi220), .Y(new_n5778));
  xor_4  g03430(.A(new_n4186), .B(new_n5778), .Y(new_n5779));
  nand_5 g03431(.A(new_n3018), .B(pi181), .Y(new_n5780));
  nand_5 g03432(.A(new_n3019), .B(new_n2874), .Y(new_n5781));
  nand_5 g03433(.A(new_n5781), .B(new_n5780), .Y(new_n5782));
  xor_4  g03434(.A(new_n5782), .B(new_n5779), .Y(po0019));
  xor_4  g03435(.A(new_n5712), .B(new_n5711), .Y(po0020));
  not_8  g03436(.A(pi499), .Y(new_n5785));
  xor_4  g03437(.A(new_n5593), .B(new_n5785), .Y(new_n5786));
  not_8  g03438(.A(new_n5786), .Y(new_n5787));
  xor_4  g03439(.A(pi799), .B(new_n5693), .Y(new_n5788));
  or_6   g03440(.A(new_n5788), .B(pi219), .Y(new_n5789));
  nor_5  g03441(.A(new_n5789), .B(new_n5787), .Y(new_n5790));
  not_8  g03442(.A(new_n5790), .Y(new_n5791));
  nand_5 g03443(.A(new_n5788), .B(pi219), .Y(new_n5792));
  not_8  g03444(.A(new_n5792), .Y(new_n5793));
  nand_5 g03445(.A(new_n5793), .B(new_n5787), .Y(new_n5794));
  nand_5 g03446(.A(new_n5794), .B(new_n5791), .Y(new_n5795));
  nand_5 g03447(.A(pi799), .B(new_n5693), .Y(new_n5796));
  not_8  g03448(.A(new_n5796), .Y(new_n5797));
  xor_4  g03449(.A(pi638), .B(new_n3922), .Y(new_n5798));
  xor_4  g03450(.A(new_n5798), .B(new_n5797), .Y(new_n5799));
  xor_4  g03451(.A(new_n5799), .B(pi528), .Y(new_n5800));
  not_8  g03452(.A(pi564), .Y(new_n5801));
  nand_5 g03453(.A(new_n5594), .B(pi499), .Y(new_n5802));
  xor_4  g03454(.A(new_n5802), .B(new_n5801), .Y(new_n5803));
  xor_4  g03455(.A(new_n5803), .B(new_n5607), .Y(new_n5804));
  xor_4  g03456(.A(new_n5804), .B(new_n5800), .Y(new_n5805));
  xor_4  g03457(.A(new_n5805), .B(new_n5795), .Y(po0021));
  nor_5  g03458(.A(pi385), .B(pi130), .Y(new_n5807));
  nor_5  g03459(.A(new_n3863), .B(new_n4886), .Y(new_n5808));
  nor_5  g03460(.A(new_n5808), .B(new_n5807), .Y(new_n5809));
  xor_4  g03461(.A(new_n5809), .B(new_n4797), .Y(new_n5810));
  nor_5  g03462(.A(new_n5810), .B(new_n3861), .Y(new_n5811));
  nor_5  g03463(.A(new_n5811), .B(new_n3748), .Y(new_n5812));
  xor_4  g03464(.A(pi672), .B(pi619), .Y(new_n5813));
  nand_5 g03465(.A(new_n5807), .B(new_n4796), .Y(new_n5814));
  nand_5 g03466(.A(new_n5808), .B(new_n4797), .Y(new_n5815));
  nand_5 g03467(.A(new_n5815), .B(new_n5814), .Y(new_n5816));
  xnor_4 g03468(.A(new_n5816), .B(new_n5813), .Y(new_n5817));
  xor_4  g03469(.A(new_n5817), .B(new_n4801), .Y(new_n5818));
  xnor_4 g03470(.A(new_n5811), .B(new_n3748), .Y(new_n5819));
  nor_5  g03471(.A(new_n5819), .B(new_n5818), .Y(new_n5820));
  or_6   g03472(.A(new_n5820), .B(new_n5812), .Y(new_n5821));
  xnor_4 g03473(.A(new_n5821), .B(new_n3753), .Y(new_n5822));
  nand_5 g03474(.A(new_n5817), .B(new_n4802), .Y(new_n5823));
  nand_5 g03475(.A(new_n5816), .B(new_n5813), .Y(new_n5824));
  nand_5 g03476(.A(new_n5813), .B(pi385), .Y(new_n5825));
  nand_5 g03477(.A(new_n5825), .B(new_n5814), .Y(new_n5826));
  nand_5 g03478(.A(new_n5826), .B(new_n5824), .Y(new_n5827));
  nand_5 g03479(.A(new_n5827), .B(new_n5823), .Y(new_n5828));
  xor_4  g03480(.A(pi796), .B(pi597), .Y(new_n5829));
  nand_5 g03481(.A(pi672), .B(pi619), .Y(new_n5830));
  and_6  g03482(.A(new_n5825), .B(new_n5830), .Y(new_n5831));
  xor_4  g03483(.A(new_n5831), .B(new_n5829), .Y(new_n5832));
  nand_5 g03484(.A(new_n5832), .B(new_n4805), .Y(new_n5833));
  or_6   g03485(.A(new_n5832), .B(new_n4805), .Y(new_n5834));
  nand_5 g03486(.A(new_n5834), .B(new_n5833), .Y(new_n5835));
  xor_4  g03487(.A(new_n5835), .B(new_n5828), .Y(new_n5836));
  xnor_4 g03488(.A(new_n5836), .B(new_n5822), .Y(po0022));
  nor_5  g03489(.A(new_n5694), .B(new_n5690), .Y(new_n5838));
  xor_4  g03490(.A(new_n5838), .B(new_n5689), .Y(po0023));
  xor_4  g03491(.A(new_n4223), .B(new_n4202), .Y(po0024));
  xor_4  g03492(.A(pi246), .B(pi106), .Y(new_n5841));
  not_8  g03493(.A(pi254), .Y(new_n5842));
  nand_5 g03494(.A(new_n4904), .B(new_n5842), .Y(new_n5843));
  xor_4  g03495(.A(pi317), .B(pi254), .Y(new_n5844));
  not_8  g03496(.A(pi399), .Y(new_n5845));
  nand_5 g03497(.A(new_n4795), .B(new_n5845), .Y(new_n5846));
  xor_4  g03498(.A(pi681), .B(pi399), .Y(new_n5847));
  not_8  g03499(.A(pi261), .Y(new_n5848));
  nor_5  g03500(.A(new_n3489), .B(new_n5848), .Y(new_n5849));
  xor_4  g03501(.A(pi361), .B(pi261), .Y(new_n5850));
  not_8  g03502(.A(new_n5850), .Y(new_n5851));
  not_8  g03503(.A(pi753), .Y(new_n5852));
  nor_5  g03504(.A(new_n3629), .B(new_n5852), .Y(new_n5853));
  xor_4  g03505(.A(pi787), .B(pi753), .Y(new_n5854));
  not_8  g03506(.A(new_n5854), .Y(new_n5855));
  nand_5 g03507(.A(pi670), .B(pi455), .Y(new_n5856));
  nor_5  g03508(.A(new_n5856), .B(new_n5855), .Y(new_n5857));
  nor_5  g03509(.A(new_n5857), .B(new_n5853), .Y(new_n5858));
  nor_5  g03510(.A(new_n5858), .B(new_n5851), .Y(new_n5859));
  nor_5  g03511(.A(new_n5859), .B(new_n5849), .Y(new_n5860));
  nand_5 g03512(.A(new_n5860), .B(new_n5847), .Y(new_n5861));
  nand_5 g03513(.A(new_n5861), .B(new_n5846), .Y(new_n5862));
  nand_5 g03514(.A(new_n5862), .B(new_n5844), .Y(new_n5863));
  nand_5 g03515(.A(new_n5863), .B(new_n5843), .Y(new_n5864));
  xor_4  g03516(.A(new_n5864), .B(new_n5841), .Y(new_n5865));
  xor_4  g03517(.A(new_n5862), .B(new_n5844), .Y(new_n5866));
  nand_5 g03518(.A(new_n5866), .B(new_n3763), .Y(new_n5867));
  xor_4  g03519(.A(new_n5866), .B(new_n3763), .Y(new_n5868));
  not_8  g03520(.A(new_n5868), .Y(new_n5869));
  xor_4  g03521(.A(new_n5860), .B(new_n5847), .Y(new_n5870));
  xor_4  g03522(.A(new_n5856), .B(new_n5855), .Y(new_n5871));
  nand_5 g03523(.A(new_n5871), .B(pi488), .Y(new_n5872));
  nand_5 g03524(.A(new_n5872), .B(new_n3746), .Y(new_n5873));
  xor_4  g03525(.A(new_n5872), .B(new_n3746), .Y(new_n5874));
  xor_4  g03526(.A(new_n5858), .B(new_n5850), .Y(new_n5875));
  nand_5 g03527(.A(new_n5875), .B(new_n5874), .Y(new_n5876));
  nand_5 g03528(.A(new_n5876), .B(new_n5873), .Y(new_n5877));
  nand_5 g03529(.A(new_n5877), .B(new_n5870), .Y(new_n5878));
  not_8  g03530(.A(new_n5878), .Y(new_n5879));
  nor_5  g03531(.A(new_n5877), .B(new_n5870), .Y(new_n5880));
  nor_5  g03532(.A(new_n5880), .B(pi157), .Y(new_n5881));
  nor_5  g03533(.A(new_n5881), .B(new_n5879), .Y(new_n5882));
  or_6   g03534(.A(new_n5882), .B(new_n5869), .Y(new_n5883));
  nand_5 g03535(.A(new_n5883), .B(new_n5867), .Y(new_n5884));
  nand_5 g03536(.A(new_n5884), .B(new_n5865), .Y(new_n5885));
  xor_4  g03537(.A(new_n5884), .B(new_n5865), .Y(new_n5886));
  nand_5 g03538(.A(new_n5886), .B(new_n4756), .Y(new_n5887));
  nand_5 g03539(.A(new_n5887), .B(new_n5885), .Y(new_n5888));
  nor_5  g03540(.A(new_n5888), .B(new_n3709), .Y(new_n5889));
  xor_4  g03541(.A(new_n5888), .B(pi793), .Y(new_n5890));
  not_8  g03542(.A(pi106), .Y(new_n5891));
  nand_5 g03543(.A(new_n3484), .B(new_n5891), .Y(new_n5892));
  nand_5 g03544(.A(new_n5864), .B(new_n5841), .Y(new_n5893));
  nand_5 g03545(.A(new_n5893), .B(new_n5892), .Y(new_n5894));
  nand_5 g03546(.A(pi441), .B(pi383), .Y(new_n5895));
  not_8  g03547(.A(pi383), .Y(new_n5896));
  nand_5 g03548(.A(new_n4828), .B(new_n5896), .Y(new_n5897));
  nand_5 g03549(.A(new_n5897), .B(new_n5895), .Y(new_n5898));
  xor_4  g03550(.A(new_n5898), .B(new_n5894), .Y(new_n5899));
  not_8  g03551(.A(new_n5899), .Y(new_n5900));
  nor_5  g03552(.A(new_n5900), .B(new_n5890), .Y(new_n5901));
  or_6   g03553(.A(new_n5901), .B(new_n5889), .Y(new_n5902));
  xor_4  g03554(.A(pi823), .B(pi616), .Y(new_n5903));
  nand_5 g03555(.A(new_n5895), .B(new_n5894), .Y(new_n5904));
  nand_5 g03556(.A(new_n5904), .B(new_n5897), .Y(new_n5905));
  xor_4  g03557(.A(new_n5905), .B(new_n5903), .Y(new_n5906));
  not_8  g03558(.A(new_n5906), .Y(new_n5907));
  nand_5 g03559(.A(new_n5907), .B(new_n5902), .Y(new_n5908));
  xor_4  g03560(.A(new_n5907), .B(new_n5902), .Y(new_n5909));
  nand_5 g03561(.A(new_n5909), .B(pi623), .Y(new_n5910));
  nand_5 g03562(.A(new_n5910), .B(new_n5908), .Y(new_n5911));
  nor_5  g03563(.A(new_n5911), .B(pi013), .Y(new_n5912));
  xor_4  g03564(.A(new_n5911), .B(new_n4838), .Y(new_n5913));
  not_8  g03565(.A(pi136), .Y(new_n5914));
  nand_5 g03566(.A(new_n3473), .B(new_n5914), .Y(new_n5915));
  nand_5 g03567(.A(pi650), .B(pi136), .Y(new_n5916));
  nand_5 g03568(.A(new_n5916), .B(new_n5915), .Y(new_n5917));
  not_8  g03569(.A(pi616), .Y(new_n5918));
  not_8  g03570(.A(pi823), .Y(new_n5919));
  nand_5 g03571(.A(new_n5919), .B(new_n5918), .Y(new_n5920));
  nand_5 g03572(.A(new_n5905), .B(new_n5903), .Y(new_n5921));
  nand_5 g03573(.A(new_n5921), .B(new_n5920), .Y(new_n5922));
  not_8  g03574(.A(new_n5922), .Y(new_n5923));
  xor_4  g03575(.A(new_n5923), .B(new_n5917), .Y(new_n5924));
  not_8  g03576(.A(new_n5924), .Y(new_n5925));
  nor_5  g03577(.A(new_n5925), .B(new_n5913), .Y(new_n5926));
  or_6   g03578(.A(new_n5926), .B(new_n5912), .Y(new_n5927));
  nand_5 g03579(.A(pi303), .B(pi207), .Y(new_n5928));
  not_8  g03580(.A(pi207), .Y(new_n5929));
  nand_5 g03581(.A(new_n3423), .B(new_n5929), .Y(new_n5930));
  nand_5 g03582(.A(new_n5930), .B(new_n5928), .Y(new_n5931));
  nand_5 g03583(.A(new_n5922), .B(new_n5916), .Y(new_n5932));
  nand_5 g03584(.A(new_n5932), .B(new_n5915), .Y(new_n5933));
  not_8  g03585(.A(new_n5933), .Y(new_n5934));
  xor_4  g03586(.A(new_n5934), .B(new_n5931), .Y(new_n5935));
  or_6   g03587(.A(new_n5935), .B(new_n5927), .Y(new_n5936));
  nand_5 g03588(.A(new_n5935), .B(new_n5927), .Y(new_n5937));
  nand_5 g03589(.A(new_n5937), .B(new_n5936), .Y(new_n5938));
  xor_4  g03590(.A(new_n5938), .B(new_n4857), .Y(new_n5939));
  not_8  g03591(.A(pi146), .Y(new_n5940));
  not_8  g03592(.A(pi143), .Y(new_n5941));
  not_8  g03593(.A(pi352), .Y(new_n5942));
  nand_5 g03594(.A(new_n5942), .B(new_n5941), .Y(new_n5943));
  nand_5 g03595(.A(pi352), .B(pi143), .Y(new_n5944));
  nand_5 g03596(.A(new_n5944), .B(new_n5943), .Y(new_n5945));
  nand_5 g03597(.A(pi177), .B(pi081), .Y(new_n5946));
  not_8  g03598(.A(pi081), .Y(new_n5947));
  nand_5 g03599(.A(new_n3805), .B(new_n5947), .Y(new_n5948));
  nand_5 g03600(.A(pi019), .B(pi012), .Y(new_n5949));
  nor_5  g03601(.A(pi628), .B(pi027), .Y(new_n5950));
  nor_5  g03602(.A(pi830), .B(pi597), .Y(new_n5951));
  xor_4  g03603(.A(pi830), .B(new_n3828), .Y(new_n5952));
  not_8  g03604(.A(pi696), .Y(new_n5953));
  nor_5  g03605(.A(new_n5953), .B(new_n3814), .Y(new_n5954));
  nor_5  g03606(.A(new_n5954), .B(new_n5952), .Y(new_n5955));
  nor_5  g03607(.A(new_n5955), .B(new_n5951), .Y(new_n5956));
  xor_4  g03608(.A(pi628), .B(new_n3811), .Y(new_n5957));
  nor_5  g03609(.A(new_n5957), .B(new_n5956), .Y(new_n5958));
  nor_5  g03610(.A(new_n5958), .B(new_n5950), .Y(new_n5959));
  xor_4  g03611(.A(pi019), .B(pi012), .Y(new_n5960));
  nand_5 g03612(.A(new_n5960), .B(new_n5959), .Y(new_n5961));
  nand_5 g03613(.A(new_n5961), .B(new_n5949), .Y(new_n5962));
  nand_5 g03614(.A(new_n5962), .B(new_n5948), .Y(new_n5963));
  nand_5 g03615(.A(new_n5963), .B(new_n5946), .Y(new_n5964));
  xor_4  g03616(.A(new_n5964), .B(new_n5945), .Y(new_n5965));
  nor_5  g03617(.A(new_n5965), .B(new_n5940), .Y(new_n5966));
  xor_4  g03618(.A(new_n5965), .B(new_n5940), .Y(new_n5967));
  not_8  g03619(.A(new_n5967), .Y(new_n5968));
  nand_5 g03620(.A(new_n5948), .B(new_n5946), .Y(new_n5969));
  xnor_4 g03621(.A(new_n5969), .B(new_n5962), .Y(new_n5970));
  or_6   g03622(.A(new_n5970), .B(pi120), .Y(new_n5971));
  xor_4  g03623(.A(new_n5970), .B(pi120), .Y(new_n5972));
  xor_4  g03624(.A(new_n5960), .B(new_n5959), .Y(new_n5973));
  nor_5  g03625(.A(new_n5973), .B(pi432), .Y(new_n5974));
  xor_4  g03626(.A(new_n5973), .B(pi432), .Y(new_n5975));
  not_8  g03627(.A(new_n5975), .Y(new_n5976));
  not_8  g03628(.A(pi645), .Y(new_n5977));
  xor_4  g03629(.A(new_n5957), .B(new_n5956), .Y(new_n5978));
  or_6   g03630(.A(new_n5978), .B(new_n5977), .Y(new_n5979));
  xor_4  g03631(.A(new_n5978), .B(new_n5977), .Y(new_n5980));
  xor_4  g03632(.A(new_n5954), .B(new_n5952), .Y(new_n5981));
  or_6   g03633(.A(new_n5981), .B(new_n4149), .Y(new_n5982));
  xor_4  g03634(.A(new_n5981), .B(new_n4149), .Y(new_n5983));
  xor_4  g03635(.A(pi696), .B(new_n3814), .Y(new_n5984));
  nor_5  g03636(.A(new_n5984), .B(new_n4152), .Y(new_n5985));
  xor_4  g03637(.A(new_n5984), .B(new_n4152), .Y(new_n5986));
  not_8  g03638(.A(new_n5986), .Y(new_n5987));
  nand_5 g03639(.A(new_n3863), .B(new_n5778), .Y(new_n5988));
  nand_5 g03640(.A(pi385), .B(pi220), .Y(new_n5989));
  nand_5 g03641(.A(new_n5989), .B(new_n4184), .Y(new_n5990));
  nand_5 g03642(.A(new_n5990), .B(new_n5988), .Y(new_n5991));
  nor_5  g03643(.A(new_n5991), .B(new_n5987), .Y(new_n5992));
  or_6   g03644(.A(new_n5992), .B(new_n5985), .Y(new_n5993));
  nand_5 g03645(.A(new_n5993), .B(new_n5983), .Y(new_n5994));
  nand_5 g03646(.A(new_n5994), .B(new_n5982), .Y(new_n5995));
  nand_5 g03647(.A(new_n5995), .B(new_n5980), .Y(new_n5996));
  nand_5 g03648(.A(new_n5996), .B(new_n5979), .Y(new_n5997));
  nor_5  g03649(.A(new_n5997), .B(new_n5976), .Y(new_n5998));
  nor_5  g03650(.A(new_n5998), .B(new_n5974), .Y(new_n5999));
  not_8  g03651(.A(new_n5999), .Y(new_n6000));
  nand_5 g03652(.A(new_n6000), .B(new_n5972), .Y(new_n6001));
  nand_5 g03653(.A(new_n6001), .B(new_n5971), .Y(new_n6002));
  nor_5  g03654(.A(new_n6002), .B(new_n5968), .Y(new_n6003));
  nor_5  g03655(.A(new_n6003), .B(new_n5966), .Y(new_n6004));
  not_8  g03656(.A(pi162), .Y(new_n6005));
  xor_4  g03657(.A(pi382), .B(new_n6005), .Y(new_n6006));
  nand_5 g03658(.A(new_n5964), .B(new_n5943), .Y(new_n6007));
  nand_5 g03659(.A(new_n6007), .B(new_n5944), .Y(new_n6008));
  xor_4  g03660(.A(new_n6008), .B(new_n6006), .Y(new_n6009));
  xor_4  g03661(.A(new_n6009), .B(pi621), .Y(new_n6010));
  xor_4  g03662(.A(new_n6010), .B(new_n6004), .Y(new_n6011));
  xor_4  g03663(.A(new_n5886), .B(new_n4756), .Y(new_n6012));
  not_8  g03664(.A(new_n6012), .Y(new_n6013));
  xor_4  g03665(.A(new_n5995), .B(new_n5980), .Y(new_n6014));
  not_8  g03666(.A(new_n6014), .Y(new_n6015));
  xor_4  g03667(.A(new_n5993), .B(new_n5983), .Y(new_n6016));
  not_8  g03668(.A(new_n6016), .Y(new_n6017));
  not_8  g03669(.A(pi488), .Y(new_n6018));
  xor_4  g03670(.A(new_n5871), .B(new_n6018), .Y(new_n6019));
  xor_4  g03671(.A(new_n5991), .B(new_n5986), .Y(new_n6020));
  not_8  g03672(.A(new_n6020), .Y(new_n6021));
  or_6   g03673(.A(new_n6021), .B(new_n6019), .Y(new_n6022));
  nand_5 g03674(.A(new_n6021), .B(new_n6019), .Y(new_n6023));
  xor_4  g03675(.A(pi670), .B(pi455), .Y(new_n6024));
  nand_5 g03676(.A(new_n6024), .B(pi631), .Y(new_n6025));
  not_8  g03677(.A(new_n6024), .Y(new_n6026));
  nand_5 g03678(.A(new_n6026), .B(new_n3860), .Y(new_n6027));
  nand_5 g03679(.A(new_n6027), .B(new_n5779), .Y(new_n6028));
  nand_5 g03680(.A(new_n6028), .B(new_n6025), .Y(new_n6029));
  nand_5 g03681(.A(new_n6029), .B(new_n6023), .Y(new_n6030));
  nand_5 g03682(.A(new_n6030), .B(new_n6022), .Y(new_n6031));
  nand_5 g03683(.A(new_n6031), .B(new_n6017), .Y(new_n6032));
  xor_4  g03684(.A(new_n6031), .B(new_n6016), .Y(new_n6033));
  xor_4  g03685(.A(new_n5875), .B(new_n5874), .Y(new_n6034));
  or_6   g03686(.A(new_n6034), .B(new_n6033), .Y(new_n6035));
  nand_5 g03687(.A(new_n6035), .B(new_n6032), .Y(new_n6036));
  nand_5 g03688(.A(new_n6036), .B(new_n6015), .Y(new_n6037));
  nor_5  g03689(.A(new_n5880), .B(new_n5879), .Y(new_n6038));
  xor_4  g03690(.A(new_n6038), .B(new_n3758), .Y(new_n6039));
  xor_4  g03691(.A(new_n6036), .B(new_n6014), .Y(new_n6040));
  or_6   g03692(.A(new_n6040), .B(new_n6039), .Y(new_n6041));
  nand_5 g03693(.A(new_n6041), .B(new_n6037), .Y(new_n6042));
  xor_4  g03694(.A(new_n5997), .B(new_n5975), .Y(new_n6043));
  not_8  g03695(.A(new_n6043), .Y(new_n6044));
  nand_5 g03696(.A(new_n6044), .B(new_n6042), .Y(new_n6045));
  xor_4  g03697(.A(new_n6043), .B(new_n6042), .Y(new_n6046));
  xor_4  g03698(.A(new_n5882), .B(new_n5869), .Y(new_n6047));
  or_6   g03699(.A(new_n6047), .B(new_n6046), .Y(new_n6048));
  nand_5 g03700(.A(new_n6048), .B(new_n6045), .Y(new_n6049));
  nand_5 g03701(.A(new_n6049), .B(new_n6013), .Y(new_n6050));
  xor_4  g03702(.A(new_n6049), .B(new_n6012), .Y(new_n6051));
  xor_4  g03703(.A(new_n5999), .B(new_n5972), .Y(new_n6052));
  or_6   g03704(.A(new_n6052), .B(new_n6051), .Y(new_n6053));
  nand_5 g03705(.A(new_n6053), .B(new_n6050), .Y(new_n6054));
  xor_4  g03706(.A(new_n6002), .B(new_n5967), .Y(new_n6055));
  nor_5  g03707(.A(new_n6055), .B(new_n6054), .Y(new_n6056));
  xor_4  g03708(.A(new_n6055), .B(new_n6054), .Y(new_n6057));
  not_8  g03709(.A(new_n6057), .Y(new_n6058));
  xor_4  g03710(.A(new_n5900), .B(new_n5890), .Y(new_n6059));
  nor_5  g03711(.A(new_n6059), .B(new_n6058), .Y(new_n6060));
  or_6   g03712(.A(new_n6060), .B(new_n6056), .Y(new_n6061));
  nor_5  g03713(.A(new_n6061), .B(new_n6011), .Y(new_n6062));
  not_8  g03714(.A(new_n6011), .Y(new_n6063));
  xor_4  g03715(.A(new_n6061), .B(new_n6063), .Y(new_n6064));
  xor_4  g03716(.A(new_n5909), .B(new_n4843), .Y(new_n6065));
  nor_5  g03717(.A(new_n6065), .B(new_n6064), .Y(new_n6066));
  or_6   g03718(.A(new_n6066), .B(new_n6062), .Y(new_n6067));
  xor_4  g03719(.A(pi185), .B(pi066), .Y(new_n6068));
  nand_5 g03720(.A(pi382), .B(pi162), .Y(new_n6069));
  not_8  g03721(.A(new_n6006), .Y(new_n6070));
  nand_5 g03722(.A(new_n6008), .B(new_n6070), .Y(new_n6071));
  nand_5 g03723(.A(new_n6071), .B(new_n6069), .Y(new_n6072));
  xor_4  g03724(.A(new_n6072), .B(new_n6068), .Y(new_n6073));
  or_6   g03725(.A(new_n6073), .B(pi092), .Y(new_n6074));
  nand_5 g03726(.A(new_n6073), .B(pi092), .Y(new_n6075));
  nand_5 g03727(.A(new_n6075), .B(new_n6074), .Y(new_n6076));
  not_8  g03728(.A(pi621), .Y(new_n6077));
  or_6   g03729(.A(new_n6009), .B(new_n6077), .Y(new_n6078));
  or_6   g03730(.A(new_n6010), .B(new_n6004), .Y(new_n6079));
  nand_5 g03731(.A(new_n6079), .B(new_n6078), .Y(new_n6080));
  xor_4  g03732(.A(new_n6080), .B(new_n6076), .Y(new_n6081));
  nand_5 g03733(.A(new_n6081), .B(new_n6067), .Y(new_n6082));
  or_6   g03734(.A(new_n6081), .B(new_n6067), .Y(new_n6083));
  xor_4  g03735(.A(new_n5924), .B(new_n5913), .Y(new_n6084));
  nand_5 g03736(.A(new_n6084), .B(new_n6083), .Y(new_n6085));
  nand_5 g03737(.A(new_n6085), .B(new_n6082), .Y(new_n6086));
  not_8  g03738(.A(new_n6080), .Y(new_n6087));
  nand_5 g03739(.A(new_n6087), .B(new_n6075), .Y(new_n6088));
  nand_5 g03740(.A(new_n6088), .B(new_n6074), .Y(new_n6089));
  not_8  g03741(.A(new_n6089), .Y(new_n6090));
  not_8  g03742(.A(pi280), .Y(new_n6091));
  xor_4  g03743(.A(pi661), .B(new_n6091), .Y(new_n6092));
  nand_5 g03744(.A(pi185), .B(pi066), .Y(new_n6093));
  nand_5 g03745(.A(new_n6072), .B(new_n6068), .Y(new_n6094));
  nand_5 g03746(.A(new_n6094), .B(new_n6093), .Y(new_n6095));
  nand_5 g03747(.A(new_n6095), .B(pi121), .Y(new_n6096));
  nor_5  g03748(.A(new_n6095), .B(pi121), .Y(new_n6097));
  not_8  g03749(.A(new_n6097), .Y(new_n6098));
  nand_5 g03750(.A(new_n6098), .B(new_n6096), .Y(new_n6099));
  xnor_4 g03751(.A(new_n6099), .B(new_n6092), .Y(new_n6100));
  xor_4  g03752(.A(new_n6100), .B(new_n6090), .Y(new_n6101));
  xor_4  g03753(.A(new_n6101), .B(new_n6086), .Y(new_n6102));
  xnor_4 g03754(.A(new_n6102), .B(new_n5939), .Y(po0025));
  xor_4  g03755(.A(pi826), .B(pi433), .Y(new_n6104));
  not_8  g03756(.A(new_n6104), .Y(new_n6105));
  not_8  g03757(.A(pi210), .Y(new_n6106));
  nand_5 g03758(.A(new_n3894), .B(new_n6106), .Y(new_n6107));
  xor_4  g03759(.A(pi568), .B(pi210), .Y(new_n6108));
  not_8  g03760(.A(pi129), .Y(new_n6109));
  nand_5 g03761(.A(new_n4005), .B(new_n6109), .Y(new_n6110));
  not_8  g03762(.A(new_n6110), .Y(new_n6111));
  xor_4  g03763(.A(pi183), .B(pi129), .Y(new_n6112));
  not_8  g03764(.A(new_n6112), .Y(new_n6113));
  nand_5 g03765(.A(new_n3933), .B(new_n4112), .Y(new_n6114));
  not_8  g03766(.A(new_n6114), .Y(new_n6115));
  nor_5  g03767(.A(new_n4113), .B(new_n4111), .Y(new_n6116));
  nor_5  g03768(.A(new_n6116), .B(new_n6115), .Y(new_n6117));
  nor_5  g03769(.A(new_n6117), .B(new_n6113), .Y(new_n6118));
  nor_5  g03770(.A(new_n6118), .B(new_n6111), .Y(new_n6119));
  not_8  g03771(.A(new_n6119), .Y(new_n6120));
  nand_5 g03772(.A(new_n6120), .B(new_n6108), .Y(new_n6121));
  nand_5 g03773(.A(new_n6121), .B(new_n6107), .Y(new_n6122));
  xor_4  g03774(.A(new_n6122), .B(new_n6105), .Y(new_n6123));
  not_8  g03775(.A(new_n6123), .Y(new_n6124));
  xor_4  g03776(.A(pi609), .B(pi271), .Y(new_n6125));
  nor_5  g03777(.A(pi356), .B(pi218), .Y(new_n6126));
  nand_5 g03778(.A(pi656), .B(pi307), .Y(new_n6127));
  not_8  g03779(.A(new_n6127), .Y(new_n6128));
  xor_4  g03780(.A(pi356), .B(new_n3976), .Y(new_n6129));
  nor_5  g03781(.A(new_n6129), .B(new_n6128), .Y(new_n6130));
  nor_5  g03782(.A(new_n6130), .B(new_n6126), .Y(new_n6131));
  xor_4  g03783(.A(new_n6131), .B(new_n6125), .Y(new_n6132));
  xor_4  g03784(.A(new_n6129), .B(new_n6127), .Y(new_n6133));
  not_8  g03785(.A(new_n6133), .Y(new_n6134));
  xor_4  g03786(.A(pi656), .B(pi307), .Y(new_n6135));
  nand_5 g03787(.A(new_n6135), .B(pi219), .Y(new_n6136));
  not_8  g03788(.A(new_n6136), .Y(new_n6137));
  nor_5  g03789(.A(new_n6135), .B(pi219), .Y(new_n6138));
  or_6   g03790(.A(new_n6138), .B(new_n6137), .Y(new_n6139));
  nand_5 g03791(.A(new_n6139), .B(new_n2572), .Y(new_n6140));
  xor_4  g03792(.A(new_n6140), .B(new_n3971), .Y(new_n6141));
  or_6   g03793(.A(new_n6141), .B(new_n6134), .Y(new_n6142));
  and_6  g03794(.A(new_n6135), .B(new_n2572), .Y(new_n6143));
  nand_5 g03795(.A(new_n6143), .B(new_n6141), .Y(new_n6144));
  nand_5 g03796(.A(new_n6144), .B(new_n6142), .Y(new_n6145));
  nand_5 g03797(.A(new_n6145), .B(new_n6132), .Y(new_n6146));
  not_8  g03798(.A(new_n6146), .Y(new_n6147));
  not_8  g03799(.A(new_n6132), .Y(new_n6148));
  xor_4  g03800(.A(new_n6145), .B(new_n6148), .Y(new_n6149));
  nor_5  g03801(.A(new_n6149), .B(new_n3968), .Y(new_n6150));
  nor_5  g03802(.A(new_n6150), .B(new_n6147), .Y(new_n6151));
  nand_5 g03803(.A(new_n6151), .B(new_n3961), .Y(new_n6152));
  xor_4  g03804(.A(pi614), .B(pi147), .Y(new_n6153));
  nand_5 g03805(.A(pi609), .B(pi271), .Y(new_n6154));
  nand_5 g03806(.A(new_n6131), .B(new_n6125), .Y(new_n6155));
  nand_5 g03807(.A(new_n6155), .B(new_n6154), .Y(new_n6156));
  xor_4  g03808(.A(new_n6156), .B(new_n6153), .Y(new_n6157));
  not_8  g03809(.A(new_n6157), .Y(new_n6158));
  xor_4  g03810(.A(new_n6151), .B(new_n3961), .Y(new_n6159));
  nand_5 g03811(.A(new_n6159), .B(new_n6158), .Y(new_n6160));
  nand_5 g03812(.A(new_n6160), .B(new_n6152), .Y(new_n6161));
  nand_5 g03813(.A(pi614), .B(pi147), .Y(new_n6162));
  nand_5 g03814(.A(new_n6156), .B(new_n6153), .Y(new_n6163));
  nand_5 g03815(.A(new_n6163), .B(new_n6162), .Y(new_n6164));
  not_8  g03816(.A(pi644), .Y(new_n6165));
  nand_5 g03817(.A(new_n6165), .B(new_n3999), .Y(new_n6166));
  nand_5 g03818(.A(pi644), .B(pi602), .Y(new_n6167));
  nand_5 g03819(.A(new_n6167), .B(new_n6166), .Y(new_n6168));
  xor_4  g03820(.A(new_n6168), .B(new_n6164), .Y(new_n6169));
  not_8  g03821(.A(new_n6169), .Y(new_n6170));
  xor_4  g03822(.A(new_n6170), .B(new_n3998), .Y(new_n6171));
  xor_4  g03823(.A(new_n6171), .B(new_n6161), .Y(new_n6172));
  xor_4  g03824(.A(new_n6119), .B(new_n6108), .Y(new_n6173));
  or_6   g03825(.A(new_n6173), .B(new_n6172), .Y(new_n6174));
  xor_4  g03826(.A(new_n6173), .B(new_n6172), .Y(new_n6175));
  xor_4  g03827(.A(new_n6159), .B(new_n6157), .Y(new_n6176));
  xor_4  g03828(.A(new_n6117), .B(new_n6112), .Y(new_n6177));
  not_8  g03829(.A(new_n6177), .Y(new_n6178));
  nor_5  g03830(.A(new_n6178), .B(new_n6176), .Y(new_n6179));
  xor_4  g03831(.A(new_n6177), .B(new_n6176), .Y(new_n6180));
  not_8  g03832(.A(new_n4114), .Y(new_n6181));
  xnor_4 g03833(.A(new_n6135), .B(new_n2572), .Y(new_n6182));
  nand_5 g03834(.A(new_n6182), .B(new_n4117), .Y(new_n6183));
  nand_5 g03835(.A(new_n6183), .B(new_n4116), .Y(new_n6184));
  nand_5 g03836(.A(new_n6184), .B(new_n4115), .Y(new_n6185));
  xor_4  g03837(.A(new_n6141), .B(new_n6133), .Y(new_n6186));
  xor_4  g03838(.A(new_n6184), .B(new_n4115), .Y(new_n6187));
  nand_5 g03839(.A(new_n6187), .B(new_n6186), .Y(new_n6188));
  nand_5 g03840(.A(new_n6188), .B(new_n6185), .Y(new_n6189));
  and_6  g03841(.A(new_n6189), .B(new_n6181), .Y(new_n6190));
  xor_4  g03842(.A(new_n6189), .B(new_n4114), .Y(new_n6191));
  xor_4  g03843(.A(new_n6149), .B(new_n3968), .Y(new_n6192));
  nor_5  g03844(.A(new_n6192), .B(new_n6191), .Y(new_n6193));
  nor_5  g03845(.A(new_n6193), .B(new_n6190), .Y(new_n6194));
  nor_5  g03846(.A(new_n6194), .B(new_n6180), .Y(new_n6195));
  or_6   g03847(.A(new_n6195), .B(new_n6179), .Y(new_n6196));
  not_8  g03848(.A(new_n6196), .Y(new_n6197));
  nand_5 g03849(.A(new_n6197), .B(new_n6175), .Y(new_n6198));
  nand_5 g03850(.A(new_n6198), .B(new_n6174), .Y(new_n6199));
  nor_5  g03851(.A(new_n6199), .B(new_n6124), .Y(new_n6200));
  not_8  g03852(.A(pi726), .Y(new_n6201));
  nand_5 g03853(.A(new_n6201), .B(new_n4060), .Y(new_n6202));
  nand_5 g03854(.A(pi726), .B(pi394), .Y(new_n6203));
  and_6  g03855(.A(new_n6203), .B(new_n6202), .Y(new_n6204));
  nand_5 g03856(.A(new_n6166), .B(new_n6164), .Y(new_n6205));
  nand_5 g03857(.A(new_n6205), .B(new_n6167), .Y(new_n6206));
  xor_4  g03858(.A(new_n6206), .B(new_n6204), .Y(new_n6207));
  xor_4  g03859(.A(new_n6207), .B(new_n4065), .Y(new_n6208));
  or_6   g03860(.A(new_n6170), .B(new_n3998), .Y(new_n6209));
  nand_5 g03861(.A(new_n6171), .B(new_n6161), .Y(new_n6210));
  nand_5 g03862(.A(new_n6210), .B(new_n6209), .Y(new_n6211));
  xnor_4 g03863(.A(new_n6211), .B(new_n6208), .Y(new_n6212));
  xor_4  g03864(.A(new_n6199), .B(new_n6123), .Y(new_n6213));
  nor_5  g03865(.A(new_n6213), .B(new_n6212), .Y(new_n6214));
  or_6   g03866(.A(new_n6214), .B(new_n6200), .Y(new_n6215));
  nand_5 g03867(.A(pi826), .B(pi433), .Y(new_n6216));
  not_8  g03868(.A(new_n6216), .Y(new_n6217));
  nor_5  g03869(.A(new_n6122), .B(new_n6105), .Y(new_n6218));
  nor_5  g03870(.A(new_n6218), .B(new_n6217), .Y(new_n6219));
  not_8  g03871(.A(pi150), .Y(new_n6220));
  not_8  g03872(.A(pi707), .Y(new_n6221));
  nand_5 g03873(.A(new_n6221), .B(new_n6220), .Y(new_n6222));
  nand_5 g03874(.A(pi707), .B(pi150), .Y(new_n6223));
  nand_5 g03875(.A(new_n6223), .B(new_n6222), .Y(new_n6224));
  xor_4  g03876(.A(new_n6224), .B(new_n6219), .Y(new_n6225));
  or_6   g03877(.A(new_n6225), .B(new_n6215), .Y(new_n6226));
  xor_4  g03878(.A(new_n6225), .B(new_n6215), .Y(new_n6227));
  or_6   g03879(.A(new_n6207), .B(new_n4065), .Y(new_n6228));
  nand_5 g03880(.A(new_n6211), .B(new_n6208), .Y(new_n6229));
  nand_5 g03881(.A(new_n6229), .B(new_n6228), .Y(new_n6230));
  xor_4  g03882(.A(pi647), .B(pi578), .Y(new_n6231));
  nand_5 g03883(.A(new_n6206), .B(new_n6202), .Y(new_n6232));
  nand_5 g03884(.A(new_n6232), .B(new_n6203), .Y(new_n6233));
  xor_4  g03885(.A(new_n6233), .B(new_n6231), .Y(new_n6234));
  xor_4  g03886(.A(new_n6234), .B(new_n6230), .Y(new_n6235));
  not_8  g03887(.A(pi418), .Y(new_n6236));
  not_8  g03888(.A(pi791), .Y(new_n6237));
  nand_5 g03889(.A(new_n3952), .B(new_n3949), .Y(new_n6238));
  nor_5  g03890(.A(new_n6238), .B(pi606), .Y(new_n6239));
  not_8  g03891(.A(new_n6239), .Y(new_n6240));
  not_8  g03892(.A(pi479), .Y(new_n6241));
  nand_5 g03893(.A(new_n6241), .B(new_n3944), .Y(new_n6242));
  nor_5  g03894(.A(new_n6242), .B(new_n6240), .Y(new_n6243));
  nand_5 g03895(.A(new_n6243), .B(new_n6237), .Y(new_n6244));
  not_8  g03896(.A(new_n6244), .Y(new_n6245));
  nand_5 g03897(.A(new_n6245), .B(new_n6236), .Y(new_n6246));
  nand_5 g03898(.A(new_n6244), .B(pi418), .Y(new_n6247));
  nand_5 g03899(.A(new_n6247), .B(new_n6246), .Y(new_n6248));
  xor_4  g03900(.A(new_n6248), .B(new_n5644), .Y(new_n6249));
  nand_5 g03901(.A(new_n6237), .B(pi613), .Y(new_n6250));
  not_8  g03902(.A(new_n6250), .Y(new_n6251));
  nor_5  g03903(.A(new_n4064), .B(new_n4063), .Y(new_n6252));
  nor_5  g03904(.A(new_n6252), .B(new_n6251), .Y(new_n6253));
  nor_5  g03905(.A(new_n6253), .B(new_n6245), .Y(new_n6254));
  xor_4  g03906(.A(new_n6254), .B(new_n6249), .Y(new_n6255));
  xnor_4 g03907(.A(new_n6255), .B(new_n6235), .Y(new_n6256));
  nand_5 g03908(.A(new_n6256), .B(new_n6227), .Y(new_n6257));
  nand_5 g03909(.A(new_n6257), .B(new_n6226), .Y(new_n6258));
  not_8  g03910(.A(pi249), .Y(new_n6259));
  not_8  g03911(.A(pi782), .Y(new_n6260));
  nand_5 g03912(.A(new_n6260), .B(new_n6259), .Y(new_n6261));
  nand_5 g03913(.A(pi782), .B(pi249), .Y(new_n6262));
  nand_5 g03914(.A(new_n6262), .B(new_n6261), .Y(new_n6263));
  not_8  g03915(.A(new_n6223), .Y(new_n6264));
  not_8  g03916(.A(new_n6222), .Y(new_n6265));
  nor_5  g03917(.A(new_n6265), .B(new_n6219), .Y(new_n6266));
  nor_5  g03918(.A(new_n6266), .B(new_n6264), .Y(new_n6267));
  not_8  g03919(.A(new_n6267), .Y(new_n6268));
  xor_4  g03920(.A(new_n6268), .B(new_n6263), .Y(new_n6269));
  nor_5  g03921(.A(new_n6269), .B(new_n6258), .Y(new_n6270));
  not_8  g03922(.A(new_n6269), .Y(new_n6271));
  xor_4  g03923(.A(new_n6271), .B(new_n6258), .Y(new_n6272));
  nand_5 g03924(.A(new_n6254), .B(new_n6249), .Y(new_n6273));
  not_8  g03925(.A(new_n6246), .Y(new_n6274));
  nor_5  g03926(.A(new_n6248), .B(new_n5644), .Y(new_n6275));
  nor_5  g03927(.A(new_n6275), .B(new_n6274), .Y(new_n6276));
  nand_5 g03928(.A(new_n6276), .B(new_n6273), .Y(new_n6277));
  xor_4  g03929(.A(new_n6277), .B(pi834), .Y(new_n6278));
  xor_4  g03930(.A(new_n6278), .B(pi054), .Y(new_n6279));
  not_8  g03931(.A(new_n6234), .Y(new_n6280));
  nand_5 g03932(.A(new_n6280), .B(new_n6230), .Y(new_n6281));
  or_6   g03933(.A(new_n6255), .B(new_n6235), .Y(new_n6282));
  nand_5 g03934(.A(new_n6282), .B(new_n6281), .Y(new_n6283));
  xor_4  g03935(.A(pi554), .B(pi205), .Y(new_n6284));
  nor_5  g03936(.A(pi647), .B(pi578), .Y(new_n6285));
  not_8  g03937(.A(new_n6231), .Y(new_n6286));
  nor_5  g03938(.A(new_n6233), .B(new_n6286), .Y(new_n6287));
  nor_5  g03939(.A(new_n6287), .B(new_n6285), .Y(new_n6288));
  xor_4  g03940(.A(new_n6288), .B(new_n6284), .Y(new_n6289));
  xor_4  g03941(.A(new_n6289), .B(new_n6283), .Y(new_n6290));
  xor_4  g03942(.A(new_n6290), .B(new_n6279), .Y(new_n6291));
  nor_5  g03943(.A(new_n6291), .B(new_n6272), .Y(new_n6292));
  or_6   g03944(.A(new_n6292), .B(new_n6270), .Y(new_n6293));
  not_8  g03945(.A(pi126), .Y(new_n6294));
  not_8  g03946(.A(pi789), .Y(new_n6295));
  nand_5 g03947(.A(new_n6295), .B(new_n6294), .Y(new_n6296));
  nand_5 g03948(.A(pi789), .B(pi126), .Y(new_n6297));
  and_6  g03949(.A(new_n6297), .B(new_n6296), .Y(new_n6298));
  nand_5 g03950(.A(new_n6268), .B(new_n6261), .Y(new_n6299));
  nand_5 g03951(.A(new_n6299), .B(new_n6262), .Y(new_n6300));
  xor_4  g03952(.A(new_n6300), .B(new_n6298), .Y(new_n6301));
  nor_5  g03953(.A(new_n6301), .B(new_n6293), .Y(new_n6302));
  nor_5  g03954(.A(pi554), .B(pi205), .Y(new_n6303));
  not_8  g03955(.A(new_n6284), .Y(new_n6304));
  nor_5  g03956(.A(new_n6288), .B(new_n6304), .Y(new_n6305));
  nor_5  g03957(.A(new_n6305), .B(new_n6303), .Y(new_n6306));
  not_8  g03958(.A(pi247), .Y(new_n6307));
  xor_4  g03959(.A(pi419), .B(new_n6307), .Y(new_n6308));
  xor_4  g03960(.A(new_n6308), .B(new_n6306), .Y(new_n6309));
  not_8  g03961(.A(new_n6309), .Y(new_n6310));
  not_8  g03962(.A(new_n6289), .Y(new_n6311));
  nor_5  g03963(.A(new_n6311), .B(new_n6283), .Y(new_n6312));
  nor_5  g03964(.A(new_n6290), .B(new_n6279), .Y(new_n6313));
  or_6   g03965(.A(new_n6313), .B(new_n6312), .Y(new_n6314));
  xor_4  g03966(.A(new_n6314), .B(new_n6310), .Y(new_n6315));
  not_8  g03967(.A(pi054), .Y(new_n6316));
  nand_5 g03968(.A(new_n6274), .B(new_n6316), .Y(new_n6317));
  xor_4  g03969(.A(new_n6317), .B(pi032), .Y(new_n6318));
  xor_4  g03970(.A(new_n6318), .B(pi472), .Y(new_n6319));
  not_8  g03971(.A(new_n6319), .Y(new_n6320));
  nand_5 g03972(.A(new_n6278), .B(pi054), .Y(new_n6321));
  nor_5  g03973(.A(new_n6277), .B(pi834), .Y(new_n6322));
  not_8  g03974(.A(new_n6317), .Y(new_n6323));
  nor_5  g03975(.A(new_n6323), .B(new_n6322), .Y(new_n6324));
  nand_5 g03976(.A(new_n6324), .B(new_n6321), .Y(new_n6325));
  xor_4  g03977(.A(new_n6325), .B(new_n6320), .Y(new_n6326));
  not_8  g03978(.A(new_n6326), .Y(new_n6327));
  xor_4  g03979(.A(new_n6327), .B(new_n6315), .Y(new_n6328));
  not_8  g03980(.A(new_n6301), .Y(new_n6329));
  xor_4  g03981(.A(new_n6329), .B(new_n6293), .Y(new_n6330));
  nor_5  g03982(.A(new_n6330), .B(new_n6328), .Y(new_n6331));
  nor_5  g03983(.A(new_n6331), .B(new_n6302), .Y(new_n6332));
  xor_4  g03984(.A(pi490), .B(pi197), .Y(new_n6333));
  nand_5 g03985(.A(new_n6300), .B(new_n6296), .Y(new_n6334));
  nand_5 g03986(.A(new_n6334), .B(new_n6297), .Y(new_n6335));
  xor_4  g03987(.A(new_n6335), .B(new_n6333), .Y(new_n6336));
  nand_5 g03988(.A(new_n6336), .B(new_n6332), .Y(new_n6337));
  not_8  g03989(.A(new_n6336), .Y(new_n6338));
  xor_4  g03990(.A(new_n6338), .B(new_n6332), .Y(new_n6339));
  or_6   g03991(.A(new_n6314), .B(new_n6310), .Y(new_n6340));
  nand_5 g03992(.A(new_n6327), .B(new_n6315), .Y(new_n6341));
  nand_5 g03993(.A(new_n6341), .B(new_n6340), .Y(new_n6342));
  xor_4  g03994(.A(pi335), .B(pi056), .Y(new_n6343));
  nor_5  g03995(.A(pi419), .B(pi247), .Y(new_n6344));
  nor_5  g03996(.A(new_n6308), .B(new_n6306), .Y(new_n6345));
  nor_5  g03997(.A(new_n6345), .B(new_n6344), .Y(new_n6346));
  xor_4  g03998(.A(new_n6346), .B(new_n6343), .Y(new_n6347));
  xor_4  g03999(.A(new_n6347), .B(new_n6342), .Y(new_n6348));
  nand_5 g04000(.A(new_n6318), .B(pi472), .Y(new_n6349));
  or_6   g04001(.A(new_n6325), .B(new_n6320), .Y(new_n6350));
  nand_5 g04002(.A(new_n6350), .B(new_n6349), .Y(new_n6351));
  not_8  g04003(.A(pi110), .Y(new_n6352));
  not_8  g04004(.A(pi032), .Y(new_n6353));
  nand_5 g04005(.A(new_n6323), .B(new_n6353), .Y(new_n6354));
  not_8  g04006(.A(new_n6354), .Y(new_n6355));
  nand_5 g04007(.A(new_n6355), .B(new_n6352), .Y(new_n6356));
  nand_5 g04008(.A(new_n6354), .B(pi110), .Y(new_n6357));
  nand_5 g04009(.A(new_n6357), .B(new_n6356), .Y(new_n6358));
  xor_4  g04010(.A(new_n6358), .B(new_n5634), .Y(new_n6359));
  xor_4  g04011(.A(new_n6359), .B(new_n6351), .Y(new_n6360));
  not_8  g04012(.A(new_n6360), .Y(new_n6361));
  xor_4  g04013(.A(new_n6361), .B(new_n6348), .Y(new_n6362));
  or_6   g04014(.A(new_n6362), .B(new_n6339), .Y(new_n6363));
  nand_5 g04015(.A(new_n6363), .B(new_n6337), .Y(new_n6364));
  not_8  g04016(.A(new_n6347), .Y(new_n6365));
  nor_5  g04017(.A(new_n6365), .B(new_n6342), .Y(new_n6366));
  nor_5  g04018(.A(new_n6361), .B(new_n6348), .Y(new_n6367));
  nor_5  g04019(.A(new_n6367), .B(new_n6366), .Y(new_n6368));
  nand_5 g04020(.A(new_n6368), .B(new_n6364), .Y(new_n6369));
  not_8  g04021(.A(new_n6369), .Y(new_n6370));
  xnor_4 g04022(.A(new_n6368), .B(new_n6364), .Y(new_n6371));
  not_8  g04023(.A(pi056), .Y(new_n6372));
  not_8  g04024(.A(pi335), .Y(new_n6373));
  nand_5 g04025(.A(new_n6373), .B(new_n6372), .Y(new_n6374));
  not_8  g04026(.A(new_n6374), .Y(new_n6375));
  not_8  g04027(.A(new_n6343), .Y(new_n6376));
  nor_5  g04028(.A(new_n6346), .B(new_n6376), .Y(new_n6377));
  nor_5  g04029(.A(new_n6377), .B(new_n6375), .Y(new_n6378));
  not_8  g04030(.A(pi197), .Y(new_n6379));
  not_8  g04031(.A(pi490), .Y(new_n6380));
  nand_5 g04032(.A(new_n6380), .B(new_n6379), .Y(new_n6381));
  not_8  g04033(.A(new_n6381), .Y(new_n6382));
  not_8  g04034(.A(new_n6333), .Y(new_n6383));
  nor_5  g04035(.A(new_n6335), .B(new_n6383), .Y(new_n6384));
  nor_5  g04036(.A(new_n6384), .B(new_n6382), .Y(new_n6385));
  not_8  g04037(.A(new_n6385), .Y(new_n6386));
  xor_4  g04038(.A(new_n6386), .B(new_n6378), .Y(new_n6387));
  nand_5 g04039(.A(new_n5634), .B(pi110), .Y(new_n6388));
  nand_5 g04040(.A(new_n6388), .B(new_n6361), .Y(new_n6389));
  nand_5 g04041(.A(pi282), .B(new_n6352), .Y(new_n6390));
  nand_5 g04042(.A(new_n6390), .B(new_n6389), .Y(new_n6391));
  not_8  g04043(.A(new_n6391), .Y(new_n6392));
  xor_4  g04044(.A(new_n6392), .B(new_n6387), .Y(new_n6393));
  nor_5  g04045(.A(new_n6393), .B(new_n6371), .Y(new_n6394));
  nor_5  g04046(.A(new_n6394), .B(new_n6370), .Y(new_n6395));
  nand_5 g04047(.A(new_n6386), .B(new_n6378), .Y(new_n6396));
  nand_5 g04048(.A(new_n6392), .B(new_n6387), .Y(new_n6397));
  nand_5 g04049(.A(new_n6397), .B(new_n6396), .Y(new_n6398));
  nor_5  g04050(.A(new_n6398), .B(new_n6395), .Y(po0026));
  not_8  g04051(.A(pi007), .Y(new_n6400));
  xor_4  g04052(.A(pi251), .B(new_n6400), .Y(new_n6401));
  not_8  g04053(.A(pi184), .Y(new_n6402));
  nand_5 g04054(.A(pi669), .B(new_n6402), .Y(new_n6403));
  xor_4  g04055(.A(pi669), .B(new_n6402), .Y(new_n6404));
  not_8  g04056(.A(pi384), .Y(new_n6405));
  nand_5 g04057(.A(pi413), .B(new_n6405), .Y(new_n6406));
  not_8  g04058(.A(pi344), .Y(new_n6407));
  nand_5 g04059(.A(pi664), .B(new_n6407), .Y(new_n6408));
  not_8  g04060(.A(new_n6408), .Y(new_n6409));
  xor_4  g04061(.A(pi664), .B(new_n6407), .Y(new_n6410));
  not_8  g04062(.A(new_n6410), .Y(new_n6411));
  not_8  g04063(.A(pi322), .Y(new_n6412));
  nand_5 g04064(.A(pi360), .B(new_n6412), .Y(new_n6413));
  not_8  g04065(.A(pi085), .Y(new_n6414));
  nand_5 g04066(.A(pi674), .B(new_n6414), .Y(new_n6415));
  or_6   g04067(.A(pi360), .B(new_n6412), .Y(new_n6416));
  nand_5 g04068(.A(new_n6416), .B(new_n6415), .Y(new_n6417));
  nand_5 g04069(.A(new_n6417), .B(new_n6413), .Y(new_n6418));
  nor_5  g04070(.A(new_n6418), .B(new_n6411), .Y(new_n6419));
  nor_5  g04071(.A(new_n6419), .B(new_n6409), .Y(new_n6420));
  xor_4  g04072(.A(pi413), .B(pi384), .Y(new_n6421));
  or_6   g04073(.A(new_n6421), .B(new_n6420), .Y(new_n6422));
  nand_5 g04074(.A(new_n6422), .B(new_n6406), .Y(new_n6423));
  nand_5 g04075(.A(new_n6423), .B(new_n6404), .Y(new_n6424));
  nand_5 g04076(.A(new_n6424), .B(new_n6403), .Y(new_n6425));
  xor_4  g04077(.A(new_n6425), .B(new_n6401), .Y(new_n6426));
  not_8  g04078(.A(pi030), .Y(new_n6427));
  xor_4  g04079(.A(pi154), .B(new_n6427), .Y(new_n6428));
  not_8  g04080(.A(pi267), .Y(new_n6429));
  nand_5 g04081(.A(pi456), .B(new_n6429), .Y(new_n6430));
  xor_4  g04082(.A(pi456), .B(new_n6429), .Y(new_n6431));
  not_8  g04083(.A(pi312), .Y(new_n6432));
  nand_5 g04084(.A(new_n6432), .B(pi098), .Y(new_n6433));
  not_8  g04085(.A(pi471), .Y(new_n6434));
  nand_5 g04086(.A(new_n6434), .B(pi188), .Y(new_n6435));
  not_8  g04087(.A(new_n6435), .Y(new_n6436));
  not_8  g04088(.A(pi188), .Y(new_n6437));
  xor_4  g04089(.A(pi471), .B(new_n6437), .Y(new_n6438));
  not_8  g04090(.A(new_n6438), .Y(new_n6439));
  not_8  g04091(.A(pi487), .Y(new_n6440));
  nand_5 g04092(.A(pi640), .B(new_n6440), .Y(new_n6441));
  not_8  g04093(.A(pi284), .Y(new_n6442));
  nand_5 g04094(.A(new_n6442), .B(pi156), .Y(new_n6443));
  not_8  g04095(.A(pi640), .Y(new_n6444));
  nand_5 g04096(.A(new_n6444), .B(pi487), .Y(new_n6445));
  nand_5 g04097(.A(new_n6445), .B(new_n6443), .Y(new_n6446));
  nand_5 g04098(.A(new_n6446), .B(new_n6441), .Y(new_n6447));
  nor_5  g04099(.A(new_n6447), .B(new_n6439), .Y(new_n6448));
  nor_5  g04100(.A(new_n6448), .B(new_n6436), .Y(new_n6449));
  xor_4  g04101(.A(pi312), .B(pi098), .Y(new_n6450));
  or_6   g04102(.A(new_n6450), .B(new_n6449), .Y(new_n6451));
  nand_5 g04103(.A(new_n6451), .B(new_n6433), .Y(new_n6452));
  nand_5 g04104(.A(new_n6452), .B(new_n6431), .Y(new_n6453));
  nand_5 g04105(.A(new_n6453), .B(new_n6430), .Y(new_n6454));
  xor_4  g04106(.A(new_n6454), .B(new_n6428), .Y(new_n6455));
  xor_4  g04107(.A(new_n6455), .B(new_n6426), .Y(new_n6456));
  xor_4  g04108(.A(new_n6423), .B(new_n6404), .Y(new_n6457));
  xor_4  g04109(.A(new_n6452), .B(new_n6431), .Y(new_n6458));
  nor_5  g04110(.A(new_n6458), .B(new_n6457), .Y(new_n6459));
  xor_4  g04111(.A(new_n6458), .B(new_n6457), .Y(new_n6460));
  not_8  g04112(.A(new_n6460), .Y(new_n6461));
  xor_4  g04113(.A(new_n6421), .B(new_n6420), .Y(new_n6462));
  xor_4  g04114(.A(new_n6450), .B(new_n6449), .Y(new_n6463));
  nor_5  g04115(.A(new_n6463), .B(new_n6462), .Y(new_n6464));
  xor_4  g04116(.A(new_n6463), .B(new_n6462), .Y(new_n6465));
  not_8  g04117(.A(new_n6465), .Y(new_n6466));
  xor_4  g04118(.A(new_n6418), .B(new_n6411), .Y(new_n6467));
  not_8  g04119(.A(new_n6467), .Y(new_n6468));
  xor_4  g04120(.A(new_n6447), .B(new_n6438), .Y(new_n6469));
  or_6   g04121(.A(new_n6469), .B(new_n6468), .Y(new_n6470));
  xor_4  g04122(.A(new_n6469), .B(new_n6468), .Y(new_n6471));
  not_8  g04123(.A(pi156), .Y(new_n6472));
  nand_5 g04124(.A(pi284), .B(new_n6472), .Y(new_n6473));
  nor_5  g04125(.A(pi674), .B(new_n6414), .Y(new_n6474));
  not_8  g04126(.A(new_n6474), .Y(new_n6475));
  nand_5 g04127(.A(new_n6475), .B(new_n6415), .Y(new_n6476));
  nand_5 g04128(.A(new_n6473), .B(new_n6443), .Y(new_n6477));
  not_8  g04129(.A(new_n6477), .Y(new_n6478));
  nand_5 g04130(.A(new_n6478), .B(new_n6476), .Y(new_n6479));
  nand_5 g04131(.A(new_n6479), .B(new_n6443), .Y(new_n6480));
  nand_5 g04132(.A(new_n6480), .B(new_n6475), .Y(new_n6481));
  not_8  g04133(.A(new_n6473), .Y(new_n6482));
  nand_5 g04134(.A(new_n6474), .B(new_n6482), .Y(new_n6483));
  nand_5 g04135(.A(new_n6483), .B(new_n6481), .Y(new_n6484));
  nand_5 g04136(.A(new_n6416), .B(new_n6413), .Y(new_n6485));
  nand_5 g04137(.A(new_n6445), .B(new_n6441), .Y(new_n6486));
  xor_4  g04138(.A(new_n6486), .B(new_n6485), .Y(new_n6487));
  xor_4  g04139(.A(new_n6487), .B(new_n6484), .Y(new_n6488));
  nor_5  g04140(.A(new_n6488), .B(new_n6473), .Y(new_n6489));
  not_8  g04141(.A(new_n6486), .Y(new_n6490));
  nand_5 g04142(.A(new_n6490), .B(new_n6443), .Y(new_n6491));
  or_6   g04143(.A(new_n6491), .B(new_n6489), .Y(new_n6492));
  nand_5 g04144(.A(new_n6486), .B(new_n6485), .Y(new_n6493));
  nor_5  g04145(.A(new_n6493), .B(new_n6481), .Y(new_n6494));
  nor_5  g04146(.A(new_n6482), .B(pi674), .Y(new_n6495));
  nand_5 g04147(.A(new_n6495), .B(new_n6486), .Y(new_n6496));
  and_6  g04148(.A(new_n6496), .B(new_n6476), .Y(new_n6497));
  nor_5  g04149(.A(new_n6497), .B(new_n6485), .Y(new_n6498));
  nor_5  g04150(.A(new_n6498), .B(new_n6494), .Y(new_n6499));
  nand_5 g04151(.A(new_n6499), .B(new_n6492), .Y(new_n6500));
  nand_5 g04152(.A(new_n6500), .B(new_n6471), .Y(new_n6501));
  nand_5 g04153(.A(new_n6501), .B(new_n6470), .Y(new_n6502));
  nor_5  g04154(.A(new_n6502), .B(new_n6466), .Y(new_n6503));
  nor_5  g04155(.A(new_n6503), .B(new_n6464), .Y(new_n6504));
  nor_5  g04156(.A(new_n6504), .B(new_n6461), .Y(new_n6505));
  or_6   g04157(.A(new_n6505), .B(new_n6459), .Y(new_n6506));
  xor_4  g04158(.A(new_n6506), .B(new_n6456), .Y(new_n6507));
  xor_4  g04159(.A(new_n6504), .B(new_n6461), .Y(new_n6508));
  not_8  g04160(.A(new_n6508), .Y(new_n6509));
  xor_4  g04161(.A(new_n6502), .B(new_n6465), .Y(new_n6510));
  xor_4  g04162(.A(new_n6478), .B(new_n6476), .Y(new_n6511));
  nand_5 g04163(.A(new_n6511), .B(new_n4567), .Y(new_n6512));
  not_8  g04164(.A(new_n6511), .Y(new_n6513));
  nand_5 g04165(.A(new_n6513), .B(new_n4595), .Y(new_n6514));
  nand_5 g04166(.A(new_n6514), .B(new_n6512), .Y(new_n6515));
  xnor_4 g04167(.A(new_n6515), .B(new_n4592), .Y(new_n6516));
  or_6   g04168(.A(new_n6516), .B(new_n6488), .Y(new_n6517));
  nand_5 g04169(.A(new_n6513), .B(new_n4598), .Y(new_n6518));
  nand_5 g04170(.A(new_n6518), .B(new_n6516), .Y(new_n6519));
  nand_5 g04171(.A(new_n6519), .B(new_n6517), .Y(new_n6520));
  nand_5 g04172(.A(new_n6520), .B(new_n4586), .Y(new_n6521));
  xnor_4 g04173(.A(new_n6500), .B(new_n6471), .Y(new_n6522));
  xor_4  g04174(.A(new_n6520), .B(new_n4585), .Y(new_n6523));
  or_6   g04175(.A(new_n6523), .B(new_n6522), .Y(new_n6524));
  nand_5 g04176(.A(new_n6524), .B(new_n6521), .Y(new_n6525));
  nand_5 g04177(.A(new_n6525), .B(new_n6510), .Y(new_n6526));
  xnor_4 g04178(.A(new_n6525), .B(new_n6510), .Y(new_n6527));
  or_6   g04179(.A(new_n6527), .B(new_n4579), .Y(new_n6528));
  nand_5 g04180(.A(new_n6528), .B(new_n6526), .Y(new_n6529));
  nand_5 g04181(.A(new_n6529), .B(new_n6509), .Y(new_n6530));
  not_8  g04182(.A(new_n6530), .Y(new_n6531));
  xor_4  g04183(.A(new_n6529), .B(new_n6508), .Y(new_n6532));
  nor_5  g04184(.A(new_n6532), .B(new_n4699), .Y(new_n6533));
  nor_5  g04185(.A(new_n6533), .B(new_n6531), .Y(new_n6534));
  nand_5 g04186(.A(new_n6534), .B(new_n6507), .Y(new_n6535));
  not_8  g04187(.A(new_n6507), .Y(new_n6536));
  xor_4  g04188(.A(new_n6534), .B(new_n6536), .Y(new_n6537));
  or_6   g04189(.A(new_n6537), .B(new_n4695), .Y(new_n6538));
  nand_5 g04190(.A(new_n6538), .B(new_n6535), .Y(new_n6539));
  not_8  g04191(.A(pi560), .Y(new_n6540));
  xor_4  g04192(.A(pi603), .B(new_n6540), .Y(new_n6541));
  nand_5 g04193(.A(new_n4693), .B(new_n4690), .Y(new_n6542));
  nand_5 g04194(.A(new_n6542), .B(new_n4692), .Y(new_n6543));
  xor_4  g04195(.A(new_n6543), .B(new_n6541), .Y(new_n6544));
  not_8  g04196(.A(new_n6544), .Y(new_n6545));
  nand_5 g04197(.A(pi251), .B(new_n6400), .Y(new_n6546));
  nand_5 g04198(.A(new_n6425), .B(new_n6401), .Y(new_n6547));
  nand_5 g04199(.A(new_n6547), .B(new_n6546), .Y(new_n6548));
  not_8  g04200(.A(pi256), .Y(new_n6549));
  or_6   g04201(.A(pi519), .B(new_n6549), .Y(new_n6550));
  nand_5 g04202(.A(pi519), .B(new_n6549), .Y(new_n6551));
  nand_5 g04203(.A(new_n6551), .B(new_n6550), .Y(new_n6552));
  xnor_4 g04204(.A(new_n6552), .B(new_n6548), .Y(new_n6553));
  not_8  g04205(.A(pi053), .Y(new_n6554));
  xor_4  g04206(.A(pi517), .B(new_n6554), .Y(new_n6555));
  not_8  g04207(.A(pi154), .Y(new_n6556));
  nand_5 g04208(.A(new_n6556), .B(pi030), .Y(new_n6557));
  nand_5 g04209(.A(new_n6454), .B(new_n6428), .Y(new_n6558));
  nand_5 g04210(.A(new_n6558), .B(new_n6557), .Y(new_n6559));
  xor_4  g04211(.A(new_n6559), .B(new_n6555), .Y(new_n6560));
  xor_4  g04212(.A(new_n6560), .B(new_n6553), .Y(new_n6561));
  or_6   g04213(.A(new_n6455), .B(new_n6426), .Y(new_n6562));
  nand_5 g04214(.A(new_n6506), .B(new_n6456), .Y(new_n6563));
  nand_5 g04215(.A(new_n6563), .B(new_n6562), .Y(new_n6564));
  xor_4  g04216(.A(new_n6564), .B(new_n6561), .Y(new_n6565));
  xor_4  g04217(.A(new_n6565), .B(new_n6545), .Y(new_n6566));
  xor_4  g04218(.A(new_n6566), .B(new_n6539), .Y(po0027));
  not_8  g04219(.A(pi318), .Y(new_n6568));
  xor_4  g04220(.A(pi448), .B(new_n6568), .Y(new_n6569));
  xor_4  g04221(.A(new_n6569), .B(pi799), .Y(new_n6570));
  xor_4  g04222(.A(new_n6570), .B(new_n5787), .Y(po0028));
  nor_5  g04223(.A(pi475), .B(pi388), .Y(new_n6572));
  nand_5 g04224(.A(pi797), .B(pi161), .Y(new_n6573));
  not_8  g04225(.A(new_n6573), .Y(new_n6574));
  not_8  g04226(.A(pi388), .Y(new_n6575));
  xor_4  g04227(.A(pi475), .B(new_n6575), .Y(new_n6576));
  nor_5  g04228(.A(new_n6576), .B(new_n6574), .Y(new_n6577));
  nor_5  g04229(.A(new_n6577), .B(new_n6572), .Y(new_n6578));
  not_8  g04230(.A(pi353), .Y(new_n6579));
  xor_4  g04231(.A(pi545), .B(new_n6579), .Y(new_n6580));
  xnor_4 g04232(.A(new_n6580), .B(new_n6578), .Y(new_n6581));
  xor_4  g04233(.A(new_n6581), .B(pi618), .Y(new_n6582));
  xor_4  g04234(.A(new_n6576), .B(new_n6573), .Y(new_n6583));
  nand_5 g04235(.A(new_n6583), .B(pi192), .Y(new_n6584));
  xor_4  g04236(.A(new_n6583), .B(pi192), .Y(new_n6585));
  xor_4  g04237(.A(pi797), .B(pi161), .Y(new_n6586));
  nor_5  g04238(.A(new_n6586), .B(pi813), .Y(new_n6587));
  nor_5  g04239(.A(pi751), .B(pi049), .Y(new_n6588));
  nor_5  g04240(.A(new_n5763), .B(pi281), .Y(new_n6589));
  nor_5  g04241(.A(new_n6589), .B(new_n6588), .Y(new_n6590));
  xnor_4 g04242(.A(new_n6586), .B(pi813), .Y(new_n6591));
  nor_5  g04243(.A(new_n6591), .B(new_n6590), .Y(new_n6592));
  nor_5  g04244(.A(new_n6592), .B(new_n6587), .Y(new_n6593));
  nand_5 g04245(.A(new_n6593), .B(new_n6585), .Y(new_n6594));
  nand_5 g04246(.A(new_n6594), .B(new_n6584), .Y(new_n6595));
  xor_4  g04247(.A(new_n6595), .B(new_n6582), .Y(new_n6596));
  xor_4  g04248(.A(new_n6593), .B(new_n6585), .Y(new_n6597));
  xor_4  g04249(.A(new_n6591), .B(new_n6590), .Y(new_n6598));
  nor_5  g04250(.A(pi781), .B(pi000), .Y(new_n6599));
  nand_5 g04251(.A(pi781), .B(pi000), .Y(new_n6600));
  not_8  g04252(.A(new_n6600), .Y(new_n6601));
  or_6   g04253(.A(new_n6601), .B(new_n6599), .Y(new_n6602));
  nor_5  g04254(.A(new_n6602), .B(pi482), .Y(new_n6603));
  nor_5  g04255(.A(new_n6603), .B(new_n6599), .Y(new_n6604));
  xor_4  g04256(.A(pi480), .B(pi422), .Y(new_n6605));
  xor_4  g04257(.A(new_n6605), .B(new_n4770), .Y(new_n6606));
  xor_4  g04258(.A(new_n6606), .B(new_n6604), .Y(new_n6607));
  not_8  g04259(.A(new_n6607), .Y(new_n6608));
  or_6   g04260(.A(new_n6608), .B(new_n6598), .Y(new_n6609));
  xor_4  g04261(.A(new_n5763), .B(pi281), .Y(new_n6610));
  not_8  g04262(.A(new_n6610), .Y(new_n6611));
  xor_4  g04263(.A(new_n6602), .B(pi482), .Y(new_n6612));
  or_6   g04264(.A(new_n6612), .B(new_n6611), .Y(new_n6613));
  xor_4  g04265(.A(new_n6608), .B(new_n6598), .Y(new_n6614));
  nand_5 g04266(.A(new_n6614), .B(new_n6613), .Y(new_n6615));
  nand_5 g04267(.A(new_n6615), .B(new_n6609), .Y(new_n6616));
  nor_5  g04268(.A(new_n6616), .B(new_n6597), .Y(new_n6617));
  xor_4  g04269(.A(pi495), .B(pi090), .Y(new_n6618));
  nor_5  g04270(.A(pi480), .B(pi422), .Y(new_n6619));
  and_6  g04271(.A(new_n6605), .B(new_n6600), .Y(new_n6620));
  nor_5  g04272(.A(new_n6620), .B(new_n6619), .Y(new_n6621));
  xor_4  g04273(.A(new_n6621), .B(new_n6618), .Y(new_n6622));
  nor_5  g04274(.A(new_n6606), .B(new_n6604), .Y(new_n6623));
  nor_5  g04275(.A(new_n6605), .B(new_n4770), .Y(new_n6624));
  nor_5  g04276(.A(new_n6620), .B(new_n6624), .Y(new_n6625));
  nor_5  g04277(.A(new_n6625), .B(new_n6623), .Y(new_n6626));
  xor_4  g04278(.A(new_n6626), .B(pi599), .Y(new_n6627));
  xor_4  g04279(.A(new_n6627), .B(new_n6622), .Y(new_n6628));
  not_8  g04280(.A(new_n6628), .Y(new_n6629));
  not_8  g04281(.A(new_n6597), .Y(new_n6630));
  xor_4  g04282(.A(new_n6616), .B(new_n6630), .Y(new_n6631));
  nor_5  g04283(.A(new_n6631), .B(new_n6629), .Y(new_n6632));
  or_6   g04284(.A(new_n6632), .B(new_n6617), .Y(new_n6633));
  xor_4  g04285(.A(new_n6633), .B(new_n6596), .Y(new_n6634));
  xor_4  g04286(.A(pi795), .B(pi343), .Y(new_n6635));
  nor_5  g04287(.A(pi495), .B(pi090), .Y(new_n6636));
  not_8  g04288(.A(new_n6618), .Y(new_n6637));
  nor_5  g04289(.A(new_n6621), .B(new_n6637), .Y(new_n6638));
  nor_5  g04290(.A(new_n6638), .B(new_n6636), .Y(new_n6639));
  xor_4  g04291(.A(new_n6639), .B(new_n6635), .Y(new_n6640));
  nand_5 g04292(.A(new_n6626), .B(pi599), .Y(new_n6641));
  nand_5 g04293(.A(new_n6627), .B(new_n6622), .Y(new_n6642));
  nand_5 g04294(.A(new_n6642), .B(new_n6641), .Y(new_n6643));
  or_6   g04295(.A(new_n6643), .B(new_n6640), .Y(new_n6644));
  nand_5 g04296(.A(new_n6643), .B(new_n6640), .Y(new_n6645));
  and_6  g04297(.A(new_n6645), .B(new_n6644), .Y(new_n6646));
  xor_4  g04298(.A(new_n6646), .B(new_n4763), .Y(new_n6647));
  not_8  g04299(.A(new_n6647), .Y(new_n6648));
  xor_4  g04300(.A(new_n6648), .B(new_n6634), .Y(po0029));
  nand_5 g04301(.A(new_n2450), .B(new_n5654), .Y(new_n6650));
  not_8  g04302(.A(pi638), .Y(new_n6651));
  xor_4  g04303(.A(new_n2394), .B(new_n6651), .Y(new_n6652));
  nor_5  g04304(.A(new_n2520), .B(pi393), .Y(new_n6653));
  nor_5  g04305(.A(new_n6653), .B(new_n2424), .Y(new_n6654));
  nand_5 g04306(.A(new_n6654), .B(new_n6652), .Y(new_n6655));
  nor_5  g04307(.A(new_n2394), .B(new_n6651), .Y(new_n6656));
  nor_5  g04308(.A(new_n6656), .B(new_n2397), .Y(new_n6657));
  nand_5 g04309(.A(new_n6657), .B(new_n6655), .Y(new_n6658));
  nand_5 g04310(.A(new_n6658), .B(pi391), .Y(new_n6659));
  xor_4  g04311(.A(new_n6658), .B(pi391), .Y(new_n6660));
  nand_5 g04312(.A(new_n6660), .B(new_n2416), .Y(new_n6661));
  nand_5 g04313(.A(new_n6661), .B(new_n6659), .Y(new_n6662));
  xor_4  g04314(.A(new_n2450), .B(pi252), .Y(new_n6663));
  or_6   g04315(.A(new_n6663), .B(new_n6662), .Y(new_n6664));
  nand_5 g04316(.A(new_n6664), .B(new_n6650), .Y(new_n6665));
  xor_4  g04317(.A(new_n2453), .B(pi242), .Y(new_n6666));
  xor_4  g04318(.A(new_n6666), .B(new_n6665), .Y(new_n6667));
  xor_4  g04319(.A(new_n6663), .B(new_n6662), .Y(new_n6668));
  xor_4  g04320(.A(new_n2520), .B(pi393), .Y(new_n6669));
  nand_5 g04321(.A(new_n6669), .B(pi077), .Y(new_n6670));
  nor_5  g04322(.A(new_n6670), .B(new_n2484), .Y(new_n6671));
  xor_4  g04323(.A(new_n6654), .B(new_n6652), .Y(new_n6672));
  xor_4  g04324(.A(new_n6670), .B(new_n2484), .Y(new_n6673));
  not_8  g04325(.A(new_n6673), .Y(new_n6674));
  nor_5  g04326(.A(new_n6674), .B(new_n6672), .Y(new_n6675));
  or_6   g04327(.A(new_n6675), .B(new_n6671), .Y(new_n6676));
  nand_5 g04328(.A(new_n6676), .B(pi501), .Y(new_n6677));
  xor_4  g04329(.A(new_n6660), .B(new_n2415), .Y(new_n6678));
  not_8  g04330(.A(new_n6678), .Y(new_n6679));
  xor_4  g04331(.A(new_n6676), .B(new_n2480), .Y(new_n6680));
  or_6   g04332(.A(new_n6680), .B(new_n6679), .Y(new_n6681));
  nand_5 g04333(.A(new_n6681), .B(new_n6677), .Y(new_n6682));
  nor_5  g04334(.A(new_n6682), .B(new_n6668), .Y(new_n6683));
  not_8  g04335(.A(new_n6668), .Y(new_n6684));
  xor_4  g04336(.A(new_n6682), .B(new_n6684), .Y(new_n6685));
  nor_5  g04337(.A(new_n6685), .B(pi831), .Y(new_n6686));
  or_6   g04338(.A(new_n6686), .B(new_n6683), .Y(new_n6687));
  nand_5 g04339(.A(new_n6687), .B(new_n6667), .Y(new_n6688));
  or_6   g04340(.A(new_n6687), .B(new_n6667), .Y(new_n6689));
  nand_5 g04341(.A(new_n6689), .B(new_n6688), .Y(new_n6690));
  xor_4  g04342(.A(new_n6690), .B(pi662), .Y(new_n6691));
  xor_4  g04343(.A(new_n6685), .B(pi831), .Y(new_n6692));
  xor_4  g04344(.A(new_n6669), .B(pi077), .Y(new_n6693));
  nor_5  g04345(.A(new_n6693), .B(new_n3342), .Y(new_n6694));
  nor_5  g04346(.A(new_n6694), .B(new_n3347), .Y(new_n6695));
  not_8  g04347(.A(new_n3350), .Y(new_n6696));
  nor_5  g04348(.A(new_n6693), .B(new_n6696), .Y(new_n6697));
  or_6   g04349(.A(new_n6697), .B(new_n6695), .Y(new_n6698));
  xor_4  g04350(.A(new_n6673), .B(new_n6672), .Y(new_n6699));
  nor_5  g04351(.A(new_n6699), .B(new_n6698), .Y(new_n6700));
  nor_5  g04352(.A(new_n6700), .B(new_n6695), .Y(new_n6701));
  or_6   g04353(.A(new_n6701), .B(new_n3357), .Y(new_n6702));
  xor_4  g04354(.A(new_n6680), .B(new_n6678), .Y(new_n6703));
  xor_4  g04355(.A(new_n6701), .B(new_n3358), .Y(new_n6704));
  or_6   g04356(.A(new_n6704), .B(new_n6703), .Y(new_n6705));
  nand_5 g04357(.A(new_n6705), .B(new_n6702), .Y(new_n6706));
  not_8  g04358(.A(new_n6706), .Y(new_n6707));
  nor_5  g04359(.A(new_n6707), .B(new_n6692), .Y(new_n6708));
  and_6  g04360(.A(new_n6707), .B(new_n6692), .Y(new_n6709));
  nor_5  g04361(.A(new_n6709), .B(new_n3367), .Y(new_n6710));
  nor_5  g04362(.A(new_n6710), .B(new_n6708), .Y(new_n6711));
  xnor_4 g04363(.A(new_n6711), .B(new_n6691), .Y(new_n6712));
  xor_4  g04364(.A(new_n6712), .B(new_n3337), .Y(po0030));
  not_8  g04365(.A(pi022), .Y(new_n6714));
  xor_4  g04366(.A(pi395), .B(new_n6714), .Y(new_n6715));
  not_8  g04367(.A(pi615), .Y(new_n6716));
  nand_5 g04368(.A(new_n6716), .B(new_n4045), .Y(new_n6717));
  nand_5 g04369(.A(pi615), .B(pi351), .Y(new_n6718));
  not_8  g04370(.A(pi579), .Y(new_n6719));
  nand_5 g04371(.A(new_n6719), .B(new_n3895), .Y(new_n6720));
  xor_4  g04372(.A(pi579), .B(new_n3895), .Y(new_n6721));
  not_8  g04373(.A(new_n6721), .Y(new_n6722));
  not_8  g04374(.A(pi483), .Y(new_n6723));
  nand_5 g04375(.A(new_n3897), .B(new_n6723), .Y(new_n6724));
  nand_5 g04376(.A(pi506), .B(pi483), .Y(new_n6725));
  not_8  g04377(.A(pi264), .Y(new_n6726));
  nand_5 g04378(.A(new_n3900), .B(new_n6726), .Y(new_n6727));
  nand_5 g04379(.A(pi374), .B(pi264), .Y(new_n6728));
  nand_5 g04380(.A(pi569), .B(pi445), .Y(new_n6729));
  nand_5 g04381(.A(pi688), .B(pi333), .Y(new_n6730));
  nand_5 g04382(.A(new_n6730), .B(new_n6729), .Y(new_n6731));
  not_8  g04383(.A(pi333), .Y(new_n6732));
  nand_5 g04384(.A(new_n3905), .B(new_n6732), .Y(new_n6733));
  nand_5 g04385(.A(new_n6733), .B(new_n6731), .Y(new_n6734));
  nand_5 g04386(.A(new_n6734), .B(new_n6728), .Y(new_n6735));
  nand_5 g04387(.A(new_n6735), .B(new_n6727), .Y(new_n6736));
  nand_5 g04388(.A(new_n6736), .B(new_n6725), .Y(new_n6737));
  nand_5 g04389(.A(new_n6737), .B(new_n6724), .Y(new_n6738));
  nand_5 g04390(.A(new_n6738), .B(new_n6722), .Y(new_n6739));
  nand_5 g04391(.A(new_n6739), .B(new_n6720), .Y(new_n6740));
  nand_5 g04392(.A(new_n6740), .B(new_n6718), .Y(new_n6741));
  nand_5 g04393(.A(new_n6741), .B(new_n6717), .Y(new_n6742));
  xnor_4 g04394(.A(new_n6742), .B(new_n6715), .Y(new_n6743));
  nand_5 g04395(.A(new_n6743), .B(new_n5460), .Y(new_n6744));
  xor_4  g04396(.A(new_n6743), .B(new_n5460), .Y(new_n6745));
  nand_5 g04397(.A(new_n6718), .B(new_n6717), .Y(new_n6746));
  xor_4  g04398(.A(new_n6746), .B(new_n6740), .Y(new_n6747));
  or_6   g04399(.A(new_n6747), .B(pi699), .Y(new_n6748));
  not_8  g04400(.A(new_n6748), .Y(new_n6749));
  xor_4  g04401(.A(new_n6747), .B(pi699), .Y(new_n6750));
  not_8  g04402(.A(new_n6750), .Y(new_n6751));
  xor_4  g04403(.A(new_n6738), .B(new_n6721), .Y(new_n6752));
  not_8  g04404(.A(new_n6752), .Y(new_n6753));
  nand_5 g04405(.A(new_n6753), .B(new_n2405), .Y(new_n6754));
  not_8  g04406(.A(new_n6754), .Y(new_n6755));
  xor_4  g04407(.A(new_n6752), .B(new_n2405), .Y(new_n6756));
  nand_5 g04408(.A(new_n6725), .B(new_n6724), .Y(new_n6757));
  xor_4  g04409(.A(new_n6757), .B(new_n6736), .Y(new_n6758));
  nand_5 g04410(.A(new_n6758), .B(pi289), .Y(new_n6759));
  or_6   g04411(.A(new_n6758), .B(pi289), .Y(new_n6760));
  nand_5 g04412(.A(new_n6728), .B(new_n6727), .Y(new_n6761));
  xor_4  g04413(.A(new_n6761), .B(new_n6734), .Y(new_n6762));
  nand_5 g04414(.A(new_n6762), .B(pi486), .Y(new_n6763));
  or_6   g04415(.A(new_n6762), .B(pi486), .Y(new_n6764));
  nand_5 g04416(.A(new_n6733), .B(new_n6730), .Y(new_n6765));
  not_8  g04417(.A(pi569), .Y(new_n6766));
  nand_5 g04418(.A(new_n6766), .B(new_n2565), .Y(new_n6767));
  nand_5 g04419(.A(new_n6767), .B(pi223), .Y(new_n6768));
  nand_5 g04420(.A(new_n6768), .B(new_n6729), .Y(new_n6769));
  xor_4  g04421(.A(new_n6769), .B(new_n6765), .Y(new_n6770));
  or_6   g04422(.A(new_n6770), .B(new_n2392), .Y(new_n6771));
  not_8  g04423(.A(new_n6729), .Y(new_n6772));
  nor_5  g04424(.A(new_n6765), .B(new_n6772), .Y(new_n6773));
  nand_5 g04425(.A(new_n6773), .B(new_n6769), .Y(new_n6774));
  nand_5 g04426(.A(new_n6774), .B(new_n6771), .Y(new_n6775));
  nand_5 g04427(.A(new_n6775), .B(new_n6764), .Y(new_n6776));
  nand_5 g04428(.A(new_n6776), .B(new_n6763), .Y(new_n6777));
  nand_5 g04429(.A(new_n6777), .B(new_n6760), .Y(new_n6778));
  nand_5 g04430(.A(new_n6778), .B(new_n6759), .Y(new_n6779));
  nor_5  g04431(.A(new_n6779), .B(new_n6756), .Y(new_n6780));
  nor_5  g04432(.A(new_n6780), .B(new_n6755), .Y(new_n6781));
  nor_5  g04433(.A(new_n6781), .B(new_n6751), .Y(new_n6782));
  nor_5  g04434(.A(new_n6782), .B(new_n6749), .Y(new_n6783));
  not_8  g04435(.A(new_n6783), .Y(new_n6784));
  nand_5 g04436(.A(new_n6784), .B(new_n6745), .Y(new_n6785));
  nand_5 g04437(.A(new_n6785), .B(new_n6744), .Y(new_n6786));
  not_8  g04438(.A(pi073), .Y(new_n6787));
  xor_4  g04439(.A(pi734), .B(new_n6787), .Y(new_n6788));
  nor_5  g04440(.A(new_n4266), .B(new_n6714), .Y(new_n6789));
  nor_5  g04441(.A(new_n6742), .B(new_n6715), .Y(new_n6790));
  nor_5  g04442(.A(new_n6790), .B(new_n6789), .Y(new_n6791));
  xor_4  g04443(.A(new_n6791), .B(new_n6788), .Y(new_n6792));
  or_6   g04444(.A(new_n6792), .B(pi319), .Y(new_n6793));
  nand_5 g04445(.A(new_n6792), .B(pi319), .Y(new_n6794));
  and_6  g04446(.A(new_n6794), .B(new_n6793), .Y(new_n6795));
  xor_4  g04447(.A(new_n6795), .B(new_n6786), .Y(new_n6796));
  not_8  g04448(.A(new_n6796), .Y(new_n6797));
  nand_5 g04449(.A(pi297), .B(pi033), .Y(new_n6798));
  not_8  g04450(.A(pi033), .Y(new_n6799));
  nand_5 g04451(.A(new_n5644), .B(new_n6799), .Y(new_n6800));
  nand_5 g04452(.A(pi613), .B(pi572), .Y(new_n6801));
  not_8  g04453(.A(pi572), .Y(new_n6802));
  nand_5 g04454(.A(new_n5646), .B(new_n6802), .Y(new_n6803));
  nand_5 g04455(.A(pi587), .B(pi250), .Y(new_n6804));
  nand_5 g04456(.A(pi779), .B(pi338), .Y(new_n6805));
  not_8  g04457(.A(new_n6805), .Y(new_n6806));
  xor_4  g04458(.A(pi779), .B(pi338), .Y(new_n6807));
  not_8  g04459(.A(new_n6807), .Y(new_n6808));
  not_8  g04460(.A(pi760), .Y(new_n6809));
  nor_5  g04461(.A(new_n6809), .B(new_n3946), .Y(new_n6810));
  nor_5  g04462(.A(new_n4082), .B(new_n4081), .Y(new_n6811));
  nor_5  g04463(.A(new_n6811), .B(new_n6810), .Y(new_n6812));
  nor_5  g04464(.A(new_n6812), .B(new_n6808), .Y(new_n6813));
  nor_5  g04465(.A(new_n6813), .B(new_n6806), .Y(new_n6814));
  nor_5  g04466(.A(pi587), .B(pi250), .Y(new_n6815));
  or_6   g04467(.A(new_n6815), .B(new_n6814), .Y(new_n6816));
  nand_5 g04468(.A(new_n6816), .B(new_n6804), .Y(new_n6817));
  nand_5 g04469(.A(new_n6817), .B(new_n6803), .Y(new_n6818));
  nand_5 g04470(.A(new_n6818), .B(new_n6801), .Y(new_n6819));
  nand_5 g04471(.A(new_n6819), .B(new_n6800), .Y(new_n6820));
  nand_5 g04472(.A(new_n6820), .B(new_n6798), .Y(new_n6821));
  not_8  g04473(.A(new_n6821), .Y(new_n6822));
  nand_5 g04474(.A(pi834), .B(pi437), .Y(new_n6823));
  not_8  g04475(.A(pi437), .Y(new_n6824));
  nand_5 g04476(.A(new_n5640), .B(new_n6824), .Y(new_n6825));
  nand_5 g04477(.A(new_n6825), .B(new_n6823), .Y(new_n6826));
  xor_4  g04478(.A(new_n6826), .B(new_n6822), .Y(new_n6827));
  not_8  g04479(.A(new_n6827), .Y(new_n6828));
  not_8  g04480(.A(pi714), .Y(new_n6829));
  xor_4  g04481(.A(pi587), .B(pi250), .Y(new_n6830));
  xor_4  g04482(.A(new_n6830), .B(new_n6814), .Y(new_n6831));
  not_8  g04483(.A(new_n6831), .Y(new_n6832));
  nand_5 g04484(.A(new_n6832), .B(pi242), .Y(new_n6833));
  nand_5 g04485(.A(new_n6831), .B(new_n5651), .Y(new_n6834));
  xor_4  g04486(.A(new_n6812), .B(new_n6807), .Y(new_n6835));
  not_8  g04487(.A(pi391), .Y(new_n6836));
  xor_4  g04488(.A(new_n4079), .B(new_n4077), .Y(new_n6837));
  not_8  g04489(.A(new_n6837), .Y(new_n6838));
  nand_5 g04490(.A(new_n6838), .B(new_n6651), .Y(new_n6839));
  nand_5 g04491(.A(new_n6837), .B(pi638), .Y(new_n6840));
  nand_5 g04492(.A(new_n4118), .B(pi393), .Y(new_n6841));
  nand_5 g04493(.A(new_n6841), .B(new_n6840), .Y(new_n6842));
  nand_5 g04494(.A(new_n6842), .B(new_n6839), .Y(new_n6843));
  nand_5 g04495(.A(new_n6843), .B(new_n6836), .Y(new_n6844));
  xor_4  g04496(.A(new_n6843), .B(pi391), .Y(new_n6845));
  or_6   g04497(.A(new_n6845), .B(new_n4083), .Y(new_n6846));
  nand_5 g04498(.A(new_n6846), .B(new_n6844), .Y(new_n6847));
  or_6   g04499(.A(new_n6847), .B(new_n6835), .Y(new_n6848));
  xor_4  g04500(.A(new_n6847), .B(new_n6835), .Y(new_n6849));
  nand_5 g04501(.A(new_n6849), .B(pi252), .Y(new_n6850));
  nand_5 g04502(.A(new_n6850), .B(new_n6848), .Y(new_n6851));
  nand_5 g04503(.A(new_n6851), .B(new_n6834), .Y(new_n6852));
  nand_5 g04504(.A(new_n6852), .B(new_n6833), .Y(new_n6853));
  nor_5  g04505(.A(new_n6853), .B(pi539), .Y(new_n6854));
  and_6  g04506(.A(new_n6801), .B(new_n6803), .Y(new_n6855));
  xor_4  g04507(.A(new_n6855), .B(new_n6817), .Y(new_n6856));
  xor_4  g04508(.A(new_n6853), .B(new_n5648), .Y(new_n6857));
  nor_5  g04509(.A(new_n6857), .B(new_n6856), .Y(new_n6858));
  or_6   g04510(.A(new_n6858), .B(new_n6854), .Y(new_n6859));
  nand_5 g04511(.A(new_n6859), .B(new_n6829), .Y(new_n6860));
  nand_5 g04512(.A(new_n6798), .B(new_n6800), .Y(new_n6861));
  xor_4  g04513(.A(new_n6861), .B(new_n6819), .Y(new_n6862));
  xor_4  g04514(.A(new_n6859), .B(new_n6829), .Y(new_n6863));
  nand_5 g04515(.A(new_n6863), .B(new_n6862), .Y(new_n6864));
  nand_5 g04516(.A(new_n6864), .B(new_n6860), .Y(new_n6865));
  nand_5 g04517(.A(new_n6865), .B(new_n6828), .Y(new_n6866));
  or_6   g04518(.A(new_n6865), .B(new_n6828), .Y(new_n6867));
  nand_5 g04519(.A(new_n6867), .B(new_n6866), .Y(new_n6868));
  xor_4  g04520(.A(new_n6868), .B(pi377), .Y(new_n6869));
  nor_5  g04521(.A(new_n6869), .B(new_n6797), .Y(new_n6870));
  xor_4  g04522(.A(new_n6869), .B(new_n6797), .Y(new_n6871));
  xor_4  g04523(.A(new_n6783), .B(new_n6745), .Y(new_n6872));
  not_8  g04524(.A(new_n6872), .Y(new_n6873));
  not_8  g04525(.A(new_n6862), .Y(new_n6874));
  xor_4  g04526(.A(new_n6863), .B(new_n6874), .Y(new_n6875));
  nor_5  g04527(.A(new_n6875), .B(new_n6873), .Y(new_n6876));
  and_6  g04528(.A(new_n6875), .B(new_n6873), .Y(new_n6877));
  xor_4  g04529(.A(new_n6781), .B(new_n6750), .Y(new_n6878));
  xor_4  g04530(.A(new_n6857), .B(new_n6856), .Y(new_n6879));
  or_6   g04531(.A(new_n6879), .B(new_n6878), .Y(new_n6880));
  xor_4  g04532(.A(new_n6879), .B(new_n6878), .Y(new_n6881));
  xor_4  g04533(.A(new_n6779), .B(new_n6756), .Y(new_n6882));
  not_8  g04534(.A(new_n6882), .Y(new_n6883));
  nand_5 g04535(.A(new_n6834), .B(new_n6833), .Y(new_n6884));
  xor_4  g04536(.A(new_n6884), .B(new_n6851), .Y(new_n6885));
  or_6   g04537(.A(new_n6885), .B(new_n6883), .Y(new_n6886));
  xor_4  g04538(.A(new_n6885), .B(new_n6883), .Y(new_n6887));
  and_6  g04539(.A(new_n6760), .B(new_n6759), .Y(new_n6888));
  xor_4  g04540(.A(new_n6888), .B(new_n6777), .Y(new_n6889));
  xor_4  g04541(.A(new_n6849), .B(new_n5654), .Y(new_n6890));
  nand_5 g04542(.A(new_n6890), .B(new_n6889), .Y(new_n6891));
  nand_5 g04543(.A(new_n6764), .B(new_n6763), .Y(new_n6892));
  xor_4  g04544(.A(new_n6892), .B(new_n6775), .Y(new_n6893));
  not_8  g04545(.A(new_n4083), .Y(new_n6894));
  xor_4  g04546(.A(new_n6845), .B(new_n6894), .Y(new_n6895));
  nor_5  g04547(.A(new_n6895), .B(new_n6893), .Y(new_n6896));
  not_8  g04548(.A(new_n6893), .Y(new_n6897));
  xor_4  g04549(.A(new_n6895), .B(new_n6897), .Y(new_n6898));
  xor_4  g04550(.A(new_n6770), .B(new_n2392), .Y(new_n6899));
  not_8  g04551(.A(new_n6899), .Y(new_n6900));
  nand_5 g04552(.A(new_n6840), .B(new_n6839), .Y(new_n6901));
  xor_4  g04553(.A(new_n5593), .B(pi569), .Y(new_n6902));
  nand_5 g04554(.A(new_n6902), .B(new_n6841), .Y(new_n6903));
  not_8  g04555(.A(new_n6902), .Y(new_n6904));
  not_8  g04556(.A(new_n4118), .Y(new_n6905));
  nand_5 g04557(.A(new_n6905), .B(new_n5693), .Y(new_n6906));
  nand_5 g04558(.A(new_n6906), .B(new_n6904), .Y(new_n6907));
  nand_5 g04559(.A(new_n6907), .B(new_n6903), .Y(new_n6908));
  xor_4  g04560(.A(new_n6908), .B(new_n6901), .Y(new_n6909));
  nor_5  g04561(.A(new_n6909), .B(new_n6900), .Y(new_n6910));
  and_6  g04562(.A(new_n6906), .B(new_n6841), .Y(new_n6911));
  nor_5  g04563(.A(new_n6911), .B(new_n6902), .Y(new_n6912));
  and_6  g04564(.A(new_n6912), .B(new_n6909), .Y(new_n6913));
  nor_5  g04565(.A(new_n6913), .B(new_n6910), .Y(new_n6914));
  nor_5  g04566(.A(new_n6914), .B(new_n6898), .Y(new_n6915));
  nor_5  g04567(.A(new_n6915), .B(new_n6896), .Y(new_n6916));
  not_8  g04568(.A(new_n6889), .Y(new_n6917));
  xor_4  g04569(.A(new_n6890), .B(new_n6917), .Y(new_n6918));
  or_6   g04570(.A(new_n6918), .B(new_n6916), .Y(new_n6919));
  nand_5 g04571(.A(new_n6919), .B(new_n6891), .Y(new_n6920));
  not_8  g04572(.A(new_n6920), .Y(new_n6921));
  nand_5 g04573(.A(new_n6921), .B(new_n6887), .Y(new_n6922));
  nand_5 g04574(.A(new_n6922), .B(new_n6886), .Y(new_n6923));
  nand_5 g04575(.A(new_n6923), .B(new_n6881), .Y(new_n6924));
  nand_5 g04576(.A(new_n6924), .B(new_n6880), .Y(new_n6925));
  nor_5  g04577(.A(new_n6925), .B(new_n6877), .Y(new_n6926));
  nor_5  g04578(.A(new_n6926), .B(new_n6876), .Y(new_n6927));
  nand_5 g04579(.A(new_n6927), .B(new_n6871), .Y(new_n6928));
  not_8  g04580(.A(new_n6928), .Y(new_n6929));
  nor_5  g04581(.A(new_n6929), .B(new_n6870), .Y(new_n6930));
  xor_4  g04582(.A(pi784), .B(pi728), .Y(new_n6931));
  nor_5  g04583(.A(new_n4262), .B(new_n6787), .Y(new_n6932));
  nor_5  g04584(.A(new_n6791), .B(new_n6788), .Y(new_n6933));
  nor_5  g04585(.A(new_n6933), .B(new_n6932), .Y(new_n6934));
  xor_4  g04586(.A(new_n6934), .B(new_n6931), .Y(new_n6935));
  xor_4  g04587(.A(new_n6935), .B(pi777), .Y(new_n6936));
  nand_5 g04588(.A(new_n6794), .B(new_n6786), .Y(new_n6937));
  nand_5 g04589(.A(new_n6937), .B(new_n6793), .Y(new_n6938));
  xor_4  g04590(.A(new_n6938), .B(new_n6936), .Y(new_n6939));
  xor_4  g04591(.A(pi666), .B(pi472), .Y(new_n6940));
  nand_5 g04592(.A(new_n6825), .B(new_n6821), .Y(new_n6941));
  nand_5 g04593(.A(new_n6941), .B(new_n6823), .Y(new_n6942));
  xor_4  g04594(.A(new_n6942), .B(new_n6940), .Y(new_n6943));
  not_8  g04595(.A(new_n6943), .Y(new_n6944));
  nand_5 g04596(.A(new_n6867), .B(new_n5642), .Y(new_n6945));
  nand_5 g04597(.A(new_n6945), .B(new_n6866), .Y(new_n6946));
  xor_4  g04598(.A(new_n6946), .B(new_n6944), .Y(new_n6947));
  xor_4  g04599(.A(new_n6947), .B(pi533), .Y(new_n6948));
  xor_4  g04600(.A(new_n6948), .B(new_n6939), .Y(new_n6949));
  xor_4  g04601(.A(new_n6949), .B(new_n6930), .Y(po0031));
  not_8  g04602(.A(pi646), .Y(new_n6951));
  xor_4  g04603(.A(pi775), .B(new_n6951), .Y(new_n6952));
  not_8  g04604(.A(pi555), .Y(new_n6953));
  nand_5 g04605(.A(new_n6953), .B(pi139), .Y(new_n6954));
  not_8  g04606(.A(pi139), .Y(new_n6955));
  xor_4  g04607(.A(pi555), .B(new_n6955), .Y(new_n6956));
  not_8  g04608(.A(pi667), .Y(new_n6957));
  nand_5 g04609(.A(pi683), .B(new_n6957), .Y(new_n6958));
  xor_4  g04610(.A(pi683), .B(new_n6957), .Y(new_n6959));
  not_8  g04611(.A(pi566), .Y(new_n6960));
  nand_5 g04612(.A(pi567), .B(new_n6960), .Y(new_n6961));
  xor_4  g04613(.A(pi567), .B(new_n6960), .Y(new_n6962));
  not_8  g04614(.A(pi145), .Y(new_n6963));
  nand_5 g04615(.A(new_n6963), .B(pi088), .Y(new_n6964));
  xor_4  g04616(.A(pi145), .B(new_n2373), .Y(new_n6965));
  not_8  g04617(.A(pi454), .Y(new_n6966));
  nand_5 g04618(.A(pi605), .B(new_n6966), .Y(new_n6967));
  xor_4  g04619(.A(pi605), .B(new_n6966), .Y(new_n6968));
  not_8  g04620(.A(pi731), .Y(new_n6969));
  nand_5 g04621(.A(new_n6969), .B(pi434), .Y(new_n6970));
  xor_4  g04622(.A(pi731), .B(new_n2357), .Y(new_n6971));
  not_8  g04623(.A(pi270), .Y(new_n6972));
  nand_5 g04624(.A(pi552), .B(new_n6972), .Y(new_n6973));
  xor_4  g04625(.A(pi552), .B(new_n6972), .Y(new_n6974));
  not_8  g04626(.A(pi367), .Y(new_n6975));
  nand_5 g04627(.A(new_n6975), .B(pi190), .Y(new_n6976));
  not_8  g04628(.A(new_n6976), .Y(new_n6977));
  nand_5 g04629(.A(new_n6977), .B(new_n6974), .Y(new_n6978));
  nand_5 g04630(.A(new_n6978), .B(new_n6973), .Y(new_n6979));
  nand_5 g04631(.A(new_n6979), .B(new_n6971), .Y(new_n6980));
  nand_5 g04632(.A(new_n6980), .B(new_n6970), .Y(new_n6981));
  nand_5 g04633(.A(new_n6981), .B(new_n6968), .Y(new_n6982));
  nand_5 g04634(.A(new_n6982), .B(new_n6967), .Y(new_n6983));
  nand_5 g04635(.A(new_n6983), .B(new_n6965), .Y(new_n6984));
  nand_5 g04636(.A(new_n6984), .B(new_n6964), .Y(new_n6985));
  nand_5 g04637(.A(new_n6985), .B(new_n6962), .Y(new_n6986));
  nand_5 g04638(.A(new_n6986), .B(new_n6961), .Y(new_n6987));
  nand_5 g04639(.A(new_n6987), .B(new_n6959), .Y(new_n6988));
  nand_5 g04640(.A(new_n6988), .B(new_n6958), .Y(new_n6989));
  nand_5 g04641(.A(new_n6989), .B(new_n6956), .Y(new_n6990));
  nand_5 g04642(.A(new_n6990), .B(new_n6954), .Y(new_n6991));
  xor_4  g04643(.A(new_n6991), .B(new_n6952), .Y(new_n6992));
  xor_4  g04644(.A(pi507), .B(pi423), .Y(new_n6993));
  nand_5 g04645(.A(pi324), .B(pi071), .Y(new_n6994));
  nand_5 g04646(.A(new_n5180), .B(new_n5179), .Y(new_n6995));
  nand_5 g04647(.A(new_n6995), .B(new_n5182), .Y(new_n6996));
  not_8  g04648(.A(pi071), .Y(new_n6997));
  xor_4  g04649(.A(pi324), .B(new_n6997), .Y(new_n6998));
  or_6   g04650(.A(new_n6998), .B(new_n6996), .Y(new_n6999));
  nand_5 g04651(.A(new_n6999), .B(new_n6994), .Y(new_n7000));
  xor_4  g04652(.A(new_n7000), .B(new_n6993), .Y(new_n7001));
  nand_5 g04653(.A(pi738), .B(pi513), .Y(new_n7002));
  not_8  g04654(.A(new_n7002), .Y(new_n7003));
  xor_4  g04655(.A(pi738), .B(pi513), .Y(new_n7004));
  not_8  g04656(.A(new_n7004), .Y(new_n7005));
  nand_5 g04657(.A(pi657), .B(pi004), .Y(new_n7006));
  not_8  g04658(.A(new_n7006), .Y(new_n7007));
  xor_4  g04659(.A(pi657), .B(pi004), .Y(new_n7008));
  not_8  g04660(.A(new_n7008), .Y(new_n7009));
  not_8  g04661(.A(pi747), .Y(new_n7010));
  nand_5 g04662(.A(new_n7010), .B(new_n4705), .Y(new_n7011));
  nand_5 g04663(.A(pi747), .B(pi743), .Y(new_n7012));
  not_8  g04664(.A(pi078), .Y(new_n7013));
  nand_5 g04665(.A(new_n4669), .B(new_n7013), .Y(new_n7014));
  xor_4  g04666(.A(pi444), .B(pi078), .Y(new_n7015));
  not_8  g04667(.A(pi294), .Y(new_n7016));
  nand_5 g04668(.A(new_n7016), .B(new_n4641), .Y(new_n7017));
  nand_5 g04669(.A(pi294), .B(pi052), .Y(new_n7018));
  not_8  g04670(.A(pi337), .Y(new_n7019));
  nand_5 g04671(.A(new_n4623), .B(new_n7019), .Y(new_n7020));
  nand_5 g04672(.A(pi386), .B(pi337), .Y(new_n7021));
  nand_5 g04673(.A(pi574), .B(pi238), .Y(new_n7022));
  nand_5 g04674(.A(new_n7022), .B(new_n7021), .Y(new_n7023));
  nand_5 g04675(.A(new_n7023), .B(new_n7020), .Y(new_n7024));
  nand_5 g04676(.A(new_n7024), .B(new_n7018), .Y(new_n7025));
  nand_5 g04677(.A(new_n7025), .B(new_n7017), .Y(new_n7026));
  nand_5 g04678(.A(new_n7026), .B(new_n7015), .Y(new_n7027));
  nand_5 g04679(.A(new_n7027), .B(new_n7014), .Y(new_n7028));
  nand_5 g04680(.A(new_n7028), .B(new_n7012), .Y(new_n7029));
  nand_5 g04681(.A(new_n7029), .B(new_n7011), .Y(new_n7030));
  nor_5  g04682(.A(new_n7030), .B(new_n7009), .Y(new_n7031));
  nor_5  g04683(.A(new_n7031), .B(new_n7007), .Y(new_n7032));
  nor_5  g04684(.A(new_n7032), .B(new_n7005), .Y(new_n7033));
  nor_5  g04685(.A(new_n7033), .B(new_n7003), .Y(new_n7034));
  xor_4  g04686(.A(pi314), .B(pi180), .Y(new_n7035));
  xor_4  g04687(.A(new_n7035), .B(new_n7034), .Y(new_n7036));
  nand_5 g04688(.A(new_n7036), .B(new_n7001), .Y(new_n7037));
  xor_4  g04689(.A(new_n7036), .B(new_n7001), .Y(new_n7038));
  xnor_4 g04690(.A(new_n6998), .B(new_n6996), .Y(new_n7039));
  xor_4  g04691(.A(new_n7032), .B(new_n7004), .Y(new_n7040));
  not_8  g04692(.A(new_n7040), .Y(new_n7041));
  nor_5  g04693(.A(new_n7041), .B(new_n7039), .Y(new_n7042));
  xor_4  g04694(.A(new_n7041), .B(new_n7039), .Y(new_n7043));
  not_8  g04695(.A(new_n7043), .Y(new_n7044));
  xor_4  g04696(.A(new_n7030), .B(new_n7009), .Y(new_n7045));
  nand_5 g04697(.A(new_n7045), .B(new_n5184), .Y(new_n7046));
  xor_4  g04698(.A(new_n7045), .B(new_n5184), .Y(new_n7047));
  xnor_4 g04699(.A(new_n7026), .B(new_n7015), .Y(new_n7048));
  or_6   g04700(.A(new_n7048), .B(new_n5094), .Y(new_n7049));
  nand_5 g04701(.A(new_n7018), .B(new_n7017), .Y(new_n7050));
  xnor_4 g04702(.A(new_n7050), .B(new_n7024), .Y(new_n7051));
  or_6   g04703(.A(new_n7051), .B(new_n5095), .Y(new_n7052));
  nand_5 g04704(.A(new_n7021), .B(new_n7020), .Y(new_n7053));
  not_8  g04705(.A(pi238), .Y(new_n7054));
  nand_5 g04706(.A(pi302), .B(new_n7054), .Y(new_n7055));
  not_8  g04707(.A(new_n7055), .Y(new_n7056));
  nor_5  g04708(.A(new_n7056), .B(new_n4637), .Y(new_n7057));
  nand_5 g04709(.A(new_n3641), .B(pi238), .Y(new_n7058));
  not_8  g04710(.A(new_n7058), .Y(new_n7059));
  or_6   g04711(.A(new_n7059), .B(new_n4627), .Y(new_n7060));
  nand_5 g04712(.A(new_n7059), .B(pi682), .Y(new_n7061));
  nand_5 g04713(.A(new_n7061), .B(new_n7060), .Y(new_n7062));
  nor_5  g04714(.A(new_n7062), .B(new_n7057), .Y(new_n7063));
  xor_4  g04715(.A(new_n7063), .B(new_n5105), .Y(new_n7064));
  or_6   g04716(.A(new_n7064), .B(new_n7053), .Y(new_n7065));
  nand_5 g04717(.A(new_n7065), .B(new_n7022), .Y(new_n7066));
  nand_5 g04718(.A(new_n7064), .B(new_n7053), .Y(new_n7067));
  nand_5 g04719(.A(new_n7067), .B(pi574), .Y(new_n7068));
  nand_5 g04720(.A(new_n7068), .B(new_n7066), .Y(new_n7069));
  nand_5 g04721(.A(new_n5087), .B(new_n5105), .Y(new_n7070));
  and_6  g04722(.A(new_n7070), .B(new_n7053), .Y(new_n7071));
  xor_4  g04723(.A(pi574), .B(new_n7054), .Y(new_n7072));
  nor_5  g04724(.A(new_n7072), .B(new_n7071), .Y(new_n7073));
  nand_5 g04725(.A(new_n5098), .B(new_n5105), .Y(new_n7074));
  nand_5 g04726(.A(new_n7074), .B(new_n5089), .Y(new_n7075));
  nor_5  g04727(.A(new_n7075), .B(new_n7073), .Y(new_n7076));
  nand_5 g04728(.A(new_n7076), .B(new_n7069), .Y(new_n7077));
  nand_5 g04729(.A(new_n7051), .B(new_n5095), .Y(new_n7078));
  nand_5 g04730(.A(new_n7078), .B(new_n7077), .Y(new_n7079));
  nand_5 g04731(.A(new_n7079), .B(new_n7052), .Y(new_n7080));
  nand_5 g04732(.A(new_n7080), .B(new_n7049), .Y(new_n7081));
  nand_5 g04733(.A(new_n7048), .B(new_n5094), .Y(new_n7082));
  nand_5 g04734(.A(new_n7082), .B(new_n7081), .Y(new_n7083));
  nand_5 g04735(.A(new_n7012), .B(new_n7011), .Y(new_n7084));
  xor_4  g04736(.A(new_n7084), .B(new_n7028), .Y(new_n7085));
  or_6   g04737(.A(new_n7085), .B(new_n5124), .Y(new_n7086));
  nand_5 g04738(.A(new_n7086), .B(new_n7083), .Y(new_n7087));
  nand_5 g04739(.A(new_n7085), .B(new_n5124), .Y(new_n7088));
  nand_5 g04740(.A(new_n7088), .B(new_n7087), .Y(new_n7089));
  nand_5 g04741(.A(new_n7089), .B(new_n7047), .Y(new_n7090));
  nand_5 g04742(.A(new_n7090), .B(new_n7046), .Y(new_n7091));
  nor_5  g04743(.A(new_n7091), .B(new_n7044), .Y(new_n7092));
  or_6   g04744(.A(new_n7092), .B(new_n7042), .Y(new_n7093));
  nand_5 g04745(.A(new_n7093), .B(new_n7038), .Y(new_n7094));
  and_6  g04746(.A(new_n7094), .B(new_n7037), .Y(new_n7095));
  nand_5 g04747(.A(pi507), .B(pi423), .Y(new_n7096));
  nand_5 g04748(.A(new_n7000), .B(new_n6993), .Y(new_n7097));
  nand_5 g04749(.A(new_n7097), .B(new_n7096), .Y(new_n7098));
  nand_5 g04750(.A(pi446), .B(pi408), .Y(new_n7099));
  not_8  g04751(.A(pi408), .Y(new_n7100));
  nand_5 g04752(.A(new_n3525), .B(new_n7100), .Y(new_n7101));
  and_6  g04753(.A(new_n7101), .B(new_n7099), .Y(new_n7102));
  xor_4  g04754(.A(new_n7102), .B(new_n7098), .Y(new_n7103));
  not_8  g04755(.A(new_n7103), .Y(new_n7104));
  nand_5 g04756(.A(pi314), .B(pi180), .Y(new_n7105));
  not_8  g04757(.A(new_n7105), .Y(new_n7106));
  not_8  g04758(.A(new_n7035), .Y(new_n7107));
  nor_5  g04759(.A(new_n7107), .B(new_n7034), .Y(new_n7108));
  nor_5  g04760(.A(new_n7108), .B(new_n7106), .Y(new_n7109));
  xor_4  g04761(.A(pi029), .B(pi009), .Y(new_n7110));
  xor_4  g04762(.A(new_n7110), .B(new_n7109), .Y(new_n7111));
  xor_4  g04763(.A(new_n7111), .B(new_n7104), .Y(new_n7112));
  xor_4  g04764(.A(new_n7112), .B(new_n7095), .Y(new_n7113));
  or_6   g04765(.A(new_n7113), .B(new_n6992), .Y(new_n7114));
  xor_4  g04766(.A(new_n7113), .B(new_n6992), .Y(new_n7115));
  xor_4  g04767(.A(new_n6989), .B(new_n6956), .Y(new_n7116));
  not_8  g04768(.A(new_n7116), .Y(new_n7117));
  xor_4  g04769(.A(new_n6985), .B(new_n6962), .Y(new_n7118));
  xor_4  g04770(.A(new_n7089), .B(new_n7047), .Y(new_n7119));
  not_8  g04771(.A(new_n7119), .Y(new_n7120));
  or_6   g04772(.A(new_n7120), .B(new_n7118), .Y(new_n7121));
  xor_4  g04773(.A(new_n6983), .B(new_n6965), .Y(new_n7122));
  not_8  g04774(.A(new_n7122), .Y(new_n7123));
  nand_5 g04775(.A(new_n7088), .B(new_n7086), .Y(new_n7124));
  xnor_4 g04776(.A(new_n7124), .B(new_n7083), .Y(new_n7125));
  nand_5 g04777(.A(new_n7125), .B(new_n7123), .Y(new_n7126));
  xor_4  g04778(.A(new_n7125), .B(new_n7122), .Y(new_n7127));
  xor_4  g04779(.A(new_n6981), .B(new_n6968), .Y(new_n7128));
  xor_4  g04780(.A(new_n6979), .B(new_n6971), .Y(new_n7129));
  not_8  g04781(.A(new_n7129), .Y(new_n7130));
  not_8  g04782(.A(new_n6978), .Y(new_n7131));
  nand_5 g04783(.A(new_n7067), .B(new_n7065), .Y(new_n7132));
  nand_5 g04784(.A(new_n7058), .B(new_n7055), .Y(new_n7133));
  xor_4  g04785(.A(new_n7133), .B(new_n4637), .Y(new_n7134));
  not_8  g04786(.A(new_n7134), .Y(new_n7135));
  nand_5 g04787(.A(new_n7135), .B(new_n7132), .Y(new_n7136));
  nand_5 g04788(.A(new_n7136), .B(new_n7131), .Y(new_n7137));
  nand_5 g04789(.A(pi367), .B(new_n2419), .Y(new_n7138));
  nor_5  g04790(.A(new_n7138), .B(new_n7135), .Y(new_n7139));
  nor_5  g04791(.A(new_n7134), .B(new_n6976), .Y(new_n7140));
  or_6   g04792(.A(new_n7140), .B(new_n7139), .Y(new_n7141));
  nor_5  g04793(.A(new_n7141), .B(new_n6974), .Y(new_n7142));
  or_6   g04794(.A(new_n7142), .B(new_n7139), .Y(new_n7143));
  xnor_4 g04795(.A(new_n7141), .B(new_n6974), .Y(new_n7144));
  nand_5 g04796(.A(new_n7144), .B(new_n7132), .Y(new_n7145));
  nand_5 g04797(.A(new_n7145), .B(new_n7143), .Y(new_n7146));
  nand_5 g04798(.A(new_n7146), .B(new_n7137), .Y(new_n7147));
  nor_5  g04799(.A(new_n7147), .B(new_n7130), .Y(new_n7148));
  xor_4  g04800(.A(new_n7147), .B(new_n7129), .Y(new_n7149));
  nand_5 g04801(.A(new_n7078), .B(new_n7052), .Y(new_n7150));
  xnor_4 g04802(.A(new_n7150), .B(new_n7077), .Y(new_n7151));
  nor_5  g04803(.A(new_n7151), .B(new_n7149), .Y(new_n7152));
  or_6   g04804(.A(new_n7152), .B(new_n7148), .Y(new_n7153));
  nand_5 g04805(.A(new_n7153), .B(new_n7128), .Y(new_n7154));
  or_6   g04806(.A(new_n7153), .B(new_n7128), .Y(new_n7155));
  nand_5 g04807(.A(new_n7082), .B(new_n7049), .Y(new_n7156));
  xor_4  g04808(.A(new_n7156), .B(new_n7080), .Y(new_n7157));
  nand_5 g04809(.A(new_n7157), .B(new_n7155), .Y(new_n7158));
  nand_5 g04810(.A(new_n7158), .B(new_n7154), .Y(new_n7159));
  or_6   g04811(.A(new_n7159), .B(new_n7127), .Y(new_n7160));
  nand_5 g04812(.A(new_n7160), .B(new_n7126), .Y(new_n7161));
  xor_4  g04813(.A(new_n7120), .B(new_n7118), .Y(new_n7162));
  nand_5 g04814(.A(new_n7162), .B(new_n7161), .Y(new_n7163));
  nand_5 g04815(.A(new_n7163), .B(new_n7121), .Y(new_n7164));
  xor_4  g04816(.A(new_n7091), .B(new_n7043), .Y(new_n7165));
  nand_5 g04817(.A(new_n7165), .B(new_n7164), .Y(new_n7166));
  xor_4  g04818(.A(new_n7165), .B(new_n7164), .Y(new_n7167));
  not_8  g04819(.A(new_n7167), .Y(new_n7168));
  xor_4  g04820(.A(new_n6987), .B(new_n6959), .Y(new_n7169));
  or_6   g04821(.A(new_n7169), .B(new_n7168), .Y(new_n7170));
  nand_5 g04822(.A(new_n7170), .B(new_n7166), .Y(new_n7171));
  nor_5  g04823(.A(new_n7171), .B(new_n7117), .Y(new_n7172));
  xor_4  g04824(.A(new_n7171), .B(new_n7116), .Y(new_n7173));
  nor_5  g04825(.A(new_n7092), .B(new_n7042), .Y(new_n7174));
  xor_4  g04826(.A(new_n7174), .B(new_n7038), .Y(new_n7175));
  nor_5  g04827(.A(new_n7175), .B(new_n7173), .Y(new_n7176));
  nor_5  g04828(.A(new_n7176), .B(new_n7172), .Y(new_n7177));
  nand_5 g04829(.A(new_n7177), .B(new_n7115), .Y(new_n7178));
  nand_5 g04830(.A(new_n7178), .B(new_n7114), .Y(new_n7179));
  not_8  g04831(.A(new_n7179), .Y(new_n7180));
  not_8  g04832(.A(pi775), .Y(new_n7181));
  nand_5 g04833(.A(new_n7181), .B(pi646), .Y(new_n7182));
  nand_5 g04834(.A(new_n6991), .B(new_n6952), .Y(new_n7183));
  nand_5 g04835(.A(new_n7183), .B(new_n7182), .Y(new_n7184));
  not_8  g04836(.A(pi833), .Y(new_n7185));
  nand_5 g04837(.A(new_n7185), .B(pi072), .Y(new_n7186));
  not_8  g04838(.A(pi072), .Y(new_n7187));
  nand_5 g04839(.A(pi833), .B(new_n7187), .Y(new_n7188));
  nand_5 g04840(.A(new_n7188), .B(new_n7186), .Y(new_n7189));
  xnor_4 g04841(.A(new_n7189), .B(new_n7184), .Y(new_n7190));
  or_6   g04842(.A(new_n7190), .B(new_n7180), .Y(new_n7191));
  xor_4  g04843(.A(new_n7190), .B(new_n7180), .Y(new_n7192));
  not_8  g04844(.A(pi272), .Y(new_n7193));
  xor_4  g04845(.A(pi293), .B(new_n7193), .Y(new_n7194));
  nand_5 g04846(.A(new_n7101), .B(new_n7098), .Y(new_n7195));
  nand_5 g04847(.A(new_n7195), .B(new_n7099), .Y(new_n7196));
  xor_4  g04848(.A(new_n7196), .B(new_n7194), .Y(new_n7197));
  xor_4  g04849(.A(pi689), .B(pi678), .Y(new_n7198));
  nand_5 g04850(.A(pi029), .B(pi009), .Y(new_n7199));
  not_8  g04851(.A(new_n7199), .Y(new_n7200));
  not_8  g04852(.A(new_n7110), .Y(new_n7201));
  nor_5  g04853(.A(new_n7201), .B(new_n7109), .Y(new_n7202));
  nor_5  g04854(.A(new_n7202), .B(new_n7200), .Y(new_n7203));
  xor_4  g04855(.A(new_n7203), .B(new_n7198), .Y(new_n7204));
  not_8  g04856(.A(new_n7204), .Y(new_n7205));
  xor_4  g04857(.A(new_n7205), .B(new_n7197), .Y(new_n7206));
  nand_5 g04858(.A(new_n7111), .B(new_n7103), .Y(new_n7207));
  not_8  g04859(.A(new_n7207), .Y(new_n7208));
  nor_5  g04860(.A(new_n7112), .B(new_n7095), .Y(new_n7209));
  nor_5  g04861(.A(new_n7209), .B(new_n7208), .Y(new_n7210));
  xor_4  g04862(.A(new_n7210), .B(new_n7206), .Y(new_n7211));
  nand_5 g04863(.A(new_n7211), .B(new_n7192), .Y(new_n7212));
  nand_5 g04864(.A(new_n7212), .B(new_n7191), .Y(new_n7213));
  nand_5 g04865(.A(new_n7186), .B(new_n7184), .Y(new_n7214));
  and_6  g04866(.A(new_n7214), .B(new_n7188), .Y(new_n7215));
  nor_5  g04867(.A(new_n7215), .B(new_n7213), .Y(new_n7216));
  and_6  g04868(.A(new_n7215), .B(new_n7213), .Y(new_n7217));
  nor_5  g04869(.A(new_n7217), .B(new_n7216), .Y(new_n7218));
  nand_5 g04870(.A(new_n3697), .B(new_n7193), .Y(new_n7219));
  not_8  g04871(.A(new_n7219), .Y(new_n7220));
  nor_5  g04872(.A(new_n7196), .B(new_n7194), .Y(new_n7221));
  nor_5  g04873(.A(new_n7221), .B(new_n7220), .Y(new_n7222));
  nand_5 g04874(.A(pi689), .B(pi678), .Y(new_n7223));
  not_8  g04875(.A(new_n7223), .Y(new_n7224));
  not_8  g04876(.A(new_n7198), .Y(new_n7225));
  nor_5  g04877(.A(new_n7203), .B(new_n7225), .Y(new_n7226));
  nor_5  g04878(.A(new_n7226), .B(new_n7224), .Y(new_n7227));
  nand_5 g04879(.A(new_n7227), .B(new_n7222), .Y(new_n7228));
  not_8  g04880(.A(new_n7228), .Y(new_n7229));
  nor_5  g04881(.A(new_n7205), .B(new_n7197), .Y(new_n7230));
  not_8  g04882(.A(new_n7206), .Y(new_n7231));
  nor_5  g04883(.A(new_n7210), .B(new_n7231), .Y(new_n7232));
  nor_5  g04884(.A(new_n7232), .B(new_n7230), .Y(new_n7233));
  not_8  g04885(.A(new_n7233), .Y(new_n7234));
  nand_5 g04886(.A(new_n7234), .B(new_n7229), .Y(new_n7235));
  nand_5 g04887(.A(new_n7233), .B(new_n7228), .Y(new_n7236));
  nor_5  g04888(.A(new_n7227), .B(new_n7222), .Y(new_n7237));
  not_8  g04889(.A(new_n7237), .Y(new_n7238));
  nand_5 g04890(.A(new_n7238), .B(new_n7236), .Y(new_n7239));
  nand_5 g04891(.A(new_n7237), .B(new_n7233), .Y(new_n7240));
  nand_5 g04892(.A(new_n7240), .B(new_n7239), .Y(new_n7241));
  nand_5 g04893(.A(new_n7241), .B(new_n7235), .Y(new_n7242));
  xor_4  g04894(.A(new_n7242), .B(new_n7218), .Y(po0032));
  not_8  g04895(.A(pi448), .Y(new_n7244));
  not_8  g04896(.A(pi642), .Y(new_n7245));
  nand_5 g04897(.A(new_n7245), .B(new_n7244), .Y(new_n7246));
  nand_5 g04898(.A(pi642), .B(pi448), .Y(new_n7247));
  and_6  g04899(.A(new_n7247), .B(new_n7246), .Y(new_n7248));
  not_8  g04900(.A(pi806), .Y(new_n7249));
  xor_4  g04901(.A(pi580), .B(new_n6766), .Y(new_n7250));
  xor_4  g04902(.A(new_n7250), .B(pi445), .Y(new_n7251));
  xor_4  g04903(.A(new_n7251), .B(new_n7249), .Y(new_n7252));
  xor_4  g04904(.A(new_n7252), .B(new_n7248), .Y(po0033));
  xor_4  g04905(.A(pi534), .B(new_n6091), .Y(new_n7254));
  not_8  g04906(.A(pi092), .Y(new_n7255));
  nand_5 g04907(.A(new_n7255), .B(pi028), .Y(new_n7256));
  not_8  g04908(.A(pi028), .Y(new_n7257));
  xor_4  g04909(.A(pi092), .B(new_n7257), .Y(new_n7258));
  nand_5 g04910(.A(pi772), .B(new_n6077), .Y(new_n7259));
  xor_4  g04911(.A(pi772), .B(new_n6077), .Y(new_n7260));
  nand_5 g04912(.A(pi332), .B(new_n5940), .Y(new_n7261));
  xor_4  g04913(.A(pi332), .B(new_n5940), .Y(new_n7262));
  not_8  g04914(.A(pi120), .Y(new_n7263));
  nand_5 g04915(.A(pi265), .B(new_n7263), .Y(new_n7264));
  xor_4  g04916(.A(pi265), .B(new_n7263), .Y(new_n7265));
  not_8  g04917(.A(pi432), .Y(new_n7266));
  nand_5 g04918(.A(pi635), .B(new_n7266), .Y(new_n7267));
  xor_4  g04919(.A(pi635), .B(new_n7266), .Y(new_n7268));
  nand_5 g04920(.A(new_n5977), .B(pi545), .Y(new_n7269));
  not_8  g04921(.A(pi545), .Y(new_n7270));
  xor_4  g04922(.A(pi645), .B(new_n7270), .Y(new_n7271));
  nand_5 g04923(.A(new_n4149), .B(pi388), .Y(new_n7272));
  xor_4  g04924(.A(pi825), .B(new_n6575), .Y(new_n7273));
  nand_5 g04925(.A(new_n4152), .B(pi161), .Y(new_n7274));
  nand_5 g04926(.A(new_n4184), .B(pi281), .Y(new_n7275));
  xor_4  g04927(.A(pi329), .B(pi161), .Y(new_n7276));
  or_6   g04928(.A(new_n7276), .B(new_n7275), .Y(new_n7277));
  nand_5 g04929(.A(new_n7277), .B(new_n7274), .Y(new_n7278));
  nand_5 g04930(.A(new_n7278), .B(new_n7273), .Y(new_n7279));
  nand_5 g04931(.A(new_n7279), .B(new_n7272), .Y(new_n7280));
  nand_5 g04932(.A(new_n7280), .B(new_n7271), .Y(new_n7281));
  nand_5 g04933(.A(new_n7281), .B(new_n7269), .Y(new_n7282));
  nand_5 g04934(.A(new_n7282), .B(new_n7268), .Y(new_n7283));
  nand_5 g04935(.A(new_n7283), .B(new_n7267), .Y(new_n7284));
  nand_5 g04936(.A(new_n7284), .B(new_n7265), .Y(new_n7285));
  nand_5 g04937(.A(new_n7285), .B(new_n7264), .Y(new_n7286));
  nand_5 g04938(.A(new_n7286), .B(new_n7262), .Y(new_n7287));
  nand_5 g04939(.A(new_n7287), .B(new_n7261), .Y(new_n7288));
  nand_5 g04940(.A(new_n7288), .B(new_n7260), .Y(new_n7289));
  nand_5 g04941(.A(new_n7289), .B(new_n7259), .Y(new_n7290));
  nand_5 g04942(.A(new_n7290), .B(new_n7258), .Y(new_n7291));
  nand_5 g04943(.A(new_n7291), .B(new_n7256), .Y(new_n7292));
  xor_4  g04944(.A(new_n7292), .B(new_n7254), .Y(new_n7293));
  nand_5 g04945(.A(new_n7185), .B(pi582), .Y(new_n7294));
  not_8  g04946(.A(pi582), .Y(new_n7295));
  nand_5 g04947(.A(pi833), .B(new_n7295), .Y(new_n7296));
  nand_5 g04948(.A(new_n7296), .B(new_n7294), .Y(new_n7297));
  nand_5 g04949(.A(new_n6951), .B(pi404), .Y(new_n7298));
  xor_4  g04950(.A(pi646), .B(new_n2978), .Y(new_n7299));
  nand_5 g04951(.A(pi527), .B(new_n6955), .Y(new_n7300));
  xor_4  g04952(.A(pi527), .B(new_n6955), .Y(new_n7301));
  nand_5 g04953(.A(new_n3801), .B(new_n3798), .Y(new_n7302));
  nand_5 g04954(.A(new_n7302), .B(new_n3800), .Y(new_n7303));
  nand_5 g04955(.A(new_n7303), .B(new_n7301), .Y(new_n7304));
  nand_5 g04956(.A(new_n7304), .B(new_n7300), .Y(new_n7305));
  nand_5 g04957(.A(new_n7305), .B(new_n7299), .Y(new_n7306));
  nand_5 g04958(.A(new_n7306), .B(new_n7298), .Y(new_n7307));
  not_8  g04959(.A(new_n7307), .Y(new_n7308));
  xor_4  g04960(.A(new_n7308), .B(new_n7297), .Y(new_n7309));
  or_6   g04961(.A(new_n7309), .B(new_n7293), .Y(new_n7310));
  xor_4  g04962(.A(new_n7309), .B(new_n7293), .Y(new_n7311));
  xor_4  g04963(.A(new_n7290), .B(new_n7258), .Y(new_n7312));
  not_8  g04964(.A(new_n7312), .Y(new_n7313));
  xnor_4 g04965(.A(new_n7305), .B(new_n7299), .Y(new_n7314));
  nor_5  g04966(.A(new_n7314), .B(new_n7313), .Y(new_n7315));
  xor_4  g04967(.A(new_n7314), .B(new_n7313), .Y(new_n7316));
  not_8  g04968(.A(new_n7316), .Y(new_n7317));
  xor_4  g04969(.A(new_n7288), .B(new_n7260), .Y(new_n7318));
  not_8  g04970(.A(new_n7318), .Y(new_n7319));
  xor_4  g04971(.A(new_n7303), .B(new_n7301), .Y(new_n7320));
  not_8  g04972(.A(new_n7320), .Y(new_n7321));
  nand_5 g04973(.A(new_n7321), .B(new_n7319), .Y(new_n7322));
  xor_4  g04974(.A(new_n7320), .B(new_n7318), .Y(new_n7323));
  xor_4  g04975(.A(new_n7286), .B(new_n7262), .Y(new_n7324));
  not_8  g04976(.A(new_n7324), .Y(new_n7325));
  nand_5 g04977(.A(new_n7325), .B(new_n3804), .Y(new_n7326));
  xor_4  g04978(.A(new_n7324), .B(new_n3803), .Y(new_n7327));
  xor_4  g04979(.A(new_n7284), .B(new_n7265), .Y(new_n7328));
  not_8  g04980(.A(new_n7328), .Y(new_n7329));
  nand_5 g04981(.A(new_n7329), .B(new_n3806), .Y(new_n7330));
  xor_4  g04982(.A(new_n7329), .B(new_n3806), .Y(new_n7331));
  xor_4  g04983(.A(new_n7282), .B(new_n7268), .Y(new_n7332));
  not_8  g04984(.A(new_n7332), .Y(new_n7333));
  nor_5  g04985(.A(new_n7333), .B(new_n3810), .Y(new_n7334));
  xor_4  g04986(.A(new_n7333), .B(new_n3810), .Y(new_n7335));
  not_8  g04987(.A(new_n7335), .Y(new_n7336));
  xor_4  g04988(.A(new_n7280), .B(new_n7271), .Y(new_n7337));
  not_8  g04989(.A(new_n7337), .Y(new_n7338));
  nand_5 g04990(.A(new_n7338), .B(new_n3813), .Y(new_n7339));
  xor_4  g04991(.A(new_n7337), .B(new_n3812), .Y(new_n7340));
  xor_4  g04992(.A(new_n7278), .B(new_n7273), .Y(new_n7341));
  or_6   g04993(.A(new_n7341), .B(new_n3827), .Y(new_n7342));
  not_8  g04994(.A(pi281), .Y(new_n7343));
  xor_4  g04995(.A(pi295), .B(new_n7343), .Y(new_n7344));
  not_8  g04996(.A(new_n7344), .Y(new_n7345));
  nor_5  g04997(.A(new_n7345), .B(new_n7276), .Y(new_n7346));
  nor_5  g04998(.A(new_n7346), .B(new_n3789), .Y(new_n7347));
  xor_4  g04999(.A(new_n7276), .B(new_n7275), .Y(new_n7348));
  not_8  g05000(.A(new_n7348), .Y(new_n7349));
  xor_4  g05001(.A(new_n7349), .B(new_n3786), .Y(new_n7350));
  nor_5  g05002(.A(new_n7344), .B(new_n3816), .Y(new_n7351));
  nor_5  g05003(.A(new_n7351), .B(new_n7350), .Y(new_n7352));
  nand_5 g05004(.A(new_n7348), .B(new_n3786), .Y(new_n7353));
  nand_5 g05005(.A(new_n7344), .B(new_n3788), .Y(new_n7354));
  nand_5 g05006(.A(new_n7354), .B(new_n7353), .Y(new_n7355));
  nor_5  g05007(.A(new_n7355), .B(new_n7352), .Y(new_n7356));
  or_6   g05008(.A(new_n7356), .B(new_n7347), .Y(new_n7357));
  xor_4  g05009(.A(new_n7341), .B(new_n3827), .Y(new_n7358));
  nand_5 g05010(.A(new_n7358), .B(new_n7357), .Y(new_n7359));
  nand_5 g05011(.A(new_n7359), .B(new_n7342), .Y(new_n7360));
  nand_5 g05012(.A(new_n7360), .B(new_n7340), .Y(new_n7361));
  nand_5 g05013(.A(new_n7361), .B(new_n7339), .Y(new_n7362));
  nor_5  g05014(.A(new_n7362), .B(new_n7336), .Y(new_n7363));
  nor_5  g05015(.A(new_n7363), .B(new_n7334), .Y(new_n7364));
  nand_5 g05016(.A(new_n7364), .B(new_n7331), .Y(new_n7365));
  nand_5 g05017(.A(new_n7365), .B(new_n7330), .Y(new_n7366));
  nand_5 g05018(.A(new_n7366), .B(new_n7327), .Y(new_n7367));
  nand_5 g05019(.A(new_n7367), .B(new_n7326), .Y(new_n7368));
  nand_5 g05020(.A(new_n7368), .B(new_n7323), .Y(new_n7369));
  nand_5 g05021(.A(new_n7369), .B(new_n7322), .Y(new_n7370));
  nor_5  g05022(.A(new_n7370), .B(new_n7317), .Y(new_n7371));
  nor_5  g05023(.A(new_n7371), .B(new_n7315), .Y(new_n7372));
  nand_5 g05024(.A(new_n7372), .B(new_n7311), .Y(new_n7373));
  nand_5 g05025(.A(new_n7373), .B(new_n7310), .Y(new_n7374));
  nand_5 g05026(.A(pi534), .B(new_n6091), .Y(new_n7375));
  nand_5 g05027(.A(new_n7292), .B(new_n7254), .Y(new_n7376));
  nand_5 g05028(.A(new_n7376), .B(new_n7375), .Y(new_n7377));
  not_8  g05029(.A(new_n7377), .Y(new_n7378));
  nand_5 g05030(.A(new_n7307), .B(new_n7296), .Y(new_n7379));
  nand_5 g05031(.A(new_n7379), .B(new_n7294), .Y(new_n7380));
  not_8  g05032(.A(new_n7380), .Y(new_n7381));
  nand_5 g05033(.A(new_n7381), .B(new_n7378), .Y(new_n7382));
  not_8  g05034(.A(new_n7382), .Y(new_n7383));
  nand_5 g05035(.A(new_n7383), .B(new_n7374), .Y(new_n7384));
  nand_5 g05036(.A(new_n7380), .B(new_n7377), .Y(new_n7385));
  not_8  g05037(.A(new_n7385), .Y(new_n7386));
  nor_5  g05038(.A(new_n7383), .B(new_n7374), .Y(new_n7387));
  nor_5  g05039(.A(new_n7387), .B(new_n7386), .Y(new_n7388));
  not_8  g05040(.A(new_n7388), .Y(new_n7389));
  nor_5  g05041(.A(new_n7385), .B(new_n7374), .Y(new_n7390));
  not_8  g05042(.A(new_n7390), .Y(new_n7391));
  nand_5 g05043(.A(new_n7391), .B(new_n7389), .Y(new_n7392));
  nand_5 g05044(.A(new_n7392), .B(new_n7384), .Y(new_n7393));
  xor_4  g05045(.A(new_n7372), .B(new_n7311), .Y(new_n7394));
  xor_4  g05046(.A(new_n7368), .B(new_n7323), .Y(new_n7395));
  xor_4  g05047(.A(new_n7366), .B(new_n7327), .Y(new_n7396));
  not_8  g05048(.A(new_n7396), .Y(new_n7397));
  xor_4  g05049(.A(pi641), .B(new_n4756), .Y(new_n7398));
  nand_5 g05050(.A(new_n3763), .B(pi201), .Y(new_n7399));
  xor_4  g05051(.A(pi298), .B(new_n3718), .Y(new_n7400));
  nand_5 g05052(.A(pi795), .B(new_n3758), .Y(new_n7401));
  nor_5  g05053(.A(new_n3723), .B(pi241), .Y(new_n7402));
  xor_4  g05054(.A(pi495), .B(new_n3746), .Y(new_n7403));
  not_8  g05055(.A(new_n7403), .Y(new_n7404));
  nand_5 g05056(.A(pi488), .B(new_n3726), .Y(new_n7405));
  nand_5 g05057(.A(new_n6018), .B(pi422), .Y(new_n7406));
  nand_5 g05058(.A(pi781), .B(new_n3860), .Y(new_n7407));
  nand_5 g05059(.A(new_n7407), .B(new_n7406), .Y(new_n7408));
  nand_5 g05060(.A(new_n7408), .B(new_n7405), .Y(new_n7409));
  nor_5  g05061(.A(new_n7409), .B(new_n7404), .Y(new_n7410));
  nor_5  g05062(.A(new_n7410), .B(new_n7402), .Y(new_n7411));
  xor_4  g05063(.A(pi795), .B(pi157), .Y(new_n7412));
  or_6   g05064(.A(new_n7412), .B(new_n7411), .Y(new_n7413));
  nand_5 g05065(.A(new_n7413), .B(new_n7401), .Y(new_n7414));
  nand_5 g05066(.A(new_n7414), .B(new_n7400), .Y(new_n7415));
  nand_5 g05067(.A(new_n7415), .B(new_n7399), .Y(new_n7416));
  xor_4  g05068(.A(new_n7416), .B(new_n7398), .Y(new_n7417));
  not_8  g05069(.A(new_n7417), .Y(new_n7418));
  xnor_4 g05070(.A(new_n7360), .B(new_n7340), .Y(new_n7419));
  xor_4  g05071(.A(new_n7412), .B(new_n7411), .Y(new_n7420));
  or_6   g05072(.A(new_n7420), .B(new_n7419), .Y(new_n7421));
  xor_4  g05073(.A(new_n7420), .B(new_n7419), .Y(new_n7422));
  not_8  g05074(.A(new_n7354), .Y(new_n7423));
  nor_5  g05075(.A(new_n7423), .B(new_n7351), .Y(new_n7424));
  xor_4  g05076(.A(new_n7424), .B(new_n7350), .Y(new_n7425));
  nand_5 g05077(.A(new_n7406), .B(new_n7405), .Y(new_n7426));
  xor_4  g05078(.A(new_n7344), .B(new_n3818), .Y(new_n7427));
  not_8  g05079(.A(new_n7427), .Y(new_n7428));
  nand_5 g05080(.A(new_n7428), .B(new_n7407), .Y(new_n7429));
  nand_5 g05081(.A(new_n4136), .B(pi631), .Y(new_n7430));
  nand_5 g05082(.A(new_n7430), .B(new_n7427), .Y(new_n7431));
  nand_5 g05083(.A(new_n7431), .B(new_n7429), .Y(new_n7432));
  xor_4  g05084(.A(new_n7432), .B(new_n7426), .Y(new_n7433));
  or_6   g05085(.A(new_n7433), .B(new_n7425), .Y(new_n7434));
  nand_5 g05086(.A(new_n7430), .B(new_n7407), .Y(new_n7435));
  nand_5 g05087(.A(new_n7435), .B(new_n7427), .Y(new_n7436));
  nand_5 g05088(.A(new_n7436), .B(new_n7433), .Y(new_n7437));
  nand_5 g05089(.A(new_n7437), .B(new_n7434), .Y(new_n7438));
  xor_4  g05090(.A(new_n7409), .B(new_n7403), .Y(new_n7439));
  not_8  g05091(.A(new_n7439), .Y(new_n7440));
  and_6  g05092(.A(new_n7440), .B(new_n7438), .Y(new_n7441));
  xor_4  g05093(.A(new_n7358), .B(new_n7357), .Y(new_n7442));
  xor_4  g05094(.A(new_n7439), .B(new_n7438), .Y(new_n7443));
  nor_5  g05095(.A(new_n7443), .B(new_n7442), .Y(new_n7444));
  nor_5  g05096(.A(new_n7444), .B(new_n7441), .Y(new_n7445));
  nand_5 g05097(.A(new_n7445), .B(new_n7422), .Y(new_n7446));
  nand_5 g05098(.A(new_n7446), .B(new_n7421), .Y(new_n7447));
  xor_4  g05099(.A(new_n7414), .B(new_n7400), .Y(new_n7448));
  not_8  g05100(.A(new_n7448), .Y(new_n7449));
  nand_5 g05101(.A(new_n7449), .B(new_n7447), .Y(new_n7450));
  xor_4  g05102(.A(new_n7362), .B(new_n7335), .Y(new_n7451));
  xor_4  g05103(.A(new_n7449), .B(new_n7447), .Y(new_n7452));
  nand_5 g05104(.A(new_n7452), .B(new_n7451), .Y(new_n7453));
  nand_5 g05105(.A(new_n7453), .B(new_n7450), .Y(new_n7454));
  nor_5  g05106(.A(new_n7454), .B(new_n7418), .Y(new_n7455));
  xor_4  g05107(.A(new_n7364), .B(new_n7331), .Y(new_n7456));
  xor_4  g05108(.A(new_n7454), .B(new_n7417), .Y(new_n7457));
  nor_5  g05109(.A(new_n7457), .B(new_n7456), .Y(new_n7458));
  or_6   g05110(.A(new_n7458), .B(new_n7455), .Y(new_n7459));
  or_6   g05111(.A(new_n7459), .B(new_n7397), .Y(new_n7460));
  xor_4  g05112(.A(pi793), .B(new_n3710), .Y(new_n7461));
  nand_5 g05113(.A(pi641), .B(new_n4756), .Y(new_n7462));
  nand_5 g05114(.A(new_n7416), .B(new_n7398), .Y(new_n7463));
  nand_5 g05115(.A(new_n7463), .B(new_n7462), .Y(new_n7464));
  xnor_4 g05116(.A(new_n7464), .B(new_n7461), .Y(new_n7465));
  xor_4  g05117(.A(new_n7459), .B(new_n7396), .Y(new_n7466));
  not_8  g05118(.A(new_n7466), .Y(new_n7467));
  nand_5 g05119(.A(new_n7467), .B(new_n7465), .Y(new_n7468));
  nand_5 g05120(.A(new_n7468), .B(new_n7460), .Y(new_n7469));
  nor_5  g05121(.A(new_n7469), .B(new_n7395), .Y(new_n7470));
  not_8  g05122(.A(pi021), .Y(new_n7471));
  xor_4  g05123(.A(pi623), .B(new_n7471), .Y(new_n7472));
  nand_5 g05124(.A(new_n3709), .B(pi064), .Y(new_n7473));
  nand_5 g05125(.A(new_n7464), .B(new_n7461), .Y(new_n7474));
  nand_5 g05126(.A(new_n7474), .B(new_n7473), .Y(new_n7475));
  xnor_4 g05127(.A(new_n7475), .B(new_n7472), .Y(new_n7476));
  xnor_4 g05128(.A(new_n7469), .B(new_n7395), .Y(new_n7477));
  nor_5  g05129(.A(new_n7477), .B(new_n7476), .Y(new_n7478));
  nor_5  g05130(.A(new_n7478), .B(new_n7470), .Y(new_n7479));
  nand_5 g05131(.A(new_n4843), .B(pi021), .Y(new_n7480));
  nand_5 g05132(.A(new_n7475), .B(new_n7472), .Y(new_n7481));
  nand_5 g05133(.A(new_n7481), .B(new_n7480), .Y(new_n7482));
  not_8  g05134(.A(pi607), .Y(new_n7483));
  nand_5 g05135(.A(new_n7483), .B(pi013), .Y(new_n7484));
  nand_5 g05136(.A(pi607), .B(new_n4838), .Y(new_n7485));
  nand_5 g05137(.A(new_n7485), .B(new_n7484), .Y(new_n7486));
  xor_4  g05138(.A(new_n7486), .B(new_n7482), .Y(new_n7487));
  nand_5 g05139(.A(new_n7487), .B(new_n7479), .Y(new_n7488));
  xor_4  g05140(.A(new_n7370), .B(new_n7316), .Y(new_n7489));
  xor_4  g05141(.A(new_n7487), .B(new_n7479), .Y(new_n7490));
  nand_5 g05142(.A(new_n7490), .B(new_n7489), .Y(new_n7491));
  nand_5 g05143(.A(new_n7491), .B(new_n7488), .Y(new_n7492));
  nand_5 g05144(.A(new_n7492), .B(new_n7394), .Y(new_n7493));
  not_8  g05145(.A(pi381), .Y(new_n7494));
  nand_5 g05146(.A(new_n7494), .B(pi097), .Y(new_n7495));
  nand_5 g05147(.A(new_n7484), .B(new_n7482), .Y(new_n7496));
  nand_5 g05148(.A(new_n7496), .B(new_n7485), .Y(new_n7497));
  nand_5 g05149(.A(new_n7497), .B(new_n7495), .Y(new_n7498));
  nand_5 g05150(.A(pi381), .B(new_n4857), .Y(new_n7499));
  nand_5 g05151(.A(new_n7499), .B(new_n7498), .Y(new_n7500));
  nor_5  g05152(.A(new_n7500), .B(new_n7493), .Y(new_n7501));
  nor_5  g05153(.A(new_n7492), .B(new_n7394), .Y(new_n7502));
  or_6   g05154(.A(new_n7497), .B(new_n7495), .Y(new_n7503));
  nor_5  g05155(.A(new_n7503), .B(new_n7502), .Y(new_n7504));
  nor_5  g05156(.A(new_n7504), .B(new_n7501), .Y(new_n7505));
  not_8  g05157(.A(new_n7505), .Y(new_n7506));
  nand_5 g05158(.A(new_n7502), .B(new_n7500), .Y(new_n7507));
  not_8  g05159(.A(new_n7497), .Y(new_n7508));
  nor_5  g05160(.A(new_n7499), .B(new_n7508), .Y(new_n7509));
  nand_5 g05161(.A(new_n7509), .B(new_n7493), .Y(new_n7510));
  nand_5 g05162(.A(new_n7510), .B(new_n7507), .Y(new_n7511));
  or_6   g05163(.A(new_n7511), .B(new_n7506), .Y(new_n7512));
  xor_4  g05164(.A(new_n7512), .B(new_n7393), .Y(po0034));
  nand_5 g05165(.A(pi430), .B(pi114), .Y(new_n7514));
  nand_5 g05166(.A(new_n5451), .B(new_n3327), .Y(new_n7515));
  nand_5 g05167(.A(pi777), .B(pi325), .Y(new_n7516));
  nand_5 g05168(.A(new_n5454), .B(new_n3262), .Y(new_n7517));
  nand_5 g05169(.A(pi637), .B(pi319), .Y(new_n7518));
  xor_4  g05170(.A(pi637), .B(pi319), .Y(new_n7519));
  nand_5 g05171(.A(pi429), .B(pi253), .Y(new_n7520));
  nand_5 g05172(.A(new_n2410), .B(new_n2381), .Y(new_n7521));
  nand_5 g05173(.A(new_n7521), .B(new_n7520), .Y(new_n7522));
  nand_5 g05174(.A(new_n7522), .B(new_n7519), .Y(new_n7523));
  nand_5 g05175(.A(new_n7523), .B(new_n7518), .Y(new_n7524));
  nand_5 g05176(.A(new_n7524), .B(new_n7517), .Y(new_n7525));
  nand_5 g05177(.A(new_n7525), .B(new_n7516), .Y(new_n7526));
  nand_5 g05178(.A(new_n7526), .B(new_n7515), .Y(new_n7527));
  nand_5 g05179(.A(new_n7527), .B(new_n7514), .Y(new_n7528));
  nand_5 g05180(.A(pi833), .B(pi697), .Y(new_n7529));
  not_8  g05181(.A(pi697), .Y(new_n7530));
  nand_5 g05182(.A(new_n7185), .B(new_n7530), .Y(new_n7531));
  nand_5 g05183(.A(pi646), .B(pi452), .Y(new_n7532));
  not_8  g05184(.A(pi452), .Y(new_n7533));
  nand_5 g05185(.A(new_n6951), .B(new_n7533), .Y(new_n7534));
  nand_5 g05186(.A(pi139), .B(pi046), .Y(new_n7535));
  xor_4  g05187(.A(pi139), .B(pi046), .Y(new_n7536));
  nand_5 g05188(.A(pi683), .B(pi439), .Y(new_n7537));
  nand_5 g05189(.A(new_n2378), .B(new_n2349), .Y(new_n7538));
  nand_5 g05190(.A(new_n7538), .B(new_n7537), .Y(new_n7539));
  nand_5 g05191(.A(new_n7539), .B(new_n7536), .Y(new_n7540));
  nand_5 g05192(.A(new_n7540), .B(new_n7535), .Y(new_n7541));
  nand_5 g05193(.A(new_n7541), .B(new_n7534), .Y(new_n7542));
  nand_5 g05194(.A(new_n7542), .B(new_n7532), .Y(new_n7543));
  nand_5 g05195(.A(new_n7543), .B(new_n7531), .Y(new_n7544));
  nand_5 g05196(.A(new_n7544), .B(new_n7529), .Y(new_n7545));
  not_8  g05197(.A(new_n7545), .Y(new_n7546));
  or_6   g05198(.A(new_n7546), .B(new_n7528), .Y(new_n7547));
  nand_5 g05199(.A(new_n7546), .B(new_n7528), .Y(new_n7548));
  nand_5 g05200(.A(new_n7531), .B(new_n7529), .Y(new_n7549));
  xor_4  g05201(.A(new_n7549), .B(new_n7543), .Y(new_n7550));
  not_8  g05202(.A(new_n7550), .Y(new_n7551));
  nand_5 g05203(.A(new_n7515), .B(new_n7514), .Y(new_n7552));
  xor_4  g05204(.A(new_n7552), .B(new_n7526), .Y(new_n7553));
  nand_5 g05205(.A(new_n7553), .B(new_n7551), .Y(new_n7554));
  xor_4  g05206(.A(new_n7553), .B(new_n7551), .Y(new_n7555));
  nand_5 g05207(.A(new_n7517), .B(new_n7516), .Y(new_n7556));
  xor_4  g05208(.A(new_n7556), .B(new_n7524), .Y(new_n7557));
  not_8  g05209(.A(new_n7557), .Y(new_n7558));
  nand_5 g05210(.A(new_n7534), .B(new_n7532), .Y(new_n7559));
  xor_4  g05211(.A(new_n7559), .B(new_n7541), .Y(new_n7560));
  or_6   g05212(.A(new_n7560), .B(new_n7558), .Y(new_n7561));
  xor_4  g05213(.A(new_n7560), .B(new_n7558), .Y(new_n7562));
  xor_4  g05214(.A(new_n7522), .B(new_n7519), .Y(new_n7563));
  xnor_4 g05215(.A(new_n7539), .B(new_n7536), .Y(new_n7564));
  nor_5  g05216(.A(new_n7564), .B(new_n7563), .Y(new_n7565));
  xor_4  g05217(.A(new_n7564), .B(new_n7563), .Y(new_n7566));
  nand_5 g05218(.A(new_n2465), .B(new_n2411), .Y(new_n7567));
  not_8  g05219(.A(new_n7567), .Y(new_n7568));
  nor_5  g05220(.A(new_n2466), .B(new_n2379), .Y(new_n7569));
  nor_5  g05221(.A(new_n7569), .B(new_n7568), .Y(new_n7570));
  nand_5 g05222(.A(new_n7570), .B(new_n7566), .Y(new_n7571));
  not_8  g05223(.A(new_n7571), .Y(new_n7572));
  nor_5  g05224(.A(new_n7572), .B(new_n7565), .Y(new_n7573));
  not_8  g05225(.A(new_n7573), .Y(new_n7574));
  nand_5 g05226(.A(new_n7574), .B(new_n7562), .Y(new_n7575));
  nand_5 g05227(.A(new_n7575), .B(new_n7561), .Y(new_n7576));
  nand_5 g05228(.A(new_n7576), .B(new_n7555), .Y(new_n7577));
  nand_5 g05229(.A(new_n7577), .B(new_n7554), .Y(new_n7578));
  nand_5 g05230(.A(new_n7578), .B(new_n7548), .Y(new_n7579));
  nand_5 g05231(.A(new_n7579), .B(new_n7547), .Y(new_n7580));
  not_8  g05232(.A(new_n7580), .Y(new_n7581));
  or_6   g05233(.A(new_n7578), .B(new_n7548), .Y(new_n7582));
  not_8  g05234(.A(new_n7578), .Y(new_n7583));
  nor_5  g05235(.A(new_n7583), .B(new_n7547), .Y(new_n7584));
  nor_5  g05236(.A(new_n7584), .B(new_n7581), .Y(new_n7585));
  not_8  g05237(.A(new_n7585), .Y(new_n7586));
  nand_5 g05238(.A(new_n7586), .B(new_n7582), .Y(new_n7587));
  xor_4  g05239(.A(new_n7576), .B(new_n7555), .Y(new_n7588));
  not_8  g05240(.A(new_n7588), .Y(new_n7589));
  not_8  g05241(.A(pi096), .Y(new_n7590));
  xor_4  g05242(.A(pi582), .B(new_n7590), .Y(new_n7591));
  not_8  g05243(.A(pi728), .Y(new_n7592));
  nand_5 g05244(.A(new_n7592), .B(pi404), .Y(new_n7593));
  xor_4  g05245(.A(pi728), .B(new_n2978), .Y(new_n7594));
  nand_5 g05246(.A(pi527), .B(new_n6787), .Y(new_n7595));
  xor_4  g05247(.A(pi527), .B(new_n6787), .Y(new_n7596));
  nand_5 g05248(.A(pi816), .B(new_n6714), .Y(new_n7597));
  nand_5 g05249(.A(pi709), .B(new_n6716), .Y(new_n7598));
  nand_5 g05250(.A(pi590), .B(new_n6719), .Y(new_n7599));
  xor_4  g05251(.A(pi590), .B(new_n6719), .Y(new_n7600));
  nand_5 g05252(.A(new_n6723), .B(pi328), .Y(new_n7601));
  xor_4  g05253(.A(pi483), .B(new_n2948), .Y(new_n7602));
  nand_5 g05254(.A(pi277), .B(new_n6726), .Y(new_n7603));
  xor_4  g05255(.A(pi277), .B(new_n6726), .Y(new_n7604));
  nand_5 g05256(.A(new_n6732), .B(pi313), .Y(new_n7605));
  xor_4  g05257(.A(pi333), .B(new_n3785), .Y(new_n7606));
  nor_5  g05258(.A(new_n3815), .B(pi569), .Y(new_n7607));
  nand_5 g05259(.A(new_n7607), .B(new_n7606), .Y(new_n7608));
  nand_5 g05260(.A(new_n7608), .B(new_n7605), .Y(new_n7609));
  nand_5 g05261(.A(new_n7609), .B(new_n7604), .Y(new_n7610));
  nand_5 g05262(.A(new_n7610), .B(new_n7603), .Y(new_n7611));
  nand_5 g05263(.A(new_n7611), .B(new_n7602), .Y(new_n7612));
  nand_5 g05264(.A(new_n7612), .B(new_n7601), .Y(new_n7613));
  nand_5 g05265(.A(new_n7613), .B(new_n7600), .Y(new_n7614));
  nand_5 g05266(.A(new_n7614), .B(new_n7599), .Y(new_n7615));
  xor_4  g05267(.A(pi709), .B(new_n6716), .Y(new_n7616));
  nand_5 g05268(.A(new_n7616), .B(new_n7615), .Y(new_n7617));
  nand_5 g05269(.A(new_n7617), .B(new_n7598), .Y(new_n7618));
  xor_4  g05270(.A(pi816), .B(new_n6714), .Y(new_n7619));
  nand_5 g05271(.A(new_n7619), .B(new_n7618), .Y(new_n7620));
  nand_5 g05272(.A(new_n7620), .B(new_n7597), .Y(new_n7621));
  nand_5 g05273(.A(new_n7621), .B(new_n7596), .Y(new_n7622));
  nand_5 g05274(.A(new_n7622), .B(new_n7595), .Y(new_n7623));
  nand_5 g05275(.A(new_n7623), .B(new_n7594), .Y(new_n7624));
  nand_5 g05276(.A(new_n7624), .B(new_n7593), .Y(new_n7625));
  xnor_4 g05277(.A(new_n7625), .B(new_n7591), .Y(new_n7626));
  nor_5  g05278(.A(new_n7626), .B(new_n7589), .Y(new_n7627));
  xor_4  g05279(.A(new_n7623), .B(new_n7594), .Y(new_n7628));
  xor_4  g05280(.A(new_n7573), .B(new_n7562), .Y(new_n7629));
  not_8  g05281(.A(new_n7629), .Y(new_n7630));
  nand_5 g05282(.A(new_n7630), .B(new_n7628), .Y(new_n7631));
  xnor_4 g05283(.A(new_n7621), .B(new_n7596), .Y(new_n7632));
  xor_4  g05284(.A(new_n7570), .B(new_n7566), .Y(new_n7633));
  not_8  g05285(.A(new_n7633), .Y(new_n7634));
  or_6   g05286(.A(new_n7634), .B(new_n7632), .Y(new_n7635));
  not_8  g05287(.A(new_n2467), .Y(new_n7636));
  xnor_4 g05288(.A(new_n7619), .B(new_n7618), .Y(new_n7637));
  nor_5  g05289(.A(new_n7637), .B(new_n7636), .Y(new_n7638));
  xor_4  g05290(.A(new_n7637), .B(new_n2467), .Y(new_n7639));
  xor_4  g05291(.A(new_n7616), .B(new_n7615), .Y(new_n7640));
  or_6   g05292(.A(new_n7640), .B(new_n2503), .Y(new_n7641));
  xor_4  g05293(.A(new_n7640), .B(new_n2503), .Y(new_n7642));
  xnor_4 g05294(.A(new_n7613), .B(new_n7600), .Y(new_n7643));
  nor_5  g05295(.A(new_n7643), .B(new_n2544), .Y(new_n7644));
  xor_4  g05296(.A(new_n7643), .B(new_n2507), .Y(new_n7645));
  xor_4  g05297(.A(new_n7611), .B(new_n7602), .Y(new_n7646));
  not_8  g05298(.A(new_n7646), .Y(new_n7647));
  nor_5  g05299(.A(new_n7647), .B(new_n2510), .Y(new_n7648));
  xor_4  g05300(.A(new_n7609), .B(new_n7604), .Y(new_n7649));
  nand_5 g05301(.A(new_n7649), .B(new_n2516), .Y(new_n7650));
  nand_5 g05302(.A(new_n3815), .B(pi569), .Y(new_n7651));
  or_6   g05303(.A(new_n7651), .B(new_n2527), .Y(new_n7652));
  nand_5 g05304(.A(new_n7652), .B(new_n7608), .Y(new_n7653));
  nand_5 g05305(.A(new_n7653), .B(new_n2522), .Y(new_n7654));
  or_6   g05306(.A(new_n7651), .B(new_n2523), .Y(new_n7655));
  nand_5 g05307(.A(new_n7607), .B(new_n2523), .Y(new_n7656));
  nand_5 g05308(.A(new_n7656), .B(new_n7655), .Y(new_n7657));
  xor_4  g05309(.A(new_n7657), .B(new_n7606), .Y(new_n7658));
  nand_5 g05310(.A(new_n7658), .B(new_n2527), .Y(new_n7659));
  nor_5  g05311(.A(new_n7659), .B(new_n7655), .Y(new_n7660));
  nor_5  g05312(.A(new_n7658), .B(new_n2527), .Y(new_n7661));
  nor_5  g05313(.A(new_n7661), .B(new_n7660), .Y(new_n7662));
  nand_5 g05314(.A(new_n7662), .B(new_n7654), .Y(new_n7663));
  nand_5 g05315(.A(new_n7663), .B(new_n7650), .Y(new_n7664));
  or_6   g05316(.A(new_n7649), .B(new_n2516), .Y(new_n7665));
  nand_5 g05317(.A(new_n7665), .B(new_n7664), .Y(new_n7666));
  xor_4  g05318(.A(new_n7646), .B(new_n2510), .Y(new_n7667));
  nor_5  g05319(.A(new_n7667), .B(new_n7666), .Y(new_n7668));
  nor_5  g05320(.A(new_n7668), .B(new_n7648), .Y(new_n7669));
  nor_5  g05321(.A(new_n7669), .B(new_n7645), .Y(new_n7670));
  nor_5  g05322(.A(new_n7670), .B(new_n7644), .Y(new_n7671));
  nand_5 g05323(.A(new_n7671), .B(new_n7642), .Y(new_n7672));
  nand_5 g05324(.A(new_n7672), .B(new_n7641), .Y(new_n7673));
  nor_5  g05325(.A(new_n7673), .B(new_n7639), .Y(new_n7674));
  or_6   g05326(.A(new_n7674), .B(new_n7638), .Y(new_n7675));
  xor_4  g05327(.A(new_n7634), .B(new_n7632), .Y(new_n7676));
  nand_5 g05328(.A(new_n7676), .B(new_n7675), .Y(new_n7677));
  nand_5 g05329(.A(new_n7677), .B(new_n7635), .Y(new_n7678));
  xor_4  g05330(.A(new_n7630), .B(new_n7628), .Y(new_n7679));
  nand_5 g05331(.A(new_n7679), .B(new_n7678), .Y(new_n7680));
  nand_5 g05332(.A(new_n7680), .B(new_n7631), .Y(new_n7681));
  xor_4  g05333(.A(new_n7626), .B(new_n7589), .Y(new_n7682));
  and_6  g05334(.A(new_n7682), .B(new_n7681), .Y(new_n7683));
  nor_5  g05335(.A(new_n7683), .B(new_n7627), .Y(new_n7684));
  nand_5 g05336(.A(new_n7684), .B(new_n7587), .Y(new_n7685));
  nand_5 g05337(.A(new_n7685), .B(new_n7581), .Y(new_n7686));
  xnor_4 g05338(.A(new_n7684), .B(new_n7587), .Y(new_n7687));
  not_8  g05339(.A(new_n7687), .Y(new_n7688));
  nand_5 g05340(.A(pi582), .B(new_n7590), .Y(new_n7689));
  nand_5 g05341(.A(new_n7625), .B(new_n7591), .Y(new_n7690));
  nand_5 g05342(.A(new_n7690), .B(new_n7689), .Y(new_n7691));
  nor_5  g05343(.A(new_n7691), .B(new_n7585), .Y(new_n7692));
  or_6   g05344(.A(new_n7692), .B(new_n7688), .Y(new_n7693));
  nand_5 g05345(.A(new_n7693), .B(new_n7686), .Y(new_n7694));
  nor_5  g05346(.A(new_n7684), .B(new_n7587), .Y(new_n7695));
  nand_5 g05347(.A(new_n7695), .B(new_n7581), .Y(new_n7696));
  nand_5 g05348(.A(new_n7696), .B(new_n7586), .Y(new_n7697));
  nand_5 g05349(.A(new_n7697), .B(new_n7691), .Y(new_n7698));
  nand_5 g05350(.A(new_n7698), .B(new_n7694), .Y(po0035));
  not_8  g05351(.A(pi121), .Y(new_n7700));
  nand_5 g05352(.A(pi769), .B(new_n7700), .Y(new_n7701));
  xor_4  g05353(.A(pi769), .B(new_n7700), .Y(new_n7702));
  not_8  g05354(.A(pi066), .Y(new_n7703));
  nand_5 g05355(.A(pi275), .B(new_n7703), .Y(new_n7704));
  xor_4  g05356(.A(pi275), .B(new_n7703), .Y(new_n7705));
  nand_5 g05357(.A(pi459), .B(new_n6005), .Y(new_n7706));
  xor_4  g05358(.A(pi459), .B(new_n6005), .Y(new_n7707));
  nand_5 g05359(.A(pi530), .B(new_n5942), .Y(new_n7708));
  xor_4  g05360(.A(pi530), .B(new_n5942), .Y(new_n7709));
  nand_5 g05361(.A(pi712), .B(new_n5947), .Y(new_n7710));
  xor_4  g05362(.A(pi712), .B(new_n5947), .Y(new_n7711));
  not_8  g05363(.A(pi019), .Y(new_n7712));
  nand_5 g05364(.A(pi511), .B(new_n7712), .Y(new_n7713));
  xor_4  g05365(.A(pi511), .B(new_n7712), .Y(new_n7714));
  not_8  g05366(.A(pi628), .Y(new_n7715));
  nand_5 g05367(.A(new_n7715), .B(pi353), .Y(new_n7716));
  not_8  g05368(.A(new_n7716), .Y(new_n7717));
  xor_4  g05369(.A(pi628), .B(new_n6579), .Y(new_n7718));
  not_8  g05370(.A(new_n7718), .Y(new_n7719));
  not_8  g05371(.A(pi475), .Y(new_n7720));
  nor_5  g05372(.A(pi830), .B(new_n7720), .Y(new_n7721));
  xor_4  g05373(.A(pi830), .B(new_n7720), .Y(new_n7722));
  not_8  g05374(.A(new_n7722), .Y(new_n7723));
  nor_5  g05375(.A(new_n5768), .B(pi696), .Y(new_n7724));
  xor_4  g05376(.A(pi797), .B(new_n5953), .Y(new_n7725));
  nand_5 g05377(.A(new_n7725), .B(pi751), .Y(new_n7726));
  nor_5  g05378(.A(new_n7726), .B(pi220), .Y(new_n7727));
  nor_5  g05379(.A(new_n7727), .B(new_n7724), .Y(new_n7728));
  nor_5  g05380(.A(new_n7728), .B(new_n7723), .Y(new_n7729));
  nor_5  g05381(.A(new_n7729), .B(new_n7721), .Y(new_n7730));
  nor_5  g05382(.A(new_n7730), .B(new_n7719), .Y(new_n7731));
  nor_5  g05383(.A(new_n7731), .B(new_n7717), .Y(new_n7732));
  not_8  g05384(.A(new_n7732), .Y(new_n7733));
  nand_5 g05385(.A(new_n7733), .B(new_n7714), .Y(new_n7734));
  nand_5 g05386(.A(new_n7734), .B(new_n7713), .Y(new_n7735));
  nand_5 g05387(.A(new_n7735), .B(new_n7711), .Y(new_n7736));
  nand_5 g05388(.A(new_n7736), .B(new_n7710), .Y(new_n7737));
  nand_5 g05389(.A(new_n7737), .B(new_n7709), .Y(new_n7738));
  nand_5 g05390(.A(new_n7738), .B(new_n7708), .Y(new_n7739));
  nand_5 g05391(.A(new_n7739), .B(new_n7707), .Y(new_n7740));
  nand_5 g05392(.A(new_n7740), .B(new_n7706), .Y(new_n7741));
  nand_5 g05393(.A(new_n7741), .B(new_n7705), .Y(new_n7742));
  nand_5 g05394(.A(new_n7742), .B(new_n7704), .Y(new_n7743));
  nand_5 g05395(.A(new_n7743), .B(new_n7702), .Y(new_n7744));
  nand_5 g05396(.A(new_n7744), .B(new_n7701), .Y(new_n7745));
  nand_5 g05397(.A(pi697), .B(new_n3697), .Y(new_n7746));
  xor_4  g05398(.A(pi697), .B(new_n3697), .Y(new_n7747));
  nand_5 g05399(.A(pi452), .B(new_n3525), .Y(new_n7748));
  xor_4  g05400(.A(pi452), .B(new_n3525), .Y(new_n7749));
  nand_5 g05401(.A(new_n3530), .B(pi046), .Y(new_n7750));
  not_8  g05402(.A(pi046), .Y(new_n7751));
  xor_4  g05403(.A(pi507), .B(new_n7751), .Y(new_n7752));
  nand_5 g05404(.A(pi439), .B(new_n2468), .Y(new_n7753));
  xor_4  g05405(.A(pi439), .B(new_n2468), .Y(new_n7754));
  nand_5 g05406(.A(pi822), .B(new_n5181), .Y(new_n7755));
  xor_4  g05407(.A(pi822), .B(new_n5181), .Y(new_n7756));
  nand_5 g05408(.A(new_n2474), .B(pi100), .Y(new_n7757));
  not_8  g05409(.A(pi100), .Y(new_n7758));
  xor_4  g05410(.A(pi316), .B(new_n7758), .Y(new_n7759));
  nand_5 g05411(.A(pi117), .B(new_n2478), .Y(new_n7760));
  nand_5 g05412(.A(pi514), .B(new_n2482), .Y(new_n7761));
  not_8  g05413(.A(new_n7761), .Y(new_n7762));
  xor_4  g05414(.A(pi514), .B(new_n2482), .Y(new_n7763));
  not_8  g05415(.A(new_n7763), .Y(new_n7764));
  nand_5 g05416(.A(pi612), .B(new_n2360), .Y(new_n7765));
  nand_5 g05417(.A(new_n3552), .B(pi369), .Y(new_n7766));
  nand_5 g05418(.A(pi438), .B(new_n3641), .Y(new_n7767));
  nand_5 g05419(.A(new_n7767), .B(new_n7766), .Y(new_n7768));
  nand_5 g05420(.A(new_n7768), .B(new_n7765), .Y(new_n7769));
  nor_5  g05421(.A(new_n7769), .B(new_n7764), .Y(new_n7770));
  nor_5  g05422(.A(new_n7770), .B(new_n7762), .Y(new_n7771));
  xor_4  g05423(.A(pi117), .B(pi102), .Y(new_n7772));
  or_6   g05424(.A(new_n7772), .B(new_n7771), .Y(new_n7773));
  nand_5 g05425(.A(new_n7773), .B(new_n7760), .Y(new_n7774));
  nand_5 g05426(.A(new_n7774), .B(new_n7759), .Y(new_n7775));
  nand_5 g05427(.A(new_n7775), .B(new_n7757), .Y(new_n7776));
  nand_5 g05428(.A(new_n7776), .B(new_n7756), .Y(new_n7777));
  nand_5 g05429(.A(new_n7777), .B(new_n7755), .Y(new_n7778));
  nand_5 g05430(.A(new_n7778), .B(new_n7754), .Y(new_n7779));
  nand_5 g05431(.A(new_n7779), .B(new_n7753), .Y(new_n7780));
  nand_5 g05432(.A(new_n7780), .B(new_n7752), .Y(new_n7781));
  nand_5 g05433(.A(new_n7781), .B(new_n7750), .Y(new_n7782));
  nand_5 g05434(.A(new_n7782), .B(new_n7749), .Y(new_n7783));
  nand_5 g05435(.A(new_n7783), .B(new_n7748), .Y(new_n7784));
  nand_5 g05436(.A(new_n7784), .B(new_n7747), .Y(new_n7785));
  nand_5 g05437(.A(new_n7785), .B(new_n7746), .Y(new_n7786));
  xor_4  g05438(.A(new_n7786), .B(new_n7745), .Y(new_n7787));
  xor_4  g05439(.A(new_n7743), .B(new_n7702), .Y(new_n7788));
  not_8  g05440(.A(new_n7788), .Y(new_n7789));
  xor_4  g05441(.A(new_n7741), .B(new_n7705), .Y(new_n7790));
  not_8  g05442(.A(new_n7790), .Y(new_n7791));
  xnor_4 g05443(.A(new_n7782), .B(new_n7749), .Y(new_n7792));
  nor_5  g05444(.A(new_n7792), .B(new_n7791), .Y(new_n7793));
  xor_4  g05445(.A(new_n7792), .B(new_n7791), .Y(new_n7794));
  not_8  g05446(.A(new_n7794), .Y(new_n7795));
  xor_4  g05447(.A(new_n7739), .B(new_n7707), .Y(new_n7796));
  not_8  g05448(.A(new_n7796), .Y(new_n7797));
  xnor_4 g05449(.A(new_n7780), .B(new_n7752), .Y(new_n7798));
  nor_5  g05450(.A(new_n7798), .B(new_n7797), .Y(new_n7799));
  xor_4  g05451(.A(new_n7798), .B(new_n7797), .Y(new_n7800));
  not_8  g05452(.A(new_n7800), .Y(new_n7801));
  xor_4  g05453(.A(new_n7737), .B(new_n7709), .Y(new_n7802));
  xor_4  g05454(.A(new_n7778), .B(new_n7754), .Y(new_n7803));
  or_6   g05455(.A(new_n7803), .B(new_n7802), .Y(new_n7804));
  xor_4  g05456(.A(new_n7803), .B(new_n7802), .Y(new_n7805));
  xor_4  g05457(.A(new_n7735), .B(new_n7711), .Y(new_n7806));
  not_8  g05458(.A(new_n7806), .Y(new_n7807));
  xor_4  g05459(.A(new_n7774), .B(new_n7759), .Y(new_n7808));
  not_8  g05460(.A(new_n7808), .Y(new_n7809));
  xor_4  g05461(.A(new_n7732), .B(new_n7714), .Y(new_n7810));
  nand_5 g05462(.A(new_n7810), .B(new_n7809), .Y(new_n7811));
  xor_4  g05463(.A(new_n7730), .B(new_n7719), .Y(new_n7812));
  not_8  g05464(.A(new_n7812), .Y(new_n7813));
  xor_4  g05465(.A(new_n7728), .B(new_n7723), .Y(new_n7814));
  xor_4  g05466(.A(new_n7769), .B(new_n7763), .Y(new_n7815));
  not_8  g05467(.A(new_n7815), .Y(new_n7816));
  nand_5 g05468(.A(new_n7816), .B(new_n7814), .Y(new_n7817));
  nand_5 g05469(.A(new_n5765), .B(pi220), .Y(new_n7818));
  xor_4  g05470(.A(pi438), .B(new_n3641), .Y(new_n7819));
  nand_5 g05471(.A(pi751), .B(new_n5778), .Y(new_n7820));
  nand_5 g05472(.A(new_n7820), .B(new_n7818), .Y(new_n7821));
  nand_5 g05473(.A(new_n7821), .B(new_n7819), .Y(new_n7822));
  nand_5 g05474(.A(new_n7822), .B(new_n7767), .Y(new_n7823));
  nand_5 g05475(.A(new_n7823), .B(new_n7818), .Y(new_n7824));
  not_8  g05476(.A(new_n7725), .Y(new_n7825));
  nand_5 g05477(.A(new_n7766), .B(new_n7765), .Y(new_n7826));
  nand_5 g05478(.A(new_n7826), .B(new_n7825), .Y(new_n7827));
  nor_5  g05479(.A(new_n7827), .B(new_n7824), .Y(new_n7828));
  nand_5 g05480(.A(new_n7820), .B(new_n7725), .Y(new_n7829));
  nor_5  g05481(.A(pi438), .B(new_n3641), .Y(new_n7830));
  not_8  g05482(.A(new_n7826), .Y(new_n7831));
  nor_5  g05483(.A(new_n7831), .B(new_n7830), .Y(new_n7832));
  nor_5  g05484(.A(new_n7832), .B(new_n7818), .Y(new_n7833));
  nor_5  g05485(.A(new_n7833), .B(new_n7829), .Y(new_n7834));
  not_8  g05486(.A(new_n7818), .Y(new_n7835));
  nand_5 g05487(.A(new_n7835), .B(new_n7825), .Y(new_n7836));
  nand_5 g05488(.A(new_n7836), .B(new_n7726), .Y(new_n7837));
  nand_5 g05489(.A(new_n7831), .B(new_n2420), .Y(new_n7838));
  nor_5  g05490(.A(new_n7838), .B(new_n7837), .Y(new_n7839));
  nand_5 g05491(.A(new_n7831), .B(new_n7819), .Y(new_n7840));
  not_8  g05492(.A(new_n7840), .Y(new_n7841));
  or_6   g05493(.A(new_n7841), .B(new_n7839), .Y(new_n7842));
  nor_5  g05494(.A(new_n7842), .B(new_n7834), .Y(new_n7843));
  not_8  g05495(.A(new_n7843), .Y(new_n7844));
  nor_5  g05496(.A(new_n7844), .B(new_n7828), .Y(new_n7845));
  xor_4  g05497(.A(new_n7815), .B(new_n7814), .Y(new_n7846));
  or_6   g05498(.A(new_n7846), .B(new_n7845), .Y(new_n7847));
  and_6  g05499(.A(new_n7847), .B(new_n7817), .Y(new_n7848));
  nand_5 g05500(.A(new_n7848), .B(new_n7813), .Y(new_n7849));
  xor_4  g05501(.A(new_n7848), .B(new_n7812), .Y(new_n7850));
  xor_4  g05502(.A(new_n7772), .B(new_n7771), .Y(new_n7851));
  or_6   g05503(.A(new_n7851), .B(new_n7850), .Y(new_n7852));
  nand_5 g05504(.A(new_n7852), .B(new_n7849), .Y(new_n7853));
  xor_4  g05505(.A(new_n7810), .B(new_n7808), .Y(new_n7854));
  not_8  g05506(.A(new_n7854), .Y(new_n7855));
  nand_5 g05507(.A(new_n7855), .B(new_n7853), .Y(new_n7856));
  nand_5 g05508(.A(new_n7856), .B(new_n7811), .Y(new_n7857));
  nand_5 g05509(.A(new_n7857), .B(new_n7807), .Y(new_n7858));
  xor_4  g05510(.A(new_n7776), .B(new_n7756), .Y(new_n7859));
  xor_4  g05511(.A(new_n7857), .B(new_n7806), .Y(new_n7860));
  or_6   g05512(.A(new_n7860), .B(new_n7859), .Y(new_n7861));
  nand_5 g05513(.A(new_n7861), .B(new_n7858), .Y(new_n7862));
  nand_5 g05514(.A(new_n7862), .B(new_n7805), .Y(new_n7863));
  nand_5 g05515(.A(new_n7863), .B(new_n7804), .Y(new_n7864));
  nor_5  g05516(.A(new_n7864), .B(new_n7801), .Y(new_n7865));
  nor_5  g05517(.A(new_n7865), .B(new_n7799), .Y(new_n7866));
  nor_5  g05518(.A(new_n7866), .B(new_n7795), .Y(new_n7867));
  nor_5  g05519(.A(new_n7867), .B(new_n7793), .Y(new_n7868));
  nand_5 g05520(.A(new_n7868), .B(new_n7789), .Y(new_n7869));
  xor_4  g05521(.A(new_n7784), .B(new_n7747), .Y(new_n7870));
  xor_4  g05522(.A(new_n7868), .B(new_n7788), .Y(new_n7871));
  or_6   g05523(.A(new_n7871), .B(new_n7870), .Y(new_n7872));
  nand_5 g05524(.A(new_n7872), .B(new_n7869), .Y(new_n7873));
  xnor_4 g05525(.A(new_n7873), .B(new_n7787), .Y(new_n7874));
  xor_4  g05526(.A(new_n7866), .B(new_n7794), .Y(new_n7875));
  nand_5 g05527(.A(new_n4839), .B(pi650), .Y(new_n7876));
  nand_5 g05528(.A(pi812), .B(new_n3473), .Y(new_n7877));
  and_6  g05529(.A(new_n7877), .B(new_n7876), .Y(new_n7878));
  nand_5 g05530(.A(new_n5918), .B(pi547), .Y(new_n7879));
  xor_4  g05531(.A(pi616), .B(new_n4842), .Y(new_n7880));
  nand_5 g05532(.A(new_n4828), .B(pi236), .Y(new_n7881));
  xor_4  g05533(.A(pi441), .B(new_n4754), .Y(new_n7882));
  nand_5 g05534(.A(pi375), .B(new_n3484), .Y(new_n7883));
  xor_4  g05535(.A(pi375), .B(new_n3484), .Y(new_n7884));
  nand_5 g05536(.A(pi427), .B(new_n4904), .Y(new_n7885));
  xor_4  g05537(.A(pi427), .B(new_n4904), .Y(new_n7886));
  nand_5 g05538(.A(new_n4795), .B(pi237), .Y(new_n7887));
  xor_4  g05539(.A(pi681), .B(new_n4763), .Y(new_n7888));
  nand_5 g05540(.A(pi599), .B(new_n3489), .Y(new_n7889));
  xor_4  g05541(.A(pi599), .B(new_n3489), .Y(new_n7890));
  nand_5 g05542(.A(new_n3629), .B(pi091), .Y(new_n7891));
  nand_5 g05543(.A(new_n3493), .B(pi482), .Y(new_n7892));
  not_8  g05544(.A(new_n7892), .Y(new_n7893));
  xor_4  g05545(.A(pi787), .B(new_n4770), .Y(new_n7894));
  nand_5 g05546(.A(new_n7894), .B(new_n7893), .Y(new_n7895));
  nand_5 g05547(.A(new_n7895), .B(new_n7891), .Y(new_n7896));
  nand_5 g05548(.A(new_n7896), .B(new_n7890), .Y(new_n7897));
  nand_5 g05549(.A(new_n7897), .B(new_n7889), .Y(new_n7898));
  nand_5 g05550(.A(new_n7898), .B(new_n7888), .Y(new_n7899));
  nand_5 g05551(.A(new_n7899), .B(new_n7887), .Y(new_n7900));
  nand_5 g05552(.A(new_n7900), .B(new_n7886), .Y(new_n7901));
  nand_5 g05553(.A(new_n7901), .B(new_n7885), .Y(new_n7902));
  nand_5 g05554(.A(new_n7902), .B(new_n7884), .Y(new_n7903));
  nand_5 g05555(.A(new_n7903), .B(new_n7883), .Y(new_n7904));
  nand_5 g05556(.A(new_n7904), .B(new_n7882), .Y(new_n7905));
  nand_5 g05557(.A(new_n7905), .B(new_n7881), .Y(new_n7906));
  nand_5 g05558(.A(new_n7906), .B(new_n7880), .Y(new_n7907));
  nand_5 g05559(.A(new_n7907), .B(new_n7879), .Y(new_n7908));
  xor_4  g05560(.A(new_n7908), .B(new_n7878), .Y(new_n7909));
  not_8  g05561(.A(new_n7909), .Y(new_n7910));
  nor_5  g05562(.A(new_n7910), .B(new_n7875), .Y(new_n7911));
  xor_4  g05563(.A(new_n7909), .B(new_n7875), .Y(new_n7912));
  xor_4  g05564(.A(new_n7906), .B(new_n7880), .Y(new_n7913));
  xor_4  g05565(.A(new_n7904), .B(new_n7882), .Y(new_n7914));
  xor_4  g05566(.A(new_n7902), .B(new_n7884), .Y(new_n7915));
  not_8  g05567(.A(new_n7915), .Y(new_n7916));
  xor_4  g05568(.A(new_n7900), .B(new_n7886), .Y(new_n7917));
  not_8  g05569(.A(new_n7917), .Y(new_n7918));
  xor_4  g05570(.A(new_n7846), .B(new_n7845), .Y(new_n7919));
  not_8  g05571(.A(new_n7919), .Y(new_n7920));
  xor_4  g05572(.A(new_n7894), .B(new_n7893), .Y(new_n7921));
  not_8  g05573(.A(new_n7921), .Y(new_n7922));
  not_8  g05574(.A(pi482), .Y(new_n7923));
  xor_4  g05575(.A(pi670), .B(new_n7923), .Y(new_n7924));
  xor_4  g05576(.A(new_n7821), .B(new_n7819), .Y(new_n7925));
  nor_5  g05577(.A(new_n7925), .B(new_n7924), .Y(new_n7926));
  nand_5 g05578(.A(new_n7926), .B(new_n7922), .Y(new_n7927));
  nand_5 g05579(.A(new_n7830), .B(new_n7835), .Y(new_n7928));
  nand_5 g05580(.A(new_n7928), .B(new_n7824), .Y(new_n7929));
  xor_4  g05581(.A(new_n7826), .B(new_n7725), .Y(new_n7930));
  xor_4  g05582(.A(new_n7930), .B(new_n7929), .Y(new_n7931));
  xor_4  g05583(.A(new_n7926), .B(new_n7921), .Y(new_n7932));
  or_6   g05584(.A(new_n7932), .B(new_n7931), .Y(new_n7933));
  nand_5 g05585(.A(new_n7933), .B(new_n7927), .Y(new_n7934));
  nand_5 g05586(.A(new_n7934), .B(new_n7920), .Y(new_n7935));
  xor_4  g05587(.A(new_n7896), .B(new_n7890), .Y(new_n7936));
  xor_4  g05588(.A(new_n7934), .B(new_n7919), .Y(new_n7937));
  or_6   g05589(.A(new_n7937), .B(new_n7936), .Y(new_n7938));
  nand_5 g05590(.A(new_n7938), .B(new_n7935), .Y(new_n7939));
  not_8  g05591(.A(new_n7851), .Y(new_n7940));
  xor_4  g05592(.A(new_n7940), .B(new_n7850), .Y(new_n7941));
  not_8  g05593(.A(new_n7941), .Y(new_n7942));
  nand_5 g05594(.A(new_n7942), .B(new_n7939), .Y(new_n7943));
  xor_4  g05595(.A(new_n7898), .B(new_n7888), .Y(new_n7944));
  not_8  g05596(.A(new_n7944), .Y(new_n7945));
  xor_4  g05597(.A(new_n7942), .B(new_n7939), .Y(new_n7946));
  nand_5 g05598(.A(new_n7946), .B(new_n7945), .Y(new_n7947));
  nand_5 g05599(.A(new_n7947), .B(new_n7943), .Y(new_n7948));
  nand_5 g05600(.A(new_n7948), .B(new_n7918), .Y(new_n7949));
  xor_4  g05601(.A(new_n7854), .B(new_n7853), .Y(new_n7950));
  xor_4  g05602(.A(new_n7948), .B(new_n7917), .Y(new_n7951));
  or_6   g05603(.A(new_n7951), .B(new_n7950), .Y(new_n7952));
  nand_5 g05604(.A(new_n7952), .B(new_n7949), .Y(new_n7953));
  nor_5  g05605(.A(new_n7953), .B(new_n7916), .Y(new_n7954));
  xor_4  g05606(.A(new_n7860), .B(new_n7859), .Y(new_n7955));
  xor_4  g05607(.A(new_n7953), .B(new_n7915), .Y(new_n7956));
  nor_5  g05608(.A(new_n7956), .B(new_n7955), .Y(new_n7957));
  or_6   g05609(.A(new_n7957), .B(new_n7954), .Y(new_n7958));
  nand_5 g05610(.A(new_n7958), .B(new_n7914), .Y(new_n7959));
  xor_4  g05611(.A(new_n7862), .B(new_n7805), .Y(new_n7960));
  xnor_4 g05612(.A(new_n7958), .B(new_n7914), .Y(new_n7961));
  or_6   g05613(.A(new_n7961), .B(new_n7960), .Y(new_n7962));
  nand_5 g05614(.A(new_n7962), .B(new_n7959), .Y(new_n7963));
  or_6   g05615(.A(new_n7963), .B(new_n7913), .Y(new_n7964));
  xor_4  g05616(.A(new_n7963), .B(new_n7913), .Y(new_n7965));
  xor_4  g05617(.A(new_n7864), .B(new_n7800), .Y(new_n7966));
  nand_5 g05618(.A(new_n7966), .B(new_n7965), .Y(new_n7967));
  nand_5 g05619(.A(new_n7967), .B(new_n7964), .Y(new_n7968));
  nor_5  g05620(.A(new_n7968), .B(new_n7912), .Y(new_n7969));
  or_6   g05621(.A(new_n7969), .B(new_n7911), .Y(new_n7970));
  xor_4  g05622(.A(new_n7871), .B(new_n7870), .Y(new_n7971));
  not_8  g05623(.A(new_n7971), .Y(new_n7972));
  nand_5 g05624(.A(new_n7972), .B(new_n7970), .Y(new_n7973));
  nand_5 g05625(.A(pi315), .B(new_n3423), .Y(new_n7974));
  and_6  g05626(.A(new_n7974), .B(new_n7973), .Y(new_n7975));
  nand_5 g05627(.A(new_n7908), .B(new_n7876), .Y(new_n7976));
  nand_5 g05628(.A(new_n7976), .B(new_n7877), .Y(new_n7977));
  not_8  g05629(.A(new_n7977), .Y(new_n7978));
  not_8  g05630(.A(new_n7974), .Y(new_n7979));
  nand_5 g05631(.A(new_n7979), .B(new_n7970), .Y(new_n7980));
  nand_5 g05632(.A(new_n7980), .B(new_n7978), .Y(new_n7981));
  nor_5  g05633(.A(new_n7981), .B(new_n7975), .Y(new_n7982));
  nor_5  g05634(.A(new_n7972), .B(new_n7970), .Y(new_n7983));
  nand_5 g05635(.A(new_n4858), .B(pi303), .Y(new_n7984));
  not_8  g05636(.A(new_n7984), .Y(new_n7985));
  or_6   g05637(.A(new_n7985), .B(new_n7983), .Y(new_n7986));
  nor_5  g05638(.A(new_n7984), .B(new_n7970), .Y(new_n7987));
  nor_5  g05639(.A(new_n7987), .B(new_n7978), .Y(new_n7988));
  nand_5 g05640(.A(new_n7988), .B(new_n7986), .Y(new_n7989));
  xor_4  g05641(.A(new_n7972), .B(new_n7970), .Y(new_n7990));
  nand_5 g05642(.A(new_n7979), .B(new_n7977), .Y(new_n7991));
  nand_5 g05643(.A(new_n7978), .B(new_n7985), .Y(new_n7992));
  nand_5 g05644(.A(new_n7992), .B(new_n7991), .Y(new_n7993));
  not_8  g05645(.A(new_n7993), .Y(new_n7994));
  nand_5 g05646(.A(new_n7994), .B(new_n7990), .Y(new_n7995));
  nand_5 g05647(.A(new_n7995), .B(new_n7989), .Y(new_n7996));
  nor_5  g05648(.A(new_n7996), .B(new_n7982), .Y(new_n7997));
  xnor_4 g05649(.A(new_n7997), .B(new_n7874), .Y(po0036));
  nand_5 g05650(.A(pi716), .B(pi465), .Y(new_n7999));
  xor_4  g05651(.A(pi716), .B(pi465), .Y(new_n8000));
  nand_5 g05652(.A(pi722), .B(pi368), .Y(new_n8001));
  xor_4  g05653(.A(pi722), .B(pi368), .Y(new_n8002));
  nand_5 g05654(.A(pi505), .B(pi336), .Y(new_n8003));
  not_8  g05655(.A(pi336), .Y(new_n8004));
  not_8  g05656(.A(pi505), .Y(new_n8005));
  nand_5 g05657(.A(new_n8005), .B(new_n8004), .Y(new_n8006));
  nand_5 g05658(.A(pi473), .B(pi470), .Y(new_n8007));
  not_8  g05659(.A(pi470), .Y(new_n8008));
  nand_5 g05660(.A(new_n4382), .B(new_n8008), .Y(new_n8009));
  nand_5 g05661(.A(pi372), .B(pi248), .Y(new_n8010));
  xor_4  g05662(.A(pi372), .B(pi248), .Y(new_n8011));
  nand_5 g05663(.A(pi125), .B(pi001), .Y(new_n8012));
  xor_4  g05664(.A(pi125), .B(pi001), .Y(new_n8013));
  not_8  g05665(.A(new_n8013), .Y(new_n8014));
  not_8  g05666(.A(pi050), .Y(new_n8015));
  nand_5 g05667(.A(new_n4395), .B(new_n8015), .Y(new_n8016));
  xor_4  g05668(.A(pi618), .B(pi050), .Y(new_n8017));
  not_8  g05669(.A(pi192), .Y(new_n8018));
  not_8  g05670(.A(pi262), .Y(new_n8019));
  nand_5 g05671(.A(new_n8019), .B(new_n8018), .Y(new_n8020));
  not_8  g05672(.A(new_n8020), .Y(new_n8021));
  xor_4  g05673(.A(pi262), .B(pi192), .Y(new_n8022));
  not_8  g05674(.A(new_n8022), .Y(new_n8023));
  nor_5  g05675(.A(pi813), .B(pi326), .Y(new_n8024));
  not_8  g05676(.A(pi122), .Y(new_n8025));
  nor_5  g05677(.A(new_n8025), .B(new_n4405), .Y(new_n8026));
  not_8  g05678(.A(pi326), .Y(new_n8027));
  xor_4  g05679(.A(pi813), .B(new_n8027), .Y(new_n8028));
  nor_5  g05680(.A(new_n8028), .B(new_n8026), .Y(new_n8029));
  nor_5  g05681(.A(new_n8029), .B(new_n8024), .Y(new_n8030));
  nor_5  g05682(.A(new_n8030), .B(new_n8023), .Y(new_n8031));
  nor_5  g05683(.A(new_n8031), .B(new_n8021), .Y(new_n8032));
  not_8  g05684(.A(new_n8032), .Y(new_n8033));
  nand_5 g05685(.A(new_n8033), .B(new_n8017), .Y(new_n8034));
  nand_5 g05686(.A(new_n8034), .B(new_n8016), .Y(new_n8035));
  or_6   g05687(.A(new_n8035), .B(new_n8014), .Y(new_n8036));
  nand_5 g05688(.A(new_n8036), .B(new_n8012), .Y(new_n8037));
  nand_5 g05689(.A(new_n8037), .B(new_n8011), .Y(new_n8038));
  nand_5 g05690(.A(new_n8038), .B(new_n8010), .Y(new_n8039));
  nand_5 g05691(.A(new_n8039), .B(new_n8009), .Y(new_n8040));
  nand_5 g05692(.A(new_n8040), .B(new_n8007), .Y(new_n8041));
  nand_5 g05693(.A(new_n8041), .B(new_n8006), .Y(new_n8042));
  nand_5 g05694(.A(new_n8042), .B(new_n8003), .Y(new_n8043));
  nand_5 g05695(.A(new_n8043), .B(new_n8002), .Y(new_n8044));
  nand_5 g05696(.A(new_n8044), .B(new_n8001), .Y(new_n8045));
  nand_5 g05697(.A(new_n8045), .B(new_n8000), .Y(new_n8046));
  nand_5 g05698(.A(new_n8046), .B(new_n7999), .Y(new_n8047));
  not_8  g05699(.A(new_n8047), .Y(new_n8048));
  xor_4  g05700(.A(new_n8045), .B(new_n8000), .Y(new_n8049));
  not_8  g05701(.A(new_n8049), .Y(new_n8050));
  nand_5 g05702(.A(new_n8050), .B(pi700), .Y(new_n8051));
  not_8  g05703(.A(pi700), .Y(new_n8052));
  xor_4  g05704(.A(new_n8049), .B(new_n8052), .Y(new_n8053));
  xor_4  g05705(.A(new_n8043), .B(new_n8002), .Y(new_n8054));
  not_8  g05706(.A(pi258), .Y(new_n8055));
  nand_5 g05707(.A(new_n8009), .B(new_n8007), .Y(new_n8056));
  xor_4  g05708(.A(new_n8056), .B(new_n8039), .Y(new_n8057));
  not_8  g05709(.A(new_n8057), .Y(new_n8058));
  xor_4  g05710(.A(new_n8037), .B(new_n8011), .Y(new_n8059));
  xor_4  g05711(.A(new_n8035), .B(new_n8014), .Y(new_n8060));
  not_8  g05712(.A(new_n8060), .Y(new_n8061));
  not_8  g05713(.A(pi698), .Y(new_n8062));
  not_8  g05714(.A(pi474), .Y(new_n8063));
  not_8  g05715(.A(new_n2553), .Y(new_n8064));
  nor_5  g05716(.A(new_n8064), .B(pi149), .Y(new_n8065));
  nand_5 g05717(.A(new_n8065), .B(new_n8063), .Y(new_n8066));
  xor_4  g05718(.A(new_n8065), .B(new_n8063), .Y(new_n8067));
  not_8  g05719(.A(new_n8067), .Y(new_n8068));
  xor_4  g05720(.A(new_n8028), .B(new_n8026), .Y(new_n8069));
  or_6   g05721(.A(new_n8069), .B(new_n8068), .Y(new_n8070));
  nand_5 g05722(.A(new_n8070), .B(new_n8066), .Y(new_n8071));
  xor_4  g05723(.A(new_n8030), .B(new_n8023), .Y(new_n8072));
  not_8  g05724(.A(new_n8072), .Y(new_n8073));
  nand_5 g05725(.A(new_n8073), .B(new_n8071), .Y(new_n8074));
  not_8  g05726(.A(pi515), .Y(new_n8075));
  or_6   g05727(.A(new_n8073), .B(new_n8071), .Y(new_n8076));
  nand_5 g05728(.A(new_n8076), .B(new_n8075), .Y(new_n8077));
  nand_5 g05729(.A(new_n8077), .B(new_n8074), .Y(new_n8078));
  or_6   g05730(.A(new_n8078), .B(new_n8062), .Y(new_n8079));
  xor_4  g05731(.A(new_n8078), .B(new_n8062), .Y(new_n8080));
  xor_4  g05732(.A(new_n8032), .B(new_n8017), .Y(new_n8081));
  not_8  g05733(.A(new_n8081), .Y(new_n8082));
  nand_5 g05734(.A(new_n8082), .B(new_n8080), .Y(new_n8083));
  nand_5 g05735(.A(new_n8083), .B(new_n8079), .Y(new_n8084));
  or_6   g05736(.A(new_n8084), .B(new_n8061), .Y(new_n8085));
  not_8  g05737(.A(pi075), .Y(new_n8086));
  xor_4  g05738(.A(new_n8084), .B(new_n8061), .Y(new_n8087));
  nand_5 g05739(.A(new_n8087), .B(new_n8086), .Y(new_n8088));
  nand_5 g05740(.A(new_n8088), .B(new_n8085), .Y(new_n8089));
  nand_5 g05741(.A(new_n8089), .B(new_n8059), .Y(new_n8090));
  not_8  g05742(.A(pi764), .Y(new_n8091));
  or_6   g05743(.A(new_n8089), .B(new_n8059), .Y(new_n8092));
  nand_5 g05744(.A(new_n8092), .B(new_n8091), .Y(new_n8093));
  nand_5 g05745(.A(new_n8093), .B(new_n8090), .Y(new_n8094));
  nor_5  g05746(.A(new_n8094), .B(new_n8058), .Y(new_n8095));
  xor_4  g05747(.A(new_n8094), .B(new_n8058), .Y(new_n8096));
  nand_5 g05748(.A(new_n8096), .B(pi516), .Y(new_n8097));
  not_8  g05749(.A(new_n8097), .Y(new_n8098));
  nor_5  g05750(.A(new_n8098), .B(new_n8095), .Y(new_n8099));
  nand_5 g05751(.A(new_n8099), .B(new_n8055), .Y(new_n8100));
  xor_4  g05752(.A(new_n8099), .B(pi258), .Y(new_n8101));
  nand_5 g05753(.A(new_n8006), .B(new_n8003), .Y(new_n8102));
  xor_4  g05754(.A(new_n8102), .B(new_n8041), .Y(new_n8103));
  or_6   g05755(.A(new_n8103), .B(new_n8101), .Y(new_n8104));
  nand_5 g05756(.A(new_n8104), .B(new_n8100), .Y(new_n8105));
  nand_5 g05757(.A(new_n8105), .B(new_n8054), .Y(new_n8106));
  not_8  g05758(.A(new_n8106), .Y(new_n8107));
  nor_5  g05759(.A(new_n8105), .B(new_n8054), .Y(new_n8108));
  nor_5  g05760(.A(new_n8108), .B(pi810), .Y(new_n8109));
  nor_5  g05761(.A(new_n8109), .B(new_n8107), .Y(new_n8110));
  nand_5 g05762(.A(new_n8110), .B(new_n8053), .Y(new_n8111));
  nand_5 g05763(.A(new_n8111), .B(new_n8051), .Y(new_n8112));
  nand_5 g05764(.A(new_n8112), .B(new_n8048), .Y(new_n8113));
  xor_4  g05765(.A(new_n8112), .B(new_n8047), .Y(new_n8114));
  xor_4  g05766(.A(pi542), .B(new_n5546), .Y(new_n8115));
  nand_5 g05767(.A(new_n5497), .B(pi748), .Y(new_n8116));
  not_8  g05768(.A(pi748), .Y(new_n8117));
  xor_4  g05769(.A(pi827), .B(new_n8117), .Y(new_n8118));
  nand_5 g05770(.A(new_n5499), .B(pi503), .Y(new_n8119));
  xor_4  g05771(.A(pi737), .B(new_n4280), .Y(new_n8120));
  nand_5 g05772(.A(pi780), .B(new_n5503), .Y(new_n8121));
  xor_4  g05773(.A(pi780), .B(new_n5503), .Y(new_n8122));
  nand_5 g05774(.A(new_n5507), .B(pi400), .Y(new_n8123));
  xor_4  g05775(.A(new_n5507), .B(pi400), .Y(new_n8124));
  nand_5 g05776(.A(new_n5511), .B(pi003), .Y(new_n8125));
  not_8  g05777(.A(pi003), .Y(new_n8126));
  xor_4  g05778(.A(pi128), .B(new_n8126), .Y(new_n8127));
  nand_5 g05779(.A(pi761), .B(new_n5513), .Y(new_n8128));
  xor_4  g05780(.A(pi761), .B(new_n5513), .Y(new_n8129));
  nand_5 g05781(.A(pi221), .B(new_n5517), .Y(new_n8130));
  xor_4  g05782(.A(pi221), .B(new_n5517), .Y(new_n8131));
  nand_5 g05783(.A(pi741), .B(new_n5520), .Y(new_n8132));
  xor_4  g05784(.A(pi741), .B(new_n5520), .Y(new_n8133));
  nand_5 g05785(.A(new_n8133), .B(new_n2557), .Y(new_n8134));
  nand_5 g05786(.A(new_n8134), .B(new_n8132), .Y(new_n8135));
  nand_5 g05787(.A(new_n8135), .B(new_n8131), .Y(new_n8136));
  nand_5 g05788(.A(new_n8136), .B(new_n8130), .Y(new_n8137));
  nand_5 g05789(.A(new_n8137), .B(new_n8129), .Y(new_n8138));
  nand_5 g05790(.A(new_n8138), .B(new_n8128), .Y(new_n8139));
  nand_5 g05791(.A(new_n8139), .B(new_n8127), .Y(new_n8140));
  nand_5 g05792(.A(new_n8140), .B(new_n8125), .Y(new_n8141));
  nand_5 g05793(.A(new_n8141), .B(new_n8124), .Y(new_n8142));
  nand_5 g05794(.A(new_n8142), .B(new_n8123), .Y(new_n8143));
  nand_5 g05795(.A(new_n8143), .B(new_n8122), .Y(new_n8144));
  nand_5 g05796(.A(new_n8144), .B(new_n8121), .Y(new_n8145));
  nand_5 g05797(.A(new_n8145), .B(new_n8120), .Y(new_n8146));
  nand_5 g05798(.A(new_n8146), .B(new_n8119), .Y(new_n8147));
  nand_5 g05799(.A(new_n8147), .B(new_n8118), .Y(new_n8148));
  nand_5 g05800(.A(new_n8148), .B(new_n8116), .Y(new_n8149));
  xor_4  g05801(.A(new_n8149), .B(new_n8115), .Y(new_n8150));
  xor_4  g05802(.A(new_n8147), .B(new_n8118), .Y(new_n8151));
  not_8  g05803(.A(pi310), .Y(new_n8152));
  not_8  g05804(.A(pi274), .Y(new_n8153));
  not_8  g05805(.A(pi398), .Y(new_n8154));
  xor_4  g05806(.A(new_n8139), .B(new_n8127), .Y(new_n8155));
  nand_5 g05807(.A(new_n8155), .B(new_n8154), .Y(new_n8156));
  xor_4  g05808(.A(new_n8155), .B(new_n8154), .Y(new_n8157));
  not_8  g05809(.A(pi639), .Y(new_n8158));
  xor_4  g05810(.A(new_n8137), .B(new_n8129), .Y(new_n8159));
  nand_5 g05811(.A(new_n8159), .B(new_n8158), .Y(new_n8160));
  xor_4  g05812(.A(new_n8159), .B(new_n8158), .Y(new_n8161));
  not_8  g05813(.A(pi754), .Y(new_n8162));
  not_8  g05814(.A(pi080), .Y(new_n8163));
  xor_4  g05815(.A(new_n8133), .B(new_n8163), .Y(new_n8164));
  not_8  g05816(.A(new_n8164), .Y(new_n8165));
  not_8  g05817(.A(pi677), .Y(new_n8166));
  nand_5 g05818(.A(new_n2557), .B(new_n8166), .Y(new_n8167));
  nand_5 g05819(.A(new_n2560), .B(pi677), .Y(new_n8168));
  nand_5 g05820(.A(new_n8168), .B(new_n8167), .Y(new_n8169));
  nand_5 g05821(.A(new_n8169), .B(new_n8165), .Y(new_n8170));
  not_8  g05822(.A(new_n8170), .Y(new_n8171));
  nor_5  g05823(.A(new_n8171), .B(new_n8134), .Y(new_n8172));
  nor_5  g05824(.A(new_n8169), .B(new_n8165), .Y(new_n8173));
  nand_5 g05825(.A(new_n8133), .B(new_n8163), .Y(new_n8174));
  nand_5 g05826(.A(new_n8167), .B(new_n8174), .Y(new_n8175));
  nor_5  g05827(.A(new_n8175), .B(new_n8173), .Y(new_n8176));
  nor_5  g05828(.A(new_n8176), .B(new_n8172), .Y(new_n8177));
  nand_5 g05829(.A(new_n8177), .B(new_n8162), .Y(new_n8178));
  xnor_4 g05830(.A(new_n8135), .B(new_n8131), .Y(new_n8179));
  xor_4  g05831(.A(new_n8177), .B(pi754), .Y(new_n8180));
  or_6   g05832(.A(new_n8180), .B(new_n8179), .Y(new_n8181));
  nand_5 g05833(.A(new_n8181), .B(new_n8178), .Y(new_n8182));
  nand_5 g05834(.A(new_n8182), .B(new_n8161), .Y(new_n8183));
  nand_5 g05835(.A(new_n8183), .B(new_n8160), .Y(new_n8184));
  nand_5 g05836(.A(new_n8184), .B(new_n8157), .Y(new_n8185));
  nand_5 g05837(.A(new_n8185), .B(new_n8156), .Y(new_n8186));
  nor_5  g05838(.A(new_n8186), .B(new_n8153), .Y(new_n8187));
  xor_4  g05839(.A(new_n8141), .B(new_n8124), .Y(new_n8188));
  xor_4  g05840(.A(new_n8186), .B(pi274), .Y(new_n8189));
  nor_5  g05841(.A(new_n8189), .B(new_n8188), .Y(new_n8190));
  or_6   g05842(.A(new_n8190), .B(new_n8187), .Y(new_n8191));
  or_6   g05843(.A(new_n8191), .B(pi031), .Y(new_n8192));
  xor_4  g05844(.A(new_n8143), .B(new_n8122), .Y(new_n8193));
  xor_4  g05845(.A(new_n8191), .B(pi031), .Y(new_n8194));
  nand_5 g05846(.A(new_n8194), .B(new_n8193), .Y(new_n8195));
  nand_5 g05847(.A(new_n8195), .B(new_n8192), .Y(new_n8196));
  nand_5 g05848(.A(new_n8196), .B(new_n8152), .Y(new_n8197));
  xor_4  g05849(.A(new_n8145), .B(new_n8120), .Y(new_n8198));
  not_8  g05850(.A(new_n8198), .Y(new_n8199));
  xor_4  g05851(.A(new_n8196), .B(pi310), .Y(new_n8200));
  or_6   g05852(.A(new_n8200), .B(new_n8199), .Y(new_n8201));
  nand_5 g05853(.A(new_n8201), .B(new_n8197), .Y(new_n8202));
  nand_5 g05854(.A(new_n8202), .B(new_n8151), .Y(new_n8203));
  not_8  g05855(.A(new_n8151), .Y(new_n8204));
  xor_4  g05856(.A(new_n8202), .B(new_n8204), .Y(new_n8205));
  or_6   g05857(.A(new_n8205), .B(pi586), .Y(new_n8206));
  nand_5 g05858(.A(new_n8206), .B(new_n8203), .Y(new_n8207));
  nand_5 g05859(.A(new_n8207), .B(new_n8150), .Y(new_n8208));
  not_8  g05860(.A(pi041), .Y(new_n8209));
  xor_4  g05861(.A(new_n8207), .B(new_n8150), .Y(new_n8210));
  nand_5 g05862(.A(new_n8210), .B(new_n8209), .Y(new_n8211));
  nand_5 g05863(.A(new_n8211), .B(new_n8208), .Y(new_n8212));
  or_6   g05864(.A(new_n8212), .B(new_n8114), .Y(new_n8213));
  nand_5 g05865(.A(new_n8213), .B(new_n8113), .Y(new_n8214));
  nand_5 g05866(.A(pi542), .B(new_n5546), .Y(new_n8215));
  nand_5 g05867(.A(new_n8149), .B(new_n8115), .Y(new_n8216));
  nand_5 g05868(.A(new_n8216), .B(new_n8215), .Y(new_n8217));
  not_8  g05869(.A(new_n8217), .Y(new_n8218));
  xnor_4 g05870(.A(new_n8212), .B(new_n8114), .Y(new_n8219));
  nor_5  g05871(.A(new_n8219), .B(new_n8218), .Y(new_n8220));
  nor_5  g05872(.A(new_n8108), .B(new_n8107), .Y(new_n8221));
  xor_4  g05873(.A(new_n8221), .B(pi810), .Y(new_n8222));
  xor_4  g05874(.A(new_n8200), .B(new_n8198), .Y(new_n8223));
  not_8  g05875(.A(new_n8103), .Y(new_n8224));
  xor_4  g05876(.A(new_n8224), .B(new_n8101), .Y(new_n8225));
  or_6   g05877(.A(new_n8225), .B(new_n8223), .Y(new_n8226));
  nand_5 g05878(.A(new_n8225), .B(new_n8223), .Y(new_n8227));
  xor_4  g05879(.A(new_n8096), .B(pi516), .Y(new_n8228));
  xor_4  g05880(.A(new_n8184), .B(new_n8157), .Y(new_n8229));
  xor_4  g05881(.A(new_n8087), .B(new_n8086), .Y(new_n8230));
  nand_5 g05882(.A(new_n8230), .B(new_n8229), .Y(new_n8231));
  not_8  g05883(.A(new_n8230), .Y(new_n8232));
  xor_4  g05884(.A(new_n8232), .B(new_n8229), .Y(new_n8233));
  xor_4  g05885(.A(new_n8182), .B(new_n8161), .Y(new_n8234));
  and_6  g05886(.A(new_n8076), .B(new_n8074), .Y(new_n8235));
  xor_4  g05887(.A(new_n8235), .B(pi515), .Y(new_n8236));
  not_8  g05888(.A(new_n8236), .Y(new_n8237));
  nor_5  g05889(.A(new_n2562), .B(new_n2554), .Y(new_n8238));
  nor_5  g05890(.A(new_n8173), .B(new_n8171), .Y(new_n8239));
  not_8  g05891(.A(new_n8239), .Y(new_n8240));
  nand_5 g05892(.A(new_n8240), .B(new_n8238), .Y(new_n8241));
  not_8  g05893(.A(new_n8241), .Y(new_n8242));
  xor_4  g05894(.A(new_n8069), .B(new_n8068), .Y(new_n8243));
  xor_4  g05895(.A(new_n8239), .B(new_n8238), .Y(new_n8244));
  nor_5  g05896(.A(new_n8244), .B(new_n8243), .Y(new_n8245));
  nor_5  g05897(.A(new_n8245), .B(new_n8242), .Y(new_n8246));
  nor_5  g05898(.A(new_n8246), .B(new_n8237), .Y(new_n8247));
  xor_4  g05899(.A(new_n8180), .B(new_n8179), .Y(new_n8248));
  xor_4  g05900(.A(new_n8246), .B(new_n8236), .Y(new_n8249));
  or_6   g05901(.A(new_n8249), .B(new_n8248), .Y(new_n8250));
  not_8  g05902(.A(new_n8250), .Y(new_n8251));
  nor_5  g05903(.A(new_n8251), .B(new_n8247), .Y(new_n8252));
  and_6  g05904(.A(new_n8252), .B(new_n8234), .Y(new_n8253));
  nor_5  g05905(.A(new_n8252), .B(new_n8234), .Y(new_n8254));
  xor_4  g05906(.A(new_n8082), .B(new_n8080), .Y(new_n8255));
  nor_5  g05907(.A(new_n8255), .B(new_n8254), .Y(new_n8256));
  nor_5  g05908(.A(new_n8256), .B(new_n8253), .Y(new_n8257));
  or_6   g05909(.A(new_n8257), .B(new_n8233), .Y(new_n8258));
  nand_5 g05910(.A(new_n8258), .B(new_n8231), .Y(new_n8259));
  nand_5 g05911(.A(new_n8092), .B(new_n8090), .Y(new_n8260));
  xor_4  g05912(.A(new_n8260), .B(pi764), .Y(new_n8261));
  or_6   g05913(.A(new_n8261), .B(new_n8259), .Y(new_n8262));
  xor_4  g05914(.A(new_n8189), .B(new_n8188), .Y(new_n8263));
  xor_4  g05915(.A(new_n8261), .B(new_n8259), .Y(new_n8264));
  nand_5 g05916(.A(new_n8264), .B(new_n8263), .Y(new_n8265));
  nand_5 g05917(.A(new_n8265), .B(new_n8262), .Y(new_n8266));
  nor_5  g05918(.A(new_n8266), .B(new_n8228), .Y(new_n8267));
  not_8  g05919(.A(new_n8228), .Y(new_n8268));
  xor_4  g05920(.A(new_n8266), .B(new_n8268), .Y(new_n8269));
  xnor_4 g05921(.A(new_n8194), .B(new_n8193), .Y(new_n8270));
  nor_5  g05922(.A(new_n8270), .B(new_n8269), .Y(new_n8271));
  or_6   g05923(.A(new_n8271), .B(new_n8267), .Y(new_n8272));
  nand_5 g05924(.A(new_n8272), .B(new_n8227), .Y(new_n8273));
  nand_5 g05925(.A(new_n8273), .B(new_n8226), .Y(new_n8274));
  not_8  g05926(.A(new_n8274), .Y(new_n8275));
  nor_5  g05927(.A(new_n8275), .B(new_n8222), .Y(new_n8276));
  not_8  g05928(.A(pi586), .Y(new_n8277));
  xor_4  g05929(.A(new_n8205), .B(new_n8277), .Y(new_n8278));
  xor_4  g05930(.A(new_n8274), .B(new_n8222), .Y(new_n8279));
  nor_5  g05931(.A(new_n8279), .B(new_n8278), .Y(new_n8280));
  or_6   g05932(.A(new_n8280), .B(new_n8276), .Y(new_n8281));
  xor_4  g05933(.A(new_n8110), .B(new_n8053), .Y(new_n8282));
  not_8  g05934(.A(new_n8282), .Y(new_n8283));
  nand_5 g05935(.A(new_n8283), .B(new_n8281), .Y(new_n8284));
  xor_4  g05936(.A(new_n8210), .B(pi041), .Y(new_n8285));
  xor_4  g05937(.A(new_n8282), .B(new_n8281), .Y(new_n8286));
  or_6   g05938(.A(new_n8286), .B(new_n8285), .Y(new_n8287));
  nand_5 g05939(.A(new_n8287), .B(new_n8284), .Y(new_n8288));
  xor_4  g05940(.A(new_n8219), .B(new_n8217), .Y(new_n8289));
  nor_5  g05941(.A(new_n8289), .B(new_n8288), .Y(new_n8290));
  or_6   g05942(.A(new_n8290), .B(new_n8220), .Y(new_n8291));
  xnor_4 g05943(.A(new_n8291), .B(new_n8214), .Y(po0037));
  xor_4  g05944(.A(new_n2532), .B(new_n2486), .Y(po0038));
  not_8  g05945(.A(pi109), .Y(new_n8294));
  xor_4  g05946(.A(pi466), .B(new_n8294), .Y(new_n8295));
  xor_4  g05947(.A(new_n8295), .B(pi009), .Y(new_n8296));
  not_8  g05948(.A(pi684), .Y(new_n8297));
  nand_5 g05949(.A(new_n8297), .B(pi553), .Y(new_n8298));
  xor_4  g05950(.A(pi684), .B(new_n4721), .Y(new_n8299));
  not_8  g05951(.A(pi742), .Y(new_n8300));
  nand_5 g05952(.A(pi757), .B(new_n8300), .Y(new_n8301));
  xor_4  g05953(.A(pi757), .B(new_n8300), .Y(new_n8302));
  nand_5 g05954(.A(pi655), .B(new_n4683), .Y(new_n8303));
  nand_5 g05955(.A(pi531), .B(new_n4679), .Y(new_n8304));
  nand_5 g05956(.A(new_n4534), .B(pi464), .Y(new_n8305));
  not_8  g05957(.A(new_n8305), .Y(new_n8306));
  xor_4  g05958(.A(pi660), .B(pi464), .Y(new_n8307));
  nand_5 g05959(.A(new_n3443), .B(pi178), .Y(new_n8308));
  nand_5 g05960(.A(pi330), .B(new_n4537), .Y(new_n8309));
  nand_5 g05961(.A(pi523), .B(new_n4540), .Y(new_n8310));
  nand_5 g05962(.A(new_n8310), .B(new_n8309), .Y(new_n8311));
  nand_5 g05963(.A(new_n8311), .B(new_n8308), .Y(new_n8312));
  nor_5  g05964(.A(new_n8312), .B(new_n8307), .Y(new_n8313));
  nor_5  g05965(.A(new_n8313), .B(new_n8306), .Y(new_n8314));
  xor_4  g05966(.A(pi531), .B(pi522), .Y(new_n8315));
  or_6   g05967(.A(new_n8315), .B(new_n8314), .Y(new_n8316));
  nand_5 g05968(.A(new_n8316), .B(new_n8304), .Y(new_n8317));
  xor_4  g05969(.A(pi655), .B(pi040), .Y(new_n8318));
  not_8  g05970(.A(new_n8318), .Y(new_n8319));
  nand_5 g05971(.A(new_n8319), .B(new_n8317), .Y(new_n8320));
  nand_5 g05972(.A(new_n8320), .B(new_n8303), .Y(new_n8321));
  nand_5 g05973(.A(new_n8321), .B(new_n8302), .Y(new_n8322));
  nand_5 g05974(.A(new_n8322), .B(new_n8301), .Y(new_n8323));
  nand_5 g05975(.A(new_n8323), .B(new_n8299), .Y(new_n8324));
  nand_5 g05976(.A(new_n8324), .B(new_n8298), .Y(new_n8325));
  nand_5 g05977(.A(new_n8325), .B(new_n8296), .Y(new_n8326));
  xor_4  g05978(.A(new_n8325), .B(new_n8296), .Y(new_n8327));
  not_8  g05979(.A(pi180), .Y(new_n8328));
  xnor_4 g05980(.A(new_n8323), .B(new_n8299), .Y(new_n8329));
  or_6   g05981(.A(new_n8329), .B(new_n8328), .Y(new_n8330));
  xor_4  g05982(.A(new_n8329), .B(new_n8328), .Y(new_n8331));
  not_8  g05983(.A(pi738), .Y(new_n8332));
  xnor_4 g05984(.A(new_n8321), .B(new_n8302), .Y(new_n8333));
  or_6   g05985(.A(new_n8333), .B(new_n8332), .Y(new_n8334));
  xor_4  g05986(.A(new_n8333), .B(new_n8332), .Y(new_n8335));
  not_8  g05987(.A(pi004), .Y(new_n8336));
  xor_4  g05988(.A(new_n8318), .B(new_n8317), .Y(new_n8337));
  nand_5 g05989(.A(new_n8337), .B(new_n8336), .Y(new_n8338));
  xor_4  g05990(.A(new_n8337), .B(new_n8336), .Y(new_n8339));
  xor_4  g05991(.A(new_n8315), .B(new_n8314), .Y(new_n8340));
  nor_5  g05992(.A(new_n8340), .B(pi747), .Y(new_n8341));
  xor_4  g05993(.A(new_n8340), .B(pi747), .Y(new_n8342));
  not_8  g05994(.A(new_n8342), .Y(new_n8343));
  xor_4  g05995(.A(new_n8312), .B(new_n8307), .Y(new_n8344));
  nand_5 g05996(.A(new_n8344), .B(pi078), .Y(new_n8345));
  xor_4  g05997(.A(new_n8344), .B(pi078), .Y(new_n8346));
  nand_5 g05998(.A(new_n8309), .B(new_n8308), .Y(new_n8347));
  xnor_4 g05999(.A(new_n8347), .B(new_n8310), .Y(new_n8348));
  or_6   g06000(.A(new_n8348), .B(new_n7016), .Y(new_n8349));
  xor_4  g06001(.A(new_n8348), .B(new_n7016), .Y(new_n8350));
  xor_4  g06002(.A(pi523), .B(new_n4540), .Y(new_n8351));
  nand_5 g06003(.A(new_n8351), .B(pi337), .Y(new_n8352));
  xor_4  g06004(.A(new_n8351), .B(new_n7019), .Y(new_n8353));
  nand_5 g06005(.A(new_n4543), .B(pi238), .Y(new_n8354));
  nand_5 g06006(.A(pi710), .B(new_n7054), .Y(new_n8355));
  nand_5 g06007(.A(new_n8355), .B(pi301), .Y(new_n8356));
  nand_5 g06008(.A(new_n8356), .B(new_n8354), .Y(new_n8357));
  not_8  g06009(.A(new_n8357), .Y(new_n8358));
  or_6   g06010(.A(new_n8358), .B(new_n8353), .Y(new_n8359));
  nand_5 g06011(.A(new_n8359), .B(new_n8352), .Y(new_n8360));
  nand_5 g06012(.A(new_n8360), .B(new_n8350), .Y(new_n8361));
  nand_5 g06013(.A(new_n8361), .B(new_n8349), .Y(new_n8362));
  nand_5 g06014(.A(new_n8362), .B(new_n8346), .Y(new_n8363));
  nand_5 g06015(.A(new_n8363), .B(new_n8345), .Y(new_n8364));
  nor_5  g06016(.A(new_n8364), .B(new_n8343), .Y(new_n8365));
  nor_5  g06017(.A(new_n8365), .B(new_n8341), .Y(new_n8366));
  not_8  g06018(.A(new_n8366), .Y(new_n8367));
  nand_5 g06019(.A(new_n8367), .B(new_n8339), .Y(new_n8368));
  and_6  g06020(.A(new_n8368), .B(new_n8338), .Y(new_n8369));
  nand_5 g06021(.A(new_n8369), .B(new_n8335), .Y(new_n8370));
  nand_5 g06022(.A(new_n8370), .B(new_n8334), .Y(new_n8371));
  nand_5 g06023(.A(new_n8371), .B(new_n8331), .Y(new_n8372));
  nand_5 g06024(.A(new_n8372), .B(new_n8330), .Y(new_n8373));
  nand_5 g06025(.A(new_n8373), .B(new_n8327), .Y(new_n8374));
  nand_5 g06026(.A(new_n8374), .B(new_n8326), .Y(new_n8375));
  nand_5 g06027(.A(pi466), .B(new_n8294), .Y(new_n8376));
  nand_5 g06028(.A(new_n8295), .B(pi009), .Y(new_n8377));
  nand_5 g06029(.A(new_n8377), .B(new_n8376), .Y(new_n8378));
  xor_4  g06030(.A(new_n8378), .B(pi118), .Y(new_n8379));
  not_8  g06031(.A(new_n8379), .Y(new_n8380));
  not_8  g06032(.A(pi034), .Y(new_n8381));
  nand_5 g06033(.A(pi689), .B(new_n8381), .Y(new_n8382));
  not_8  g06034(.A(pi689), .Y(new_n8383));
  nand_5 g06035(.A(new_n8383), .B(pi034), .Y(new_n8384));
  and_6  g06036(.A(new_n8384), .B(new_n8382), .Y(new_n8385));
  or_6   g06037(.A(new_n8385), .B(new_n8380), .Y(new_n8386));
  nand_5 g06038(.A(new_n8385), .B(new_n8380), .Y(new_n8387));
  nand_5 g06039(.A(new_n8387), .B(new_n8386), .Y(new_n8388));
  xor_4  g06040(.A(new_n8388), .B(new_n8375), .Y(new_n8389));
  or_6   g06041(.A(new_n8389), .B(new_n3706), .Y(new_n8390));
  xnor_4 g06042(.A(new_n8373), .B(new_n8327), .Y(new_n8391));
  nor_5  g06043(.A(new_n8391), .B(new_n3620), .Y(new_n8392));
  xor_4  g06044(.A(new_n8371), .B(new_n8331), .Y(new_n8393));
  nand_5 g06045(.A(new_n8393), .B(new_n3623), .Y(new_n8394));
  xnor_4 g06046(.A(new_n8393), .B(new_n3623), .Y(new_n8395));
  xor_4  g06047(.A(new_n8369), .B(new_n8335), .Y(new_n8396));
  or_6   g06048(.A(new_n8396), .B(new_n3675), .Y(new_n8397));
  xor_4  g06049(.A(new_n8396), .B(new_n3675), .Y(new_n8398));
  xor_4  g06050(.A(new_n8366), .B(new_n8339), .Y(new_n8399));
  or_6   g06051(.A(new_n8399), .B(new_n3669), .Y(new_n8400));
  xor_4  g06052(.A(new_n8399), .B(new_n3669), .Y(new_n8401));
  xor_4  g06053(.A(new_n8364), .B(new_n8342), .Y(new_n8402));
  not_8  g06054(.A(new_n8402), .Y(new_n8403));
  nor_5  g06055(.A(new_n8403), .B(new_n3624), .Y(new_n8404));
  xor_4  g06056(.A(new_n8402), .B(new_n3624), .Y(new_n8405));
  xnor_4 g06057(.A(new_n8362), .B(new_n8346), .Y(new_n8406));
  nor_5  g06058(.A(new_n8406), .B(new_n3659), .Y(new_n8407));
  xor_4  g06059(.A(new_n8406), .B(new_n3658), .Y(new_n8408));
  xor_4  g06060(.A(new_n8360), .B(new_n8350), .Y(new_n8409));
  not_8  g06061(.A(new_n8409), .Y(new_n8410));
  nor_5  g06062(.A(new_n8410), .B(new_n3648), .Y(new_n8411));
  xor_4  g06063(.A(new_n8409), .B(new_n3648), .Y(new_n8412));
  xor_4  g06064(.A(new_n8357), .B(new_n8353), .Y(new_n8413));
  nor_5  g06065(.A(new_n8413), .B(new_n3627), .Y(new_n8414));
  xor_4  g06066(.A(new_n8413), .B(new_n3628), .Y(new_n8415));
  nand_5 g06067(.A(new_n8354), .B(new_n8355), .Y(new_n8416));
  xor_4  g06068(.A(new_n8416), .B(new_n3638), .Y(new_n8417));
  or_6   g06069(.A(new_n8417), .B(new_n3642), .Y(new_n8418));
  nand_5 g06070(.A(new_n8417), .B(pi559), .Y(new_n8419));
  nand_5 g06071(.A(new_n8419), .B(new_n8418), .Y(new_n8420));
  nor_5  g06072(.A(new_n8420), .B(new_n8415), .Y(new_n8421));
  nor_5  g06073(.A(new_n8421), .B(new_n8414), .Y(new_n8422));
  nor_5  g06074(.A(new_n8422), .B(new_n8412), .Y(new_n8423));
  nor_5  g06075(.A(new_n8423), .B(new_n8411), .Y(new_n8424));
  nor_5  g06076(.A(new_n8424), .B(new_n8408), .Y(new_n8425));
  nor_5  g06077(.A(new_n8425), .B(new_n8407), .Y(new_n8426));
  nor_5  g06078(.A(new_n8426), .B(new_n8405), .Y(new_n8427));
  nor_5  g06079(.A(new_n8427), .B(new_n8404), .Y(new_n8428));
  nand_5 g06080(.A(new_n8428), .B(new_n8401), .Y(new_n8429));
  nand_5 g06081(.A(new_n8429), .B(new_n8400), .Y(new_n8430));
  nand_5 g06082(.A(new_n8430), .B(new_n8398), .Y(new_n8431));
  nand_5 g06083(.A(new_n8431), .B(new_n8397), .Y(new_n8432));
  or_6   g06084(.A(new_n8432), .B(new_n8395), .Y(new_n8433));
  nand_5 g06085(.A(new_n8433), .B(new_n8394), .Y(new_n8434));
  xor_4  g06086(.A(new_n8391), .B(new_n3620), .Y(new_n8435));
  and_6  g06087(.A(new_n8435), .B(new_n8434), .Y(new_n8436));
  nor_5  g06088(.A(new_n8436), .B(new_n8392), .Y(new_n8437));
  xor_4  g06089(.A(new_n8389), .B(new_n3706), .Y(new_n8438));
  nand_5 g06090(.A(new_n8438), .B(new_n8437), .Y(new_n8439));
  nand_5 g06091(.A(new_n8439), .B(new_n8390), .Y(new_n8440));
  not_8  g06092(.A(pi807), .Y(new_n8441));
  nor_5  g06093(.A(new_n3704), .B(new_n8441), .Y(new_n8442));
  nor_5  g06094(.A(new_n8442), .B(new_n3703), .Y(new_n8443));
  nand_5 g06095(.A(new_n3701), .B(new_n3696), .Y(new_n8444));
  nand_5 g06096(.A(new_n8444), .B(new_n3698), .Y(new_n8445));
  xor_4  g06097(.A(new_n8445), .B(new_n8443), .Y(new_n8446));
  not_8  g06098(.A(new_n8446), .Y(new_n8447));
  nand_5 g06099(.A(new_n8388), .B(new_n8375), .Y(new_n8448));
  nand_5 g06100(.A(new_n8378), .B(pi118), .Y(new_n8449));
  nand_5 g06101(.A(new_n8387), .B(new_n8384), .Y(new_n8450));
  and_6  g06102(.A(new_n8450), .B(new_n8449), .Y(new_n8451));
  nand_5 g06103(.A(new_n8451), .B(new_n8448), .Y(new_n8452));
  nand_5 g06104(.A(new_n8386), .B(new_n8449), .Y(new_n8453));
  and_6  g06105(.A(new_n8453), .B(new_n8384), .Y(new_n8454));
  and_6  g06106(.A(new_n8454), .B(new_n8375), .Y(new_n8455));
  nor_5  g06107(.A(new_n8382), .B(new_n8449), .Y(new_n8456));
  nor_5  g06108(.A(new_n8456), .B(new_n8455), .Y(new_n8457));
  nand_5 g06109(.A(new_n8457), .B(new_n8452), .Y(new_n8458));
  xor_4  g06110(.A(new_n8458), .B(new_n8447), .Y(new_n8459));
  xor_4  g06111(.A(new_n8459), .B(new_n8440), .Y(po0039));
  xor_4  g06112(.A(pi153), .B(new_n2373), .Y(new_n8461));
  nand_5 g06113(.A(new_n2386), .B(pi605), .Y(new_n8462));
  xor_4  g06114(.A(pi749), .B(new_n3779), .Y(new_n8463));
  nand_5 g06115(.A(new_n2389), .B(pi434), .Y(new_n8464));
  xor_4  g06116(.A(pi755), .B(new_n2357), .Y(new_n8465));
  nand_5 g06117(.A(pi552), .B(new_n2391), .Y(new_n8466));
  xor_4  g06118(.A(pi552), .B(new_n2391), .Y(new_n8467));
  nand_5 g06119(.A(new_n2429), .B(pi190), .Y(new_n8468));
  not_8  g06120(.A(new_n8468), .Y(new_n8469));
  nand_5 g06121(.A(new_n8469), .B(new_n8467), .Y(new_n8470));
  nand_5 g06122(.A(new_n8470), .B(new_n8466), .Y(new_n8471));
  nand_5 g06123(.A(new_n8471), .B(new_n8465), .Y(new_n8472));
  nand_5 g06124(.A(new_n8472), .B(new_n8464), .Y(new_n8473));
  nand_5 g06125(.A(new_n8473), .B(new_n8463), .Y(new_n8474));
  nand_5 g06126(.A(new_n8474), .B(new_n8462), .Y(new_n8475));
  xor_4  g06127(.A(new_n8475), .B(new_n8461), .Y(new_n8476));
  xnor_4 g06128(.A(new_n8476), .B(new_n5126), .Y(new_n8477));
  not_8  g06129(.A(new_n5147), .Y(new_n8478));
  xnor_4 g06130(.A(new_n8473), .B(new_n8463), .Y(new_n8479));
  nor_5  g06131(.A(new_n8479), .B(new_n8478), .Y(new_n8480));
  xor_4  g06132(.A(new_n8479), .B(new_n5147), .Y(new_n8481));
  xor_4  g06133(.A(new_n8471), .B(new_n8465), .Y(new_n8482));
  or_6   g06134(.A(new_n8482), .B(new_n5152), .Y(new_n8483));
  nand_5 g06135(.A(new_n8482), .B(new_n5152), .Y(new_n8484));
  not_8  g06136(.A(new_n8470), .Y(new_n8485));
  nand_5 g06137(.A(new_n8485), .B(new_n5159), .Y(new_n8486));
  nor_5  g06138(.A(new_n2429), .B(pi190), .Y(new_n8487));
  nand_5 g06139(.A(new_n8487), .B(new_n5161), .Y(new_n8488));
  nor_5  g06140(.A(new_n8488), .B(new_n8467), .Y(new_n8489));
  nand_5 g06141(.A(new_n8469), .B(new_n5157), .Y(new_n8490));
  nand_5 g06142(.A(new_n8490), .B(new_n8488), .Y(new_n8491));
  xor_4  g06143(.A(new_n8491), .B(new_n8467), .Y(new_n8492));
  nor_5  g06144(.A(new_n8492), .B(new_n5158), .Y(new_n8493));
  nor_5  g06145(.A(new_n8493), .B(new_n8489), .Y(new_n8494));
  nand_5 g06146(.A(new_n8494), .B(new_n8486), .Y(new_n8495));
  nand_5 g06147(.A(new_n8495), .B(new_n8484), .Y(new_n8496));
  nand_5 g06148(.A(new_n8496), .B(new_n8483), .Y(new_n8497));
  nor_5  g06149(.A(new_n8497), .B(new_n8481), .Y(new_n8498));
  nor_5  g06150(.A(new_n8498), .B(new_n8480), .Y(new_n8499));
  xnor_4 g06151(.A(new_n8499), .B(new_n8477), .Y(po0040));
  nor_5  g06152(.A(new_n6602), .B(new_n4204), .Y(new_n8501));
  xor_4  g06153(.A(new_n6602), .B(new_n4204), .Y(new_n8502));
  not_8  g06154(.A(new_n8502), .Y(new_n8503));
  xor_4  g06155(.A(new_n2553), .B(pi281), .Y(new_n8504));
  nor_5  g06156(.A(new_n8504), .B(new_n8503), .Y(new_n8505));
  or_6   g06157(.A(new_n8505), .B(new_n8501), .Y(new_n8506));
  xor_4  g06158(.A(new_n6605), .B(new_n6601), .Y(new_n8507));
  xor_4  g06159(.A(new_n8507), .B(new_n4139), .Y(new_n8508));
  not_8  g06160(.A(new_n8508), .Y(new_n8509));
  nand_5 g06161(.A(new_n8509), .B(new_n8506), .Y(new_n8510));
  not_8  g06162(.A(pi161), .Y(new_n8511));
  nor_5  g06163(.A(new_n8064), .B(new_n7343), .Y(new_n8512));
  xor_4  g06164(.A(new_n8512), .B(new_n8511), .Y(new_n8513));
  xor_4  g06165(.A(new_n8513), .B(new_n8069), .Y(new_n8514));
  xor_4  g06166(.A(new_n8508), .B(new_n8506), .Y(new_n8515));
  or_6   g06167(.A(new_n8515), .B(new_n8514), .Y(new_n8516));
  nand_5 g06168(.A(new_n8516), .B(new_n8510), .Y(new_n8517));
  nand_5 g06169(.A(new_n8512), .B(pi161), .Y(new_n8518));
  or_6   g06170(.A(new_n8513), .B(new_n8069), .Y(new_n8519));
  nand_5 g06171(.A(new_n8519), .B(new_n8518), .Y(new_n8520));
  xor_4  g06172(.A(new_n8072), .B(pi388), .Y(new_n8521));
  xor_4  g06173(.A(new_n8521), .B(new_n8520), .Y(new_n8522));
  or_6   g06174(.A(new_n8522), .B(new_n8517), .Y(new_n8523));
  nand_5 g06175(.A(new_n8522), .B(new_n8517), .Y(new_n8524));
  nand_5 g06176(.A(new_n8507), .B(pi215), .Y(new_n8525));
  not_8  g06177(.A(new_n8525), .Y(new_n8526));
  or_6   g06178(.A(new_n8526), .B(new_n6622), .Y(new_n8527));
  nand_5 g06179(.A(new_n8526), .B(new_n6622), .Y(new_n8528));
  nand_5 g06180(.A(new_n8528), .B(new_n8527), .Y(new_n8529));
  xor_4  g06181(.A(new_n8529), .B(pi460), .Y(new_n8530));
  nand_5 g06182(.A(new_n8530), .B(new_n8524), .Y(new_n8531));
  nand_5 g06183(.A(new_n8531), .B(new_n8523), .Y(new_n8532));
  nand_5 g06184(.A(new_n8072), .B(new_n6575), .Y(new_n8533));
  or_6   g06185(.A(new_n8521), .B(new_n8520), .Y(new_n8534));
  nand_5 g06186(.A(new_n8534), .B(new_n8533), .Y(new_n8535));
  xor_4  g06187(.A(new_n8081), .B(pi545), .Y(new_n8536));
  xor_4  g06188(.A(new_n8536), .B(new_n8535), .Y(new_n8537));
  xor_4  g06189(.A(new_n8537), .B(new_n8532), .Y(new_n8538));
  nand_5 g06190(.A(new_n8528), .B(new_n4133), .Y(new_n8539));
  nand_5 g06191(.A(new_n8539), .B(new_n8527), .Y(new_n8540));
  not_8  g06192(.A(new_n8540), .Y(new_n8541));
  or_6   g06193(.A(new_n8541), .B(new_n6640), .Y(new_n8542));
  nand_5 g06194(.A(new_n8541), .B(new_n6640), .Y(new_n8543));
  nand_5 g06195(.A(new_n8543), .B(new_n8542), .Y(new_n8544));
  xor_4  g06196(.A(new_n8544), .B(pi524), .Y(new_n8545));
  not_8  g06197(.A(new_n8545), .Y(new_n8546));
  xor_4  g06198(.A(new_n8546), .B(new_n8538), .Y(po0041));
  xor_4  g06199(.A(new_n5965), .B(new_n4879), .Y(new_n8548));
  or_6   g06200(.A(new_n5970), .B(pi676), .Y(new_n8549));
  xor_4  g06201(.A(new_n5970), .B(pi676), .Y(new_n8550));
  nor_5  g06202(.A(new_n5973), .B(pi634), .Y(new_n8551));
  nand_5 g06203(.A(new_n5978), .B(new_n4900), .Y(new_n8552));
  not_8  g06204(.A(new_n8552), .Y(new_n8553));
  not_8  g06205(.A(pi796), .Y(new_n8554));
  nor_5  g06206(.A(new_n5981), .B(new_n8554), .Y(new_n8555));
  xor_4  g06207(.A(new_n5981), .B(new_n8554), .Y(new_n8556));
  not_8  g06208(.A(new_n8556), .Y(new_n8557));
  nand_5 g06209(.A(new_n5984), .B(new_n4884), .Y(new_n8558));
  xor_4  g06210(.A(new_n5984), .B(new_n4884), .Y(new_n8559));
  not_8  g06211(.A(new_n8559), .Y(new_n8560));
  nand_5 g06212(.A(new_n5988), .B(pi130), .Y(new_n8561));
  nand_5 g06213(.A(new_n8561), .B(new_n5989), .Y(new_n8562));
  or_6   g06214(.A(new_n8562), .B(new_n8560), .Y(new_n8563));
  nand_5 g06215(.A(new_n8563), .B(new_n8558), .Y(new_n8564));
  nor_5  g06216(.A(new_n8564), .B(new_n8557), .Y(new_n8565));
  or_6   g06217(.A(new_n8565), .B(new_n8555), .Y(new_n8566));
  xor_4  g06218(.A(new_n5978), .B(pi232), .Y(new_n8567));
  nor_5  g06219(.A(new_n8567), .B(new_n8566), .Y(new_n8568));
  nor_5  g06220(.A(new_n8568), .B(new_n8553), .Y(new_n8569));
  xor_4  g06221(.A(new_n5973), .B(new_n4908), .Y(new_n8570));
  nor_5  g06222(.A(new_n8570), .B(new_n8569), .Y(new_n8571));
  or_6   g06223(.A(new_n8571), .B(new_n8551), .Y(new_n8572));
  nand_5 g06224(.A(new_n8572), .B(new_n8550), .Y(new_n8573));
  nand_5 g06225(.A(new_n8573), .B(new_n8549), .Y(new_n8574));
  xor_4  g06226(.A(new_n8574), .B(new_n8548), .Y(new_n8575));
  not_8  g06227(.A(pi228), .Y(new_n8576));
  nand_5 g06228(.A(new_n3016), .B(new_n5031), .Y(new_n8577));
  nand_5 g06229(.A(new_n3017), .B(pi617), .Y(new_n8578));
  nand_5 g06230(.A(new_n3018), .B(pi396), .Y(new_n8579));
  nand_5 g06231(.A(new_n8579), .B(new_n8578), .Y(new_n8580));
  nand_5 g06232(.A(new_n8580), .B(new_n8577), .Y(new_n8581));
  nand_5 g06233(.A(new_n8581), .B(new_n5021), .Y(new_n8582));
  xor_4  g06234(.A(new_n8581), .B(pi276), .Y(new_n8583));
  or_6   g06235(.A(new_n8583), .B(new_n3010), .Y(new_n8584));
  nand_5 g06236(.A(new_n8584), .B(new_n8582), .Y(new_n8585));
  or_6   g06237(.A(new_n8585), .B(new_n8576), .Y(new_n8586));
  xor_4  g06238(.A(new_n8585), .B(new_n8576), .Y(new_n8587));
  nand_5 g06239(.A(new_n8587), .B(new_n3008), .Y(new_n8588));
  nand_5 g06240(.A(new_n8588), .B(new_n8586), .Y(new_n8589));
  nand_5 g06241(.A(new_n8589), .B(pi557), .Y(new_n8590));
  not_8  g06242(.A(pi557), .Y(new_n8591));
  xor_4  g06243(.A(new_n8589), .B(new_n8591), .Y(new_n8592));
  or_6   g06244(.A(new_n8592), .B(new_n3034), .Y(new_n8593));
  nand_5 g06245(.A(new_n8593), .B(new_n8590), .Y(new_n8594));
  xor_4  g06246(.A(new_n8594), .B(new_n2993), .Y(new_n8595));
  xor_4  g06247(.A(new_n8595), .B(pi026), .Y(new_n8596));
  not_8  g06248(.A(new_n8596), .Y(new_n8597));
  xor_4  g06249(.A(new_n8570), .B(new_n8569), .Y(new_n8598));
  not_8  g06250(.A(new_n8598), .Y(new_n8599));
  xor_4  g06251(.A(new_n8567), .B(new_n8566), .Y(new_n8600));
  not_8  g06252(.A(new_n8600), .Y(new_n8601));
  xor_4  g06253(.A(new_n8587), .B(new_n3005), .Y(new_n8602));
  nand_5 g06254(.A(new_n8602), .B(new_n8601), .Y(new_n8603));
  xor_4  g06255(.A(new_n8564), .B(new_n8556), .Y(new_n8604));
  not_8  g06256(.A(new_n8604), .Y(new_n8605));
  xor_4  g06257(.A(new_n8583), .B(new_n3010), .Y(new_n8606));
  or_6   g06258(.A(new_n8606), .B(new_n8605), .Y(new_n8607));
  xor_4  g06259(.A(new_n8606), .B(new_n8605), .Y(new_n8608));
  xor_4  g06260(.A(pi220), .B(new_n4886), .Y(new_n8609));
  xor_4  g06261(.A(new_n8609), .B(pi385), .Y(new_n8610));
  nand_5 g06262(.A(new_n3019), .B(new_n5058), .Y(new_n8611));
  and_6  g06263(.A(new_n8611), .B(new_n8579), .Y(new_n8612));
  nor_5  g06264(.A(new_n8612), .B(new_n8610), .Y(new_n8613));
  nand_5 g06265(.A(new_n8577), .B(new_n8578), .Y(new_n8614));
  not_8  g06266(.A(new_n8610), .Y(new_n8615));
  nand_5 g06267(.A(new_n8611), .B(new_n8615), .Y(new_n8616));
  nand_5 g06268(.A(new_n8610), .B(new_n8579), .Y(new_n8617));
  nand_5 g06269(.A(new_n8617), .B(new_n8616), .Y(new_n8618));
  xor_4  g06270(.A(new_n8618), .B(new_n8614), .Y(new_n8619));
  and_6  g06271(.A(new_n8619), .B(new_n8613), .Y(new_n8620));
  xor_4  g06272(.A(new_n8562), .B(new_n8560), .Y(new_n8621));
  nor_5  g06273(.A(new_n8621), .B(new_n8619), .Y(new_n8622));
  nor_5  g06274(.A(new_n8622), .B(new_n8620), .Y(new_n8623));
  nand_5 g06275(.A(new_n8623), .B(new_n8608), .Y(new_n8624));
  nand_5 g06276(.A(new_n8624), .B(new_n8607), .Y(new_n8625));
  xor_4  g06277(.A(new_n8602), .B(new_n8600), .Y(new_n8626));
  or_6   g06278(.A(new_n8626), .B(new_n8625), .Y(new_n8627));
  nand_5 g06279(.A(new_n8627), .B(new_n8603), .Y(new_n8628));
  nand_5 g06280(.A(new_n8628), .B(new_n8599), .Y(new_n8629));
  xor_4  g06281(.A(new_n8628), .B(new_n8598), .Y(new_n8630));
  xor_4  g06282(.A(new_n8592), .B(new_n3034), .Y(new_n8631));
  or_6   g06283(.A(new_n8631), .B(new_n8630), .Y(new_n8632));
  nand_5 g06284(.A(new_n8632), .B(new_n8629), .Y(new_n8633));
  nor_5  g06285(.A(new_n8633), .B(new_n8597), .Y(new_n8634));
  xor_4  g06286(.A(new_n8572), .B(new_n8550), .Y(new_n8635));
  not_8  g06287(.A(new_n8635), .Y(new_n8636));
  xor_4  g06288(.A(new_n8633), .B(new_n8596), .Y(new_n8637));
  nor_5  g06289(.A(new_n8637), .B(new_n8636), .Y(new_n8638));
  or_6   g06290(.A(new_n8638), .B(new_n8634), .Y(new_n8639));
  xor_4  g06291(.A(new_n8639), .B(new_n8575), .Y(new_n8640));
  not_8  g06292(.A(pi768), .Y(new_n8641));
  xor_4  g06293(.A(new_n2987), .B(new_n8641), .Y(new_n8642));
  nand_5 g06294(.A(new_n8594), .B(new_n2993), .Y(new_n8643));
  nand_5 g06295(.A(new_n8595), .B(pi026), .Y(new_n8644));
  nand_5 g06296(.A(new_n8644), .B(new_n8643), .Y(new_n8645));
  xor_4  g06297(.A(new_n8645), .B(new_n8642), .Y(new_n8646));
  xor_4  g06298(.A(new_n8646), .B(new_n8640), .Y(po0042));
  not_8  g06299(.A(new_n6667), .Y(new_n8648));
  xor_4  g06300(.A(pi563), .B(new_n6723), .Y(new_n8649));
  nand_5 g06301(.A(new_n3234), .B(pi264), .Y(new_n8650));
  xor_4  g06302(.A(pi457), .B(new_n6726), .Y(new_n8651));
  nand_5 g06303(.A(new_n3238), .B(pi333), .Y(new_n8652));
  xor_4  g06304(.A(pi633), .B(new_n6732), .Y(new_n8653));
  nand_5 g06305(.A(new_n3340), .B(pi569), .Y(new_n8654));
  not_8  g06306(.A(new_n8654), .Y(new_n8655));
  nand_5 g06307(.A(new_n8655), .B(new_n8653), .Y(new_n8656));
  nand_5 g06308(.A(new_n8656), .B(new_n8652), .Y(new_n8657));
  nand_5 g06309(.A(new_n8657), .B(new_n8651), .Y(new_n8658));
  nand_5 g06310(.A(new_n8658), .B(new_n8650), .Y(new_n8659));
  xor_4  g06311(.A(new_n8659), .B(new_n8649), .Y(new_n8660));
  not_8  g06312(.A(new_n8660), .Y(new_n8661));
  nand_5 g06313(.A(new_n8661), .B(pi779), .Y(new_n8662));
  xnor_4 g06314(.A(new_n8657), .B(new_n8651), .Y(new_n8663));
  nand_5 g06315(.A(new_n8663), .B(pi760), .Y(new_n8664));
  or_6   g06316(.A(new_n8663), .B(new_n6809), .Y(new_n8665));
  nand_5 g06317(.A(new_n8663), .B(new_n6809), .Y(new_n8666));
  nand_5 g06318(.A(new_n8666), .B(new_n8665), .Y(new_n8667));
  xor_4  g06319(.A(new_n8653), .B(new_n4075), .Y(new_n8668));
  nand_5 g06320(.A(pi718), .B(new_n6766), .Y(new_n8669));
  nand_5 g06321(.A(new_n8669), .B(pi708), .Y(new_n8670));
  not_8  g06322(.A(pi708), .Y(new_n8671));
  nand_5 g06323(.A(new_n8654), .B(new_n8671), .Y(new_n8672));
  nand_5 g06324(.A(new_n8672), .B(new_n8670), .Y(new_n8673));
  xor_4  g06325(.A(new_n8673), .B(new_n8668), .Y(new_n8674));
  nor_5  g06326(.A(new_n8655), .B(new_n8653), .Y(new_n8675));
  nand_5 g06327(.A(new_n8675), .B(new_n8674), .Y(new_n8676));
  nand_5 g06328(.A(pi837), .B(pi708), .Y(new_n8677));
  nand_5 g06329(.A(new_n8669), .B(new_n8654), .Y(new_n8678));
  not_8  g06330(.A(new_n8678), .Y(new_n8679));
  nor_5  g06331(.A(new_n8679), .B(new_n8677), .Y(new_n8680));
  not_8  g06332(.A(new_n8656), .Y(new_n8681));
  nand_5 g06333(.A(new_n4075), .B(new_n8671), .Y(new_n8682));
  and_6  g06334(.A(new_n8682), .B(new_n8681), .Y(new_n8683));
  nor_5  g06335(.A(new_n8683), .B(new_n8680), .Y(new_n8684));
  nand_5 g06336(.A(new_n8684), .B(new_n8676), .Y(new_n8685));
  nand_5 g06337(.A(new_n8685), .B(new_n8667), .Y(new_n8686));
  nand_5 g06338(.A(new_n8686), .B(new_n8664), .Y(new_n8687));
  xor_4  g06339(.A(new_n8660), .B(pi779), .Y(new_n8688));
  not_8  g06340(.A(new_n8688), .Y(new_n8689));
  nand_5 g06341(.A(new_n8689), .B(new_n8687), .Y(new_n8690));
  nand_5 g06342(.A(new_n8690), .B(new_n8662), .Y(new_n8691));
  xor_4  g06343(.A(pi649), .B(new_n6719), .Y(new_n8692));
  nand_5 g06344(.A(new_n3231), .B(pi483), .Y(new_n8693));
  nand_5 g06345(.A(new_n8659), .B(new_n8649), .Y(new_n8694));
  nand_5 g06346(.A(new_n8694), .B(new_n8693), .Y(new_n8695));
  xor_4  g06347(.A(new_n8695), .B(new_n8692), .Y(new_n8696));
  xor_4  g06348(.A(new_n8696), .B(pi587), .Y(new_n8697));
  not_8  g06349(.A(new_n8697), .Y(new_n8698));
  xor_4  g06350(.A(new_n8698), .B(new_n8691), .Y(new_n8699));
  xor_4  g06351(.A(new_n8688), .B(new_n8687), .Y(new_n8700));
  nand_5 g06352(.A(new_n8700), .B(new_n6668), .Y(new_n8701));
  xor_4  g06353(.A(new_n8700), .B(new_n6684), .Y(new_n8702));
  xor_4  g06354(.A(new_n8678), .B(new_n8671), .Y(new_n8703));
  nor_5  g06355(.A(new_n8703), .B(new_n6669), .Y(new_n8704));
  not_8  g06356(.A(new_n8704), .Y(new_n8705));
  nand_5 g06357(.A(new_n8705), .B(new_n8674), .Y(new_n8706));
  xor_4  g06358(.A(new_n8704), .B(new_n8674), .Y(new_n8707));
  or_6   g06359(.A(new_n8707), .B(new_n6672), .Y(new_n8708));
  nand_5 g06360(.A(new_n8708), .B(new_n8706), .Y(new_n8709));
  and_6  g06361(.A(new_n8709), .B(new_n6678), .Y(new_n8710));
  nor_5  g06362(.A(new_n8709), .B(new_n6678), .Y(new_n8711));
  xor_4  g06363(.A(new_n8685), .B(new_n8667), .Y(new_n8712));
  nor_5  g06364(.A(new_n8712), .B(new_n8711), .Y(new_n8713));
  nor_5  g06365(.A(new_n8713), .B(new_n8710), .Y(new_n8714));
  or_6   g06366(.A(new_n8714), .B(new_n8702), .Y(new_n8715));
  nand_5 g06367(.A(new_n8715), .B(new_n8701), .Y(new_n8716));
  xor_4  g06368(.A(new_n8716), .B(new_n8699), .Y(new_n8717));
  xor_4  g06369(.A(new_n8717), .B(new_n8648), .Y(po0043));
  nand_5 g06370(.A(pi551), .B(new_n6787), .Y(new_n8719));
  xor_4  g06371(.A(pi551), .B(new_n6787), .Y(new_n8720));
  nand_5 g06372(.A(pi420), .B(new_n6714), .Y(new_n8721));
  xor_4  g06373(.A(pi420), .B(new_n6714), .Y(new_n8722));
  nand_5 g06374(.A(new_n6716), .B(pi115), .Y(new_n8723));
  not_8  g06375(.A(pi115), .Y(new_n8724));
  xor_4  g06376(.A(pi615), .B(new_n8724), .Y(new_n8725));
  nand_5 g06377(.A(new_n6719), .B(pi173), .Y(new_n8726));
  not_8  g06378(.A(pi173), .Y(new_n8727));
  xor_4  g06379(.A(pi579), .B(new_n8727), .Y(new_n8728));
  nand_5 g06380(.A(pi535), .B(new_n6723), .Y(new_n8729));
  xor_4  g06381(.A(pi535), .B(new_n6723), .Y(new_n8730));
  nand_5 g06382(.A(pi719), .B(new_n6726), .Y(new_n8731));
  xor_4  g06383(.A(pi719), .B(new_n6726), .Y(new_n8732));
  nand_5 g06384(.A(new_n6732), .B(pi024), .Y(new_n8733));
  nand_5 g06385(.A(pi580), .B(new_n6766), .Y(new_n8734));
  not_8  g06386(.A(new_n8734), .Y(new_n8735));
  xor_4  g06387(.A(pi333), .B(new_n2638), .Y(new_n8736));
  nand_5 g06388(.A(new_n8736), .B(new_n8735), .Y(new_n8737));
  nand_5 g06389(.A(new_n8737), .B(new_n8733), .Y(new_n8738));
  nand_5 g06390(.A(new_n8738), .B(new_n8732), .Y(new_n8739));
  nand_5 g06391(.A(new_n8739), .B(new_n8731), .Y(new_n8740));
  nand_5 g06392(.A(new_n8740), .B(new_n8730), .Y(new_n8741));
  nand_5 g06393(.A(new_n8741), .B(new_n8729), .Y(new_n8742));
  nand_5 g06394(.A(new_n8742), .B(new_n8728), .Y(new_n8743));
  nand_5 g06395(.A(new_n8743), .B(new_n8726), .Y(new_n8744));
  nand_5 g06396(.A(new_n8744), .B(new_n8725), .Y(new_n8745));
  nand_5 g06397(.A(new_n8745), .B(new_n8723), .Y(new_n8746));
  nand_5 g06398(.A(new_n8746), .B(new_n8722), .Y(new_n8747));
  nand_5 g06399(.A(new_n8747), .B(new_n8721), .Y(new_n8748));
  nand_5 g06400(.A(new_n8748), .B(new_n8720), .Y(new_n8749));
  nand_5 g06401(.A(new_n8749), .B(new_n8719), .Y(new_n8750));
  not_8  g06402(.A(pi592), .Y(new_n8751));
  nand_5 g06403(.A(pi728), .B(new_n8751), .Y(new_n8752));
  nand_5 g06404(.A(new_n7592), .B(pi592), .Y(new_n8753));
  and_6  g06405(.A(new_n8753), .B(new_n8752), .Y(new_n8754));
  xor_4  g06406(.A(new_n8754), .B(new_n8750), .Y(new_n8755));
  not_8  g06407(.A(new_n8755), .Y(new_n8756));
  nand_5 g06408(.A(new_n8055), .B(pi123), .Y(new_n8757));
  not_8  g06409(.A(new_n8757), .Y(new_n8758));
  not_8  g06410(.A(pi123), .Y(new_n8759));
  xor_4  g06411(.A(pi258), .B(new_n8759), .Y(new_n8760));
  not_8  g06412(.A(new_n8760), .Y(new_n8761));
  not_8  g06413(.A(pi516), .Y(new_n8762));
  nand_5 g06414(.A(pi811), .B(new_n8762), .Y(new_n8763));
  not_8  g06415(.A(new_n8763), .Y(new_n8764));
  xor_4  g06416(.A(pi811), .B(new_n8762), .Y(new_n8765));
  not_8  g06417(.A(new_n8765), .Y(new_n8766));
  not_8  g06418(.A(pi804), .Y(new_n8767));
  nand_5 g06419(.A(new_n8767), .B(pi764), .Y(new_n8768));
  xor_4  g06420(.A(pi804), .B(new_n8091), .Y(new_n8769));
  not_8  g06421(.A(pi573), .Y(new_n8770));
  nand_5 g06422(.A(new_n8770), .B(pi075), .Y(new_n8771));
  nand_5 g06423(.A(pi573), .B(new_n8086), .Y(new_n8772));
  not_8  g06424(.A(pi273), .Y(new_n8773));
  nand_5 g06425(.A(pi698), .B(new_n8773), .Y(new_n8774));
  nand_5 g06426(.A(pi576), .B(new_n8075), .Y(new_n8775));
  xor_4  g06427(.A(pi576), .B(new_n8075), .Y(new_n8776));
  nand_5 g06428(.A(new_n8063), .B(pi401), .Y(new_n8777));
  not_8  g06429(.A(pi401), .Y(new_n8778));
  nand_5 g06430(.A(pi474), .B(new_n8778), .Y(new_n8779));
  nand_5 g06431(.A(new_n8779), .B(pi435), .Y(new_n8780));
  nand_5 g06432(.A(new_n8780), .B(new_n8777), .Y(new_n8781));
  nand_5 g06433(.A(new_n8781), .B(new_n8776), .Y(new_n8782));
  nand_5 g06434(.A(new_n8782), .B(new_n8775), .Y(new_n8783));
  xor_4  g06435(.A(pi698), .B(new_n8773), .Y(new_n8784));
  not_8  g06436(.A(new_n8784), .Y(new_n8785));
  or_6   g06437(.A(new_n8785), .B(new_n8783), .Y(new_n8786));
  nand_5 g06438(.A(new_n8786), .B(new_n8774), .Y(new_n8787));
  nand_5 g06439(.A(new_n8787), .B(new_n8772), .Y(new_n8788));
  nand_5 g06440(.A(new_n8788), .B(new_n8771), .Y(new_n8789));
  nand_5 g06441(.A(new_n8789), .B(new_n8769), .Y(new_n8790));
  nand_5 g06442(.A(new_n8790), .B(new_n8768), .Y(new_n8791));
  nor_5  g06443(.A(new_n8791), .B(new_n8766), .Y(new_n8792));
  nor_5  g06444(.A(new_n8792), .B(new_n8764), .Y(new_n8793));
  nor_5  g06445(.A(new_n8793), .B(new_n8761), .Y(new_n8794));
  nor_5  g06446(.A(new_n8794), .B(new_n8758), .Y(new_n8795));
  not_8  g06447(.A(pi469), .Y(new_n8796));
  nand_5 g06448(.A(pi810), .B(new_n8796), .Y(new_n8797));
  not_8  g06449(.A(pi810), .Y(new_n8798));
  nand_5 g06450(.A(new_n8798), .B(pi469), .Y(new_n8799));
  nand_5 g06451(.A(new_n8799), .B(new_n8797), .Y(new_n8800));
  xor_4  g06452(.A(new_n8800), .B(new_n8795), .Y(new_n8801));
  xor_4  g06453(.A(new_n8801), .B(new_n8756), .Y(new_n8802));
  not_8  g06454(.A(new_n8802), .Y(new_n8803));
  xor_4  g06455(.A(new_n8748), .B(new_n8720), .Y(new_n8804));
  xor_4  g06456(.A(new_n8793), .B(new_n8760), .Y(new_n8805));
  or_6   g06457(.A(new_n8805), .B(new_n8804), .Y(new_n8806));
  xor_4  g06458(.A(new_n8805), .B(new_n8804), .Y(new_n8807));
  xor_4  g06459(.A(new_n8746), .B(new_n8722), .Y(new_n8808));
  xor_4  g06460(.A(new_n8791), .B(new_n8765), .Y(new_n8809));
  or_6   g06461(.A(new_n8809), .B(new_n8808), .Y(new_n8810));
  xor_4  g06462(.A(new_n8809), .B(new_n8808), .Y(new_n8811));
  xor_4  g06463(.A(new_n8744), .B(new_n8725), .Y(new_n8812));
  xor_4  g06464(.A(new_n8789), .B(new_n8769), .Y(new_n8813));
  nor_5  g06465(.A(new_n8813), .B(new_n8812), .Y(new_n8814));
  xor_4  g06466(.A(new_n8742), .B(new_n8728), .Y(new_n8815));
  nand_5 g06467(.A(new_n8772), .B(new_n8771), .Y(new_n8816));
  xnor_4 g06468(.A(new_n8816), .B(new_n8787), .Y(new_n8817));
  or_6   g06469(.A(new_n8817), .B(new_n8815), .Y(new_n8818));
  xor_4  g06470(.A(new_n8817), .B(new_n8815), .Y(new_n8819));
  xor_4  g06471(.A(new_n8740), .B(new_n8730), .Y(new_n8820));
  xor_4  g06472(.A(new_n8785), .B(new_n8783), .Y(new_n8821));
  nor_5  g06473(.A(new_n8821), .B(new_n8820), .Y(new_n8822));
  xor_4  g06474(.A(new_n8821), .B(new_n8820), .Y(new_n8823));
  not_8  g06475(.A(new_n8823), .Y(new_n8824));
  xor_4  g06476(.A(new_n8738), .B(new_n8732), .Y(new_n8825));
  xnor_4 g06477(.A(new_n8781), .B(new_n8776), .Y(new_n8826));
  nand_5 g06478(.A(new_n8826), .B(new_n8825), .Y(new_n8827));
  or_6   g06479(.A(new_n8826), .B(new_n8825), .Y(new_n8828));
  nand_5 g06480(.A(new_n7250), .B(pi149), .Y(new_n8829));
  not_8  g06481(.A(new_n8829), .Y(new_n8830));
  nand_5 g06482(.A(new_n8830), .B(new_n8736), .Y(new_n8831));
  nand_5 g06483(.A(new_n8777), .B(new_n8779), .Y(new_n8832));
  xor_4  g06484(.A(new_n8736), .B(new_n8735), .Y(new_n8833));
  not_8  g06485(.A(new_n8833), .Y(new_n8834));
  not_8  g06486(.A(pi435), .Y(new_n8835));
  nor_5  g06487(.A(new_n7250), .B(pi149), .Y(new_n8836));
  nor_5  g06488(.A(new_n8836), .B(new_n8835), .Y(new_n8837));
  nor_5  g06489(.A(new_n8830), .B(pi435), .Y(new_n8838));
  or_6   g06490(.A(new_n8838), .B(new_n8837), .Y(new_n8839));
  xor_4  g06491(.A(new_n8839), .B(new_n8832), .Y(new_n8840));
  xor_4  g06492(.A(new_n8840), .B(new_n8834), .Y(new_n8841));
  nand_5 g06493(.A(new_n8841), .B(new_n8832), .Y(new_n8842));
  nor_5  g06494(.A(new_n8832), .B(pi435), .Y(new_n8843));
  nand_5 g06495(.A(new_n8834), .B(new_n8829), .Y(new_n8844));
  nor_5  g06496(.A(new_n8844), .B(new_n8837), .Y(new_n8845));
  nor_5  g06497(.A(new_n8845), .B(new_n8843), .Y(new_n8846));
  nand_5 g06498(.A(new_n8846), .B(new_n8842), .Y(new_n8847));
  nand_5 g06499(.A(new_n8847), .B(new_n8831), .Y(new_n8848));
  nand_5 g06500(.A(new_n8848), .B(new_n8828), .Y(new_n8849));
  nand_5 g06501(.A(new_n8849), .B(new_n8827), .Y(new_n8850));
  nor_5  g06502(.A(new_n8850), .B(new_n8824), .Y(new_n8851));
  or_6   g06503(.A(new_n8851), .B(new_n8822), .Y(new_n8852));
  nand_5 g06504(.A(new_n8852), .B(new_n8819), .Y(new_n8853));
  nand_5 g06505(.A(new_n8853), .B(new_n8818), .Y(new_n8854));
  not_8  g06506(.A(new_n8854), .Y(new_n8855));
  xnor_4 g06507(.A(new_n8813), .B(new_n8812), .Y(new_n8856));
  nor_5  g06508(.A(new_n8856), .B(new_n8855), .Y(new_n8857));
  or_6   g06509(.A(new_n8857), .B(new_n8814), .Y(new_n8858));
  nand_5 g06510(.A(new_n8858), .B(new_n8811), .Y(new_n8859));
  nand_5 g06511(.A(new_n8859), .B(new_n8810), .Y(new_n8860));
  nand_5 g06512(.A(new_n8860), .B(new_n8807), .Y(new_n8861));
  nand_5 g06513(.A(new_n8861), .B(new_n8806), .Y(new_n8862));
  xor_4  g06514(.A(new_n8862), .B(new_n8803), .Y(new_n8863));
  not_8  g06515(.A(new_n8863), .Y(new_n8864));
  not_8  g06516(.A(pi205), .Y(new_n8865));
  nand_5 g06517(.A(pi437), .B(new_n8865), .Y(new_n8866));
  xor_4  g06518(.A(pi437), .B(new_n8865), .Y(new_n8867));
  not_8  g06519(.A(pi578), .Y(new_n8868));
  nand_5 g06520(.A(new_n8868), .B(pi033), .Y(new_n8869));
  xor_4  g06521(.A(pi578), .B(new_n6799), .Y(new_n8870));
  nand_5 g06522(.A(new_n6201), .B(pi572), .Y(new_n8871));
  nand_5 g06523(.A(new_n6165), .B(pi587), .Y(new_n8872));
  not_8  g06524(.A(pi587), .Y(new_n8873));
  xor_4  g06525(.A(pi644), .B(new_n8873), .Y(new_n8874));
  not_8  g06526(.A(pi147), .Y(new_n8875));
  nand_5 g06527(.A(pi779), .B(new_n8875), .Y(new_n8876));
  not_8  g06528(.A(new_n8876), .Y(new_n8877));
  xor_4  g06529(.A(pi779), .B(new_n8875), .Y(new_n8878));
  not_8  g06530(.A(new_n8878), .Y(new_n8879));
  nor_5  g06531(.A(new_n6809), .B(pi609), .Y(new_n8880));
  xor_4  g06532(.A(pi760), .B(pi609), .Y(new_n8881));
  nand_5 g06533(.A(new_n8677), .B(pi356), .Y(new_n8882));
  nand_5 g06534(.A(new_n8882), .B(new_n8682), .Y(new_n8883));
  nor_5  g06535(.A(new_n8883), .B(new_n8881), .Y(new_n8884));
  nor_5  g06536(.A(new_n8884), .B(new_n8880), .Y(new_n8885));
  nor_5  g06537(.A(new_n8885), .B(new_n8879), .Y(new_n8886));
  nor_5  g06538(.A(new_n8886), .B(new_n8877), .Y(new_n8887));
  not_8  g06539(.A(new_n8887), .Y(new_n8888));
  nand_5 g06540(.A(new_n8888), .B(new_n8874), .Y(new_n8889));
  nand_5 g06541(.A(new_n8889), .B(new_n8872), .Y(new_n8890));
  xor_4  g06542(.A(pi726), .B(pi572), .Y(new_n8891));
  not_8  g06543(.A(new_n8891), .Y(new_n8892));
  nand_5 g06544(.A(new_n8892), .B(new_n8890), .Y(new_n8893));
  nand_5 g06545(.A(new_n8893), .B(new_n8871), .Y(new_n8894));
  nand_5 g06546(.A(new_n8894), .B(new_n8870), .Y(new_n8895));
  nand_5 g06547(.A(new_n8895), .B(new_n8869), .Y(new_n8896));
  nand_5 g06548(.A(new_n8896), .B(new_n8867), .Y(new_n8897));
  nand_5 g06549(.A(new_n8897), .B(new_n8866), .Y(new_n8898));
  xor_4  g06550(.A(pi666), .B(new_n6307), .Y(new_n8899));
  xor_4  g06551(.A(new_n8899), .B(new_n8898), .Y(new_n8900));
  nor_5  g06552(.A(new_n8900), .B(new_n8864), .Y(new_n8901));
  xor_4  g06553(.A(new_n8896), .B(new_n8867), .Y(new_n8902));
  xor_4  g06554(.A(new_n8860), .B(new_n8807), .Y(new_n8903));
  nor_5  g06555(.A(new_n8903), .B(new_n8902), .Y(new_n8904));
  xor_4  g06556(.A(new_n8858), .B(new_n8811), .Y(new_n8905));
  not_8  g06557(.A(new_n8905), .Y(new_n8906));
  xnor_4 g06558(.A(new_n8894), .B(new_n8870), .Y(new_n8907));
  nor_5  g06559(.A(new_n8907), .B(new_n8906), .Y(new_n8908));
  xor_4  g06560(.A(new_n8892), .B(new_n8890), .Y(new_n8909));
  xor_4  g06561(.A(new_n8856), .B(new_n8854), .Y(new_n8910));
  not_8  g06562(.A(new_n8910), .Y(new_n8911));
  nor_5  g06563(.A(new_n8911), .B(new_n8909), .Y(new_n8912));
  xnor_4 g06564(.A(new_n8852), .B(new_n8819), .Y(new_n8913));
  xor_4  g06565(.A(new_n8887), .B(new_n8874), .Y(new_n8914));
  or_6   g06566(.A(new_n8914), .B(new_n8913), .Y(new_n8915));
  xor_4  g06567(.A(new_n8885), .B(new_n8878), .Y(new_n8916));
  xor_4  g06568(.A(new_n8850), .B(new_n8823), .Y(new_n8917));
  or_6   g06569(.A(new_n8917), .B(new_n8916), .Y(new_n8918));
  xor_4  g06570(.A(new_n8917), .B(new_n8916), .Y(new_n8919));
  xor_4  g06571(.A(new_n8883), .B(new_n8881), .Y(new_n8920));
  nand_5 g06572(.A(new_n8828), .B(new_n8827), .Y(new_n8921));
  xor_4  g06573(.A(new_n8921), .B(new_n8848), .Y(new_n8922));
  nor_5  g06574(.A(new_n8922), .B(new_n8920), .Y(new_n8923));
  xnor_4 g06575(.A(new_n8922), .B(new_n8920), .Y(new_n8924));
  xor_4  g06576(.A(pi837), .B(new_n4086), .Y(new_n8925));
  xor_4  g06577(.A(new_n8925), .B(new_n8841), .Y(new_n8926));
  nor_5  g06578(.A(new_n8836), .B(new_n8830), .Y(new_n8927));
  xor_4  g06579(.A(new_n8927), .B(pi435), .Y(new_n8928));
  nor_5  g06580(.A(pi708), .B(new_n4088), .Y(new_n8929));
  nand_5 g06581(.A(new_n8929), .B(new_n8928), .Y(new_n8930));
  nand_5 g06582(.A(pi708), .B(new_n4088), .Y(new_n8931));
  nor_5  g06583(.A(new_n8931), .B(new_n8928), .Y(new_n8932));
  not_8  g06584(.A(new_n8932), .Y(new_n8933));
  nand_5 g06585(.A(new_n8933), .B(new_n8930), .Y(new_n8934));
  xor_4  g06586(.A(new_n8934), .B(new_n8926), .Y(po1281));
  nand_5 g06587(.A(po1281), .B(new_n8841), .Y(new_n8936));
  nor_5  g06588(.A(new_n8930), .B(new_n8925), .Y(new_n8937));
  nor_5  g06589(.A(new_n8925), .B(new_n8841), .Y(new_n8938));
  nand_5 g06590(.A(new_n8933), .B(pi708), .Y(new_n8939));
  nor_5  g06591(.A(new_n8939), .B(new_n8938), .Y(new_n8940));
  nor_5  g06592(.A(new_n8940), .B(new_n8937), .Y(new_n8941));
  and_6  g06593(.A(new_n8941), .B(new_n8936), .Y(new_n8942));
  nor_5  g06594(.A(new_n8942), .B(new_n8924), .Y(new_n8943));
  or_6   g06595(.A(new_n8943), .B(new_n8923), .Y(new_n8944));
  not_8  g06596(.A(new_n8944), .Y(new_n8945));
  nand_5 g06597(.A(new_n8945), .B(new_n8919), .Y(new_n8946));
  nand_5 g06598(.A(new_n8946), .B(new_n8918), .Y(new_n8947));
  xor_4  g06599(.A(new_n8914), .B(new_n8913), .Y(new_n8948));
  nand_5 g06600(.A(new_n8948), .B(new_n8947), .Y(new_n8949));
  nand_5 g06601(.A(new_n8949), .B(new_n8915), .Y(new_n8950));
  xor_4  g06602(.A(new_n8910), .B(new_n8909), .Y(new_n8951));
  nor_5  g06603(.A(new_n8951), .B(new_n8950), .Y(new_n8952));
  or_6   g06604(.A(new_n8952), .B(new_n8912), .Y(new_n8953));
  xor_4  g06605(.A(new_n8907), .B(new_n8905), .Y(new_n8954));
  nor_5  g06606(.A(new_n8954), .B(new_n8953), .Y(new_n8955));
  or_6   g06607(.A(new_n8955), .B(new_n8908), .Y(new_n8956));
  not_8  g06608(.A(new_n8903), .Y(new_n8957));
  xor_4  g06609(.A(new_n8957), .B(new_n8902), .Y(new_n8958));
  nor_5  g06610(.A(new_n8958), .B(new_n8956), .Y(new_n8959));
  nor_5  g06611(.A(new_n8959), .B(new_n8904), .Y(new_n8960));
  xor_4  g06612(.A(new_n8900), .B(new_n8863), .Y(new_n8961));
  nor_5  g06613(.A(new_n8961), .B(new_n8960), .Y(new_n8962));
  or_6   g06614(.A(new_n8962), .B(new_n8901), .Y(new_n8963));
  or_6   g06615(.A(new_n8801), .B(new_n8756), .Y(new_n8964));
  or_6   g06616(.A(new_n8862), .B(new_n8803), .Y(new_n8965));
  nand_5 g06617(.A(new_n8965), .B(new_n8964), .Y(new_n8966));
  xor_4  g06618(.A(pi610), .B(new_n7590), .Y(new_n8967));
  nand_5 g06619(.A(new_n8752), .B(new_n8750), .Y(new_n8968));
  nand_5 g06620(.A(new_n8968), .B(new_n8753), .Y(new_n8969));
  xor_4  g06621(.A(new_n8969), .B(new_n8967), .Y(new_n8970));
  not_8  g06622(.A(new_n8970), .Y(new_n8971));
  not_8  g06623(.A(new_n8799), .Y(new_n8972));
  not_8  g06624(.A(new_n8797), .Y(new_n8973));
  nor_5  g06625(.A(new_n8973), .B(new_n8795), .Y(new_n8974));
  nor_5  g06626(.A(new_n8974), .B(new_n8972), .Y(new_n8975));
  not_8  g06627(.A(new_n8975), .Y(new_n8976));
  nand_5 g06628(.A(new_n8976), .B(new_n8971), .Y(new_n8977));
  nand_5 g06629(.A(new_n8975), .B(new_n8970), .Y(new_n8978));
  nand_5 g06630(.A(new_n8978), .B(new_n8977), .Y(new_n8979));
  nand_5 g06631(.A(new_n8052), .B(pi397), .Y(new_n8980));
  not_8  g06632(.A(pi397), .Y(new_n8981));
  nand_5 g06633(.A(pi700), .B(new_n8981), .Y(new_n8982));
  nand_5 g06634(.A(new_n8982), .B(new_n8980), .Y(new_n8983));
  xor_4  g06635(.A(new_n8983), .B(new_n8979), .Y(new_n8984));
  xor_4  g06636(.A(new_n8984), .B(new_n8966), .Y(new_n8985));
  not_8  g06637(.A(pi800), .Y(new_n8986));
  nand_5 g06638(.A(new_n8986), .B(pi335), .Y(new_n8987));
  nand_5 g06639(.A(pi800), .B(new_n6373), .Y(new_n8988));
  nand_5 g06640(.A(new_n8988), .B(new_n8987), .Y(new_n8989));
  nand_5 g06641(.A(pi666), .B(new_n6307), .Y(new_n8990));
  nand_5 g06642(.A(new_n8899), .B(new_n8898), .Y(new_n8991));
  nand_5 g06643(.A(new_n8991), .B(new_n8990), .Y(new_n8992));
  xor_4  g06644(.A(new_n8992), .B(new_n8989), .Y(new_n8993));
  xor_4  g06645(.A(new_n8993), .B(new_n8985), .Y(new_n8994));
  xnor_4 g06646(.A(new_n8994), .B(new_n8963), .Y(po0044));
  xor_4  g06647(.A(new_n7250), .B(pi622), .Y(new_n8996));
  or_6   g06648(.A(pi806), .B(pi745), .Y(new_n8997));
  nand_5 g06649(.A(pi806), .B(pi745), .Y(new_n8998));
  nand_5 g06650(.A(new_n8998), .B(new_n8997), .Y(new_n8999));
  xor_4  g06651(.A(new_n8999), .B(pi642), .Y(new_n9000));
  xor_4  g06652(.A(new_n9000), .B(new_n8996), .Y(po0045));
  not_8  g06653(.A(new_n7745), .Y(new_n9002));
  nand_5 g06654(.A(new_n9002), .B(new_n4516), .Y(new_n9003));
  nand_5 g06655(.A(new_n7789), .B(new_n4373), .Y(new_n9004));
  xor_4  g06656(.A(new_n7789), .B(new_n4373), .Y(new_n9005));
  or_6   g06657(.A(new_n7790), .B(new_n4376), .Y(new_n9006));
  xor_4  g06658(.A(new_n7790), .B(new_n4376), .Y(new_n9007));
  nor_5  g06659(.A(new_n7797), .B(new_n4379), .Y(new_n9008));
  nor_5  g06660(.A(new_n7802), .B(new_n4383), .Y(new_n9009));
  xor_4  g06661(.A(new_n7802), .B(new_n4383), .Y(new_n9010));
  not_8  g06662(.A(new_n9010), .Y(new_n9011));
  or_6   g06663(.A(new_n7807), .B(new_n4386), .Y(new_n9012));
  xor_4  g06664(.A(new_n7807), .B(new_n4386), .Y(new_n9013));
  or_6   g06665(.A(new_n7810), .B(new_n4390), .Y(new_n9014));
  xor_4  g06666(.A(new_n7810), .B(new_n4390), .Y(new_n9015));
  nand_5 g06667(.A(new_n7812), .B(new_n4396), .Y(new_n9016));
  xor_4  g06668(.A(new_n7812), .B(new_n4396), .Y(new_n9017));
  not_8  g06669(.A(new_n7814), .Y(new_n9018));
  or_6   g06670(.A(new_n9018), .B(new_n4398), .Y(new_n9019));
  xor_4  g06671(.A(new_n9018), .B(new_n4398), .Y(new_n9020));
  xor_4  g06672(.A(new_n7821), .B(new_n4411), .Y(new_n9021));
  not_8  g06673(.A(new_n9021), .Y(new_n9022));
  xor_4  g06674(.A(new_n7725), .B(new_n4401), .Y(new_n9023));
  or_6   g06675(.A(new_n7821), .B(new_n4411), .Y(new_n9024));
  not_8  g06676(.A(new_n9024), .Y(new_n9025));
  nand_5 g06677(.A(new_n7818), .B(new_n4403), .Y(new_n9026));
  nor_5  g06678(.A(new_n9026), .B(new_n9025), .Y(new_n9027));
  nor_5  g06679(.A(new_n7818), .B(new_n4403), .Y(new_n9028));
  or_6   g06680(.A(new_n9028), .B(new_n9027), .Y(new_n9029));
  xor_4  g06681(.A(new_n9029), .B(new_n9023), .Y(new_n9030));
  not_8  g06682(.A(new_n9030), .Y(new_n9031));
  nand_5 g06683(.A(new_n9031), .B(new_n9022), .Y(new_n9032));
  not_8  g06684(.A(new_n9032), .Y(new_n9033));
  nor_5  g06685(.A(new_n9033), .B(new_n7829), .Y(new_n9034));
  nor_5  g06686(.A(new_n7725), .B(new_n4401), .Y(new_n9035));
  nand_5 g06687(.A(new_n9027), .B(new_n9035), .Y(new_n9036));
  nand_5 g06688(.A(new_n7837), .B(new_n4402), .Y(new_n9037));
  and_6  g06689(.A(new_n4401), .B(new_n4350), .Y(new_n9038));
  nand_5 g06690(.A(new_n9038), .B(new_n9037), .Y(new_n9039));
  nand_5 g06691(.A(new_n9039), .B(new_n9036), .Y(new_n9040));
  or_6   g06692(.A(new_n9040), .B(new_n9034), .Y(new_n9041));
  nand_5 g06693(.A(new_n9041), .B(new_n9020), .Y(new_n9042));
  nand_5 g06694(.A(new_n9042), .B(new_n9019), .Y(new_n9043));
  nand_5 g06695(.A(new_n9043), .B(new_n9017), .Y(new_n9044));
  nand_5 g06696(.A(new_n9044), .B(new_n9016), .Y(new_n9045));
  nand_5 g06697(.A(new_n9045), .B(new_n9015), .Y(new_n9046));
  nand_5 g06698(.A(new_n9046), .B(new_n9014), .Y(new_n9047));
  nand_5 g06699(.A(new_n9047), .B(new_n9013), .Y(new_n9048));
  nand_5 g06700(.A(new_n9048), .B(new_n9012), .Y(new_n9049));
  nor_5  g06701(.A(new_n9049), .B(new_n9011), .Y(new_n9050));
  nor_5  g06702(.A(new_n9050), .B(new_n9009), .Y(new_n9051));
  xor_4  g06703(.A(new_n7796), .B(new_n4379), .Y(new_n9052));
  not_8  g06704(.A(new_n9052), .Y(new_n9053));
  nand_5 g06705(.A(new_n9053), .B(new_n9051), .Y(new_n9054));
  not_8  g06706(.A(new_n9054), .Y(new_n9055));
  nor_5  g06707(.A(new_n9055), .B(new_n9008), .Y(new_n9056));
  nand_5 g06708(.A(new_n9056), .B(new_n9007), .Y(new_n9057));
  nand_5 g06709(.A(new_n9057), .B(new_n9006), .Y(new_n9058));
  nand_5 g06710(.A(new_n9058), .B(new_n9005), .Y(new_n9059));
  nand_5 g06711(.A(new_n9059), .B(new_n9004), .Y(new_n9060));
  not_8  g06712(.A(new_n9060), .Y(new_n9061));
  nor_5  g06713(.A(new_n9061), .B(new_n9003), .Y(new_n9062));
  nand_5 g06714(.A(new_n7745), .B(new_n4510), .Y(new_n9063));
  nor_5  g06715(.A(new_n9063), .B(new_n9060), .Y(new_n9064));
  nand_5 g06716(.A(new_n9063), .B(new_n9060), .Y(new_n9065));
  nand_5 g06717(.A(new_n9065), .B(new_n9003), .Y(new_n9066));
  nor_5  g06718(.A(new_n9066), .B(new_n9064), .Y(new_n9067));
  nor_5  g06719(.A(new_n9067), .B(new_n9062), .Y(new_n9068));
  xor_4  g06720(.A(new_n9058), .B(new_n9005), .Y(new_n9069));
  not_8  g06721(.A(new_n9069), .Y(new_n9070));
  xor_4  g06722(.A(pi724), .B(new_n5505), .Y(new_n9071));
  or_6   g06723(.A(pi756), .B(new_n5509), .Y(new_n9072));
  xor_4  g06724(.A(pi756), .B(new_n5509), .Y(new_n9073));
  nand_5 g06725(.A(pi492), .B(new_n2908), .Y(new_n9074));
  xor_4  g06726(.A(pi492), .B(new_n2908), .Y(new_n9075));
  nand_5 g06727(.A(new_n2913), .B(pi200), .Y(new_n9076));
  not_8  g06728(.A(pi550), .Y(new_n9077));
  nand_5 g06729(.A(pi836), .B(new_n9077), .Y(new_n9078));
  xor_4  g06730(.A(pi836), .B(new_n9077), .Y(new_n9079));
  nand_5 g06731(.A(pi839), .B(new_n5026), .Y(new_n9080));
  not_8  g06732(.A(pi491), .Y(new_n9081));
  nand_5 g06733(.A(new_n9081), .B(pi214), .Y(new_n9082));
  not_8  g06734(.A(new_n9082), .Y(new_n9083));
  xor_4  g06735(.A(pi839), .B(new_n5026), .Y(new_n9084));
  nand_5 g06736(.A(new_n9084), .B(new_n9083), .Y(new_n9085));
  nand_5 g06737(.A(new_n9085), .B(new_n9080), .Y(new_n9086));
  nand_5 g06738(.A(new_n9086), .B(new_n9079), .Y(new_n9087));
  nand_5 g06739(.A(new_n9087), .B(new_n9078), .Y(new_n9088));
  xor_4  g06740(.A(pi414), .B(pi200), .Y(new_n9089));
  not_8  g06741(.A(new_n9089), .Y(new_n9090));
  nand_5 g06742(.A(new_n9090), .B(new_n9088), .Y(new_n9091));
  nand_5 g06743(.A(new_n9091), .B(new_n9076), .Y(new_n9092));
  nand_5 g06744(.A(new_n9092), .B(new_n9075), .Y(new_n9093));
  nand_5 g06745(.A(new_n9093), .B(new_n9074), .Y(new_n9094));
  nand_5 g06746(.A(new_n9094), .B(new_n9073), .Y(new_n9095));
  nand_5 g06747(.A(new_n9095), .B(new_n9072), .Y(new_n9096));
  xnor_4 g06748(.A(new_n9096), .B(new_n9071), .Y(new_n9097));
  xnor_4 g06749(.A(new_n9094), .B(new_n9073), .Y(new_n9098));
  xor_4  g06750(.A(new_n9045), .B(new_n9015), .Y(new_n9099));
  xor_4  g06751(.A(new_n9092), .B(new_n9075), .Y(new_n9100));
  or_6   g06752(.A(new_n9100), .B(new_n9099), .Y(new_n9101));
  xor_4  g06753(.A(new_n9086), .B(new_n9079), .Y(new_n9102));
  nor_5  g06754(.A(new_n9085), .B(new_n9033), .Y(new_n9103));
  nor_5  g06755(.A(new_n9081), .B(pi214), .Y(new_n9104));
  nand_5 g06756(.A(new_n9104), .B(new_n9021), .Y(new_n9105));
  nand_5 g06757(.A(new_n9083), .B(new_n9022), .Y(new_n9106));
  nand_5 g06758(.A(new_n9106), .B(new_n9105), .Y(new_n9107));
  xor_4  g06759(.A(new_n9107), .B(new_n9084), .Y(new_n9108));
  not_8  g06760(.A(new_n9108), .Y(new_n9109));
  nand_5 g06761(.A(new_n9109), .B(new_n9030), .Y(new_n9110));
  or_6   g06762(.A(new_n9105), .B(new_n9084), .Y(new_n9111));
  nand_5 g06763(.A(new_n9111), .B(new_n9110), .Y(new_n9112));
  nor_5  g06764(.A(new_n9112), .B(new_n9103), .Y(new_n9113));
  nand_5 g06765(.A(new_n9113), .B(new_n9102), .Y(new_n9114));
  not_8  g06766(.A(new_n9114), .Y(new_n9115));
  xnor_4 g06767(.A(new_n9041), .B(new_n9020), .Y(new_n9116));
  xnor_4 g06768(.A(new_n9113), .B(new_n9102), .Y(new_n9117));
  nor_5  g06769(.A(new_n9117), .B(new_n9116), .Y(new_n9118));
  nor_5  g06770(.A(new_n9118), .B(new_n9115), .Y(new_n9119));
  xor_4  g06771(.A(new_n9090), .B(new_n9088), .Y(new_n9120));
  not_8  g06772(.A(new_n9120), .Y(new_n9121));
  nand_5 g06773(.A(new_n9121), .B(new_n9119), .Y(new_n9122));
  xnor_4 g06774(.A(new_n9043), .B(new_n9017), .Y(new_n9123));
  xor_4  g06775(.A(new_n9120), .B(new_n9119), .Y(new_n9124));
  not_8  g06776(.A(new_n9124), .Y(new_n9125));
  nand_5 g06777(.A(new_n9125), .B(new_n9123), .Y(new_n9126));
  nand_5 g06778(.A(new_n9126), .B(new_n9122), .Y(new_n9127));
  xor_4  g06779(.A(new_n9100), .B(new_n9099), .Y(new_n9128));
  nand_5 g06780(.A(new_n9128), .B(new_n9127), .Y(new_n9129));
  nand_5 g06781(.A(new_n9129), .B(new_n9101), .Y(new_n9130));
  nand_5 g06782(.A(new_n9130), .B(new_n9098), .Y(new_n9131));
  xnor_4 g06783(.A(new_n9047), .B(new_n9013), .Y(new_n9132));
  xor_4  g06784(.A(new_n9130), .B(new_n9098), .Y(new_n9133));
  nand_5 g06785(.A(new_n9133), .B(new_n9132), .Y(new_n9134));
  nand_5 g06786(.A(new_n9134), .B(new_n9131), .Y(new_n9135));
  nand_5 g06787(.A(new_n9135), .B(new_n9097), .Y(new_n9136));
  xor_4  g06788(.A(new_n9049), .B(new_n9010), .Y(new_n9137));
  not_8  g06789(.A(new_n9137), .Y(new_n9138));
  xor_4  g06790(.A(new_n9135), .B(new_n9097), .Y(new_n9139));
  nand_5 g06791(.A(new_n9139), .B(new_n9138), .Y(new_n9140));
  nand_5 g06792(.A(new_n9140), .B(new_n9136), .Y(new_n9141));
  xor_4  g06793(.A(pi600), .B(new_n5501), .Y(new_n9142));
  not_8  g06794(.A(pi724), .Y(new_n9143));
  nand_5 g06795(.A(new_n9143), .B(pi549), .Y(new_n9144));
  nand_5 g06796(.A(new_n9096), .B(new_n9071), .Y(new_n9145));
  nand_5 g06797(.A(new_n9145), .B(new_n9144), .Y(new_n9146));
  xor_4  g06798(.A(new_n9146), .B(new_n9142), .Y(new_n9147));
  not_8  g06799(.A(new_n9147), .Y(new_n9148));
  nor_5  g06800(.A(new_n9148), .B(new_n9141), .Y(new_n9149));
  xor_4  g06801(.A(new_n9052), .B(new_n9051), .Y(new_n9150));
  xor_4  g06802(.A(new_n9147), .B(new_n9141), .Y(new_n9151));
  nor_5  g06803(.A(new_n9151), .B(new_n9150), .Y(new_n9152));
  or_6   g06804(.A(new_n9152), .B(new_n9149), .Y(new_n9153));
  not_8  g06805(.A(pi224), .Y(new_n9154));
  xor_4  g06806(.A(pi334), .B(new_n9154), .Y(new_n9155));
  nand_5 g06807(.A(pi600), .B(new_n5501), .Y(new_n9156));
  not_8  g06808(.A(new_n9156), .Y(new_n9157));
  not_8  g06809(.A(new_n9142), .Y(new_n9158));
  nor_5  g06810(.A(new_n9146), .B(new_n9158), .Y(new_n9159));
  nor_5  g06811(.A(new_n9159), .B(new_n9157), .Y(new_n9160));
  xor_4  g06812(.A(new_n9160), .B(new_n9155), .Y(new_n9161));
  nand_5 g06813(.A(new_n9161), .B(new_n9153), .Y(new_n9162));
  xor_4  g06814(.A(new_n9056), .B(new_n9007), .Y(new_n9163));
  xnor_4 g06815(.A(new_n9161), .B(new_n9153), .Y(new_n9164));
  or_6   g06816(.A(new_n9164), .B(new_n9163), .Y(new_n9165));
  nand_5 g06817(.A(new_n9165), .B(new_n9162), .Y(new_n9166));
  nand_5 g06818(.A(new_n9166), .B(new_n9070), .Y(new_n9167));
  not_8  g06819(.A(new_n9167), .Y(new_n9168));
  not_8  g06820(.A(pi512), .Y(new_n9169));
  nand_5 g06821(.A(new_n9169), .B(pi403), .Y(new_n9170));
  not_8  g06822(.A(new_n9170), .Y(new_n9171));
  nand_5 g06823(.A(new_n9171), .B(new_n9168), .Y(new_n9172));
  nor_5  g06824(.A(new_n9169), .B(pi403), .Y(new_n9173));
  not_8  g06825(.A(pi334), .Y(new_n9174));
  nand_5 g06826(.A(new_n9174), .B(pi224), .Y(new_n9175));
  not_8  g06827(.A(new_n9175), .Y(new_n9176));
  not_8  g06828(.A(new_n9155), .Y(new_n9177));
  nor_5  g06829(.A(new_n9160), .B(new_n9177), .Y(new_n9178));
  nor_5  g06830(.A(new_n9178), .B(new_n9176), .Y(new_n9179));
  nor_5  g06831(.A(new_n9179), .B(new_n9171), .Y(new_n9180));
  nor_5  g06832(.A(new_n9180), .B(new_n9173), .Y(new_n9181));
  nor_5  g06833(.A(new_n9181), .B(new_n9167), .Y(new_n9182));
  nor_5  g06834(.A(new_n9166), .B(new_n9070), .Y(new_n9183));
  nor_5  g06835(.A(new_n9183), .B(new_n9168), .Y(new_n9184));
  not_8  g06836(.A(new_n9184), .Y(new_n9185));
  not_8  g06837(.A(new_n9179), .Y(new_n9186));
  nand_5 g06838(.A(new_n9186), .B(new_n9173), .Y(new_n9187));
  nand_5 g06839(.A(new_n9179), .B(new_n9171), .Y(new_n9188));
  nand_5 g06840(.A(new_n9188), .B(new_n9187), .Y(new_n9189));
  nor_5  g06841(.A(new_n9189), .B(new_n9185), .Y(new_n9190));
  nor_5  g06842(.A(new_n9190), .B(new_n9182), .Y(new_n9191));
  nor_5  g06843(.A(new_n9183), .B(new_n9186), .Y(new_n9192));
  nand_5 g06844(.A(new_n9192), .B(new_n9191), .Y(new_n9193));
  nand_5 g06845(.A(new_n9193), .B(new_n9172), .Y(new_n9194));
  nand_5 g06846(.A(new_n9194), .B(new_n9068), .Y(new_n9195));
  nor_5  g06847(.A(new_n9191), .B(new_n9068), .Y(new_n9196));
  not_8  g06848(.A(new_n9068), .Y(new_n9197));
  nor_5  g06849(.A(new_n9189), .B(new_n9183), .Y(new_n9198));
  nor_5  g06850(.A(new_n9198), .B(new_n9181), .Y(new_n9199));
  nor_5  g06851(.A(new_n9199), .B(new_n9197), .Y(new_n9200));
  nand_5 g06852(.A(new_n9183), .B(new_n9181), .Y(new_n9201));
  nand_5 g06853(.A(new_n9201), .B(new_n9197), .Y(new_n9202));
  nand_5 g06854(.A(new_n9202), .B(new_n9167), .Y(new_n9203));
  nor_5  g06855(.A(new_n9203), .B(new_n9200), .Y(new_n9204));
  nor_5  g06856(.A(new_n9204), .B(new_n9196), .Y(new_n9205));
  nand_5 g06857(.A(new_n9205), .B(new_n9195), .Y(po0046));
  not_8  g06858(.A(pi141), .Y(new_n9207));
  xor_4  g06859(.A(pi713), .B(new_n9207), .Y(new_n9208));
  not_8  g06860(.A(new_n9208), .Y(new_n9209));
  not_8  g06861(.A(pi341), .Y(new_n9210));
  nor_5  g06862(.A(pi748), .B(new_n9210), .Y(new_n9211));
  nor_5  g06863(.A(new_n8117), .B(pi341), .Y(new_n9212));
  not_8  g06864(.A(pi203), .Y(new_n9213));
  nor_5  g06865(.A(pi503), .B(new_n9213), .Y(new_n9214));
  xor_4  g06866(.A(pi503), .B(new_n9213), .Y(new_n9215));
  not_8  g06867(.A(new_n9215), .Y(new_n9216));
  not_8  g06868(.A(pi451), .Y(new_n9217));
  nand_5 g06869(.A(pi780), .B(new_n9217), .Y(new_n9218));
  xor_4  g06870(.A(pi780), .B(new_n9217), .Y(new_n9219));
  not_8  g06871(.A(pi363), .Y(new_n9220));
  nand_5 g06872(.A(pi400), .B(new_n9220), .Y(new_n9221));
  xor_4  g06873(.A(pi400), .B(new_n9220), .Y(new_n9222));
  not_8  g06874(.A(pi104), .Y(new_n9223));
  nand_5 g06875(.A(new_n9223), .B(pi003), .Y(new_n9224));
  xor_4  g06876(.A(pi104), .B(new_n8126), .Y(new_n9225));
  not_8  g06877(.A(pi343), .Y(new_n9226));
  nand_5 g06878(.A(pi761), .B(new_n9226), .Y(new_n9227));
  xor_4  g06879(.A(pi761), .B(new_n9226), .Y(new_n9228));
  not_8  g06880(.A(pi090), .Y(new_n9229));
  nand_5 g06881(.A(pi221), .B(new_n9229), .Y(new_n9230));
  xor_4  g06882(.A(pi221), .B(new_n9229), .Y(new_n9231));
  not_8  g06883(.A(pi480), .Y(new_n9232));
  nand_5 g06884(.A(pi741), .B(new_n9232), .Y(new_n9233));
  xor_4  g06885(.A(pi741), .B(new_n9232), .Y(new_n9234));
  not_8  g06886(.A(pi000), .Y(new_n9235));
  nand_5 g06887(.A(pi702), .B(new_n9235), .Y(new_n9236));
  not_8  g06888(.A(new_n9236), .Y(new_n9237));
  nand_5 g06889(.A(new_n9237), .B(new_n9234), .Y(new_n9238));
  nand_5 g06890(.A(new_n9238), .B(new_n9233), .Y(new_n9239));
  nand_5 g06891(.A(new_n9239), .B(new_n9231), .Y(new_n9240));
  nand_5 g06892(.A(new_n9240), .B(new_n9230), .Y(new_n9241));
  nand_5 g06893(.A(new_n9241), .B(new_n9228), .Y(new_n9242));
  nand_5 g06894(.A(new_n9242), .B(new_n9227), .Y(new_n9243));
  nand_5 g06895(.A(new_n9243), .B(new_n9225), .Y(new_n9244));
  nand_5 g06896(.A(new_n9244), .B(new_n9224), .Y(new_n9245));
  nand_5 g06897(.A(new_n9245), .B(new_n9222), .Y(new_n9246));
  nand_5 g06898(.A(new_n9246), .B(new_n9221), .Y(new_n9247));
  nand_5 g06899(.A(new_n9247), .B(new_n9219), .Y(new_n9248));
  nand_5 g06900(.A(new_n9248), .B(new_n9218), .Y(new_n9249));
  nor_5  g06901(.A(new_n9249), .B(new_n9216), .Y(new_n9250));
  nor_5  g06902(.A(new_n9250), .B(new_n9214), .Y(new_n9251));
  nor_5  g06903(.A(new_n9251), .B(new_n9212), .Y(new_n9252));
  nor_5  g06904(.A(new_n9252), .B(new_n9211), .Y(new_n9253));
  xor_4  g06905(.A(new_n9253), .B(pi542), .Y(new_n9254));
  xor_4  g06906(.A(new_n9254), .B(new_n9209), .Y(new_n9255));
  xor_4  g06907(.A(new_n9247), .B(new_n9219), .Y(new_n9256));
  not_8  g06908(.A(new_n9256), .Y(new_n9257));
  xor_4  g06909(.A(new_n9245), .B(new_n9222), .Y(new_n9258));
  not_8  g06910(.A(new_n9258), .Y(new_n9259));
  xor_4  g06911(.A(new_n9243), .B(new_n9225), .Y(new_n9260));
  not_8  g06912(.A(pi048), .Y(new_n9261));
  xnor_4 g06913(.A(new_n9239), .B(new_n9231), .Y(new_n9262));
  not_8  g06914(.A(new_n9234), .Y(new_n9263));
  nand_5 g06915(.A(new_n2558), .B(pi000), .Y(new_n9264));
  nand_5 g06916(.A(new_n9264), .B(pi828), .Y(new_n9265));
  nand_5 g06917(.A(new_n9265), .B(new_n9263), .Y(new_n9266));
  or_6   g06918(.A(new_n9266), .B(new_n9237), .Y(new_n9267));
  not_8  g06919(.A(new_n9238), .Y(new_n9268));
  nor_5  g06920(.A(new_n9265), .B(new_n9263), .Y(new_n9269));
  nor_5  g06921(.A(new_n9269), .B(pi235), .Y(new_n9270));
  nor_5  g06922(.A(new_n9270), .B(new_n9268), .Y(new_n9271));
  nand_5 g06923(.A(new_n9271), .B(new_n9267), .Y(new_n9272));
  or_6   g06924(.A(new_n9272), .B(new_n9262), .Y(new_n9273));
  nand_5 g06925(.A(new_n9273), .B(new_n9261), .Y(new_n9274));
  nand_5 g06926(.A(new_n9272), .B(new_n9262), .Y(new_n9275));
  nand_5 g06927(.A(new_n9275), .B(new_n9274), .Y(new_n9276));
  xor_4  g06928(.A(new_n9241), .B(new_n9228), .Y(new_n9277));
  not_8  g06929(.A(new_n9277), .Y(new_n9278));
  nor_5  g06930(.A(new_n9278), .B(new_n9276), .Y(new_n9279));
  not_8  g06931(.A(pi087), .Y(new_n9280));
  xor_4  g06932(.A(new_n9277), .B(new_n9276), .Y(new_n9281));
  nor_5  g06933(.A(new_n9281), .B(new_n9280), .Y(new_n9282));
  or_6   g06934(.A(new_n9282), .B(new_n9279), .Y(new_n9283));
  or_6   g06935(.A(new_n9283), .B(new_n9260), .Y(new_n9284));
  not_8  g06936(.A(pi083), .Y(new_n9285));
  nand_5 g06937(.A(new_n9283), .B(new_n9260), .Y(new_n9286));
  nand_5 g06938(.A(new_n9286), .B(new_n9285), .Y(new_n9287));
  nand_5 g06939(.A(new_n9287), .B(new_n9284), .Y(new_n9288));
  nand_5 g06940(.A(new_n9288), .B(new_n9259), .Y(new_n9289));
  xor_4  g06941(.A(new_n9288), .B(new_n9258), .Y(new_n9290));
  or_6   g06942(.A(new_n9290), .B(pi099), .Y(new_n9291));
  nand_5 g06943(.A(new_n9291), .B(new_n9289), .Y(new_n9292));
  nor_5  g06944(.A(new_n9292), .B(new_n9257), .Y(new_n9293));
  not_8  g06945(.A(pi462), .Y(new_n9294));
  xor_4  g06946(.A(new_n9292), .B(new_n9256), .Y(new_n9295));
  nor_5  g06947(.A(new_n9295), .B(new_n9294), .Y(new_n9296));
  or_6   g06948(.A(new_n9296), .B(new_n9293), .Y(new_n9297));
  xor_4  g06949(.A(new_n9249), .B(new_n9215), .Y(new_n9298));
  or_6   g06950(.A(new_n9298), .B(new_n9297), .Y(new_n9299));
  nand_5 g06951(.A(new_n9299), .B(pi442), .Y(new_n9300));
  nand_5 g06952(.A(new_n9298), .B(new_n9297), .Y(new_n9301));
  nand_5 g06953(.A(new_n9301), .B(new_n9300), .Y(new_n9302));
  nand_5 g06954(.A(new_n9302), .B(pi108), .Y(new_n9303));
  xor_4  g06955(.A(new_n9302), .B(pi108), .Y(new_n9304));
  nor_5  g06956(.A(new_n9212), .B(new_n9211), .Y(new_n9305));
  xor_4  g06957(.A(new_n9305), .B(new_n9251), .Y(new_n9306));
  nand_5 g06958(.A(new_n9306), .B(new_n9304), .Y(new_n9307));
  nand_5 g06959(.A(new_n9307), .B(new_n9303), .Y(new_n9308));
  xnor_4 g06960(.A(new_n9308), .B(new_n9255), .Y(new_n9309));
  xor_4  g06961(.A(new_n9309), .B(new_n4432), .Y(new_n9310));
  not_8  g06962(.A(new_n9306), .Y(new_n9311));
  xor_4  g06963(.A(new_n9311), .B(new_n9304), .Y(new_n9312));
  nor_5  g06964(.A(new_n9312), .B(new_n4439), .Y(new_n9313));
  xor_4  g06965(.A(new_n9312), .B(new_n4502), .Y(new_n9314));
  nand_5 g06966(.A(new_n9301), .B(new_n9299), .Y(new_n9315));
  xor_4  g06967(.A(new_n9315), .B(pi442), .Y(new_n9316));
  nand_5 g06968(.A(new_n9316), .B(new_n4444), .Y(new_n9317));
  xor_4  g06969(.A(new_n9295), .B(pi462), .Y(new_n9318));
  nor_5  g06970(.A(new_n9318), .B(new_n4448), .Y(new_n9319));
  xor_4  g06971(.A(new_n9318), .B(new_n4449), .Y(new_n9320));
  not_8  g06972(.A(new_n4490), .Y(new_n9321));
  not_8  g06973(.A(pi099), .Y(new_n9322));
  xor_4  g06974(.A(new_n9290), .B(new_n9322), .Y(new_n9323));
  and_6  g06975(.A(new_n9323), .B(new_n9321), .Y(new_n9324));
  xor_4  g06976(.A(new_n9323), .B(new_n4490), .Y(new_n9325));
  nand_5 g06977(.A(new_n9286), .B(new_n9284), .Y(new_n9326));
  xor_4  g06978(.A(new_n9326), .B(pi083), .Y(new_n9327));
  nor_5  g06979(.A(new_n9327), .B(new_n4487), .Y(new_n9328));
  xor_4  g06980(.A(new_n9281), .B(pi087), .Y(new_n9329));
  nand_5 g06981(.A(new_n9329), .B(new_n4454), .Y(new_n9330));
  nand_5 g06982(.A(new_n9275), .B(new_n9273), .Y(new_n9331));
  xor_4  g06983(.A(new_n9331), .B(pi048), .Y(new_n9332));
  or_6   g06984(.A(new_n9332), .B(new_n4460), .Y(new_n9333));
  xor_4  g06985(.A(new_n4468), .B(pi828), .Y(new_n9334));
  nor_5  g06986(.A(new_n9237), .B(new_n9263), .Y(new_n9335));
  nand_5 g06987(.A(new_n9335), .B(new_n9334), .Y(new_n9336));
  nor_5  g06988(.A(new_n4468), .B(pi828), .Y(new_n9337));
  nand_5 g06989(.A(new_n9237), .B(new_n9263), .Y(new_n9338));
  nor_5  g06990(.A(new_n9338), .B(new_n9337), .Y(new_n9339));
  xor_4  g06991(.A(new_n9264), .B(new_n9263), .Y(new_n9340));
  nand_5 g06992(.A(new_n9340), .B(new_n9337), .Y(new_n9341));
  nand_5 g06993(.A(new_n9264), .B(new_n9234), .Y(new_n9342));
  nand_5 g06994(.A(new_n9342), .B(new_n9266), .Y(new_n9343));
  or_6   g06995(.A(new_n9343), .B(new_n4465), .Y(new_n9344));
  nand_5 g06996(.A(new_n9344), .B(new_n9341), .Y(new_n9345));
  nor_5  g06997(.A(new_n9345), .B(new_n9339), .Y(new_n9346));
  nand_5 g06998(.A(new_n9346), .B(new_n9336), .Y(new_n9347));
  xor_4  g06999(.A(new_n9347), .B(pi235), .Y(new_n9348));
  or_6   g07000(.A(new_n9348), .B(new_n4463), .Y(new_n9349));
  nand_5 g07001(.A(new_n9264), .B(new_n9236), .Y(new_n9350));
  not_8  g07002(.A(new_n9350), .Y(new_n9351));
  xor_4  g07003(.A(new_n9351), .B(new_n9334), .Y(po1271));
  or_6   g07004(.A(po1271), .B(new_n4468), .Y(new_n9353));
  nand_5 g07005(.A(new_n9353), .B(new_n9348), .Y(new_n9354));
  nand_5 g07006(.A(new_n9354), .B(new_n9349), .Y(new_n9355));
  xor_4  g07007(.A(new_n9332), .B(new_n4460), .Y(new_n9356));
  nand_5 g07008(.A(new_n9356), .B(new_n9355), .Y(new_n9357));
  nand_5 g07009(.A(new_n9357), .B(new_n9333), .Y(new_n9358));
  xor_4  g07010(.A(new_n9329), .B(new_n4453), .Y(new_n9359));
  or_6   g07011(.A(new_n9359), .B(new_n9358), .Y(new_n9360));
  nand_5 g07012(.A(new_n9360), .B(new_n9330), .Y(new_n9361));
  xnor_4 g07013(.A(new_n9327), .B(new_n4487), .Y(new_n9362));
  nor_5  g07014(.A(new_n9362), .B(new_n9361), .Y(new_n9363));
  nor_5  g07015(.A(new_n9363), .B(new_n9328), .Y(new_n9364));
  nor_5  g07016(.A(new_n9364), .B(new_n9325), .Y(new_n9365));
  nor_5  g07017(.A(new_n9365), .B(new_n9324), .Y(new_n9366));
  nor_5  g07018(.A(new_n9366), .B(new_n9320), .Y(new_n9367));
  or_6   g07019(.A(new_n9367), .B(new_n9319), .Y(new_n9368));
  xor_4  g07020(.A(new_n9316), .B(new_n4443), .Y(new_n9369));
  or_6   g07021(.A(new_n9369), .B(new_n9368), .Y(new_n9370));
  nand_5 g07022(.A(new_n9370), .B(new_n9317), .Y(new_n9371));
  nor_5  g07023(.A(new_n9371), .B(new_n9314), .Y(new_n9372));
  nor_5  g07024(.A(new_n9372), .B(new_n9313), .Y(new_n9373));
  xor_4  g07025(.A(new_n9373), .B(new_n9310), .Y(po0047));
  xnor_4 g07026(.A(new_n9366), .B(new_n9320), .Y(po0048));
  xor_4  g07027(.A(new_n3398), .B(new_n3397), .Y(po0049));
  xnor_4 g07028(.A(new_n4036), .B(new_n4035), .Y(po0050));
  xor_4  g07029(.A(pi645), .B(pi353), .Y(new_n9378));
  nor_5  g07030(.A(pi825), .B(pi475), .Y(new_n9379));
  nor_5  g07031(.A(pi797), .B(pi329), .Y(new_n9380));
  xor_4  g07032(.A(pi797), .B(pi329), .Y(new_n9381));
  nand_5 g07033(.A(pi751), .B(pi295), .Y(new_n9382));
  nand_5 g07034(.A(new_n9382), .B(new_n9381), .Y(new_n9383));
  not_8  g07035(.A(new_n9383), .Y(new_n9384));
  nor_5  g07036(.A(new_n9384), .B(new_n9380), .Y(new_n9385));
  xor_4  g07037(.A(pi825), .B(new_n7720), .Y(new_n9386));
  nor_5  g07038(.A(new_n9386), .B(new_n9385), .Y(new_n9387));
  nor_5  g07039(.A(new_n9387), .B(new_n9379), .Y(new_n9388));
  xor_4  g07040(.A(new_n9388), .B(new_n9378), .Y(new_n9389));
  nor_5  g07041(.A(new_n9381), .B(new_n5953), .Y(new_n9390));
  nor_5  g07042(.A(new_n9390), .B(new_n9384), .Y(new_n9391));
  xor_4  g07043(.A(new_n9381), .B(new_n5953), .Y(new_n9392));
  nor_5  g07044(.A(pi751), .B(pi295), .Y(new_n9393));
  not_8  g07045(.A(new_n9382), .Y(new_n9394));
  nor_5  g07046(.A(new_n9393), .B(new_n9394), .Y(new_n9395));
  not_8  g07047(.A(new_n9395), .Y(new_n9396));
  nor_5  g07048(.A(new_n9396), .B(pi220), .Y(new_n9397));
  nor_5  g07049(.A(new_n9397), .B(new_n9393), .Y(new_n9398));
  nor_5  g07050(.A(new_n9398), .B(new_n9392), .Y(new_n9399));
  nor_5  g07051(.A(new_n9399), .B(new_n9391), .Y(new_n9400));
  nand_5 g07052(.A(new_n9400), .B(pi830), .Y(new_n9401));
  xnor_4 g07053(.A(new_n9400), .B(pi830), .Y(new_n9402));
  xor_4  g07054(.A(new_n9386), .B(new_n9385), .Y(new_n9403));
  or_6   g07055(.A(new_n9403), .B(new_n9402), .Y(new_n9404));
  nand_5 g07056(.A(new_n9404), .B(new_n9401), .Y(new_n9405));
  or_6   g07057(.A(new_n9405), .B(new_n9389), .Y(new_n9406));
  nand_5 g07058(.A(new_n9405), .B(new_n9389), .Y(new_n9407));
  and_6  g07059(.A(new_n9407), .B(new_n9406), .Y(new_n9408));
  xor_4  g07060(.A(new_n9408), .B(pi628), .Y(new_n9409));
  nand_5 g07061(.A(pi214), .B(pi181), .Y(new_n9410));
  not_8  g07062(.A(new_n9410), .Y(new_n9411));
  xor_4  g07063(.A(pi839), .B(new_n2872), .Y(new_n9412));
  xor_4  g07064(.A(new_n9412), .B(new_n9411), .Y(new_n9413));
  not_8  g07065(.A(new_n9413), .Y(new_n9414));
  nand_5 g07066(.A(new_n9414), .B(pi209), .Y(new_n9415));
  xor_4  g07067(.A(pi214), .B(pi181), .Y(new_n9416));
  nand_5 g07068(.A(new_n9416), .B(pi491), .Y(new_n9417));
  not_8  g07069(.A(new_n9417), .Y(new_n9418));
  xor_4  g07070(.A(new_n9413), .B(new_n5026), .Y(new_n9419));
  nand_5 g07071(.A(new_n9419), .B(new_n9418), .Y(new_n9420));
  nand_5 g07072(.A(new_n9420), .B(new_n9415), .Y(new_n9421));
  xor_4  g07073(.A(pi836), .B(pi570), .Y(new_n9422));
  nand_5 g07074(.A(new_n5522), .B(new_n2872), .Y(new_n9423));
  not_8  g07075(.A(new_n9423), .Y(new_n9424));
  nor_5  g07076(.A(new_n9412), .B(new_n9411), .Y(new_n9425));
  nor_5  g07077(.A(new_n9425), .B(new_n9424), .Y(new_n9426));
  xor_4  g07078(.A(new_n9426), .B(new_n9422), .Y(new_n9427));
  or_6   g07079(.A(new_n9427), .B(new_n9421), .Y(new_n9428));
  nand_5 g07080(.A(new_n9428), .B(pi550), .Y(new_n9429));
  nand_5 g07081(.A(new_n9427), .B(new_n9421), .Y(new_n9430));
  nand_5 g07082(.A(new_n9430), .B(new_n9429), .Y(new_n9431));
  xor_4  g07083(.A(new_n9431), .B(new_n2913), .Y(new_n9432));
  xor_4  g07084(.A(pi200), .B(pi151), .Y(new_n9433));
  not_8  g07085(.A(pi836), .Y(new_n9434));
  nand_5 g07086(.A(new_n9434), .B(new_n5246), .Y(new_n9435));
  not_8  g07087(.A(new_n9435), .Y(new_n9436));
  not_8  g07088(.A(new_n9422), .Y(new_n9437));
  nor_5  g07089(.A(new_n9426), .B(new_n9437), .Y(new_n9438));
  nor_5  g07090(.A(new_n9438), .B(new_n9436), .Y(new_n9439));
  xor_4  g07091(.A(new_n9439), .B(new_n9433), .Y(new_n9440));
  xor_4  g07092(.A(new_n9440), .B(new_n9432), .Y(new_n9441));
  nand_5 g07093(.A(new_n9441), .B(new_n9409), .Y(new_n9442));
  xor_4  g07094(.A(new_n9403), .B(new_n9402), .Y(new_n9443));
  xor_4  g07095(.A(new_n9398), .B(new_n9392), .Y(new_n9444));
  not_8  g07096(.A(new_n9444), .Y(new_n9445));
  xor_4  g07097(.A(new_n9395), .B(new_n5778), .Y(new_n9446));
  not_8  g07098(.A(new_n9416), .Y(new_n9447));
  nand_5 g07099(.A(new_n9447), .B(new_n9081), .Y(new_n9448));
  and_6  g07100(.A(new_n9448), .B(new_n9417), .Y(new_n9449));
  nor_5  g07101(.A(new_n9449), .B(new_n9446), .Y(new_n9450));
  nand_5 g07102(.A(new_n9450), .B(new_n9445), .Y(new_n9451));
  nand_5 g07103(.A(new_n9451), .B(new_n9420), .Y(new_n9452));
  nand_5 g07104(.A(new_n9446), .B(new_n9444), .Y(new_n9453));
  nand_5 g07105(.A(new_n9453), .B(new_n9452), .Y(new_n9454));
  nand_5 g07106(.A(new_n9446), .B(new_n9417), .Y(new_n9455));
  not_8  g07107(.A(new_n9446), .Y(new_n9456));
  nand_5 g07108(.A(new_n9448), .B(new_n9456), .Y(new_n9457));
  nand_5 g07109(.A(new_n9457), .B(new_n9455), .Y(new_n9458));
  nand_5 g07110(.A(new_n9458), .B(new_n9444), .Y(new_n9459));
  nor_5  g07111(.A(new_n9419), .B(new_n9418), .Y(new_n9460));
  nand_5 g07112(.A(new_n9460), .B(new_n9459), .Y(new_n9461));
  nand_5 g07113(.A(new_n9461), .B(new_n9454), .Y(new_n9462));
  or_6   g07114(.A(new_n9462), .B(new_n9443), .Y(new_n9463));
  nand_5 g07115(.A(new_n9430), .B(new_n9428), .Y(new_n9464));
  xor_4  g07116(.A(new_n9464), .B(new_n9077), .Y(new_n9465));
  xor_4  g07117(.A(new_n9462), .B(new_n9443), .Y(new_n9466));
  nand_5 g07118(.A(new_n9466), .B(new_n9465), .Y(new_n9467));
  nand_5 g07119(.A(new_n9467), .B(new_n9463), .Y(new_n9468));
  xnor_4 g07120(.A(new_n9441), .B(new_n9409), .Y(new_n9469));
  or_6   g07121(.A(new_n9469), .B(new_n9468), .Y(new_n9470));
  nand_5 g07122(.A(new_n9470), .B(new_n9442), .Y(new_n9471));
  nand_5 g07123(.A(new_n9407), .B(new_n7715), .Y(new_n9472));
  nand_5 g07124(.A(new_n9472), .B(new_n9406), .Y(new_n9473));
  xor_4  g07125(.A(new_n9473), .B(new_n7712), .Y(new_n9474));
  not_8  g07126(.A(new_n9474), .Y(new_n9475));
  xor_4  g07127(.A(pi511), .B(pi432), .Y(new_n9476));
  nand_5 g07128(.A(pi645), .B(pi353), .Y(new_n9477));
  nand_5 g07129(.A(new_n9388), .B(new_n9378), .Y(new_n9478));
  nand_5 g07130(.A(new_n9478), .B(new_n9477), .Y(new_n9479));
  xor_4  g07131(.A(new_n9479), .B(new_n9476), .Y(new_n9480));
  xor_4  g07132(.A(new_n9480), .B(new_n9475), .Y(new_n9481));
  not_8  g07133(.A(new_n9481), .Y(new_n9482));
  nand_5 g07134(.A(new_n5515), .B(new_n2883), .Y(new_n9483));
  not_8  g07135(.A(new_n9483), .Y(new_n9484));
  not_8  g07136(.A(new_n9433), .Y(new_n9485));
  nor_5  g07137(.A(new_n9439), .B(new_n9485), .Y(new_n9486));
  nor_5  g07138(.A(new_n9486), .B(new_n9484), .Y(new_n9487));
  not_8  g07139(.A(pi172), .Y(new_n9488));
  xor_4  g07140(.A(pi492), .B(new_n9488), .Y(new_n9489));
  xor_4  g07141(.A(new_n9489), .B(new_n9487), .Y(new_n9490));
  not_8  g07142(.A(new_n9490), .Y(new_n9491));
  nand_5 g07143(.A(new_n9431), .B(pi414), .Y(new_n9492));
  not_8  g07144(.A(new_n9440), .Y(new_n9493));
  or_6   g07145(.A(new_n9493), .B(new_n9432), .Y(new_n9494));
  nand_5 g07146(.A(new_n9494), .B(new_n9492), .Y(new_n9495));
  nand_5 g07147(.A(new_n9495), .B(new_n9491), .Y(new_n9496));
  or_6   g07148(.A(new_n9495), .B(new_n9491), .Y(new_n9497));
  nand_5 g07149(.A(new_n9497), .B(new_n9496), .Y(new_n9498));
  xor_4  g07150(.A(new_n9498), .B(pi171), .Y(new_n9499));
  or_6   g07151(.A(new_n9499), .B(new_n9482), .Y(new_n9500));
  nand_5 g07152(.A(new_n9500), .B(new_n9471), .Y(new_n9501));
  nand_5 g07153(.A(new_n9499), .B(new_n9482), .Y(new_n9502));
  nand_5 g07154(.A(new_n9502), .B(new_n9501), .Y(new_n9503));
  nand_5 g07155(.A(new_n9473), .B(new_n7712), .Y(new_n9504));
  or_6   g07156(.A(new_n9480), .B(new_n9475), .Y(new_n9505));
  nand_5 g07157(.A(new_n9505), .B(new_n9504), .Y(new_n9506));
  nand_5 g07158(.A(pi511), .B(pi432), .Y(new_n9507));
  nand_5 g07159(.A(new_n9479), .B(new_n9476), .Y(new_n9508));
  nand_5 g07160(.A(new_n9508), .B(new_n9507), .Y(new_n9509));
  not_8  g07161(.A(new_n9509), .Y(new_n9510));
  nand_5 g07162(.A(pi712), .B(pi120), .Y(new_n9511));
  not_8  g07163(.A(pi712), .Y(new_n9512));
  nand_5 g07164(.A(new_n9512), .B(new_n7263), .Y(new_n9513));
  nand_5 g07165(.A(new_n9513), .B(new_n9511), .Y(new_n9514));
  xor_4  g07166(.A(new_n9514), .B(new_n9510), .Y(new_n9515));
  not_8  g07167(.A(new_n9515), .Y(new_n9516));
  nand_5 g07168(.A(new_n9516), .B(new_n9506), .Y(new_n9517));
  or_6   g07169(.A(new_n9516), .B(new_n9506), .Y(new_n9518));
  and_6  g07170(.A(new_n9518), .B(new_n9517), .Y(new_n9519));
  xor_4  g07171(.A(new_n9519), .B(new_n5947), .Y(new_n9520));
  not_8  g07172(.A(new_n9520), .Y(new_n9521));
  nor_5  g07173(.A(new_n9521), .B(new_n9503), .Y(new_n9522));
  xor_4  g07174(.A(new_n9521), .B(new_n9503), .Y(new_n9523));
  not_8  g07175(.A(new_n9523), .Y(new_n9524));
  xor_4  g07176(.A(pi373), .B(pi061), .Y(new_n9525));
  not_8  g07177(.A(pi492), .Y(new_n9526));
  nand_5 g07178(.A(new_n9526), .B(new_n9488), .Y(new_n9527));
  or_6   g07179(.A(new_n9489), .B(new_n9487), .Y(new_n9528));
  nand_5 g07180(.A(new_n9528), .B(new_n9527), .Y(new_n9529));
  xnor_4 g07181(.A(new_n9529), .B(new_n9525), .Y(new_n9530));
  nand_5 g07182(.A(new_n9497), .B(pi171), .Y(new_n9531));
  nand_5 g07183(.A(new_n9531), .B(new_n9496), .Y(new_n9532));
  xor_4  g07184(.A(new_n9532), .B(pi756), .Y(new_n9533));
  not_8  g07185(.A(new_n9533), .Y(new_n9534));
  xor_4  g07186(.A(new_n9534), .B(new_n9530), .Y(new_n9535));
  nor_5  g07187(.A(new_n9535), .B(new_n9524), .Y(new_n9536));
  nor_5  g07188(.A(new_n9536), .B(new_n9522), .Y(new_n9537));
  xor_4  g07189(.A(pi549), .B(pi410), .Y(new_n9538));
  nand_5 g07190(.A(new_n5509), .B(new_n2862), .Y(new_n9539));
  nand_5 g07191(.A(new_n9529), .B(new_n9525), .Y(new_n9540));
  nand_5 g07192(.A(new_n9540), .B(new_n9539), .Y(new_n9541));
  xor_4  g07193(.A(new_n9541), .B(new_n9538), .Y(new_n9542));
  nor_5  g07194(.A(new_n9532), .B(pi756), .Y(new_n9543));
  nor_5  g07195(.A(new_n9534), .B(new_n9530), .Y(new_n9544));
  or_6   g07196(.A(new_n9544), .B(new_n9543), .Y(new_n9545));
  or_6   g07197(.A(new_n9545), .B(new_n9542), .Y(new_n9546));
  nand_5 g07198(.A(new_n9545), .B(new_n9542), .Y(new_n9547));
  nand_5 g07199(.A(new_n9547), .B(new_n9546), .Y(new_n9548));
  xor_4  g07200(.A(new_n9548), .B(pi724), .Y(new_n9549));
  nand_5 g07201(.A(new_n9513), .B(new_n9509), .Y(new_n9550));
  nand_5 g07202(.A(new_n9550), .B(new_n9511), .Y(new_n9551));
  not_8  g07203(.A(new_n9551), .Y(new_n9552));
  nand_5 g07204(.A(pi530), .B(pi146), .Y(new_n9553));
  not_8  g07205(.A(pi530), .Y(new_n9554));
  nand_5 g07206(.A(new_n9554), .B(new_n5940), .Y(new_n9555));
  nand_5 g07207(.A(new_n9555), .B(new_n9553), .Y(new_n9556));
  xor_4  g07208(.A(new_n9556), .B(new_n9552), .Y(new_n9557));
  not_8  g07209(.A(new_n9557), .Y(new_n9558));
  nand_5 g07210(.A(new_n9518), .B(new_n5947), .Y(new_n9559));
  nand_5 g07211(.A(new_n9559), .B(new_n9517), .Y(new_n9560));
  nand_5 g07212(.A(new_n9560), .B(new_n9558), .Y(new_n9561));
  or_6   g07213(.A(new_n9560), .B(new_n9558), .Y(new_n9562));
  nand_5 g07214(.A(new_n9562), .B(new_n9561), .Y(new_n9563));
  xor_4  g07215(.A(new_n9563), .B(pi352), .Y(new_n9564));
  xor_4  g07216(.A(new_n9564), .B(new_n9549), .Y(new_n9565));
  xor_4  g07217(.A(new_n9565), .B(new_n9537), .Y(po0051));
  xor_4  g07218(.A(pi830), .B(pi796), .Y(new_n9567));
  nand_5 g07219(.A(new_n5953), .B(pi619), .Y(new_n9568));
  nand_5 g07220(.A(pi220), .B(new_n4886), .Y(new_n9569));
  nand_5 g07221(.A(pi696), .B(new_n4884), .Y(new_n9570));
  nand_5 g07222(.A(new_n9570), .B(new_n9569), .Y(new_n9571));
  nand_5 g07223(.A(new_n9571), .B(new_n9568), .Y(new_n9572));
  xor_4  g07224(.A(new_n9572), .B(new_n9567), .Y(new_n9573));
  and_6  g07225(.A(new_n9570), .B(new_n9568), .Y(new_n9574));
  xor_4  g07226(.A(new_n9574), .B(new_n9569), .Y(new_n9575));
  not_8  g07227(.A(new_n9575), .Y(new_n9576));
  nand_5 g07228(.A(new_n9576), .B(new_n5760), .Y(new_n9577));
  nor_5  g07229(.A(new_n8609), .B(new_n5762), .Y(new_n9578));
  xor_4  g07230(.A(new_n9575), .B(new_n5760), .Y(new_n9579));
  or_6   g07231(.A(new_n9579), .B(new_n9578), .Y(new_n9580));
  nand_5 g07232(.A(new_n9580), .B(new_n9577), .Y(new_n9581));
  nor_5  g07233(.A(new_n9581), .B(new_n9573), .Y(new_n9582));
  xor_4  g07234(.A(pi514), .B(new_n4347), .Y(new_n9583));
  nand_5 g07235(.A(new_n2360), .B(pi309), .Y(new_n9584));
  nand_5 g07236(.A(new_n5759), .B(new_n5758), .Y(new_n9585));
  nand_5 g07237(.A(new_n9585), .B(new_n9584), .Y(new_n9586));
  xor_4  g07238(.A(new_n9586), .B(new_n9583), .Y(new_n9587));
  not_8  g07239(.A(new_n9573), .Y(new_n9588));
  xor_4  g07240(.A(new_n9581), .B(new_n9588), .Y(new_n9589));
  nor_5  g07241(.A(new_n9589), .B(new_n9587), .Y(new_n9590));
  or_6   g07242(.A(new_n9590), .B(new_n9582), .Y(new_n9591));
  xor_4  g07243(.A(pi628), .B(new_n4900), .Y(new_n9592));
  nand_5 g07244(.A(pi830), .B(new_n8554), .Y(new_n9593));
  not_8  g07245(.A(new_n9593), .Y(new_n9594));
  nor_5  g07246(.A(new_n9572), .B(new_n9567), .Y(new_n9595));
  nor_5  g07247(.A(new_n9595), .B(new_n9594), .Y(new_n9596));
  xor_4  g07248(.A(new_n9596), .B(new_n9592), .Y(new_n9597));
  xor_4  g07249(.A(new_n9597), .B(new_n9591), .Y(new_n9598));
  xor_4  g07250(.A(pi766), .B(pi117), .Y(new_n9599));
  nand_5 g07251(.A(new_n2358), .B(pi504), .Y(new_n9600));
  nand_5 g07252(.A(new_n9586), .B(new_n9583), .Y(new_n9601));
  nand_5 g07253(.A(new_n9601), .B(new_n9600), .Y(new_n9602));
  xor_4  g07254(.A(new_n9602), .B(new_n9599), .Y(new_n9603));
  xor_4  g07255(.A(new_n9603), .B(new_n9598), .Y(new_n9604));
  xor_4  g07256(.A(pi414), .B(new_n8576), .Y(new_n9605));
  nand_5 g07257(.A(pi550), .B(new_n5021), .Y(new_n9606));
  not_8  g07258(.A(new_n9606), .Y(new_n9607));
  xor_4  g07259(.A(pi550), .B(new_n5021), .Y(new_n9608));
  not_8  g07260(.A(new_n9608), .Y(new_n9609));
  nand_5 g07261(.A(pi617), .B(new_n5026), .Y(new_n9610));
  nand_5 g07262(.A(new_n5031), .B(pi209), .Y(new_n9611));
  nand_5 g07263(.A(pi491), .B(new_n5058), .Y(new_n9612));
  nand_5 g07264(.A(new_n9612), .B(new_n9611), .Y(new_n9613));
  nand_5 g07265(.A(new_n9613), .B(new_n9610), .Y(new_n9614));
  nor_5  g07266(.A(new_n9614), .B(new_n9609), .Y(new_n9615));
  nor_5  g07267(.A(new_n9615), .B(new_n9607), .Y(new_n9616));
  xor_4  g07268(.A(new_n9616), .B(new_n9605), .Y(new_n9617));
  xnor_4 g07269(.A(new_n9617), .B(new_n9604), .Y(new_n9618));
  not_8  g07270(.A(new_n9587), .Y(new_n9619));
  xor_4  g07271(.A(new_n9589), .B(new_n9619), .Y(new_n9620));
  xor_4  g07272(.A(new_n9614), .B(new_n9609), .Y(new_n9621));
  or_6   g07273(.A(new_n9621), .B(new_n9620), .Y(new_n9622));
  xor_4  g07274(.A(new_n9621), .B(new_n9620), .Y(new_n9623));
  xor_4  g07275(.A(new_n9579), .B(new_n9578), .Y(new_n9624));
  nand_5 g07276(.A(new_n9611), .B(new_n9610), .Y(new_n9625));
  xor_4  g07277(.A(new_n8609), .B(new_n5762), .Y(new_n9626));
  nand_5 g07278(.A(new_n9081), .B(pi396), .Y(new_n9627));
  nand_5 g07279(.A(new_n9627), .B(new_n9626), .Y(new_n9628));
  not_8  g07280(.A(new_n9626), .Y(new_n9629));
  nand_5 g07281(.A(new_n9629), .B(new_n9612), .Y(new_n9630));
  nand_5 g07282(.A(new_n9630), .B(new_n9628), .Y(new_n9631));
  xnor_4 g07283(.A(new_n9631), .B(new_n9625), .Y(new_n9632));
  nand_5 g07284(.A(new_n9632), .B(new_n9624), .Y(new_n9633));
  not_8  g07285(.A(new_n9632), .Y(new_n9634));
  nand_5 g07286(.A(new_n9627), .B(new_n9612), .Y(new_n9635));
  nand_5 g07287(.A(new_n9635), .B(new_n9626), .Y(new_n9636));
  nand_5 g07288(.A(new_n9636), .B(new_n9634), .Y(new_n9637));
  and_6  g07289(.A(new_n9637), .B(new_n9633), .Y(new_n9638));
  nand_5 g07290(.A(new_n9638), .B(new_n9623), .Y(new_n9639));
  nand_5 g07291(.A(new_n9639), .B(new_n9622), .Y(new_n9640));
  xnor_4 g07292(.A(new_n9640), .B(new_n9618), .Y(po0052));
  xnor_4 g07293(.A(new_n3389), .B(new_n3387), .Y(po0053));
  xor_4  g07294(.A(pi320), .B(pi133), .Y(new_n9643));
  nor_5  g07295(.A(pi371), .B(pi042), .Y(new_n9644));
  xor_4  g07296(.A(pi371), .B(pi042), .Y(new_n9645));
  not_8  g07297(.A(new_n9645), .Y(new_n9646));
  nor_5  g07298(.A(pi824), .B(pi658), .Y(new_n9647));
  not_8  g07299(.A(pi658), .Y(new_n9648));
  xor_4  g07300(.A(pi824), .B(new_n9648), .Y(new_n9649));
  not_8  g07301(.A(pi255), .Y(new_n9650));
  not_8  g07302(.A(pi821), .Y(new_n9651));
  nor_5  g07303(.A(new_n9651), .B(new_n9650), .Y(new_n9652));
  nor_5  g07304(.A(new_n9652), .B(new_n9649), .Y(new_n9653));
  nor_5  g07305(.A(new_n9653), .B(new_n9647), .Y(new_n9654));
  nor_5  g07306(.A(new_n9654), .B(new_n9646), .Y(new_n9655));
  nor_5  g07307(.A(new_n9655), .B(new_n9644), .Y(new_n9656));
  xor_4  g07308(.A(new_n9656), .B(new_n9643), .Y(new_n9657));
  nor_5  g07309(.A(new_n6758), .B(pi535), .Y(new_n9658));
  not_8  g07310(.A(pi535), .Y(new_n9659));
  xor_4  g07311(.A(new_n6758), .B(new_n9659), .Y(new_n9660));
  nand_5 g07312(.A(new_n6762), .B(pi719), .Y(new_n9661));
  or_6   g07313(.A(new_n6762), .B(pi719), .Y(new_n9662));
  nand_5 g07314(.A(new_n6767), .B(pi580), .Y(new_n9663));
  nand_5 g07315(.A(new_n9663), .B(new_n6729), .Y(new_n9664));
  xor_4  g07316(.A(new_n9664), .B(new_n6765), .Y(new_n9665));
  or_6   g07317(.A(new_n9665), .B(new_n2638), .Y(new_n9666));
  nand_5 g07318(.A(new_n9664), .B(new_n6773), .Y(new_n9667));
  nand_5 g07319(.A(new_n9667), .B(new_n9666), .Y(new_n9668));
  nand_5 g07320(.A(new_n9668), .B(new_n9662), .Y(new_n9669));
  nand_5 g07321(.A(new_n9669), .B(new_n9661), .Y(new_n9670));
  nor_5  g07322(.A(new_n9670), .B(new_n9660), .Y(new_n9671));
  nor_5  g07323(.A(new_n9671), .B(new_n9658), .Y(new_n9672));
  nand_5 g07324(.A(new_n6753), .B(new_n8727), .Y(new_n9673));
  nand_5 g07325(.A(new_n6752), .B(pi173), .Y(new_n9674));
  nand_5 g07326(.A(new_n9674), .B(new_n9673), .Y(new_n9675));
  xor_4  g07327(.A(new_n9675), .B(new_n9672), .Y(new_n9676));
  xor_4  g07328(.A(new_n9676), .B(pi594), .Y(new_n9677));
  not_8  g07329(.A(pi694), .Y(new_n9678));
  nand_5 g07330(.A(new_n7251), .B(pi806), .Y(new_n9679));
  or_6   g07331(.A(new_n9679), .B(new_n9678), .Y(new_n9680));
  xor_4  g07332(.A(new_n9665), .B(new_n2638), .Y(new_n9681));
  not_8  g07333(.A(new_n9681), .Y(new_n9682));
  xor_4  g07334(.A(new_n9679), .B(new_n9678), .Y(new_n9683));
  nand_5 g07335(.A(new_n9683), .B(new_n9682), .Y(new_n9684));
  nand_5 g07336(.A(new_n9684), .B(new_n9680), .Y(new_n9685));
  nand_5 g07337(.A(new_n9685), .B(pi529), .Y(new_n9686));
  nand_5 g07338(.A(new_n9662), .B(new_n9661), .Y(new_n9687));
  xor_4  g07339(.A(new_n9687), .B(new_n9668), .Y(new_n9688));
  not_8  g07340(.A(new_n9688), .Y(new_n9689));
  not_8  g07341(.A(pi529), .Y(new_n9690));
  xor_4  g07342(.A(new_n9685), .B(new_n9690), .Y(new_n9691));
  or_6   g07343(.A(new_n9691), .B(new_n9689), .Y(new_n9692));
  nand_5 g07344(.A(new_n9692), .B(new_n9686), .Y(new_n9693));
  nor_5  g07345(.A(new_n9693), .B(pi478), .Y(new_n9694));
  xor_4  g07346(.A(new_n9670), .B(new_n9660), .Y(new_n9695));
  not_8  g07347(.A(pi478), .Y(new_n9696));
  xor_4  g07348(.A(new_n9693), .B(new_n9696), .Y(new_n9697));
  nor_5  g07349(.A(new_n9697), .B(new_n9695), .Y(new_n9698));
  or_6   g07350(.A(new_n9698), .B(new_n9694), .Y(new_n9699));
  xnor_4 g07351(.A(new_n9699), .B(new_n9677), .Y(new_n9700));
  xor_4  g07352(.A(new_n9700), .B(new_n9657), .Y(new_n9701));
  not_8  g07353(.A(new_n9701), .Y(new_n9702));
  xor_4  g07354(.A(new_n9652), .B(new_n9649), .Y(new_n9703));
  xor_4  g07355(.A(pi821), .B(pi255), .Y(new_n9704));
  not_8  g07356(.A(new_n9704), .Y(new_n9705));
  nand_5 g07357(.A(new_n7252), .B(new_n7248), .Y(new_n9706));
  nand_5 g07358(.A(new_n9706), .B(new_n7246), .Y(new_n9707));
  nand_5 g07359(.A(new_n9707), .B(new_n9705), .Y(new_n9708));
  xor_4  g07360(.A(new_n9683), .B(new_n9681), .Y(new_n9709));
  xor_4  g07361(.A(new_n9707), .B(new_n9705), .Y(new_n9710));
  nand_5 g07362(.A(new_n9710), .B(new_n9709), .Y(new_n9711));
  nand_5 g07363(.A(new_n9711), .B(new_n9708), .Y(new_n9712));
  nand_5 g07364(.A(new_n9712), .B(new_n9703), .Y(new_n9713));
  xor_4  g07365(.A(new_n9712), .B(new_n9703), .Y(new_n9714));
  xor_4  g07366(.A(new_n9691), .B(new_n9688), .Y(new_n9715));
  nand_5 g07367(.A(new_n9715), .B(new_n9714), .Y(new_n9716));
  nand_5 g07368(.A(new_n9716), .B(new_n9713), .Y(new_n9717));
  xor_4  g07369(.A(new_n9654), .B(new_n9645), .Y(new_n9718));
  not_8  g07370(.A(new_n9718), .Y(new_n9719));
  nor_5  g07371(.A(new_n9719), .B(new_n9717), .Y(new_n9720));
  xor_4  g07372(.A(new_n9718), .B(new_n9717), .Y(new_n9721));
  xor_4  g07373(.A(new_n9697), .B(new_n9695), .Y(new_n9722));
  nor_5  g07374(.A(new_n9722), .B(new_n9721), .Y(new_n9723));
  or_6   g07375(.A(new_n9723), .B(new_n9720), .Y(new_n9724));
  xor_4  g07376(.A(new_n9724), .B(new_n9702), .Y(po0054));
  xor_4  g07377(.A(new_n2615), .B(pi784), .Y(new_n9726));
  or_6   g07378(.A(new_n2620), .B(pi734), .Y(new_n9727));
  not_8  g07379(.A(new_n9727), .Y(new_n9728));
  xor_4  g07380(.A(new_n2620), .B(pi734), .Y(new_n9729));
  not_8  g07381(.A(new_n9729), .Y(new_n9730));
  nand_5 g07382(.A(new_n2623), .B(pi395), .Y(new_n9731));
  or_6   g07383(.A(new_n2626), .B(pi351), .Y(new_n9732));
  not_8  g07384(.A(new_n9732), .Y(new_n9733));
  xor_4  g07385(.A(new_n2626), .B(pi351), .Y(new_n9734));
  not_8  g07386(.A(new_n9734), .Y(new_n9735));
  nand_5 g07387(.A(new_n2629), .B(pi497), .Y(new_n9736));
  xor_4  g07388(.A(new_n2629), .B(pi497), .Y(new_n9737));
  nand_5 g07389(.A(new_n2632), .B(pi506), .Y(new_n9738));
  or_6   g07390(.A(new_n2632), .B(pi506), .Y(new_n9739));
  nand_5 g07391(.A(new_n2634), .B(pi374), .Y(new_n9740));
  xor_4  g07392(.A(new_n2634), .B(pi374), .Y(new_n9741));
  nor_5  g07393(.A(new_n2639), .B(new_n3905), .Y(new_n9742));
  xor_4  g07394(.A(new_n2639), .B(new_n3905), .Y(new_n9743));
  not_8  g07395(.A(new_n9743), .Y(new_n9744));
  nand_5 g07396(.A(new_n2643), .B(new_n2565), .Y(new_n9745));
  nand_5 g07397(.A(new_n9745), .B(new_n2644), .Y(new_n9746));
  nor_5  g07398(.A(new_n9746), .B(new_n9744), .Y(new_n9747));
  or_6   g07399(.A(new_n9747), .B(new_n9742), .Y(new_n9748));
  nand_5 g07400(.A(new_n9748), .B(new_n9741), .Y(new_n9749));
  nand_5 g07401(.A(new_n9749), .B(new_n9740), .Y(new_n9750));
  nand_5 g07402(.A(new_n9750), .B(new_n9739), .Y(new_n9751));
  nand_5 g07403(.A(new_n9751), .B(new_n9738), .Y(new_n9752));
  nand_5 g07404(.A(new_n9752), .B(new_n9737), .Y(new_n9753));
  nand_5 g07405(.A(new_n9753), .B(new_n9736), .Y(new_n9754));
  nor_5  g07406(.A(new_n9754), .B(new_n9735), .Y(new_n9755));
  nor_5  g07407(.A(new_n9755), .B(new_n9733), .Y(new_n9756));
  xor_4  g07408(.A(new_n2623), .B(new_n4266), .Y(new_n9757));
  not_8  g07409(.A(new_n9757), .Y(new_n9758));
  nand_5 g07410(.A(new_n9758), .B(new_n9756), .Y(new_n9759));
  nand_5 g07411(.A(new_n9759), .B(new_n9731), .Y(new_n9760));
  nor_5  g07412(.A(new_n9760), .B(new_n9730), .Y(new_n9761));
  nor_5  g07413(.A(new_n9761), .B(new_n9728), .Y(new_n9762));
  xor_4  g07414(.A(new_n9762), .B(new_n9726), .Y(new_n9763));
  not_8  g07415(.A(new_n9763), .Y(new_n9764));
  nand_5 g07416(.A(new_n2737), .B(pi380), .Y(new_n9765));
  not_8  g07417(.A(new_n2699), .Y(new_n9766));
  nand_5 g07418(.A(new_n2716), .B(new_n2949), .Y(new_n9767));
  xor_4  g07419(.A(new_n2716), .B(pi766), .Y(new_n9768));
  nand_5 g07420(.A(new_n2707), .B(pi309), .Y(new_n9769));
  or_6   g07421(.A(new_n9769), .B(new_n4347), .Y(new_n9770));
  nand_5 g07422(.A(new_n9769), .B(new_n4347), .Y(new_n9771));
  nand_5 g07423(.A(new_n9771), .B(new_n2711), .Y(new_n9772));
  nand_5 g07424(.A(new_n9772), .B(new_n9770), .Y(new_n9773));
  or_6   g07425(.A(new_n9773), .B(new_n9768), .Y(new_n9774));
  nand_5 g07426(.A(new_n9774), .B(new_n9767), .Y(new_n9775));
  or_6   g07427(.A(new_n9775), .B(new_n2966), .Y(new_n9776));
  xor_4  g07428(.A(new_n9775), .B(new_n2966), .Y(new_n9777));
  nand_5 g07429(.A(new_n9777), .B(new_n2702), .Y(new_n9778));
  nand_5 g07430(.A(new_n9778), .B(new_n9776), .Y(new_n9779));
  nand_5 g07431(.A(new_n9779), .B(new_n9766), .Y(new_n9780));
  nor_5  g07432(.A(new_n9779), .B(new_n9766), .Y(new_n9781));
  not_8  g07433(.A(new_n9781), .Y(new_n9782));
  nand_5 g07434(.A(new_n9782), .B(pi636), .Y(new_n9783));
  and_6  g07435(.A(new_n9783), .B(new_n9780), .Y(new_n9784));
  nor_5  g07436(.A(new_n9784), .B(new_n2696), .Y(new_n9785));
  xor_4  g07437(.A(new_n9784), .B(new_n2697), .Y(new_n9786));
  nor_5  g07438(.A(new_n9786), .B(new_n2943), .Y(new_n9787));
  or_6   g07439(.A(new_n9787), .B(new_n9785), .Y(new_n9788));
  xor_4  g07440(.A(new_n2737), .B(pi380), .Y(new_n9789));
  nand_5 g07441(.A(new_n9789), .B(new_n9788), .Y(new_n9790));
  nand_5 g07442(.A(new_n9790), .B(new_n9765), .Y(new_n9791));
  xor_4  g07443(.A(new_n2820), .B(new_n4335), .Y(new_n9792));
  xor_4  g07444(.A(new_n9792), .B(new_n9791), .Y(new_n9793));
  xor_4  g07445(.A(new_n9793), .B(new_n9764), .Y(new_n9794));
  xor_4  g07446(.A(new_n9789), .B(new_n9788), .Y(new_n9795));
  xor_4  g07447(.A(new_n9760), .B(new_n9729), .Y(new_n9796));
  not_8  g07448(.A(new_n9796), .Y(new_n9797));
  and_6  g07449(.A(new_n9797), .B(new_n9795), .Y(new_n9798));
  xor_4  g07450(.A(new_n9796), .B(new_n9795), .Y(new_n9799));
  xor_4  g07451(.A(new_n9777), .B(new_n2702), .Y(new_n9800));
  xor_4  g07452(.A(new_n9748), .B(new_n9741), .Y(new_n9801));
  not_8  g07453(.A(new_n9801), .Y(new_n9802));
  xor_4  g07454(.A(new_n9746), .B(new_n9744), .Y(new_n9803));
  nand_5 g07455(.A(new_n2748), .B(new_n3020), .Y(new_n9804));
  xor_4  g07456(.A(new_n2748), .B(pi062), .Y(new_n9805));
  not_8  g07457(.A(new_n9805), .Y(new_n9806));
  xor_4  g07458(.A(new_n2566), .B(pi580), .Y(new_n9807));
  not_8  g07459(.A(new_n9807), .Y(new_n9808));
  nand_5 g07460(.A(new_n9808), .B(new_n9806), .Y(new_n9809));
  nand_5 g07461(.A(new_n9809), .B(new_n9804), .Y(new_n9810));
  nor_5  g07462(.A(new_n9810), .B(new_n9803), .Y(new_n9811));
  and_6  g07463(.A(new_n9810), .B(new_n9803), .Y(new_n9812));
  xor_4  g07464(.A(new_n2706), .B(pi309), .Y(new_n9813));
  nor_5  g07465(.A(new_n9813), .B(new_n9812), .Y(new_n9814));
  or_6   g07466(.A(new_n9814), .B(new_n9811), .Y(new_n9815));
  or_6   g07467(.A(new_n9815), .B(new_n9802), .Y(new_n9816));
  xor_4  g07468(.A(new_n9815), .B(new_n9802), .Y(new_n9817));
  nand_5 g07469(.A(new_n9771), .B(new_n9770), .Y(new_n9818));
  xor_4  g07470(.A(new_n9818), .B(new_n2711), .Y(new_n9819));
  nand_5 g07471(.A(new_n9819), .B(new_n9817), .Y(new_n9820));
  nand_5 g07472(.A(new_n9820), .B(new_n9816), .Y(new_n9821));
  and_6  g07473(.A(new_n9739), .B(new_n9738), .Y(new_n9822));
  xor_4  g07474(.A(new_n9822), .B(new_n9750), .Y(new_n9823));
  nand_5 g07475(.A(new_n9823), .B(new_n9821), .Y(new_n9824));
  xor_4  g07476(.A(new_n9773), .B(new_n9768), .Y(new_n9825));
  xor_4  g07477(.A(new_n9823), .B(new_n9821), .Y(new_n9826));
  nand_5 g07478(.A(new_n9826), .B(new_n9825), .Y(new_n9827));
  and_6  g07479(.A(new_n9827), .B(new_n9824), .Y(new_n9828));
  nand_5 g07480(.A(new_n9828), .B(new_n9800), .Y(new_n9829));
  xor_4  g07481(.A(new_n9752), .B(new_n9737), .Y(new_n9830));
  not_8  g07482(.A(new_n9830), .Y(new_n9831));
  xor_4  g07483(.A(new_n9828), .B(new_n9800), .Y(new_n9832));
  nand_5 g07484(.A(new_n9832), .B(new_n9831), .Y(new_n9833));
  nand_5 g07485(.A(new_n9833), .B(new_n9829), .Y(new_n9834));
  xor_4  g07486(.A(new_n9754), .B(new_n9734), .Y(new_n9835));
  not_8  g07487(.A(new_n9835), .Y(new_n9836));
  nand_5 g07488(.A(new_n9836), .B(new_n9834), .Y(new_n9837));
  xor_4  g07489(.A(new_n9835), .B(new_n9834), .Y(new_n9838));
  nand_5 g07490(.A(new_n9780), .B(new_n9782), .Y(new_n9839));
  xor_4  g07491(.A(new_n9839), .B(pi636), .Y(new_n9840));
  or_6   g07492(.A(new_n9840), .B(new_n9838), .Y(new_n9841));
  nand_5 g07493(.A(new_n9841), .B(new_n9837), .Y(new_n9842));
  xor_4  g07494(.A(new_n9757), .B(new_n9756), .Y(new_n9843));
  nor_5  g07495(.A(new_n9843), .B(new_n9842), .Y(new_n9844));
  xor_4  g07496(.A(new_n9843), .B(new_n9842), .Y(new_n9845));
  not_8  g07497(.A(new_n9845), .Y(new_n9846));
  xor_4  g07498(.A(new_n9786), .B(new_n2943), .Y(new_n9847));
  nor_5  g07499(.A(new_n9847), .B(new_n9846), .Y(new_n9848));
  or_6   g07500(.A(new_n9848), .B(new_n9844), .Y(new_n9849));
  nor_5  g07501(.A(new_n9849), .B(new_n9799), .Y(new_n9850));
  nor_5  g07502(.A(new_n9850), .B(new_n9798), .Y(new_n9851));
  xnor_4 g07503(.A(new_n9851), .B(new_n9794), .Y(po0055));
  xor_4  g07504(.A(new_n7946), .B(new_n7945), .Y(po0056));
  nand_5 g07505(.A(new_n3491), .B(pi130), .Y(new_n9854));
  nand_5 g07506(.A(pi301), .B(new_n4886), .Y(new_n9855));
  nand_5 g07507(.A(new_n9855), .B(new_n9854), .Y(new_n9856));
  not_8  g07508(.A(new_n9856), .Y(new_n9857));
  xor_4  g07509(.A(new_n9857), .B(new_n7819), .Y(new_n9858));
  nand_5 g07510(.A(pi396), .B(new_n7054), .Y(new_n9859));
  nand_5 g07511(.A(new_n5058), .B(pi238), .Y(new_n9860));
  nand_5 g07512(.A(new_n9860), .B(new_n9859), .Y(new_n9861));
  xor_4  g07513(.A(new_n9861), .B(new_n9858), .Y(po0057));
  xor_4  g07514(.A(pi501), .B(pi486), .Y(new_n9863));
  nand_5 g07515(.A(new_n2392), .B(pi589), .Y(new_n9864));
  nand_5 g07516(.A(pi611), .B(new_n2484), .Y(new_n9865));
  nand_5 g07517(.A(new_n9865), .B(new_n2428), .Y(new_n9866));
  nand_5 g07518(.A(new_n9866), .B(new_n9864), .Y(new_n9867));
  xor_4  g07519(.A(new_n9867), .B(new_n9863), .Y(new_n9868));
  xor_4  g07520(.A(new_n9868), .B(new_n7920), .Y(new_n9869));
  not_8  g07521(.A(new_n7931), .Y(new_n9870));
  nand_5 g07522(.A(new_n9864), .B(new_n9865), .Y(new_n9871));
  not_8  g07523(.A(new_n9871), .Y(new_n9872));
  nor_5  g07524(.A(new_n2428), .B(pi077), .Y(new_n9873));
  nand_5 g07525(.A(new_n9873), .B(new_n7925), .Y(new_n9874));
  nand_5 g07526(.A(new_n2428), .B(pi077), .Y(new_n9875));
  or_6   g07527(.A(new_n9875), .B(new_n7925), .Y(new_n9876));
  nand_5 g07528(.A(new_n9876), .B(new_n9874), .Y(new_n9877));
  xor_4  g07529(.A(new_n9877), .B(new_n9872), .Y(new_n9878));
  nor_5  g07530(.A(new_n9878), .B(new_n9870), .Y(new_n9879));
  or_6   g07531(.A(new_n9877), .B(new_n9871), .Y(new_n9880));
  nor_5  g07532(.A(new_n9880), .B(pi223), .Y(new_n9881));
  nor_5  g07533(.A(new_n9874), .B(new_n9872), .Y(new_n9882));
  or_6   g07534(.A(new_n9882), .B(new_n9881), .Y(new_n9883));
  nor_5  g07535(.A(new_n9883), .B(new_n9879), .Y(new_n9884));
  xnor_4 g07536(.A(new_n9884), .B(new_n9869), .Y(po0058));
  not_8  g07537(.A(new_n5753), .Y(new_n9886));
  xor_4  g07538(.A(new_n9886), .B(new_n5752), .Y(po0059));
  not_8  g07539(.A(pi186), .Y(new_n9888));
  xor_4  g07540(.A(pi470), .B(new_n9888), .Y(new_n9889));
  not_8  g07541(.A(new_n9889), .Y(new_n9890));
  nand_5 g07542(.A(pi372), .B(pi134), .Y(new_n9891));
  not_8  g07543(.A(pi134), .Y(new_n9892));
  or_6   g07544(.A(pi372), .B(new_n9892), .Y(new_n9893));
  nand_5 g07545(.A(pi372), .B(new_n9892), .Y(new_n9894));
  nand_5 g07546(.A(new_n9894), .B(new_n9893), .Y(new_n9895));
  nand_5 g07547(.A(pi723), .B(pi001), .Y(new_n9896));
  xor_4  g07548(.A(pi723), .B(pi001), .Y(new_n9897));
  nor_5  g07549(.A(pi206), .B(pi050), .Y(new_n9898));
  xor_4  g07550(.A(pi206), .B(pi050), .Y(new_n9899));
  not_8  g07551(.A(new_n9899), .Y(new_n9900));
  nor_5  g07552(.A(pi262), .B(pi212), .Y(new_n9901));
  xor_4  g07553(.A(pi262), .B(pi212), .Y(new_n9902));
  nand_5 g07554(.A(pi620), .B(pi326), .Y(new_n9903));
  and_6  g07555(.A(new_n9903), .B(new_n9902), .Y(new_n9904));
  nor_5  g07556(.A(new_n9904), .B(new_n9901), .Y(new_n9905));
  nor_5  g07557(.A(new_n9905), .B(new_n9900), .Y(new_n9906));
  nor_5  g07558(.A(new_n9906), .B(new_n9898), .Y(new_n9907));
  nand_5 g07559(.A(new_n9907), .B(new_n9897), .Y(new_n9908));
  nand_5 g07560(.A(new_n9908), .B(new_n9896), .Y(new_n9909));
  nand_5 g07561(.A(new_n9909), .B(new_n9895), .Y(new_n9910));
  nand_5 g07562(.A(new_n9910), .B(new_n9891), .Y(new_n9911));
  xor_4  g07563(.A(new_n9911), .B(new_n9890), .Y(new_n9912));
  xor_4  g07564(.A(new_n9912), .B(pi780), .Y(new_n9913));
  xor_4  g07565(.A(new_n9909), .B(new_n9895), .Y(new_n9914));
  or_6   g07566(.A(new_n9914), .B(pi400), .Y(new_n9915));
  xor_4  g07567(.A(new_n9914), .B(pi400), .Y(new_n9916));
  xor_4  g07568(.A(new_n9907), .B(new_n9897), .Y(new_n9917));
  or_6   g07569(.A(new_n9917), .B(pi003), .Y(new_n9918));
  xor_4  g07570(.A(new_n9917), .B(pi003), .Y(new_n9919));
  xor_4  g07571(.A(new_n9905), .B(new_n9899), .Y(new_n9920));
  and_6  g07572(.A(new_n9920), .B(pi761), .Y(new_n9921));
  xor_4  g07573(.A(new_n9920), .B(pi761), .Y(new_n9922));
  not_8  g07574(.A(new_n9922), .Y(new_n9923));
  xor_4  g07575(.A(new_n9903), .B(new_n9902), .Y(new_n9924));
  nand_5 g07576(.A(new_n9924), .B(new_n4288), .Y(new_n9925));
  xor_4  g07577(.A(pi620), .B(pi326), .Y(new_n9926));
  not_8  g07578(.A(new_n9926), .Y(new_n9927));
  nor_5  g07579(.A(new_n9927), .B(new_n4282), .Y(new_n9928));
  xor_4  g07580(.A(new_n9926), .B(pi741), .Y(new_n9929));
  not_8  g07581(.A(new_n9929), .Y(new_n9930));
  nand_5 g07582(.A(pi494), .B(new_n8025), .Y(new_n9931));
  not_8  g07583(.A(pi494), .Y(new_n9932));
  nand_5 g07584(.A(new_n9932), .B(pi122), .Y(new_n9933));
  nand_5 g07585(.A(new_n9933), .B(new_n9931), .Y(new_n9934));
  not_8  g07586(.A(new_n9934), .Y(new_n9935));
  nor_5  g07587(.A(new_n9935), .B(new_n2558), .Y(new_n9936));
  nor_5  g07588(.A(new_n9932), .B(new_n8025), .Y(new_n9937));
  nor_5  g07589(.A(new_n9937), .B(new_n9936), .Y(new_n9938));
  nor_5  g07590(.A(new_n9938), .B(new_n9930), .Y(new_n9939));
  nor_5  g07591(.A(new_n9939), .B(new_n9928), .Y(new_n9940));
  xor_4  g07592(.A(new_n9924), .B(pi221), .Y(new_n9941));
  not_8  g07593(.A(new_n9941), .Y(new_n9942));
  nand_5 g07594(.A(new_n9942), .B(new_n9940), .Y(new_n9943));
  nand_5 g07595(.A(new_n9943), .B(new_n9925), .Y(new_n9944));
  nor_5  g07596(.A(new_n9944), .B(new_n9923), .Y(new_n9945));
  nor_5  g07597(.A(new_n9945), .B(new_n9921), .Y(new_n9946));
  nand_5 g07598(.A(new_n9946), .B(new_n9919), .Y(new_n9947));
  nand_5 g07599(.A(new_n9947), .B(new_n9918), .Y(new_n9948));
  nand_5 g07600(.A(new_n9948), .B(new_n9916), .Y(new_n9949));
  nand_5 g07601(.A(new_n9949), .B(new_n9915), .Y(new_n9950));
  xor_4  g07602(.A(new_n9950), .B(new_n9913), .Y(new_n9951));
  xor_4  g07603(.A(pi764), .B(pi274), .Y(new_n9952));
  nor_5  g07604(.A(pi398), .B(pi075), .Y(new_n9953));
  nor_5  g07605(.A(pi698), .B(pi639), .Y(new_n9954));
  nor_5  g07606(.A(pi754), .B(pi515), .Y(new_n9955));
  nand_5 g07607(.A(pi474), .B(pi080), .Y(new_n9956));
  not_8  g07608(.A(new_n9956), .Y(new_n9957));
  xor_4  g07609(.A(pi754), .B(new_n8075), .Y(new_n9958));
  nor_5  g07610(.A(new_n9958), .B(new_n9957), .Y(new_n9959));
  nor_5  g07611(.A(new_n9959), .B(new_n9955), .Y(new_n9960));
  xor_4  g07612(.A(pi698), .B(new_n8158), .Y(new_n9961));
  nor_5  g07613(.A(new_n9961), .B(new_n9960), .Y(new_n9962));
  nor_5  g07614(.A(new_n9962), .B(new_n9954), .Y(new_n9963));
  xor_4  g07615(.A(pi398), .B(new_n8086), .Y(new_n9964));
  nor_5  g07616(.A(new_n9964), .B(new_n9963), .Y(new_n9965));
  or_6   g07617(.A(new_n9965), .B(new_n9953), .Y(new_n9966));
  xnor_4 g07618(.A(new_n9966), .B(new_n9952), .Y(new_n9967));
  xor_4  g07619(.A(new_n9967), .B(pi222), .Y(new_n9968));
  not_8  g07620(.A(pi704), .Y(new_n9969));
  xor_4  g07621(.A(new_n9964), .B(new_n9963), .Y(new_n9970));
  or_6   g07622(.A(new_n9970), .B(new_n9969), .Y(new_n9971));
  xnor_4 g07623(.A(new_n9961), .B(new_n9960), .Y(new_n9972));
  nand_5 g07624(.A(new_n9972), .B(pi065), .Y(new_n9973));
  xor_4  g07625(.A(new_n9972), .B(pi065), .Y(new_n9974));
  xor_4  g07626(.A(new_n9958), .B(new_n9956), .Y(new_n9975));
  nand_5 g07627(.A(new_n9975), .B(pi195), .Y(new_n9976));
  xor_4  g07628(.A(new_n9975), .B(pi195), .Y(new_n9977));
  not_8  g07629(.A(pi379), .Y(new_n9978));
  xor_4  g07630(.A(pi474), .B(new_n8163), .Y(new_n9979));
  or_6   g07631(.A(new_n9979), .B(new_n9978), .Y(new_n9980));
  xor_4  g07632(.A(new_n9979), .B(new_n9978), .Y(new_n9981));
  nor_5  g07633(.A(pi838), .B(pi149), .Y(new_n9982));
  nand_5 g07634(.A(pi838), .B(new_n2552), .Y(new_n9983));
  or_6   g07635(.A(pi838), .B(new_n2552), .Y(new_n9984));
  and_6  g07636(.A(new_n9984), .B(new_n9983), .Y(new_n9985));
  nor_5  g07637(.A(new_n9985), .B(pi677), .Y(new_n9986));
  nor_5  g07638(.A(new_n9986), .B(new_n9982), .Y(new_n9987));
  nand_5 g07639(.A(new_n9987), .B(new_n9981), .Y(new_n9988));
  nand_5 g07640(.A(new_n9988), .B(new_n9980), .Y(new_n9989));
  nand_5 g07641(.A(new_n9989), .B(new_n9977), .Y(new_n9990));
  nand_5 g07642(.A(new_n9990), .B(new_n9976), .Y(new_n9991));
  nand_5 g07643(.A(new_n9991), .B(new_n9974), .Y(new_n9992));
  nand_5 g07644(.A(new_n9992), .B(new_n9973), .Y(new_n9993));
  xor_4  g07645(.A(new_n9970), .B(new_n9969), .Y(new_n9994));
  nand_5 g07646(.A(new_n9994), .B(new_n9993), .Y(new_n9995));
  nand_5 g07647(.A(new_n9995), .B(new_n9971), .Y(new_n9996));
  xnor_4 g07648(.A(new_n9996), .B(new_n9968), .Y(new_n9997));
  xor_4  g07649(.A(new_n9946), .B(new_n9919), .Y(new_n9998));
  xor_4  g07650(.A(new_n9994), .B(new_n9993), .Y(new_n9999));
  nor_5  g07651(.A(new_n9999), .B(new_n9998), .Y(new_n10000));
  not_8  g07652(.A(new_n9998), .Y(new_n10001));
  xor_4  g07653(.A(new_n9999), .B(new_n10001), .Y(new_n10002));
  xor_4  g07654(.A(new_n9989), .B(new_n9977), .Y(new_n10003));
  xor_4  g07655(.A(new_n9987), .B(new_n9981), .Y(new_n10004));
  xor_4  g07656(.A(new_n9938), .B(new_n9929), .Y(new_n10005));
  nand_5 g07657(.A(new_n10005), .B(new_n10004), .Y(new_n10006));
  xor_4  g07658(.A(new_n9934), .B(pi702), .Y(new_n10007));
  not_8  g07659(.A(new_n10007), .Y(new_n10008));
  xor_4  g07660(.A(new_n9985), .B(new_n8166), .Y(new_n10009));
  or_6   g07661(.A(new_n10009), .B(new_n10008), .Y(new_n10010));
  xor_4  g07662(.A(new_n10005), .B(new_n10004), .Y(new_n10011));
  nand_5 g07663(.A(new_n10011), .B(new_n10010), .Y(new_n10012));
  nand_5 g07664(.A(new_n10012), .B(new_n10006), .Y(new_n10013));
  nor_5  g07665(.A(new_n10013), .B(new_n10003), .Y(new_n10014));
  xnor_4 g07666(.A(new_n10013), .B(new_n10003), .Y(new_n10015));
  xor_4  g07667(.A(new_n9941), .B(new_n9940), .Y(new_n10016));
  not_8  g07668(.A(new_n10016), .Y(new_n10017));
  nor_5  g07669(.A(new_n10017), .B(new_n10015), .Y(new_n10018));
  or_6   g07670(.A(new_n10018), .B(new_n10014), .Y(new_n10019));
  xnor_4 g07671(.A(new_n9991), .B(new_n9974), .Y(new_n10020));
  or_6   g07672(.A(new_n10020), .B(new_n10019), .Y(new_n10021));
  xor_4  g07673(.A(new_n10020), .B(new_n10019), .Y(new_n10022));
  xor_4  g07674(.A(new_n9944), .B(new_n9922), .Y(new_n10023));
  nand_5 g07675(.A(new_n10023), .B(new_n10022), .Y(new_n10024));
  nand_5 g07676(.A(new_n10024), .B(new_n10021), .Y(new_n10025));
  nor_5  g07677(.A(new_n10025), .B(new_n10002), .Y(new_n10026));
  or_6   g07678(.A(new_n10026), .B(new_n10000), .Y(new_n10027));
  or_6   g07679(.A(new_n10027), .B(new_n9997), .Y(new_n10028));
  xor_4  g07680(.A(new_n9948), .B(new_n9916), .Y(new_n10029));
  xor_4  g07681(.A(new_n10027), .B(new_n9997), .Y(new_n10030));
  nand_5 g07682(.A(new_n10030), .B(new_n10029), .Y(new_n10031));
  nand_5 g07683(.A(new_n10031), .B(new_n10028), .Y(new_n10032));
  nor_5  g07684(.A(new_n10032), .B(new_n9951), .Y(new_n10033));
  nand_5 g07685(.A(new_n9967), .B(pi222), .Y(new_n10034));
  nand_5 g07686(.A(new_n9996), .B(new_n9968), .Y(new_n10035));
  nand_5 g07687(.A(new_n10035), .B(new_n10034), .Y(new_n10036));
  xor_4  g07688(.A(pi798), .B(new_n8762), .Y(new_n10037));
  not_8  g07689(.A(new_n10037), .Y(new_n10038));
  not_8  g07690(.A(pi031), .Y(new_n10039));
  nand_5 g07691(.A(new_n8091), .B(new_n8153), .Y(new_n10040));
  nand_5 g07692(.A(new_n9966), .B(new_n9952), .Y(new_n10041));
  nand_5 g07693(.A(new_n10041), .B(new_n10040), .Y(new_n10042));
  nand_5 g07694(.A(new_n10042), .B(new_n10039), .Y(new_n10043));
  not_8  g07695(.A(new_n10043), .Y(new_n10044));
  nor_5  g07696(.A(new_n10042), .B(new_n10039), .Y(new_n10045));
  nor_5  g07697(.A(new_n10045), .B(new_n10044), .Y(new_n10046));
  xor_4  g07698(.A(new_n10046), .B(new_n10038), .Y(new_n10047));
  xor_4  g07699(.A(new_n10047), .B(new_n10036), .Y(new_n10048));
  not_8  g07700(.A(new_n9951), .Y(new_n10049));
  xor_4  g07701(.A(new_n10032), .B(new_n10049), .Y(new_n10050));
  nor_5  g07702(.A(new_n10050), .B(new_n10048), .Y(new_n10051));
  or_6   g07703(.A(new_n10051), .B(new_n10033), .Y(new_n10052));
  not_8  g07704(.A(new_n10047), .Y(new_n10053));
  nor_5  g07705(.A(new_n10053), .B(new_n10036), .Y(new_n10054));
  nor_5  g07706(.A(new_n10047), .B(pi798), .Y(new_n10055));
  nor_5  g07707(.A(new_n10055), .B(new_n10054), .Y(new_n10056));
  not_8  g07708(.A(pi705), .Y(new_n10057));
  nor_5  g07709(.A(new_n10045), .B(pi516), .Y(new_n10058));
  nor_5  g07710(.A(new_n10058), .B(new_n10044), .Y(new_n10059));
  nand_5 g07711(.A(pi310), .B(pi258), .Y(new_n10060));
  nand_5 g07712(.A(new_n8152), .B(new_n8055), .Y(new_n10061));
  nand_5 g07713(.A(new_n10061), .B(new_n10060), .Y(new_n10062));
  xor_4  g07714(.A(new_n10062), .B(new_n10059), .Y(new_n10063));
  nand_5 g07715(.A(new_n10063), .B(new_n10057), .Y(new_n10064));
  not_8  g07716(.A(new_n10064), .Y(new_n10065));
  nor_5  g07717(.A(new_n10063), .B(new_n10057), .Y(new_n10066));
  or_6   g07718(.A(new_n10066), .B(new_n10065), .Y(new_n10067));
  xor_4  g07719(.A(new_n10067), .B(new_n10056), .Y(new_n10068));
  nand_5 g07720(.A(new_n10068), .B(new_n10052), .Y(new_n10069));
  xnor_4 g07721(.A(new_n10068), .B(new_n10052), .Y(new_n10070));
  or_6   g07722(.A(new_n9912), .B(pi780), .Y(new_n10071));
  nand_5 g07723(.A(new_n9950), .B(new_n9913), .Y(new_n10072));
  nand_5 g07724(.A(new_n10072), .B(new_n10071), .Y(new_n10073));
  nand_5 g07725(.A(new_n8008), .B(new_n9888), .Y(new_n10074));
  or_6   g07726(.A(new_n9911), .B(new_n9889), .Y(new_n10075));
  nand_5 g07727(.A(new_n10075), .B(new_n10074), .Y(new_n10076));
  nand_5 g07728(.A(new_n10076), .B(new_n10073), .Y(new_n10077));
  not_8  g07729(.A(new_n10077), .Y(new_n10078));
  nor_5  g07730(.A(new_n10076), .B(new_n10073), .Y(new_n10079));
  nor_5  g07731(.A(new_n10079), .B(new_n10078), .Y(new_n10080));
  nor_5  g07732(.A(pi686), .B(new_n8004), .Y(new_n10081));
  not_8  g07733(.A(pi686), .Y(new_n10082));
  nor_5  g07734(.A(new_n10082), .B(pi336), .Y(new_n10083));
  nor_5  g07735(.A(new_n10083), .B(new_n10081), .Y(new_n10084));
  nor_5  g07736(.A(new_n10084), .B(pi503), .Y(new_n10085));
  nand_5 g07737(.A(new_n10084), .B(pi503), .Y(new_n10086));
  not_8  g07738(.A(new_n10086), .Y(new_n10087));
  nor_5  g07739(.A(new_n10087), .B(new_n10085), .Y(new_n10088));
  xor_4  g07740(.A(new_n10088), .B(new_n10080), .Y(new_n10089));
  or_6   g07741(.A(new_n10089), .B(new_n10070), .Y(new_n10090));
  nand_5 g07742(.A(new_n10090), .B(new_n10069), .Y(new_n10091));
  not_8  g07743(.A(pi665), .Y(new_n10092));
  nand_5 g07744(.A(pi810), .B(new_n10092), .Y(new_n10093));
  nand_5 g07745(.A(new_n8798), .B(pi665), .Y(new_n10094));
  nand_5 g07746(.A(new_n10094), .B(new_n10093), .Y(new_n10095));
  xor_4  g07747(.A(new_n10095), .B(new_n8277), .Y(new_n10096));
  not_8  g07748(.A(new_n10061), .Y(new_n10097));
  not_8  g07749(.A(new_n10060), .Y(new_n10098));
  nor_5  g07750(.A(new_n10098), .B(new_n10059), .Y(new_n10099));
  nor_5  g07751(.A(new_n10099), .B(new_n10097), .Y(new_n10100));
  not_8  g07752(.A(new_n10100), .Y(new_n10101));
  nand_5 g07753(.A(new_n10101), .B(new_n10096), .Y(new_n10102));
  or_6   g07754(.A(new_n10101), .B(new_n10096), .Y(new_n10103));
  nand_5 g07755(.A(new_n10103), .B(new_n10102), .Y(new_n10104));
  nor_5  g07756(.A(new_n10066), .B(new_n10056), .Y(new_n10105));
  nor_5  g07757(.A(new_n10105), .B(new_n10065), .Y(new_n10106));
  xnor_4 g07758(.A(new_n10106), .B(new_n10104), .Y(new_n10107));
  not_8  g07759(.A(new_n10107), .Y(new_n10108));
  nand_5 g07760(.A(new_n10108), .B(new_n10091), .Y(new_n10109));
  not_8  g07761(.A(new_n10109), .Y(new_n10110));
  nor_5  g07762(.A(new_n10108), .B(new_n10091), .Y(new_n10111));
  xor_4  g07763(.A(pi722), .B(pi278), .Y(new_n10112));
  xor_4  g07764(.A(new_n10112), .B(pi748), .Y(new_n10113));
  not_8  g07765(.A(new_n10079), .Y(new_n10114));
  nand_5 g07766(.A(new_n10082), .B(new_n8004), .Y(new_n10115));
  not_8  g07767(.A(new_n10115), .Y(new_n10116));
  nor_5  g07768(.A(new_n10116), .B(new_n10085), .Y(new_n10117));
  nor_5  g07769(.A(new_n10115), .B(pi503), .Y(new_n10118));
  nor_5  g07770(.A(new_n10118), .B(new_n10078), .Y(new_n10119));
  nor_5  g07771(.A(new_n10119), .B(new_n10117), .Y(new_n10120));
  nand_5 g07772(.A(new_n10120), .B(new_n10114), .Y(new_n10121));
  nand_5 g07773(.A(new_n10087), .B(pi336), .Y(new_n10122));
  nor_5  g07774(.A(new_n10122), .B(new_n10078), .Y(new_n10123));
  not_8  g07775(.A(new_n10123), .Y(new_n10124));
  nand_5 g07776(.A(new_n10124), .B(new_n10121), .Y(new_n10125));
  nand_5 g07777(.A(new_n10125), .B(new_n10113), .Y(new_n10126));
  xor_4  g07778(.A(new_n10117), .B(new_n10113), .Y(new_n10127));
  nor_5  g07779(.A(new_n10127), .B(new_n10114), .Y(new_n10128));
  nor_5  g07780(.A(new_n10113), .B(new_n10079), .Y(new_n10129));
  nand_5 g07781(.A(new_n10129), .B(new_n10124), .Y(new_n10130));
  nor_5  g07782(.A(new_n10130), .B(new_n10120), .Y(new_n10131));
  nor_5  g07783(.A(new_n10131), .B(new_n10128), .Y(new_n10132));
  nand_5 g07784(.A(new_n10132), .B(new_n10126), .Y(new_n10133));
  not_8  g07785(.A(new_n10133), .Y(new_n10134));
  nor_5  g07786(.A(new_n10134), .B(new_n10111), .Y(new_n10135));
  nor_5  g07787(.A(new_n10135), .B(new_n10110), .Y(new_n10136));
  nand_5 g07788(.A(pi700), .B(pi079), .Y(new_n10137));
  not_8  g07789(.A(pi079), .Y(new_n10138));
  nand_5 g07790(.A(new_n8052), .B(new_n10138), .Y(new_n10139));
  nand_5 g07791(.A(new_n10139), .B(new_n10137), .Y(new_n10140));
  not_8  g07792(.A(new_n10140), .Y(new_n10141));
  not_8  g07793(.A(new_n10102), .Y(new_n10142));
  nand_5 g07794(.A(new_n10092), .B(new_n8277), .Y(new_n10143));
  nand_5 g07795(.A(pi665), .B(pi586), .Y(new_n10144));
  nand_5 g07796(.A(new_n10144), .B(new_n8798), .Y(new_n10145));
  nand_5 g07797(.A(new_n10145), .B(new_n10143), .Y(new_n10146));
  nor_5  g07798(.A(new_n10146), .B(new_n10142), .Y(new_n10147));
  nand_5 g07799(.A(new_n10147), .B(new_n10106), .Y(new_n10148));
  nor_5  g07800(.A(new_n10144), .B(new_n8798), .Y(new_n10149));
  nand_5 g07801(.A(new_n10149), .B(new_n10100), .Y(new_n10150));
  nand_5 g07802(.A(new_n10150), .B(new_n10148), .Y(new_n10151));
  not_8  g07803(.A(new_n10151), .Y(new_n10152));
  nand_5 g07804(.A(new_n10146), .B(new_n10103), .Y(new_n10153));
  nor_5  g07805(.A(new_n10153), .B(new_n10106), .Y(new_n10154));
  nor_5  g07806(.A(new_n10143), .B(pi810), .Y(new_n10155));
  nand_5 g07807(.A(new_n10155), .B(new_n10101), .Y(new_n10156));
  not_8  g07808(.A(new_n10156), .Y(new_n10157));
  nor_5  g07809(.A(new_n10157), .B(new_n10154), .Y(new_n10158));
  nand_5 g07810(.A(new_n10158), .B(new_n10152), .Y(new_n10159));
  xor_4  g07811(.A(new_n10159), .B(pi041), .Y(new_n10160));
  xor_4  g07812(.A(new_n10160), .B(new_n10141), .Y(new_n10161));
  not_8  g07813(.A(new_n10161), .Y(new_n10162));
  nand_5 g07814(.A(new_n10162), .B(new_n10136), .Y(new_n10163));
  xor_4  g07815(.A(new_n10161), .B(new_n10136), .Y(new_n10164));
  not_8  g07816(.A(pi431), .Y(new_n10165));
  not_8  g07817(.A(pi465), .Y(new_n10166));
  nand_5 g07818(.A(new_n10166), .B(new_n10165), .Y(new_n10167));
  nand_5 g07819(.A(pi465), .B(pi431), .Y(new_n10168));
  nand_5 g07820(.A(new_n10168), .B(new_n10167), .Y(new_n10169));
  xor_4  g07821(.A(new_n10169), .B(pi542), .Y(new_n10170));
  or_6   g07822(.A(pi722), .B(pi278), .Y(new_n10171));
  nand_5 g07823(.A(new_n10112), .B(new_n8117), .Y(new_n10172));
  nand_5 g07824(.A(new_n10172), .B(new_n10171), .Y(new_n10173));
  or_6   g07825(.A(new_n10117), .B(new_n10113), .Y(new_n10174));
  nand_5 g07826(.A(new_n10174), .B(new_n10121), .Y(new_n10175));
  or_6   g07827(.A(new_n10175), .B(new_n10131), .Y(new_n10176));
  nor_5  g07828(.A(new_n10176), .B(new_n10173), .Y(new_n10177));
  nand_5 g07829(.A(new_n10176), .B(new_n10173), .Y(new_n10178));
  not_8  g07830(.A(new_n10178), .Y(new_n10179));
  nor_5  g07831(.A(new_n10179), .B(new_n10177), .Y(new_n10180));
  xor_4  g07832(.A(new_n10180), .B(new_n10170), .Y(new_n10181));
  not_8  g07833(.A(new_n10181), .Y(new_n10182));
  or_6   g07834(.A(new_n10182), .B(new_n10164), .Y(new_n10183));
  nand_5 g07835(.A(new_n10183), .B(new_n10163), .Y(new_n10184));
  or_6   g07836(.A(new_n10152), .B(new_n10137), .Y(new_n10185));
  not_8  g07837(.A(new_n10185), .Y(new_n10186));
  nand_5 g07838(.A(new_n10152), .B(new_n10137), .Y(new_n10187));
  not_8  g07839(.A(new_n10187), .Y(new_n10188));
  nand_5 g07840(.A(new_n10139), .B(pi041), .Y(new_n10189));
  not_8  g07841(.A(new_n10189), .Y(new_n10190));
  nand_5 g07842(.A(new_n10190), .B(new_n10158), .Y(new_n10191));
  nor_5  g07843(.A(new_n10191), .B(new_n10188), .Y(new_n10192));
  nor_5  g07844(.A(new_n10192), .B(new_n10186), .Y(new_n10193));
  nor_5  g07845(.A(new_n10139), .B(pi041), .Y(new_n10194));
  nand_5 g07846(.A(new_n10194), .B(new_n10152), .Y(new_n10195));
  not_8  g07847(.A(new_n10195), .Y(new_n10196));
  nand_5 g07848(.A(new_n10189), .B(new_n10137), .Y(new_n10197));
  nor_5  g07849(.A(new_n10197), .B(new_n10158), .Y(new_n10198));
  nor_5  g07850(.A(new_n10198), .B(new_n10196), .Y(new_n10199));
  nand_5 g07851(.A(new_n10199), .B(new_n10193), .Y(new_n10200));
  not_8  g07852(.A(new_n10200), .Y(new_n10201));
  nor_5  g07853(.A(new_n10201), .B(new_n10184), .Y(new_n10202));
  xor_4  g07854(.A(new_n10200), .B(new_n10184), .Y(new_n10203));
  nand_5 g07855(.A(new_n10182), .B(new_n4327), .Y(new_n10204));
  not_8  g07856(.A(new_n10204), .Y(new_n10205));
  nand_5 g07857(.A(new_n10177), .B(new_n10167), .Y(new_n10206));
  not_8  g07858(.A(new_n10206), .Y(new_n10207));
  nor_5  g07859(.A(new_n10179), .B(new_n10168), .Y(new_n10208));
  nor_5  g07860(.A(new_n10208), .B(new_n10207), .Y(new_n10209));
  nor_5  g07861(.A(new_n10209), .B(new_n10205), .Y(new_n10210));
  not_8  g07862(.A(new_n10210), .Y(new_n10211));
  not_8  g07863(.A(new_n10167), .Y(new_n10212));
  nand_5 g07864(.A(new_n10212), .B(new_n4327), .Y(new_n10213));
  nor_5  g07865(.A(new_n10213), .B(new_n10177), .Y(new_n10214));
  nor_5  g07866(.A(new_n10169), .B(pi542), .Y(new_n10215));
  nor_5  g07867(.A(new_n10215), .B(new_n10212), .Y(new_n10216));
  nor_5  g07868(.A(new_n10216), .B(new_n10178), .Y(new_n10217));
  nor_5  g07869(.A(new_n10217), .B(new_n10214), .Y(new_n10218));
  nand_5 g07870(.A(new_n10218), .B(new_n10211), .Y(new_n10219));
  nor_5  g07871(.A(new_n10219), .B(new_n10203), .Y(new_n10220));
  or_6   g07872(.A(new_n10220), .B(new_n10202), .Y(new_n10221));
  xor_4  g07873(.A(new_n10210), .B(new_n10193), .Y(new_n10222));
  xnor_4 g07874(.A(new_n10222), .B(new_n10221), .Y(po0060));
  xor_4  g07875(.A(pi443), .B(new_n8981), .Y(new_n10224));
  nor_5  g07876(.A(pi701), .B(new_n8796), .Y(new_n10225));
  xor_4  g07877(.A(pi701), .B(new_n8796), .Y(new_n10226));
  not_8  g07878(.A(new_n10226), .Y(new_n10227));
  nor_5  g07879(.A(pi279), .B(new_n8759), .Y(new_n10228));
  not_8  g07880(.A(pi811), .Y(new_n10229));
  nand_5 g07881(.A(new_n10229), .B(pi786), .Y(new_n10230));
  xor_4  g07882(.A(new_n10229), .B(pi786), .Y(new_n10231));
  nand_5 g07883(.A(new_n8767), .B(pi187), .Y(new_n10232));
  not_8  g07884(.A(pi187), .Y(new_n10233));
  xor_4  g07885(.A(pi804), .B(new_n10233), .Y(new_n10234));
  nand_5 g07886(.A(pi720), .B(new_n8770), .Y(new_n10235));
  xor_4  g07887(.A(pi720), .B(new_n8770), .Y(new_n10236));
  nand_5 g07888(.A(pi339), .B(new_n8773), .Y(new_n10237));
  xor_4  g07889(.A(pi339), .B(new_n8773), .Y(new_n10238));
  not_8  g07890(.A(pi576), .Y(new_n10239));
  nand_5 g07891(.A(new_n10239), .B(pi521), .Y(new_n10240));
  xor_4  g07892(.A(pi576), .B(new_n2705), .Y(new_n10241));
  nand_5 g07893(.A(new_n8778), .B(pi370), .Y(new_n10242));
  not_8  g07894(.A(pi370), .Y(new_n10243));
  xor_4  g07895(.A(pi401), .B(new_n10243), .Y(new_n10244));
  nand_5 g07896(.A(pi544), .B(new_n8835), .Y(new_n10245));
  not_8  g07897(.A(new_n10245), .Y(new_n10246));
  nand_5 g07898(.A(new_n10246), .B(new_n10244), .Y(new_n10247));
  nand_5 g07899(.A(new_n10247), .B(new_n10242), .Y(new_n10248));
  nand_5 g07900(.A(new_n10248), .B(new_n10241), .Y(new_n10249));
  nand_5 g07901(.A(new_n10249), .B(new_n10240), .Y(new_n10250));
  nand_5 g07902(.A(new_n10250), .B(new_n10238), .Y(new_n10251));
  nand_5 g07903(.A(new_n10251), .B(new_n10237), .Y(new_n10252));
  nand_5 g07904(.A(new_n10252), .B(new_n10236), .Y(new_n10253));
  nand_5 g07905(.A(new_n10253), .B(new_n10235), .Y(new_n10254));
  nand_5 g07906(.A(new_n10254), .B(new_n10234), .Y(new_n10255));
  nand_5 g07907(.A(new_n10255), .B(new_n10232), .Y(new_n10256));
  nand_5 g07908(.A(new_n10256), .B(new_n10231), .Y(new_n10257));
  nand_5 g07909(.A(new_n10257), .B(new_n10230), .Y(new_n10258));
  xor_4  g07910(.A(pi279), .B(pi123), .Y(new_n10259));
  nor_5  g07911(.A(new_n10259), .B(new_n10258), .Y(new_n10260));
  nor_5  g07912(.A(new_n10260), .B(new_n10228), .Y(new_n10261));
  nor_5  g07913(.A(new_n10261), .B(new_n10227), .Y(new_n10262));
  nor_5  g07914(.A(new_n10262), .B(new_n10225), .Y(new_n10263));
  xor_4  g07915(.A(new_n10263), .B(new_n10224), .Y(new_n10264));
  xor_4  g07916(.A(pi403), .B(pi358), .Y(new_n10265));
  not_8  g07917(.A(pi687), .Y(new_n10266));
  nand_5 g07918(.A(new_n10266), .B(new_n9174), .Y(new_n10267));
  xor_4  g07919(.A(pi687), .B(pi334), .Y(new_n10268));
  nand_5 g07920(.A(new_n5501), .B(new_n2855), .Y(new_n10269));
  xor_4  g07921(.A(pi342), .B(pi047), .Y(new_n10270));
  nand_5 g07922(.A(new_n5505), .B(new_n2859), .Y(new_n10271));
  nand_5 g07923(.A(new_n9541), .B(new_n9538), .Y(new_n10272));
  nand_5 g07924(.A(new_n10272), .B(new_n10271), .Y(new_n10273));
  nand_5 g07925(.A(new_n10273), .B(new_n10270), .Y(new_n10274));
  nand_5 g07926(.A(new_n10274), .B(new_n10269), .Y(new_n10275));
  nand_5 g07927(.A(new_n10275), .B(new_n10268), .Y(new_n10276));
  nand_5 g07928(.A(new_n10276), .B(new_n10267), .Y(new_n10277));
  xor_4  g07929(.A(new_n10277), .B(new_n10265), .Y(new_n10278));
  not_8  g07930(.A(new_n2820), .Y(new_n10279));
  xor_4  g07931(.A(new_n10273), .B(new_n10270), .Y(new_n10280));
  not_8  g07932(.A(new_n10280), .Y(new_n10281));
  nand_5 g07933(.A(new_n10281), .B(new_n2738), .Y(new_n10282));
  xor_4  g07934(.A(new_n10280), .B(new_n2737), .Y(new_n10283));
  not_8  g07935(.A(new_n9427), .Y(new_n10284));
  nand_5 g07936(.A(new_n9447), .B(new_n2750), .Y(new_n10285));
  not_8  g07937(.A(new_n10285), .Y(new_n10286));
  nand_5 g07938(.A(new_n10286), .B(new_n2684), .Y(new_n10287));
  nand_5 g07939(.A(new_n10285), .B(new_n2706), .Y(new_n10288));
  and_6  g07940(.A(new_n10288), .B(new_n10287), .Y(new_n10289));
  nand_5 g07941(.A(new_n10289), .B(new_n9413), .Y(new_n10290));
  nand_5 g07942(.A(new_n10290), .B(new_n10287), .Y(new_n10291));
  or_6   g07943(.A(new_n10291), .B(new_n10284), .Y(new_n10292));
  xor_4  g07944(.A(new_n10291), .B(new_n10284), .Y(new_n10293));
  nand_5 g07945(.A(new_n10293), .B(new_n2712), .Y(new_n10294));
  nand_5 g07946(.A(new_n10294), .B(new_n10292), .Y(new_n10295));
  or_6   g07947(.A(new_n10295), .B(new_n9440), .Y(new_n10296));
  not_8  g07948(.A(new_n2716), .Y(new_n10297));
  xor_4  g07949(.A(new_n10295), .B(new_n9440), .Y(new_n10298));
  nand_5 g07950(.A(new_n10298), .B(new_n10297), .Y(new_n10299));
  nand_5 g07951(.A(new_n10299), .B(new_n10296), .Y(new_n10300));
  or_6   g07952(.A(new_n10300), .B(new_n2702), .Y(new_n10301));
  xor_4  g07953(.A(new_n10300), .B(new_n2702), .Y(new_n10302));
  nand_5 g07954(.A(new_n10302), .B(new_n9491), .Y(new_n10303));
  nand_5 g07955(.A(new_n10303), .B(new_n10301), .Y(new_n10304));
  nor_5  g07956(.A(new_n10304), .B(new_n2699), .Y(new_n10305));
  xor_4  g07957(.A(new_n10304), .B(new_n2699), .Y(new_n10306));
  not_8  g07958(.A(new_n10306), .Y(new_n10307));
  nor_5  g07959(.A(new_n10307), .B(new_n9530), .Y(new_n10308));
  or_6   g07960(.A(new_n10308), .B(new_n10305), .Y(new_n10309));
  nand_5 g07961(.A(new_n10309), .B(new_n9542), .Y(new_n10310));
  not_8  g07962(.A(new_n9542), .Y(new_n10311));
  xor_4  g07963(.A(new_n10309), .B(new_n10311), .Y(new_n10312));
  or_6   g07964(.A(new_n10312), .B(new_n2696), .Y(new_n10313));
  nand_5 g07965(.A(new_n10313), .B(new_n10310), .Y(new_n10314));
  not_8  g07966(.A(new_n10314), .Y(new_n10315));
  nand_5 g07967(.A(new_n10315), .B(new_n10283), .Y(new_n10316));
  nand_5 g07968(.A(new_n10316), .B(new_n10282), .Y(new_n10317));
  or_6   g07969(.A(new_n10317), .B(new_n10279), .Y(new_n10318));
  xor_4  g07970(.A(new_n10275), .B(new_n10268), .Y(new_n10319));
  xor_4  g07971(.A(new_n10317), .B(new_n10279), .Y(new_n10320));
  nand_5 g07972(.A(new_n10320), .B(new_n10319), .Y(new_n10321));
  nand_5 g07973(.A(new_n10321), .B(new_n10318), .Y(new_n10322));
  xor_4  g07974(.A(new_n10322), .B(new_n10278), .Y(new_n10323));
  xor_4  g07975(.A(new_n10323), .B(new_n2847), .Y(new_n10324));
  not_8  g07976(.A(new_n10324), .Y(new_n10325));
  or_6   g07977(.A(new_n10325), .B(new_n10264), .Y(new_n10326));
  xor_4  g07978(.A(new_n10325), .B(new_n10264), .Y(new_n10327));
  xor_4  g07979(.A(new_n10261), .B(new_n10226), .Y(new_n10328));
  xor_4  g07980(.A(new_n10320), .B(new_n10319), .Y(new_n10329));
  or_6   g07981(.A(new_n10329), .B(new_n10328), .Y(new_n10330));
  xor_4  g07982(.A(new_n10329), .B(new_n10328), .Y(new_n10331));
  xor_4  g07983(.A(new_n10259), .B(new_n10258), .Y(new_n10332));
  xor_4  g07984(.A(new_n10314), .B(new_n10283), .Y(new_n10333));
  not_8  g07985(.A(new_n10333), .Y(new_n10334));
  nor_5  g07986(.A(new_n10334), .B(new_n10332), .Y(new_n10335));
  nand_5 g07987(.A(new_n10334), .B(new_n10332), .Y(new_n10336));
  xor_4  g07988(.A(new_n10256), .B(new_n10231), .Y(new_n10337));
  not_8  g07989(.A(new_n10337), .Y(new_n10338));
  xor_4  g07990(.A(new_n10312), .B(new_n2697), .Y(new_n10339));
  nor_5  g07991(.A(new_n10339), .B(new_n10338), .Y(new_n10340));
  xor_4  g07992(.A(new_n10339), .B(new_n10337), .Y(new_n10341));
  xor_4  g07993(.A(new_n10307), .B(new_n9530), .Y(new_n10342));
  xor_4  g07994(.A(new_n10252), .B(new_n10236), .Y(new_n10343));
  xor_4  g07995(.A(new_n10302), .B(new_n9490), .Y(new_n10344));
  nand_5 g07996(.A(new_n10344), .B(new_n10343), .Y(new_n10345));
  xnor_4 g07997(.A(new_n10344), .B(new_n10343), .Y(new_n10346));
  xor_4  g07998(.A(new_n10250), .B(new_n10238), .Y(new_n10347));
  not_8  g07999(.A(new_n10347), .Y(new_n10348));
  xor_4  g08000(.A(new_n10298), .B(new_n2716), .Y(new_n10349));
  nor_5  g08001(.A(new_n10349), .B(new_n10348), .Y(new_n10350));
  xor_4  g08002(.A(new_n10349), .B(new_n10347), .Y(new_n10351));
  xor_4  g08003(.A(new_n10248), .B(new_n10241), .Y(new_n10352));
  not_8  g08004(.A(new_n10352), .Y(new_n10353));
  xor_4  g08005(.A(new_n10293), .B(new_n2712), .Y(new_n10354));
  nand_5 g08006(.A(new_n10354), .B(new_n10353), .Y(new_n10355));
  or_6   g08007(.A(new_n10354), .B(new_n10353), .Y(new_n10356));
  xor_4  g08008(.A(new_n10289), .B(new_n9414), .Y(new_n10357));
  not_8  g08009(.A(new_n10357), .Y(new_n10358));
  xor_4  g08010(.A(new_n9416), .B(new_n2748), .Y(new_n10359));
  nand_5 g08011(.A(new_n10359), .B(new_n10358), .Y(new_n10360));
  not_8  g08012(.A(new_n10360), .Y(new_n10361));
  or_6   g08013(.A(new_n10361), .B(new_n10247), .Y(new_n10362));
  not_8  g08014(.A(new_n10359), .Y(new_n10363));
  nor_5  g08015(.A(pi544), .B(new_n8835), .Y(new_n10364));
  nand_5 g08016(.A(new_n10364), .B(new_n10363), .Y(new_n10365));
  nand_5 g08017(.A(new_n10359), .B(new_n10246), .Y(new_n10366));
  nand_5 g08018(.A(new_n10366), .B(new_n10365), .Y(new_n10367));
  xor_4  g08019(.A(new_n10367), .B(new_n10244), .Y(new_n10368));
  nor_5  g08020(.A(new_n10368), .B(new_n10358), .Y(new_n10369));
  nor_5  g08021(.A(new_n10365), .B(new_n10244), .Y(new_n10370));
  nor_5  g08022(.A(new_n10370), .B(new_n10369), .Y(new_n10371));
  nand_5 g08023(.A(new_n10371), .B(new_n10362), .Y(new_n10372));
  nand_5 g08024(.A(new_n10372), .B(new_n10356), .Y(new_n10373));
  nand_5 g08025(.A(new_n10373), .B(new_n10355), .Y(new_n10374));
  nor_5  g08026(.A(new_n10374), .B(new_n10351), .Y(new_n10375));
  nor_5  g08027(.A(new_n10375), .B(new_n10350), .Y(new_n10376));
  or_6   g08028(.A(new_n10376), .B(new_n10346), .Y(new_n10377));
  nand_5 g08029(.A(new_n10377), .B(new_n10345), .Y(new_n10378));
  nand_5 g08030(.A(new_n10378), .B(new_n10342), .Y(new_n10379));
  xor_4  g08031(.A(new_n10254), .B(new_n10234), .Y(new_n10380));
  xor_4  g08032(.A(new_n10378), .B(new_n10342), .Y(new_n10381));
  nand_5 g08033(.A(new_n10381), .B(new_n10380), .Y(new_n10382));
  and_6  g08034(.A(new_n10382), .B(new_n10379), .Y(new_n10383));
  nor_5  g08035(.A(new_n10383), .B(new_n10341), .Y(new_n10384));
  or_6   g08036(.A(new_n10384), .B(new_n10340), .Y(new_n10385));
  and_6  g08037(.A(new_n10385), .B(new_n10336), .Y(new_n10386));
  nor_5  g08038(.A(new_n10386), .B(new_n10335), .Y(new_n10387));
  nand_5 g08039(.A(new_n10387), .B(new_n10331), .Y(new_n10388));
  nand_5 g08040(.A(new_n10388), .B(new_n10330), .Y(new_n10389));
  nand_5 g08041(.A(new_n10389), .B(new_n10327), .Y(new_n10390));
  nand_5 g08042(.A(new_n10390), .B(new_n10326), .Y(new_n10391));
  nand_5 g08043(.A(new_n2846), .B(pi397), .Y(new_n10392));
  not_8  g08044(.A(new_n10263), .Y(new_n10393));
  nand_5 g08045(.A(new_n10393), .B(new_n10224), .Y(new_n10394));
  nand_5 g08046(.A(new_n10394), .B(new_n10392), .Y(new_n10395));
  nand_5 g08047(.A(new_n10395), .B(new_n10391), .Y(new_n10396));
  not_8  g08048(.A(new_n10396), .Y(new_n10397));
  nor_5  g08049(.A(new_n10395), .B(new_n10391), .Y(new_n10398));
  nor_5  g08050(.A(new_n10398), .B(new_n10397), .Y(new_n10399));
  not_8  g08051(.A(pi358), .Y(new_n10400));
  nand_5 g08052(.A(new_n5545), .B(new_n10400), .Y(new_n10401));
  nand_5 g08053(.A(new_n10277), .B(new_n10265), .Y(new_n10402));
  nand_5 g08054(.A(new_n10402), .B(new_n10401), .Y(new_n10403));
  not_8  g08055(.A(new_n10403), .Y(new_n10404));
  not_8  g08056(.A(pi095), .Y(new_n10405));
  nand_5 g08057(.A(new_n4329), .B(new_n10405), .Y(new_n10406));
  not_8  g08058(.A(new_n10406), .Y(new_n10407));
  not_8  g08059(.A(new_n2836), .Y(new_n10408));
  nor_5  g08060(.A(new_n2843), .B(new_n10408), .Y(new_n10409));
  nor_5  g08061(.A(new_n10409), .B(new_n10407), .Y(new_n10410));
  not_8  g08062(.A(new_n10410), .Y(new_n10411));
  nand_5 g08063(.A(new_n10411), .B(new_n10404), .Y(new_n10412));
  nand_5 g08064(.A(new_n10322), .B(new_n10278), .Y(new_n10413));
  nand_5 g08065(.A(new_n10323), .B(new_n2844), .Y(new_n10414));
  nand_5 g08066(.A(new_n10414), .B(new_n10413), .Y(new_n10415));
  or_6   g08067(.A(new_n10415), .B(new_n10412), .Y(new_n10416));
  nand_5 g08068(.A(new_n10410), .B(new_n10403), .Y(new_n10417));
  nand_5 g08069(.A(new_n10415), .B(new_n10412), .Y(new_n10418));
  nand_5 g08070(.A(new_n10418), .B(new_n10417), .Y(new_n10419));
  not_8  g08071(.A(new_n10419), .Y(new_n10420));
  nand_5 g08072(.A(new_n10420), .B(new_n10416), .Y(new_n10421));
  not_8  g08073(.A(new_n10415), .Y(new_n10422));
  nor_5  g08074(.A(new_n10417), .B(new_n10422), .Y(new_n10423));
  not_8  g08075(.A(new_n10423), .Y(new_n10424));
  nand_5 g08076(.A(new_n10424), .B(new_n10421), .Y(new_n10425));
  xor_4  g08077(.A(new_n10425), .B(new_n10399), .Y(po0061));
  not_8  g08078(.A(pi461), .Y(new_n10427));
  not_8  g08079(.A(new_n5555), .Y(new_n10428));
  not_8  g08080(.A(new_n5560), .Y(new_n10429));
  nand_5 g08081(.A(new_n10429), .B(pi137), .Y(new_n10430));
  xor_4  g08082(.A(new_n10429), .B(pi137), .Y(new_n10431));
  not_8  g08083(.A(new_n5565), .Y(new_n10432));
  not_8  g08084(.A(new_n5573), .Y(new_n10433));
  not_8  g08085(.A(new_n5577), .Y(new_n10434));
  nand_5 g08086(.A(new_n10434), .B(pi562), .Y(new_n10435));
  xor_4  g08087(.A(new_n10434), .B(pi562), .Y(new_n10436));
  nand_5 g08088(.A(new_n5802), .B(new_n5801), .Y(new_n10437));
  nand_5 g08089(.A(new_n5803), .B(new_n5607), .Y(new_n10438));
  nand_5 g08090(.A(new_n10438), .B(new_n10437), .Y(new_n10439));
  or_6   g08091(.A(new_n10439), .B(new_n5588), .Y(new_n10440));
  nand_5 g08092(.A(new_n10439), .B(new_n5588), .Y(new_n10441));
  nand_5 g08093(.A(new_n10441), .B(pi416), .Y(new_n10442));
  nand_5 g08094(.A(new_n10442), .B(new_n10440), .Y(new_n10443));
  nand_5 g08095(.A(new_n10443), .B(pi387), .Y(new_n10444));
  xnor_4 g08096(.A(new_n10443), .B(pi387), .Y(new_n10445));
  or_6   g08097(.A(new_n10445), .B(new_n5583), .Y(new_n10446));
  nand_5 g08098(.A(new_n10446), .B(new_n10444), .Y(new_n10447));
  nand_5 g08099(.A(new_n10447), .B(new_n10436), .Y(new_n10448));
  nand_5 g08100(.A(new_n10448), .B(new_n10435), .Y(new_n10449));
  or_6   g08101(.A(new_n10449), .B(new_n10433), .Y(new_n10450));
  nand_5 g08102(.A(new_n10450), .B(pi357), .Y(new_n10451));
  nand_5 g08103(.A(new_n10449), .B(new_n10433), .Y(new_n10452));
  and_6  g08104(.A(new_n10452), .B(new_n10451), .Y(new_n10453));
  nand_5 g08105(.A(new_n10453), .B(new_n5569), .Y(new_n10454));
  nand_5 g08106(.A(new_n10454), .B(pi489), .Y(new_n10455));
  or_6   g08107(.A(new_n10453), .B(new_n5569), .Y(new_n10456));
  nand_5 g08108(.A(new_n10456), .B(new_n10455), .Y(new_n10457));
  nand_5 g08109(.A(new_n10457), .B(new_n10432), .Y(new_n10458));
  not_8  g08110(.A(pi668), .Y(new_n10459));
  xor_4  g08111(.A(new_n10457), .B(new_n5565), .Y(new_n10460));
  or_6   g08112(.A(new_n10460), .B(new_n10459), .Y(new_n10461));
  nand_5 g08113(.A(new_n10461), .B(new_n10458), .Y(new_n10462));
  nand_5 g08114(.A(new_n10462), .B(new_n10431), .Y(new_n10463));
  nand_5 g08115(.A(new_n10463), .B(new_n10430), .Y(new_n10464));
  nor_5  g08116(.A(new_n10464), .B(new_n10428), .Y(new_n10465));
  nor_5  g08117(.A(new_n10465), .B(new_n10427), .Y(new_n10466));
  and_6  g08118(.A(new_n10464), .B(new_n10428), .Y(new_n10467));
  nor_5  g08119(.A(new_n10467), .B(new_n10466), .Y(new_n10468));
  nor_5  g08120(.A(new_n10468), .B(new_n5496), .Y(new_n10469));
  not_8  g08121(.A(pi533), .Y(new_n10470));
  xor_4  g08122(.A(pi789), .B(new_n10470), .Y(new_n10471));
  nand_5 g08123(.A(new_n5642), .B(pi249), .Y(new_n10472));
  xor_4  g08124(.A(pi377), .B(new_n6259), .Y(new_n10473));
  nand_5 g08125(.A(new_n6829), .B(pi707), .Y(new_n10474));
  xor_4  g08126(.A(pi714), .B(new_n6221), .Y(new_n10475));
  nand_5 g08127(.A(new_n5648), .B(pi433), .Y(new_n10476));
  not_8  g08128(.A(pi433), .Y(new_n10477));
  xor_4  g08129(.A(pi539), .B(new_n10477), .Y(new_n10478));
  nand_5 g08130(.A(pi568), .B(new_n5651), .Y(new_n10479));
  xor_4  g08131(.A(pi568), .B(new_n5651), .Y(new_n10480));
  nand_5 g08132(.A(new_n5654), .B(pi183), .Y(new_n10481));
  xor_4  g08133(.A(pi252), .B(new_n4005), .Y(new_n10482));
  nand_5 g08134(.A(new_n6836), .B(pi176), .Y(new_n10483));
  xor_4  g08135(.A(pi391), .B(new_n3933), .Y(new_n10484));
  nand_5 g08136(.A(new_n6651), .B(pi245), .Y(new_n10485));
  nand_5 g08137(.A(new_n5798), .B(new_n5797), .Y(new_n10486));
  nand_5 g08138(.A(new_n10486), .B(new_n10485), .Y(new_n10487));
  nand_5 g08139(.A(new_n10487), .B(new_n10484), .Y(new_n10488));
  nand_5 g08140(.A(new_n10488), .B(new_n10483), .Y(new_n10489));
  nand_5 g08141(.A(new_n10489), .B(new_n10482), .Y(new_n10490));
  nand_5 g08142(.A(new_n10490), .B(new_n10481), .Y(new_n10491));
  nand_5 g08143(.A(new_n10491), .B(new_n10480), .Y(new_n10492));
  nand_5 g08144(.A(new_n10492), .B(new_n10479), .Y(new_n10493));
  nand_5 g08145(.A(new_n10493), .B(new_n10478), .Y(new_n10494));
  nand_5 g08146(.A(new_n10494), .B(new_n10476), .Y(new_n10495));
  nand_5 g08147(.A(new_n10495), .B(new_n10475), .Y(new_n10496));
  nand_5 g08148(.A(new_n10496), .B(new_n10474), .Y(new_n10497));
  nand_5 g08149(.A(new_n10497), .B(new_n10473), .Y(new_n10498));
  nand_5 g08150(.A(new_n10498), .B(new_n10472), .Y(new_n10499));
  xor_4  g08151(.A(new_n10499), .B(new_n10471), .Y(new_n10500));
  not_8  g08152(.A(new_n10500), .Y(new_n10501));
  xor_4  g08153(.A(new_n10497), .B(new_n10473), .Y(new_n10502));
  not_8  g08154(.A(new_n10502), .Y(new_n10503));
  xor_4  g08155(.A(new_n10495), .B(new_n10475), .Y(new_n10504));
  not_8  g08156(.A(new_n10504), .Y(new_n10505));
  xor_4  g08157(.A(new_n10493), .B(new_n10478), .Y(new_n10506));
  not_8  g08158(.A(new_n10506), .Y(new_n10507));
  xor_4  g08159(.A(new_n10491), .B(new_n10480), .Y(new_n10508));
  not_8  g08160(.A(new_n10508), .Y(new_n10509));
  xor_4  g08161(.A(new_n10489), .B(new_n10482), .Y(new_n10510));
  xor_4  g08162(.A(new_n10487), .B(new_n10484), .Y(new_n10511));
  nand_5 g08163(.A(new_n5799), .B(pi528), .Y(new_n10512));
  nand_5 g08164(.A(new_n5800), .B(new_n5793), .Y(new_n10513));
  nand_5 g08165(.A(new_n10513), .B(new_n10512), .Y(new_n10514));
  nand_5 g08166(.A(new_n10514), .B(new_n10511), .Y(new_n10515));
  xor_4  g08167(.A(new_n10514), .B(new_n10511), .Y(new_n10516));
  nand_5 g08168(.A(new_n10516), .B(pi362), .Y(new_n10517));
  nand_5 g08169(.A(new_n10517), .B(new_n10515), .Y(new_n10518));
  nor_5  g08170(.A(new_n10518), .B(new_n10510), .Y(new_n10519));
  not_8  g08171(.A(new_n10510), .Y(new_n10520));
  xor_4  g08172(.A(new_n10518), .B(new_n10520), .Y(new_n10521));
  nor_5  g08173(.A(new_n10521), .B(pi338), .Y(new_n10522));
  or_6   g08174(.A(new_n10522), .B(new_n10519), .Y(new_n10523));
  nand_5 g08175(.A(new_n10523), .B(new_n10509), .Y(new_n10524));
  xor_4  g08176(.A(new_n10523), .B(new_n10508), .Y(new_n10525));
  or_6   g08177(.A(new_n10525), .B(pi250), .Y(new_n10526));
  nand_5 g08178(.A(new_n10526), .B(new_n10524), .Y(new_n10527));
  nand_5 g08179(.A(new_n10527), .B(new_n10507), .Y(new_n10528));
  xor_4  g08180(.A(new_n10527), .B(new_n10506), .Y(new_n10529));
  or_6   g08181(.A(new_n10529), .B(pi613), .Y(new_n10530));
  nand_5 g08182(.A(new_n10530), .B(new_n10528), .Y(new_n10531));
  nand_5 g08183(.A(new_n10531), .B(new_n10505), .Y(new_n10532));
  xor_4  g08184(.A(new_n10531), .B(new_n10504), .Y(new_n10533));
  or_6   g08185(.A(new_n10533), .B(pi297), .Y(new_n10534));
  nand_5 g08186(.A(new_n10534), .B(new_n10532), .Y(new_n10535));
  nand_5 g08187(.A(new_n10535), .B(new_n10503), .Y(new_n10536));
  xor_4  g08188(.A(new_n10535), .B(new_n10502), .Y(new_n10537));
  or_6   g08189(.A(new_n10537), .B(pi834), .Y(new_n10538));
  nand_5 g08190(.A(new_n10538), .B(new_n10536), .Y(new_n10539));
  nand_5 g08191(.A(new_n10539), .B(new_n10501), .Y(new_n10540));
  xor_4  g08192(.A(new_n10539), .B(new_n10500), .Y(new_n10541));
  or_6   g08193(.A(new_n10541), .B(pi472), .Y(new_n10542));
  nand_5 g08194(.A(new_n10542), .B(new_n10540), .Y(new_n10543));
  nor_5  g08195(.A(new_n10543), .B(new_n5634), .Y(new_n10544));
  xor_4  g08196(.A(new_n10543), .B(new_n5634), .Y(new_n10545));
  not_8  g08197(.A(new_n10545), .Y(new_n10546));
  xor_4  g08198(.A(pi735), .B(new_n6380), .Y(new_n10547));
  nand_5 g08199(.A(pi789), .B(new_n10470), .Y(new_n10548));
  nand_5 g08200(.A(new_n10499), .B(new_n10471), .Y(new_n10549));
  nand_5 g08201(.A(new_n10549), .B(new_n10548), .Y(new_n10550));
  xnor_4 g08202(.A(new_n10550), .B(new_n10547), .Y(new_n10551));
  nor_5  g08203(.A(new_n10551), .B(new_n10546), .Y(new_n10552));
  nor_5  g08204(.A(new_n10552), .B(new_n10544), .Y(new_n10553));
  not_8  g08205(.A(pi735), .Y(new_n10554));
  nand_5 g08206(.A(new_n10554), .B(pi490), .Y(new_n10555));
  nand_5 g08207(.A(new_n10550), .B(new_n10547), .Y(new_n10556));
  nand_5 g08208(.A(new_n10556), .B(new_n10555), .Y(new_n10557));
  or_6   g08209(.A(new_n10557), .B(new_n10553), .Y(new_n10558));
  and_6  g08210(.A(new_n10558), .B(new_n10469), .Y(new_n10559));
  nor_5  g08211(.A(new_n10558), .B(new_n10469), .Y(new_n10560));
  nor_5  g08212(.A(new_n10560), .B(new_n10559), .Y(new_n10561));
  xor_4  g08213(.A(new_n10468), .B(new_n5496), .Y(new_n10562));
  not_8  g08214(.A(new_n10557), .Y(new_n10563));
  xor_4  g08215(.A(new_n10563), .B(new_n10553), .Y(new_n10564));
  nand_5 g08216(.A(new_n10564), .B(new_n10562), .Y(new_n10565));
  not_8  g08217(.A(new_n10565), .Y(new_n10566));
  or_6   g08218(.A(new_n10467), .B(new_n10465), .Y(new_n10567));
  xor_4  g08219(.A(new_n10567), .B(new_n10427), .Y(new_n10568));
  xor_4  g08220(.A(new_n10551), .B(new_n10545), .Y(new_n10569));
  nor_5  g08221(.A(new_n10569), .B(new_n10568), .Y(new_n10570));
  not_8  g08222(.A(new_n10568), .Y(new_n10571));
  xor_4  g08223(.A(new_n10569), .B(new_n10571), .Y(new_n10572));
  xor_4  g08224(.A(new_n10462), .B(new_n10431), .Y(new_n10573));
  not_8  g08225(.A(new_n10573), .Y(new_n10574));
  xor_4  g08226(.A(new_n10541), .B(new_n5636), .Y(new_n10575));
  and_6  g08227(.A(new_n10575), .B(new_n10574), .Y(new_n10576));
  xor_4  g08228(.A(new_n10537), .B(new_n5640), .Y(new_n10577));
  xor_4  g08229(.A(new_n10460), .B(pi668), .Y(new_n10578));
  nor_5  g08230(.A(new_n10578), .B(new_n10577), .Y(new_n10579));
  xnor_4 g08231(.A(new_n10578), .B(new_n10577), .Y(new_n10580));
  xor_4  g08232(.A(new_n10533), .B(new_n5644), .Y(new_n10581));
  nand_5 g08233(.A(new_n10456), .B(new_n10454), .Y(new_n10582));
  xor_4  g08234(.A(new_n10582), .B(pi489), .Y(new_n10583));
  nand_5 g08235(.A(new_n10583), .B(new_n10581), .Y(new_n10584));
  xnor_4 g08236(.A(new_n10583), .B(new_n10581), .Y(new_n10585));
  xor_4  g08237(.A(new_n10529), .B(new_n5646), .Y(new_n10586));
  nand_5 g08238(.A(new_n10452), .B(new_n10450), .Y(new_n10587));
  xor_4  g08239(.A(new_n10587), .B(pi357), .Y(new_n10588));
  and_6  g08240(.A(new_n10588), .B(new_n10586), .Y(new_n10589));
  xnor_4 g08241(.A(new_n10588), .B(new_n10586), .Y(new_n10590));
  xor_4  g08242(.A(new_n10447), .B(new_n10436), .Y(new_n10591));
  not_8  g08243(.A(new_n10591), .Y(new_n10592));
  xor_4  g08244(.A(new_n10525), .B(new_n3991), .Y(new_n10593));
  nor_5  g08245(.A(new_n10593), .B(new_n10592), .Y(new_n10594));
  xor_4  g08246(.A(new_n10521), .B(new_n3993), .Y(new_n10595));
  xor_4  g08247(.A(new_n10445), .B(new_n5582), .Y(new_n10596));
  nand_5 g08248(.A(new_n10596), .B(new_n10595), .Y(new_n10597));
  nand_5 g08249(.A(new_n10441), .B(new_n10440), .Y(new_n10598));
  xor_4  g08250(.A(new_n10598), .B(pi416), .Y(new_n10599));
  not_8  g08251(.A(new_n10599), .Y(new_n10600));
  xor_4  g08252(.A(new_n10516), .B(new_n3946), .Y(new_n10601));
  nand_5 g08253(.A(new_n10601), .B(new_n10600), .Y(new_n10602));
  xor_4  g08254(.A(new_n10601), .B(new_n10600), .Y(new_n10603));
  nand_5 g08255(.A(new_n5804), .B(new_n5800), .Y(new_n10604));
  nor_5  g08256(.A(new_n5792), .B(new_n5787), .Y(new_n10605));
  nor_5  g08257(.A(new_n10605), .B(new_n10604), .Y(new_n10606));
  nor_5  g08258(.A(new_n5805), .B(new_n5795), .Y(new_n10607));
  nand_5 g08259(.A(new_n10513), .B(new_n5791), .Y(new_n10608));
  nor_5  g08260(.A(new_n10608), .B(new_n10607), .Y(new_n10609));
  nor_5  g08261(.A(new_n10609), .B(new_n10606), .Y(new_n10610));
  nand_5 g08262(.A(new_n10610), .B(new_n10603), .Y(new_n10611));
  nand_5 g08263(.A(new_n10611), .B(new_n10602), .Y(new_n10612));
  xnor_4 g08264(.A(new_n10596), .B(new_n10595), .Y(new_n10613));
  or_6   g08265(.A(new_n10613), .B(new_n10612), .Y(new_n10614));
  nand_5 g08266(.A(new_n10614), .B(new_n10597), .Y(new_n10615));
  xor_4  g08267(.A(new_n10593), .B(new_n10591), .Y(new_n10616));
  nor_5  g08268(.A(new_n10616), .B(new_n10615), .Y(new_n10617));
  or_6   g08269(.A(new_n10617), .B(new_n10594), .Y(new_n10618));
  nor_5  g08270(.A(new_n10618), .B(new_n10590), .Y(new_n10619));
  nor_5  g08271(.A(new_n10619), .B(new_n10589), .Y(new_n10620));
  or_6   g08272(.A(new_n10620), .B(new_n10585), .Y(new_n10621));
  nand_5 g08273(.A(new_n10621), .B(new_n10584), .Y(new_n10622));
  nor_5  g08274(.A(new_n10622), .B(new_n10580), .Y(new_n10623));
  or_6   g08275(.A(new_n10623), .B(new_n10579), .Y(new_n10624));
  xor_4  g08276(.A(new_n10575), .B(new_n10573), .Y(new_n10625));
  nor_5  g08277(.A(new_n10625), .B(new_n10624), .Y(new_n10626));
  nor_5  g08278(.A(new_n10626), .B(new_n10576), .Y(new_n10627));
  nor_5  g08279(.A(new_n10627), .B(new_n10572), .Y(new_n10628));
  or_6   g08280(.A(new_n10628), .B(new_n10570), .Y(new_n10629));
  not_8  g08281(.A(new_n10562), .Y(new_n10630));
  xor_4  g08282(.A(new_n10564), .B(new_n10630), .Y(new_n10631));
  nor_5  g08283(.A(new_n10631), .B(new_n10629), .Y(new_n10632));
  nor_5  g08284(.A(new_n10632), .B(new_n10566), .Y(new_n10633));
  xor_4  g08285(.A(new_n10633), .B(new_n10561), .Y(po0062));
  nand_5 g08286(.A(new_n8082), .B(new_n7270), .Y(new_n10635));
  nand_5 g08287(.A(new_n8536), .B(new_n8535), .Y(new_n10636));
  nand_5 g08288(.A(new_n10636), .B(new_n10635), .Y(new_n10637));
  or_6   g08289(.A(new_n10637), .B(new_n8061), .Y(new_n10638));
  nand_5 g08290(.A(new_n10637), .B(new_n8061), .Y(new_n10639));
  nand_5 g08291(.A(new_n10639), .B(pi635), .Y(new_n10640));
  nand_5 g08292(.A(new_n10640), .B(new_n10638), .Y(new_n10641));
  nand_5 g08293(.A(new_n10641), .B(new_n8059), .Y(new_n10642));
  xor_4  g08294(.A(new_n10641), .B(new_n8059), .Y(new_n10643));
  nand_5 g08295(.A(new_n10643), .B(pi265), .Y(new_n10644));
  nand_5 g08296(.A(new_n10644), .B(new_n10642), .Y(new_n10645));
  or_6   g08297(.A(new_n10645), .B(new_n8058), .Y(new_n10646));
  not_8  g08298(.A(pi332), .Y(new_n10647));
  xor_4  g08299(.A(new_n10645), .B(new_n8058), .Y(new_n10648));
  nand_5 g08300(.A(new_n10648), .B(new_n10647), .Y(new_n10649));
  nand_5 g08301(.A(new_n10649), .B(new_n10646), .Y(new_n10650));
  xor_4  g08302(.A(new_n10650), .B(new_n8103), .Y(new_n10651));
  xor_4  g08303(.A(new_n10651), .B(pi772), .Y(new_n10652));
  xor_4  g08304(.A(new_n10648), .B(new_n10647), .Y(new_n10653));
  xor_4  g08305(.A(new_n10643), .B(pi265), .Y(new_n10654));
  not_8  g08306(.A(pi604), .Y(new_n10655));
  xor_4  g08307(.A(pi201), .B(pi104), .Y(new_n10656));
  nand_5 g08308(.A(pi795), .B(pi343), .Y(new_n10657));
  nand_5 g08309(.A(new_n6639), .B(new_n6635), .Y(new_n10658));
  nand_5 g08310(.A(new_n10658), .B(new_n10657), .Y(new_n10659));
  xor_4  g08311(.A(new_n10659), .B(new_n10656), .Y(new_n10660));
  nand_5 g08312(.A(new_n8543), .B(new_n4130), .Y(new_n10661));
  nand_5 g08313(.A(new_n10661), .B(new_n8542), .Y(new_n10662));
  not_8  g08314(.A(new_n10662), .Y(new_n10663));
  or_6   g08315(.A(new_n10663), .B(new_n10660), .Y(new_n10664));
  nand_5 g08316(.A(new_n10663), .B(new_n10660), .Y(new_n10665));
  nand_5 g08317(.A(new_n10665), .B(new_n10664), .Y(new_n10666));
  xor_4  g08318(.A(new_n10666), .B(new_n10655), .Y(new_n10667));
  nand_5 g08319(.A(new_n10639), .B(new_n10638), .Y(new_n10668));
  xor_4  g08320(.A(new_n10668), .B(pi635), .Y(new_n10669));
  nor_5  g08321(.A(new_n10669), .B(new_n10667), .Y(new_n10670));
  xnor_4 g08322(.A(new_n10669), .B(new_n10667), .Y(new_n10671));
  not_8  g08323(.A(new_n8537), .Y(new_n10672));
  nor_5  g08324(.A(new_n10672), .B(new_n8532), .Y(new_n10673));
  nor_5  g08325(.A(new_n8545), .B(new_n8538), .Y(new_n10674));
  or_6   g08326(.A(new_n10674), .B(new_n10673), .Y(new_n10675));
  nor_5  g08327(.A(new_n10675), .B(new_n10671), .Y(new_n10676));
  or_6   g08328(.A(new_n10676), .B(new_n10670), .Y(new_n10677));
  nor_5  g08329(.A(new_n10677), .B(new_n10654), .Y(new_n10678));
  xnor_4 g08330(.A(new_n10677), .B(new_n10654), .Y(new_n10679));
  xor_4  g08331(.A(pi641), .B(pi363), .Y(new_n10680));
  nand_5 g08332(.A(pi201), .B(pi104), .Y(new_n10681));
  nand_5 g08333(.A(new_n10659), .B(new_n10656), .Y(new_n10682));
  nand_5 g08334(.A(new_n10682), .B(new_n10681), .Y(new_n10683));
  xor_4  g08335(.A(new_n10683), .B(new_n10680), .Y(new_n10684));
  nand_5 g08336(.A(new_n10665), .B(new_n10655), .Y(new_n10685));
  nand_5 g08337(.A(new_n10685), .B(new_n10664), .Y(new_n10686));
  not_8  g08338(.A(new_n10686), .Y(new_n10687));
  or_6   g08339(.A(new_n10687), .B(new_n10684), .Y(new_n10688));
  nand_5 g08340(.A(new_n10687), .B(new_n10684), .Y(new_n10689));
  nand_5 g08341(.A(new_n10689), .B(new_n10688), .Y(new_n10690));
  xor_4  g08342(.A(new_n10690), .B(pi814), .Y(new_n10691));
  nor_5  g08343(.A(new_n10691), .B(new_n10679), .Y(new_n10692));
  or_6   g08344(.A(new_n10692), .B(new_n10678), .Y(new_n10693));
  nand_5 g08345(.A(new_n10693), .B(new_n10653), .Y(new_n10694));
  xnor_4 g08346(.A(new_n10693), .B(new_n10653), .Y(new_n10695));
  xor_4  g08347(.A(pi451), .B(pi064), .Y(new_n10696));
  nand_5 g08348(.A(pi641), .B(pi363), .Y(new_n10697));
  nand_5 g08349(.A(new_n10683), .B(new_n10680), .Y(new_n10698));
  nand_5 g08350(.A(new_n10698), .B(new_n10697), .Y(new_n10699));
  xor_4  g08351(.A(new_n10699), .B(new_n10696), .Y(new_n10700));
  not_8  g08352(.A(pi814), .Y(new_n10701));
  nand_5 g08353(.A(new_n10689), .B(new_n10701), .Y(new_n10702));
  nand_5 g08354(.A(new_n10702), .B(new_n10688), .Y(new_n10703));
  not_8  g08355(.A(new_n10703), .Y(new_n10704));
  or_6   g08356(.A(new_n10704), .B(new_n10700), .Y(new_n10705));
  nand_5 g08357(.A(new_n10704), .B(new_n10700), .Y(new_n10706));
  nand_5 g08358(.A(new_n10706), .B(new_n10705), .Y(new_n10707));
  xor_4  g08359(.A(new_n10707), .B(pi484), .Y(new_n10708));
  or_6   g08360(.A(new_n10708), .B(new_n10695), .Y(new_n10709));
  nand_5 g08361(.A(new_n10709), .B(new_n10694), .Y(new_n10710));
  not_8  g08362(.A(pi164), .Y(new_n10711));
  xor_4  g08363(.A(pi203), .B(pi021), .Y(new_n10712));
  nand_5 g08364(.A(pi451), .B(pi064), .Y(new_n10713));
  nand_5 g08365(.A(new_n10699), .B(new_n10696), .Y(new_n10714));
  nand_5 g08366(.A(new_n10714), .B(new_n10713), .Y(new_n10715));
  xnor_4 g08367(.A(new_n10715), .B(new_n10712), .Y(new_n10716));
  xor_4  g08368(.A(new_n10716), .B(new_n10711), .Y(new_n10717));
  not_8  g08369(.A(pi484), .Y(new_n10718));
  nand_5 g08370(.A(new_n10706), .B(new_n10718), .Y(new_n10719));
  nand_5 g08371(.A(new_n10719), .B(new_n10705), .Y(new_n10720));
  xor_4  g08372(.A(new_n10720), .B(new_n10717), .Y(new_n10721));
  xor_4  g08373(.A(new_n10721), .B(new_n10710), .Y(new_n10722));
  xnor_4 g08374(.A(new_n10722), .B(new_n10652), .Y(po0063));
  xor_4  g08375(.A(pi439), .B(new_n2943), .Y(new_n10724));
  and_6  g08376(.A(pi822), .B(new_n4341), .Y(new_n10725));
  nor_5  g08377(.A(pi822), .B(new_n4341), .Y(new_n10726));
  nor_5  g08378(.A(pi263), .B(new_n7758), .Y(new_n10727));
  nor_5  g08379(.A(new_n2966), .B(pi100), .Y(new_n10728));
  not_8  g08380(.A(pi117), .Y(new_n10729));
  nor_5  g08381(.A(pi766), .B(new_n10729), .Y(new_n10730));
  nor_5  g08382(.A(new_n9602), .B(new_n9599), .Y(new_n10731));
  nor_5  g08383(.A(new_n10731), .B(new_n10730), .Y(new_n10732));
  nor_5  g08384(.A(new_n10732), .B(new_n10728), .Y(new_n10733));
  nor_5  g08385(.A(new_n10733), .B(new_n10727), .Y(new_n10734));
  nor_5  g08386(.A(new_n10734), .B(new_n10726), .Y(new_n10735));
  nor_5  g08387(.A(new_n10735), .B(new_n10725), .Y(new_n10736));
  xor_4  g08388(.A(new_n10736), .B(new_n10724), .Y(new_n10737));
  xor_4  g08389(.A(pi530), .B(new_n4382), .Y(new_n10738));
  nand_5 g08390(.A(new_n9512), .B(pi248), .Y(new_n10739));
  not_8  g08391(.A(pi248), .Y(new_n10740));
  xor_4  g08392(.A(pi712), .B(new_n10740), .Y(new_n10741));
  not_8  g08393(.A(pi511), .Y(new_n10742));
  nand_5 g08394(.A(new_n10742), .B(pi125), .Y(new_n10743));
  not_8  g08395(.A(pi125), .Y(new_n10744));
  xor_4  g08396(.A(pi511), .B(new_n10744), .Y(new_n10745));
  nand_5 g08397(.A(pi618), .B(new_n6579), .Y(new_n10746));
  xor_4  g08398(.A(pi618), .B(new_n6579), .Y(new_n10747));
  nand_5 g08399(.A(new_n7720), .B(pi192), .Y(new_n10748));
  xor_4  g08400(.A(pi475), .B(new_n8018), .Y(new_n10749));
  nand_5 g08401(.A(pi813), .B(new_n5768), .Y(new_n10750));
  nand_5 g08402(.A(new_n5769), .B(new_n5767), .Y(new_n10751));
  nand_5 g08403(.A(new_n10751), .B(new_n10750), .Y(new_n10752));
  nand_5 g08404(.A(new_n10752), .B(new_n10749), .Y(new_n10753));
  nand_5 g08405(.A(new_n10753), .B(new_n10748), .Y(new_n10754));
  nand_5 g08406(.A(new_n10754), .B(new_n10747), .Y(new_n10755));
  nand_5 g08407(.A(new_n10755), .B(new_n10746), .Y(new_n10756));
  nand_5 g08408(.A(new_n10756), .B(new_n10745), .Y(new_n10757));
  nand_5 g08409(.A(new_n10757), .B(new_n10743), .Y(new_n10758));
  nand_5 g08410(.A(new_n10758), .B(new_n10741), .Y(new_n10759));
  nand_5 g08411(.A(new_n10759), .B(new_n10739), .Y(new_n10760));
  xor_4  g08412(.A(new_n10760), .B(new_n10738), .Y(new_n10761));
  xor_4  g08413(.A(new_n10761), .B(new_n10737), .Y(new_n10762));
  nor_5  g08414(.A(new_n10726), .B(new_n10725), .Y(new_n10763));
  xor_4  g08415(.A(new_n10763), .B(new_n10734), .Y(new_n10764));
  xor_4  g08416(.A(new_n10758), .B(new_n10741), .Y(new_n10765));
  nand_5 g08417(.A(new_n10765), .B(new_n10764), .Y(new_n10766));
  xor_4  g08418(.A(new_n10756), .B(new_n10745), .Y(new_n10767));
  xor_4  g08419(.A(new_n10752), .B(new_n10749), .Y(new_n10768));
  not_8  g08420(.A(new_n5770), .Y(new_n10769));
  nor_5  g08421(.A(new_n10769), .B(new_n5764), .Y(new_n10770));
  nor_5  g08422(.A(new_n5771), .B(new_n5761), .Y(new_n10771));
  or_6   g08423(.A(new_n10771), .B(new_n10770), .Y(new_n10772));
  nor_5  g08424(.A(new_n10772), .B(new_n10768), .Y(new_n10773));
  not_8  g08425(.A(new_n10768), .Y(new_n10774));
  xor_4  g08426(.A(new_n10772), .B(new_n10774), .Y(new_n10775));
  nor_5  g08427(.A(new_n10775), .B(new_n9587), .Y(new_n10776));
  or_6   g08428(.A(new_n10776), .B(new_n10773), .Y(new_n10777));
  nor_5  g08429(.A(new_n10754), .B(new_n10747), .Y(new_n10778));
  not_8  g08430(.A(new_n10778), .Y(new_n10779));
  nand_5 g08431(.A(new_n10779), .B(new_n10755), .Y(new_n10780));
  nor_5  g08432(.A(new_n10780), .B(new_n10777), .Y(new_n10781));
  not_8  g08433(.A(new_n10780), .Y(new_n10782));
  xor_4  g08434(.A(new_n10782), .B(new_n10777), .Y(new_n10783));
  nor_5  g08435(.A(new_n10783), .B(new_n9603), .Y(new_n10784));
  or_6   g08436(.A(new_n10784), .B(new_n10781), .Y(new_n10785));
  nand_5 g08437(.A(new_n10785), .B(new_n10767), .Y(new_n10786));
  not_8  g08438(.A(new_n10786), .Y(new_n10787));
  nor_5  g08439(.A(new_n10728), .B(new_n10727), .Y(new_n10788));
  xor_4  g08440(.A(new_n10788), .B(new_n10732), .Y(new_n10789));
  not_8  g08441(.A(new_n10789), .Y(new_n10790));
  not_8  g08442(.A(new_n10767), .Y(new_n10791));
  xor_4  g08443(.A(new_n10785), .B(new_n10791), .Y(new_n10792));
  nor_5  g08444(.A(new_n10792), .B(new_n10790), .Y(new_n10793));
  nor_5  g08445(.A(new_n10793), .B(new_n10787), .Y(new_n10794));
  not_8  g08446(.A(new_n10765), .Y(new_n10795));
  xor_4  g08447(.A(new_n10795), .B(new_n10764), .Y(new_n10796));
  or_6   g08448(.A(new_n10796), .B(new_n10794), .Y(new_n10797));
  nand_5 g08449(.A(new_n10797), .B(new_n10766), .Y(new_n10798));
  xor_4  g08450(.A(new_n10798), .B(new_n10762), .Y(new_n10799));
  xor_4  g08451(.A(new_n10792), .B(new_n10789), .Y(new_n10800));
  nand_5 g08452(.A(new_n10800), .B(new_n10434), .Y(new_n10801));
  xor_4  g08453(.A(new_n10783), .B(new_n9603), .Y(new_n10802));
  xor_4  g08454(.A(new_n10775), .B(new_n9619), .Y(new_n10803));
  nand_5 g08455(.A(new_n10803), .B(new_n5588), .Y(new_n10804));
  xor_4  g08456(.A(new_n10803), .B(new_n5587), .Y(new_n10805));
  nand_5 g08457(.A(new_n5774), .B(new_n5606), .Y(new_n10806));
  or_6   g08458(.A(new_n5776), .B(new_n5772), .Y(new_n10807));
  nand_5 g08459(.A(new_n10807), .B(new_n10806), .Y(new_n10808));
  or_6   g08460(.A(new_n10808), .B(new_n10805), .Y(new_n10809));
  nand_5 g08461(.A(new_n10809), .B(new_n10804), .Y(new_n10810));
  or_6   g08462(.A(new_n10810), .B(new_n10802), .Y(new_n10811));
  xor_4  g08463(.A(new_n10810), .B(new_n10802), .Y(new_n10812));
  nand_5 g08464(.A(new_n10812), .B(new_n5582), .Y(new_n10813));
  nand_5 g08465(.A(new_n10813), .B(new_n10811), .Y(new_n10814));
  xor_4  g08466(.A(new_n10800), .B(new_n10434), .Y(new_n10815));
  nand_5 g08467(.A(new_n10815), .B(new_n10814), .Y(new_n10816));
  nand_5 g08468(.A(new_n10816), .B(new_n10801), .Y(new_n10817));
  nor_5  g08469(.A(new_n10817), .B(new_n10433), .Y(new_n10818));
  not_8  g08470(.A(new_n10796), .Y(new_n10819));
  xor_4  g08471(.A(new_n10819), .B(new_n10794), .Y(new_n10820));
  xor_4  g08472(.A(new_n10817), .B(new_n5573), .Y(new_n10821));
  nor_5  g08473(.A(new_n10821), .B(new_n10820), .Y(new_n10822));
  or_6   g08474(.A(new_n10822), .B(new_n10818), .Y(new_n10823));
  xnor_4 g08475(.A(new_n10823), .B(new_n10799), .Y(new_n10824));
  xor_4  g08476(.A(new_n10824), .B(new_n5569), .Y(po0064));
  xor_4  g08477(.A(pi484), .B(pi462), .Y(new_n10826));
  nand_5 g08478(.A(new_n10701), .B(new_n9322), .Y(new_n10827));
  xor_4  g08479(.A(pi814), .B(pi099), .Y(new_n10828));
  nand_5 g08480(.A(new_n10655), .B(new_n9285), .Y(new_n10829));
  nand_5 g08481(.A(new_n4130), .B(new_n9280), .Y(new_n10830));
  not_8  g08482(.A(new_n10830), .Y(new_n10831));
  xor_4  g08483(.A(pi524), .B(pi087), .Y(new_n10832));
  not_8  g08484(.A(new_n10832), .Y(new_n10833));
  nand_5 g08485(.A(new_n4133), .B(new_n9261), .Y(new_n10834));
  not_8  g08486(.A(new_n10834), .Y(new_n10835));
  xor_4  g08487(.A(pi460), .B(pi048), .Y(new_n10836));
  not_8  g08488(.A(new_n10836), .Y(new_n10837));
  not_8  g08489(.A(pi235), .Y(new_n10838));
  nand_5 g08490(.A(new_n10838), .B(new_n4139), .Y(new_n10839));
  not_8  g08491(.A(new_n10839), .Y(new_n10840));
  nand_5 g08492(.A(pi828), .B(pi758), .Y(new_n10841));
  not_8  g08493(.A(new_n10841), .Y(new_n10842));
  xor_4  g08494(.A(pi235), .B(new_n4139), .Y(new_n10843));
  nor_5  g08495(.A(new_n10843), .B(new_n10842), .Y(new_n10844));
  nor_5  g08496(.A(new_n10844), .B(new_n10840), .Y(new_n10845));
  nor_5  g08497(.A(new_n10845), .B(new_n10837), .Y(new_n10846));
  nor_5  g08498(.A(new_n10846), .B(new_n10835), .Y(new_n10847));
  nor_5  g08499(.A(new_n10847), .B(new_n10833), .Y(new_n10848));
  nor_5  g08500(.A(new_n10848), .B(new_n10831), .Y(new_n10849));
  xor_4  g08501(.A(pi604), .B(new_n9285), .Y(new_n10850));
  or_6   g08502(.A(new_n10850), .B(new_n10849), .Y(new_n10851));
  nand_5 g08503(.A(new_n10851), .B(new_n10829), .Y(new_n10852));
  nand_5 g08504(.A(new_n10852), .B(new_n10828), .Y(new_n10853));
  nand_5 g08505(.A(new_n10853), .B(new_n10827), .Y(new_n10854));
  xor_4  g08506(.A(new_n10854), .B(new_n10826), .Y(new_n10855));
  not_8  g08507(.A(new_n10855), .Y(new_n10856));
  xor_4  g08508(.A(new_n10850), .B(new_n10849), .Y(new_n10857));
  xor_4  g08509(.A(new_n10845), .B(new_n10836), .Y(new_n10858));
  not_8  g08510(.A(new_n10858), .Y(new_n10859));
  nand_5 g08511(.A(new_n10859), .B(new_n8073), .Y(new_n10860));
  xor_4  g08512(.A(pi828), .B(pi758), .Y(new_n10861));
  nand_5 g08513(.A(new_n10861), .B(new_n8064), .Y(new_n10862));
  xor_4  g08514(.A(new_n10843), .B(new_n10842), .Y(new_n10863));
  nand_5 g08515(.A(new_n10863), .B(new_n10862), .Y(new_n10864));
  or_6   g08516(.A(new_n10862), .B(new_n10843), .Y(new_n10865));
  nand_5 g08517(.A(new_n10865), .B(new_n10864), .Y(new_n10866));
  or_6   g08518(.A(new_n10866), .B(new_n8069), .Y(new_n10867));
  nand_5 g08519(.A(new_n10867), .B(new_n10864), .Y(new_n10868));
  xor_4  g08520(.A(new_n10858), .B(new_n8072), .Y(new_n10869));
  nand_5 g08521(.A(new_n10869), .B(new_n10868), .Y(new_n10870));
  nand_5 g08522(.A(new_n10870), .B(new_n10860), .Y(new_n10871));
  xor_4  g08523(.A(new_n10847), .B(new_n10832), .Y(new_n10872));
  not_8  g08524(.A(new_n10872), .Y(new_n10873));
  nand_5 g08525(.A(new_n10873), .B(new_n10871), .Y(new_n10874));
  xor_4  g08526(.A(new_n10873), .B(new_n10871), .Y(new_n10875));
  nand_5 g08527(.A(new_n10875), .B(new_n8081), .Y(new_n10876));
  nand_5 g08528(.A(new_n10876), .B(new_n10874), .Y(new_n10877));
  or_6   g08529(.A(new_n10877), .B(new_n10857), .Y(new_n10878));
  xor_4  g08530(.A(new_n10877), .B(new_n10857), .Y(new_n10879));
  nand_5 g08531(.A(new_n10879), .B(new_n8061), .Y(new_n10880));
  nand_5 g08532(.A(new_n10880), .B(new_n10878), .Y(new_n10881));
  xor_4  g08533(.A(new_n10852), .B(new_n10828), .Y(new_n10882));
  not_8  g08534(.A(new_n10882), .Y(new_n10883));
  nand_5 g08535(.A(new_n10883), .B(new_n10881), .Y(new_n10884));
  xor_4  g08536(.A(new_n10883), .B(new_n10881), .Y(new_n10885));
  not_8  g08537(.A(new_n10885), .Y(new_n10886));
  or_6   g08538(.A(new_n10886), .B(new_n8059), .Y(new_n10887));
  nand_5 g08539(.A(new_n10887), .B(new_n10884), .Y(new_n10888));
  nand_5 g08540(.A(new_n10888), .B(new_n10856), .Y(new_n10889));
  xor_4  g08541(.A(new_n10888), .B(new_n10856), .Y(new_n10890));
  nand_5 g08542(.A(new_n10890), .B(new_n8057), .Y(new_n10891));
  nand_5 g08543(.A(new_n10891), .B(new_n10889), .Y(new_n10892));
  xor_4  g08544(.A(pi442), .B(pi164), .Y(new_n10893));
  nand_5 g08545(.A(new_n10718), .B(new_n9294), .Y(new_n10894));
  nand_5 g08546(.A(new_n10854), .B(new_n10826), .Y(new_n10895));
  nand_5 g08547(.A(new_n10895), .B(new_n10894), .Y(new_n10896));
  xor_4  g08548(.A(new_n10896), .B(new_n10893), .Y(new_n10897));
  not_8  g08549(.A(new_n10897), .Y(new_n10898));
  nor_5  g08550(.A(new_n10898), .B(new_n10892), .Y(new_n10899));
  xor_4  g08551(.A(new_n10897), .B(new_n10892), .Y(new_n10900));
  nor_5  g08552(.A(new_n10900), .B(new_n8103), .Y(new_n10901));
  or_6   g08553(.A(new_n10901), .B(new_n10899), .Y(new_n10902));
  xor_4  g08554(.A(pi541), .B(pi108), .Y(new_n10903));
  or_6   g08555(.A(pi442), .B(pi164), .Y(new_n10904));
  nand_5 g08556(.A(new_n10896), .B(new_n10893), .Y(new_n10905));
  nand_5 g08557(.A(new_n10905), .B(new_n10904), .Y(new_n10906));
  xor_4  g08558(.A(new_n10906), .B(new_n10903), .Y(new_n10907));
  xor_4  g08559(.A(new_n10907), .B(new_n10902), .Y(new_n10908));
  xor_4  g08560(.A(new_n10908), .B(new_n8054), .Y(new_n10909));
  nand_5 g08561(.A(new_n10909), .B(new_n9306), .Y(new_n10910));
  not_8  g08562(.A(new_n10910), .Y(new_n10911));
  xor_4  g08563(.A(new_n10909), .B(new_n9311), .Y(new_n10912));
  not_8  g08564(.A(new_n9298), .Y(new_n10913));
  xor_4  g08565(.A(new_n10900), .B(new_n8224), .Y(new_n10914));
  nand_5 g08566(.A(new_n10914), .B(new_n10913), .Y(new_n10915));
  xor_4  g08567(.A(new_n10914), .B(new_n9298), .Y(new_n10916));
  xor_4  g08568(.A(new_n10890), .B(new_n8058), .Y(new_n10917));
  nor_5  g08569(.A(new_n10917), .B(new_n9256), .Y(new_n10918));
  xor_4  g08570(.A(new_n10885), .B(new_n8059), .Y(new_n10919));
  nor_5  g08571(.A(new_n10919), .B(new_n9258), .Y(new_n10920));
  xor_4  g08572(.A(new_n10919), .B(new_n9259), .Y(new_n10921));
  xor_4  g08573(.A(new_n10879), .B(new_n8060), .Y(new_n10922));
  nor_5  g08574(.A(new_n10922), .B(new_n9260), .Y(new_n10923));
  xnor_4 g08575(.A(new_n10922), .B(new_n9260), .Y(new_n10924));
  xor_4  g08576(.A(new_n10875), .B(new_n8082), .Y(new_n10925));
  and_6  g08577(.A(new_n10925), .B(new_n9278), .Y(new_n10926));
  xnor_4 g08578(.A(new_n10869), .B(new_n10868), .Y(new_n10927));
  or_6   g08579(.A(new_n10927), .B(new_n9262), .Y(new_n10928));
  not_8  g08580(.A(new_n10861), .Y(new_n10929));
  xor_4  g08581(.A(new_n10929), .B(new_n2553), .Y(new_n10930));
  nand_5 g08582(.A(new_n10930), .B(new_n9350), .Y(new_n10931));
  nand_5 g08583(.A(new_n10930), .B(new_n9264), .Y(new_n10932));
  or_6   g08584(.A(new_n10930), .B(new_n9237), .Y(new_n10933));
  nand_5 g08585(.A(new_n10933), .B(new_n10932), .Y(new_n10934));
  xor_4  g08586(.A(new_n10934), .B(new_n9234), .Y(new_n10935));
  nor_5  g08587(.A(new_n10935), .B(new_n10931), .Y(new_n10936));
  not_8  g08588(.A(new_n10935), .Y(new_n10937));
  xor_4  g08589(.A(new_n10866), .B(new_n8069), .Y(new_n10938));
  nor_5  g08590(.A(new_n10938), .B(new_n10937), .Y(new_n10939));
  nor_5  g08591(.A(new_n10939), .B(new_n10936), .Y(new_n10940));
  xor_4  g08592(.A(new_n10927), .B(new_n9262), .Y(new_n10941));
  nand_5 g08593(.A(new_n10941), .B(new_n10940), .Y(new_n10942));
  nand_5 g08594(.A(new_n10942), .B(new_n10928), .Y(new_n10943));
  xor_4  g08595(.A(new_n10925), .B(new_n9277), .Y(new_n10944));
  nor_5  g08596(.A(new_n10944), .B(new_n10943), .Y(new_n10945));
  nor_5  g08597(.A(new_n10945), .B(new_n10926), .Y(new_n10946));
  nor_5  g08598(.A(new_n10946), .B(new_n10924), .Y(new_n10947));
  nor_5  g08599(.A(new_n10947), .B(new_n10923), .Y(new_n10948));
  nor_5  g08600(.A(new_n10948), .B(new_n10921), .Y(new_n10949));
  nor_5  g08601(.A(new_n10949), .B(new_n10920), .Y(new_n10950));
  xor_4  g08602(.A(new_n10917), .B(new_n9257), .Y(new_n10951));
  nor_5  g08603(.A(new_n10951), .B(new_n10950), .Y(new_n10952));
  nor_5  g08604(.A(new_n10952), .B(new_n10918), .Y(new_n10953));
  or_6   g08605(.A(new_n10953), .B(new_n10916), .Y(new_n10954));
  nand_5 g08606(.A(new_n10954), .B(new_n10915), .Y(new_n10955));
  nor_5  g08607(.A(new_n10955), .B(new_n10912), .Y(new_n10956));
  nor_5  g08608(.A(new_n10956), .B(new_n10911), .Y(new_n10957));
  not_8  g08609(.A(new_n10957), .Y(new_n10958));
  xor_4  g08610(.A(new_n9254), .B(pi713), .Y(new_n10959));
  not_8  g08611(.A(new_n10959), .Y(new_n10960));
  nand_5 g08612(.A(new_n10960), .B(new_n8049), .Y(new_n10961));
  nand_5 g08613(.A(new_n10959), .B(new_n8050), .Y(new_n10962));
  nand_5 g08614(.A(new_n10962), .B(new_n10961), .Y(new_n10963));
  xor_4  g08615(.A(pi292), .B(pi141), .Y(new_n10964));
  not_8  g08616(.A(pi108), .Y(new_n10965));
  not_8  g08617(.A(pi541), .Y(new_n10966));
  nand_5 g08618(.A(new_n10966), .B(new_n10965), .Y(new_n10967));
  nand_5 g08619(.A(new_n10906), .B(new_n10903), .Y(new_n10968));
  nand_5 g08620(.A(new_n10968), .B(new_n10967), .Y(new_n10969));
  xor_4  g08621(.A(new_n10969), .B(new_n10964), .Y(new_n10970));
  or_6   g08622(.A(new_n10907), .B(new_n10902), .Y(new_n10971));
  not_8  g08623(.A(new_n8054), .Y(new_n10972));
  nand_5 g08624(.A(new_n10908), .B(new_n10972), .Y(new_n10973));
  nand_5 g08625(.A(new_n10973), .B(new_n10971), .Y(new_n10974));
  xor_4  g08626(.A(new_n10974), .B(new_n10970), .Y(new_n10975));
  xor_4  g08627(.A(new_n10975), .B(new_n10963), .Y(new_n10976));
  xor_4  g08628(.A(new_n10976), .B(new_n10958), .Y(po0065));
  not_8  g08629(.A(pi299), .Y(new_n10978));
  xor_4  g08630(.A(pi631), .B(new_n10978), .Y(new_n10979));
  xor_4  g08631(.A(new_n10979), .B(new_n6024), .Y(new_n10980));
  xor_4  g08632(.A(new_n10980), .B(new_n4988), .Y(po0066));
  nand_5 g08633(.A(pi320), .B(pi133), .Y(new_n10982));
  nand_5 g08634(.A(new_n9656), .B(new_n9643), .Y(new_n10983));
  nand_5 g08635(.A(new_n10983), .B(new_n10982), .Y(new_n10984));
  nand_5 g08636(.A(pi819), .B(pi643), .Y(new_n10985));
  not_8  g08637(.A(pi643), .Y(new_n10986));
  not_8  g08638(.A(pi819), .Y(new_n10987));
  nand_5 g08639(.A(new_n10987), .B(new_n10986), .Y(new_n10988));
  nand_5 g08640(.A(new_n10988), .B(new_n10985), .Y(new_n10989));
  xnor_4 g08641(.A(new_n10989), .B(new_n10984), .Y(new_n10990));
  not_8  g08642(.A(pi767), .Y(new_n10991));
  not_8  g08643(.A(pi366), .Y(new_n10992));
  not_8  g08644(.A(pi651), .Y(new_n10993));
  nand_5 g08645(.A(new_n10993), .B(new_n10992), .Y(new_n10994));
  not_8  g08646(.A(pi169), .Y(new_n10995));
  not_8  g08647(.A(pi481), .Y(new_n10996));
  nand_5 g08648(.A(new_n10996), .B(new_n10995), .Y(new_n10997));
  nor_5  g08649(.A(new_n10997), .B(new_n10994), .Y(new_n10998));
  xor_4  g08650(.A(new_n10998), .B(new_n10991), .Y(new_n10999));
  or_6   g08651(.A(new_n10999), .B(new_n9830), .Y(new_n11000));
  xor_4  g08652(.A(new_n10999), .B(new_n9830), .Y(new_n11001));
  not_8  g08653(.A(new_n9823), .Y(new_n11002));
  nand_5 g08654(.A(new_n9803), .B(new_n10992), .Y(new_n11003));
  not_8  g08655(.A(new_n9803), .Y(new_n11004));
  nand_5 g08656(.A(new_n11004), .B(pi366), .Y(new_n11005));
  nand_5 g08657(.A(new_n9807), .B(pi481), .Y(new_n11006));
  nand_5 g08658(.A(new_n11006), .B(new_n11005), .Y(new_n11007));
  nand_5 g08659(.A(new_n11007), .B(new_n11003), .Y(new_n11008));
  or_6   g08660(.A(new_n11008), .B(new_n9801), .Y(new_n11009));
  nand_5 g08661(.A(new_n11008), .B(new_n9801), .Y(new_n11010));
  nand_5 g08662(.A(new_n11010), .B(pi169), .Y(new_n11011));
  nand_5 g08663(.A(new_n11011), .B(new_n11009), .Y(new_n11012));
  xor_4  g08664(.A(new_n11012), .B(pi651), .Y(new_n11013));
  nand_5 g08665(.A(new_n11013), .B(new_n11002), .Y(new_n11014));
  not_8  g08666(.A(new_n10998), .Y(new_n11015));
  nand_5 g08667(.A(new_n11012), .B(pi651), .Y(new_n11016));
  and_6  g08668(.A(new_n11016), .B(new_n11015), .Y(new_n11017));
  nand_5 g08669(.A(new_n11017), .B(new_n11014), .Y(new_n11018));
  nand_5 g08670(.A(new_n11018), .B(new_n11001), .Y(new_n11019));
  nand_5 g08671(.A(new_n11019), .B(new_n11000), .Y(new_n11020));
  not_8  g08672(.A(pi043), .Y(new_n11021));
  nand_5 g08673(.A(new_n10998), .B(new_n10991), .Y(new_n11022));
  not_8  g08674(.A(new_n11022), .Y(new_n11023));
  nand_5 g08675(.A(new_n11023), .B(new_n11021), .Y(new_n11024));
  not_8  g08676(.A(new_n11024), .Y(new_n11025));
  nor_5  g08677(.A(new_n11023), .B(new_n11021), .Y(new_n11026));
  nor_5  g08678(.A(new_n11026), .B(new_n11025), .Y(new_n11027));
  xor_4  g08679(.A(new_n11027), .B(new_n9835), .Y(new_n11028));
  xor_4  g08680(.A(new_n11028), .B(new_n11020), .Y(new_n11029));
  or_6   g08681(.A(new_n11029), .B(new_n10990), .Y(new_n11030));
  xor_4  g08682(.A(new_n11029), .B(new_n10990), .Y(new_n11031));
  not_8  g08683(.A(new_n11031), .Y(new_n11032));
  not_8  g08684(.A(new_n9657), .Y(new_n11033));
  xnor_4 g08685(.A(new_n11018), .B(new_n11001), .Y(new_n11034));
  nor_5  g08686(.A(new_n11034), .B(new_n11033), .Y(new_n11035));
  xor_4  g08687(.A(new_n11013), .B(new_n11002), .Y(new_n11036));
  or_6   g08688(.A(new_n11036), .B(new_n9718), .Y(new_n11037));
  xor_4  g08689(.A(new_n11036), .B(new_n9718), .Y(new_n11038));
  nand_5 g08690(.A(new_n11010), .B(new_n11009), .Y(new_n11039));
  xor_4  g08691(.A(new_n11039), .B(pi169), .Y(new_n11040));
  nor_5  g08692(.A(new_n11040), .B(new_n9703), .Y(new_n11041));
  xor_4  g08693(.A(new_n11040), .B(new_n9703), .Y(new_n11042));
  not_8  g08694(.A(new_n11006), .Y(new_n11043));
  nand_5 g08695(.A(new_n11043), .B(new_n7247), .Y(new_n11044));
  xor_4  g08696(.A(pi481), .B(new_n7244), .Y(new_n11045));
  xor_4  g08697(.A(new_n11045), .B(pi642), .Y(new_n11046));
  xor_4  g08698(.A(new_n11046), .B(new_n9807), .Y(po1322));
  nand_5 g08699(.A(po1322), .B(new_n7246), .Y(new_n11048));
  nand_5 g08700(.A(new_n11048), .B(new_n7247), .Y(new_n11049));
  nand_5 g08701(.A(new_n11049), .B(new_n11006), .Y(new_n11050));
  nand_5 g08702(.A(new_n11050), .B(new_n11044), .Y(new_n11051));
  nand_5 g08703(.A(new_n11003), .B(new_n11005), .Y(new_n11052));
  xor_4  g08704(.A(new_n11052), .B(new_n9704), .Y(new_n11053));
  xor_4  g08705(.A(new_n11053), .B(new_n11051), .Y(po1489));
  nand_5 g08706(.A(po1489), .B(new_n9704), .Y(new_n11055));
  or_6   g08707(.A(po1489), .B(new_n9704), .Y(new_n11056));
  nand_5 g08708(.A(new_n11056), .B(new_n11049), .Y(new_n11057));
  nand_5 g08709(.A(new_n11057), .B(new_n11055), .Y(new_n11058));
  and_6  g08710(.A(new_n11058), .B(new_n11042), .Y(new_n11059));
  nor_5  g08711(.A(new_n11059), .B(new_n11041), .Y(new_n11060));
  nand_5 g08712(.A(new_n11060), .B(new_n11038), .Y(new_n11061));
  nand_5 g08713(.A(new_n11061), .B(new_n11037), .Y(new_n11062));
  xor_4  g08714(.A(new_n11034), .B(new_n9657), .Y(new_n11063));
  nor_5  g08715(.A(new_n11063), .B(new_n11062), .Y(new_n11064));
  or_6   g08716(.A(new_n11064), .B(new_n11035), .Y(new_n11065));
  or_6   g08717(.A(new_n11065), .B(new_n11032), .Y(new_n11066));
  nand_5 g08718(.A(new_n11066), .B(new_n11030), .Y(new_n11067));
  nand_5 g08719(.A(new_n10988), .B(new_n10984), .Y(new_n11068));
  nand_5 g08720(.A(new_n11068), .B(new_n10985), .Y(new_n11069));
  nand_5 g08721(.A(pi627), .B(pi113), .Y(new_n11070));
  not_8  g08722(.A(pi113), .Y(new_n11071));
  not_8  g08723(.A(pi627), .Y(new_n11072));
  nand_5 g08724(.A(new_n11072), .B(new_n11071), .Y(new_n11073));
  and_6  g08725(.A(new_n11073), .B(new_n11070), .Y(new_n11074));
  xor_4  g08726(.A(new_n11074), .B(new_n11069), .Y(new_n11075));
  not_8  g08727(.A(new_n11075), .Y(new_n11076));
  not_8  g08728(.A(pi015), .Y(new_n11077));
  xor_4  g08729(.A(new_n11024), .B(new_n11077), .Y(new_n11078));
  xor_4  g08730(.A(new_n11078), .B(new_n9843), .Y(new_n11079));
  not_8  g08731(.A(new_n11079), .Y(new_n11080));
  or_6   g08732(.A(new_n11027), .B(new_n9835), .Y(new_n11081));
  nand_5 g08733(.A(new_n11028), .B(new_n11020), .Y(new_n11082));
  nand_5 g08734(.A(new_n11082), .B(new_n11081), .Y(new_n11083));
  xor_4  g08735(.A(new_n11083), .B(new_n11080), .Y(new_n11084));
  xor_4  g08736(.A(new_n11084), .B(new_n11076), .Y(new_n11085));
  xor_4  g08737(.A(new_n11085), .B(new_n11067), .Y(po0067));
  nand_5 g08738(.A(pi610), .B(new_n7590), .Y(new_n11087));
  nand_5 g08739(.A(new_n8969), .B(new_n8967), .Y(new_n11088));
  nand_5 g08740(.A(new_n11088), .B(new_n11087), .Y(new_n11089));
  not_8  g08741(.A(new_n11089), .Y(new_n11090));
  not_8  g08742(.A(pi534), .Y(new_n11091));
  nand_5 g08743(.A(new_n11091), .B(pi465), .Y(new_n11092));
  xor_4  g08744(.A(pi534), .B(new_n10166), .Y(new_n11093));
  nand_5 g08745(.A(pi722), .B(new_n7257), .Y(new_n11094));
  xor_4  g08746(.A(pi722), .B(new_n7257), .Y(new_n11095));
  not_8  g08747(.A(pi772), .Y(new_n11096));
  nand_5 g08748(.A(new_n11096), .B(pi336), .Y(new_n11097));
  xor_4  g08749(.A(pi772), .B(new_n8004), .Y(new_n11098));
  nand_5 g08750(.A(pi470), .B(new_n10647), .Y(new_n11099));
  xor_4  g08751(.A(pi470), .B(new_n10647), .Y(new_n11100));
  not_8  g08752(.A(pi265), .Y(new_n11101));
  nand_5 g08753(.A(pi372), .B(new_n11101), .Y(new_n11102));
  xor_4  g08754(.A(pi372), .B(new_n11101), .Y(new_n11103));
  not_8  g08755(.A(pi001), .Y(new_n11104));
  or_6   g08756(.A(pi635), .B(new_n11104), .Y(new_n11105));
  xor_4  g08757(.A(pi635), .B(new_n11104), .Y(new_n11106));
  nand_5 g08758(.A(new_n7270), .B(pi050), .Y(new_n11107));
  xor_4  g08759(.A(pi545), .B(new_n8015), .Y(new_n11108));
  nand_5 g08760(.A(new_n6575), .B(pi262), .Y(new_n11109));
  not_8  g08761(.A(new_n11109), .Y(new_n11110));
  xor_4  g08762(.A(pi388), .B(new_n8019), .Y(new_n11111));
  not_8  g08763(.A(new_n11111), .Y(new_n11112));
  nand_5 g08764(.A(new_n8027), .B(pi161), .Y(new_n11113));
  nand_5 g08765(.A(pi326), .B(new_n8511), .Y(new_n11114));
  nand_5 g08766(.A(new_n7343), .B(pi122), .Y(new_n11115));
  nand_5 g08767(.A(new_n11115), .B(new_n11114), .Y(new_n11116));
  nand_5 g08768(.A(new_n11116), .B(new_n11113), .Y(new_n11117));
  nor_5  g08769(.A(new_n11117), .B(new_n11112), .Y(new_n11118));
  nor_5  g08770(.A(new_n11118), .B(new_n11110), .Y(new_n11119));
  not_8  g08771(.A(new_n11119), .Y(new_n11120));
  nand_5 g08772(.A(new_n11120), .B(new_n11108), .Y(new_n11121));
  nand_5 g08773(.A(new_n11121), .B(new_n11107), .Y(new_n11122));
  nand_5 g08774(.A(new_n11122), .B(new_n11106), .Y(new_n11123));
  nand_5 g08775(.A(new_n11123), .B(new_n11105), .Y(new_n11124));
  nand_5 g08776(.A(new_n11124), .B(new_n11103), .Y(new_n11125));
  nand_5 g08777(.A(new_n11125), .B(new_n11102), .Y(new_n11126));
  nand_5 g08778(.A(new_n11126), .B(new_n11100), .Y(new_n11127));
  nand_5 g08779(.A(new_n11127), .B(new_n11099), .Y(new_n11128));
  nand_5 g08780(.A(new_n11128), .B(new_n11098), .Y(new_n11129));
  nand_5 g08781(.A(new_n11129), .B(new_n11097), .Y(new_n11130));
  nand_5 g08782(.A(new_n11130), .B(new_n11095), .Y(new_n11131));
  nand_5 g08783(.A(new_n11131), .B(new_n11094), .Y(new_n11132));
  nand_5 g08784(.A(new_n11132), .B(new_n11093), .Y(new_n11133));
  nand_5 g08785(.A(new_n11133), .B(new_n11092), .Y(new_n11134));
  nand_5 g08786(.A(pi582), .B(new_n10405), .Y(new_n11135));
  not_8  g08787(.A(new_n11135), .Y(new_n11136));
  nand_5 g08788(.A(new_n2978), .B(pi016), .Y(new_n11137));
  xor_4  g08789(.A(pi404), .B(new_n2837), .Y(new_n11138));
  nand_5 g08790(.A(new_n2940), .B(pi233), .Y(new_n11139));
  xor_4  g08791(.A(pi527), .B(new_n2814), .Y(new_n11140));
  nand_5 g08792(.A(new_n2944), .B(pi691), .Y(new_n11141));
  xor_4  g08793(.A(pi816), .B(new_n2857), .Y(new_n11142));
  not_8  g08794(.A(pi709), .Y(new_n11143));
  nand_5 g08795(.A(new_n11143), .B(pi407), .Y(new_n11144));
  xor_4  g08796(.A(pi709), .B(new_n2675), .Y(new_n11145));
  or_6   g08797(.A(pi590), .B(new_n2864), .Y(new_n11146));
  nand_5 g08798(.A(new_n4237), .B(new_n4233), .Y(new_n11147));
  nand_5 g08799(.A(new_n11147), .B(new_n11146), .Y(new_n11148));
  nand_5 g08800(.A(new_n11148), .B(new_n11145), .Y(new_n11149));
  nand_5 g08801(.A(new_n11149), .B(new_n11144), .Y(new_n11150));
  nand_5 g08802(.A(new_n11150), .B(new_n11142), .Y(new_n11151));
  nand_5 g08803(.A(new_n11151), .B(new_n11141), .Y(new_n11152));
  nand_5 g08804(.A(new_n11152), .B(new_n11140), .Y(new_n11153));
  nand_5 g08805(.A(new_n11153), .B(new_n11139), .Y(new_n11154));
  nand_5 g08806(.A(new_n11154), .B(new_n11138), .Y(new_n11155));
  nand_5 g08807(.A(new_n11155), .B(new_n11137), .Y(new_n11156));
  xor_4  g08808(.A(pi582), .B(pi095), .Y(new_n11157));
  nor_5  g08809(.A(new_n11157), .B(new_n11156), .Y(new_n11158));
  nor_5  g08810(.A(new_n11158), .B(new_n11136), .Y(new_n11159));
  xor_4  g08811(.A(new_n11159), .B(new_n11134), .Y(new_n11160));
  xor_4  g08812(.A(new_n11132), .B(new_n11093), .Y(new_n11161));
  not_8  g08813(.A(new_n11161), .Y(new_n11162));
  xor_4  g08814(.A(new_n11157), .B(new_n11156), .Y(new_n11163));
  nor_5  g08815(.A(new_n11163), .B(new_n11162), .Y(new_n11164));
  xor_4  g08816(.A(new_n11163), .B(new_n11162), .Y(new_n11165));
  not_8  g08817(.A(new_n11165), .Y(new_n11166));
  xor_4  g08818(.A(new_n11130), .B(new_n11095), .Y(new_n11167));
  xor_4  g08819(.A(new_n11154), .B(new_n11138), .Y(new_n11168));
  or_6   g08820(.A(new_n11168), .B(new_n11167), .Y(new_n11169));
  xor_4  g08821(.A(new_n11128), .B(new_n11098), .Y(new_n11170));
  xor_4  g08822(.A(new_n11152), .B(new_n11140), .Y(new_n11171));
  or_6   g08823(.A(new_n11171), .B(new_n11170), .Y(new_n11172));
  xor_4  g08824(.A(new_n11171), .B(new_n11170), .Y(new_n11173));
  xor_4  g08825(.A(new_n11126), .B(new_n11100), .Y(new_n11174));
  not_8  g08826(.A(new_n11174), .Y(new_n11175));
  xor_4  g08827(.A(new_n11150), .B(new_n11142), .Y(new_n11176));
  not_8  g08828(.A(new_n11176), .Y(new_n11177));
  nand_5 g08829(.A(new_n11177), .B(new_n11175), .Y(new_n11178));
  xor_4  g08830(.A(new_n11176), .B(new_n11174), .Y(new_n11179));
  not_8  g08831(.A(new_n11179), .Y(new_n11180));
  xor_4  g08832(.A(new_n11124), .B(new_n11103), .Y(new_n11181));
  xor_4  g08833(.A(new_n11148), .B(new_n11145), .Y(new_n11182));
  nor_5  g08834(.A(new_n11182), .B(new_n11181), .Y(new_n11183));
  xor_4  g08835(.A(new_n11182), .B(new_n11181), .Y(new_n11184));
  not_8  g08836(.A(new_n11184), .Y(new_n11185));
  xor_4  g08837(.A(new_n11122), .B(new_n11106), .Y(new_n11186));
  nand_5 g08838(.A(new_n11186), .B(new_n4238), .Y(new_n11187));
  xor_4  g08839(.A(new_n11186), .B(new_n4238), .Y(new_n11188));
  xor_4  g08840(.A(new_n11119), .B(new_n11108), .Y(new_n11189));
  or_6   g08841(.A(new_n11189), .B(new_n4173), .Y(new_n11190));
  xor_4  g08842(.A(new_n11117), .B(new_n11111), .Y(new_n11191));
  nand_5 g08843(.A(new_n11191), .B(new_n4177), .Y(new_n11192));
  not_8  g08844(.A(new_n11192), .Y(new_n11193));
  xor_4  g08845(.A(new_n11191), .B(new_n4178), .Y(new_n11194));
  and_6  g08846(.A(new_n11114), .B(new_n11113), .Y(new_n11195));
  xnor_4 g08847(.A(new_n11195), .B(new_n11115), .Y(new_n11196));
  nand_5 g08848(.A(new_n11196), .B(new_n4188), .Y(new_n11197));
  nand_5 g08849(.A(pi281), .B(new_n8025), .Y(new_n11198));
  xor_4  g08850(.A(new_n11198), .B(new_n11195), .Y(new_n11199));
  or_6   g08851(.A(new_n11199), .B(new_n4188), .Y(new_n11200));
  nand_5 g08852(.A(new_n11200), .B(new_n11197), .Y(new_n11201));
  nor_5  g08853(.A(new_n11201), .B(new_n4194), .Y(new_n11202));
  nand_5 g08854(.A(new_n11198), .B(new_n11115), .Y(new_n11203));
  not_8  g08855(.A(new_n11203), .Y(new_n11204));
  nor_5  g08856(.A(new_n11204), .B(new_n11200), .Y(new_n11205));
  nor_5  g08857(.A(new_n11205), .B(new_n11202), .Y(new_n11206));
  nor_5  g08858(.A(new_n11206), .B(new_n11194), .Y(new_n11207));
  nor_5  g08859(.A(new_n11207), .B(new_n11193), .Y(new_n11208));
  xor_4  g08860(.A(new_n11189), .B(new_n4173), .Y(new_n11209));
  nand_5 g08861(.A(new_n11209), .B(new_n11208), .Y(new_n11210));
  nand_5 g08862(.A(new_n11210), .B(new_n11190), .Y(new_n11211));
  nand_5 g08863(.A(new_n11211), .B(new_n11188), .Y(new_n11212));
  nand_5 g08864(.A(new_n11212), .B(new_n11187), .Y(new_n11213));
  nor_5  g08865(.A(new_n11213), .B(new_n11185), .Y(new_n11214));
  nor_5  g08866(.A(new_n11214), .B(new_n11183), .Y(new_n11215));
  or_6   g08867(.A(new_n11215), .B(new_n11180), .Y(new_n11216));
  nand_5 g08868(.A(new_n11216), .B(new_n11178), .Y(new_n11217));
  nand_5 g08869(.A(new_n11217), .B(new_n11173), .Y(new_n11218));
  nand_5 g08870(.A(new_n11218), .B(new_n11172), .Y(new_n11219));
  not_8  g08871(.A(new_n11168), .Y(new_n11220));
  xor_4  g08872(.A(new_n11220), .B(new_n11167), .Y(new_n11221));
  not_8  g08873(.A(new_n11221), .Y(new_n11222));
  nand_5 g08874(.A(new_n11222), .B(new_n11219), .Y(new_n11223));
  nand_5 g08875(.A(new_n11223), .B(new_n11169), .Y(new_n11224));
  nor_5  g08876(.A(new_n11224), .B(new_n11166), .Y(new_n11225));
  nor_5  g08877(.A(new_n11225), .B(new_n11164), .Y(new_n11226));
  xor_4  g08878(.A(new_n11226), .B(new_n11160), .Y(new_n11227));
  not_8  g08879(.A(new_n11227), .Y(new_n11228));
  nand_5 g08880(.A(new_n11228), .B(new_n11090), .Y(new_n11229));
  xor_4  g08881(.A(new_n11227), .B(new_n11090), .Y(new_n11230));
  xor_4  g08882(.A(new_n11217), .B(new_n11173), .Y(new_n11231));
  xor_4  g08883(.A(new_n11215), .B(new_n11180), .Y(new_n11232));
  not_8  g08884(.A(new_n8815), .Y(new_n11233));
  xor_4  g08885(.A(new_n11204), .B(new_n4188), .Y(new_n11234));
  not_8  g08886(.A(new_n11234), .Y(new_n11235));
  nor_5  g08887(.A(new_n11235), .B(new_n7250), .Y(new_n11236));
  nor_5  g08888(.A(new_n11236), .B(new_n8834), .Y(new_n11237));
  xor_4  g08889(.A(new_n11201), .B(new_n4194), .Y(new_n11238));
  xor_4  g08890(.A(new_n11236), .B(new_n8833), .Y(new_n11239));
  nor_5  g08891(.A(new_n11239), .B(new_n11238), .Y(new_n11240));
  or_6   g08892(.A(new_n11240), .B(new_n11237), .Y(new_n11241));
  nand_5 g08893(.A(new_n11241), .B(new_n8825), .Y(new_n11242));
  xnor_4 g08894(.A(new_n11241), .B(new_n8825), .Y(new_n11243));
  xor_4  g08895(.A(new_n11206), .B(new_n11194), .Y(new_n11244));
  or_6   g08896(.A(new_n11244), .B(new_n11243), .Y(new_n11245));
  nand_5 g08897(.A(new_n11245), .B(new_n11242), .Y(new_n11246));
  or_6   g08898(.A(new_n11246), .B(new_n8820), .Y(new_n11247));
  xor_4  g08899(.A(new_n11209), .B(new_n11208), .Y(new_n11248));
  not_8  g08900(.A(new_n11248), .Y(new_n11249));
  xor_4  g08901(.A(new_n11246), .B(new_n8820), .Y(new_n11250));
  nand_5 g08902(.A(new_n11250), .B(new_n11249), .Y(new_n11251));
  nand_5 g08903(.A(new_n11251), .B(new_n11247), .Y(new_n11252));
  nor_5  g08904(.A(new_n11252), .B(new_n11233), .Y(new_n11253));
  xor_4  g08905(.A(new_n11252), .B(new_n8815), .Y(new_n11254));
  xor_4  g08906(.A(new_n11211), .B(new_n11188), .Y(new_n11255));
  not_8  g08907(.A(new_n11255), .Y(new_n11256));
  nor_5  g08908(.A(new_n11256), .B(new_n11254), .Y(new_n11257));
  or_6   g08909(.A(new_n11257), .B(new_n11253), .Y(new_n11258));
  xor_4  g08910(.A(new_n11213), .B(new_n11184), .Y(new_n11259));
  nor_5  g08911(.A(new_n11259), .B(new_n11258), .Y(new_n11260));
  not_8  g08912(.A(new_n11259), .Y(new_n11261));
  xor_4  g08913(.A(new_n11261), .B(new_n11258), .Y(new_n11262));
  nor_5  g08914(.A(new_n11262), .B(new_n8812), .Y(new_n11263));
  or_6   g08915(.A(new_n11263), .B(new_n11260), .Y(new_n11264));
  nand_5 g08916(.A(new_n11264), .B(new_n11232), .Y(new_n11265));
  not_8  g08917(.A(new_n11232), .Y(new_n11266));
  xor_4  g08918(.A(new_n11264), .B(new_n11266), .Y(new_n11267));
  or_6   g08919(.A(new_n11267), .B(new_n8808), .Y(new_n11268));
  nand_5 g08920(.A(new_n11268), .B(new_n11265), .Y(new_n11269));
  nand_5 g08921(.A(new_n11269), .B(new_n11231), .Y(new_n11270));
  xor_4  g08922(.A(new_n11269), .B(new_n11231), .Y(new_n11271));
  not_8  g08923(.A(new_n11271), .Y(new_n11272));
  or_6   g08924(.A(new_n11272), .B(new_n8804), .Y(new_n11273));
  nand_5 g08925(.A(new_n11273), .B(new_n11270), .Y(new_n11274));
  xor_4  g08926(.A(new_n11221), .B(new_n11219), .Y(new_n11275));
  not_8  g08927(.A(new_n11275), .Y(new_n11276));
  nor_5  g08928(.A(new_n11276), .B(new_n11274), .Y(new_n11277));
  xor_4  g08929(.A(new_n11275), .B(new_n11274), .Y(new_n11278));
  nor_5  g08930(.A(new_n11278), .B(new_n8756), .Y(new_n11279));
  nor_5  g08931(.A(new_n11279), .B(new_n11277), .Y(new_n11280));
  nand_5 g08932(.A(new_n11280), .B(new_n8971), .Y(new_n11281));
  xor_4  g08933(.A(new_n11280), .B(new_n8971), .Y(new_n11282));
  xor_4  g08934(.A(new_n11224), .B(new_n11165), .Y(new_n11283));
  nand_5 g08935(.A(new_n11283), .B(new_n11282), .Y(new_n11284));
  nand_5 g08936(.A(new_n11284), .B(new_n11281), .Y(new_n11285));
  or_6   g08937(.A(new_n11285), .B(new_n11230), .Y(new_n11286));
  nand_5 g08938(.A(new_n11286), .B(new_n11229), .Y(new_n11287));
  or_6   g08939(.A(new_n11159), .B(new_n11134), .Y(new_n11288));
  nand_5 g08940(.A(new_n11226), .B(new_n11160), .Y(new_n11289));
  nand_5 g08941(.A(new_n11289), .B(new_n11288), .Y(new_n11290));
  xor_4  g08942(.A(new_n11290), .B(new_n11090), .Y(new_n11291));
  xnor_4 g08943(.A(new_n11291), .B(new_n11287), .Y(po0068));
  not_8  g08944(.A(new_n7966), .Y(new_n11293));
  not_8  g08945(.A(pi348), .Y(new_n11294));
  nand_5 g08946(.A(pi429), .B(new_n11294), .Y(new_n11295));
  xor_4  g08947(.A(pi429), .B(new_n11294), .Y(new_n11296));
  nand_5 g08948(.A(pi699), .B(new_n2470), .Y(new_n11297));
  xor_4  g08949(.A(pi699), .B(new_n2470), .Y(new_n11298));
  nand_5 g08950(.A(new_n2472), .B(pi055), .Y(new_n11299));
  xor_4  g08951(.A(pi662), .B(new_n2405), .Y(new_n11300));
  nand_5 g08952(.A(new_n2476), .B(pi289), .Y(new_n11301));
  xor_4  g08953(.A(pi831), .B(new_n2385), .Y(new_n11302));
  nand_5 g08954(.A(new_n2480), .B(pi486), .Y(new_n11303));
  or_6   g08955(.A(new_n9867), .B(new_n9863), .Y(new_n11304));
  nand_5 g08956(.A(new_n11304), .B(new_n11303), .Y(new_n11305));
  nand_5 g08957(.A(new_n11305), .B(new_n11302), .Y(new_n11306));
  nand_5 g08958(.A(new_n11306), .B(new_n11301), .Y(new_n11307));
  nand_5 g08959(.A(new_n11307), .B(new_n11300), .Y(new_n11308));
  nand_5 g08960(.A(new_n11308), .B(new_n11299), .Y(new_n11309));
  nand_5 g08961(.A(new_n11309), .B(new_n11298), .Y(new_n11310));
  nand_5 g08962(.A(new_n11310), .B(new_n11297), .Y(new_n11311));
  nand_5 g08963(.A(new_n11311), .B(new_n11296), .Y(new_n11312));
  nand_5 g08964(.A(new_n11312), .B(new_n11295), .Y(new_n11313));
  xor_4  g08965(.A(pi417), .B(new_n5457), .Y(new_n11314));
  xor_4  g08966(.A(new_n11314), .B(new_n11313), .Y(new_n11315));
  nor_5  g08967(.A(new_n11315), .B(new_n11293), .Y(new_n11316));
  xor_4  g08968(.A(new_n11315), .B(new_n11293), .Y(new_n11317));
  xnor_4 g08969(.A(new_n11311), .B(new_n11296), .Y(new_n11318));
  or_6   g08970(.A(new_n11318), .B(new_n7960), .Y(new_n11319));
  not_8  g08971(.A(new_n7955), .Y(new_n11320));
  xor_4  g08972(.A(new_n11309), .B(new_n11298), .Y(new_n11321));
  nand_5 g08973(.A(new_n11321), .B(new_n11320), .Y(new_n11322));
  xor_4  g08974(.A(new_n11321), .B(new_n7955), .Y(new_n11323));
  xor_4  g08975(.A(new_n11307), .B(new_n11300), .Y(new_n11324));
  or_6   g08976(.A(new_n11324), .B(new_n7950), .Y(new_n11325));
  xor_4  g08977(.A(new_n11324), .B(new_n7950), .Y(new_n11326));
  xnor_4 g08978(.A(new_n11305), .B(new_n11302), .Y(new_n11327));
  nor_5  g08979(.A(new_n11327), .B(new_n7942), .Y(new_n11328));
  xor_4  g08980(.A(new_n11327), .B(new_n7941), .Y(new_n11329));
  and_6  g08981(.A(new_n9868), .B(new_n7919), .Y(new_n11330));
  nor_5  g08982(.A(new_n9884), .B(new_n9869), .Y(new_n11331));
  nor_5  g08983(.A(new_n11331), .B(new_n11330), .Y(new_n11332));
  nor_5  g08984(.A(new_n11332), .B(new_n11329), .Y(new_n11333));
  nor_5  g08985(.A(new_n11333), .B(new_n11328), .Y(new_n11334));
  nand_5 g08986(.A(new_n11334), .B(new_n11326), .Y(new_n11335));
  nand_5 g08987(.A(new_n11335), .B(new_n11325), .Y(new_n11336));
  or_6   g08988(.A(new_n11336), .B(new_n11323), .Y(new_n11337));
  nand_5 g08989(.A(new_n11337), .B(new_n11322), .Y(new_n11338));
  xor_4  g08990(.A(new_n11318), .B(new_n7960), .Y(new_n11339));
  nand_5 g08991(.A(new_n11339), .B(new_n11338), .Y(new_n11340));
  nand_5 g08992(.A(new_n11340), .B(new_n11319), .Y(new_n11341));
  not_8  g08993(.A(new_n11341), .Y(new_n11342));
  and_6  g08994(.A(new_n11342), .B(new_n11317), .Y(new_n11343));
  nor_5  g08995(.A(new_n11343), .B(new_n11316), .Y(new_n11344));
  not_8  g08996(.A(pi417), .Y(new_n11345));
  nand_5 g08997(.A(new_n11345), .B(pi319), .Y(new_n11346));
  nand_5 g08998(.A(new_n11314), .B(new_n11313), .Y(new_n11347));
  nand_5 g08999(.A(new_n11347), .B(new_n11346), .Y(new_n11348));
  not_8  g09000(.A(pi721), .Y(new_n11349));
  nand_5 g09001(.A(pi777), .B(new_n11349), .Y(new_n11350));
  nand_5 g09002(.A(new_n5454), .B(pi721), .Y(new_n11351));
  nand_5 g09003(.A(new_n11351), .B(new_n11350), .Y(new_n11352));
  xor_4  g09004(.A(new_n11352), .B(new_n11348), .Y(new_n11353));
  xor_4  g09005(.A(new_n11353), .B(new_n7875), .Y(new_n11354));
  xnor_4 g09006(.A(new_n11354), .B(new_n11344), .Y(po0069));
  nand_5 g09007(.A(new_n7344), .B(pi569), .Y(new_n11356));
  nand_5 g09008(.A(new_n7345), .B(new_n6766), .Y(new_n11357));
  nand_5 g09009(.A(new_n11357), .B(new_n11356), .Y(new_n11358));
  or_6   g09010(.A(new_n8487), .B(new_n8469), .Y(new_n11359));
  nor_5  g09011(.A(new_n11359), .B(new_n3818), .Y(new_n11360));
  nor_5  g09012(.A(new_n11360), .B(new_n11358), .Y(new_n11361));
  nand_5 g09013(.A(new_n3816), .B(new_n2429), .Y(new_n11362));
  nand_5 g09014(.A(new_n11362), .B(new_n3787), .Y(new_n11363));
  not_8  g09015(.A(new_n11363), .Y(new_n11364));
  nor_5  g09016(.A(new_n11364), .B(new_n11357), .Y(new_n11365));
  nor_5  g09017(.A(new_n11363), .B(new_n11356), .Y(new_n11366));
  or_6   g09018(.A(new_n11366), .B(new_n11365), .Y(new_n11367));
  nor_5  g09019(.A(new_n11367), .B(new_n11361), .Y(new_n11368));
  xor_4  g09020(.A(new_n11368), .B(new_n7350), .Y(new_n11369));
  nand_5 g09021(.A(new_n6732), .B(pi132), .Y(new_n11370));
  nand_5 g09022(.A(pi333), .B(new_n2391), .Y(new_n11371));
  nand_5 g09023(.A(new_n11371), .B(new_n11370), .Y(new_n11372));
  xnor_4 g09024(.A(new_n11372), .B(new_n11369), .Y(po0070));
  nand_5 g09025(.A(pi331), .B(new_n8294), .Y(new_n11374));
  xor_4  g09026(.A(pi331), .B(new_n8294), .Y(new_n11375));
  nand_5 g09027(.A(new_n8297), .B(pi428), .Y(new_n11376));
  xor_4  g09028(.A(pi684), .B(new_n3533), .Y(new_n11377));
  nand_5 g09029(.A(new_n8300), .B(pi196), .Y(new_n11378));
  xor_4  g09030(.A(pi742), .B(new_n3536), .Y(new_n11379));
  nand_5 g09031(.A(new_n4685), .B(new_n4682), .Y(new_n11380));
  nand_5 g09032(.A(new_n11380), .B(new_n4684), .Y(new_n11381));
  nand_5 g09033(.A(new_n11381), .B(new_n11379), .Y(new_n11382));
  nand_5 g09034(.A(new_n11382), .B(new_n11378), .Y(new_n11383));
  nand_5 g09035(.A(new_n11383), .B(new_n11377), .Y(new_n11384));
  nand_5 g09036(.A(new_n11384), .B(new_n11376), .Y(new_n11385));
  nand_5 g09037(.A(new_n11385), .B(new_n11375), .Y(new_n11386));
  nand_5 g09038(.A(new_n11386), .B(new_n11374), .Y(new_n11387));
  nand_5 g09039(.A(pi785), .B(new_n8381), .Y(new_n11388));
  nand_5 g09040(.A(new_n3695), .B(pi034), .Y(new_n11389));
  and_6  g09041(.A(new_n11389), .B(new_n11388), .Y(new_n11390));
  xor_4  g09042(.A(new_n11390), .B(new_n11387), .Y(new_n11391));
  not_8  g09043(.A(new_n11391), .Y(new_n11392));
  not_8  g09044(.A(pi729), .Y(new_n11393));
  xor_4  g09045(.A(pi773), .B(new_n11393), .Y(new_n11394));
  not_8  g09046(.A(pi257), .Y(new_n11395));
  nand_5 g09047(.A(pi608), .B(new_n11395), .Y(new_n11396));
  xor_4  g09048(.A(pi608), .B(new_n11395), .Y(new_n11397));
  not_8  g09049(.A(pi035), .Y(new_n11398));
  or_6   g09050(.A(pi182), .B(new_n11398), .Y(new_n11399));
  xor_4  g09051(.A(pi182), .B(new_n11398), .Y(new_n11400));
  nand_5 g09052(.A(pi603), .B(new_n6540), .Y(new_n11401));
  nand_5 g09053(.A(new_n6543), .B(new_n6541), .Y(new_n11402));
  nand_5 g09054(.A(new_n11402), .B(new_n11401), .Y(new_n11403));
  nand_5 g09055(.A(new_n11403), .B(new_n11400), .Y(new_n11404));
  nand_5 g09056(.A(new_n11404), .B(new_n11399), .Y(new_n11405));
  nand_5 g09057(.A(new_n11405), .B(new_n11397), .Y(new_n11406));
  nand_5 g09058(.A(new_n11406), .B(new_n11396), .Y(new_n11407));
  xnor_4 g09059(.A(new_n11407), .B(new_n11394), .Y(new_n11408));
  xor_4  g09060(.A(new_n11408), .B(new_n11392), .Y(new_n11409));
  xnor_4 g09061(.A(new_n11385), .B(new_n11375), .Y(new_n11410));
  xor_4  g09062(.A(new_n11405), .B(new_n11397), .Y(new_n11411));
  not_8  g09063(.A(new_n11411), .Y(new_n11412));
  or_6   g09064(.A(new_n11412), .B(new_n11410), .Y(new_n11413));
  xor_4  g09065(.A(new_n11412), .B(new_n11410), .Y(new_n11414));
  xor_4  g09066(.A(new_n11383), .B(new_n11377), .Y(new_n11415));
  xor_4  g09067(.A(new_n11403), .B(new_n11400), .Y(new_n11416));
  nor_5  g09068(.A(new_n11416), .B(new_n11415), .Y(new_n11417));
  xor_4  g09069(.A(new_n11416), .B(new_n11415), .Y(new_n11418));
  not_8  g09070(.A(new_n11418), .Y(new_n11419));
  xnor_4 g09071(.A(new_n11381), .B(new_n11379), .Y(new_n11420));
  or_6   g09072(.A(new_n11420), .B(new_n6545), .Y(new_n11421));
  xor_4  g09073(.A(new_n11420), .B(new_n6545), .Y(new_n11422));
  or_6   g09074(.A(new_n4696), .B(new_n4687), .Y(new_n11423));
  nand_5 g09075(.A(new_n4703), .B(new_n4697), .Y(new_n11424));
  nand_5 g09076(.A(new_n11424), .B(new_n11423), .Y(new_n11425));
  nand_5 g09077(.A(new_n11425), .B(new_n11422), .Y(new_n11426));
  nand_5 g09078(.A(new_n11426), .B(new_n11421), .Y(new_n11427));
  nor_5  g09079(.A(new_n11427), .B(new_n11419), .Y(new_n11428));
  nor_5  g09080(.A(new_n11428), .B(new_n11417), .Y(new_n11429));
  nand_5 g09081(.A(new_n11429), .B(new_n11414), .Y(new_n11430));
  nand_5 g09082(.A(new_n11430), .B(new_n11413), .Y(new_n11431));
  xor_4  g09083(.A(new_n11431), .B(new_n11409), .Y(new_n11432));
  not_8  g09084(.A(pi039), .Y(new_n11433));
  xor_4  g09085(.A(pi593), .B(new_n11433), .Y(new_n11434));
  not_8  g09086(.A(pi266), .Y(new_n11435));
  nand_5 g09087(.A(pi744), .B(new_n11435), .Y(new_n11436));
  or_6   g09088(.A(pi744), .B(new_n11435), .Y(new_n11437));
  not_8  g09089(.A(pi706), .Y(new_n11438));
  or_6   g09090(.A(pi727), .B(new_n11438), .Y(new_n11439));
  xor_4  g09091(.A(pi727), .B(new_n11438), .Y(new_n11440));
  nand_5 g09092(.A(new_n6551), .B(new_n6548), .Y(new_n11441));
  nand_5 g09093(.A(new_n11441), .B(new_n6550), .Y(new_n11442));
  nand_5 g09094(.A(new_n11442), .B(new_n11440), .Y(new_n11443));
  nand_5 g09095(.A(new_n11443), .B(new_n11439), .Y(new_n11444));
  nand_5 g09096(.A(new_n11444), .B(new_n11437), .Y(new_n11445));
  nand_5 g09097(.A(new_n11445), .B(new_n11436), .Y(new_n11446));
  xor_4  g09098(.A(new_n11446), .B(new_n11434), .Y(new_n11447));
  xor_4  g09099(.A(new_n11447), .B(new_n11432), .Y(new_n11448));
  xor_4  g09100(.A(new_n11429), .B(new_n11414), .Y(new_n11449));
  and_6  g09101(.A(new_n11437), .B(new_n11436), .Y(new_n11450));
  xor_4  g09102(.A(new_n11450), .B(new_n11444), .Y(new_n11451));
  nand_5 g09103(.A(new_n11451), .B(new_n11449), .Y(new_n11452));
  xor_4  g09104(.A(new_n11427), .B(new_n11419), .Y(new_n11453));
  xor_4  g09105(.A(new_n11442), .B(new_n11440), .Y(new_n11454));
  not_8  g09106(.A(new_n11454), .Y(new_n11455));
  nor_5  g09107(.A(new_n11455), .B(new_n11453), .Y(new_n11456));
  xor_4  g09108(.A(new_n11454), .B(new_n11453), .Y(new_n11457));
  xor_4  g09109(.A(new_n11425), .B(new_n11422), .Y(new_n11458));
  or_6   g09110(.A(new_n11458), .B(new_n6553), .Y(new_n11459));
  nand_5 g09111(.A(new_n11458), .B(new_n6553), .Y(new_n11460));
  not_8  g09112(.A(new_n6426), .Y(new_n11461));
  nand_5 g09113(.A(new_n6475), .B(new_n4628), .Y(new_n11462));
  nand_5 g09114(.A(new_n6415), .B(new_n4630), .Y(new_n11463));
  nand_5 g09115(.A(new_n11463), .B(new_n11462), .Y(new_n11464));
  xor_4  g09116(.A(new_n11464), .B(new_n6485), .Y(new_n11465));
  or_6   g09117(.A(new_n11465), .B(new_n4603), .Y(new_n11466));
  nand_5 g09118(.A(new_n6476), .B(new_n4628), .Y(new_n11467));
  nand_5 g09119(.A(new_n11467), .B(new_n11465), .Y(new_n11468));
  nand_5 g09120(.A(new_n11468), .B(new_n11466), .Y(new_n11469));
  nand_5 g09121(.A(new_n11469), .B(new_n6467), .Y(new_n11470));
  xor_4  g09122(.A(new_n11469), .B(new_n6468), .Y(new_n11471));
  or_6   g09123(.A(new_n11471), .B(new_n4648), .Y(new_n11472));
  nand_5 g09124(.A(new_n11472), .B(new_n11470), .Y(new_n11473));
  nand_5 g09125(.A(new_n11473), .B(new_n6462), .Y(new_n11474));
  xnor_4 g09126(.A(new_n11473), .B(new_n6462), .Y(new_n11475));
  or_6   g09127(.A(new_n11475), .B(new_n4662), .Y(new_n11476));
  nand_5 g09128(.A(new_n11476), .B(new_n11474), .Y(new_n11477));
  nand_5 g09129(.A(new_n11477), .B(new_n6457), .Y(new_n11478));
  not_8  g09130(.A(new_n11478), .Y(new_n11479));
  xnor_4 g09131(.A(new_n11477), .B(new_n6457), .Y(new_n11480));
  nor_5  g09132(.A(new_n11480), .B(new_n4675), .Y(new_n11481));
  nor_5  g09133(.A(new_n11481), .B(new_n11479), .Y(new_n11482));
  nand_5 g09134(.A(new_n11482), .B(new_n11461), .Y(new_n11483));
  xor_4  g09135(.A(new_n11482), .B(new_n11461), .Y(new_n11484));
  nand_5 g09136(.A(new_n11484), .B(new_n4704), .Y(new_n11485));
  nand_5 g09137(.A(new_n11485), .B(new_n11483), .Y(new_n11486));
  nand_5 g09138(.A(new_n11486), .B(new_n11460), .Y(new_n11487));
  nand_5 g09139(.A(new_n11487), .B(new_n11459), .Y(new_n11488));
  nor_5  g09140(.A(new_n11488), .B(new_n11457), .Y(new_n11489));
  nor_5  g09141(.A(new_n11489), .B(new_n11456), .Y(new_n11490));
  not_8  g09142(.A(new_n11449), .Y(new_n11491));
  xor_4  g09143(.A(new_n11451), .B(new_n11491), .Y(new_n11492));
  or_6   g09144(.A(new_n11492), .B(new_n11490), .Y(new_n11493));
  nand_5 g09145(.A(new_n11493), .B(new_n11452), .Y(new_n11494));
  xnor_4 g09146(.A(new_n11494), .B(new_n11448), .Y(po0071));
  xnor_4 g09147(.A(new_n7667), .B(new_n7666), .Y(po0072));
  xnor_4 g09148(.A(new_n2827), .B(new_n2825), .Y(po0073));
  xnor_4 g09149(.A(new_n11492), .B(new_n11490), .Y(po0074));
  not_8  g09150(.A(pi148), .Y(new_n11499));
  not_8  g09151(.A(pi340), .Y(new_n11500));
  nand_5 g09152(.A(new_n11500), .B(new_n11499), .Y(new_n11501));
  not_8  g09153(.A(new_n11501), .Y(new_n11502));
  nand_5 g09154(.A(pi340), .B(pi148), .Y(new_n11503));
  not_8  g09155(.A(new_n11503), .Y(new_n11504));
  not_8  g09156(.A(pi135), .Y(new_n11505));
  not_8  g09157(.A(pi561), .Y(new_n11506));
  nand_5 g09158(.A(new_n11506), .B(new_n11505), .Y(new_n11507));
  not_8  g09159(.A(new_n11507), .Y(new_n11508));
  nand_5 g09160(.A(pi561), .B(pi135), .Y(new_n11509));
  not_8  g09161(.A(new_n11509), .Y(new_n11510));
  not_8  g09162(.A(pi199), .Y(new_n11511));
  not_8  g09163(.A(pi598), .Y(new_n11512));
  nand_5 g09164(.A(new_n11512), .B(new_n11511), .Y(new_n11513));
  not_8  g09165(.A(new_n11513), .Y(new_n11514));
  xor_4  g09166(.A(pi598), .B(pi199), .Y(new_n11515));
  not_8  g09167(.A(new_n11515), .Y(new_n11516));
  nand_5 g09168(.A(new_n11073), .B(new_n11069), .Y(new_n11517));
  nand_5 g09169(.A(new_n11517), .B(new_n11070), .Y(new_n11518));
  nor_5  g09170(.A(new_n11518), .B(new_n11516), .Y(new_n11519));
  nor_5  g09171(.A(new_n11519), .B(new_n11514), .Y(new_n11520));
  nor_5  g09172(.A(new_n11520), .B(new_n11510), .Y(new_n11521));
  nor_5  g09173(.A(new_n11521), .B(new_n11508), .Y(new_n11522));
  nor_5  g09174(.A(new_n11522), .B(new_n11504), .Y(new_n11523));
  nor_5  g09175(.A(new_n11523), .B(new_n11502), .Y(new_n11524));
  xor_4  g09176(.A(pi565), .B(pi096), .Y(new_n11525));
  not_8  g09177(.A(pi784), .Y(new_n11526));
  nand_5 g09178(.A(new_n11526), .B(new_n7592), .Y(new_n11527));
  nand_5 g09179(.A(new_n6934), .B(new_n6931), .Y(new_n11528));
  nand_5 g09180(.A(new_n11528), .B(new_n11527), .Y(new_n11529));
  xor_4  g09181(.A(new_n11529), .B(new_n11525), .Y(new_n11530));
  or_6   g09182(.A(new_n11530), .B(new_n2608), .Y(new_n11531));
  xor_4  g09183(.A(new_n11530), .B(new_n2608), .Y(new_n11532));
  or_6   g09184(.A(new_n6935), .B(new_n8751), .Y(new_n11533));
  xor_4  g09185(.A(new_n6935), .B(new_n8751), .Y(new_n11534));
  nand_5 g09186(.A(new_n6792), .B(pi551), .Y(new_n11535));
  xor_4  g09187(.A(new_n6792), .B(pi551), .Y(new_n11536));
  not_8  g09188(.A(pi420), .Y(new_n11537));
  or_6   g09189(.A(new_n6743), .B(new_n11537), .Y(new_n11538));
  xor_4  g09190(.A(new_n6743), .B(new_n11537), .Y(new_n11539));
  nand_5 g09191(.A(new_n6747), .B(pi115), .Y(new_n11540));
  xor_4  g09192(.A(new_n6747), .B(pi115), .Y(new_n11541));
  nand_5 g09193(.A(new_n9673), .B(new_n9672), .Y(new_n11542));
  nand_5 g09194(.A(new_n11542), .B(new_n9674), .Y(new_n11543));
  nand_5 g09195(.A(new_n11543), .B(new_n11541), .Y(new_n11544));
  nand_5 g09196(.A(new_n11544), .B(new_n11540), .Y(new_n11545));
  nand_5 g09197(.A(new_n11545), .B(new_n11539), .Y(new_n11546));
  nand_5 g09198(.A(new_n11546), .B(new_n11538), .Y(new_n11547));
  nand_5 g09199(.A(new_n11547), .B(new_n11536), .Y(new_n11548));
  nand_5 g09200(.A(new_n11548), .B(new_n11535), .Y(new_n11549));
  nand_5 g09201(.A(new_n11549), .B(new_n11534), .Y(new_n11550));
  nand_5 g09202(.A(new_n11550), .B(new_n11533), .Y(new_n11551));
  nand_5 g09203(.A(new_n11551), .B(new_n11532), .Y(new_n11552));
  nand_5 g09204(.A(new_n11552), .B(new_n11531), .Y(new_n11553));
  or_6   g09205(.A(pi565), .B(pi096), .Y(new_n11554));
  nand_5 g09206(.A(new_n11529), .B(new_n11525), .Y(new_n11555));
  nand_5 g09207(.A(new_n11555), .B(new_n11554), .Y(new_n11556));
  not_8  g09208(.A(new_n11556), .Y(new_n11557));
  nand_5 g09209(.A(new_n11557), .B(new_n11553), .Y(new_n11558));
  nor_5  g09210(.A(new_n11557), .B(new_n11553), .Y(new_n11559));
  not_8  g09211(.A(new_n11559), .Y(new_n11560));
  nand_5 g09212(.A(new_n11560), .B(new_n11558), .Y(new_n11561));
  not_8  g09213(.A(new_n11561), .Y(new_n11562));
  xor_4  g09214(.A(new_n11551), .B(new_n11532), .Y(new_n11563));
  not_8  g09215(.A(new_n11563), .Y(new_n11564));
  xor_4  g09216(.A(new_n11547), .B(new_n11536), .Y(new_n11565));
  not_8  g09217(.A(new_n11565), .Y(new_n11566));
  nand_5 g09218(.A(new_n11566), .B(pi179), .Y(new_n11567));
  not_8  g09219(.A(pi179), .Y(new_n11568));
  xor_4  g09220(.A(new_n11565), .B(new_n11568), .Y(new_n11569));
  xor_4  g09221(.A(new_n11543), .B(new_n11541), .Y(new_n11570));
  or_6   g09222(.A(new_n9676), .B(pi594), .Y(new_n11571));
  nand_5 g09223(.A(new_n9699), .B(new_n9677), .Y(new_n11572));
  nand_5 g09224(.A(new_n11572), .B(new_n11571), .Y(new_n11573));
  and_6  g09225(.A(new_n11573), .B(new_n11570), .Y(new_n11574));
  nor_5  g09226(.A(new_n11573), .B(new_n11570), .Y(new_n11575));
  nor_5  g09227(.A(new_n11575), .B(pi817), .Y(new_n11576));
  nor_5  g09228(.A(new_n11576), .B(new_n11574), .Y(new_n11577));
  nand_5 g09229(.A(new_n11577), .B(pi808), .Y(new_n11578));
  xor_4  g09230(.A(new_n11545), .B(new_n11539), .Y(new_n11579));
  not_8  g09231(.A(pi808), .Y(new_n11580));
  xor_4  g09232(.A(new_n11577), .B(new_n11580), .Y(new_n11581));
  or_6   g09233(.A(new_n11581), .B(new_n11579), .Y(new_n11582));
  nand_5 g09234(.A(new_n11582), .B(new_n11578), .Y(new_n11583));
  nand_5 g09235(.A(new_n11583), .B(new_n11569), .Y(new_n11584));
  nand_5 g09236(.A(new_n11584), .B(new_n11567), .Y(new_n11585));
  nand_5 g09237(.A(new_n11585), .B(pi525), .Y(new_n11586));
  xor_4  g09238(.A(new_n11549), .B(new_n11534), .Y(new_n11587));
  not_8  g09239(.A(pi525), .Y(new_n11588));
  xor_4  g09240(.A(new_n11585), .B(new_n11588), .Y(new_n11589));
  or_6   g09241(.A(new_n11589), .B(new_n11587), .Y(new_n11590));
  nand_5 g09242(.A(new_n11590), .B(new_n11586), .Y(new_n11591));
  nand_5 g09243(.A(new_n11591), .B(new_n11564), .Y(new_n11592));
  not_8  g09244(.A(new_n11592), .Y(new_n11593));
  not_8  g09245(.A(pi243), .Y(new_n11594));
  xor_4  g09246(.A(new_n11591), .B(new_n11563), .Y(new_n11595));
  nor_5  g09247(.A(new_n11595), .B(new_n11594), .Y(new_n11596));
  nor_5  g09248(.A(new_n11596), .B(new_n11593), .Y(new_n11597));
  xor_4  g09249(.A(new_n11597), .B(new_n11562), .Y(new_n11598));
  xor_4  g09250(.A(new_n11598), .B(new_n11524), .Y(new_n11599));
  not_8  g09251(.A(new_n11599), .Y(new_n11600));
  xor_4  g09252(.A(new_n11583), .B(new_n11569), .Y(new_n11601));
  xor_4  g09253(.A(new_n11518), .B(new_n11515), .Y(new_n11602));
  nand_5 g09254(.A(new_n11602), .B(new_n11601), .Y(new_n11603));
  xor_4  g09255(.A(new_n11581), .B(new_n11579), .Y(new_n11604));
  nor_5  g09256(.A(new_n9700), .B(new_n9657), .Y(new_n11605));
  nor_5  g09257(.A(new_n9724), .B(new_n9702), .Y(new_n11606));
  nor_5  g09258(.A(new_n11606), .B(new_n11605), .Y(new_n11607));
  nand_5 g09259(.A(new_n11607), .B(new_n10990), .Y(new_n11608));
  not_8  g09260(.A(pi817), .Y(new_n11609));
  nor_5  g09261(.A(new_n11575), .B(new_n11574), .Y(new_n11610));
  xor_4  g09262(.A(new_n11610), .B(new_n11609), .Y(new_n11611));
  xnor_4 g09263(.A(new_n11607), .B(new_n10990), .Y(new_n11612));
  or_6   g09264(.A(new_n11612), .B(new_n11611), .Y(new_n11613));
  nand_5 g09265(.A(new_n11613), .B(new_n11608), .Y(new_n11614));
  nand_5 g09266(.A(new_n11614), .B(new_n11604), .Y(new_n11615));
  xnor_4 g09267(.A(new_n11614), .B(new_n11604), .Y(new_n11616));
  or_6   g09268(.A(new_n11616), .B(new_n11076), .Y(new_n11617));
  nand_5 g09269(.A(new_n11617), .B(new_n11615), .Y(new_n11618));
  xor_4  g09270(.A(new_n11602), .B(new_n11601), .Y(new_n11619));
  nand_5 g09271(.A(new_n11619), .B(new_n11618), .Y(new_n11620));
  nand_5 g09272(.A(new_n11620), .B(new_n11603), .Y(new_n11621));
  nor_5  g09273(.A(new_n11510), .B(new_n11508), .Y(new_n11622));
  xor_4  g09274(.A(new_n11622), .B(new_n11520), .Y(new_n11623));
  or_6   g09275(.A(new_n11623), .B(new_n11621), .Y(new_n11624));
  xor_4  g09276(.A(new_n11623), .B(new_n11621), .Y(new_n11625));
  not_8  g09277(.A(new_n11587), .Y(new_n11626));
  xor_4  g09278(.A(new_n11589), .B(new_n11626), .Y(new_n11627));
  nand_5 g09279(.A(new_n11627), .B(new_n11625), .Y(new_n11628));
  nand_5 g09280(.A(new_n11628), .B(new_n11624), .Y(new_n11629));
  nand_5 g09281(.A(new_n11503), .B(new_n11501), .Y(new_n11630));
  xor_4  g09282(.A(new_n11630), .B(new_n11522), .Y(new_n11631));
  nand_5 g09283(.A(new_n11631), .B(new_n11629), .Y(new_n11632));
  not_8  g09284(.A(new_n11632), .Y(new_n11633));
  xor_4  g09285(.A(new_n11631), .B(new_n11629), .Y(new_n11634));
  not_8  g09286(.A(new_n11634), .Y(new_n11635));
  xor_4  g09287(.A(new_n11595), .B(new_n11594), .Y(new_n11636));
  nor_5  g09288(.A(new_n11636), .B(new_n11635), .Y(new_n11637));
  nor_5  g09289(.A(new_n11637), .B(new_n11633), .Y(new_n11638));
  xor_4  g09290(.A(new_n11638), .B(new_n11600), .Y(po0075));
  not_8  g09291(.A(new_n4320), .Y(new_n11640));
  nand_5 g09292(.A(new_n11640), .B(pi490), .Y(new_n11641));
  xor_4  g09293(.A(new_n4320), .B(new_n6380), .Y(new_n11642));
  not_8  g09294(.A(new_n4304), .Y(new_n11643));
  nand_5 g09295(.A(new_n4055), .B(pi433), .Y(new_n11644));
  nand_5 g09296(.A(new_n11644), .B(new_n4056), .Y(new_n11645));
  nand_5 g09297(.A(new_n11645), .B(new_n11643), .Y(new_n11646));
  xor_4  g09298(.A(new_n11645), .B(new_n4304), .Y(new_n11647));
  or_6   g09299(.A(new_n11647), .B(new_n6221), .Y(new_n11648));
  nand_5 g09300(.A(new_n11648), .B(new_n11646), .Y(new_n11649));
  or_6   g09301(.A(new_n11649), .B(new_n4441), .Y(new_n11650));
  nand_5 g09302(.A(new_n11649), .B(new_n4441), .Y(new_n11651));
  nand_5 g09303(.A(new_n11651), .B(new_n6259), .Y(new_n11652));
  nand_5 g09304(.A(new_n11652), .B(new_n11650), .Y(new_n11653));
  and_6  g09305(.A(new_n11653), .B(new_n4317), .Y(new_n11654));
  nor_5  g09306(.A(new_n11653), .B(new_n4317), .Y(new_n11655));
  nor_5  g09307(.A(new_n11655), .B(pi789), .Y(new_n11656));
  nor_5  g09308(.A(new_n11656), .B(new_n11654), .Y(new_n11657));
  nand_5 g09309(.A(new_n11657), .B(new_n11642), .Y(new_n11658));
  nand_5 g09310(.A(new_n11658), .B(new_n11641), .Y(new_n11659));
  nand_5 g09311(.A(new_n11659), .B(new_n4278), .Y(new_n11660));
  not_8  g09312(.A(new_n11660), .Y(new_n11661));
  nand_5 g09313(.A(new_n6318), .B(pi135), .Y(new_n11662));
  xor_4  g09314(.A(new_n6318), .B(pi135), .Y(new_n11663));
  xor_4  g09315(.A(new_n6246), .B(pi054), .Y(new_n11664));
  not_8  g09316(.A(new_n11664), .Y(new_n11665));
  nand_5 g09317(.A(new_n6248), .B(new_n11071), .Y(new_n11666));
  nand_5 g09318(.A(new_n6247), .B(pi113), .Y(new_n11667));
  nand_5 g09319(.A(pi819), .B(new_n6237), .Y(new_n11668));
  xor_4  g09320(.A(pi819), .B(new_n6237), .Y(new_n11669));
  not_8  g09321(.A(new_n11669), .Y(new_n11670));
  not_8  g09322(.A(pi133), .Y(new_n11671));
  nand_5 g09323(.A(pi479), .B(new_n11671), .Y(new_n11672));
  xor_4  g09324(.A(pi479), .B(new_n11671), .Y(new_n11673));
  not_8  g09325(.A(pi371), .Y(new_n11674));
  nand_5 g09326(.A(new_n11674), .B(pi058), .Y(new_n11675));
  not_8  g09327(.A(new_n11675), .Y(new_n11676));
  xor_4  g09328(.A(pi371), .B(new_n3944), .Y(new_n11677));
  not_8  g09329(.A(new_n11677), .Y(new_n11678));
  nand_5 g09330(.A(pi824), .B(new_n3949), .Y(new_n11679));
  not_8  g09331(.A(pi824), .Y(new_n11680));
  nand_5 g09332(.A(new_n11680), .B(pi305), .Y(new_n11681));
  nand_5 g09333(.A(new_n9651), .B(pi350), .Y(new_n11682));
  nand_5 g09334(.A(new_n11682), .B(new_n11681), .Y(new_n11683));
  nand_5 g09335(.A(new_n11683), .B(new_n11679), .Y(new_n11684));
  nor_5  g09336(.A(new_n11684), .B(new_n11678), .Y(new_n11685));
  nor_5  g09337(.A(new_n11685), .B(new_n11676), .Y(new_n11686));
  not_8  g09338(.A(new_n11686), .Y(new_n11687));
  nand_5 g09339(.A(new_n11687), .B(new_n11673), .Y(new_n11688));
  nand_5 g09340(.A(new_n11688), .B(new_n11672), .Y(new_n11689));
  or_6   g09341(.A(new_n11689), .B(new_n11670), .Y(new_n11690));
  nand_5 g09342(.A(new_n11690), .B(new_n11668), .Y(new_n11691));
  nand_5 g09343(.A(new_n11691), .B(new_n6244), .Y(new_n11692));
  nand_5 g09344(.A(new_n11692), .B(new_n11667), .Y(new_n11693));
  nand_5 g09345(.A(new_n11693), .B(new_n11666), .Y(new_n11694));
  and_6  g09346(.A(new_n11694), .B(new_n11665), .Y(new_n11695));
  nor_5  g09347(.A(new_n11694), .B(pi054), .Y(new_n11696));
  or_6   g09348(.A(new_n11696), .B(new_n11695), .Y(new_n11697));
  or_6   g09349(.A(new_n11697), .B(new_n11512), .Y(new_n11698));
  nand_5 g09350(.A(new_n11696), .B(new_n6246), .Y(new_n11699));
  nand_5 g09351(.A(new_n11699), .B(new_n11698), .Y(new_n11700));
  nand_5 g09352(.A(new_n11700), .B(new_n11663), .Y(new_n11701));
  nand_5 g09353(.A(new_n11701), .B(new_n11662), .Y(new_n11702));
  not_8  g09354(.A(new_n11702), .Y(new_n11703));
  nand_5 g09355(.A(new_n6354), .B(new_n11499), .Y(new_n11704));
  nand_5 g09356(.A(new_n11704), .B(new_n6357), .Y(new_n11705));
  nand_5 g09357(.A(new_n11705), .B(new_n11703), .Y(new_n11706));
  nand_5 g09358(.A(new_n11499), .B(pi110), .Y(new_n11707));
  nand_5 g09359(.A(new_n11707), .B(new_n11706), .Y(new_n11708));
  not_8  g09360(.A(new_n11708), .Y(new_n11709));
  xor_4  g09361(.A(new_n11697), .B(pi598), .Y(new_n11710));
  xor_4  g09362(.A(new_n11686), .B(new_n11673), .Y(new_n11711));
  xor_4  g09363(.A(new_n11684), .B(new_n11678), .Y(new_n11712));
  xor_4  g09364(.A(pi821), .B(pi350), .Y(new_n11713));
  or_6   g09365(.A(new_n11713), .B(new_n10992), .Y(new_n11714));
  nand_5 g09366(.A(new_n11713), .B(new_n10992), .Y(new_n11715));
  nand_5 g09367(.A(new_n2570), .B(new_n10996), .Y(new_n11716));
  nand_5 g09368(.A(new_n11716), .B(new_n11715), .Y(new_n11717));
  nand_5 g09369(.A(new_n11717), .B(new_n11714), .Y(new_n11718));
  and_6  g09370(.A(new_n11681), .B(new_n11679), .Y(new_n11719));
  xor_4  g09371(.A(new_n11719), .B(new_n11682), .Y(new_n11720));
  not_8  g09372(.A(new_n11720), .Y(new_n11721));
  nand_5 g09373(.A(new_n11721), .B(new_n11718), .Y(new_n11722));
  xor_4  g09374(.A(new_n11720), .B(new_n11718), .Y(new_n11723));
  or_6   g09375(.A(new_n11723), .B(new_n10995), .Y(new_n11724));
  nand_5 g09376(.A(new_n11724), .B(new_n11722), .Y(new_n11725));
  and_6  g09377(.A(new_n11725), .B(new_n11712), .Y(new_n11726));
  nor_5  g09378(.A(new_n11725), .B(new_n11712), .Y(new_n11727));
  nor_5  g09379(.A(new_n11727), .B(new_n10993), .Y(new_n11728));
  nor_5  g09380(.A(new_n11728), .B(new_n11726), .Y(new_n11729));
  or_6   g09381(.A(new_n11729), .B(new_n11711), .Y(new_n11730));
  xor_4  g09382(.A(new_n11729), .B(new_n11711), .Y(new_n11731));
  nand_5 g09383(.A(new_n11731), .B(pi767), .Y(new_n11732));
  nand_5 g09384(.A(new_n11732), .B(new_n11730), .Y(new_n11733));
  xor_4  g09385(.A(new_n11689), .B(new_n11669), .Y(new_n11734));
  or_6   g09386(.A(new_n11734), .B(new_n11733), .Y(new_n11735));
  nand_5 g09387(.A(new_n11735), .B(pi043), .Y(new_n11736));
  nand_5 g09388(.A(new_n11734), .B(new_n11733), .Y(new_n11737));
  nand_5 g09389(.A(new_n11737), .B(new_n11736), .Y(new_n11738));
  nand_5 g09390(.A(new_n11738), .B(pi015), .Y(new_n11739));
  xor_4  g09391(.A(new_n11738), .B(new_n11077), .Y(new_n11740));
  xor_4  g09392(.A(new_n6248), .B(pi113), .Y(new_n11741));
  xor_4  g09393(.A(new_n11741), .B(new_n11692), .Y(new_n11742));
  or_6   g09394(.A(new_n11742), .B(new_n11740), .Y(new_n11743));
  nand_5 g09395(.A(new_n11743), .B(new_n11739), .Y(new_n11744));
  or_6   g09396(.A(new_n11744), .B(new_n11710), .Y(new_n11745));
  nand_5 g09397(.A(new_n11745), .B(pi069), .Y(new_n11746));
  nand_5 g09398(.A(new_n11744), .B(new_n11710), .Y(new_n11747));
  nand_5 g09399(.A(new_n11747), .B(new_n11746), .Y(new_n11748));
  nand_5 g09400(.A(new_n11748), .B(pi415), .Y(new_n11749));
  nor_5  g09401(.A(new_n11748), .B(pi415), .Y(new_n11750));
  xor_4  g09402(.A(new_n11700), .B(new_n11663), .Y(new_n11751));
  or_6   g09403(.A(new_n11751), .B(new_n11750), .Y(new_n11752));
  nand_5 g09404(.A(new_n11752), .B(new_n11749), .Y(new_n11753));
  nor_5  g09405(.A(new_n11753), .B(pi736), .Y(new_n11754));
  nand_5 g09406(.A(new_n11754), .B(new_n11709), .Y(new_n11755));
  not_8  g09407(.A(new_n11755), .Y(new_n11756));
  nor_5  g09408(.A(new_n11705), .B(new_n11703), .Y(new_n11757));
  not_8  g09409(.A(new_n6356), .Y(new_n11758));
  xor_4  g09410(.A(new_n11702), .B(pi148), .Y(new_n11759));
  nand_5 g09411(.A(new_n11759), .B(new_n11758), .Y(new_n11760));
  not_8  g09412(.A(new_n11760), .Y(new_n11761));
  nor_5  g09413(.A(new_n11761), .B(new_n11757), .Y(new_n11762));
  nand_5 g09414(.A(new_n11753), .B(pi736), .Y(new_n11763));
  not_8  g09415(.A(new_n11763), .Y(new_n11764));
  nor_5  g09416(.A(new_n11764), .B(new_n11762), .Y(new_n11765));
  nor_5  g09417(.A(new_n11765), .B(new_n11756), .Y(new_n11766));
  xor_4  g09418(.A(new_n11766), .B(new_n11661), .Y(new_n11767));
  xor_4  g09419(.A(new_n11659), .B(new_n4278), .Y(new_n11768));
  nor_5  g09420(.A(new_n11763), .B(new_n11709), .Y(new_n11769));
  not_8  g09421(.A(new_n6357), .Y(new_n11770));
  nand_5 g09422(.A(new_n11770), .B(new_n11499), .Y(new_n11771));
  nor_5  g09423(.A(new_n11771), .B(new_n11702), .Y(new_n11772));
  nor_5  g09424(.A(new_n11772), .B(new_n11769), .Y(new_n11773));
  or_6   g09425(.A(new_n11773), .B(new_n11754), .Y(new_n11774));
  and_6  g09426(.A(new_n11774), .B(new_n11766), .Y(new_n11775));
  nand_5 g09427(.A(new_n11775), .B(new_n11768), .Y(new_n11776));
  xor_4  g09428(.A(new_n11657), .B(new_n11642), .Y(new_n11777));
  nor_5  g09429(.A(new_n11764), .B(new_n11754), .Y(new_n11778));
  not_8  g09430(.A(new_n6358), .Y(new_n11779));
  xor_4  g09431(.A(new_n11759), .B(new_n11779), .Y(new_n11780));
  xor_4  g09432(.A(new_n11780), .B(new_n11778), .Y(new_n11781));
  nor_5  g09433(.A(new_n11781), .B(new_n11777), .Y(new_n11782));
  nor_5  g09434(.A(new_n11655), .B(new_n11654), .Y(new_n11783));
  xor_4  g09435(.A(new_n11783), .B(new_n6295), .Y(new_n11784));
  xor_4  g09436(.A(new_n11748), .B(pi415), .Y(new_n11785));
  xor_4  g09437(.A(new_n11785), .B(new_n11751), .Y(new_n11786));
  not_8  g09438(.A(new_n11786), .Y(new_n11787));
  or_6   g09439(.A(new_n11787), .B(new_n11784), .Y(new_n11788));
  not_8  g09440(.A(pi069), .Y(new_n11789));
  nand_5 g09441(.A(new_n11747), .B(new_n11745), .Y(new_n11790));
  xor_4  g09442(.A(new_n11790), .B(new_n11789), .Y(new_n11791));
  nand_5 g09443(.A(new_n11651), .B(new_n11650), .Y(new_n11792));
  xor_4  g09444(.A(new_n11792), .B(new_n6259), .Y(new_n11793));
  not_8  g09445(.A(new_n11793), .Y(new_n11794));
  or_6   g09446(.A(new_n11794), .B(new_n11791), .Y(new_n11795));
  xor_4  g09447(.A(new_n11647), .B(pi707), .Y(new_n11796));
  xor_4  g09448(.A(new_n11742), .B(new_n11740), .Y(new_n11797));
  nor_5  g09449(.A(new_n11797), .B(new_n11796), .Y(new_n11798));
  xnor_4 g09450(.A(new_n11797), .B(new_n11796), .Y(new_n11799));
  nand_5 g09451(.A(new_n11737), .B(new_n11735), .Y(new_n11800));
  xor_4  g09452(.A(new_n11800), .B(new_n11021), .Y(new_n11801));
  nand_5 g09453(.A(new_n11801), .B(new_n4058), .Y(new_n11802));
  xor_4  g09454(.A(new_n11801), .B(new_n4059), .Y(new_n11803));
  xor_4  g09455(.A(new_n11731), .B(pi767), .Y(new_n11804));
  and_6  g09456(.A(new_n11804), .B(new_n3943), .Y(new_n11805));
  xor_4  g09457(.A(new_n11804), .B(new_n3942), .Y(new_n11806));
  nor_5  g09458(.A(new_n11727), .B(new_n11726), .Y(new_n11807));
  xor_4  g09459(.A(new_n11807), .B(new_n10993), .Y(new_n11808));
  nand_5 g09460(.A(new_n11808), .B(new_n4006), .Y(new_n11809));
  xnor_4 g09461(.A(new_n11808), .B(new_n4006), .Y(new_n11810));
  not_8  g09462(.A(new_n4011), .Y(new_n11811));
  xor_4  g09463(.A(new_n11723), .B(pi169), .Y(new_n11812));
  nor_5  g09464(.A(new_n11812), .B(new_n11811), .Y(new_n11813));
  xor_4  g09465(.A(new_n11045), .B(pi606), .Y(new_n11814));
  nor_5  g09466(.A(new_n11814), .B(new_n2567), .Y(new_n11815));
  and_6  g09467(.A(new_n11814), .B(new_n7244), .Y(new_n11816));
  nor_5  g09468(.A(new_n11816), .B(new_n11815), .Y(new_n11817));
  nand_5 g09469(.A(new_n11715), .B(new_n11714), .Y(new_n11818));
  not_8  g09470(.A(new_n2567), .Y(new_n11819));
  nor_5  g09471(.A(new_n11819), .B(new_n7244), .Y(new_n11820));
  or_6   g09472(.A(new_n11820), .B(new_n11716), .Y(new_n11821));
  nand_5 g09473(.A(new_n11817), .B(new_n11716), .Y(new_n11822));
  nand_5 g09474(.A(new_n11822), .B(new_n11821), .Y(new_n11823));
  xor_4  g09475(.A(new_n11823), .B(new_n11818), .Y(new_n11824));
  not_8  g09476(.A(new_n11824), .Y(new_n11825));
  nor_5  g09477(.A(new_n11825), .B(new_n11817), .Y(new_n11826));
  and_6  g09478(.A(new_n11825), .B(new_n4016), .Y(new_n11827));
  nor_5  g09479(.A(new_n11827), .B(new_n11826), .Y(new_n11828));
  xor_4  g09480(.A(new_n11812), .B(new_n4011), .Y(new_n11829));
  nor_5  g09481(.A(new_n11829), .B(new_n11828), .Y(new_n11830));
  or_6   g09482(.A(new_n11830), .B(new_n11813), .Y(new_n11831));
  or_6   g09483(.A(new_n11831), .B(new_n11810), .Y(new_n11832));
  nand_5 g09484(.A(new_n11832), .B(new_n11809), .Y(new_n11833));
  nor_5  g09485(.A(new_n11833), .B(new_n11806), .Y(new_n11834));
  nor_5  g09486(.A(new_n11834), .B(new_n11805), .Y(new_n11835));
  or_6   g09487(.A(new_n11835), .B(new_n11803), .Y(new_n11836));
  nand_5 g09488(.A(new_n11836), .B(new_n11802), .Y(new_n11837));
  nor_5  g09489(.A(new_n11837), .B(new_n11799), .Y(new_n11838));
  nor_5  g09490(.A(new_n11838), .B(new_n11798), .Y(new_n11839));
  not_8  g09491(.A(new_n11839), .Y(new_n11840));
  xor_4  g09492(.A(new_n11794), .B(new_n11791), .Y(new_n11841));
  nand_5 g09493(.A(new_n11841), .B(new_n11840), .Y(new_n11842));
  nand_5 g09494(.A(new_n11842), .B(new_n11795), .Y(new_n11843));
  xor_4  g09495(.A(new_n11786), .B(new_n11784), .Y(new_n11844));
  not_8  g09496(.A(new_n11844), .Y(new_n11845));
  nand_5 g09497(.A(new_n11845), .B(new_n11843), .Y(new_n11846));
  nand_5 g09498(.A(new_n11846), .B(new_n11788), .Y(new_n11847));
  not_8  g09499(.A(new_n11777), .Y(new_n11848));
  xor_4  g09500(.A(new_n11781), .B(new_n11848), .Y(new_n11849));
  nor_5  g09501(.A(new_n11849), .B(new_n11847), .Y(new_n11850));
  or_6   g09502(.A(new_n11850), .B(new_n11782), .Y(new_n11851));
  not_8  g09503(.A(new_n11851), .Y(new_n11852));
  xor_4  g09504(.A(new_n11775), .B(new_n11768), .Y(new_n11853));
  nand_5 g09505(.A(new_n11853), .B(new_n11852), .Y(new_n11854));
  nand_5 g09506(.A(new_n11854), .B(new_n11776), .Y(new_n11855));
  xor_4  g09507(.A(new_n11855), .B(new_n11767), .Y(po0076));
  not_8  g09508(.A(new_n3888), .Y(new_n11857));
  xor_4  g09509(.A(new_n3889), .B(new_n11857), .Y(po0077));
  xor_4  g09510(.A(new_n4503), .B(new_n4501), .Y(po0078));
  or_6   g09511(.A(new_n9064), .B(new_n9062), .Y(new_n11860));
  nor_5  g09512(.A(new_n9168), .B(new_n9068), .Y(new_n11861));
  nand_5 g09513(.A(new_n11861), .B(new_n9199), .Y(new_n11862));
  nand_5 g09514(.A(new_n11862), .B(new_n9195), .Y(new_n11863));
  not_8  g09515(.A(new_n11863), .Y(new_n11864));
  nor_5  g09516(.A(new_n11864), .B(new_n11860), .Y(po0079));
  xor_4  g09517(.A(new_n4033), .B(new_n4015), .Y(po0080));
  xor_4  g09518(.A(new_n3344), .B(new_n3343), .Y(po0081));
  not_8  g09519(.A(new_n7786), .Y(new_n11868));
  nand_5 g09520(.A(new_n11868), .B(new_n9002), .Y(new_n11869));
  nand_5 g09521(.A(new_n7873), .B(new_n7787), .Y(new_n11870));
  nand_5 g09522(.A(new_n11870), .B(new_n11869), .Y(new_n11871));
  xor_4  g09523(.A(pi430), .B(pi142), .Y(new_n11872));
  nand_5 g09524(.A(new_n11351), .B(new_n11348), .Y(new_n11873));
  nand_5 g09525(.A(new_n11873), .B(new_n11350), .Y(new_n11874));
  xor_4  g09526(.A(new_n11874), .B(new_n11872), .Y(new_n11875));
  or_6   g09527(.A(new_n11875), .B(new_n7971), .Y(new_n11876));
  nor_5  g09528(.A(new_n11353), .B(new_n7875), .Y(new_n11877));
  and_6  g09529(.A(new_n11354), .B(new_n11344), .Y(new_n11878));
  nor_5  g09530(.A(new_n11878), .B(new_n11877), .Y(new_n11879));
  xor_4  g09531(.A(new_n11875), .B(new_n7972), .Y(new_n11880));
  or_6   g09532(.A(new_n11880), .B(new_n11879), .Y(new_n11881));
  nand_5 g09533(.A(new_n11881), .B(new_n11876), .Y(new_n11882));
  nand_5 g09534(.A(new_n5451), .B(pi142), .Y(new_n11883));
  not_8  g09535(.A(new_n11883), .Y(new_n11884));
  nor_5  g09536(.A(new_n11874), .B(new_n11872), .Y(new_n11885));
  nor_5  g09537(.A(new_n11885), .B(new_n11884), .Y(new_n11886));
  or_6   g09538(.A(new_n11886), .B(new_n7874), .Y(new_n11887));
  nor_5  g09539(.A(new_n11887), .B(new_n11882), .Y(new_n11888));
  nor_5  g09540(.A(new_n11888), .B(new_n11871), .Y(new_n11889));
  not_8  g09541(.A(new_n11871), .Y(new_n11890));
  not_8  g09542(.A(new_n11882), .Y(new_n11891));
  nand_5 g09543(.A(new_n11886), .B(new_n7874), .Y(new_n11892));
  nor_5  g09544(.A(new_n11892), .B(new_n11891), .Y(new_n11893));
  nor_5  g09545(.A(new_n11893), .B(new_n11890), .Y(new_n11894));
  nor_5  g09546(.A(new_n11894), .B(new_n11889), .Y(po0082));
  xor_4  g09547(.A(new_n6911), .B(new_n6904), .Y(po0083));
  xor_4  g09548(.A(pi323), .B(pi068), .Y(new_n11897));
  nand_5 g09549(.A(pi775), .B(pi556), .Y(new_n11898));
  not_8  g09550(.A(pi349), .Y(new_n11899));
  nand_5 g09551(.A(pi809), .B(pi555), .Y(new_n11900));
  not_8  g09552(.A(pi809), .Y(new_n11901));
  nand_5 g09553(.A(new_n11901), .B(new_n6953), .Y(new_n11902));
  nand_5 g09554(.A(pi667), .B(pi583), .Y(new_n11903));
  nand_5 g09555(.A(new_n6957), .B(new_n4724), .Y(new_n11904));
  nand_5 g09556(.A(pi695), .B(pi566), .Y(new_n11905));
  nand_5 g09557(.A(new_n3712), .B(new_n6960), .Y(new_n11906));
  nand_5 g09558(.A(pi805), .B(pi145), .Y(new_n11907));
  nand_5 g09559(.A(new_n3716), .B(new_n6963), .Y(new_n11908));
  nand_5 g09560(.A(pi454), .B(pi006), .Y(new_n11909));
  xor_4  g09561(.A(pi454), .B(pi006), .Y(new_n11910));
  nand_5 g09562(.A(pi818), .B(pi731), .Y(new_n11911));
  xor_4  g09563(.A(pi818), .B(pi731), .Y(new_n11912));
  nor_5  g09564(.A(pi270), .B(pi158), .Y(new_n11913));
  nand_5 g09565(.A(pi367), .B(pi259), .Y(new_n11914));
  not_8  g09566(.A(new_n11914), .Y(new_n11915));
  xor_4  g09567(.A(pi270), .B(new_n3728), .Y(new_n11916));
  nor_5  g09568(.A(new_n11916), .B(new_n11915), .Y(new_n11917));
  nor_5  g09569(.A(new_n11917), .B(new_n11913), .Y(new_n11918));
  nand_5 g09570(.A(new_n11918), .B(new_n11912), .Y(new_n11919));
  nand_5 g09571(.A(new_n11919), .B(new_n11911), .Y(new_n11920));
  nand_5 g09572(.A(new_n11920), .B(new_n11910), .Y(new_n11921));
  nand_5 g09573(.A(new_n11921), .B(new_n11909), .Y(new_n11922));
  nand_5 g09574(.A(new_n11922), .B(new_n11908), .Y(new_n11923));
  nand_5 g09575(.A(new_n11923), .B(new_n11907), .Y(new_n11924));
  nand_5 g09576(.A(new_n11924), .B(new_n11906), .Y(new_n11925));
  nand_5 g09577(.A(new_n11925), .B(new_n11905), .Y(new_n11926));
  nand_5 g09578(.A(new_n11926), .B(new_n11904), .Y(new_n11927));
  nand_5 g09579(.A(new_n11927), .B(new_n11903), .Y(new_n11928));
  nand_5 g09580(.A(new_n11928), .B(new_n11902), .Y(new_n11929));
  nand_5 g09581(.A(new_n11929), .B(new_n11900), .Y(new_n11930));
  nand_5 g09582(.A(new_n11930), .B(new_n11899), .Y(new_n11931));
  nand_5 g09583(.A(new_n11931), .B(new_n11898), .Y(new_n11932));
  not_8  g09584(.A(new_n11932), .Y(new_n11933));
  not_8  g09585(.A(pi556), .Y(new_n11934));
  nand_5 g09586(.A(new_n7181), .B(new_n11934), .Y(new_n11935));
  nand_5 g09587(.A(new_n11935), .B(new_n11898), .Y(new_n11936));
  nor_5  g09588(.A(new_n11930), .B(new_n11899), .Y(new_n11937));
  not_8  g09589(.A(new_n11937), .Y(new_n11938));
  nand_5 g09590(.A(new_n11938), .B(new_n11931), .Y(new_n11939));
  nand_5 g09591(.A(new_n11939), .B(new_n11936), .Y(new_n11940));
  xor_4  g09592(.A(new_n11939), .B(new_n11936), .Y(new_n11941));
  not_8  g09593(.A(new_n11941), .Y(new_n11942));
  nand_5 g09594(.A(new_n11902), .B(new_n11900), .Y(new_n11943));
  xnor_4 g09595(.A(new_n11943), .B(new_n11928), .Y(new_n11944));
  nand_5 g09596(.A(new_n11944), .B(new_n2897), .Y(new_n11945));
  or_6   g09597(.A(new_n11944), .B(new_n2897), .Y(new_n11946));
  xnor_4 g09598(.A(new_n11920), .B(new_n11910), .Y(new_n11947));
  xor_4  g09599(.A(new_n11918), .B(new_n11912), .Y(new_n11948));
  xor_4  g09600(.A(pi367), .B(new_n3730), .Y(new_n11949));
  nand_5 g09601(.A(new_n11949), .B(pi038), .Y(new_n11950));
  xor_4  g09602(.A(new_n11916), .B(new_n11915), .Y(new_n11951));
  nand_5 g09603(.A(new_n11951), .B(pi044), .Y(new_n11952));
  nand_5 g09604(.A(new_n11952), .B(new_n11950), .Y(new_n11953));
  or_6   g09605(.A(new_n11951), .B(pi044), .Y(new_n11954));
  nand_5 g09606(.A(new_n11954), .B(new_n11953), .Y(new_n11955));
  or_6   g09607(.A(new_n11955), .B(new_n11948), .Y(new_n11956));
  nand_5 g09608(.A(new_n11955), .B(new_n11948), .Y(new_n11957));
  nand_5 g09609(.A(new_n11957), .B(pi801), .Y(new_n11958));
  nand_5 g09610(.A(new_n11958), .B(new_n11956), .Y(new_n11959));
  nand_5 g09611(.A(new_n11959), .B(new_n11947), .Y(new_n11960));
  xnor_4 g09612(.A(new_n11959), .B(new_n11947), .Y(new_n11961));
  or_6   g09613(.A(new_n11961), .B(new_n2912), .Y(new_n11962));
  nand_5 g09614(.A(new_n11962), .B(new_n11960), .Y(new_n11963));
  nand_5 g09615(.A(new_n11908), .B(new_n11907), .Y(new_n11964));
  xor_4  g09616(.A(new_n11964), .B(new_n11922), .Y(new_n11965));
  nand_5 g09617(.A(new_n11965), .B(new_n11963), .Y(new_n11966));
  xnor_4 g09618(.A(new_n11965), .B(new_n11963), .Y(new_n11967));
  or_6   g09619(.A(new_n11967), .B(new_n2909), .Y(new_n11968));
  nand_5 g09620(.A(new_n11968), .B(new_n11966), .Y(new_n11969));
  nand_5 g09621(.A(new_n11906), .B(new_n11905), .Y(new_n11970));
  xor_4  g09622(.A(new_n11970), .B(new_n11924), .Y(new_n11971));
  nand_5 g09623(.A(new_n11971), .B(new_n11969), .Y(new_n11972));
  xor_4  g09624(.A(new_n11971), .B(new_n11969), .Y(new_n11973));
  nand_5 g09625(.A(new_n11973), .B(pi229), .Y(new_n11974));
  nand_5 g09626(.A(new_n11974), .B(new_n11972), .Y(new_n11975));
  nand_5 g09627(.A(new_n11904), .B(new_n11903), .Y(new_n11976));
  xor_4  g09628(.A(new_n11976), .B(new_n11926), .Y(new_n11977));
  or_6   g09629(.A(new_n11977), .B(new_n11975), .Y(new_n11978));
  xor_4  g09630(.A(new_n11977), .B(new_n11975), .Y(new_n11979));
  nand_5 g09631(.A(new_n11979), .B(new_n2932), .Y(new_n11980));
  nand_5 g09632(.A(new_n11980), .B(new_n11978), .Y(new_n11981));
  nand_5 g09633(.A(new_n11981), .B(new_n11946), .Y(new_n11982));
  nand_5 g09634(.A(new_n11982), .B(new_n11945), .Y(new_n11983));
  nor_5  g09635(.A(new_n11983), .B(new_n11942), .Y(new_n11984));
  not_8  g09636(.A(new_n11984), .Y(new_n11985));
  nand_5 g09637(.A(new_n11985), .B(new_n11940), .Y(new_n11986));
  nand_5 g09638(.A(new_n11986), .B(new_n11933), .Y(new_n11987));
  nand_5 g09639(.A(new_n11938), .B(new_n11935), .Y(new_n11988));
  nor_5  g09640(.A(new_n11988), .B(new_n11933), .Y(new_n11989));
  nand_5 g09641(.A(new_n11989), .B(new_n11985), .Y(new_n11990));
  nand_5 g09642(.A(new_n11990), .B(new_n11987), .Y(new_n11991));
  xor_4  g09643(.A(new_n11991), .B(new_n7187), .Y(new_n11992));
  xor_4  g09644(.A(new_n11992), .B(new_n11897), .Y(new_n11993));
  not_8  g09645(.A(pi661), .Y(new_n11994));
  not_8  g09646(.A(pi185), .Y(new_n11995));
  nand_5 g09647(.A(new_n7314), .B(new_n11995), .Y(new_n11996));
  xor_4  g09648(.A(new_n7314), .B(new_n11995), .Y(new_n11997));
  nand_5 g09649(.A(new_n3843), .B(pi143), .Y(new_n11998));
  nand_5 g09650(.A(new_n11998), .B(new_n3842), .Y(new_n11999));
  nand_5 g09651(.A(new_n11999), .B(new_n7320), .Y(new_n12000));
  not_8  g09652(.A(new_n12000), .Y(new_n12001));
  not_8  g09653(.A(pi382), .Y(new_n12002));
  xor_4  g09654(.A(new_n11999), .B(new_n7321), .Y(new_n12003));
  nor_5  g09655(.A(new_n12003), .B(new_n12002), .Y(new_n12004));
  nor_5  g09656(.A(new_n12004), .B(new_n12001), .Y(new_n12005));
  nand_5 g09657(.A(new_n12005), .B(new_n11997), .Y(new_n12006));
  nand_5 g09658(.A(new_n12006), .B(new_n11996), .Y(new_n12007));
  or_6   g09659(.A(new_n12007), .B(new_n11994), .Y(new_n12008));
  nand_5 g09660(.A(new_n12007), .B(new_n11994), .Y(new_n12009));
  nand_5 g09661(.A(new_n12009), .B(new_n12008), .Y(new_n12010));
  xor_4  g09662(.A(new_n12010), .B(new_n7309), .Y(new_n12011));
  xor_4  g09663(.A(new_n12011), .B(new_n11993), .Y(new_n12012));
  xor_4  g09664(.A(new_n11983), .B(new_n11941), .Y(new_n12013));
  xor_4  g09665(.A(new_n12005), .B(new_n11997), .Y(new_n12014));
  nor_5  g09666(.A(new_n12014), .B(new_n12013), .Y(new_n12015));
  xor_4  g09667(.A(new_n12003), .B(pi382), .Y(new_n12016));
  nand_5 g09668(.A(new_n11946), .B(new_n11945), .Y(new_n12017));
  xor_4  g09669(.A(new_n12017), .B(new_n11981), .Y(new_n12018));
  not_8  g09670(.A(new_n12018), .Y(new_n12019));
  nor_5  g09671(.A(new_n12019), .B(new_n12016), .Y(new_n12020));
  xor_4  g09672(.A(new_n12018), .B(new_n12016), .Y(new_n12021));
  not_8  g09673(.A(new_n3845), .Y(new_n12022));
  xor_4  g09674(.A(new_n11979), .B(pi632), .Y(new_n12023));
  and_6  g09675(.A(new_n12023), .B(new_n12022), .Y(new_n12024));
  xor_4  g09676(.A(new_n12023), .B(new_n3845), .Y(new_n12025));
  xor_4  g09677(.A(new_n11973), .B(pi229), .Y(new_n12026));
  nand_5 g09678(.A(new_n12026), .B(new_n11857), .Y(new_n12027));
  or_6   g09679(.A(new_n12026), .B(new_n11857), .Y(new_n12028));
  xor_4  g09680(.A(new_n11967), .B(new_n2909), .Y(new_n12029));
  nand_5 g09681(.A(new_n12029), .B(new_n3847), .Y(new_n12030));
  xnor_4 g09682(.A(new_n12029), .B(new_n3847), .Y(new_n12031));
  xor_4  g09683(.A(new_n11961), .B(new_n2912), .Y(new_n12032));
  not_8  g09684(.A(new_n12032), .Y(new_n12033));
  nor_5  g09685(.A(new_n12033), .B(new_n3879), .Y(new_n12034));
  xor_4  g09686(.A(new_n12032), .B(new_n3879), .Y(new_n12035));
  nand_5 g09687(.A(new_n11957), .B(new_n11956), .Y(new_n12036));
  xor_4  g09688(.A(new_n12036), .B(pi801), .Y(new_n12037));
  nor_5  g09689(.A(new_n12037), .B(new_n3873), .Y(new_n12038));
  not_8  g09690(.A(new_n3873), .Y(new_n12039));
  xor_4  g09691(.A(new_n12037), .B(new_n12039), .Y(new_n12040));
  xor_4  g09692(.A(new_n11949), .B(pi038), .Y(new_n12041));
  not_8  g09693(.A(new_n12041), .Y(new_n12042));
  nand_5 g09694(.A(new_n12042), .B(new_n3864), .Y(new_n12043));
  nor_5  g09695(.A(new_n11949), .B(pi038), .Y(new_n12044));
  nor_5  g09696(.A(new_n12044), .B(new_n11915), .Y(new_n12045));
  xor_4  g09697(.A(new_n11916), .B(new_n2920), .Y(new_n12046));
  xor_4  g09698(.A(new_n12046), .B(new_n12045), .Y(new_n12047));
  xor_4  g09699(.A(new_n12047), .B(new_n12043), .Y(new_n12048));
  nand_5 g09700(.A(new_n12048), .B(new_n3857), .Y(new_n12049));
  nand_5 g09701(.A(new_n12042), .B(new_n3865), .Y(new_n12050));
  or_6   g09702(.A(new_n12050), .B(new_n12048), .Y(new_n12051));
  nand_5 g09703(.A(new_n12051), .B(new_n12049), .Y(new_n12052));
  nor_5  g09704(.A(new_n12052), .B(new_n12040), .Y(new_n12053));
  nor_5  g09705(.A(new_n12053), .B(new_n12038), .Y(new_n12054));
  nor_5  g09706(.A(new_n12054), .B(new_n12035), .Y(new_n12055));
  nor_5  g09707(.A(new_n12055), .B(new_n12034), .Y(new_n12056));
  or_6   g09708(.A(new_n12056), .B(new_n12031), .Y(new_n12057));
  nand_5 g09709(.A(new_n12057), .B(new_n12030), .Y(new_n12058));
  nand_5 g09710(.A(new_n12058), .B(new_n12028), .Y(new_n12059));
  nand_5 g09711(.A(new_n12059), .B(new_n12027), .Y(new_n12060));
  not_8  g09712(.A(new_n12060), .Y(new_n12061));
  nor_5  g09713(.A(new_n12061), .B(new_n12025), .Y(new_n12062));
  nor_5  g09714(.A(new_n12062), .B(new_n12024), .Y(new_n12063));
  nor_5  g09715(.A(new_n12063), .B(new_n12021), .Y(new_n12064));
  or_6   g09716(.A(new_n12064), .B(new_n12020), .Y(new_n12065));
  xor_4  g09717(.A(new_n12014), .B(new_n12013), .Y(new_n12066));
  and_6  g09718(.A(new_n12066), .B(new_n12065), .Y(new_n12067));
  nor_5  g09719(.A(new_n12067), .B(new_n12015), .Y(new_n12068));
  xnor_4 g09720(.A(new_n12068), .B(new_n12012), .Y(po0084));
  xnor_4 g09721(.A(new_n5174), .B(new_n5146), .Y(po0085));
  nand_5 g09722(.A(new_n8986), .B(new_n5634), .Y(new_n12071));
  not_8  g09723(.A(new_n12071), .Y(new_n12072));
  not_8  g09724(.A(pi666), .Y(new_n12073));
  nand_5 g09725(.A(new_n12073), .B(new_n5636), .Y(new_n12074));
  not_8  g09726(.A(new_n12074), .Y(new_n12075));
  not_8  g09727(.A(new_n6940), .Y(new_n12076));
  nor_5  g09728(.A(new_n6942), .B(new_n12076), .Y(new_n12077));
  nor_5  g09729(.A(new_n12077), .B(new_n12075), .Y(new_n12078));
  nand_5 g09730(.A(pi800), .B(pi282), .Y(new_n12079));
  not_8  g09731(.A(new_n12079), .Y(new_n12080));
  nor_5  g09732(.A(new_n12080), .B(new_n12078), .Y(new_n12081));
  nor_5  g09733(.A(new_n12081), .B(new_n12072), .Y(new_n12082));
  not_8  g09734(.A(new_n12082), .Y(new_n12083));
  nor_5  g09735(.A(new_n12080), .B(new_n12072), .Y(new_n12084));
  xor_4  g09736(.A(new_n12084), .B(new_n12078), .Y(new_n12085));
  not_8  g09737(.A(new_n12085), .Y(new_n12086));
  nand_5 g09738(.A(new_n6832), .B(pi644), .Y(new_n12087));
  nand_5 g09739(.A(new_n6831), .B(new_n6165), .Y(new_n12088));
  nand_5 g09740(.A(new_n6837), .B(pi356), .Y(new_n12089));
  xor_4  g09741(.A(new_n6837), .B(pi356), .Y(new_n12090));
  nand_5 g09742(.A(new_n4118), .B(pi307), .Y(new_n12091));
  not_8  g09743(.A(new_n12091), .Y(new_n12092));
  nand_5 g09744(.A(new_n12092), .B(new_n12090), .Y(new_n12093));
  nand_5 g09745(.A(new_n12093), .B(new_n12089), .Y(new_n12094));
  nor_5  g09746(.A(new_n12094), .B(pi609), .Y(new_n12095));
  not_8  g09747(.A(pi609), .Y(new_n12096));
  xor_4  g09748(.A(new_n12094), .B(new_n12096), .Y(new_n12097));
  nor_5  g09749(.A(new_n12097), .B(new_n4083), .Y(new_n12098));
  or_6   g09750(.A(new_n12098), .B(new_n12095), .Y(new_n12099));
  or_6   g09751(.A(new_n12099), .B(new_n6835), .Y(new_n12100));
  xor_4  g09752(.A(new_n12099), .B(new_n6835), .Y(new_n12101));
  nand_5 g09753(.A(new_n12101), .B(pi147), .Y(new_n12102));
  nand_5 g09754(.A(new_n12102), .B(new_n12100), .Y(new_n12103));
  nand_5 g09755(.A(new_n12103), .B(new_n12088), .Y(new_n12104));
  nand_5 g09756(.A(new_n12104), .B(new_n12087), .Y(new_n12105));
  or_6   g09757(.A(new_n12105), .B(new_n6856), .Y(new_n12106));
  nand_5 g09758(.A(new_n12105), .B(new_n6856), .Y(new_n12107));
  nand_5 g09759(.A(new_n12107), .B(new_n6201), .Y(new_n12108));
  nand_5 g09760(.A(new_n12108), .B(new_n12106), .Y(new_n12109));
  nand_5 g09761(.A(new_n12109), .B(new_n6862), .Y(new_n12110));
  xor_4  g09762(.A(new_n12109), .B(new_n6874), .Y(new_n12111));
  or_6   g09763(.A(new_n12111), .B(pi578), .Y(new_n12112));
  nand_5 g09764(.A(new_n12112), .B(new_n12110), .Y(new_n12113));
  or_6   g09765(.A(new_n12113), .B(new_n6828), .Y(new_n12114));
  xor_4  g09766(.A(new_n12113), .B(new_n6828), .Y(new_n12115));
  nand_5 g09767(.A(new_n12115), .B(pi205), .Y(new_n12116));
  nand_5 g09768(.A(new_n12116), .B(new_n12114), .Y(new_n12117));
  or_6   g09769(.A(new_n12117), .B(new_n6943), .Y(new_n12118));
  xor_4  g09770(.A(new_n12117), .B(new_n6943), .Y(new_n12119));
  nand_5 g09771(.A(new_n12119), .B(new_n6307), .Y(new_n12120));
  nand_5 g09772(.A(new_n12120), .B(new_n12118), .Y(new_n12121));
  nand_5 g09773(.A(new_n12121), .B(new_n12086), .Y(new_n12122));
  or_6   g09774(.A(new_n12121), .B(new_n12086), .Y(new_n12123));
  nand_5 g09775(.A(new_n12123), .B(new_n6373), .Y(new_n12124));
  nand_5 g09776(.A(new_n12124), .B(new_n12122), .Y(new_n12125));
  nand_5 g09777(.A(new_n12125), .B(new_n12083), .Y(new_n12126));
  nand_5 g09778(.A(new_n12126), .B(new_n11558), .Y(new_n12127));
  nor_5  g09779(.A(new_n12125), .B(new_n12083), .Y(new_n12128));
  nor_5  g09780(.A(new_n12128), .B(new_n11559), .Y(new_n12129));
  nor_5  g09781(.A(new_n12129), .B(new_n12127), .Y(new_n12130));
  nand_5 g09782(.A(new_n12123), .B(new_n12122), .Y(new_n12131));
  xor_4  g09783(.A(new_n12131), .B(pi335), .Y(new_n12132));
  nor_5  g09784(.A(new_n12132), .B(new_n11563), .Y(new_n12133));
  xor_4  g09785(.A(new_n12132), .B(new_n11563), .Y(new_n12134));
  not_8  g09786(.A(new_n12134), .Y(new_n12135));
  xor_4  g09787(.A(new_n12119), .B(pi247), .Y(new_n12136));
  nand_5 g09788(.A(new_n12136), .B(new_n11626), .Y(new_n12137));
  not_8  g09789(.A(new_n12137), .Y(new_n12138));
  xor_4  g09790(.A(new_n12136), .B(new_n11587), .Y(new_n12139));
  xor_4  g09791(.A(new_n12115), .B(new_n8865), .Y(new_n12140));
  nand_5 g09792(.A(new_n12140), .B(new_n11565), .Y(new_n12141));
  xor_4  g09793(.A(new_n12140), .B(new_n11566), .Y(new_n12142));
  not_8  g09794(.A(new_n11579), .Y(new_n12143));
  xor_4  g09795(.A(new_n12111), .B(new_n8868), .Y(new_n12144));
  nor_5  g09796(.A(new_n12144), .B(new_n12143), .Y(new_n12145));
  nand_5 g09797(.A(new_n12106), .B(new_n12107), .Y(new_n12146));
  xor_4  g09798(.A(new_n12146), .B(pi726), .Y(new_n12147));
  and_6  g09799(.A(new_n12147), .B(new_n11570), .Y(new_n12148));
  nand_5 g09800(.A(new_n12088), .B(new_n12087), .Y(new_n12149));
  xor_4  g09801(.A(new_n12149), .B(new_n12103), .Y(new_n12150));
  not_8  g09802(.A(new_n12150), .Y(new_n12151));
  nor_5  g09803(.A(new_n12151), .B(new_n9676), .Y(new_n12152));
  not_8  g09804(.A(new_n9695), .Y(new_n12153));
  xor_4  g09805(.A(new_n12101), .B(new_n8875), .Y(new_n12154));
  or_6   g09806(.A(new_n12154), .B(new_n12153), .Y(new_n12155));
  xor_4  g09807(.A(new_n12154), .B(new_n12153), .Y(new_n12156));
  xor_4  g09808(.A(new_n12097), .B(new_n6894), .Y(new_n12157));
  nor_5  g09809(.A(new_n12157), .B(new_n9688), .Y(new_n12158));
  xor_4  g09810(.A(new_n12157), .B(new_n9689), .Y(new_n12159));
  xor_4  g09811(.A(new_n12090), .B(new_n9682), .Y(new_n12160));
  nand_5 g09812(.A(new_n12092), .B(new_n7251), .Y(new_n12161));
  not_8  g09813(.A(new_n12161), .Y(new_n12162));
  nand_5 g09814(.A(new_n6905), .B(new_n4088), .Y(new_n12163));
  nor_5  g09815(.A(new_n12163), .B(new_n7251), .Y(new_n12164));
  nor_5  g09816(.A(new_n12164), .B(new_n12162), .Y(new_n12165));
  nor_5  g09817(.A(new_n12165), .B(new_n12160), .Y(new_n12166));
  nor_5  g09818(.A(new_n12166), .B(new_n12093), .Y(new_n12167));
  and_6  g09819(.A(new_n12165), .B(new_n12160), .Y(new_n12168));
  nand_5 g09820(.A(new_n12090), .B(new_n9682), .Y(new_n12169));
  nand_5 g09821(.A(new_n12161), .B(new_n12169), .Y(new_n12170));
  nor_5  g09822(.A(new_n12170), .B(new_n12168), .Y(new_n12171));
  nor_5  g09823(.A(new_n12171), .B(new_n12167), .Y(new_n12172));
  nor_5  g09824(.A(new_n12172), .B(new_n12159), .Y(new_n12173));
  nor_5  g09825(.A(new_n12173), .B(new_n12158), .Y(new_n12174));
  nand_5 g09826(.A(new_n12174), .B(new_n12156), .Y(new_n12175));
  nand_5 g09827(.A(new_n12175), .B(new_n12155), .Y(new_n12176));
  xor_4  g09828(.A(new_n12150), .B(new_n9676), .Y(new_n12177));
  nor_5  g09829(.A(new_n12177), .B(new_n12176), .Y(new_n12178));
  nor_5  g09830(.A(new_n12178), .B(new_n12152), .Y(new_n12179));
  not_8  g09831(.A(new_n11570), .Y(new_n12180));
  xor_4  g09832(.A(new_n12147), .B(new_n12180), .Y(new_n12181));
  nor_5  g09833(.A(new_n12181), .B(new_n12179), .Y(new_n12182));
  nor_5  g09834(.A(new_n12182), .B(new_n12148), .Y(new_n12183));
  xor_4  g09835(.A(new_n12144), .B(new_n11579), .Y(new_n12184));
  nor_5  g09836(.A(new_n12184), .B(new_n12183), .Y(new_n12185));
  nor_5  g09837(.A(new_n12185), .B(new_n12145), .Y(new_n12186));
  or_6   g09838(.A(new_n12186), .B(new_n12142), .Y(new_n12187));
  nand_5 g09839(.A(new_n12187), .B(new_n12141), .Y(new_n12188));
  nor_5  g09840(.A(new_n12188), .B(new_n12139), .Y(new_n12189));
  nor_5  g09841(.A(new_n12189), .B(new_n12138), .Y(new_n12190));
  nor_5  g09842(.A(new_n12190), .B(new_n12135), .Y(new_n12191));
  nor_5  g09843(.A(new_n12191), .B(new_n12133), .Y(new_n12192));
  xor_4  g09844(.A(new_n12125), .B(new_n12083), .Y(new_n12193));
  or_6   g09845(.A(new_n12193), .B(new_n11562), .Y(new_n12194));
  nand_5 g09846(.A(new_n12194), .B(new_n12127), .Y(new_n12195));
  xor_4  g09847(.A(new_n12193), .B(new_n11561), .Y(new_n12196));
  not_8  g09848(.A(new_n12192), .Y(new_n12197));
  nor_5  g09849(.A(new_n12082), .B(new_n11558), .Y(new_n12198));
  nor_5  g09850(.A(new_n12198), .B(new_n12130), .Y(new_n12199));
  xor_4  g09851(.A(new_n12199), .B(new_n12197), .Y(new_n12200));
  nand_5 g09852(.A(new_n12200), .B(new_n12196), .Y(new_n12201));
  nand_5 g09853(.A(new_n12201), .B(new_n12195), .Y(po0915));
  nor_5  g09854(.A(po0915), .B(new_n12192), .Y(new_n12203));
  nor_5  g09855(.A(new_n12203), .B(new_n12130), .Y(po0086));
  xor_4  g09856(.A(new_n5383), .B(new_n10229), .Y(new_n12205));
  or_6   g09857(.A(new_n5320), .B(new_n8767), .Y(new_n12206));
  xor_4  g09858(.A(new_n5320), .B(new_n8767), .Y(new_n12207));
  nor_5  g09859(.A(new_n5325), .B(new_n8770), .Y(new_n12208));
  nand_5 g09860(.A(new_n5331), .B(pi273), .Y(new_n12209));
  xor_4  g09861(.A(new_n5331), .B(new_n8773), .Y(new_n12210));
  or_6   g09862(.A(new_n5335), .B(new_n10239), .Y(new_n12211));
  nand_5 g09863(.A(new_n5335), .B(new_n10239), .Y(new_n12212));
  nand_5 g09864(.A(new_n5251), .B(new_n8835), .Y(new_n12213));
  nand_5 g09865(.A(new_n5356), .B(pi435), .Y(new_n12214));
  nand_5 g09866(.A(new_n12214), .B(new_n12213), .Y(new_n12215));
  xor_4  g09867(.A(new_n12215), .B(new_n5249), .Y(new_n12216));
  nand_5 g09868(.A(new_n12216), .B(pi401), .Y(new_n12217));
  nand_5 g09869(.A(new_n5372), .B(pi435), .Y(new_n12218));
  nand_5 g09870(.A(new_n12218), .B(new_n12217), .Y(new_n12219));
  nand_5 g09871(.A(new_n12219), .B(new_n12212), .Y(new_n12220));
  nand_5 g09872(.A(new_n12220), .B(new_n12211), .Y(new_n12221));
  not_8  g09873(.A(new_n12221), .Y(new_n12222));
  or_6   g09874(.A(new_n12222), .B(new_n12210), .Y(new_n12223));
  nand_5 g09875(.A(new_n12223), .B(new_n12209), .Y(new_n12224));
  not_8  g09876(.A(new_n12224), .Y(new_n12225));
  xor_4  g09877(.A(new_n5325), .B(pi573), .Y(new_n12226));
  nor_5  g09878(.A(new_n12226), .B(new_n12225), .Y(new_n12227));
  or_6   g09879(.A(new_n12227), .B(new_n12208), .Y(new_n12228));
  nand_5 g09880(.A(new_n12228), .B(new_n12207), .Y(new_n12229));
  nand_5 g09881(.A(new_n12229), .B(new_n12206), .Y(new_n12230));
  xor_4  g09882(.A(new_n12230), .B(new_n12205), .Y(new_n12231));
  not_8  g09883(.A(new_n12231), .Y(new_n12232));
  xor_4  g09884(.A(new_n12226), .B(new_n12224), .Y(new_n12233));
  not_8  g09885(.A(new_n12233), .Y(new_n12234));
  nand_5 g09886(.A(new_n7349), .B(new_n6732), .Y(new_n12235));
  nand_5 g09887(.A(new_n7348), .B(pi333), .Y(new_n12236));
  nand_5 g09888(.A(new_n12236), .B(new_n11356), .Y(new_n12237));
  nand_5 g09889(.A(new_n12237), .B(new_n12235), .Y(new_n12238));
  nand_5 g09890(.A(new_n12238), .B(new_n6726), .Y(new_n12239));
  nor_5  g09891(.A(new_n12238), .B(new_n6726), .Y(new_n12240));
  or_6   g09892(.A(new_n12240), .B(new_n7341), .Y(new_n12241));
  nand_5 g09893(.A(new_n12241), .B(new_n12239), .Y(new_n12242));
  nor_5  g09894(.A(new_n12242), .B(new_n7338), .Y(new_n12243));
  xor_4  g09895(.A(new_n12242), .B(new_n7337), .Y(new_n12244));
  nor_5  g09896(.A(new_n12244), .B(new_n6723), .Y(new_n12245));
  or_6   g09897(.A(new_n12245), .B(new_n12243), .Y(new_n12246));
  xor_4  g09898(.A(new_n12246), .B(new_n6719), .Y(new_n12247));
  xor_4  g09899(.A(new_n12247), .B(new_n7333), .Y(new_n12248));
  or_6   g09900(.A(new_n12248), .B(new_n12234), .Y(new_n12249));
  xor_4  g09901(.A(new_n12248), .B(new_n12234), .Y(new_n12250));
  xor_4  g09902(.A(new_n12244), .B(new_n6723), .Y(new_n12251));
  xor_4  g09903(.A(new_n12216), .B(pi401), .Y(new_n12252));
  nand_5 g09904(.A(new_n12236), .B(new_n12235), .Y(new_n12253));
  nor_5  g09905(.A(pi435), .B(new_n2874), .Y(new_n12254));
  nand_5 g09906(.A(pi435), .B(new_n2874), .Y(new_n12255));
  not_8  g09907(.A(new_n12255), .Y(new_n12256));
  nor_5  g09908(.A(new_n12256), .B(new_n12254), .Y(new_n12257));
  xor_4  g09909(.A(new_n12257), .B(pi390), .Y(new_n12258));
  nand_5 g09910(.A(new_n12258), .B(new_n11356), .Y(new_n12259));
  not_8  g09911(.A(new_n12258), .Y(new_n12260));
  nand_5 g09912(.A(new_n12260), .B(new_n11357), .Y(new_n12261));
  nand_5 g09913(.A(new_n12261), .B(new_n12259), .Y(new_n12262));
  xnor_4 g09914(.A(new_n12262), .B(new_n12253), .Y(new_n12263));
  nand_5 g09915(.A(new_n12263), .B(new_n12252), .Y(new_n12264));
  and_6  g09916(.A(new_n12260), .B(new_n11358), .Y(new_n12265));
  or_6   g09917(.A(new_n12265), .B(new_n12263), .Y(new_n12266));
  nand_5 g09918(.A(new_n12266), .B(new_n12264), .Y(new_n12267));
  xor_4  g09919(.A(new_n12238), .B(new_n6726), .Y(new_n12268));
  xor_4  g09920(.A(new_n12268), .B(new_n7341), .Y(new_n12269));
  nand_5 g09921(.A(new_n12269), .B(new_n12267), .Y(new_n12270));
  nand_5 g09922(.A(new_n12212), .B(new_n12211), .Y(new_n12271));
  xor_4  g09923(.A(new_n12271), .B(new_n12219), .Y(new_n12272));
  not_8  g09924(.A(new_n12272), .Y(new_n12273));
  or_6   g09925(.A(new_n12269), .B(new_n12267), .Y(new_n12274));
  nand_5 g09926(.A(new_n12274), .B(new_n12273), .Y(new_n12275));
  nand_5 g09927(.A(new_n12275), .B(new_n12270), .Y(new_n12276));
  or_6   g09928(.A(new_n12276), .B(new_n12251), .Y(new_n12277));
  xor_4  g09929(.A(new_n12221), .B(new_n12210), .Y(new_n12278));
  xor_4  g09930(.A(new_n12276), .B(new_n12251), .Y(new_n12279));
  nand_5 g09931(.A(new_n12279), .B(new_n12278), .Y(new_n12280));
  nand_5 g09932(.A(new_n12280), .B(new_n12277), .Y(new_n12281));
  nand_5 g09933(.A(new_n12281), .B(new_n12250), .Y(new_n12282));
  nand_5 g09934(.A(new_n12282), .B(new_n12249), .Y(new_n12283));
  nor_5  g09935(.A(new_n12246), .B(pi579), .Y(new_n12284));
  nor_5  g09936(.A(new_n12247), .B(new_n7332), .Y(new_n12285));
  or_6   g09937(.A(new_n12285), .B(new_n12284), .Y(new_n12286));
  nand_5 g09938(.A(new_n12286), .B(new_n7329), .Y(new_n12287));
  or_6   g09939(.A(new_n12286), .B(new_n7329), .Y(new_n12288));
  nand_5 g09940(.A(new_n12288), .B(new_n12287), .Y(new_n12289));
  xor_4  g09941(.A(new_n12289), .B(pi615), .Y(new_n12290));
  nor_5  g09942(.A(new_n12290), .B(new_n12283), .Y(new_n12291));
  xor_4  g09943(.A(new_n12228), .B(new_n12207), .Y(new_n12292));
  not_8  g09944(.A(new_n12292), .Y(new_n12293));
  xnor_4 g09945(.A(new_n12290), .B(new_n12283), .Y(new_n12294));
  nor_5  g09946(.A(new_n12294), .B(new_n12293), .Y(new_n12295));
  or_6   g09947(.A(new_n12295), .B(new_n12291), .Y(new_n12296));
  nand_5 g09948(.A(new_n12287), .B(pi615), .Y(new_n12297));
  nand_5 g09949(.A(new_n12297), .B(new_n12288), .Y(new_n12298));
  or_6   g09950(.A(new_n12298), .B(new_n7324), .Y(new_n12299));
  nand_5 g09951(.A(new_n12298), .B(new_n7324), .Y(new_n12300));
  nand_5 g09952(.A(new_n12300), .B(new_n12299), .Y(new_n12301));
  xor_4  g09953(.A(new_n12301), .B(new_n6714), .Y(new_n12302));
  xor_4  g09954(.A(new_n12302), .B(new_n12296), .Y(new_n12303));
  xor_4  g09955(.A(new_n12303), .B(new_n12232), .Y(po0087));
  nand_5 g09956(.A(new_n3952), .B(pi218), .Y(new_n12305));
  nand_5 g09957(.A(pi350), .B(new_n3976), .Y(new_n12306));
  nand_5 g09958(.A(new_n12306), .B(new_n12305), .Y(new_n12307));
  nand_5 g09959(.A(new_n3979), .B(pi606), .Y(new_n12308));
  nand_5 g09960(.A(new_n6511), .B(new_n12308), .Y(new_n12309));
  nand_5 g09961(.A(pi656), .B(new_n2570), .Y(new_n12310));
  nand_5 g09962(.A(new_n12310), .B(new_n6513), .Y(new_n12311));
  nand_5 g09963(.A(new_n12311), .B(new_n12309), .Y(new_n12312));
  xor_4  g09964(.A(new_n12312), .B(new_n12307), .Y(new_n12313));
  or_6   g09965(.A(new_n12313), .B(new_n6488), .Y(new_n12314));
  nand_5 g09966(.A(new_n12310), .B(new_n12308), .Y(new_n12315));
  nand_5 g09967(.A(new_n12315), .B(new_n6513), .Y(new_n12316));
  nand_5 g09968(.A(new_n12316), .B(new_n12313), .Y(new_n12317));
  nand_5 g09969(.A(new_n12317), .B(new_n12314), .Y(new_n12318));
  xor_4  g09970(.A(pi305), .B(new_n3963), .Y(new_n12319));
  nand_5 g09971(.A(new_n12306), .B(new_n12308), .Y(new_n12320));
  nand_5 g09972(.A(new_n12320), .B(new_n12305), .Y(new_n12321));
  xor_4  g09973(.A(new_n12321), .B(new_n12319), .Y(new_n12322));
  not_8  g09974(.A(new_n12322), .Y(new_n12323));
  nand_5 g09975(.A(new_n12323), .B(new_n12318), .Y(new_n12324));
  xor_4  g09976(.A(new_n12322), .B(new_n12318), .Y(new_n12325));
  or_6   g09977(.A(new_n12325), .B(new_n6522), .Y(new_n12326));
  nand_5 g09978(.A(new_n12326), .B(new_n12324), .Y(new_n12327));
  xor_4  g09979(.A(pi614), .B(new_n3944), .Y(new_n12328));
  nand_5 g09980(.A(pi305), .B(new_n3963), .Y(new_n12329));
  not_8  g09981(.A(new_n12329), .Y(new_n12330));
  not_8  g09982(.A(new_n12319), .Y(new_n12331));
  nor_5  g09983(.A(new_n12321), .B(new_n12331), .Y(new_n12332));
  nor_5  g09984(.A(new_n12332), .B(new_n12330), .Y(new_n12333));
  xor_4  g09985(.A(new_n12333), .B(new_n12328), .Y(new_n12334));
  xor_4  g09986(.A(new_n12334), .B(new_n12327), .Y(new_n12335));
  xor_4  g09987(.A(new_n12335), .B(new_n6510), .Y(po0088));
  xor_4  g09988(.A(new_n7671), .B(new_n7642), .Y(po0089));
  xnor_4 g09989(.A(new_n6362), .B(new_n6339), .Y(po0090));
  not_8  g09990(.A(new_n11134), .Y(new_n12339));
  nand_5 g09991(.A(new_n8980), .B(new_n8966), .Y(new_n12340));
  nand_5 g09992(.A(new_n12340), .B(new_n8982), .Y(new_n12341));
  not_8  g09993(.A(new_n12341), .Y(new_n12342));
  nor_5  g09994(.A(new_n12342), .B(new_n8978), .Y(new_n12343));
  not_8  g09995(.A(new_n8966), .Y(new_n12344));
  not_8  g09996(.A(new_n8982), .Y(new_n12345));
  nand_5 g09997(.A(new_n12345), .B(new_n8977), .Y(new_n12346));
  nor_5  g09998(.A(new_n12346), .B(new_n12344), .Y(new_n12347));
  nor_5  g09999(.A(new_n12347), .B(new_n12343), .Y(new_n12348));
  nand_5 g10000(.A(new_n12348), .B(new_n11090), .Y(new_n12349));
  not_8  g10001(.A(new_n8978), .Y(new_n12350));
  nor_5  g10002(.A(new_n8980), .B(new_n12350), .Y(new_n12351));
  nand_5 g10003(.A(new_n12351), .B(new_n12344), .Y(new_n12352));
  nand_5 g10004(.A(new_n12352), .B(new_n8977), .Y(new_n12353));
  nand_5 g10005(.A(new_n12353), .B(new_n12342), .Y(new_n12354));
  nand_5 g10006(.A(new_n12354), .B(new_n11089), .Y(new_n12355));
  nand_5 g10007(.A(new_n12355), .B(new_n12349), .Y(new_n12356));
  or_6   g10008(.A(new_n12356), .B(new_n12339), .Y(new_n12357));
  nand_5 g10009(.A(new_n11186), .B(new_n8913), .Y(new_n12358));
  or_6   g10010(.A(new_n11199), .B(new_n8928), .Y(new_n12359));
  nand_5 g10011(.A(new_n11196), .B(new_n8928), .Y(new_n12360));
  nand_5 g10012(.A(new_n12360), .B(new_n12359), .Y(new_n12361));
  nor_5  g10013(.A(new_n12361), .B(new_n8841), .Y(new_n12362));
  nor_5  g10014(.A(new_n12359), .B(new_n11204), .Y(new_n12363));
  or_6   g10015(.A(new_n12363), .B(new_n12362), .Y(new_n12364));
  nand_5 g10016(.A(new_n12364), .B(new_n11191), .Y(new_n12365));
  xor_4  g10017(.A(new_n12364), .B(new_n11191), .Y(new_n12366));
  nand_5 g10018(.A(new_n12366), .B(new_n8922), .Y(new_n12367));
  nand_5 g10019(.A(new_n12367), .B(new_n12365), .Y(new_n12368));
  nand_5 g10020(.A(new_n12368), .B(new_n11189), .Y(new_n12369));
  xor_4  g10021(.A(new_n12368), .B(new_n11189), .Y(new_n12370));
  not_8  g10022(.A(new_n12370), .Y(new_n12371));
  or_6   g10023(.A(new_n12371), .B(new_n8917), .Y(new_n12372));
  nand_5 g10024(.A(new_n12372), .B(new_n12369), .Y(new_n12373));
  xnor_4 g10025(.A(new_n11186), .B(new_n8913), .Y(new_n12374));
  or_6   g10026(.A(new_n12374), .B(new_n12373), .Y(new_n12375));
  nand_5 g10027(.A(new_n12375), .B(new_n12358), .Y(new_n12376));
  nand_5 g10028(.A(new_n12376), .B(new_n11181), .Y(new_n12377));
  xnor_4 g10029(.A(new_n12376), .B(new_n11181), .Y(new_n12378));
  or_6   g10030(.A(new_n12378), .B(new_n8911), .Y(new_n12379));
  nand_5 g10031(.A(new_n12379), .B(new_n12377), .Y(new_n12380));
  nand_5 g10032(.A(new_n12380), .B(new_n11174), .Y(new_n12381));
  xor_4  g10033(.A(new_n12380), .B(new_n11175), .Y(new_n12382));
  or_6   g10034(.A(new_n12382), .B(new_n8905), .Y(new_n12383));
  nand_5 g10035(.A(new_n12383), .B(new_n12381), .Y(new_n12384));
  nand_5 g10036(.A(new_n12384), .B(new_n8957), .Y(new_n12385));
  not_8  g10037(.A(new_n11170), .Y(new_n12386));
  xor_4  g10038(.A(new_n12384), .B(new_n8903), .Y(new_n12387));
  or_6   g10039(.A(new_n12387), .B(new_n12386), .Y(new_n12388));
  nand_5 g10040(.A(new_n12388), .B(new_n12385), .Y(new_n12389));
  or_6   g10041(.A(new_n12389), .B(new_n11167), .Y(new_n12390));
  xor_4  g10042(.A(new_n12389), .B(new_n11167), .Y(new_n12391));
  nand_5 g10043(.A(new_n12391), .B(new_n8864), .Y(new_n12392));
  nand_5 g10044(.A(new_n12392), .B(new_n12390), .Y(new_n12393));
  or_6   g10045(.A(new_n12393), .B(new_n11162), .Y(new_n12394));
  nand_5 g10046(.A(new_n12393), .B(new_n11162), .Y(new_n12395));
  nand_5 g10047(.A(new_n12395), .B(new_n8985), .Y(new_n12396));
  nand_5 g10048(.A(new_n12396), .B(new_n12394), .Y(new_n12397));
  nand_5 g10049(.A(new_n12397), .B(new_n12339), .Y(new_n12398));
  xor_4  g10050(.A(new_n12397), .B(new_n12339), .Y(new_n12399));
  nand_5 g10051(.A(new_n12354), .B(new_n11090), .Y(new_n12400));
  nand_5 g10052(.A(new_n12400), .B(new_n12348), .Y(new_n12401));
  not_8  g10053(.A(new_n12401), .Y(new_n12402));
  nand_5 g10054(.A(new_n12402), .B(new_n12356), .Y(new_n12403));
  not_8  g10055(.A(new_n12403), .Y(new_n12404));
  not_8  g10056(.A(new_n12355), .Y(new_n12405));
  nor_5  g10057(.A(new_n12405), .B(new_n12348), .Y(new_n12406));
  nor_5  g10058(.A(new_n12406), .B(new_n12404), .Y(new_n12407));
  nand_5 g10059(.A(new_n12407), .B(new_n12399), .Y(new_n12408));
  nand_5 g10060(.A(new_n12408), .B(new_n12398), .Y(new_n12409));
  xor_4  g10061(.A(new_n12356), .B(new_n12339), .Y(new_n12410));
  nand_5 g10062(.A(new_n12410), .B(new_n12409), .Y(new_n12411));
  nand_5 g10063(.A(new_n12411), .B(new_n12357), .Y(po0091));
  nand_5 g10064(.A(new_n12394), .B(new_n12395), .Y(new_n12413));
  xor_4  g10065(.A(new_n12413), .B(new_n8985), .Y(po0092));
  not_8  g10066(.A(pi517), .Y(new_n12415));
  xor_4  g10067(.A(new_n6243), .B(new_n6237), .Y(new_n12416));
  nand_5 g10068(.A(new_n12416), .B(new_n6427), .Y(new_n12417));
  nand_5 g10069(.A(new_n3949), .B(new_n6437), .Y(new_n12418));
  nand_5 g10070(.A(new_n2570), .B(new_n6472), .Y(new_n12419));
  nand_5 g10071(.A(new_n6440), .B(new_n3952), .Y(new_n12420));
  nor_5  g10072(.A(new_n12420), .B(new_n12419), .Y(new_n12421));
  or_6   g10073(.A(new_n12421), .B(new_n12418), .Y(new_n12422));
  not_8  g10074(.A(new_n12422), .Y(new_n12423));
  xor_4  g10075(.A(pi305), .B(pi188), .Y(new_n12424));
  not_8  g10076(.A(new_n12419), .Y(new_n12425));
  nand_5 g10077(.A(pi487), .B(pi350), .Y(new_n12426));
  nor_5  g10078(.A(new_n12426), .B(new_n12425), .Y(new_n12427));
  or_6   g10079(.A(new_n12427), .B(new_n12421), .Y(new_n12428));
  nor_5  g10080(.A(new_n12428), .B(new_n12424), .Y(new_n12429));
  not_8  g10081(.A(new_n12427), .Y(new_n12430));
  nand_5 g10082(.A(new_n12430), .B(new_n12418), .Y(new_n12431));
  nor_5  g10083(.A(new_n12431), .B(new_n12429), .Y(new_n12432));
  nor_5  g10084(.A(new_n12432), .B(new_n12423), .Y(new_n12433));
  not_8  g10085(.A(new_n12433), .Y(new_n12434));
  nor_5  g10086(.A(new_n12434), .B(new_n6240), .Y(new_n12435));
  not_8  g10087(.A(pi098), .Y(new_n12436));
  nand_5 g10088(.A(new_n12436), .B(new_n3944), .Y(new_n12437));
  not_8  g10089(.A(new_n12437), .Y(new_n12438));
  xor_4  g10090(.A(new_n12438), .B(new_n12435), .Y(new_n12439));
  xor_4  g10091(.A(pi098), .B(new_n3944), .Y(new_n12440));
  or_6   g10092(.A(new_n12440), .B(new_n12433), .Y(new_n12441));
  not_8  g10093(.A(new_n12441), .Y(new_n12442));
  nor_5  g10094(.A(new_n12442), .B(new_n12439), .Y(new_n12443));
  not_8  g10095(.A(pi456), .Y(new_n12444));
  xor_4  g10096(.A(pi479), .B(new_n12444), .Y(new_n12445));
  nor_5  g10097(.A(new_n12445), .B(new_n12443), .Y(new_n12446));
  nand_5 g10098(.A(new_n12438), .B(new_n12435), .Y(new_n12447));
  nand_5 g10099(.A(new_n12447), .B(pi479), .Y(new_n12448));
  nor_5  g10100(.A(new_n12448), .B(new_n12446), .Y(new_n12449));
  xor_4  g10101(.A(new_n12433), .B(new_n6240), .Y(new_n12450));
  nor_5  g10102(.A(new_n12450), .B(new_n12436), .Y(new_n12451));
  or_6   g10103(.A(new_n12451), .B(new_n6243), .Y(new_n12452));
  nand_5 g10104(.A(new_n12452), .B(pi456), .Y(new_n12453));
  nand_5 g10105(.A(new_n12450), .B(new_n12436), .Y(new_n12454));
  nand_5 g10106(.A(pi456), .B(pi058), .Y(new_n12455));
  nor_5  g10107(.A(new_n12455), .B(new_n6239), .Y(new_n12456));
  or_6   g10108(.A(new_n12456), .B(new_n6243), .Y(new_n12457));
  nand_5 g10109(.A(new_n12457), .B(new_n12454), .Y(new_n12458));
  nand_5 g10110(.A(new_n12458), .B(new_n12453), .Y(new_n12459));
  or_6   g10111(.A(new_n12459), .B(new_n12449), .Y(new_n12460));
  nand_5 g10112(.A(new_n12460), .B(new_n12417), .Y(new_n12461));
  or_6   g10113(.A(new_n12416), .B(new_n6427), .Y(new_n12462));
  nand_5 g10114(.A(new_n12462), .B(new_n12461), .Y(new_n12463));
  xor_4  g10115(.A(new_n12463), .B(new_n12415), .Y(new_n12464));
  xor_4  g10116(.A(new_n12464), .B(new_n6248), .Y(new_n12465));
  nor_5  g10117(.A(new_n12465), .B(new_n6234), .Y(new_n12466));
  xor_4  g10118(.A(new_n12465), .B(new_n6280), .Y(new_n12467));
  xor_4  g10119(.A(new_n12440), .B(new_n12433), .Y(new_n12468));
  or_6   g10120(.A(new_n12468), .B(new_n6157), .Y(new_n12469));
  xor_4  g10121(.A(new_n12468), .B(new_n6157), .Y(new_n12470));
  xor_4  g10122(.A(new_n12428), .B(new_n12424), .Y(new_n12471));
  nand_5 g10123(.A(new_n12471), .B(new_n6148), .Y(new_n12472));
  xor_4  g10124(.A(new_n12471), .B(new_n6148), .Y(new_n12473));
  nand_5 g10125(.A(new_n12426), .B(new_n12420), .Y(new_n12474));
  nand_5 g10126(.A(pi606), .B(pi156), .Y(new_n12475));
  nand_5 g10127(.A(new_n12475), .B(new_n12419), .Y(new_n12476));
  or_6   g10128(.A(new_n12476), .B(new_n6135), .Y(new_n12477));
  nand_5 g10129(.A(new_n12477), .B(new_n12475), .Y(new_n12478));
  xor_4  g10130(.A(new_n12478), .B(new_n6134), .Y(new_n12479));
  not_8  g10131(.A(new_n12479), .Y(new_n12480));
  nor_5  g10132(.A(new_n12480), .B(new_n12474), .Y(new_n12481));
  nand_5 g10133(.A(new_n12478), .B(new_n6134), .Y(new_n12482));
  nand_5 g10134(.A(new_n12474), .B(new_n12425), .Y(new_n12483));
  nand_5 g10135(.A(new_n12483), .B(new_n12482), .Y(new_n12484));
  or_6   g10136(.A(new_n12484), .B(new_n12481), .Y(new_n12485));
  nand_5 g10137(.A(new_n12485), .B(new_n12473), .Y(new_n12486));
  nand_5 g10138(.A(new_n12486), .B(new_n12472), .Y(new_n12487));
  nand_5 g10139(.A(new_n12487), .B(new_n12470), .Y(new_n12488));
  nand_5 g10140(.A(new_n12488), .B(new_n12469), .Y(new_n12489));
  nand_5 g10141(.A(new_n12489), .B(new_n6169), .Y(new_n12490));
  xor_4  g10142(.A(new_n12489), .B(new_n6170), .Y(new_n12491));
  xor_4  g10143(.A(new_n12445), .B(new_n12443), .Y(new_n12492));
  or_6   g10144(.A(new_n12492), .B(new_n12491), .Y(new_n12493));
  nand_5 g10145(.A(new_n12493), .B(new_n12490), .Y(new_n12494));
  nand_5 g10146(.A(new_n12462), .B(new_n12417), .Y(new_n12495));
  xor_4  g10147(.A(new_n12495), .B(new_n12460), .Y(new_n12496));
  not_8  g10148(.A(new_n12496), .Y(new_n12497));
  or_6   g10149(.A(new_n12497), .B(new_n12494), .Y(new_n12498));
  xor_4  g10150(.A(new_n12497), .B(new_n12494), .Y(new_n12499));
  nand_5 g10151(.A(new_n12499), .B(new_n6207), .Y(new_n12500));
  nand_5 g10152(.A(new_n12500), .B(new_n12498), .Y(new_n12501));
  nor_5  g10153(.A(new_n12501), .B(new_n12467), .Y(new_n12502));
  or_6   g10154(.A(new_n12502), .B(new_n12466), .Y(new_n12503));
  nand_5 g10155(.A(new_n12503), .B(new_n6311), .Y(new_n12504));
  not_8  g10156(.A(new_n12504), .Y(new_n12505));
  nor_5  g10157(.A(new_n12503), .B(new_n6311), .Y(new_n12506));
  nand_5 g10158(.A(new_n12463), .B(pi517), .Y(new_n12507));
  nor_5  g10159(.A(new_n12507), .B(new_n6274), .Y(new_n12508));
  nor_5  g10160(.A(new_n12463), .B(pi517), .Y(new_n12509));
  nor_5  g10161(.A(new_n12509), .B(new_n6247), .Y(new_n12510));
  nor_5  g10162(.A(new_n12510), .B(new_n12508), .Y(new_n12511));
  xor_4  g10163(.A(pi119), .B(pi054), .Y(new_n12512));
  not_8  g10164(.A(new_n12512), .Y(new_n12513));
  nor_5  g10165(.A(new_n12513), .B(new_n12511), .Y(new_n12514));
  nor_5  g10166(.A(new_n12512), .B(new_n12509), .Y(new_n12515));
  nand_5 g10167(.A(new_n12515), .B(new_n12511), .Y(new_n12516));
  nand_5 g10168(.A(new_n11665), .B(pi119), .Y(new_n12517));
  not_8  g10169(.A(pi119), .Y(new_n12518));
  nand_5 g10170(.A(new_n11664), .B(new_n12518), .Y(new_n12519));
  nand_5 g10171(.A(new_n12519), .B(new_n12517), .Y(new_n12520));
  nand_5 g10172(.A(new_n12520), .B(new_n12509), .Y(new_n12521));
  nand_5 g10173(.A(new_n12521), .B(new_n12516), .Y(new_n12522));
  or_6   g10174(.A(new_n12522), .B(new_n12514), .Y(new_n12523));
  nor_5  g10175(.A(new_n12523), .B(new_n12506), .Y(new_n12524));
  nor_5  g10176(.A(new_n12524), .B(new_n12505), .Y(new_n12525));
  nand_5 g10177(.A(new_n12525), .B(new_n6310), .Y(new_n12526));
  xor_4  g10178(.A(new_n6318), .B(pi070), .Y(new_n12527));
  nand_5 g10179(.A(new_n12523), .B(new_n12519), .Y(new_n12528));
  nand_5 g10180(.A(new_n12528), .B(new_n12517), .Y(new_n12529));
  xor_4  g10181(.A(new_n12529), .B(new_n12527), .Y(new_n12530));
  xor_4  g10182(.A(new_n12525), .B(new_n6310), .Y(new_n12531));
  nand_5 g10183(.A(new_n12531), .B(new_n12530), .Y(new_n12532));
  nand_5 g10184(.A(new_n12532), .B(new_n12526), .Y(new_n12533));
  not_8  g10185(.A(pi327), .Y(new_n12534));
  not_8  g10186(.A(pi070), .Y(new_n12535));
  nand_5 g10187(.A(new_n6318), .B(new_n12535), .Y(new_n12536));
  or_6   g10188(.A(new_n12529), .B(new_n12527), .Y(new_n12537));
  nand_5 g10189(.A(new_n12537), .B(new_n12536), .Y(new_n12538));
  xor_4  g10190(.A(new_n12538), .B(new_n12534), .Y(new_n12539));
  xor_4  g10191(.A(new_n12539), .B(new_n11779), .Y(new_n12540));
  nand_5 g10192(.A(new_n12540), .B(new_n12533), .Y(new_n12541));
  xor_4  g10193(.A(new_n12540), .B(new_n12533), .Y(new_n12542));
  nand_5 g10194(.A(new_n12542), .B(new_n6347), .Y(new_n12543));
  nand_5 g10195(.A(new_n12543), .B(new_n12541), .Y(new_n12544));
  nand_5 g10196(.A(new_n12544), .B(new_n6378), .Y(new_n12545));
  nand_5 g10197(.A(new_n12538), .B(new_n12534), .Y(new_n12546));
  not_8  g10198(.A(new_n12546), .Y(new_n12547));
  nor_5  g10199(.A(new_n12539), .B(new_n6358), .Y(new_n12548));
  nor_5  g10200(.A(new_n12548), .B(new_n11770), .Y(new_n12549));
  nor_5  g10201(.A(new_n12549), .B(new_n12547), .Y(new_n12550));
  not_8  g10202(.A(new_n12550), .Y(new_n12551));
  not_8  g10203(.A(new_n6378), .Y(new_n12552));
  xor_4  g10204(.A(new_n12544), .B(new_n12552), .Y(new_n12553));
  nand_5 g10205(.A(new_n12547), .B(new_n11758), .Y(new_n12554));
  nand_5 g10206(.A(new_n12554), .B(new_n12551), .Y(new_n12555));
  not_8  g10207(.A(new_n12555), .Y(new_n12556));
  nand_5 g10208(.A(new_n12556), .B(new_n12553), .Y(new_n12557));
  nand_5 g10209(.A(new_n12557), .B(new_n12551), .Y(new_n12558));
  nand_5 g10210(.A(new_n12558), .B(new_n12545), .Y(new_n12559));
  not_8  g10211(.A(pi198), .Y(new_n12560));
  nand_5 g10212(.A(new_n12560), .B(pi126), .Y(new_n12561));
  xor_4  g10213(.A(pi198), .B(new_n6294), .Y(new_n12562));
  not_8  g10214(.A(pi112), .Y(new_n12563));
  nand_5 g10215(.A(pi782), .B(new_n12563), .Y(new_n12564));
  nand_5 g10216(.A(new_n6260), .B(pi112), .Y(new_n12565));
  nand_5 g10217(.A(pi150), .B(new_n6554), .Y(new_n12566));
  xor_4  g10218(.A(pi150), .B(new_n6554), .Y(new_n12567));
  nand_5 g10219(.A(pi826), .B(new_n6556), .Y(new_n12568));
  xor_4  g10220(.A(pi826), .B(new_n6556), .Y(new_n12569));
  nand_5 g10221(.A(new_n6429), .B(pi210), .Y(new_n12570));
  xor_4  g10222(.A(pi267), .B(new_n6106), .Y(new_n12571));
  nand_5 g10223(.A(new_n6432), .B(pi129), .Y(new_n12572));
  xor_4  g10224(.A(pi312), .B(new_n6109), .Y(new_n12573));
  nand_5 g10225(.A(new_n6434), .B(pi017), .Y(new_n12574));
  xor_4  g10226(.A(pi471), .B(new_n4112), .Y(new_n12575));
  nand_5 g10227(.A(pi774), .B(new_n6444), .Y(new_n12576));
  nand_5 g10228(.A(pi622), .B(new_n6442), .Y(new_n12577));
  not_8  g10229(.A(new_n12577), .Y(new_n12578));
  xor_4  g10230(.A(pi774), .B(new_n6444), .Y(new_n12579));
  nand_5 g10231(.A(new_n12579), .B(new_n12578), .Y(new_n12580));
  nand_5 g10232(.A(new_n12580), .B(new_n12576), .Y(new_n12581));
  nand_5 g10233(.A(new_n12581), .B(new_n12575), .Y(new_n12582));
  nand_5 g10234(.A(new_n12582), .B(new_n12574), .Y(new_n12583));
  nand_5 g10235(.A(new_n12583), .B(new_n12573), .Y(new_n12584));
  nand_5 g10236(.A(new_n12584), .B(new_n12572), .Y(new_n12585));
  nand_5 g10237(.A(new_n12585), .B(new_n12571), .Y(new_n12586));
  nand_5 g10238(.A(new_n12586), .B(new_n12570), .Y(new_n12587));
  nand_5 g10239(.A(new_n12587), .B(new_n12569), .Y(new_n12588));
  nand_5 g10240(.A(new_n12588), .B(new_n12568), .Y(new_n12589));
  nand_5 g10241(.A(new_n12589), .B(new_n12567), .Y(new_n12590));
  nand_5 g10242(.A(new_n12590), .B(new_n12566), .Y(new_n12591));
  nand_5 g10243(.A(new_n12591), .B(new_n12565), .Y(new_n12592));
  nand_5 g10244(.A(new_n12592), .B(new_n12564), .Y(new_n12593));
  nand_5 g10245(.A(new_n12593), .B(new_n12562), .Y(new_n12594));
  nand_5 g10246(.A(new_n12594), .B(new_n12561), .Y(new_n12595));
  nand_5 g10247(.A(new_n12595), .B(pi197), .Y(new_n12596));
  not_8  g10248(.A(pi170), .Y(new_n12597));
  xor_4  g10249(.A(new_n12595), .B(pi197), .Y(new_n12598));
  nand_5 g10250(.A(new_n12598), .B(new_n12597), .Y(new_n12599));
  nand_5 g10251(.A(new_n12599), .B(new_n12596), .Y(new_n12600));
  xor_4  g10252(.A(new_n12542), .B(new_n6347), .Y(new_n12601));
  not_8  g10253(.A(new_n12601), .Y(new_n12602));
  xor_4  g10254(.A(new_n12501), .B(new_n12467), .Y(new_n12603));
  xnor_4 g10255(.A(new_n12585), .B(new_n12571), .Y(new_n12604));
  xor_4  g10256(.A(new_n12583), .B(new_n12573), .Y(new_n12605));
  xor_4  g10257(.A(new_n12581), .B(new_n12575), .Y(new_n12606));
  not_8  g10258(.A(new_n12606), .Y(new_n12607));
  xor_4  g10259(.A(new_n12476), .B(new_n6135), .Y(new_n12608));
  or_6   g10260(.A(pi622), .B(new_n6442), .Y(new_n12609));
  nor_5  g10261(.A(new_n12609), .B(new_n12608), .Y(new_n12610));
  not_8  g10262(.A(new_n12579), .Y(new_n12611));
  xor_4  g10263(.A(new_n12479), .B(new_n12474), .Y(new_n12612));
  or_6   g10264(.A(new_n12612), .B(new_n12611), .Y(new_n12613));
  nand_5 g10265(.A(new_n12613), .B(new_n12610), .Y(new_n12614));
  nand_5 g10266(.A(new_n12612), .B(new_n12611), .Y(new_n12615));
  nand_5 g10267(.A(new_n12615), .B(new_n12580), .Y(new_n12616));
  nand_5 g10268(.A(new_n12608), .B(new_n12578), .Y(new_n12617));
  not_8  g10269(.A(new_n12580), .Y(new_n12618));
  and_6  g10270(.A(new_n12612), .B(new_n12618), .Y(new_n12619));
  or_6   g10271(.A(new_n12619), .B(new_n12617), .Y(new_n12620));
  nand_5 g10272(.A(new_n12620), .B(new_n12616), .Y(new_n12621));
  nand_5 g10273(.A(new_n12621), .B(new_n12614), .Y(new_n12622));
  nor_5  g10274(.A(new_n12622), .B(new_n12607), .Y(new_n12623));
  xnor_4 g10275(.A(new_n12485), .B(new_n12473), .Y(new_n12624));
  xor_4  g10276(.A(new_n12622), .B(new_n12606), .Y(new_n12625));
  nor_5  g10277(.A(new_n12625), .B(new_n12624), .Y(new_n12626));
  or_6   g10278(.A(new_n12626), .B(new_n12623), .Y(new_n12627));
  or_6   g10279(.A(new_n12627), .B(new_n12605), .Y(new_n12628));
  xor_4  g10280(.A(new_n12627), .B(new_n12605), .Y(new_n12629));
  xnor_4 g10281(.A(new_n12487), .B(new_n12470), .Y(new_n12630));
  nand_5 g10282(.A(new_n12630), .B(new_n12629), .Y(new_n12631));
  nand_5 g10283(.A(new_n12631), .B(new_n12628), .Y(new_n12632));
  nand_5 g10284(.A(new_n12632), .B(new_n12604), .Y(new_n12633));
  xor_4  g10285(.A(new_n12632), .B(new_n12604), .Y(new_n12634));
  xnor_4 g10286(.A(new_n12492), .B(new_n12491), .Y(new_n12635));
  nand_5 g10287(.A(new_n12635), .B(new_n12634), .Y(new_n12636));
  nand_5 g10288(.A(new_n12636), .B(new_n12633), .Y(new_n12637));
  xnor_4 g10289(.A(new_n12587), .B(new_n12569), .Y(new_n12638));
  nor_5  g10290(.A(new_n12638), .B(new_n12637), .Y(new_n12639));
  and_6  g10291(.A(new_n12638), .B(new_n12637), .Y(new_n12640));
  xor_4  g10292(.A(new_n12499), .B(new_n6207), .Y(new_n12641));
  nor_5  g10293(.A(new_n12641), .B(new_n12640), .Y(new_n12642));
  or_6   g10294(.A(new_n12642), .B(new_n12639), .Y(new_n12643));
  or_6   g10295(.A(new_n12643), .B(new_n12603), .Y(new_n12644));
  xor_4  g10296(.A(new_n12589), .B(new_n12567), .Y(new_n12645));
  not_8  g10297(.A(new_n12645), .Y(new_n12646));
  xor_4  g10298(.A(new_n12643), .B(new_n12603), .Y(new_n12647));
  nand_5 g10299(.A(new_n12647), .B(new_n12646), .Y(new_n12648));
  nand_5 g10300(.A(new_n12648), .B(new_n12644), .Y(new_n12649));
  nand_5 g10301(.A(new_n12565), .B(new_n12564), .Y(new_n12650));
  xor_4  g10302(.A(new_n12650), .B(new_n12591), .Y(new_n12651));
  nor_5  g10303(.A(new_n12651), .B(new_n12649), .Y(new_n12652));
  not_8  g10304(.A(new_n12651), .Y(new_n12653));
  xor_4  g10305(.A(new_n12653), .B(new_n12649), .Y(new_n12654));
  nor_5  g10306(.A(new_n12506), .B(new_n12505), .Y(new_n12655));
  xor_4  g10307(.A(new_n12655), .B(new_n12523), .Y(new_n12656));
  nor_5  g10308(.A(new_n12656), .B(new_n12654), .Y(new_n12657));
  or_6   g10309(.A(new_n12657), .B(new_n12652), .Y(new_n12658));
  xor_4  g10310(.A(new_n12593), .B(new_n12562), .Y(new_n12659));
  nand_5 g10311(.A(new_n12659), .B(new_n12658), .Y(new_n12660));
  xnor_4 g10312(.A(new_n12659), .B(new_n12658), .Y(new_n12661));
  xor_4  g10313(.A(new_n12531), .B(new_n12530), .Y(new_n12662));
  or_6   g10314(.A(new_n12662), .B(new_n12661), .Y(new_n12663));
  nand_5 g10315(.A(new_n12663), .B(new_n12660), .Y(new_n12664));
  or_6   g10316(.A(new_n12664), .B(new_n12602), .Y(new_n12665));
  xor_4  g10317(.A(new_n12598), .B(new_n12597), .Y(new_n12666));
  not_8  g10318(.A(new_n12666), .Y(new_n12667));
  xor_4  g10319(.A(new_n12664), .B(new_n12602), .Y(new_n12668));
  nand_5 g10320(.A(new_n12668), .B(new_n12667), .Y(new_n12669));
  nand_5 g10321(.A(new_n12669), .B(new_n12665), .Y(new_n12670));
  nand_5 g10322(.A(new_n12670), .B(new_n12600), .Y(new_n12671));
  xor_4  g10323(.A(new_n12556), .B(new_n12553), .Y(new_n12672));
  not_8  g10324(.A(new_n12672), .Y(new_n12673));
  xor_4  g10325(.A(new_n12670), .B(new_n12600), .Y(new_n12674));
  nand_5 g10326(.A(new_n12674), .B(new_n12673), .Y(new_n12675));
  nand_5 g10327(.A(new_n12675), .B(new_n12671), .Y(new_n12676));
  nor_5  g10328(.A(new_n12676), .B(new_n12559), .Y(po0093));
  xnor_4 g10329(.A(new_n8942), .B(new_n8924), .Y(po0094));
  xor_4  g10330(.A(new_n11410), .B(new_n7113), .Y(new_n12679));
  not_8  g10331(.A(new_n7175), .Y(new_n12680));
  or_6   g10332(.A(new_n11415), .B(new_n12680), .Y(new_n12681));
  xor_4  g10333(.A(new_n11415), .B(new_n12680), .Y(new_n12682));
  nor_5  g10334(.A(new_n11420), .B(new_n7165), .Y(new_n12683));
  xnor_4 g10335(.A(new_n11420), .B(new_n7165), .Y(new_n12684));
  nor_5  g10336(.A(new_n7119), .B(new_n4687), .Y(new_n12685));
  nor_5  g10337(.A(new_n7125), .B(new_n4698), .Y(new_n12686));
  and_6  g10338(.A(new_n7157), .B(new_n4577), .Y(new_n12687));
  xor_4  g10339(.A(new_n7157), .B(new_n4578), .Y(new_n12688));
  nand_5 g10340(.A(new_n7151), .B(new_n4588), .Y(new_n12689));
  or_6   g10341(.A(new_n7151), .B(new_n4588), .Y(new_n12690));
  nand_5 g10342(.A(new_n7132), .B(new_n4542), .Y(new_n12691));
  nand_5 g10343(.A(new_n7134), .B(new_n4609), .Y(new_n12692));
  xor_4  g10344(.A(new_n7132), .B(new_n4542), .Y(new_n12693));
  nand_5 g10345(.A(new_n7135), .B(new_n4545), .Y(new_n12694));
  nand_5 g10346(.A(new_n12694), .B(new_n12692), .Y(new_n12695));
  or_6   g10347(.A(new_n12695), .B(new_n12693), .Y(new_n12696));
  nand_5 g10348(.A(new_n12696), .B(new_n12692), .Y(new_n12697));
  nand_5 g10349(.A(new_n12697), .B(new_n12691), .Y(new_n12698));
  not_8  g10350(.A(new_n4546), .Y(new_n12699));
  nand_5 g10351(.A(new_n7136), .B(new_n12699), .Y(new_n12700));
  nand_5 g10352(.A(new_n12700), .B(new_n12698), .Y(new_n12701));
  nand_5 g10353(.A(new_n12701), .B(new_n12690), .Y(new_n12702));
  nand_5 g10354(.A(new_n12702), .B(new_n12689), .Y(new_n12703));
  nor_5  g10355(.A(new_n12703), .B(new_n12688), .Y(new_n12704));
  nor_5  g10356(.A(new_n12704), .B(new_n12687), .Y(new_n12705));
  xor_4  g10357(.A(new_n7125), .B(new_n4552), .Y(new_n12706));
  nor_5  g10358(.A(new_n12706), .B(new_n12705), .Y(new_n12707));
  nor_5  g10359(.A(new_n12707), .B(new_n12686), .Y(new_n12708));
  xor_4  g10360(.A(new_n7120), .B(new_n4687), .Y(new_n12709));
  nor_5  g10361(.A(new_n12709), .B(new_n12708), .Y(new_n12710));
  nor_5  g10362(.A(new_n12710), .B(new_n12685), .Y(new_n12711));
  nor_5  g10363(.A(new_n12711), .B(new_n12684), .Y(new_n12712));
  or_6   g10364(.A(new_n12712), .B(new_n12683), .Y(new_n12713));
  not_8  g10365(.A(new_n12713), .Y(new_n12714));
  nand_5 g10366(.A(new_n12714), .B(new_n12682), .Y(new_n12715));
  nand_5 g10367(.A(new_n12715), .B(new_n12681), .Y(new_n12716));
  xnor_4 g10368(.A(new_n12716), .B(new_n12679), .Y(po0095));
  xor_4  g10369(.A(pi657), .B(pi493), .Y(new_n12718));
  nor_5  g10370(.A(pi743), .B(pi536), .Y(new_n12719));
  not_8  g10371(.A(pi536), .Y(new_n12720));
  nor_5  g10372(.A(new_n4705), .B(new_n12720), .Y(new_n12721));
  nor_5  g10373(.A(pi450), .B(pi444), .Y(new_n12722));
  xor_4  g10374(.A(pi450), .B(pi444), .Y(new_n12723));
  not_8  g10375(.A(new_n12723), .Y(new_n12724));
  nand_5 g10376(.A(pi094), .B(pi052), .Y(new_n12725));
  nor_5  g10377(.A(pi386), .B(pi020), .Y(new_n12726));
  nand_5 g10378(.A(pi574), .B(pi299), .Y(new_n12727));
  not_8  g10379(.A(new_n12727), .Y(new_n12728));
  not_8  g10380(.A(pi020), .Y(new_n12729));
  xor_4  g10381(.A(pi386), .B(new_n12729), .Y(new_n12730));
  or_6   g10382(.A(new_n12730), .B(new_n12728), .Y(new_n12731));
  not_8  g10383(.A(new_n12731), .Y(new_n12732));
  nor_5  g10384(.A(new_n12732), .B(new_n12726), .Y(new_n12733));
  xor_4  g10385(.A(pi094), .B(new_n4641), .Y(new_n12734));
  not_8  g10386(.A(new_n12734), .Y(new_n12735));
  nand_5 g10387(.A(new_n12735), .B(new_n12733), .Y(new_n12736));
  nand_5 g10388(.A(new_n12736), .B(new_n12725), .Y(new_n12737));
  nor_5  g10389(.A(new_n12737), .B(new_n12724), .Y(new_n12738));
  nor_5  g10390(.A(new_n12738), .B(new_n12722), .Y(new_n12739));
  nor_5  g10391(.A(new_n12739), .B(new_n12721), .Y(new_n12740));
  nor_5  g10392(.A(new_n12740), .B(new_n12719), .Y(new_n12741));
  xnor_4 g10393(.A(new_n12741), .B(new_n12718), .Y(new_n12742));
  nand_5 g10394(.A(new_n4631), .B(pi367), .Y(new_n12743));
  not_8  g10395(.A(new_n12743), .Y(new_n12744));
  nand_5 g10396(.A(new_n12744), .B(pi270), .Y(new_n12745));
  nand_5 g10397(.A(new_n12730), .B(new_n12728), .Y(new_n12746));
  nand_5 g10398(.A(new_n12746), .B(pi270), .Y(new_n12747));
  nand_5 g10399(.A(new_n12747), .B(new_n6975), .Y(new_n12748));
  nand_5 g10400(.A(new_n12730), .B(new_n6972), .Y(new_n12749));
  nor_5  g10401(.A(new_n12749), .B(new_n4631), .Y(new_n12750));
  nor_5  g10402(.A(new_n12750), .B(new_n12732), .Y(new_n12751));
  nand_5 g10403(.A(new_n12751), .B(new_n12748), .Y(new_n12752));
  nand_5 g10404(.A(new_n12752), .B(new_n12745), .Y(new_n12753));
  xor_4  g10405(.A(new_n12734), .B(new_n12733), .Y(new_n12754));
  nor_5  g10406(.A(new_n12754), .B(new_n12753), .Y(new_n12755));
  xor_4  g10407(.A(new_n12754), .B(new_n12753), .Y(new_n12756));
  nand_5 g10408(.A(new_n12756), .B(new_n6969), .Y(new_n12757));
  not_8  g10409(.A(new_n12757), .Y(new_n12758));
  nor_5  g10410(.A(new_n12758), .B(new_n12755), .Y(new_n12759));
  nand_5 g10411(.A(new_n12759), .B(pi454), .Y(new_n12760));
  xor_4  g10412(.A(new_n12737), .B(new_n12724), .Y(new_n12761));
  not_8  g10413(.A(new_n12761), .Y(new_n12762));
  xor_4  g10414(.A(new_n12759), .B(new_n6966), .Y(new_n12763));
  or_6   g10415(.A(new_n12763), .B(new_n12762), .Y(new_n12764));
  nand_5 g10416(.A(new_n12764), .B(new_n12760), .Y(new_n12765));
  or_6   g10417(.A(new_n12721), .B(new_n12719), .Y(new_n12766));
  xor_4  g10418(.A(new_n12766), .B(new_n12739), .Y(new_n12767));
  nand_5 g10419(.A(new_n12767), .B(new_n12765), .Y(new_n12768));
  or_6   g10420(.A(new_n12767), .B(new_n12765), .Y(new_n12769));
  nand_5 g10421(.A(new_n12769), .B(pi145), .Y(new_n12770));
  nand_5 g10422(.A(new_n12770), .B(new_n12768), .Y(new_n12771));
  nand_5 g10423(.A(new_n12771), .B(new_n12742), .Y(new_n12772));
  xor_4  g10424(.A(new_n12771), .B(new_n12742), .Y(new_n12773));
  nand_5 g10425(.A(new_n12773), .B(pi566), .Y(new_n12774));
  nand_5 g10426(.A(new_n12774), .B(new_n12772), .Y(new_n12775));
  not_8  g10427(.A(pi513), .Y(new_n12776));
  not_8  g10428(.A(pi526), .Y(new_n12777));
  nor_5  g10429(.A(new_n12777), .B(new_n12776), .Y(new_n12778));
  nor_5  g10430(.A(pi526), .B(pi513), .Y(new_n12779));
  nor_5  g10431(.A(new_n12779), .B(new_n12778), .Y(new_n12780));
  nand_5 g10432(.A(pi657), .B(pi493), .Y(new_n12781));
  nand_5 g10433(.A(new_n12741), .B(new_n12718), .Y(new_n12782));
  nand_5 g10434(.A(new_n12782), .B(new_n12781), .Y(new_n12783));
  not_8  g10435(.A(new_n12783), .Y(new_n12784));
  xor_4  g10436(.A(new_n12784), .B(new_n12780), .Y(new_n12785));
  nand_5 g10437(.A(new_n12785), .B(new_n12775), .Y(new_n12786));
  xor_4  g10438(.A(new_n12785), .B(new_n12775), .Y(new_n12787));
  nand_5 g10439(.A(new_n12787), .B(pi667), .Y(new_n12788));
  nand_5 g10440(.A(new_n12788), .B(new_n12786), .Y(new_n12789));
  nor_5  g10441(.A(new_n12784), .B(new_n12779), .Y(new_n12790));
  nor_5  g10442(.A(new_n12790), .B(new_n12778), .Y(new_n12791));
  nand_5 g10443(.A(new_n12791), .B(new_n12789), .Y(new_n12792));
  nand_5 g10444(.A(pi624), .B(pi314), .Y(new_n12793));
  not_8  g10445(.A(pi314), .Y(new_n12794));
  not_8  g10446(.A(pi624), .Y(new_n12795));
  nand_5 g10447(.A(new_n12795), .B(new_n12794), .Y(new_n12796));
  nand_5 g10448(.A(new_n12796), .B(new_n12793), .Y(new_n12797));
  or_6   g10449(.A(new_n12797), .B(pi555), .Y(new_n12798));
  nand_5 g10450(.A(new_n12798), .B(new_n12793), .Y(new_n12799));
  nor_5  g10451(.A(new_n12799), .B(new_n12792), .Y(new_n12800));
  nor_5  g10452(.A(new_n12791), .B(new_n12789), .Y(new_n12801));
  or_6   g10453(.A(new_n12796), .B(new_n6953), .Y(new_n12802));
  nor_5  g10454(.A(new_n12802), .B(new_n12801), .Y(new_n12803));
  or_6   g10455(.A(new_n12803), .B(new_n12800), .Y(new_n12804));
  nor_5  g10456(.A(new_n12804), .B(pi775), .Y(new_n12805));
  nand_5 g10457(.A(new_n12801), .B(new_n12799), .Y(new_n12806));
  nor_5  g10458(.A(new_n12793), .B(pi555), .Y(new_n12807));
  nand_5 g10459(.A(new_n12807), .B(new_n12792), .Y(new_n12808));
  nand_5 g10460(.A(new_n12808), .B(new_n12806), .Y(new_n12809));
  nor_5  g10461(.A(new_n12809), .B(new_n12805), .Y(new_n12810));
  not_8  g10462(.A(pi029), .Y(new_n12811));
  not_8  g10463(.A(pi412), .Y(new_n12812));
  nand_5 g10464(.A(new_n12812), .B(new_n12811), .Y(new_n12813));
  xor_4  g10465(.A(pi412), .B(pi029), .Y(new_n12814));
  not_8  g10466(.A(new_n12814), .Y(new_n12815));
  nor_5  g10467(.A(new_n12809), .B(new_n12804), .Y(new_n12816));
  xor_4  g10468(.A(new_n12816), .B(new_n7181), .Y(new_n12817));
  or_6   g10469(.A(new_n12817), .B(new_n12815), .Y(new_n12818));
  nand_5 g10470(.A(new_n12818), .B(new_n12813), .Y(new_n12819));
  xor_4  g10471(.A(new_n12819), .B(new_n12810), .Y(new_n12820));
  xor_4  g10472(.A(pi678), .B(pi345), .Y(new_n12821));
  and_6  g10473(.A(new_n12821), .B(new_n7187), .Y(new_n12822));
  nor_5  g10474(.A(new_n12821), .B(new_n7187), .Y(new_n12823));
  nor_5  g10475(.A(new_n12823), .B(new_n12822), .Y(new_n12824));
  xor_4  g10476(.A(new_n12824), .B(new_n12820), .Y(new_n12825));
  nand_5 g10477(.A(new_n6951), .B(pi408), .Y(new_n12826));
  xor_4  g10478(.A(pi646), .B(new_n7100), .Y(new_n12827));
  nor_5  g10479(.A(pi423), .B(new_n6955), .Y(new_n12828));
  xor_4  g10480(.A(pi423), .B(pi139), .Y(new_n12829));
  nand_5 g10481(.A(new_n3799), .B(pi071), .Y(new_n12830));
  xor_4  g10482(.A(pi683), .B(new_n6997), .Y(new_n12831));
  nand_5 g10483(.A(new_n4709), .B(pi567), .Y(new_n12832));
  not_8  g10484(.A(new_n12832), .Y(new_n12833));
  xor_4  g10485(.A(pi630), .B(new_n3774), .Y(new_n12834));
  not_8  g10486(.A(new_n12834), .Y(new_n12835));
  nand_5 g10487(.A(new_n4667), .B(pi088), .Y(new_n12836));
  not_8  g10488(.A(new_n12836), .Y(new_n12837));
  xor_4  g10489(.A(pi498), .B(new_n2373), .Y(new_n12838));
  not_8  g10490(.A(new_n12838), .Y(new_n12839));
  nand_5 g10491(.A(pi605), .B(new_n4652), .Y(new_n12840));
  not_8  g10492(.A(new_n12840), .Y(new_n12841));
  xor_4  g10493(.A(pi605), .B(pi191), .Y(new_n12842));
  nand_5 g10494(.A(pi546), .B(new_n2357), .Y(new_n12843));
  nand_5 g10495(.A(new_n5083), .B(pi434), .Y(new_n12844));
  nand_5 g10496(.A(pi765), .B(new_n2361), .Y(new_n12845));
  nand_5 g10497(.A(new_n4626), .B(pi190), .Y(new_n12846));
  nand_5 g10498(.A(new_n4621), .B(pi552), .Y(new_n12847));
  nand_5 g10499(.A(new_n12847), .B(new_n12846), .Y(new_n12848));
  nand_5 g10500(.A(new_n12848), .B(new_n12845), .Y(new_n12849));
  nand_5 g10501(.A(new_n12849), .B(new_n12844), .Y(new_n12850));
  nand_5 g10502(.A(new_n12850), .B(new_n12843), .Y(new_n12851));
  nor_5  g10503(.A(new_n12851), .B(new_n12842), .Y(new_n12852));
  nor_5  g10504(.A(new_n12852), .B(new_n12841), .Y(new_n12853));
  nor_5  g10505(.A(new_n12853), .B(new_n12839), .Y(new_n12854));
  nor_5  g10506(.A(new_n12854), .B(new_n12837), .Y(new_n12855));
  nor_5  g10507(.A(new_n12855), .B(new_n12835), .Y(new_n12856));
  nor_5  g10508(.A(new_n12856), .B(new_n12833), .Y(new_n12857));
  nand_5 g10509(.A(new_n12857), .B(new_n12831), .Y(new_n12858));
  nand_5 g10510(.A(new_n12858), .B(new_n12830), .Y(new_n12859));
  nor_5  g10511(.A(new_n12859), .B(new_n12829), .Y(new_n12860));
  nor_5  g10512(.A(new_n12860), .B(new_n12828), .Y(new_n12861));
  nand_5 g10513(.A(new_n12861), .B(new_n12827), .Y(new_n12862));
  nand_5 g10514(.A(new_n12862), .B(new_n12826), .Y(new_n12863));
  nand_5 g10515(.A(new_n7185), .B(pi272), .Y(new_n12864));
  nand_5 g10516(.A(pi833), .B(new_n7193), .Y(new_n12865));
  nand_5 g10517(.A(new_n12865), .B(new_n12864), .Y(new_n12866));
  not_8  g10518(.A(new_n12866), .Y(new_n12867));
  xor_4  g10519(.A(new_n12867), .B(new_n12863), .Y(new_n12868));
  xor_4  g10520(.A(new_n12861), .B(new_n12827), .Y(new_n12869));
  not_8  g10521(.A(new_n12869), .Y(new_n12870));
  xor_4  g10522(.A(new_n12859), .B(new_n12829), .Y(new_n12871));
  xor_4  g10523(.A(new_n12857), .B(new_n12831), .Y(new_n12872));
  not_8  g10524(.A(new_n12872), .Y(new_n12873));
  xor_4  g10525(.A(new_n12853), .B(new_n12838), .Y(new_n12874));
  not_8  g10526(.A(new_n12874), .Y(new_n12875));
  xor_4  g10527(.A(new_n12851), .B(new_n12842), .Y(new_n12876));
  nand_5 g10528(.A(pi682), .B(new_n2419), .Y(new_n12877));
  and_6  g10529(.A(new_n12877), .B(new_n12846), .Y(new_n12878));
  nand_5 g10530(.A(new_n12878), .B(pi259), .Y(new_n12879));
  nand_5 g10531(.A(new_n12879), .B(new_n12846), .Y(new_n12880));
  nand_5 g10532(.A(new_n12847), .B(new_n12845), .Y(new_n12881));
  nor_5  g10533(.A(new_n12881), .B(new_n3728), .Y(new_n12882));
  nor_5  g10534(.A(new_n12882), .B(new_n12880), .Y(new_n12883));
  nand_5 g10535(.A(new_n12881), .B(new_n3728), .Y(new_n12884));
  not_8  g10536(.A(new_n12846), .Y(new_n12885));
  not_8  g10537(.A(new_n12881), .Y(new_n12886));
  nand_5 g10538(.A(new_n12886), .B(new_n12885), .Y(new_n12887));
  nand_5 g10539(.A(new_n12887), .B(new_n12884), .Y(new_n12888));
  nor_5  g10540(.A(new_n12888), .B(new_n12883), .Y(new_n12889));
  nand_5 g10541(.A(new_n12889), .B(pi818), .Y(new_n12890));
  and_6  g10542(.A(new_n12844), .B(new_n12843), .Y(new_n12891));
  xor_4  g10543(.A(new_n12891), .B(new_n12849), .Y(new_n12892));
  xnor_4 g10544(.A(new_n12889), .B(pi818), .Y(new_n12893));
  or_6   g10545(.A(new_n12893), .B(new_n12892), .Y(new_n12894));
  nand_5 g10546(.A(new_n12894), .B(new_n12890), .Y(new_n12895));
  nand_5 g10547(.A(new_n12895), .B(new_n12876), .Y(new_n12896));
  or_6   g10548(.A(new_n12895), .B(new_n12876), .Y(new_n12897));
  nand_5 g10549(.A(new_n12897), .B(pi006), .Y(new_n12898));
  nand_5 g10550(.A(new_n12898), .B(new_n12896), .Y(new_n12899));
  nand_5 g10551(.A(new_n12899), .B(new_n12875), .Y(new_n12900));
  xor_4  g10552(.A(new_n12899), .B(new_n12874), .Y(new_n12901));
  or_6   g10553(.A(new_n12901), .B(new_n3716), .Y(new_n12902));
  nand_5 g10554(.A(new_n12902), .B(new_n12900), .Y(new_n12903));
  nand_5 g10555(.A(new_n12903), .B(pi695), .Y(new_n12904));
  xor_4  g10556(.A(new_n12855), .B(new_n12834), .Y(new_n12905));
  not_8  g10557(.A(new_n12905), .Y(new_n12906));
  xor_4  g10558(.A(new_n12903), .B(pi695), .Y(new_n12907));
  nand_5 g10559(.A(new_n12907), .B(new_n12906), .Y(new_n12908));
  nand_5 g10560(.A(new_n12908), .B(new_n12904), .Y(new_n12909));
  or_6   g10561(.A(new_n12909), .B(new_n12873), .Y(new_n12910));
  nand_5 g10562(.A(new_n12910), .B(pi583), .Y(new_n12911));
  nand_5 g10563(.A(new_n12909), .B(new_n12873), .Y(new_n12912));
  nand_5 g10564(.A(new_n12912), .B(new_n12911), .Y(new_n12913));
  nand_5 g10565(.A(new_n12913), .B(new_n12871), .Y(new_n12914));
  or_6   g10566(.A(new_n12913), .B(new_n12871), .Y(new_n12915));
  nand_5 g10567(.A(new_n12915), .B(pi809), .Y(new_n12916));
  nand_5 g10568(.A(new_n12916), .B(new_n12914), .Y(new_n12917));
  nand_5 g10569(.A(new_n12917), .B(new_n12870), .Y(new_n12918));
  or_6   g10570(.A(new_n12917), .B(new_n12870), .Y(new_n12919));
  nand_5 g10571(.A(new_n12919), .B(pi556), .Y(new_n12920));
  nand_5 g10572(.A(new_n12920), .B(new_n12918), .Y(new_n12921));
  nand_5 g10573(.A(new_n12921), .B(pi323), .Y(new_n12922));
  nor_5  g10574(.A(new_n12921), .B(pi323), .Y(new_n12923));
  not_8  g10575(.A(new_n12923), .Y(new_n12924));
  nand_5 g10576(.A(new_n12924), .B(new_n12922), .Y(new_n12925));
  xor_4  g10577(.A(new_n12925), .B(new_n12868), .Y(new_n12926));
  not_8  g10578(.A(new_n12926), .Y(new_n12927));
  nor_5  g10579(.A(new_n12927), .B(new_n12825), .Y(new_n12928));
  xor_4  g10580(.A(new_n12926), .B(new_n12825), .Y(new_n12929));
  and_6  g10581(.A(new_n12915), .B(new_n12914), .Y(new_n12930));
  xor_4  g10582(.A(new_n12930), .B(new_n11901), .Y(new_n12931));
  xor_4  g10583(.A(new_n12791), .B(new_n12789), .Y(new_n12932));
  xor_4  g10584(.A(new_n12797), .B(pi555), .Y(new_n12933));
  xor_4  g10585(.A(new_n12933), .B(new_n12932), .Y(new_n12934));
  nor_5  g10586(.A(new_n12934), .B(new_n12931), .Y(new_n12935));
  not_8  g10587(.A(new_n12931), .Y(new_n12936));
  xor_4  g10588(.A(new_n12934), .B(new_n12936), .Y(new_n12937));
  and_6  g10589(.A(new_n12912), .B(new_n12910), .Y(new_n12938));
  xor_4  g10590(.A(new_n12938), .B(new_n4724), .Y(new_n12939));
  xor_4  g10591(.A(new_n12787), .B(new_n6957), .Y(new_n12940));
  nor_5  g10592(.A(new_n12940), .B(new_n12939), .Y(new_n12941));
  nand_5 g10593(.A(new_n12940), .B(new_n12939), .Y(new_n12942));
  xor_4  g10594(.A(new_n12773), .B(new_n6960), .Y(new_n12943));
  xor_4  g10595(.A(new_n12907), .B(new_n12905), .Y(new_n12944));
  nor_5  g10596(.A(new_n12944), .B(new_n12943), .Y(new_n12945));
  nand_5 g10597(.A(new_n12768), .B(new_n12769), .Y(new_n12946));
  xor_4  g10598(.A(new_n12946), .B(pi145), .Y(new_n12947));
  xor_4  g10599(.A(new_n12901), .B(pi805), .Y(new_n12948));
  nor_5  g10600(.A(new_n12948), .B(new_n12947), .Y(new_n12949));
  not_8  g10601(.A(new_n12948), .Y(new_n12950));
  xor_4  g10602(.A(new_n12950), .B(new_n12947), .Y(new_n12951));
  xor_4  g10603(.A(new_n12763), .B(new_n12761), .Y(new_n12952));
  and_6  g10604(.A(new_n12897), .B(new_n12896), .Y(new_n12953));
  xor_4  g10605(.A(new_n12953), .B(new_n3720), .Y(new_n12954));
  nor_5  g10606(.A(new_n12954), .B(new_n12952), .Y(new_n12955));
  not_8  g10607(.A(new_n12954), .Y(new_n12956));
  xor_4  g10608(.A(new_n12956), .B(new_n12952), .Y(new_n12957));
  not_8  g10609(.A(new_n12892), .Y(new_n12958));
  xor_4  g10610(.A(new_n12893), .B(new_n12958), .Y(new_n12959));
  xor_4  g10611(.A(new_n12756), .B(pi731), .Y(new_n12960));
  not_8  g10612(.A(new_n12960), .Y(new_n12961));
  nand_5 g10613(.A(new_n12961), .B(new_n12959), .Y(new_n12962));
  or_6   g10614(.A(new_n12961), .B(new_n12959), .Y(new_n12963));
  xor_4  g10615(.A(new_n12878), .B(pi259), .Y(new_n12964));
  nand_5 g10616(.A(new_n12728), .B(new_n6975), .Y(new_n12965));
  nand_5 g10617(.A(new_n12965), .B(new_n12743), .Y(new_n12966));
  not_8  g10618(.A(new_n12966), .Y(new_n12967));
  nand_5 g10619(.A(new_n12967), .B(new_n12964), .Y(new_n12968));
  xor_4  g10620(.A(new_n12964), .B(new_n10978), .Y(new_n12969));
  nand_5 g10621(.A(new_n12969), .B(new_n4631), .Y(new_n12970));
  not_8  g10622(.A(new_n12970), .Y(new_n12971));
  nand_5 g10623(.A(new_n12727), .B(pi367), .Y(new_n12972));
  nor_5  g10624(.A(new_n12972), .B(new_n12964), .Y(new_n12973));
  nor_5  g10625(.A(new_n12973), .B(new_n12971), .Y(new_n12974));
  nand_5 g10626(.A(new_n12974), .B(new_n12968), .Y(new_n12975));
  xor_4  g10627(.A(new_n12881), .B(new_n3728), .Y(new_n12976));
  xor_4  g10628(.A(new_n12976), .B(new_n12880), .Y(new_n12977));
  or_6   g10629(.A(new_n12977), .B(new_n12975), .Y(new_n12978));
  nand_5 g10630(.A(new_n12964), .B(new_n10978), .Y(new_n12979));
  nand_5 g10631(.A(new_n12979), .B(new_n12744), .Y(new_n12980));
  nand_5 g10632(.A(new_n12980), .B(new_n12978), .Y(new_n12981));
  xor_4  g10633(.A(new_n12730), .B(pi270), .Y(new_n12982));
  nand_5 g10634(.A(new_n12982), .B(new_n12981), .Y(new_n12983));
  nand_5 g10635(.A(new_n12977), .B(new_n12975), .Y(new_n12984));
  and_6  g10636(.A(new_n12974), .B(new_n12966), .Y(new_n12985));
  nor_5  g10637(.A(new_n12985), .B(new_n12982), .Y(new_n12986));
  nand_5 g10638(.A(new_n12986), .B(new_n12984), .Y(new_n12987));
  nand_5 g10639(.A(new_n12987), .B(new_n12983), .Y(new_n12988));
  nand_5 g10640(.A(new_n12988), .B(new_n12963), .Y(new_n12989));
  nand_5 g10641(.A(new_n12989), .B(new_n12962), .Y(new_n12990));
  nor_5  g10642(.A(new_n12990), .B(new_n12957), .Y(new_n12991));
  nor_5  g10643(.A(new_n12991), .B(new_n12955), .Y(new_n12992));
  nor_5  g10644(.A(new_n12992), .B(new_n12951), .Y(new_n12993));
  nor_5  g10645(.A(new_n12993), .B(new_n12949), .Y(new_n12994));
  not_8  g10646(.A(new_n12944), .Y(new_n12995));
  xor_4  g10647(.A(new_n12995), .B(new_n12943), .Y(new_n12996));
  nor_5  g10648(.A(new_n12996), .B(new_n12994), .Y(new_n12997));
  or_6   g10649(.A(new_n12997), .B(new_n12945), .Y(new_n12998));
  and_6  g10650(.A(new_n12998), .B(new_n12942), .Y(new_n12999));
  nor_5  g10651(.A(new_n12999), .B(new_n12941), .Y(new_n13000));
  nor_5  g10652(.A(new_n13000), .B(new_n12937), .Y(new_n13001));
  or_6   g10653(.A(new_n13001), .B(new_n12935), .Y(new_n13002));
  and_6  g10654(.A(new_n12919), .B(new_n12918), .Y(new_n13003));
  xor_4  g10655(.A(new_n13003), .B(new_n11934), .Y(new_n13004));
  not_8  g10656(.A(new_n13004), .Y(new_n13005));
  and_6  g10657(.A(new_n13005), .B(new_n13002), .Y(new_n13006));
  xor_4  g10658(.A(new_n13004), .B(new_n13002), .Y(new_n13007));
  xor_4  g10659(.A(new_n12817), .B(new_n12814), .Y(new_n13008));
  nor_5  g10660(.A(new_n13008), .B(new_n13007), .Y(new_n13009));
  nor_5  g10661(.A(new_n13009), .B(new_n13006), .Y(new_n13010));
  nor_5  g10662(.A(new_n13010), .B(new_n12929), .Y(new_n13011));
  or_6   g10663(.A(new_n13011), .B(new_n12928), .Y(new_n13012));
  nand_5 g10664(.A(new_n12867), .B(new_n12863), .Y(new_n13013));
  nand_5 g10665(.A(new_n13013), .B(new_n12864), .Y(new_n13014));
  or_6   g10666(.A(new_n13014), .B(new_n12922), .Y(new_n13015));
  nor_5  g10667(.A(new_n12865), .B(new_n12863), .Y(new_n13016));
  nand_5 g10668(.A(new_n13016), .B(new_n12924), .Y(new_n13017));
  not_8  g10669(.A(new_n13017), .Y(new_n13018));
  not_8  g10670(.A(new_n12863), .Y(new_n13019));
  nor_5  g10671(.A(new_n12864), .B(new_n13019), .Y(new_n13020));
  nand_5 g10672(.A(new_n13020), .B(new_n12922), .Y(new_n13021));
  nand_5 g10673(.A(new_n13014), .B(new_n12923), .Y(new_n13022));
  nand_5 g10674(.A(new_n13022), .B(new_n13021), .Y(new_n13023));
  nor_5  g10675(.A(new_n13023), .B(new_n13018), .Y(new_n13024));
  nand_5 g10676(.A(new_n13024), .B(new_n13015), .Y(new_n13025));
  not_8  g10677(.A(new_n13025), .Y(new_n13026));
  and_6  g10678(.A(new_n12819), .B(new_n12810), .Y(new_n13027));
  nor_5  g10679(.A(new_n12823), .B(new_n13027), .Y(new_n13028));
  or_6   g10680(.A(new_n12819), .B(new_n12810), .Y(new_n13029));
  not_8  g10681(.A(pi345), .Y(new_n13030));
  not_8  g10682(.A(pi678), .Y(new_n13031));
  nor_5  g10683(.A(new_n13031), .B(new_n13030), .Y(new_n13032));
  nor_5  g10684(.A(new_n12822), .B(new_n13032), .Y(new_n13033));
  nand_5 g10685(.A(new_n13033), .B(new_n13029), .Y(new_n13034));
  nor_5  g10686(.A(new_n13034), .B(new_n13028), .Y(new_n13035));
  not_8  g10687(.A(new_n12824), .Y(new_n13036));
  nand_5 g10688(.A(new_n13036), .B(new_n12820), .Y(new_n13037));
  nor_5  g10689(.A(new_n13033), .B(new_n13027), .Y(new_n13038));
  and_6  g10690(.A(new_n13038), .B(new_n13037), .Y(new_n13039));
  or_6   g10691(.A(new_n13039), .B(new_n13035), .Y(new_n13040));
  xor_4  g10692(.A(new_n13040), .B(new_n13026), .Y(new_n13041));
  nand_5 g10693(.A(new_n13041), .B(new_n13012), .Y(new_n13042));
  not_8  g10694(.A(new_n13042), .Y(new_n13043));
  nand_5 g10695(.A(new_n13024), .B(new_n13014), .Y(new_n13044));
  not_8  g10696(.A(new_n13044), .Y(new_n13045));
  xor_4  g10697(.A(new_n13045), .B(new_n13035), .Y(new_n13046));
  nand_5 g10698(.A(new_n13046), .B(new_n13043), .Y(new_n13047));
  nor_5  g10699(.A(new_n13040), .B(new_n13026), .Y(new_n13048));
  nor_5  g10700(.A(new_n13046), .B(new_n13048), .Y(new_n13049));
  nand_5 g10701(.A(new_n13049), .B(new_n13042), .Y(new_n13050));
  nand_5 g10702(.A(new_n13050), .B(new_n13047), .Y(po0096));
  xor_4  g10703(.A(new_n11484), .B(new_n4704), .Y(po0097));
  not_8  g10704(.A(pi292), .Y(new_n13053));
  xor_4  g10705(.A(pi713), .B(new_n13053), .Y(new_n13054));
  xor_4  g10706(.A(pi607), .B(pi341), .Y(new_n13055));
  nand_5 g10707(.A(pi203), .B(pi021), .Y(new_n13056));
  nand_5 g10708(.A(new_n10715), .B(new_n10712), .Y(new_n13057));
  nand_5 g10709(.A(new_n13057), .B(new_n13056), .Y(new_n13058));
  xor_4  g10710(.A(new_n13058), .B(new_n13055), .Y(new_n13059));
  or_6   g10711(.A(new_n10716), .B(new_n10711), .Y(new_n13060));
  not_8  g10712(.A(new_n10720), .Y(new_n13061));
  nand_5 g10713(.A(new_n13061), .B(new_n10717), .Y(new_n13062));
  nand_5 g10714(.A(new_n13062), .B(new_n13060), .Y(new_n13063));
  nor_5  g10715(.A(new_n13063), .B(new_n13059), .Y(new_n13064));
  nand_5 g10716(.A(new_n13063), .B(new_n13059), .Y(new_n13065));
  nand_5 g10717(.A(new_n13065), .B(new_n10966), .Y(new_n13066));
  not_8  g10718(.A(new_n13066), .Y(new_n13067));
  nor_5  g10719(.A(new_n13067), .B(new_n13064), .Y(new_n13068));
  nand_5 g10720(.A(pi607), .B(pi341), .Y(new_n13069));
  nand_5 g10721(.A(new_n13058), .B(new_n13055), .Y(new_n13070));
  nand_5 g10722(.A(new_n13070), .B(new_n13069), .Y(new_n13071));
  nand_5 g10723(.A(new_n13071), .B(pi381), .Y(new_n13072));
  not_8  g10724(.A(new_n13072), .Y(new_n13073));
  nor_5  g10725(.A(new_n13071), .B(pi381), .Y(new_n13074));
  nor_5  g10726(.A(new_n13074), .B(new_n13073), .Y(new_n13075));
  xor_4  g10727(.A(new_n13075), .B(new_n13068), .Y(new_n13076));
  xor_4  g10728(.A(new_n13076), .B(new_n13054), .Y(new_n13077));
  not_8  g10729(.A(new_n6101), .Y(new_n13078));
  xor_4  g10730(.A(new_n13063), .B(new_n13059), .Y(new_n13079));
  xor_4  g10731(.A(new_n13079), .B(new_n10966), .Y(new_n13080));
  not_8  g10732(.A(new_n10721), .Y(new_n13081));
  nand_5 g10733(.A(new_n8508), .B(new_n6021), .Y(new_n13082));
  xor_4  g10734(.A(new_n8509), .B(new_n6020), .Y(new_n13083));
  not_8  g10735(.A(new_n5779), .Y(new_n13084));
  nor_5  g10736(.A(new_n8503), .B(new_n13084), .Y(new_n13085));
  nor_5  g10737(.A(new_n13085), .B(new_n8501), .Y(new_n13086));
  nand_5 g10738(.A(new_n13086), .B(new_n13083), .Y(new_n13087));
  nand_5 g10739(.A(new_n13087), .B(new_n13082), .Y(new_n13088));
  nor_5  g10740(.A(new_n13088), .B(new_n6016), .Y(new_n13089));
  xor_4  g10741(.A(new_n13088), .B(new_n6017), .Y(new_n13090));
  nor_5  g10742(.A(new_n13090), .B(new_n8530), .Y(new_n13091));
  or_6   g10743(.A(new_n13091), .B(new_n13089), .Y(new_n13092));
  nand_5 g10744(.A(new_n13092), .B(new_n8546), .Y(new_n13093));
  xor_4  g10745(.A(new_n13092), .B(new_n8545), .Y(new_n13094));
  or_6   g10746(.A(new_n13094), .B(new_n6014), .Y(new_n13095));
  nand_5 g10747(.A(new_n13095), .B(new_n13093), .Y(new_n13096));
  or_6   g10748(.A(new_n13096), .B(new_n10667), .Y(new_n13097));
  xor_4  g10749(.A(new_n13096), .B(new_n10667), .Y(new_n13098));
  nand_5 g10750(.A(new_n13098), .B(new_n6043), .Y(new_n13099));
  nand_5 g10751(.A(new_n13099), .B(new_n13097), .Y(new_n13100));
  nand_5 g10752(.A(new_n13100), .B(new_n10691), .Y(new_n13101));
  not_8  g10753(.A(new_n6052), .Y(new_n13102));
  not_8  g10754(.A(new_n10691), .Y(new_n13103));
  xor_4  g10755(.A(new_n13100), .B(new_n13103), .Y(new_n13104));
  or_6   g10756(.A(new_n13104), .B(new_n13102), .Y(new_n13105));
  nand_5 g10757(.A(new_n13105), .B(new_n13101), .Y(new_n13106));
  nor_5  g10758(.A(new_n13106), .B(new_n10708), .Y(new_n13107));
  not_8  g10759(.A(new_n6055), .Y(new_n13108));
  not_8  g10760(.A(new_n10708), .Y(new_n13109));
  xor_4  g10761(.A(new_n13106), .B(new_n13109), .Y(new_n13110));
  nor_5  g10762(.A(new_n13110), .B(new_n13108), .Y(new_n13111));
  or_6   g10763(.A(new_n13111), .B(new_n13107), .Y(new_n13112));
  nor_5  g10764(.A(new_n13112), .B(new_n13081), .Y(new_n13113));
  xor_4  g10765(.A(new_n13112), .B(new_n10721), .Y(new_n13114));
  nor_5  g10766(.A(new_n13114), .B(new_n6063), .Y(new_n13115));
  or_6   g10767(.A(new_n13115), .B(new_n13113), .Y(new_n13116));
  nor_5  g10768(.A(new_n13116), .B(new_n13080), .Y(new_n13117));
  not_8  g10769(.A(new_n6081), .Y(new_n13118));
  not_8  g10770(.A(new_n13080), .Y(new_n13119));
  xor_4  g10771(.A(new_n13116), .B(new_n13119), .Y(new_n13120));
  nor_5  g10772(.A(new_n13120), .B(new_n13118), .Y(new_n13121));
  or_6   g10773(.A(new_n13121), .B(new_n13117), .Y(new_n13122));
  xor_4  g10774(.A(new_n13122), .B(new_n13078), .Y(new_n13123));
  xnor_4 g10775(.A(new_n13123), .B(new_n13077), .Y(po0098));
  xor_4  g10776(.A(new_n2784), .B(new_n2783), .Y(po0099));
  xor_4  g10777(.A(new_n10622), .B(new_n10580), .Y(po0100));
  xor_4  g10778(.A(new_n5773), .B(new_n5594), .Y(po0101));
  not_8  g10779(.A(new_n11238), .Y(new_n13128));
  nand_5 g10780(.A(new_n11234), .B(new_n4206), .Y(new_n13129));
  nor_5  g10781(.A(new_n13129), .B(new_n13128), .Y(new_n13130));
  xor_4  g10782(.A(new_n13129), .B(new_n11238), .Y(new_n13131));
  nor_5  g10783(.A(new_n13131), .B(new_n4210), .Y(new_n13132));
  nor_5  g10784(.A(new_n13132), .B(new_n13130), .Y(new_n13133));
  nand_5 g10785(.A(new_n13133), .B(new_n4203), .Y(new_n13134));
  xnor_4 g10786(.A(new_n13133), .B(new_n4203), .Y(new_n13135));
  or_6   g10787(.A(new_n13135), .B(new_n11244), .Y(new_n13136));
  nand_5 g10788(.A(new_n13136), .B(new_n13134), .Y(new_n13137));
  nor_5  g10789(.A(new_n13137), .B(new_n11248), .Y(new_n13138));
  xor_4  g10790(.A(new_n13137), .B(new_n11249), .Y(new_n13139));
  nor_5  g10791(.A(new_n13139), .B(new_n4145), .Y(new_n13140));
  or_6   g10792(.A(new_n13140), .B(new_n13138), .Y(new_n13141));
  xor_4  g10793(.A(new_n13141), .B(new_n11256), .Y(new_n13142));
  xor_4  g10794(.A(new_n13142), .B(new_n4232), .Y(po0102));
  xor_4  g10795(.A(new_n11255), .B(new_n11254), .Y(po0103));
  xor_4  g10796(.A(new_n5723), .B(new_n5722), .Y(po0104));
  nor_5  g10797(.A(new_n6581), .B(pi618), .Y(new_n13146));
  not_8  g10798(.A(new_n6582), .Y(new_n13147));
  nor_5  g10799(.A(new_n6595), .B(new_n13147), .Y(new_n13148));
  nor_5  g10800(.A(new_n13148), .B(new_n13146), .Y(new_n13149));
  not_8  g10801(.A(new_n10745), .Y(new_n13150));
  nor_5  g10802(.A(pi545), .B(pi353), .Y(new_n13151));
  nor_5  g10803(.A(new_n6580), .B(new_n6578), .Y(new_n13152));
  nor_5  g10804(.A(new_n13152), .B(new_n13151), .Y(new_n13153));
  xor_4  g10805(.A(new_n13153), .B(pi635), .Y(new_n13154));
  xor_4  g10806(.A(new_n13154), .B(new_n13150), .Y(new_n13155));
  not_8  g10807(.A(new_n13155), .Y(new_n13156));
  xor_4  g10808(.A(new_n13156), .B(new_n13149), .Y(new_n13157));
  not_8  g10809(.A(new_n6596), .Y(new_n13158));
  nand_5 g10810(.A(new_n6633), .B(new_n13158), .Y(new_n13159));
  or_6   g10811(.A(new_n6647), .B(new_n6634), .Y(new_n13160));
  nand_5 g10812(.A(new_n13160), .B(new_n13159), .Y(new_n13161));
  xnor_4 g10813(.A(new_n13161), .B(new_n13157), .Y(new_n13162));
  nand_5 g10814(.A(new_n6644), .B(pi237), .Y(new_n13163));
  nand_5 g10815(.A(new_n13163), .B(new_n6645), .Y(new_n13164));
  or_6   g10816(.A(new_n13164), .B(new_n10660), .Y(new_n13165));
  nand_5 g10817(.A(new_n13164), .B(new_n10660), .Y(new_n13166));
  and_6  g10818(.A(new_n13166), .B(new_n13165), .Y(new_n13167));
  xor_4  g10819(.A(new_n13167), .B(new_n4760), .Y(new_n13168));
  not_8  g10820(.A(new_n13168), .Y(new_n13169));
  xor_4  g10821(.A(new_n13169), .B(new_n13162), .Y(po0105));
  not_8  g10822(.A(new_n3642), .Y(new_n13171));
  xor_4  g10823(.A(new_n13171), .B(new_n3639), .Y(po0106));
  xor_4  g10824(.A(new_n4494), .B(new_n4493), .Y(po0107));
  not_8  g10825(.A(new_n4818), .Y(new_n13174));
  xor_4  g10826(.A(pi634), .B(pi012), .Y(new_n13175));
  nand_5 g10827(.A(new_n4900), .B(new_n3811), .Y(new_n13176));
  nor_5  g10828(.A(new_n8554), .B(new_n3828), .Y(new_n13177));
  not_8  g10829(.A(new_n5829), .Y(new_n13178));
  nor_5  g10830(.A(new_n5831), .B(new_n13178), .Y(new_n13179));
  nor_5  g10831(.A(new_n13179), .B(new_n13177), .Y(new_n13180));
  xor_4  g10832(.A(pi232), .B(pi027), .Y(new_n13181));
  nand_5 g10833(.A(new_n13181), .B(new_n13180), .Y(new_n13182));
  nand_5 g10834(.A(new_n13182), .B(new_n13176), .Y(new_n13183));
  xor_4  g10835(.A(new_n13183), .B(new_n13175), .Y(new_n13184));
  xor_4  g10836(.A(new_n13184), .B(new_n13174), .Y(new_n13185));
  xnor_4 g10837(.A(new_n13181), .B(new_n13180), .Y(new_n13186));
  or_6   g10838(.A(new_n13186), .B(new_n4812), .Y(new_n13187));
  xor_4  g10839(.A(new_n13186), .B(new_n4812), .Y(new_n13188));
  nand_5 g10840(.A(new_n5834), .B(new_n5828), .Y(new_n13189));
  nand_5 g10841(.A(new_n13189), .B(new_n5833), .Y(new_n13190));
  nand_5 g10842(.A(new_n13190), .B(new_n13188), .Y(new_n13191));
  nand_5 g10843(.A(new_n13191), .B(new_n13187), .Y(new_n13192));
  xor_4  g10844(.A(new_n13192), .B(new_n13185), .Y(new_n13193));
  nand_5 g10845(.A(new_n5821), .B(new_n3753), .Y(new_n13194));
  or_6   g10846(.A(new_n5836), .B(new_n5822), .Y(new_n13195));
  nand_5 g10847(.A(new_n13195), .B(new_n13194), .Y(new_n13196));
  not_8  g10848(.A(new_n13196), .Y(new_n13197));
  xnor_4 g10849(.A(new_n13190), .B(new_n13188), .Y(new_n13198));
  nand_5 g10850(.A(new_n13198), .B(new_n13197), .Y(new_n13199));
  xor_4  g10851(.A(new_n13198), .B(new_n13197), .Y(new_n13200));
  nand_5 g10852(.A(new_n13200), .B(new_n3756), .Y(new_n13201));
  nand_5 g10853(.A(new_n13201), .B(new_n13199), .Y(new_n13202));
  xor_4  g10854(.A(new_n13202), .B(new_n13193), .Y(new_n13203));
  xor_4  g10855(.A(new_n13203), .B(new_n3744), .Y(po0108));
  not_8  g10856(.A(new_n5393), .Y(new_n13205));
  nor_5  g10857(.A(new_n13205), .B(new_n5233), .Y(new_n13206));
  nor_5  g10858(.A(new_n5449), .B(new_n5394), .Y(new_n13207));
  or_6   g10859(.A(new_n13207), .B(new_n13206), .Y(new_n13208));
  nand_5 g10860(.A(new_n3209), .B(pi160), .Y(new_n13209));
  nand_5 g10861(.A(pi244), .B(new_n3146), .Y(new_n13210));
  nand_5 g10862(.A(new_n13210), .B(new_n13209), .Y(new_n13211));
  nand_5 g10863(.A(new_n3147), .B(pi005), .Y(new_n13212));
  nand_5 g10864(.A(new_n5232), .B(new_n5203), .Y(new_n13213));
  nand_5 g10865(.A(new_n13213), .B(new_n13212), .Y(new_n13214));
  xnor_4 g10866(.A(new_n13214), .B(new_n13211), .Y(new_n13215));
  xor_4  g10867(.A(new_n13215), .B(new_n13208), .Y(new_n13216));
  not_8  g10868(.A(new_n13216), .Y(new_n13217));
  nand_5 g10869(.A(pi234), .B(pi068), .Y(new_n13218));
  or_6   g10870(.A(pi234), .B(pi068), .Y(new_n13219));
  nand_5 g10871(.A(new_n13219), .B(new_n13218), .Y(new_n13220));
  not_8  g10872(.A(pi189), .Y(new_n13221));
  nand_5 g10873(.A(new_n11899), .B(new_n13221), .Y(new_n13222));
  nand_5 g10874(.A(new_n5311), .B(new_n5271), .Y(new_n13223));
  nand_5 g10875(.A(new_n13223), .B(new_n13222), .Y(new_n13224));
  not_8  g10876(.A(new_n13224), .Y(new_n13225));
  xor_4  g10877(.A(new_n13225), .B(new_n13220), .Y(new_n13226));
  nand_5 g10878(.A(pi687), .B(pi325), .Y(new_n13227));
  nand_5 g10879(.A(new_n5268), .B(new_n5234), .Y(new_n13228));
  nand_5 g10880(.A(new_n13228), .B(new_n13227), .Y(new_n13229));
  nor_5  g10881(.A(new_n13229), .B(pi114), .Y(new_n13230));
  nand_5 g10882(.A(new_n13229), .B(pi114), .Y(new_n13231));
  not_8  g10883(.A(new_n13231), .Y(new_n13232));
  nor_5  g10884(.A(new_n13232), .B(new_n13230), .Y(new_n13233));
  xor_4  g10885(.A(new_n13233), .B(new_n10400), .Y(new_n13234));
  xor_4  g10886(.A(new_n13234), .B(new_n13226), .Y(new_n13235));
  nand_5 g10887(.A(new_n5392), .B(new_n5313), .Y(new_n13236));
  nand_5 g10888(.A(new_n13236), .B(new_n5314), .Y(new_n13237));
  xor_4  g10889(.A(new_n13237), .B(new_n13235), .Y(new_n13238));
  xor_4  g10890(.A(new_n13238), .B(new_n13217), .Y(po0109));
  xnor_4 g10891(.A(new_n11619), .B(new_n11618), .Y(po0110));
  not_8  g10892(.A(new_n5063), .Y(new_n13241));
  xor_4  g10893(.A(new_n13241), .B(new_n3269), .Y(po0111));
  not_8  g10894(.A(new_n12977), .Y(new_n13243));
  nand_5 g10895(.A(new_n12964), .B(new_n10979), .Y(new_n13244));
  nand_5 g10896(.A(new_n13244), .B(pi455), .Y(new_n13245));
  or_6   g10897(.A(new_n12964), .B(new_n10979), .Y(new_n13246));
  nand_5 g10898(.A(new_n13246), .B(new_n13245), .Y(new_n13247));
  nor_5  g10899(.A(new_n13247), .B(new_n13243), .Y(new_n13248));
  xor_4  g10900(.A(new_n13247), .B(new_n12977), .Y(new_n13249));
  nand_5 g10901(.A(pi631), .B(new_n10978), .Y(new_n13250));
  not_8  g10902(.A(new_n13250), .Y(new_n13251));
  xor_4  g10903(.A(pi488), .B(new_n12729), .Y(new_n13252));
  xor_4  g10904(.A(new_n13252), .B(new_n13251), .Y(new_n13253));
  xor_4  g10905(.A(new_n13253), .B(new_n5852), .Y(new_n13254));
  nor_5  g10906(.A(new_n13254), .B(new_n13249), .Y(new_n13255));
  or_6   g10907(.A(new_n13255), .B(new_n13248), .Y(new_n13256));
  not_8  g10908(.A(pi094), .Y(new_n13257));
  xor_4  g10909(.A(pi241), .B(new_n13257), .Y(new_n13258));
  nand_5 g10910(.A(pi488), .B(new_n12729), .Y(new_n13259));
  nand_5 g10911(.A(new_n13252), .B(new_n13251), .Y(new_n13260));
  nand_5 g10912(.A(new_n13260), .B(new_n13259), .Y(new_n13261));
  xor_4  g10913(.A(new_n13261), .B(new_n13258), .Y(new_n13262));
  or_6   g10914(.A(new_n13253), .B(new_n5852), .Y(new_n13263));
  xor_4  g10915(.A(new_n13263), .B(pi261), .Y(new_n13264));
  xor_4  g10916(.A(new_n13264), .B(new_n13262), .Y(new_n13265));
  nand_5 g10917(.A(new_n13265), .B(new_n12959), .Y(new_n13266));
  nand_5 g10918(.A(new_n13266), .B(new_n13256), .Y(new_n13267));
  or_6   g10919(.A(new_n13265), .B(new_n12959), .Y(new_n13268));
  nand_5 g10920(.A(new_n13268), .B(new_n13267), .Y(new_n13269));
  nor_5  g10921(.A(new_n13263), .B(new_n5848), .Y(new_n13270));
  nor_5  g10922(.A(new_n13264), .B(new_n13262), .Y(new_n13271));
  or_6   g10923(.A(new_n13271), .B(new_n13270), .Y(new_n13272));
  xor_4  g10924(.A(pi450), .B(new_n3758), .Y(new_n13273));
  nand_5 g10925(.A(pi241), .B(new_n13257), .Y(new_n13274));
  nand_5 g10926(.A(new_n13261), .B(new_n13258), .Y(new_n13275));
  nand_5 g10927(.A(new_n13275), .B(new_n13274), .Y(new_n13276));
  xnor_4 g10928(.A(new_n13276), .B(new_n13273), .Y(new_n13277));
  xor_4  g10929(.A(new_n13277), .B(new_n5845), .Y(new_n13278));
  xor_4  g10930(.A(new_n13278), .B(new_n13272), .Y(new_n13279));
  xnor_4 g10931(.A(new_n13279), .B(new_n13269), .Y(new_n13280));
  xor_4  g10932(.A(new_n13280), .B(new_n12956), .Y(po0112));
  xnor_4 g10933(.A(new_n10951), .B(new_n10950), .Y(po0113));
  or_6   g10934(.A(new_n7197), .B(new_n3202), .Y(new_n13283));
  nand_5 g10935(.A(new_n7197), .B(new_n3202), .Y(new_n13284));
  or_6   g10936(.A(new_n5184), .B(new_n3162), .Y(new_n13285));
  not_8  g10937(.A(new_n13285), .Y(new_n13286));
  not_8  g10938(.A(new_n5185), .Y(new_n13287));
  nor_5  g10939(.A(new_n5189), .B(new_n13287), .Y(new_n13288));
  nor_5  g10940(.A(new_n13288), .B(new_n13286), .Y(new_n13289));
  nor_5  g10941(.A(new_n13289), .B(new_n7039), .Y(new_n13290));
  xnor_4 g10942(.A(new_n13289), .B(new_n7039), .Y(new_n13291));
  nor_5  g10943(.A(new_n13291), .B(new_n3158), .Y(new_n13292));
  or_6   g10944(.A(new_n13292), .B(new_n13290), .Y(new_n13293));
  nor_5  g10945(.A(new_n13293), .B(new_n3153), .Y(new_n13294));
  xor_4  g10946(.A(new_n13293), .B(new_n3152), .Y(new_n13295));
  nor_5  g10947(.A(new_n13295), .B(new_n7001), .Y(new_n13296));
  nor_5  g10948(.A(new_n13296), .B(new_n13294), .Y(new_n13297));
  nand_5 g10949(.A(new_n13297), .B(new_n7103), .Y(new_n13298));
  xor_4  g10950(.A(new_n13297), .B(new_n7104), .Y(new_n13299));
  or_6   g10951(.A(new_n13299), .B(new_n3148), .Y(new_n13300));
  nand_5 g10952(.A(new_n13300), .B(new_n13298), .Y(new_n13301));
  nand_5 g10953(.A(new_n13301), .B(new_n13284), .Y(new_n13302));
  nand_5 g10954(.A(new_n13302), .B(new_n13283), .Y(new_n13303));
  nand_5 g10955(.A(new_n13303), .B(new_n3145), .Y(new_n13304));
  not_8  g10956(.A(new_n13304), .Y(new_n13305));
  not_8  g10957(.A(new_n7222), .Y(new_n13306));
  nor_5  g10958(.A(new_n13303), .B(new_n3145), .Y(new_n13307));
  or_6   g10959(.A(new_n13307), .B(new_n13305), .Y(new_n13308));
  nor_5  g10960(.A(new_n13308), .B(new_n13306), .Y(new_n13309));
  nor_5  g10961(.A(new_n13309), .B(new_n13305), .Y(new_n13310));
  nand_5 g10962(.A(pi833), .B(new_n3327), .Y(new_n13311));
  xor_4  g10963(.A(pi833), .B(new_n3327), .Y(new_n13312));
  nand_5 g10964(.A(pi646), .B(new_n3262), .Y(new_n13313));
  xor_4  g10965(.A(pi646), .B(new_n3262), .Y(new_n13314));
  nand_5 g10966(.A(new_n3303), .B(pi139), .Y(new_n13315));
  xor_4  g10967(.A(pi637), .B(new_n6955), .Y(new_n13316));
  nand_5 g10968(.A(pi683), .B(new_n3333), .Y(new_n13317));
  xor_4  g10969(.A(pi683), .B(new_n3333), .Y(new_n13318));
  nand_5 g10970(.A(new_n3264), .B(pi567), .Y(new_n13319));
  xor_4  g10971(.A(pi829), .B(new_n3774), .Y(new_n13320));
  nand_5 g10972(.A(new_n5259), .B(pi088), .Y(new_n13321));
  nand_5 g10973(.A(new_n8475), .B(new_n8461), .Y(new_n13322));
  nand_5 g10974(.A(new_n13322), .B(new_n13321), .Y(new_n13323));
  nand_5 g10975(.A(new_n13323), .B(new_n13320), .Y(new_n13324));
  nand_5 g10976(.A(new_n13324), .B(new_n13319), .Y(new_n13325));
  nand_5 g10977(.A(new_n13325), .B(new_n13318), .Y(new_n13326));
  nand_5 g10978(.A(new_n13326), .B(new_n13317), .Y(new_n13327));
  nand_5 g10979(.A(new_n13327), .B(new_n13316), .Y(new_n13328));
  nand_5 g10980(.A(new_n13328), .B(new_n13315), .Y(new_n13329));
  nand_5 g10981(.A(new_n13329), .B(new_n13314), .Y(new_n13330));
  nand_5 g10982(.A(new_n13330), .B(new_n13313), .Y(new_n13331));
  nand_5 g10983(.A(new_n13331), .B(new_n13312), .Y(new_n13332));
  nand_5 g10984(.A(new_n13332), .B(new_n13311), .Y(new_n13333));
  xnor_4 g10985(.A(new_n13331), .B(new_n13312), .Y(new_n13334));
  nand_5 g10986(.A(new_n13284), .B(new_n13283), .Y(new_n13335));
  xor_4  g10987(.A(new_n13335), .B(new_n13301), .Y(new_n13336));
  or_6   g10988(.A(new_n13336), .B(new_n13334), .Y(new_n13337));
  xor_4  g10989(.A(new_n13329), .B(new_n13314), .Y(new_n13338));
  not_8  g10990(.A(new_n13338), .Y(new_n13339));
  xnor_4 g10991(.A(new_n13299), .B(new_n3148), .Y(new_n13340));
  nor_5  g10992(.A(new_n13340), .B(new_n13339), .Y(new_n13341));
  xor_4  g10993(.A(new_n13340), .B(new_n13338), .Y(new_n13342));
  xnor_4 g10994(.A(new_n13295), .B(new_n7001), .Y(new_n13343));
  xor_4  g10995(.A(new_n13327), .B(new_n13316), .Y(new_n13344));
  and_6  g10996(.A(new_n13344), .B(new_n13343), .Y(new_n13345));
  xor_4  g10997(.A(new_n13323), .B(new_n13320), .Y(new_n13346));
  or_6   g10998(.A(new_n13346), .B(new_n5191), .Y(new_n13347));
  xor_4  g10999(.A(new_n13346), .B(new_n5191), .Y(new_n13348));
  nand_5 g11000(.A(new_n8476), .B(new_n5126), .Y(new_n13349));
  or_6   g11001(.A(new_n8499), .B(new_n8477), .Y(new_n13350));
  nand_5 g11002(.A(new_n13350), .B(new_n13349), .Y(new_n13351));
  not_8  g11003(.A(new_n13351), .Y(new_n13352));
  nand_5 g11004(.A(new_n13352), .B(new_n13348), .Y(new_n13353));
  nand_5 g11005(.A(new_n13353), .B(new_n13347), .Y(new_n13354));
  xor_4  g11006(.A(new_n13325), .B(new_n13318), .Y(new_n13355));
  xor_4  g11007(.A(new_n13291), .B(new_n3158), .Y(new_n13356));
  nand_5 g11008(.A(new_n13356), .B(new_n13355), .Y(new_n13357));
  nand_5 g11009(.A(new_n13357), .B(new_n13354), .Y(new_n13358));
  or_6   g11010(.A(new_n13356), .B(new_n13355), .Y(new_n13359));
  nand_5 g11011(.A(new_n13359), .B(new_n13358), .Y(new_n13360));
  xnor_4 g11012(.A(new_n13344), .B(new_n13343), .Y(new_n13361));
  nor_5  g11013(.A(new_n13361), .B(new_n13360), .Y(new_n13362));
  nor_5  g11014(.A(new_n13362), .B(new_n13345), .Y(new_n13363));
  nor_5  g11015(.A(new_n13363), .B(new_n13342), .Y(new_n13364));
  or_6   g11016(.A(new_n13364), .B(new_n13341), .Y(new_n13365));
  xor_4  g11017(.A(new_n13336), .B(new_n13334), .Y(new_n13366));
  nand_5 g11018(.A(new_n13366), .B(new_n13365), .Y(new_n13367));
  nand_5 g11019(.A(new_n13367), .B(new_n13337), .Y(new_n13368));
  xor_4  g11020(.A(new_n13308), .B(new_n7222), .Y(new_n13369));
  not_8  g11021(.A(new_n13369), .Y(new_n13370));
  nor_5  g11022(.A(new_n13370), .B(new_n13368), .Y(new_n13371));
  or_6   g11023(.A(new_n13371), .B(new_n13333), .Y(new_n13372));
  nand_5 g11024(.A(new_n13370), .B(new_n13368), .Y(new_n13373));
  nand_5 g11025(.A(new_n13373), .B(new_n13333), .Y(new_n13374));
  nand_5 g11026(.A(new_n13374), .B(new_n13372), .Y(new_n13375));
  xor_4  g11027(.A(new_n13375), .B(new_n13310), .Y(po0114));
  not_8  g11028(.A(pi531), .Y(new_n13377));
  nand_5 g11029(.A(pi634), .B(new_n13377), .Y(new_n13378));
  xor_4  g11030(.A(pi634), .B(new_n13377), .Y(new_n13379));
  nor_5  g11031(.A(pi464), .B(new_n4900), .Y(new_n13380));
  nor_5  g11032(.A(new_n8554), .B(pi330), .Y(new_n13381));
  xor_4  g11033(.A(pi796), .B(pi330), .Y(new_n13382));
  nand_5 g11034(.A(pi619), .B(new_n4983), .Y(new_n13383));
  nand_5 g11035(.A(new_n13383), .B(new_n9854), .Y(new_n13384));
  nand_5 g11036(.A(new_n4884), .B(pi523), .Y(new_n13385));
  nand_5 g11037(.A(new_n13385), .B(new_n13384), .Y(new_n13386));
  nor_5  g11038(.A(new_n13386), .B(new_n13382), .Y(new_n13387));
  nor_5  g11039(.A(new_n13387), .B(new_n13381), .Y(new_n13388));
  xor_4  g11040(.A(pi464), .B(pi232), .Y(new_n13389));
  nor_5  g11041(.A(new_n13389), .B(new_n13388), .Y(new_n13390));
  or_6   g11042(.A(new_n13390), .B(new_n13380), .Y(new_n13391));
  nand_5 g11043(.A(new_n13391), .B(new_n13379), .Y(new_n13392));
  nand_5 g11044(.A(new_n13392), .B(new_n13378), .Y(new_n13393));
  xor_4  g11045(.A(pi676), .B(pi655), .Y(new_n13394));
  xor_4  g11046(.A(new_n13394), .B(new_n13393), .Y(new_n13395));
  not_8  g11047(.A(new_n13395), .Y(new_n13396));
  xor_4  g11048(.A(new_n13396), .B(new_n7859), .Y(new_n13397));
  xnor_4 g11049(.A(new_n13391), .B(new_n13379), .Y(new_n13398));
  nor_5  g11050(.A(new_n13398), .B(new_n7809), .Y(new_n13399));
  xor_4  g11051(.A(new_n13389), .B(new_n13388), .Y(new_n13400));
  or_6   g11052(.A(new_n13400), .B(new_n7851), .Y(new_n13401));
  xor_4  g11053(.A(new_n13400), .B(new_n7851), .Y(new_n13402));
  not_8  g11054(.A(new_n13402), .Y(new_n13403));
  xor_4  g11055(.A(new_n13386), .B(new_n13382), .Y(new_n13404));
  nand_5 g11056(.A(new_n13404), .B(new_n7816), .Y(new_n13405));
  nand_5 g11057(.A(new_n9857), .B(new_n7819), .Y(new_n13406));
  xor_4  g11058(.A(new_n9855), .B(new_n7830), .Y(new_n13407));
  nand_5 g11059(.A(new_n13407), .B(new_n13406), .Y(new_n13408));
  xor_4  g11060(.A(new_n13408), .B(new_n7826), .Y(new_n13409));
  and_6  g11061(.A(new_n13385), .B(new_n13383), .Y(new_n13410));
  xor_4  g11062(.A(new_n13410), .B(new_n13409), .Y(new_n13411));
  not_8  g11063(.A(new_n13411), .Y(new_n13412));
  nand_5 g11064(.A(new_n9856), .B(new_n7838), .Y(new_n13413));
  nor_5  g11065(.A(new_n13413), .B(new_n7832), .Y(new_n13414));
  nor_5  g11066(.A(new_n13414), .B(new_n13412), .Y(new_n13415));
  nand_5 g11067(.A(new_n13409), .B(new_n9857), .Y(new_n13416));
  nand_5 g11068(.A(new_n13416), .B(new_n7840), .Y(new_n13417));
  or_6   g11069(.A(new_n13417), .B(new_n13415), .Y(new_n13418));
  xor_4  g11070(.A(new_n13404), .B(new_n7815), .Y(new_n13419));
  not_8  g11071(.A(new_n13419), .Y(new_n13420));
  nand_5 g11072(.A(new_n13420), .B(new_n13418), .Y(new_n13421));
  nand_5 g11073(.A(new_n13421), .B(new_n13405), .Y(new_n13422));
  or_6   g11074(.A(new_n13422), .B(new_n13403), .Y(new_n13423));
  nand_5 g11075(.A(new_n13423), .B(new_n13401), .Y(new_n13424));
  xor_4  g11076(.A(new_n13398), .B(new_n7808), .Y(new_n13425));
  or_6   g11077(.A(new_n13425), .B(new_n13424), .Y(new_n13426));
  not_8  g11078(.A(new_n13426), .Y(new_n13427));
  nor_5  g11079(.A(new_n13427), .B(new_n13399), .Y(new_n13428));
  xor_4  g11080(.A(new_n13428), .B(new_n13397), .Y(new_n13429));
  not_8  g11081(.A(new_n13429), .Y(new_n13430));
  not_8  g11082(.A(new_n13425), .Y(new_n13431));
  xor_4  g11083(.A(new_n13431), .B(new_n13424), .Y(new_n13432));
  xor_4  g11084(.A(pi747), .B(new_n8591), .Y(new_n13433));
  nand_5 g11085(.A(pi228), .B(new_n7013), .Y(new_n13434));
  xor_4  g11086(.A(pi228), .B(new_n7013), .Y(new_n13435));
  nand_5 g11087(.A(new_n7016), .B(pi276), .Y(new_n13436));
  nand_5 g11088(.A(pi617), .B(new_n7019), .Y(new_n13437));
  not_8  g11089(.A(new_n9859), .Y(new_n13438));
  xor_4  g11090(.A(pi617), .B(new_n7019), .Y(new_n13439));
  nand_5 g11091(.A(new_n13439), .B(new_n13438), .Y(new_n13440));
  nand_5 g11092(.A(new_n13440), .B(new_n13437), .Y(new_n13441));
  xor_4  g11093(.A(pi294), .B(pi276), .Y(new_n13442));
  not_8  g11094(.A(new_n13442), .Y(new_n13443));
  nand_5 g11095(.A(new_n13443), .B(new_n13441), .Y(new_n13444));
  nand_5 g11096(.A(new_n13444), .B(new_n13436), .Y(new_n13445));
  nand_5 g11097(.A(new_n13445), .B(new_n13435), .Y(new_n13446));
  nand_5 g11098(.A(new_n13446), .B(new_n13434), .Y(new_n13447));
  xnor_4 g11099(.A(new_n13447), .B(new_n13433), .Y(new_n13448));
  nor_5  g11100(.A(new_n13448), .B(new_n13432), .Y(new_n13449));
  xor_4  g11101(.A(new_n13422), .B(new_n13402), .Y(new_n13450));
  not_8  g11102(.A(new_n13450), .Y(new_n13451));
  xnor_4 g11103(.A(new_n13445), .B(new_n13435), .Y(new_n13452));
  nor_5  g11104(.A(new_n13452), .B(new_n13451), .Y(new_n13453));
  xor_4  g11105(.A(new_n13452), .B(new_n13450), .Y(new_n13454));
  xor_4  g11106(.A(new_n13442), .B(new_n13441), .Y(new_n13455));
  not_8  g11107(.A(new_n9858), .Y(new_n13456));
  nor_5  g11108(.A(new_n9859), .B(new_n13456), .Y(new_n13457));
  nand_5 g11109(.A(new_n13439), .B(new_n13412), .Y(new_n13458));
  nor_5  g11110(.A(new_n13458), .B(new_n13457), .Y(new_n13459));
  nor_5  g11111(.A(new_n9860), .B(new_n13456), .Y(new_n13460));
  not_8  g11112(.A(new_n13460), .Y(new_n13461));
  nand_5 g11113(.A(new_n13438), .B(new_n13456), .Y(new_n13462));
  nand_5 g11114(.A(new_n13462), .B(new_n13461), .Y(new_n13463));
  not_8  g11115(.A(new_n13463), .Y(new_n13464));
  xor_4  g11116(.A(new_n13439), .B(new_n13411), .Y(new_n13465));
  and_6  g11117(.A(new_n13465), .B(new_n13464), .Y(new_n13466));
  nand_5 g11118(.A(new_n13461), .B(new_n13440), .Y(new_n13467));
  nor_5  g11119(.A(new_n13467), .B(new_n13466), .Y(new_n13468));
  nor_5  g11120(.A(new_n13468), .B(new_n13459), .Y(new_n13469));
  nand_5 g11121(.A(new_n13469), .B(new_n13455), .Y(new_n13470));
  xor_4  g11122(.A(new_n13419), .B(new_n13418), .Y(new_n13471));
  xor_4  g11123(.A(new_n13469), .B(new_n13455), .Y(new_n13472));
  nand_5 g11124(.A(new_n13472), .B(new_n13471), .Y(new_n13473));
  nand_5 g11125(.A(new_n13473), .B(new_n13470), .Y(new_n13474));
  nor_5  g11126(.A(new_n13474), .B(new_n13454), .Y(new_n13475));
  nor_5  g11127(.A(new_n13475), .B(new_n13453), .Y(new_n13476));
  not_8  g11128(.A(new_n13432), .Y(new_n13477));
  xor_4  g11129(.A(new_n13448), .B(new_n13477), .Y(new_n13478));
  nor_5  g11130(.A(new_n13478), .B(new_n13476), .Y(new_n13479));
  or_6   g11131(.A(new_n13479), .B(new_n13449), .Y(new_n13480));
  nand_5 g11132(.A(new_n7010), .B(pi557), .Y(new_n13481));
  nand_5 g11133(.A(new_n13447), .B(new_n13433), .Y(new_n13482));
  nand_5 g11134(.A(new_n13482), .B(new_n13481), .Y(new_n13483));
  nand_5 g11135(.A(pi026), .B(new_n8336), .Y(new_n13484));
  not_8  g11136(.A(pi026), .Y(new_n13485));
  nand_5 g11137(.A(new_n13485), .B(pi004), .Y(new_n13486));
  nand_5 g11138(.A(new_n13486), .B(new_n13484), .Y(new_n13487));
  xnor_4 g11139(.A(new_n13487), .B(new_n13483), .Y(new_n13488));
  xnor_4 g11140(.A(new_n13488), .B(new_n13480), .Y(new_n13489));
  xor_4  g11141(.A(new_n13489), .B(new_n13430), .Y(po0115));
  nand_5 g11142(.A(new_n3026), .B(pi447), .Y(new_n13491));
  or_6   g11143(.A(new_n13491), .B(new_n2869), .Y(new_n13492));
  xor_4  g11144(.A(new_n13491), .B(new_n2869), .Y(new_n13493));
  nand_5 g11145(.A(new_n13493), .B(new_n3014), .Y(new_n13494));
  nand_5 g11146(.A(new_n13494), .B(new_n13492), .Y(new_n13495));
  nand_5 g11147(.A(new_n13495), .B(new_n3006), .Y(new_n13496));
  xor_4  g11148(.A(new_n13495), .B(new_n3006), .Y(new_n13497));
  nand_5 g11149(.A(new_n13497), .B(pi558), .Y(new_n13498));
  nand_5 g11150(.A(new_n13498), .B(new_n13496), .Y(new_n13499));
  nor_5  g11151(.A(new_n13499), .B(new_n3000), .Y(new_n13500));
  xor_4  g11152(.A(new_n13499), .B(new_n3001), .Y(new_n13501));
  nor_5  g11153(.A(new_n13501), .B(pi116), .Y(new_n13502));
  or_6   g11154(.A(new_n13502), .B(new_n13500), .Y(new_n13503));
  xor_4  g11155(.A(new_n13503), .B(new_n2995), .Y(new_n13504));
  xor_4  g11156(.A(new_n13504), .B(pi407), .Y(new_n13505));
  xor_4  g11157(.A(new_n13505), .B(new_n11570), .Y(new_n13506));
  xor_4  g11158(.A(new_n13501), .B(new_n2864), .Y(new_n13507));
  and_6  g11159(.A(new_n13507), .B(new_n9676), .Y(new_n13508));
  xnor_4 g11160(.A(new_n13507), .B(new_n9676), .Y(new_n13509));
  nand_5 g11161(.A(new_n3021), .B(new_n2747), .Y(new_n13510));
  xor_4  g11162(.A(new_n3021), .B(pi025), .Y(new_n13511));
  or_6   g11163(.A(new_n13511), .B(new_n7251), .Y(new_n13512));
  nand_5 g11164(.A(new_n13512), .B(new_n13510), .Y(new_n13513));
  xor_4  g11165(.A(new_n3025), .B(new_n2875), .Y(new_n13514));
  not_8  g11166(.A(new_n13514), .Y(new_n13515));
  nor_5  g11167(.A(new_n13515), .B(new_n13513), .Y(new_n13516));
  xor_4  g11168(.A(new_n13514), .B(new_n13513), .Y(new_n13517));
  nor_5  g11169(.A(new_n13517), .B(new_n9681), .Y(new_n13518));
  or_6   g11170(.A(new_n13518), .B(new_n13516), .Y(new_n13519));
  xor_4  g11171(.A(new_n13493), .B(new_n3011), .Y(new_n13520));
  not_8  g11172(.A(new_n13520), .Y(new_n13521));
  nor_5  g11173(.A(new_n13521), .B(new_n13519), .Y(new_n13522));
  xor_4  g11174(.A(new_n13520), .B(new_n13519), .Y(new_n13523));
  nor_5  g11175(.A(new_n13523), .B(new_n9688), .Y(new_n13524));
  or_6   g11176(.A(new_n13524), .B(new_n13522), .Y(new_n13525));
  xor_4  g11177(.A(new_n13497), .B(new_n2867), .Y(new_n13526));
  nand_5 g11178(.A(new_n13526), .B(new_n13525), .Y(new_n13527));
  xor_4  g11179(.A(new_n13526), .B(new_n13525), .Y(new_n13528));
  nand_5 g11180(.A(new_n13528), .B(new_n12153), .Y(new_n13529));
  nand_5 g11181(.A(new_n13529), .B(new_n13527), .Y(new_n13530));
  nor_5  g11182(.A(new_n13530), .B(new_n13509), .Y(new_n13531));
  nor_5  g11183(.A(new_n13531), .B(new_n13508), .Y(new_n13532));
  xnor_4 g11184(.A(new_n13532), .B(new_n13506), .Y(po0116));
  xnor_4 g11185(.A(new_n12056), .B(new_n12031), .Y(po0117));
  not_8  g11186(.A(new_n10005), .Y(new_n13535));
  nand_5 g11187(.A(new_n10861), .B(pi411), .Y(new_n13536));
  not_8  g11188(.A(pi411), .Y(new_n13537));
  nand_5 g11189(.A(new_n10929), .B(new_n13537), .Y(new_n13538));
  nand_5 g11190(.A(new_n13538), .B(new_n13536), .Y(new_n13539));
  not_8  g11191(.A(new_n13539), .Y(new_n13540));
  nand_5 g11192(.A(new_n13540), .B(new_n10008), .Y(new_n13541));
  not_8  g11193(.A(new_n13541), .Y(new_n13542));
  not_8  g11194(.A(new_n13536), .Y(new_n13543));
  not_8  g11195(.A(pi389), .Y(new_n13544));
  xor_4  g11196(.A(new_n10863), .B(new_n13544), .Y(new_n13545));
  xor_4  g11197(.A(new_n13545), .B(new_n13543), .Y(new_n13546));
  xor_4  g11198(.A(new_n13546), .B(new_n13542), .Y(new_n13547));
  xor_4  g11199(.A(new_n13547), .B(new_n13535), .Y(po0118));
  nand_5 g11200(.A(pi118), .B(new_n3424), .Y(new_n13549));
  nand_5 g11201(.A(new_n3469), .B(new_n3425), .Y(new_n13550));
  nand_5 g11202(.A(new_n13550), .B(new_n13549), .Y(new_n13551));
  not_8  g11203(.A(new_n13551), .Y(new_n13552));
  not_8  g11204(.A(new_n5875), .Y(new_n13553));
  xor_4  g11205(.A(pi458), .B(pi094), .Y(new_n13554));
  or_6   g11206(.A(pi288), .B(pi020), .Y(new_n13555));
  not_8  g11207(.A(pi559), .Y(new_n13556));
  nand_5 g11208(.A(pi288), .B(pi020), .Y(new_n13557));
  nand_5 g11209(.A(new_n13557), .B(new_n13556), .Y(new_n13558));
  nand_5 g11210(.A(new_n13558), .B(new_n13555), .Y(new_n13559));
  xor_4  g11211(.A(new_n13559), .B(new_n13554), .Y(new_n13560));
  or_6   g11212(.A(new_n13560), .B(new_n13553), .Y(new_n13561));
  nand_5 g11213(.A(new_n13560), .B(new_n13553), .Y(new_n13562));
  nor_5  g11214(.A(pi559), .B(pi299), .Y(new_n13563));
  nand_5 g11215(.A(new_n13563), .B(new_n6024), .Y(new_n13564));
  nor_5  g11216(.A(new_n13556), .B(new_n10978), .Y(new_n13565));
  nand_5 g11217(.A(new_n13565), .B(new_n6026), .Y(new_n13566));
  nand_5 g11218(.A(new_n13566), .B(new_n13564), .Y(new_n13567));
  and_6  g11219(.A(new_n13557), .B(new_n13555), .Y(new_n13568));
  xor_4  g11220(.A(new_n13568), .B(new_n5871), .Y(new_n13569));
  or_6   g11221(.A(new_n13569), .B(new_n13567), .Y(new_n13570));
  nand_5 g11222(.A(new_n13570), .B(new_n5871), .Y(new_n13571));
  nor_5  g11223(.A(new_n13567), .B(new_n13556), .Y(new_n13572));
  nor_5  g11224(.A(new_n13568), .B(new_n13564), .Y(new_n13573));
  nor_5  g11225(.A(new_n13573), .B(new_n13572), .Y(new_n13574));
  nand_5 g11226(.A(new_n13574), .B(new_n13571), .Y(new_n13575));
  xor_4  g11227(.A(new_n13569), .B(new_n13567), .Y(new_n13576));
  or_6   g11228(.A(new_n13568), .B(new_n13556), .Y(new_n13577));
  or_6   g11229(.A(new_n13577), .B(new_n13576), .Y(new_n13578));
  nand_5 g11230(.A(new_n13578), .B(new_n13575), .Y(new_n13579));
  nand_5 g11231(.A(new_n13579), .B(new_n13562), .Y(new_n13580));
  nand_5 g11232(.A(new_n13580), .B(new_n13561), .Y(new_n13581));
  not_8  g11233(.A(new_n5870), .Y(new_n13582));
  xor_4  g11234(.A(pi450), .B(pi152), .Y(new_n13583));
  nand_5 g11235(.A(new_n3581), .B(new_n13257), .Y(new_n13584));
  nand_5 g11236(.A(new_n13559), .B(new_n13554), .Y(new_n13585));
  nand_5 g11237(.A(new_n13585), .B(new_n13584), .Y(new_n13586));
  xor_4  g11238(.A(new_n13586), .B(new_n13583), .Y(new_n13587));
  nand_5 g11239(.A(new_n13587), .B(new_n13582), .Y(new_n13588));
  or_6   g11240(.A(new_n13587), .B(new_n13582), .Y(new_n13589));
  nand_5 g11241(.A(new_n13589), .B(new_n13588), .Y(new_n13590));
  xor_4  g11242(.A(new_n13590), .B(new_n13581), .Y(new_n13591));
  not_8  g11243(.A(new_n13591), .Y(new_n13592));
  nor_5  g11244(.A(new_n13592), .B(new_n3488), .Y(new_n13593));
  xor_4  g11245(.A(new_n13591), .B(new_n3488), .Y(new_n13594));
  not_8  g11246(.A(new_n3490), .Y(new_n13595));
  nand_5 g11247(.A(new_n3492), .B(new_n3449), .Y(new_n13596));
  nor_5  g11248(.A(new_n13565), .B(new_n13563), .Y(new_n13597));
  xor_4  g11249(.A(new_n13597), .B(new_n6026), .Y(new_n13598));
  nand_5 g11250(.A(new_n13598), .B(new_n13596), .Y(new_n13599));
  nand_5 g11251(.A(new_n13599), .B(new_n13595), .Y(new_n13600));
  xor_4  g11252(.A(new_n13599), .B(new_n13595), .Y(new_n13601));
  nand_5 g11253(.A(new_n13601), .B(new_n13576), .Y(new_n13602));
  nand_5 g11254(.A(new_n13602), .B(new_n13600), .Y(new_n13603));
  nand_5 g11255(.A(new_n13603), .B(new_n3501), .Y(new_n13604));
  nand_5 g11256(.A(new_n13562), .B(new_n13561), .Y(new_n13605));
  xnor_4 g11257(.A(new_n13605), .B(new_n13579), .Y(new_n13606));
  xor_4  g11258(.A(new_n13603), .B(new_n3501), .Y(new_n13607));
  nand_5 g11259(.A(new_n13607), .B(new_n13606), .Y(new_n13608));
  nand_5 g11260(.A(new_n13608), .B(new_n13604), .Y(new_n13609));
  nor_5  g11261(.A(new_n13609), .B(new_n13594), .Y(new_n13610));
  or_6   g11262(.A(new_n13610), .B(new_n13593), .Y(new_n13611));
  nand_5 g11263(.A(new_n13588), .B(new_n13581), .Y(new_n13612));
  nand_5 g11264(.A(new_n13612), .B(new_n13589), .Y(new_n13613));
  xor_4  g11265(.A(pi536), .B(pi037), .Y(new_n13614));
  not_8  g11266(.A(pi450), .Y(new_n13615));
  nand_5 g11267(.A(new_n13615), .B(new_n3656), .Y(new_n13616));
  nand_5 g11268(.A(new_n13586), .B(new_n13583), .Y(new_n13617));
  nand_5 g11269(.A(new_n13617), .B(new_n13616), .Y(new_n13618));
  xnor_4 g11270(.A(new_n13618), .B(new_n13614), .Y(new_n13619));
  xor_4  g11271(.A(new_n13619), .B(new_n5866), .Y(new_n13620));
  xnor_4 g11272(.A(new_n13620), .B(new_n13613), .Y(new_n13621));
  nor_5  g11273(.A(new_n13621), .B(new_n13611), .Y(new_n13622));
  or_6   g11274(.A(new_n13622), .B(new_n3487), .Y(new_n13623));
  nand_5 g11275(.A(new_n13621), .B(new_n13611), .Y(new_n13624));
  nand_5 g11276(.A(new_n13624), .B(new_n13623), .Y(new_n13625));
  not_8  g11277(.A(new_n5865), .Y(new_n13626));
  xor_4  g11278(.A(pi585), .B(pi493), .Y(new_n13627));
  nand_5 g11279(.A(new_n12720), .B(new_n3598), .Y(new_n13628));
  nand_5 g11280(.A(new_n13618), .B(new_n13614), .Y(new_n13629));
  nand_5 g11281(.A(new_n13629), .B(new_n13628), .Y(new_n13630));
  xor_4  g11282(.A(new_n13630), .B(new_n13627), .Y(new_n13631));
  xor_4  g11283(.A(new_n13631), .B(new_n13626), .Y(new_n13632));
  nand_5 g11284(.A(new_n13619), .B(new_n5866), .Y(new_n13633));
  nand_5 g11285(.A(new_n13620), .B(new_n13613), .Y(new_n13634));
  nand_5 g11286(.A(new_n13634), .B(new_n13633), .Y(new_n13635));
  xor_4  g11287(.A(new_n13635), .B(new_n13632), .Y(new_n13636));
  not_8  g11288(.A(new_n13636), .Y(new_n13637));
  nand_5 g11289(.A(new_n13637), .B(new_n13625), .Y(new_n13638));
  xor_4  g11290(.A(new_n13636), .B(new_n13625), .Y(new_n13639));
  or_6   g11291(.A(new_n13639), .B(new_n3482), .Y(new_n13640));
  nand_5 g11292(.A(new_n13640), .B(new_n13638), .Y(new_n13641));
  xor_4  g11293(.A(pi717), .B(pi526), .Y(new_n13642));
  not_8  g11294(.A(pi493), .Y(new_n13643));
  nand_5 g11295(.A(new_n3604), .B(new_n13643), .Y(new_n13644));
  nand_5 g11296(.A(new_n13630), .B(new_n13627), .Y(new_n13645));
  nand_5 g11297(.A(new_n13645), .B(new_n13644), .Y(new_n13646));
  xnor_4 g11298(.A(new_n13646), .B(new_n13642), .Y(new_n13647));
  xor_4  g11299(.A(new_n13647), .B(new_n5900), .Y(new_n13648));
  nand_5 g11300(.A(new_n13631), .B(new_n13626), .Y(new_n13649));
  not_8  g11301(.A(new_n13649), .Y(new_n13650));
  not_8  g11302(.A(new_n13632), .Y(new_n13651));
  nor_5  g11303(.A(new_n13635), .B(new_n13651), .Y(new_n13652));
  nor_5  g11304(.A(new_n13652), .B(new_n13650), .Y(new_n13653));
  xor_4  g11305(.A(new_n13653), .B(new_n13648), .Y(new_n13654));
  not_8  g11306(.A(new_n13654), .Y(new_n13655));
  or_6   g11307(.A(new_n13655), .B(new_n13641), .Y(new_n13656));
  xor_4  g11308(.A(new_n13655), .B(new_n13641), .Y(new_n13657));
  nand_5 g11309(.A(new_n13657), .B(new_n3480), .Y(new_n13658));
  nand_5 g11310(.A(new_n13658), .B(new_n13656), .Y(new_n13659));
  xor_4  g11311(.A(pi624), .B(pi409), .Y(new_n13660));
  nand_5 g11312(.A(new_n3611), .B(new_n12777), .Y(new_n13661));
  nand_5 g11313(.A(new_n13646), .B(new_n13642), .Y(new_n13662));
  nand_5 g11314(.A(new_n13662), .B(new_n13661), .Y(new_n13663));
  xor_4  g11315(.A(new_n13663), .B(new_n13660), .Y(new_n13664));
  xor_4  g11316(.A(new_n13664), .B(new_n5907), .Y(new_n13665));
  or_6   g11317(.A(new_n13647), .B(new_n5900), .Y(new_n13666));
  not_8  g11318(.A(new_n13653), .Y(new_n13667));
  nand_5 g11319(.A(new_n13667), .B(new_n13648), .Y(new_n13668));
  nand_5 g11320(.A(new_n13668), .B(new_n13666), .Y(new_n13669));
  xor_4  g11321(.A(new_n13669), .B(new_n13665), .Y(new_n13670));
  not_8  g11322(.A(new_n13670), .Y(new_n13671));
  nor_5  g11323(.A(new_n13671), .B(new_n13659), .Y(new_n13672));
  xor_4  g11324(.A(new_n13670), .B(new_n13659), .Y(new_n13673));
  nor_5  g11325(.A(new_n13673), .B(new_n3477), .Y(new_n13674));
  or_6   g11326(.A(new_n13674), .B(new_n13672), .Y(new_n13675));
  nand_5 g11327(.A(new_n13675), .B(new_n3475), .Y(new_n13676));
  xor_4  g11328(.A(new_n13675), .B(new_n3474), .Y(new_n13677));
  nand_5 g11329(.A(new_n13664), .B(new_n5907), .Y(new_n13678));
  nand_5 g11330(.A(new_n13669), .B(new_n13665), .Y(new_n13679));
  nand_5 g11331(.A(new_n13679), .B(new_n13678), .Y(new_n13680));
  xor_4  g11332(.A(pi740), .B(pi412), .Y(new_n13681));
  nand_5 g11333(.A(new_n12795), .B(new_n3622), .Y(new_n13682));
  nand_5 g11334(.A(new_n13663), .B(new_n13660), .Y(new_n13683));
  nand_5 g11335(.A(new_n13683), .B(new_n13682), .Y(new_n13684));
  xor_4  g11336(.A(new_n13684), .B(new_n13681), .Y(new_n13685));
  xor_4  g11337(.A(new_n13685), .B(new_n5924), .Y(new_n13686));
  xor_4  g11338(.A(new_n13686), .B(new_n13680), .Y(new_n13687));
  or_6   g11339(.A(new_n13687), .B(new_n13677), .Y(new_n13688));
  nand_5 g11340(.A(new_n13688), .B(new_n13676), .Y(new_n13689));
  nor_5  g11341(.A(new_n13689), .B(new_n3470), .Y(new_n13690));
  nor_5  g11342(.A(new_n13685), .B(new_n5925), .Y(new_n13691));
  or_6   g11343(.A(new_n13686), .B(new_n13680), .Y(new_n13692));
  not_8  g11344(.A(new_n13692), .Y(new_n13693));
  nor_5  g11345(.A(new_n13693), .B(new_n13691), .Y(new_n13694));
  xor_4  g11346(.A(new_n13694), .B(new_n5935), .Y(new_n13695));
  nand_5 g11347(.A(new_n3524), .B(new_n12812), .Y(new_n13696));
  nand_5 g11348(.A(new_n13684), .B(new_n13681), .Y(new_n13697));
  nand_5 g11349(.A(new_n13697), .B(new_n13696), .Y(new_n13698));
  nand_5 g11350(.A(pi807), .B(pi345), .Y(new_n13699));
  nand_5 g11351(.A(new_n8441), .B(new_n13030), .Y(new_n13700));
  nand_5 g11352(.A(new_n13700), .B(new_n13699), .Y(new_n13701));
  xor_4  g11353(.A(new_n13701), .B(new_n13698), .Y(new_n13702));
  xor_4  g11354(.A(new_n13702), .B(new_n13695), .Y(new_n13703));
  xor_4  g11355(.A(new_n13689), .B(new_n3470), .Y(new_n13704));
  not_8  g11356(.A(new_n13704), .Y(new_n13705));
  nor_5  g11357(.A(new_n13705), .B(new_n13703), .Y(new_n13706));
  or_6   g11358(.A(new_n13706), .B(new_n13690), .Y(new_n13707));
  nor_5  g11359(.A(new_n13707), .B(new_n13552), .Y(new_n13708));
  xor_4  g11360(.A(new_n13707), .B(new_n13551), .Y(new_n13709));
  not_8  g11361(.A(new_n5935), .Y(new_n13710));
  nand_5 g11362(.A(new_n13694), .B(new_n13710), .Y(new_n13711));
  not_8  g11363(.A(new_n13711), .Y(new_n13712));
  nor_5  g11364(.A(new_n13702), .B(new_n13695), .Y(new_n13713));
  nor_5  g11365(.A(new_n13713), .B(new_n13712), .Y(new_n13714));
  nand_5 g11366(.A(new_n13699), .B(new_n13698), .Y(new_n13715));
  nand_5 g11367(.A(new_n13715), .B(new_n13700), .Y(new_n13716));
  nand_5 g11368(.A(new_n5933), .B(new_n5928), .Y(new_n13717));
  nand_5 g11369(.A(new_n13717), .B(new_n5930), .Y(new_n13718));
  not_8  g11370(.A(new_n13718), .Y(new_n13719));
  xor_4  g11371(.A(new_n13719), .B(new_n13716), .Y(new_n13720));
  xor_4  g11372(.A(new_n13720), .B(new_n13714), .Y(new_n13721));
  nor_5  g11373(.A(new_n13721), .B(new_n13709), .Y(new_n13722));
  nor_5  g11374(.A(new_n13722), .B(new_n13708), .Y(new_n13723));
  or_6   g11375(.A(new_n13719), .B(new_n13716), .Y(new_n13724));
  nand_5 g11376(.A(new_n13720), .B(new_n13714), .Y(new_n13725));
  nand_5 g11377(.A(new_n13725), .B(new_n13724), .Y(new_n13726));
  xor_4  g11378(.A(new_n13726), .B(new_n13723), .Y(po0119));
  xor_4  g11379(.A(new_n8492), .B(new_n5158), .Y(po0120));
  nand_5 g11380(.A(new_n8019), .B(pi212), .Y(new_n13729));
  not_8  g11381(.A(new_n9902), .Y(new_n13730));
  nand_5 g11382(.A(pi620), .B(new_n8027), .Y(new_n13731));
  not_8  g11383(.A(new_n9931), .Y(new_n13732));
  nand_5 g11384(.A(new_n13732), .B(new_n9927), .Y(new_n13733));
  nand_5 g11385(.A(new_n13733), .B(new_n13731), .Y(new_n13734));
  nand_5 g11386(.A(new_n13734), .B(new_n13730), .Y(new_n13735));
  nand_5 g11387(.A(new_n13735), .B(new_n13729), .Y(new_n13736));
  xor_4  g11388(.A(new_n13736), .B(new_n9899), .Y(new_n13737));
  xor_4  g11389(.A(pi558), .B(new_n2718), .Y(new_n13738));
  nand_5 g11390(.A(pi521), .B(new_n2869), .Y(new_n13739));
  not_8  g11391(.A(new_n13739), .Y(new_n13740));
  xor_4  g11392(.A(pi521), .B(pi231), .Y(new_n13741));
  nand_5 g11393(.A(pi447), .B(new_n10243), .Y(new_n13742));
  nand_5 g11394(.A(new_n2875), .B(pi370), .Y(new_n13743));
  nand_5 g11395(.A(pi544), .B(new_n2747), .Y(new_n13744));
  nand_5 g11396(.A(new_n13744), .B(new_n13743), .Y(new_n13745));
  nand_5 g11397(.A(new_n13745), .B(new_n13742), .Y(new_n13746));
  nor_5  g11398(.A(new_n13746), .B(new_n13741), .Y(new_n13747));
  nor_5  g11399(.A(new_n13747), .B(new_n13740), .Y(new_n13748));
  xor_4  g11400(.A(new_n13748), .B(new_n13738), .Y(new_n13749));
  xor_4  g11401(.A(new_n13749), .B(new_n13737), .Y(new_n13750));
  xor_4  g11402(.A(new_n13734), .B(new_n9902), .Y(new_n13751));
  not_8  g11403(.A(new_n13751), .Y(new_n13752));
  xor_4  g11404(.A(new_n13746), .B(new_n13741), .Y(new_n13753));
  nand_5 g11405(.A(new_n13753), .B(new_n13752), .Y(new_n13754));
  nand_5 g11406(.A(new_n2746), .B(pi025), .Y(new_n13755));
  and_6  g11407(.A(new_n13743), .B(new_n13742), .Y(new_n13756));
  nor_5  g11408(.A(new_n13756), .B(new_n13755), .Y(new_n13757));
  nand_5 g11409(.A(new_n13756), .B(new_n13755), .Y(new_n13758));
  nand_5 g11410(.A(new_n13758), .B(new_n9932), .Y(new_n13759));
  nor_5  g11411(.A(new_n13759), .B(new_n13757), .Y(new_n13760));
  nor_5  g11412(.A(new_n13760), .B(new_n9935), .Y(new_n13761));
  nor_5  g11413(.A(new_n13761), .B(new_n9926), .Y(new_n13762));
  nand_5 g11414(.A(new_n13755), .B(new_n13744), .Y(new_n13763));
  nand_5 g11415(.A(new_n13763), .B(new_n9935), .Y(new_n13764));
  nand_5 g11416(.A(new_n13764), .B(new_n9931), .Y(new_n13765));
  nand_5 g11417(.A(new_n13765), .B(new_n13755), .Y(new_n13766));
  or_6   g11418(.A(new_n13756), .B(new_n9927), .Y(new_n13767));
  or_6   g11419(.A(new_n13767), .B(new_n13766), .Y(new_n13768));
  nand_5 g11420(.A(new_n9933), .B(new_n2746), .Y(new_n13769));
  or_6   g11421(.A(new_n13769), .B(new_n9927), .Y(new_n13770));
  nand_5 g11422(.A(new_n13770), .B(new_n13763), .Y(new_n13771));
  nand_5 g11423(.A(new_n13771), .B(new_n13756), .Y(new_n13772));
  nand_5 g11424(.A(new_n13772), .B(new_n13768), .Y(new_n13773));
  or_6   g11425(.A(new_n13773), .B(new_n13762), .Y(new_n13774));
  xor_4  g11426(.A(new_n13753), .B(new_n13751), .Y(new_n13775));
  not_8  g11427(.A(new_n13775), .Y(new_n13776));
  nand_5 g11428(.A(new_n13776), .B(new_n13774), .Y(new_n13777));
  nand_5 g11429(.A(new_n13777), .B(new_n13754), .Y(new_n13778));
  xor_4  g11430(.A(new_n13778), .B(new_n13750), .Y(new_n13779));
  and_6  g11431(.A(pi693), .B(new_n4133), .Y(new_n13780));
  xor_4  g11432(.A(pi693), .B(new_n4133), .Y(new_n13781));
  not_8  g11433(.A(new_n13781), .Y(new_n13782));
  nand_5 g11434(.A(new_n13544), .B(pi215), .Y(new_n13783));
  nand_5 g11435(.A(pi389), .B(new_n4139), .Y(new_n13784));
  nand_5 g11436(.A(new_n4204), .B(pi411), .Y(new_n13785));
  nand_5 g11437(.A(new_n13785), .B(new_n13784), .Y(new_n13786));
  nand_5 g11438(.A(new_n13786), .B(new_n13783), .Y(new_n13787));
  nor_5  g11439(.A(new_n13787), .B(new_n13782), .Y(new_n13788));
  nor_5  g11440(.A(new_n13788), .B(new_n13780), .Y(new_n13789));
  xor_4  g11441(.A(pi591), .B(pi524), .Y(new_n13790));
  xor_4  g11442(.A(new_n13790), .B(new_n13789), .Y(new_n13791));
  xor_4  g11443(.A(new_n13791), .B(new_n13779), .Y(new_n13792));
  xor_4  g11444(.A(new_n13776), .B(new_n13774), .Y(new_n13793));
  xor_4  g11445(.A(new_n13787), .B(new_n13781), .Y(new_n13794));
  not_8  g11446(.A(new_n13794), .Y(new_n13795));
  or_6   g11447(.A(new_n13795), .B(new_n13793), .Y(new_n13796));
  xor_4  g11448(.A(new_n13795), .B(new_n13793), .Y(new_n13797));
  not_8  g11449(.A(new_n13763), .Y(new_n13798));
  xor_4  g11450(.A(new_n13798), .B(new_n9934), .Y(new_n13799));
  xor_4  g11451(.A(pi758), .B(new_n13537), .Y(new_n13800));
  nor_5  g11452(.A(new_n13800), .B(new_n13799), .Y(new_n13801));
  and_6  g11453(.A(new_n13784), .B(new_n13783), .Y(new_n13802));
  xor_4  g11454(.A(new_n13802), .B(new_n13785), .Y(new_n13803));
  nor_5  g11455(.A(new_n13803), .B(new_n13801), .Y(new_n13804));
  or_6   g11456(.A(new_n13755), .B(new_n9933), .Y(new_n13805));
  nand_5 g11457(.A(new_n13805), .B(new_n13766), .Y(new_n13806));
  xor_4  g11458(.A(new_n13756), .B(new_n9927), .Y(new_n13807));
  xor_4  g11459(.A(new_n13807), .B(new_n13806), .Y(new_n13808));
  not_8  g11460(.A(new_n13803), .Y(new_n13809));
  xor_4  g11461(.A(new_n13809), .B(new_n13801), .Y(new_n13810));
  nor_5  g11462(.A(new_n13810), .B(new_n13808), .Y(new_n13811));
  nor_5  g11463(.A(new_n13811), .B(new_n13804), .Y(new_n13812));
  nand_5 g11464(.A(new_n13812), .B(new_n13797), .Y(new_n13813));
  nand_5 g11465(.A(new_n13813), .B(new_n13796), .Y(new_n13814));
  xor_4  g11466(.A(new_n13814), .B(new_n13792), .Y(po0121));
  nand_5 g11467(.A(new_n7974), .B(new_n7984), .Y(new_n13816));
  xor_4  g11468(.A(new_n13816), .B(new_n7977), .Y(new_n13817));
  not_8  g11469(.A(new_n13817), .Y(new_n13818));
  nand_5 g11470(.A(new_n13818), .B(new_n7974), .Y(new_n13819));
  nand_5 g11471(.A(new_n13819), .B(new_n7984), .Y(new_n13820));
  not_8  g11472(.A(new_n13820), .Y(new_n13821));
  nand_5 g11473(.A(new_n13821), .B(new_n11890), .Y(new_n13822));
  nand_5 g11474(.A(new_n13820), .B(new_n11871), .Y(new_n13823));
  nand_5 g11475(.A(new_n7997), .B(new_n7874), .Y(new_n13824));
  nand_5 g11476(.A(new_n7978), .B(new_n4858), .Y(new_n13825));
  nor_5  g11477(.A(new_n13825), .B(new_n7973), .Y(new_n13826));
  nor_5  g11478(.A(new_n13819), .B(new_n7983), .Y(new_n13827));
  nor_5  g11479(.A(new_n13827), .B(new_n13826), .Y(new_n13828));
  nand_5 g11480(.A(new_n13828), .B(new_n13824), .Y(new_n13829));
  nand_5 g11481(.A(new_n13829), .B(new_n13823), .Y(new_n13830));
  nand_5 g11482(.A(new_n13830), .B(new_n13822), .Y(po0122));
  xor_4  g11483(.A(new_n4221), .B(new_n4219), .Y(po0123));
  nand_5 g11484(.A(new_n2566), .B(pi677), .Y(new_n13833));
  nor_5  g11485(.A(new_n13833), .B(new_n8163), .Y(new_n13834));
  xor_4  g11486(.A(new_n13833), .B(new_n8163), .Y(new_n13835));
  not_8  g11487(.A(new_n13835), .Y(new_n13836));
  nor_5  g11488(.A(new_n13836), .B(new_n3927), .Y(new_n13837));
  or_6   g11489(.A(new_n13837), .B(new_n13834), .Y(new_n13838));
  nor_5  g11490(.A(new_n13838), .B(new_n3921), .Y(new_n13839));
  xor_4  g11491(.A(new_n13838), .B(new_n3920), .Y(new_n13840));
  nor_5  g11492(.A(new_n13840), .B(pi754), .Y(new_n13841));
  or_6   g11493(.A(new_n13841), .B(new_n13839), .Y(new_n13842));
  nand_5 g11494(.A(new_n13842), .B(new_n8158), .Y(new_n13843));
  xor_4  g11495(.A(new_n13842), .B(new_n8158), .Y(new_n13844));
  nand_5 g11496(.A(new_n13844), .B(new_n3918), .Y(new_n13845));
  nand_5 g11497(.A(new_n13845), .B(new_n13843), .Y(new_n13846));
  or_6   g11498(.A(new_n13846), .B(new_n4051), .Y(new_n13847));
  nand_5 g11499(.A(new_n13847), .B(new_n8154), .Y(new_n13848));
  nand_5 g11500(.A(new_n13846), .B(new_n4051), .Y(new_n13849));
  nand_5 g11501(.A(new_n13849), .B(new_n13848), .Y(new_n13850));
  xor_4  g11502(.A(new_n13850), .B(new_n4049), .Y(new_n13851));
  xor_4  g11503(.A(new_n13851), .B(new_n8153), .Y(new_n13852));
  xor_4  g11504(.A(new_n8133), .B(new_n2556), .Y(new_n13853));
  nand_5 g11505(.A(new_n13853), .B(pi813), .Y(new_n13854));
  nand_5 g11506(.A(new_n13854), .B(new_n8018), .Y(new_n13855));
  xor_4  g11507(.A(new_n13854), .B(new_n8018), .Y(new_n13856));
  not_8  g11508(.A(new_n13856), .Y(new_n13857));
  or_6   g11509(.A(new_n13857), .B(new_n8179), .Y(new_n13858));
  nand_5 g11510(.A(new_n13858), .B(new_n13855), .Y(new_n13859));
  nand_5 g11511(.A(new_n13859), .B(new_n8159), .Y(new_n13860));
  or_6   g11512(.A(new_n13859), .B(new_n8159), .Y(new_n13861));
  nand_5 g11513(.A(new_n13861), .B(new_n4395), .Y(new_n13862));
  nand_5 g11514(.A(new_n13862), .B(new_n13860), .Y(new_n13863));
  nand_5 g11515(.A(new_n13863), .B(new_n8155), .Y(new_n13864));
  or_6   g11516(.A(new_n13863), .B(new_n8155), .Y(new_n13865));
  nand_5 g11517(.A(new_n13865), .B(new_n10744), .Y(new_n13866));
  nand_5 g11518(.A(new_n13866), .B(new_n13864), .Y(new_n13867));
  nand_5 g11519(.A(new_n13867), .B(new_n8188), .Y(new_n13868));
  or_6   g11520(.A(new_n13867), .B(new_n8188), .Y(new_n13869));
  nand_5 g11521(.A(new_n13869), .B(new_n13868), .Y(new_n13870));
  xor_4  g11522(.A(new_n13870), .B(pi248), .Y(new_n13871));
  xnor_4 g11523(.A(new_n13871), .B(new_n13852), .Y(new_n13872));
  nand_5 g11524(.A(new_n13849), .B(new_n13847), .Y(new_n13873));
  xor_4  g11525(.A(new_n13873), .B(pi398), .Y(new_n13874));
  nand_5 g11526(.A(new_n13865), .B(new_n13864), .Y(new_n13875));
  xor_4  g11527(.A(new_n13875), .B(pi125), .Y(new_n13876));
  not_8  g11528(.A(new_n13876), .Y(new_n13877));
  nand_5 g11529(.A(new_n13877), .B(new_n13874), .Y(new_n13878));
  xor_4  g11530(.A(new_n13876), .B(new_n13874), .Y(new_n13879));
  xor_4  g11531(.A(new_n13844), .B(new_n3919), .Y(new_n13880));
  nand_5 g11532(.A(new_n13861), .B(new_n13860), .Y(new_n13881));
  xor_4  g11533(.A(new_n13881), .B(pi618), .Y(new_n13882));
  nand_5 g11534(.A(new_n13882), .B(new_n13880), .Y(new_n13883));
  xnor_4 g11535(.A(new_n13882), .B(new_n13880), .Y(new_n13884));
  xor_4  g11536(.A(new_n13840), .B(new_n8162), .Y(new_n13885));
  xor_4  g11537(.A(new_n13856), .B(new_n8179), .Y(new_n13886));
  not_8  g11538(.A(new_n13886), .Y(new_n13887));
  nor_5  g11539(.A(new_n13887), .B(new_n13885), .Y(new_n13888));
  xor_4  g11540(.A(new_n2566), .B(pi677), .Y(new_n13889));
  nand_5 g11541(.A(new_n13889), .B(new_n4405), .Y(new_n13890));
  xor_4  g11542(.A(new_n13889), .B(new_n4405), .Y(new_n13891));
  nand_5 g11543(.A(new_n13891), .B(new_n2561), .Y(new_n13892));
  nand_5 g11544(.A(new_n13892), .B(new_n13890), .Y(new_n13893));
  xor_4  g11545(.A(new_n8133), .B(pi813), .Y(new_n13894));
  nand_5 g11546(.A(new_n13890), .B(new_n2557), .Y(new_n13895));
  nand_5 g11547(.A(new_n13893), .B(new_n2556), .Y(new_n13896));
  nand_5 g11548(.A(new_n13896), .B(new_n13895), .Y(new_n13897));
  xor_4  g11549(.A(new_n13897), .B(new_n13894), .Y(new_n13898));
  not_8  g11550(.A(new_n13898), .Y(new_n13899));
  nand_5 g11551(.A(new_n13899), .B(new_n13893), .Y(new_n13900));
  xor_4  g11552(.A(new_n13836), .B(new_n3927), .Y(new_n13901));
  nand_5 g11553(.A(new_n13901), .B(new_n13898), .Y(new_n13902));
  nand_5 g11554(.A(new_n13902), .B(new_n13900), .Y(new_n13903));
  xor_4  g11555(.A(new_n13886), .B(new_n13885), .Y(new_n13904));
  nor_5  g11556(.A(new_n13904), .B(new_n13903), .Y(new_n13905));
  or_6   g11557(.A(new_n13905), .B(new_n13888), .Y(new_n13906));
  or_6   g11558(.A(new_n13906), .B(new_n13884), .Y(new_n13907));
  nand_5 g11559(.A(new_n13907), .B(new_n13883), .Y(new_n13908));
  or_6   g11560(.A(new_n13908), .B(new_n13879), .Y(new_n13909));
  nand_5 g11561(.A(new_n13909), .B(new_n13878), .Y(new_n13910));
  xnor_4 g11562(.A(new_n13910), .B(new_n13872), .Y(po0124));
  nand_5 g11563(.A(new_n13030), .B(pi097), .Y(new_n13912));
  xor_4  g11564(.A(pi345), .B(new_n4857), .Y(new_n13913));
  nand_5 g11565(.A(new_n12812), .B(pi013), .Y(new_n13914));
  xor_4  g11566(.A(pi412), .B(new_n4838), .Y(new_n13915));
  nand_5 g11567(.A(new_n12795), .B(pi623), .Y(new_n13916));
  xor_4  g11568(.A(pi624), .B(new_n4843), .Y(new_n13917));
  nand_5 g11569(.A(pi793), .B(new_n12777), .Y(new_n13918));
  nand_5 g11570(.A(new_n13643), .B(pi103), .Y(new_n13919));
  xor_4  g11571(.A(pi493), .B(new_n4756), .Y(new_n13920));
  nand_5 g11572(.A(new_n12720), .B(pi298), .Y(new_n13921));
  xor_4  g11573(.A(pi536), .B(new_n3763), .Y(new_n13922));
  nand_5 g11574(.A(new_n13615), .B(pi157), .Y(new_n13923));
  nand_5 g11575(.A(new_n13276), .B(new_n13273), .Y(new_n13924));
  nand_5 g11576(.A(new_n13924), .B(new_n13923), .Y(new_n13925));
  nand_5 g11577(.A(new_n13925), .B(new_n13922), .Y(new_n13926));
  nand_5 g11578(.A(new_n13926), .B(new_n13921), .Y(new_n13927));
  nand_5 g11579(.A(new_n13927), .B(new_n13920), .Y(new_n13928));
  nand_5 g11580(.A(new_n13928), .B(new_n13919), .Y(new_n13929));
  xor_4  g11581(.A(pi793), .B(pi526), .Y(new_n13930));
  not_8  g11582(.A(new_n13930), .Y(new_n13931));
  nand_5 g11583(.A(new_n13931), .B(new_n13929), .Y(new_n13932));
  nand_5 g11584(.A(new_n13932), .B(new_n13918), .Y(new_n13933));
  nand_5 g11585(.A(new_n13933), .B(new_n13917), .Y(new_n13934));
  nand_5 g11586(.A(new_n13934), .B(new_n13916), .Y(new_n13935));
  nand_5 g11587(.A(new_n13935), .B(new_n13915), .Y(new_n13936));
  nand_5 g11588(.A(new_n13936), .B(new_n13914), .Y(new_n13937));
  nand_5 g11589(.A(new_n13937), .B(new_n13913), .Y(new_n13938));
  nand_5 g11590(.A(new_n13938), .B(new_n13912), .Y(new_n13939));
  xor_4  g11591(.A(new_n13937), .B(new_n13913), .Y(new_n13940));
  not_8  g11592(.A(new_n13940), .Y(new_n13941));
  xor_4  g11593(.A(new_n13935), .B(new_n13915), .Y(new_n13942));
  not_8  g11594(.A(new_n13942), .Y(new_n13943));
  xor_4  g11595(.A(new_n13933), .B(new_n13917), .Y(new_n13944));
  not_8  g11596(.A(new_n13944), .Y(new_n13945));
  nand_5 g11597(.A(new_n13945), .B(pi823), .Y(new_n13946));
  xor_4  g11598(.A(new_n13944), .B(new_n5919), .Y(new_n13947));
  xor_4  g11599(.A(new_n13930), .B(new_n13929), .Y(new_n13948));
  not_8  g11600(.A(new_n13948), .Y(new_n13949));
  xor_4  g11601(.A(new_n13925), .B(new_n13922), .Y(new_n13950));
  nor_5  g11602(.A(new_n13277), .B(pi399), .Y(new_n13951));
  nor_5  g11603(.A(new_n13278), .B(new_n13272), .Y(new_n13952));
  or_6   g11604(.A(new_n13952), .B(new_n13951), .Y(new_n13953));
  or_6   g11605(.A(new_n13953), .B(new_n13950), .Y(new_n13954));
  xor_4  g11606(.A(new_n13953), .B(new_n13950), .Y(new_n13955));
  nand_5 g11607(.A(new_n13955), .B(pi254), .Y(new_n13956));
  nand_5 g11608(.A(new_n13956), .B(new_n13954), .Y(new_n13957));
  nor_5  g11609(.A(new_n13957), .B(pi106), .Y(new_n13958));
  xnor_4 g11610(.A(new_n13927), .B(new_n13920), .Y(new_n13959));
  xor_4  g11611(.A(new_n13957), .B(pi106), .Y(new_n13960));
  not_8  g11612(.A(new_n13960), .Y(new_n13961));
  nor_5  g11613(.A(new_n13961), .B(new_n13959), .Y(new_n13962));
  or_6   g11614(.A(new_n13962), .B(new_n13958), .Y(new_n13963));
  nand_5 g11615(.A(new_n13963), .B(new_n13949), .Y(new_n13964));
  not_8  g11616(.A(new_n13964), .Y(new_n13965));
  nor_5  g11617(.A(new_n13963), .B(new_n13949), .Y(new_n13966));
  nor_5  g11618(.A(new_n13966), .B(pi383), .Y(new_n13967));
  nor_5  g11619(.A(new_n13967), .B(new_n13965), .Y(new_n13968));
  nand_5 g11620(.A(new_n13968), .B(new_n13947), .Y(new_n13969));
  nand_5 g11621(.A(new_n13969), .B(new_n13946), .Y(new_n13970));
  or_6   g11622(.A(new_n13970), .B(new_n13943), .Y(new_n13971));
  nand_5 g11623(.A(new_n13971), .B(pi136), .Y(new_n13972));
  nand_5 g11624(.A(new_n13970), .B(new_n13943), .Y(new_n13973));
  nand_5 g11625(.A(new_n13973), .B(new_n13972), .Y(new_n13974));
  nand_5 g11626(.A(new_n13974), .B(new_n13941), .Y(new_n13975));
  or_6   g11627(.A(new_n13974), .B(new_n13941), .Y(new_n13976));
  nand_5 g11628(.A(new_n13976), .B(pi207), .Y(new_n13977));
  nand_5 g11629(.A(new_n13977), .B(new_n13975), .Y(new_n13978));
  nand_5 g11630(.A(new_n13978), .B(new_n13939), .Y(new_n13979));
  and_6  g11631(.A(new_n13979), .B(new_n13044), .Y(new_n13980));
  xor_4  g11632(.A(new_n13978), .B(new_n13939), .Y(new_n13981));
  nor_5  g11633(.A(new_n13981), .B(new_n13026), .Y(new_n13982));
  xor_4  g11634(.A(new_n13981), .B(new_n13026), .Y(new_n13983));
  nand_5 g11635(.A(new_n13976), .B(new_n13975), .Y(new_n13984));
  xor_4  g11636(.A(new_n13984), .B(pi207), .Y(new_n13985));
  xor_4  g11637(.A(new_n13968), .B(new_n13947), .Y(new_n13986));
  not_8  g11638(.A(new_n13986), .Y(new_n13987));
  not_8  g11639(.A(new_n12939), .Y(new_n13988));
  xor_4  g11640(.A(new_n13961), .B(new_n13959), .Y(new_n13989));
  xor_4  g11641(.A(new_n13955), .B(pi254), .Y(new_n13990));
  not_8  g11642(.A(new_n13990), .Y(new_n13991));
  nand_5 g11643(.A(new_n13279), .B(new_n13269), .Y(new_n13992));
  or_6   g11644(.A(new_n13280), .B(new_n12954), .Y(new_n13993));
  nand_5 g11645(.A(new_n13993), .B(new_n13992), .Y(new_n13994));
  nand_5 g11646(.A(new_n13994), .B(new_n13991), .Y(new_n13995));
  xor_4  g11647(.A(new_n13994), .B(new_n13990), .Y(new_n13996));
  or_6   g11648(.A(new_n13996), .B(new_n12948), .Y(new_n13997));
  nand_5 g11649(.A(new_n13997), .B(new_n13995), .Y(new_n13998));
  nand_5 g11650(.A(new_n13998), .B(new_n13989), .Y(new_n13999));
  xnor_4 g11651(.A(new_n13998), .B(new_n13989), .Y(new_n14000));
  or_6   g11652(.A(new_n14000), .B(new_n12944), .Y(new_n14001));
  nand_5 g11653(.A(new_n14001), .B(new_n13999), .Y(new_n14002));
  nand_5 g11654(.A(new_n14002), .B(new_n13988), .Y(new_n14003));
  nor_5  g11655(.A(new_n14002), .B(new_n13988), .Y(new_n14004));
  nor_5  g11656(.A(new_n13966), .B(new_n13965), .Y(new_n14005));
  xor_4  g11657(.A(new_n14005), .B(pi383), .Y(new_n14006));
  or_6   g11658(.A(new_n14006), .B(new_n14004), .Y(new_n14007));
  nand_5 g11659(.A(new_n14007), .B(new_n14003), .Y(new_n14008));
  nand_5 g11660(.A(new_n14008), .B(new_n13987), .Y(new_n14009));
  xor_4  g11661(.A(new_n14008), .B(new_n13986), .Y(new_n14010));
  or_6   g11662(.A(new_n14010), .B(new_n12931), .Y(new_n14011));
  nand_5 g11663(.A(new_n14011), .B(new_n14009), .Y(new_n14012));
  nand_5 g11664(.A(new_n13973), .B(new_n13971), .Y(new_n14013));
  xor_4  g11665(.A(new_n14013), .B(pi136), .Y(new_n14014));
  nand_5 g11666(.A(new_n14014), .B(new_n14012), .Y(new_n14015));
  xnor_4 g11667(.A(new_n14014), .B(new_n14012), .Y(new_n14016));
  or_6   g11668(.A(new_n14016), .B(new_n13004), .Y(new_n14017));
  nand_5 g11669(.A(new_n14017), .B(new_n14015), .Y(new_n14018));
  nand_5 g11670(.A(new_n14018), .B(new_n13985), .Y(new_n14019));
  or_6   g11671(.A(new_n14018), .B(new_n13985), .Y(new_n14020));
  nand_5 g11672(.A(new_n14020), .B(new_n12926), .Y(new_n14021));
  nand_5 g11673(.A(new_n14021), .B(new_n14019), .Y(new_n14022));
  nand_5 g11674(.A(new_n14022), .B(new_n13983), .Y(new_n14023));
  not_8  g11675(.A(new_n14023), .Y(new_n14024));
  nor_5  g11676(.A(new_n14024), .B(new_n13982), .Y(new_n14025));
  xor_4  g11677(.A(new_n13979), .B(new_n13045), .Y(new_n14026));
  nor_5  g11678(.A(new_n14026), .B(new_n14025), .Y(new_n14027));
  nor_5  g11679(.A(new_n14027), .B(new_n13980), .Y(po0125));
  xnor_4 g11680(.A(new_n11244), .B(new_n11243), .Y(po0126));
  xor_4  g11681(.A(new_n13749), .B(new_n7338), .Y(new_n14030));
  or_6   g11682(.A(new_n13753), .B(new_n7341), .Y(new_n14031));
  xor_4  g11683(.A(new_n13753), .B(new_n7341), .Y(new_n14032));
  nand_5 g11684(.A(new_n13744), .B(new_n7344), .Y(new_n14033));
  nand_5 g11685(.A(new_n13755), .B(new_n7345), .Y(new_n14034));
  nand_5 g11686(.A(new_n14034), .B(new_n14033), .Y(new_n14035));
  xor_4  g11687(.A(new_n14035), .B(new_n13756), .Y(new_n14036));
  nand_5 g11688(.A(new_n14036), .B(new_n7349), .Y(new_n14037));
  nand_5 g11689(.A(new_n13763), .B(new_n7345), .Y(new_n14038));
  or_6   g11690(.A(new_n14038), .B(new_n14036), .Y(new_n14039));
  nand_5 g11691(.A(new_n14039), .B(new_n14037), .Y(new_n14040));
  nand_5 g11692(.A(new_n14040), .B(new_n14032), .Y(new_n14041));
  nand_5 g11693(.A(new_n14041), .B(new_n14031), .Y(new_n14042));
  xnor_4 g11694(.A(new_n14042), .B(new_n14030), .Y(new_n14043));
  nand_5 g11695(.A(pi576), .B(new_n5246), .Y(new_n14044));
  xor_4  g11696(.A(pi576), .B(new_n5246), .Y(new_n14045));
  nand_5 g11697(.A(pi401), .B(new_n2872), .Y(new_n14046));
  xor_4  g11698(.A(pi401), .B(new_n2872), .Y(new_n14047));
  nand_5 g11699(.A(new_n14047), .B(new_n12256), .Y(new_n14048));
  nand_5 g11700(.A(new_n14048), .B(new_n14046), .Y(new_n14049));
  nand_5 g11701(.A(new_n14049), .B(new_n14045), .Y(new_n14050));
  nand_5 g11702(.A(new_n14050), .B(new_n14044), .Y(new_n14051));
  xor_4  g11703(.A(pi273), .B(new_n2883), .Y(new_n14052));
  xor_4  g11704(.A(new_n14052), .B(new_n14051), .Y(new_n14053));
  xor_4  g11705(.A(new_n14053), .B(new_n14043), .Y(new_n14054));
  xor_4  g11706(.A(new_n14040), .B(new_n14032), .Y(new_n14055));
  not_8  g11707(.A(new_n14055), .Y(new_n14056));
  xor_4  g11708(.A(new_n14049), .B(new_n14045), .Y(new_n14057));
  and_6  g11709(.A(new_n14057), .B(new_n14056), .Y(new_n14058));
  nor_5  g11710(.A(new_n14057), .B(new_n14056), .Y(new_n14059));
  xor_4  g11711(.A(new_n13798), .B(new_n7344), .Y(new_n14060));
  not_8  g11712(.A(new_n14060), .Y(new_n14061));
  xor_4  g11713(.A(new_n14036), .B(new_n7348), .Y(new_n14062));
  and_6  g11714(.A(new_n14062), .B(new_n14061), .Y(new_n14063));
  or_6   g11715(.A(new_n14063), .B(new_n14048), .Y(new_n14064));
  nand_5 g11716(.A(new_n14060), .B(new_n12254), .Y(new_n14065));
  nor_5  g11717(.A(new_n14065), .B(new_n14047), .Y(new_n14066));
  nand_5 g11718(.A(new_n14061), .B(new_n12256), .Y(new_n14067));
  nand_5 g11719(.A(new_n14067), .B(new_n14065), .Y(new_n14068));
  xor_4  g11720(.A(new_n14068), .B(new_n14047), .Y(new_n14069));
  nor_5  g11721(.A(new_n14069), .B(new_n14062), .Y(new_n14070));
  nor_5  g11722(.A(new_n14070), .B(new_n14066), .Y(new_n14071));
  nand_5 g11723(.A(new_n14071), .B(new_n14064), .Y(new_n14072));
  nor_5  g11724(.A(new_n14072), .B(new_n14059), .Y(new_n14073));
  nor_5  g11725(.A(new_n14073), .B(new_n14058), .Y(new_n14074));
  xor_4  g11726(.A(new_n14074), .B(new_n14054), .Y(po0127));
  xor_4  g11727(.A(new_n13094), .B(new_n6015), .Y(po0128));
  xor_4  g11728(.A(pi419), .B(new_n6353), .Y(new_n14077));
  not_8  g11729(.A(pi554), .Y(new_n14078));
  nand_5 g11730(.A(new_n14078), .B(pi054), .Y(new_n14079));
  not_8  g11731(.A(pi647), .Y(new_n14080));
  nand_5 g11732(.A(new_n14080), .B(pi418), .Y(new_n14081));
  xor_4  g11733(.A(pi647), .B(new_n6236), .Y(new_n14082));
  nand_5 g11734(.A(pi791), .B(new_n4060), .Y(new_n14083));
  xor_4  g11735(.A(pi791), .B(new_n4060), .Y(new_n14084));
  nand_5 g11736(.A(new_n3999), .B(pi479), .Y(new_n14085));
  nand_5 g11737(.A(new_n3962), .B(pi058), .Y(new_n14086));
  not_8  g11738(.A(new_n12333), .Y(new_n14087));
  nand_5 g11739(.A(new_n14087), .B(new_n12328), .Y(new_n14088));
  nand_5 g11740(.A(new_n14088), .B(new_n14086), .Y(new_n14089));
  xor_4  g11741(.A(pi602), .B(new_n6241), .Y(new_n14090));
  nand_5 g11742(.A(new_n14090), .B(new_n14089), .Y(new_n14091));
  nand_5 g11743(.A(new_n14091), .B(new_n14085), .Y(new_n14092));
  nand_5 g11744(.A(new_n14092), .B(new_n14084), .Y(new_n14093));
  nand_5 g11745(.A(new_n14093), .B(new_n14083), .Y(new_n14094));
  nand_5 g11746(.A(new_n14094), .B(new_n14082), .Y(new_n14095));
  nand_5 g11747(.A(new_n14095), .B(new_n14081), .Y(new_n14096));
  xor_4  g11748(.A(pi554), .B(pi054), .Y(new_n14097));
  not_8  g11749(.A(new_n14097), .Y(new_n14098));
  nand_5 g11750(.A(new_n14098), .B(new_n14096), .Y(new_n14099));
  nand_5 g11751(.A(new_n14099), .B(new_n14079), .Y(new_n14100));
  xor_4  g11752(.A(new_n14100), .B(new_n14077), .Y(new_n14101));
  not_8  g11753(.A(new_n14101), .Y(new_n14102));
  xor_4  g11754(.A(new_n14097), .B(new_n14096), .Y(new_n14103));
  or_6   g11755(.A(new_n6560), .B(new_n6553), .Y(new_n14104));
  nand_5 g11756(.A(new_n6564), .B(new_n6561), .Y(new_n14105));
  nand_5 g11757(.A(new_n14105), .B(new_n14104), .Y(new_n14106));
  xor_4  g11758(.A(pi119), .B(new_n12563), .Y(new_n14107));
  nor_5  g11759(.A(pi517), .B(new_n6554), .Y(new_n14108));
  not_8  g11760(.A(new_n6555), .Y(new_n14109));
  nor_5  g11761(.A(new_n6559), .B(new_n14109), .Y(new_n14110));
  nor_5  g11762(.A(new_n14110), .B(new_n14108), .Y(new_n14111));
  xnor_4 g11763(.A(new_n14111), .B(new_n14107), .Y(new_n14112));
  nand_5 g11764(.A(new_n14112), .B(new_n11455), .Y(new_n14113));
  or_6   g11765(.A(new_n14112), .B(new_n11455), .Y(new_n14114));
  nand_5 g11766(.A(new_n14114), .B(new_n14113), .Y(new_n14115));
  xor_4  g11767(.A(new_n14115), .B(new_n14106), .Y(new_n14116));
  not_8  g11768(.A(new_n14116), .Y(new_n14117));
  nand_5 g11769(.A(new_n14117), .B(new_n14103), .Y(new_n14118));
  xor_4  g11770(.A(new_n14094), .B(new_n14082), .Y(new_n14119));
  xor_4  g11771(.A(new_n14092), .B(new_n14084), .Y(new_n14120));
  xor_4  g11772(.A(new_n14090), .B(new_n14089), .Y(new_n14121));
  nor_5  g11773(.A(new_n14121), .B(new_n6509), .Y(new_n14122));
  not_8  g11774(.A(new_n12334), .Y(new_n14123));
  nor_5  g11775(.A(new_n14123), .B(new_n12327), .Y(new_n14124));
  nor_5  g11776(.A(new_n12335), .B(new_n6510), .Y(new_n14125));
  nor_5  g11777(.A(new_n14125), .B(new_n14124), .Y(new_n14126));
  xor_4  g11778(.A(new_n14121), .B(new_n6508), .Y(new_n14127));
  or_6   g11779(.A(new_n14127), .B(new_n14126), .Y(new_n14128));
  not_8  g11780(.A(new_n14128), .Y(new_n14129));
  nor_5  g11781(.A(new_n14129), .B(new_n14122), .Y(new_n14130));
  or_6   g11782(.A(new_n14130), .B(new_n14120), .Y(new_n14131));
  not_8  g11783(.A(new_n14131), .Y(new_n14132));
  xnor_4 g11784(.A(new_n14130), .B(new_n14120), .Y(new_n14133));
  nor_5  g11785(.A(new_n14133), .B(new_n6536), .Y(new_n14134));
  nor_5  g11786(.A(new_n14134), .B(new_n14132), .Y(new_n14135));
  or_6   g11787(.A(new_n14135), .B(new_n14119), .Y(new_n14136));
  xnor_4 g11788(.A(new_n14135), .B(new_n14119), .Y(new_n14137));
  not_8  g11789(.A(new_n14137), .Y(new_n14138));
  nand_5 g11790(.A(new_n14138), .B(new_n6565), .Y(new_n14139));
  nand_5 g11791(.A(new_n14139), .B(new_n14136), .Y(new_n14140));
  xor_4  g11792(.A(new_n14116), .B(new_n14103), .Y(new_n14141));
  not_8  g11793(.A(new_n14141), .Y(new_n14142));
  nand_5 g11794(.A(new_n14142), .B(new_n14140), .Y(new_n14143));
  nand_5 g11795(.A(new_n14143), .B(new_n14118), .Y(new_n14144));
  nand_5 g11796(.A(new_n14144), .B(new_n14102), .Y(new_n14145));
  not_8  g11797(.A(new_n14145), .Y(new_n14146));
  xor_4  g11798(.A(pi198), .B(new_n12535), .Y(new_n14147));
  nand_5 g11799(.A(pi119), .B(new_n12563), .Y(new_n14148));
  nand_5 g11800(.A(new_n14111), .B(new_n14107), .Y(new_n14149));
  nand_5 g11801(.A(new_n14149), .B(new_n14148), .Y(new_n14150));
  xor_4  g11802(.A(new_n14150), .B(new_n14147), .Y(new_n14151));
  xor_4  g11803(.A(new_n14151), .B(new_n11451), .Y(new_n14152));
  nand_5 g11804(.A(new_n14114), .B(new_n14106), .Y(new_n14153));
  nand_5 g11805(.A(new_n14153), .B(new_n14113), .Y(new_n14154));
  xor_4  g11806(.A(new_n14154), .B(new_n14152), .Y(new_n14155));
  not_8  g11807(.A(new_n14155), .Y(new_n14156));
  xor_4  g11808(.A(new_n14144), .B(new_n14101), .Y(new_n14157));
  nor_5  g11809(.A(new_n14157), .B(new_n14156), .Y(new_n14158));
  nor_5  g11810(.A(new_n14158), .B(new_n14146), .Y(new_n14159));
  not_8  g11811(.A(new_n11447), .Y(new_n14160));
  xor_4  g11812(.A(pi327), .B(new_n12597), .Y(new_n14161));
  nand_5 g11813(.A(new_n12560), .B(pi070), .Y(new_n14162));
  nand_5 g11814(.A(new_n14150), .B(new_n14147), .Y(new_n14163));
  nand_5 g11815(.A(new_n14163), .B(new_n14162), .Y(new_n14164));
  xnor_4 g11816(.A(new_n14164), .B(new_n14161), .Y(new_n14165));
  xor_4  g11817(.A(new_n14165), .B(new_n14160), .Y(new_n14166));
  nor_5  g11818(.A(new_n14151), .B(new_n11451), .Y(new_n14167));
  and_6  g11819(.A(new_n14154), .B(new_n14152), .Y(new_n14168));
  nor_5  g11820(.A(new_n14168), .B(new_n14167), .Y(new_n14169));
  xor_4  g11821(.A(new_n14169), .B(new_n14166), .Y(new_n14170));
  or_6   g11822(.A(new_n14170), .B(new_n14159), .Y(new_n14171));
  not_8  g11823(.A(new_n14171), .Y(new_n14172));
  xor_4  g11824(.A(pi110), .B(new_n6372), .Y(new_n14173));
  not_8  g11825(.A(pi419), .Y(new_n14174));
  nand_5 g11826(.A(new_n14174), .B(pi032), .Y(new_n14175));
  nand_5 g11827(.A(new_n14100), .B(new_n14077), .Y(new_n14176));
  nand_5 g11828(.A(new_n14176), .B(new_n14175), .Y(new_n14177));
  xor_4  g11829(.A(new_n14177), .B(new_n14173), .Y(new_n14178));
  not_8  g11830(.A(new_n14170), .Y(new_n14179));
  xor_4  g11831(.A(new_n14179), .B(new_n14159), .Y(new_n14180));
  nor_5  g11832(.A(new_n14180), .B(new_n14178), .Y(new_n14181));
  nor_5  g11833(.A(new_n14181), .B(new_n14172), .Y(new_n14182));
  nand_5 g11834(.A(pi110), .B(new_n6372), .Y(new_n14183));
  nand_5 g11835(.A(new_n14177), .B(new_n14173), .Y(new_n14184));
  nand_5 g11836(.A(new_n14184), .B(new_n14183), .Y(new_n14185));
  nand_5 g11837(.A(new_n14185), .B(new_n14182), .Y(new_n14186));
  nor_5  g11838(.A(new_n14185), .B(new_n14182), .Y(new_n14187));
  not_8  g11839(.A(new_n14187), .Y(new_n14188));
  or_6   g11840(.A(new_n14165), .B(new_n14160), .Y(new_n14189));
  nand_5 g11841(.A(new_n14169), .B(new_n14166), .Y(new_n14190));
  nand_5 g11842(.A(new_n14190), .B(new_n14189), .Y(new_n14191));
  nand_5 g11843(.A(new_n14191), .B(new_n14188), .Y(new_n14192));
  nand_5 g11844(.A(new_n14192), .B(new_n14186), .Y(new_n14193));
  nand_5 g11845(.A(pi327), .B(new_n12597), .Y(new_n14194));
  nand_5 g11846(.A(new_n14164), .B(new_n14161), .Y(new_n14195));
  nand_5 g11847(.A(new_n14195), .B(new_n14194), .Y(new_n14196));
  nand_5 g11848(.A(pi593), .B(new_n11433), .Y(new_n14197));
  nand_5 g11849(.A(new_n11446), .B(new_n11434), .Y(new_n14198));
  nand_5 g11850(.A(new_n14198), .B(new_n14197), .Y(new_n14199));
  not_8  g11851(.A(new_n14199), .Y(new_n14200));
  nand_5 g11852(.A(new_n14200), .B(new_n14196), .Y(new_n14201));
  not_8  g11853(.A(new_n14201), .Y(new_n14202));
  nand_5 g11854(.A(new_n14188), .B(new_n14186), .Y(new_n14203));
  not_8  g11855(.A(new_n14203), .Y(new_n14204));
  nor_5  g11856(.A(new_n14200), .B(new_n14196), .Y(new_n14205));
  not_8  g11857(.A(new_n14205), .Y(new_n14206));
  nand_5 g11858(.A(new_n14206), .B(new_n14201), .Y(new_n14207));
  nor_5  g11859(.A(new_n14207), .B(new_n14192), .Y(new_n14208));
  not_8  g11860(.A(new_n14191), .Y(new_n14209));
  nand_5 g11861(.A(new_n14209), .B(new_n14187), .Y(new_n14210));
  and_6  g11862(.A(new_n14202), .B(new_n14192), .Y(new_n14211));
  and_6  g11863(.A(new_n14211), .B(new_n14210), .Y(new_n14212));
  nor_5  g11864(.A(new_n14212), .B(new_n14208), .Y(new_n14213));
  nor_5  g11865(.A(new_n14213), .B(new_n14204), .Y(po1243));
  or_6   g11866(.A(po1243), .B(new_n14202), .Y(new_n14215));
  nand_5 g11867(.A(new_n14215), .B(new_n14193), .Y(new_n14216));
  nor_5  g11868(.A(new_n14210), .B(new_n14202), .Y(new_n14217));
  nor_5  g11869(.A(new_n14206), .B(new_n14193), .Y(new_n14218));
  nor_5  g11870(.A(new_n14218), .B(new_n14217), .Y(new_n14219));
  nand_5 g11871(.A(new_n14219), .B(new_n14216), .Y(po0129));
  xor_4  g11872(.A(pi090), .B(new_n9261), .Y(new_n14221));
  nand_5 g11873(.A(new_n9232), .B(pi235), .Y(new_n14222));
  xor_4  g11874(.A(pi480), .B(new_n10838), .Y(new_n14223));
  nand_5 g11875(.A(pi828), .B(new_n9235), .Y(new_n14224));
  not_8  g11876(.A(new_n14224), .Y(new_n14225));
  nand_5 g11877(.A(new_n14225), .B(new_n14223), .Y(new_n14226));
  nand_5 g11878(.A(new_n14226), .B(new_n14222), .Y(new_n14227));
  xor_4  g11879(.A(new_n14227), .B(new_n14221), .Y(new_n14228));
  not_8  g11880(.A(new_n14228), .Y(new_n14229));
  nor_5  g11881(.A(new_n14223), .B(new_n9031), .Y(new_n14230));
  nand_5 g11882(.A(new_n14225), .B(new_n9022), .Y(new_n14231));
  nand_5 g11883(.A(new_n14231), .B(new_n14230), .Y(new_n14232));
  nor_5  g11884(.A(pi828), .B(new_n9235), .Y(new_n14233));
  nand_5 g11885(.A(new_n14233), .B(new_n9021), .Y(new_n14234));
  nand_5 g11886(.A(new_n14234), .B(new_n14232), .Y(new_n14235));
  nand_5 g11887(.A(new_n14223), .B(new_n9031), .Y(new_n14236));
  nand_5 g11888(.A(new_n14236), .B(new_n14235), .Y(new_n14237));
  or_6   g11889(.A(new_n14226), .B(new_n9033), .Y(new_n14238));
  nand_5 g11890(.A(new_n14238), .B(new_n14237), .Y(new_n14239));
  nor_5  g11891(.A(new_n14239), .B(new_n14229), .Y(new_n14240));
  xor_4  g11892(.A(new_n14239), .B(new_n14228), .Y(new_n14241));
  nor_5  g11893(.A(new_n14241), .B(new_n9116), .Y(new_n14242));
  or_6   g11894(.A(new_n14242), .B(new_n14240), .Y(new_n14243));
  nand_5 g11895(.A(new_n9229), .B(pi048), .Y(new_n14244));
  nand_5 g11896(.A(new_n14227), .B(new_n14221), .Y(new_n14245));
  nand_5 g11897(.A(new_n14245), .B(new_n14244), .Y(new_n14246));
  xor_4  g11898(.A(pi343), .B(pi087), .Y(new_n14247));
  xor_4  g11899(.A(new_n14247), .B(new_n14246), .Y(new_n14248));
  xor_4  g11900(.A(new_n14248), .B(new_n14243), .Y(new_n14249));
  not_8  g11901(.A(new_n14249), .Y(new_n14250));
  xor_4  g11902(.A(new_n14250), .B(new_n9123), .Y(po0130));
  not_8  g11903(.A(pi769), .Y(new_n14252));
  nand_5 g11904(.A(new_n14252), .B(new_n6091), .Y(new_n14253));
  not_8  g11905(.A(new_n14253), .Y(new_n14254));
  xor_4  g11906(.A(pi769), .B(pi280), .Y(new_n14255));
  not_8  g11907(.A(new_n14255), .Y(new_n14256));
  nand_5 g11908(.A(pi275), .B(pi092), .Y(new_n14257));
  not_8  g11909(.A(pi275), .Y(new_n14258));
  nand_5 g11910(.A(new_n14258), .B(new_n7255), .Y(new_n14259));
  nand_5 g11911(.A(pi621), .B(pi459), .Y(new_n14260));
  not_8  g11912(.A(pi459), .Y(new_n14261));
  nand_5 g11913(.A(new_n6077), .B(new_n14261), .Y(new_n14262));
  nand_5 g11914(.A(new_n9555), .B(new_n9551), .Y(new_n14263));
  nand_5 g11915(.A(new_n14263), .B(new_n9553), .Y(new_n14264));
  nand_5 g11916(.A(new_n14264), .B(new_n14262), .Y(new_n14265));
  nand_5 g11917(.A(new_n14265), .B(new_n14260), .Y(new_n14266));
  nand_5 g11918(.A(new_n14266), .B(new_n14259), .Y(new_n14267));
  nand_5 g11919(.A(new_n14267), .B(new_n14257), .Y(new_n14268));
  nor_5  g11920(.A(new_n14268), .B(new_n14256), .Y(new_n14269));
  nor_5  g11921(.A(new_n14269), .B(new_n14254), .Y(new_n14270));
  not_8  g11922(.A(new_n14270), .Y(new_n14271));
  xor_4  g11923(.A(new_n14268), .B(new_n14255), .Y(new_n14272));
  not_8  g11924(.A(new_n14272), .Y(new_n14273));
  nand_5 g11925(.A(new_n14273), .B(new_n11091), .Y(new_n14274));
  xor_4  g11926(.A(new_n14272), .B(pi534), .Y(new_n14275));
  nand_5 g11927(.A(new_n14257), .B(new_n14259), .Y(new_n14276));
  xor_4  g11928(.A(new_n14276), .B(new_n14266), .Y(new_n14277));
  nand_5 g11929(.A(new_n14277), .B(new_n7257), .Y(new_n14278));
  not_8  g11930(.A(new_n14277), .Y(new_n14279));
  nand_5 g11931(.A(new_n14279), .B(pi028), .Y(new_n14280));
  nand_5 g11932(.A(new_n14260), .B(new_n14262), .Y(new_n14281));
  xor_4  g11933(.A(new_n14281), .B(new_n14264), .Y(new_n14282));
  nand_5 g11934(.A(new_n14282), .B(new_n11096), .Y(new_n14283));
  xor_4  g11935(.A(new_n14282), .B(new_n11096), .Y(new_n14284));
  nand_5 g11936(.A(new_n9558), .B(new_n10647), .Y(new_n14285));
  nand_5 g11937(.A(new_n9557), .B(pi332), .Y(new_n14286));
  nand_5 g11938(.A(new_n9516), .B(new_n11101), .Y(new_n14287));
  xor_4  g11939(.A(new_n9515), .B(pi265), .Y(new_n14288));
  or_6   g11940(.A(new_n9480), .B(pi635), .Y(new_n14289));
  or_6   g11941(.A(new_n9389), .B(pi545), .Y(new_n14290));
  xor_4  g11942(.A(new_n9389), .B(pi545), .Y(new_n14291));
  nand_5 g11943(.A(new_n9403), .B(new_n6575), .Y(new_n14292));
  xor_4  g11944(.A(new_n9403), .B(new_n6575), .Y(new_n14293));
  not_8  g11945(.A(new_n14293), .Y(new_n14294));
  nand_5 g11946(.A(new_n9395), .B(pi281), .Y(new_n14295));
  nand_5 g11947(.A(new_n14295), .B(new_n9382), .Y(new_n14296));
  xor_4  g11948(.A(new_n7276), .B(new_n5768), .Y(new_n14297));
  nor_5  g11949(.A(new_n14297), .B(new_n14296), .Y(new_n14298));
  and_6  g11950(.A(new_n14297), .B(new_n14296), .Y(new_n14299));
  nor_5  g11951(.A(new_n14299), .B(new_n8511), .Y(new_n14300));
  nor_5  g11952(.A(new_n14300), .B(new_n9384), .Y(new_n14301));
  nor_5  g11953(.A(new_n14301), .B(new_n14298), .Y(new_n14302));
  or_6   g11954(.A(new_n14302), .B(new_n14294), .Y(new_n14303));
  nand_5 g11955(.A(new_n14303), .B(new_n14292), .Y(new_n14304));
  nand_5 g11956(.A(new_n14304), .B(new_n14291), .Y(new_n14305));
  nand_5 g11957(.A(new_n14305), .B(new_n14290), .Y(new_n14306));
  xor_4  g11958(.A(new_n9480), .B(pi635), .Y(new_n14307));
  nand_5 g11959(.A(new_n14307), .B(new_n14306), .Y(new_n14308));
  nand_5 g11960(.A(new_n14308), .B(new_n14289), .Y(new_n14309));
  nand_5 g11961(.A(new_n14309), .B(new_n14288), .Y(new_n14310));
  nand_5 g11962(.A(new_n14310), .B(new_n14287), .Y(new_n14311));
  nand_5 g11963(.A(new_n14311), .B(new_n14286), .Y(new_n14312));
  nand_5 g11964(.A(new_n14312), .B(new_n14285), .Y(new_n14313));
  nand_5 g11965(.A(new_n14313), .B(new_n14284), .Y(new_n14314));
  nand_5 g11966(.A(new_n14314), .B(new_n14283), .Y(new_n14315));
  nand_5 g11967(.A(new_n14315), .B(new_n14280), .Y(new_n14316));
  nand_5 g11968(.A(new_n14316), .B(new_n14278), .Y(new_n14317));
  nand_5 g11969(.A(new_n14317), .B(new_n14275), .Y(new_n14318));
  nand_5 g11970(.A(new_n14318), .B(new_n14274), .Y(new_n14319));
  nor_5  g11971(.A(new_n14319), .B(new_n14271), .Y(new_n14320));
  not_8  g11972(.A(new_n14320), .Y(new_n14321));
  xor_4  g11973(.A(new_n14317), .B(new_n14275), .Y(new_n14322));
  not_8  g11974(.A(new_n14322), .Y(new_n14323));
  nand_5 g11975(.A(new_n4136), .B(new_n3726), .Y(new_n14324));
  not_8  g11976(.A(new_n14324), .Y(new_n14325));
  nand_5 g11977(.A(new_n14325), .B(new_n3723), .Y(new_n14326));
  nor_5  g11978(.A(new_n14326), .B(pi795), .Y(new_n14327));
  nand_5 g11979(.A(new_n14327), .B(new_n3718), .Y(new_n14328));
  nor_5  g11980(.A(new_n14328), .B(pi641), .Y(new_n14329));
  nand_5 g11981(.A(new_n14329), .B(new_n3710), .Y(new_n14330));
  nor_5  g11982(.A(new_n14330), .B(pi021), .Y(new_n14331));
  nand_5 g11983(.A(new_n14331), .B(new_n7483), .Y(new_n14332));
  xor_4  g11984(.A(new_n14332), .B(new_n7494), .Y(new_n14333));
  xor_4  g11985(.A(new_n14333), .B(new_n4864), .Y(new_n14334));
  xor_4  g11986(.A(new_n14331), .B(new_n7483), .Y(new_n14335));
  nor_5  g11987(.A(new_n14335), .B(new_n4848), .Y(new_n14336));
  xor_4  g11988(.A(new_n14329), .B(new_n3710), .Y(new_n14337));
  nand_5 g11989(.A(new_n14337), .B(new_n4829), .Y(new_n14338));
  xor_4  g11990(.A(new_n14337), .B(new_n4829), .Y(new_n14339));
  xor_4  g11991(.A(new_n14328), .B(pi641), .Y(new_n14340));
  nand_5 g11992(.A(new_n14340), .B(new_n4793), .Y(new_n14341));
  or_6   g11993(.A(new_n14340), .B(new_n4793), .Y(new_n14342));
  xor_4  g11994(.A(new_n14324), .B(pi495), .Y(new_n14343));
  not_8  g11995(.A(new_n14343), .Y(new_n14344));
  nand_5 g11996(.A(new_n4801), .B(new_n4797), .Y(new_n14345));
  nand_5 g11997(.A(new_n14345), .B(new_n14325), .Y(new_n14346));
  nand_5 g11998(.A(new_n4797), .B(new_n4136), .Y(new_n14347));
  nand_5 g11999(.A(new_n14347), .B(pi422), .Y(new_n14348));
  or_6   g12000(.A(new_n14348), .B(new_n4801), .Y(new_n14349));
  nand_5 g12001(.A(new_n14349), .B(new_n14346), .Y(new_n14350));
  nor_5  g12002(.A(new_n14350), .B(new_n14344), .Y(new_n14351));
  xor_4  g12003(.A(new_n14350), .B(new_n14344), .Y(new_n14352));
  not_8  g12004(.A(new_n14352), .Y(new_n14353));
  nor_5  g12005(.A(new_n14353), .B(new_n4805), .Y(new_n14354));
  nor_5  g12006(.A(new_n14354), .B(new_n14351), .Y(new_n14355));
  xor_4  g12007(.A(new_n14326), .B(new_n4227), .Y(new_n14356));
  nand_5 g12008(.A(new_n14356), .B(new_n14355), .Y(new_n14357));
  xnor_4 g12009(.A(new_n14356), .B(new_n14355), .Y(new_n14358));
  or_6   g12010(.A(new_n14358), .B(new_n4812), .Y(new_n14359));
  nand_5 g12011(.A(new_n14359), .B(new_n14357), .Y(new_n14360));
  nor_5  g12012(.A(new_n14360), .B(new_n13174), .Y(new_n14361));
  xor_4  g12013(.A(new_n14360), .B(new_n13174), .Y(new_n14362));
  not_8  g12014(.A(new_n14362), .Y(new_n14363));
  xor_4  g12015(.A(new_n14327), .B(pi201), .Y(new_n14364));
  nor_5  g12016(.A(new_n14364), .B(new_n14363), .Y(new_n14365));
  or_6   g12017(.A(new_n14365), .B(new_n14361), .Y(new_n14366));
  nand_5 g12018(.A(new_n14366), .B(new_n14342), .Y(new_n14367));
  nand_5 g12019(.A(new_n14367), .B(new_n14341), .Y(new_n14368));
  nand_5 g12020(.A(new_n14368), .B(new_n14339), .Y(new_n14369));
  nand_5 g12021(.A(new_n14369), .B(new_n14338), .Y(new_n14370));
  nor_5  g12022(.A(new_n14370), .B(new_n4790), .Y(new_n14371));
  xor_4  g12023(.A(new_n14330), .B(pi021), .Y(new_n14372));
  xor_4  g12024(.A(new_n14370), .B(new_n4790), .Y(new_n14373));
  not_8  g12025(.A(new_n14373), .Y(new_n14374));
  nor_5  g12026(.A(new_n14374), .B(new_n14372), .Y(new_n14375));
  or_6   g12027(.A(new_n14375), .B(new_n14371), .Y(new_n14376));
  xor_4  g12028(.A(new_n14335), .B(new_n4848), .Y(new_n14377));
  nand_5 g12029(.A(new_n14377), .B(new_n14376), .Y(new_n14378));
  not_8  g12030(.A(new_n14378), .Y(new_n14379));
  nor_5  g12031(.A(new_n14379), .B(new_n14336), .Y(new_n14380));
  xor_4  g12032(.A(new_n14380), .B(new_n14334), .Y(new_n14381));
  nor_5  g12033(.A(new_n14381), .B(new_n14323), .Y(new_n14382));
  nand_5 g12034(.A(new_n14278), .B(new_n14280), .Y(new_n14383));
  xnor_4 g12035(.A(new_n14383), .B(new_n14315), .Y(new_n14384));
  xor_4  g12036(.A(new_n14377), .B(new_n14376), .Y(new_n14385));
  nor_5  g12037(.A(new_n14385), .B(new_n14384), .Y(new_n14386));
  xor_4  g12038(.A(new_n14385), .B(new_n14384), .Y(new_n14387));
  not_8  g12039(.A(new_n14387), .Y(new_n14388));
  xor_4  g12040(.A(new_n14313), .B(new_n14284), .Y(new_n14389));
  not_8  g12041(.A(new_n14389), .Y(new_n14390));
  xor_4  g12042(.A(new_n14373), .B(new_n14372), .Y(new_n14391));
  nor_5  g12043(.A(new_n14391), .B(new_n14390), .Y(new_n14392));
  and_6  g12044(.A(new_n14286), .B(new_n14285), .Y(new_n14393));
  xor_4  g12045(.A(new_n14393), .B(new_n14311), .Y(new_n14394));
  not_8  g12046(.A(new_n14394), .Y(new_n14395));
  xor_4  g12047(.A(new_n14368), .B(new_n14339), .Y(new_n14396));
  nor_5  g12048(.A(new_n14396), .B(new_n14395), .Y(new_n14397));
  xor_4  g12049(.A(new_n14396), .B(new_n14394), .Y(new_n14398));
  xor_4  g12050(.A(new_n14309), .B(new_n14288), .Y(new_n14399));
  nand_5 g12051(.A(new_n14342), .B(new_n14341), .Y(new_n14400));
  xor_4  g12052(.A(new_n14400), .B(new_n14366), .Y(new_n14401));
  or_6   g12053(.A(new_n14401), .B(new_n14399), .Y(new_n14402));
  xor_4  g12054(.A(new_n14307), .B(new_n14306), .Y(new_n14403));
  xor_4  g12055(.A(new_n14364), .B(new_n14362), .Y(new_n14404));
  nor_5  g12056(.A(new_n14404), .B(new_n14403), .Y(new_n14405));
  xor_4  g12057(.A(new_n14404), .B(new_n14403), .Y(new_n14406));
  not_8  g12058(.A(new_n14406), .Y(new_n14407));
  xor_4  g12059(.A(new_n14304), .B(new_n14291), .Y(new_n14408));
  not_8  g12060(.A(new_n14408), .Y(new_n14409));
  xor_4  g12061(.A(new_n14358), .B(new_n4813), .Y(new_n14410));
  nand_5 g12062(.A(new_n14410), .B(new_n14409), .Y(new_n14411));
  not_8  g12063(.A(new_n14411), .Y(new_n14412));
  xor_4  g12064(.A(new_n14410), .B(new_n14408), .Y(new_n14413));
  xor_4  g12065(.A(new_n14302), .B(new_n14294), .Y(new_n14414));
  xor_4  g12066(.A(new_n14352), .B(new_n4805), .Y(new_n14415));
  nand_5 g12067(.A(new_n14415), .B(new_n14414), .Y(new_n14416));
  not_8  g12068(.A(new_n14414), .Y(new_n14417));
  xor_4  g12069(.A(new_n14415), .B(new_n14417), .Y(new_n14418));
  nor_5  g12070(.A(new_n14299), .B(new_n14298), .Y(new_n14419));
  xor_4  g12071(.A(new_n9395), .B(pi281), .Y(new_n14420));
  xor_4  g12072(.A(new_n4796), .B(pi781), .Y(new_n14421));
  nand_5 g12073(.A(new_n14421), .B(new_n14420), .Y(new_n14422));
  not_8  g12074(.A(new_n14422), .Y(new_n14423));
  not_8  g12075(.A(new_n14297), .Y(new_n14424));
  xor_4  g12076(.A(new_n14347), .B(new_n14295), .Y(new_n14425));
  nor_5  g12077(.A(new_n14425), .B(new_n14423), .Y(new_n14426));
  xor_4  g12078(.A(new_n9394), .B(new_n4801), .Y(new_n14427));
  xor_4  g12079(.A(new_n14427), .B(new_n14426), .Y(new_n14428));
  xor_4  g12080(.A(new_n14428), .B(pi422), .Y(new_n14429));
  xor_4  g12081(.A(new_n14429), .B(new_n14424), .Y(new_n14430));
  nand_5 g12082(.A(new_n14430), .B(new_n14423), .Y(new_n14431));
  nand_5 g12083(.A(new_n14431), .B(new_n14419), .Y(new_n14432));
  not_8  g12084(.A(new_n14430), .Y(po0150));
  nand_5 g12085(.A(po0150), .B(new_n14422), .Y(new_n14434));
  and_6  g12086(.A(new_n14434), .B(new_n14432), .Y(new_n14435));
  or_6   g12087(.A(new_n14435), .B(new_n14418), .Y(new_n14436));
  nand_5 g12088(.A(new_n14436), .B(new_n14416), .Y(new_n14437));
  nor_5  g12089(.A(new_n14437), .B(new_n14413), .Y(new_n14438));
  nor_5  g12090(.A(new_n14438), .B(new_n14412), .Y(new_n14439));
  nor_5  g12091(.A(new_n14439), .B(new_n14407), .Y(new_n14440));
  or_6   g12092(.A(new_n14440), .B(new_n14405), .Y(new_n14441));
  xor_4  g12093(.A(new_n14401), .B(new_n14399), .Y(new_n14442));
  nand_5 g12094(.A(new_n14442), .B(new_n14441), .Y(new_n14443));
  nand_5 g12095(.A(new_n14443), .B(new_n14402), .Y(new_n14444));
  nor_5  g12096(.A(new_n14444), .B(new_n14398), .Y(new_n14445));
  nor_5  g12097(.A(new_n14445), .B(new_n14397), .Y(new_n14446));
  xor_4  g12098(.A(new_n14391), .B(new_n14389), .Y(new_n14447));
  nor_5  g12099(.A(new_n14447), .B(new_n14446), .Y(new_n14448));
  or_6   g12100(.A(new_n14448), .B(new_n14392), .Y(new_n14449));
  nor_5  g12101(.A(new_n14449), .B(new_n14388), .Y(new_n14450));
  nor_5  g12102(.A(new_n14450), .B(new_n14386), .Y(new_n14451));
  or_6   g12103(.A(new_n14451), .B(new_n14382), .Y(new_n14452));
  nand_5 g12104(.A(new_n14381), .B(new_n14323), .Y(new_n14453));
  nand_5 g12105(.A(new_n14453), .B(new_n14452), .Y(new_n14454));
  xor_4  g12106(.A(new_n14319), .B(new_n14271), .Y(new_n14455));
  not_8  g12107(.A(new_n14455), .Y(new_n14456));
  nand_5 g12108(.A(new_n14333), .B(new_n4864), .Y(new_n14457));
  not_8  g12109(.A(new_n14380), .Y(new_n14458));
  nand_5 g12110(.A(new_n14458), .B(new_n14334), .Y(new_n14459));
  nand_5 g12111(.A(new_n14459), .B(new_n14457), .Y(new_n14460));
  nor_5  g12112(.A(new_n14332), .B(pi381), .Y(new_n14461));
  or_6   g12113(.A(new_n14461), .B(new_n4868), .Y(new_n14462));
  nand_5 g12114(.A(new_n14461), .B(new_n4868), .Y(new_n14463));
  nand_5 g12115(.A(new_n14463), .B(new_n14462), .Y(new_n14464));
  xor_4  g12116(.A(new_n14464), .B(new_n14460), .Y(new_n14465));
  xor_4  g12117(.A(new_n14465), .B(new_n14456), .Y(new_n14466));
  nand_5 g12118(.A(new_n14466), .B(new_n14454), .Y(new_n14467));
  nor_5  g12119(.A(new_n14467), .B(new_n14321), .Y(new_n14468));
  not_8  g12120(.A(new_n14460), .Y(new_n14469));
  nor_5  g12121(.A(new_n14462), .B(new_n14469), .Y(new_n14470));
  nor_5  g12122(.A(new_n14463), .B(new_n14460), .Y(new_n14471));
  nor_5  g12123(.A(new_n14471), .B(new_n14470), .Y(new_n14472));
  or_6   g12124(.A(new_n14465), .B(new_n14456), .Y(new_n14473));
  xor_4  g12125(.A(new_n14467), .B(new_n14320), .Y(new_n14474));
  nand_5 g12126(.A(new_n14474), .B(new_n14473), .Y(new_n14475));
  xor_4  g12127(.A(new_n14475), .B(new_n14472), .Y(po0762));
  and_6  g12128(.A(po0762), .B(new_n14321), .Y(new_n14477));
  nor_5  g12129(.A(new_n14477), .B(new_n14470), .Y(new_n14478));
  nor_5  g12130(.A(new_n14478), .B(new_n14468), .Y(po0131));
  xor_4  g12131(.A(pi162), .B(new_n4922), .Y(new_n14480));
  nand_5 g12132(.A(new_n4879), .B(pi352), .Y(new_n14481));
  xor_4  g12133(.A(pi752), .B(new_n5942), .Y(new_n14482));
  nand_5 g12134(.A(new_n4881), .B(pi081), .Y(new_n14483));
  xor_4  g12135(.A(pi676), .B(new_n5947), .Y(new_n14484));
  nand_5 g12136(.A(new_n4908), .B(pi019), .Y(new_n14485));
  xor_4  g12137(.A(pi634), .B(new_n7712), .Y(new_n14486));
  nand_5 g12138(.A(pi628), .B(new_n4900), .Y(new_n14487));
  not_8  g12139(.A(new_n9596), .Y(new_n14488));
  nand_5 g12140(.A(new_n14488), .B(new_n9592), .Y(new_n14489));
  nand_5 g12141(.A(new_n14489), .B(new_n14487), .Y(new_n14490));
  nand_5 g12142(.A(new_n14490), .B(new_n14486), .Y(new_n14491));
  nand_5 g12143(.A(new_n14491), .B(new_n14485), .Y(new_n14492));
  nand_5 g12144(.A(new_n14492), .B(new_n14484), .Y(new_n14493));
  nand_5 g12145(.A(new_n14493), .B(new_n14483), .Y(new_n14494));
  nand_5 g12146(.A(new_n14494), .B(new_n14482), .Y(new_n14495));
  nand_5 g12147(.A(new_n14495), .B(new_n14481), .Y(new_n14496));
  xor_4  g12148(.A(new_n14496), .B(new_n14480), .Y(new_n14497));
  xor_4  g12149(.A(new_n14497), .B(new_n3578), .Y(new_n14498));
  xor_4  g12150(.A(new_n14494), .B(new_n14482), .Y(new_n14499));
  not_8  g12151(.A(new_n14499), .Y(new_n14500));
  nand_5 g12152(.A(new_n14500), .B(new_n3612), .Y(new_n14501));
  xor_4  g12153(.A(new_n14499), .B(new_n3609), .Y(new_n14502));
  xor_4  g12154(.A(new_n14492), .B(new_n14484), .Y(new_n14503));
  or_6   g12155(.A(new_n14503), .B(new_n3602), .Y(new_n14504));
  xor_4  g12156(.A(new_n14490), .B(new_n14486), .Y(new_n14505));
  nor_5  g12157(.A(new_n14505), .B(new_n3579), .Y(new_n14506));
  xor_4  g12158(.A(new_n14505), .B(new_n3579), .Y(new_n14507));
  not_8  g12159(.A(new_n14507), .Y(new_n14508));
  not_8  g12160(.A(new_n9597), .Y(new_n14509));
  nand_5 g12161(.A(new_n14509), .B(new_n3580), .Y(new_n14510));
  xor_4  g12162(.A(new_n9597), .B(new_n3580), .Y(new_n14511));
  nand_5 g12163(.A(new_n9588), .B(new_n3589), .Y(new_n14512));
  xor_4  g12164(.A(new_n9588), .B(new_n3588), .Y(new_n14513));
  not_8  g12165(.A(new_n8609), .Y(new_n14514));
  nand_5 g12166(.A(new_n14514), .B(new_n13171), .Y(new_n14515));
  not_8  g12167(.A(new_n14515), .Y(new_n14516));
  or_6   g12168(.A(new_n14516), .B(new_n3583), .Y(new_n14517));
  nand_5 g12169(.A(new_n14516), .B(new_n3583), .Y(new_n14518));
  nand_5 g12170(.A(new_n14518), .B(new_n9576), .Y(new_n14519));
  nand_5 g12171(.A(new_n14519), .B(new_n14517), .Y(new_n14520));
  or_6   g12172(.A(new_n14520), .B(new_n14513), .Y(new_n14521));
  nand_5 g12173(.A(new_n14521), .B(new_n14512), .Y(new_n14522));
  or_6   g12174(.A(new_n14522), .B(new_n14511), .Y(new_n14523));
  nand_5 g12175(.A(new_n14523), .B(new_n14510), .Y(new_n14524));
  nor_5  g12176(.A(new_n14524), .B(new_n14508), .Y(new_n14525));
  or_6   g12177(.A(new_n14525), .B(new_n14506), .Y(new_n14526));
  not_8  g12178(.A(new_n14503), .Y(new_n14527));
  xor_4  g12179(.A(new_n14527), .B(new_n3602), .Y(new_n14528));
  not_8  g12180(.A(new_n14528), .Y(new_n14529));
  nand_5 g12181(.A(new_n14529), .B(new_n14526), .Y(new_n14530));
  nand_5 g12182(.A(new_n14530), .B(new_n14504), .Y(new_n14531));
  nand_5 g12183(.A(new_n14531), .B(new_n14502), .Y(new_n14532));
  nand_5 g12184(.A(new_n14532), .B(new_n14501), .Y(new_n14533));
  xor_4  g12185(.A(new_n14533), .B(new_n14498), .Y(new_n14534));
  not_8  g12186(.A(new_n14534), .Y(new_n14535));
  nand_5 g12187(.A(pi441), .B(new_n3432), .Y(new_n14536));
  xor_4  g12188(.A(pi441), .B(new_n3432), .Y(new_n14537));
  or_6   g12189(.A(pi300), .B(new_n3484), .Y(new_n14538));
  nand_5 g12190(.A(pi317), .B(new_n3435), .Y(new_n14539));
  nand_5 g12191(.A(pi681), .B(new_n3438), .Y(new_n14540));
  xor_4  g12192(.A(pi681), .B(new_n3438), .Y(new_n14541));
  nand_5 g12193(.A(new_n3441), .B(pi361), .Y(new_n14542));
  xor_4  g12194(.A(pi518), .B(new_n3489), .Y(new_n14543));
  nand_5 g12195(.A(pi787), .B(new_n3445), .Y(new_n14544));
  not_8  g12196(.A(new_n3635), .Y(new_n14545));
  xor_4  g12197(.A(pi787), .B(new_n3445), .Y(new_n14546));
  nand_5 g12198(.A(new_n14546), .B(new_n14545), .Y(new_n14547));
  nand_5 g12199(.A(new_n14547), .B(new_n14544), .Y(new_n14548));
  nand_5 g12200(.A(new_n14548), .B(new_n14543), .Y(new_n14549));
  nand_5 g12201(.A(new_n14549), .B(new_n14542), .Y(new_n14550));
  nand_5 g12202(.A(new_n14550), .B(new_n14541), .Y(new_n14551));
  nand_5 g12203(.A(new_n14551), .B(new_n14540), .Y(new_n14552));
  xor_4  g12204(.A(pi317), .B(new_n3435), .Y(new_n14553));
  nand_5 g12205(.A(new_n14553), .B(new_n14552), .Y(new_n14554));
  nand_5 g12206(.A(new_n14554), .B(new_n14539), .Y(new_n14555));
  nand_5 g12207(.A(new_n14555), .B(new_n3485), .Y(new_n14556));
  nand_5 g12208(.A(new_n14556), .B(new_n14538), .Y(new_n14557));
  nand_5 g12209(.A(new_n14557), .B(new_n14537), .Y(new_n14558));
  nand_5 g12210(.A(new_n14558), .B(new_n14536), .Y(new_n14559));
  xor_4  g12211(.A(pi616), .B(new_n3429), .Y(new_n14560));
  xor_4  g12212(.A(new_n14560), .B(new_n14559), .Y(new_n14561));
  or_6   g12213(.A(new_n14561), .B(new_n14535), .Y(new_n14562));
  xor_4  g12214(.A(new_n14561), .B(new_n14535), .Y(new_n14563));
  xor_4  g12215(.A(new_n14531), .B(new_n14502), .Y(new_n14564));
  xnor_4 g12216(.A(new_n14557), .B(new_n14537), .Y(new_n14565));
  nor_5  g12217(.A(new_n14565), .B(new_n14564), .Y(new_n14566));
  xnor_4 g12218(.A(new_n14555), .B(new_n3485), .Y(new_n14567));
  xor_4  g12219(.A(new_n14528), .B(new_n14526), .Y(new_n14568));
  not_8  g12220(.A(new_n14568), .Y(new_n14569));
  or_6   g12221(.A(new_n14569), .B(new_n14567), .Y(new_n14570));
  xor_4  g12222(.A(new_n14524), .B(new_n14507), .Y(new_n14571));
  xor_4  g12223(.A(new_n14553), .B(new_n14552), .Y(new_n14572));
  nor_5  g12224(.A(new_n14572), .B(new_n14571), .Y(new_n14573));
  xor_4  g12225(.A(new_n14572), .B(new_n14571), .Y(new_n14574));
  xnor_4 g12226(.A(new_n14522), .B(new_n14511), .Y(new_n14575));
  xnor_4 g12227(.A(new_n14550), .B(new_n14541), .Y(new_n14576));
  or_6   g12228(.A(new_n14576), .B(new_n14575), .Y(new_n14577));
  xor_4  g12229(.A(new_n14548), .B(new_n14543), .Y(new_n14578));
  xnor_4 g12230(.A(new_n14520), .B(new_n14513), .Y(new_n14579));
  nor_5  g12231(.A(new_n14579), .B(new_n14578), .Y(new_n14580));
  xor_4  g12232(.A(new_n14579), .B(new_n14578), .Y(new_n14581));
  xor_4  g12233(.A(new_n8609), .B(new_n3642), .Y(new_n14582));
  not_8  g12234(.A(new_n14582), .Y(new_n14583));
  nor_5  g12235(.A(new_n14583), .B(new_n3635), .Y(new_n14584));
  nand_5 g12236(.A(new_n14518), .B(new_n14517), .Y(new_n14585));
  xor_4  g12237(.A(new_n14585), .B(new_n9575), .Y(new_n14586));
  nand_5 g12238(.A(new_n14586), .B(new_n14546), .Y(new_n14587));
  nor_5  g12239(.A(new_n14587), .B(new_n14584), .Y(new_n14588));
  nor_5  g12240(.A(new_n14583), .B(new_n3634), .Y(new_n14589));
  not_8  g12241(.A(new_n14589), .Y(new_n14590));
  nand_5 g12242(.A(new_n14583), .B(new_n14545), .Y(new_n14591));
  nand_5 g12243(.A(new_n14591), .B(new_n14590), .Y(new_n14592));
  not_8  g12244(.A(new_n14586), .Y(new_n14593));
  xor_4  g12245(.A(new_n14593), .B(new_n14546), .Y(new_n14594));
  not_8  g12246(.A(new_n14594), .Y(new_n14595));
  nor_5  g12247(.A(new_n14595), .B(new_n14592), .Y(new_n14596));
  nand_5 g12248(.A(new_n14590), .B(new_n14547), .Y(new_n14597));
  nor_5  g12249(.A(new_n14597), .B(new_n14596), .Y(new_n14598));
  nor_5  g12250(.A(new_n14598), .B(new_n14588), .Y(new_n14599));
  and_6  g12251(.A(new_n14599), .B(new_n14581), .Y(new_n14600));
  nor_5  g12252(.A(new_n14600), .B(new_n14580), .Y(new_n14601));
  xor_4  g12253(.A(new_n14576), .B(new_n14575), .Y(new_n14602));
  nand_5 g12254(.A(new_n14602), .B(new_n14601), .Y(new_n14603));
  nand_5 g12255(.A(new_n14603), .B(new_n14577), .Y(new_n14604));
  not_8  g12256(.A(new_n14604), .Y(new_n14605));
  and_6  g12257(.A(new_n14605), .B(new_n14574), .Y(new_n14606));
  nor_5  g12258(.A(new_n14606), .B(new_n14573), .Y(new_n14607));
  xor_4  g12259(.A(new_n14569), .B(new_n14567), .Y(new_n14608));
  nand_5 g12260(.A(new_n14608), .B(new_n14607), .Y(new_n14609));
  nand_5 g12261(.A(new_n14609), .B(new_n14570), .Y(new_n14610));
  xor_4  g12262(.A(new_n14565), .B(new_n14564), .Y(new_n14611));
  nand_5 g12263(.A(new_n14611), .B(new_n14610), .Y(new_n14612));
  not_8  g12264(.A(new_n14612), .Y(new_n14613));
  nor_5  g12265(.A(new_n14613), .B(new_n14566), .Y(new_n14614));
  nand_5 g12266(.A(new_n14614), .B(new_n14563), .Y(new_n14615));
  nand_5 g12267(.A(new_n14615), .B(new_n14562), .Y(new_n14616));
  xor_4  g12268(.A(pi650), .B(new_n3426), .Y(new_n14617));
  nand_5 g12269(.A(pi616), .B(new_n3429), .Y(new_n14618));
  nand_5 g12270(.A(new_n14560), .B(new_n14559), .Y(new_n14619));
  nand_5 g12271(.A(new_n14619), .B(new_n14618), .Y(new_n14620));
  xor_4  g12272(.A(new_n14620), .B(new_n14617), .Y(new_n14621));
  xor_4  g12273(.A(pi093), .B(new_n7703), .Y(new_n14622));
  nand_5 g12274(.A(pi162), .B(new_n4922), .Y(new_n14623));
  nand_5 g12275(.A(new_n14496), .B(new_n14480), .Y(new_n14624));
  nand_5 g12276(.A(new_n14624), .B(new_n14623), .Y(new_n14625));
  xor_4  g12277(.A(new_n14625), .B(new_n14622), .Y(new_n14626));
  xor_4  g12278(.A(new_n14626), .B(new_n3576), .Y(new_n14627));
  or_6   g12279(.A(new_n14497), .B(new_n3578), .Y(new_n14628));
  nand_5 g12280(.A(new_n14533), .B(new_n14498), .Y(new_n14629));
  nand_5 g12281(.A(new_n14629), .B(new_n14628), .Y(new_n14630));
  xor_4  g12282(.A(new_n14630), .B(new_n14627), .Y(new_n14631));
  xor_4  g12283(.A(new_n14631), .B(new_n14621), .Y(new_n14632));
  xnor_4 g12284(.A(new_n14632), .B(new_n14616), .Y(po0132));
  not_8  g12285(.A(pi260), .Y(new_n14634));
  xor_4  g12286(.A(pi707), .B(new_n14634), .Y(new_n14635));
  or_6   g12287(.A(pi532), .B(new_n10477), .Y(new_n14636));
  xor_4  g12288(.A(pi532), .B(new_n10477), .Y(new_n14637));
  not_8  g12289(.A(pi060), .Y(new_n14638));
  nand_5 g12290(.A(pi568), .B(new_n14638), .Y(new_n14639));
  xor_4  g12291(.A(pi568), .B(new_n14638), .Y(new_n14640));
  nor_5  g12292(.A(pi730), .B(new_n4005), .Y(new_n14641));
  xor_4  g12293(.A(pi730), .B(pi183), .Y(new_n14642));
  not_8  g12294(.A(pi685), .Y(new_n14643));
  nand_5 g12295(.A(new_n14643), .B(pi245), .Y(new_n14644));
  nand_5 g12296(.A(new_n14644), .B(new_n3933), .Y(new_n14645));
  or_6   g12297(.A(new_n14644), .B(new_n3933), .Y(new_n14646));
  nand_5 g12298(.A(new_n14646), .B(pi577), .Y(new_n14647));
  nand_5 g12299(.A(new_n14647), .B(new_n14645), .Y(new_n14648));
  nor_5  g12300(.A(new_n14648), .B(new_n14642), .Y(new_n14649));
  or_6   g12301(.A(new_n14649), .B(new_n14641), .Y(new_n14650));
  nand_5 g12302(.A(new_n14650), .B(new_n14640), .Y(new_n14651));
  nand_5 g12303(.A(new_n14651), .B(new_n14639), .Y(new_n14652));
  nand_5 g12304(.A(new_n14652), .B(new_n14637), .Y(new_n14653));
  nand_5 g12305(.A(new_n14653), .B(new_n14636), .Y(new_n14654));
  xor_4  g12306(.A(new_n14654), .B(new_n14635), .Y(new_n14655));
  or_6   g12307(.A(new_n14655), .B(pi113), .Y(new_n14656));
  xor_4  g12308(.A(new_n14655), .B(pi113), .Y(new_n14657));
  xnor_4 g12309(.A(new_n14652), .B(new_n14637), .Y(new_n14658));
  or_6   g12310(.A(new_n14658), .B(new_n10987), .Y(new_n14659));
  xor_4  g12311(.A(new_n14658), .B(new_n10987), .Y(new_n14660));
  not_8  g12312(.A(new_n14660), .Y(new_n14661));
  xnor_4 g12313(.A(new_n14650), .B(new_n14640), .Y(new_n14662));
  nand_5 g12314(.A(new_n14662), .B(new_n11671), .Y(new_n14663));
  nor_5  g12315(.A(new_n14662), .B(new_n11671), .Y(new_n14664));
  xor_4  g12316(.A(new_n14648), .B(new_n14642), .Y(new_n14665));
  nor_5  g12317(.A(new_n14665), .B(pi371), .Y(new_n14666));
  nand_5 g12318(.A(new_n14646), .B(new_n14645), .Y(new_n14667));
  xor_4  g12319(.A(pi824), .B(pi577), .Y(new_n14668));
  xor_4  g12320(.A(new_n14668), .B(new_n14667), .Y(new_n14669));
  not_8  g12321(.A(new_n14669), .Y(new_n14670));
  xor_4  g12322(.A(pi685), .B(new_n3922), .Y(new_n14671));
  or_6   g12323(.A(new_n14671), .B(pi821), .Y(new_n14672));
  nand_5 g12324(.A(new_n14671), .B(pi821), .Y(new_n14673));
  nand_5 g12325(.A(new_n2564), .B(new_n7244), .Y(new_n14674));
  not_8  g12326(.A(new_n14674), .Y(new_n14675));
  nand_5 g12327(.A(new_n14675), .B(new_n14673), .Y(new_n14676));
  nand_5 g12328(.A(new_n14676), .B(new_n14672), .Y(new_n14677));
  or_6   g12329(.A(new_n14677), .B(new_n14670), .Y(new_n14678));
  nand_5 g12330(.A(new_n14670), .B(pi824), .Y(new_n14679));
  nand_5 g12331(.A(new_n14679), .B(new_n14678), .Y(new_n14680));
  xor_4  g12332(.A(new_n14665), .B(new_n11674), .Y(new_n14681));
  nor_5  g12333(.A(new_n14681), .B(new_n14680), .Y(new_n14682));
  nor_5  g12334(.A(new_n14682), .B(new_n14666), .Y(new_n14683));
  or_6   g12335(.A(new_n14683), .B(new_n14664), .Y(new_n14684));
  nand_5 g12336(.A(new_n14684), .B(new_n14663), .Y(new_n14685));
  or_6   g12337(.A(new_n14685), .B(new_n14661), .Y(new_n14686));
  nand_5 g12338(.A(new_n14686), .B(new_n14659), .Y(new_n14687));
  not_8  g12339(.A(new_n14687), .Y(new_n14688));
  nand_5 g12340(.A(new_n14688), .B(new_n14657), .Y(new_n14689));
  nand_5 g12341(.A(new_n14689), .B(new_n14656), .Y(new_n14690));
  nand_5 g12342(.A(pi707), .B(new_n14634), .Y(new_n14691));
  nand_5 g12343(.A(new_n14654), .B(new_n14635), .Y(new_n14692));
  nand_5 g12344(.A(new_n14692), .B(new_n14691), .Y(new_n14693));
  not_8  g12345(.A(new_n14693), .Y(new_n14694));
  nand_5 g12346(.A(new_n14694), .B(new_n14690), .Y(new_n14695));
  xor_4  g12347(.A(new_n14694), .B(new_n14690), .Y(new_n14696));
  xor_4  g12348(.A(pi803), .B(new_n11512), .Y(new_n14697));
  xor_4  g12349(.A(new_n14697), .B(new_n6259), .Y(new_n14698));
  nand_5 g12350(.A(new_n14698), .B(new_n14696), .Y(new_n14699));
  nand_5 g12351(.A(new_n14699), .B(new_n14695), .Y(new_n14700));
  not_8  g12352(.A(pi803), .Y(new_n14701));
  nand_5 g12353(.A(new_n14701), .B(pi598), .Y(new_n14702));
  nand_5 g12354(.A(new_n14697), .B(pi249), .Y(new_n14703));
  and_6  g12355(.A(new_n14703), .B(new_n14702), .Y(new_n14704));
  nand_5 g12356(.A(new_n14704), .B(new_n14700), .Y(new_n14705));
  not_8  g12357(.A(new_n14705), .Y(new_n14706));
  nand_5 g12358(.A(pi794), .B(new_n6295), .Y(new_n14707));
  not_8  g12359(.A(pi794), .Y(new_n14708));
  nand_5 g12360(.A(new_n14708), .B(pi789), .Y(new_n14709));
  nand_5 g12361(.A(new_n14709), .B(new_n11505), .Y(new_n14710));
  nand_5 g12362(.A(new_n14710), .B(new_n14707), .Y(new_n14711));
  nand_5 g12363(.A(new_n14711), .B(new_n14706), .Y(new_n14712));
  nor_5  g12364(.A(new_n14704), .B(new_n14700), .Y(new_n14713));
  not_8  g12365(.A(new_n14713), .Y(new_n14714));
  nor_5  g12366(.A(new_n14707), .B(pi135), .Y(new_n14715));
  nand_5 g12367(.A(new_n14715), .B(new_n14714), .Y(new_n14716));
  nand_5 g12368(.A(new_n14716), .B(new_n14712), .Y(new_n14717));
  not_8  g12369(.A(new_n14717), .Y(new_n14718));
  nor_5  g12370(.A(new_n14714), .B(new_n14711), .Y(new_n14719));
  nor_5  g12371(.A(new_n14709), .B(new_n11505), .Y(new_n14720));
  nand_5 g12372(.A(new_n14720), .B(new_n14705), .Y(new_n14721));
  not_8  g12373(.A(new_n14721), .Y(new_n14722));
  nor_5  g12374(.A(new_n14722), .B(new_n14719), .Y(new_n14723));
  nand_5 g12375(.A(new_n14723), .B(new_n14718), .Y(new_n14724));
  xor_4  g12376(.A(pi788), .B(new_n11499), .Y(new_n14725));
  xor_4  g12377(.A(new_n14725), .B(new_n6380), .Y(new_n14726));
  xor_4  g12378(.A(new_n14726), .B(new_n14724), .Y(new_n14727));
  nand_5 g12379(.A(new_n14727), .B(new_n10571), .Y(new_n14728));
  xnor_4 g12380(.A(new_n14698), .B(new_n14696), .Y(new_n14729));
  or_6   g12381(.A(new_n14729), .B(new_n10578), .Y(new_n14730));
  xor_4  g12382(.A(new_n14687), .B(new_n14657), .Y(new_n14731));
  or_6   g12383(.A(new_n14731), .B(new_n10583), .Y(new_n14732));
  xor_4  g12384(.A(new_n14731), .B(new_n10583), .Y(new_n14733));
  xor_4  g12385(.A(new_n14685), .B(new_n14660), .Y(new_n14734));
  not_8  g12386(.A(new_n14734), .Y(new_n14735));
  and_6  g12387(.A(new_n14735), .B(new_n10588), .Y(new_n14736));
  xor_4  g12388(.A(new_n14734), .B(new_n10588), .Y(new_n14737));
  xor_4  g12389(.A(new_n14662), .B(new_n11671), .Y(new_n14738));
  xor_4  g12390(.A(new_n14738), .B(new_n14683), .Y(new_n14739));
  nor_5  g12391(.A(new_n14739), .B(new_n10592), .Y(new_n14740));
  xor_4  g12392(.A(new_n14739), .B(new_n10591), .Y(new_n14741));
  xor_4  g12393(.A(new_n14681), .B(new_n14680), .Y(new_n14742));
  not_8  g12394(.A(new_n14742), .Y(new_n14743));
  nor_5  g12395(.A(new_n14743), .B(new_n10596), .Y(new_n14744));
  xor_4  g12396(.A(new_n14677), .B(new_n14670), .Y(new_n14745));
  not_8  g12397(.A(new_n14745), .Y(new_n14746));
  nand_5 g12398(.A(new_n14746), .B(new_n10600), .Y(new_n14747));
  xor_4  g12399(.A(new_n14746), .B(new_n10599), .Y(new_n14748));
  nor_5  g12400(.A(new_n6570), .B(new_n5786), .Y(new_n14749));
  nand_5 g12401(.A(new_n14749), .B(new_n6568), .Y(new_n14750));
  not_8  g12402(.A(new_n14750), .Y(new_n14751));
  nand_5 g12403(.A(new_n5786), .B(pi318), .Y(new_n14752));
  not_8  g12404(.A(new_n14752), .Y(new_n14753));
  nand_5 g12405(.A(pi799), .B(pi448), .Y(new_n14754));
  nor_5  g12406(.A(new_n14754), .B(new_n14753), .Y(new_n14755));
  nor_5  g12407(.A(new_n14755), .B(new_n14751), .Y(new_n14756));
  nand_5 g12408(.A(new_n14753), .B(new_n14675), .Y(new_n14757));
  nand_5 g12409(.A(new_n14757), .B(new_n14756), .Y(new_n14758));
  nand_5 g12410(.A(new_n14672), .B(new_n14673), .Y(new_n14759));
  xnor_4 g12411(.A(new_n14759), .B(new_n5804), .Y(new_n14760));
  xor_4  g12412(.A(new_n14760), .B(new_n14758), .Y(po1324));
  nand_5 g12413(.A(po1324), .B(new_n5804), .Y(new_n14762));
  nor_5  g12414(.A(new_n14759), .B(new_n5804), .Y(new_n14763));
  nor_5  g12415(.A(new_n14763), .B(new_n14756), .Y(new_n14764));
  nor_5  g12416(.A(new_n14752), .B(new_n5804), .Y(new_n14765));
  or_6   g12417(.A(new_n14759), .B(new_n14674), .Y(new_n14766));
  nor_5  g12418(.A(new_n14766), .B(new_n14765), .Y(new_n14767));
  nor_5  g12419(.A(new_n14767), .B(new_n14764), .Y(new_n14768));
  nand_5 g12420(.A(new_n14768), .B(new_n14762), .Y(new_n14769));
  or_6   g12421(.A(new_n14769), .B(new_n14748), .Y(new_n14770));
  nand_5 g12422(.A(new_n14770), .B(new_n14747), .Y(new_n14771));
  xor_4  g12423(.A(new_n14743), .B(new_n10596), .Y(new_n14772));
  and_6  g12424(.A(new_n14772), .B(new_n14771), .Y(new_n14773));
  nor_5  g12425(.A(new_n14773), .B(new_n14744), .Y(new_n14774));
  nor_5  g12426(.A(new_n14774), .B(new_n14741), .Y(new_n14775));
  or_6   g12427(.A(new_n14775), .B(new_n14740), .Y(new_n14776));
  nor_5  g12428(.A(new_n14776), .B(new_n14737), .Y(new_n14777));
  nor_5  g12429(.A(new_n14777), .B(new_n14736), .Y(new_n14778));
  nand_5 g12430(.A(new_n14778), .B(new_n14733), .Y(new_n14779));
  nand_5 g12431(.A(new_n14779), .B(new_n14732), .Y(new_n14780));
  xor_4  g12432(.A(new_n14729), .B(new_n10578), .Y(new_n14781));
  nand_5 g12433(.A(new_n14781), .B(new_n14780), .Y(new_n14782));
  nand_5 g12434(.A(new_n14782), .B(new_n14730), .Y(new_n14783));
  nand_5 g12435(.A(new_n14709), .B(new_n14707), .Y(new_n14784));
  nand_5 g12436(.A(new_n14714), .B(new_n14705), .Y(new_n14785));
  xor_4  g12437(.A(new_n14785), .B(new_n11505), .Y(new_n14786));
  xor_4  g12438(.A(new_n14786), .B(new_n14784), .Y(new_n14787));
  nor_5  g12439(.A(new_n14787), .B(new_n14783), .Y(new_n14788));
  xnor_4 g12440(.A(new_n14787), .B(new_n14783), .Y(new_n14789));
  nor_5  g12441(.A(new_n14789), .B(new_n10573), .Y(new_n14790));
  or_6   g12442(.A(new_n14790), .B(new_n14788), .Y(new_n14791));
  xor_4  g12443(.A(new_n14727), .B(new_n10571), .Y(new_n14792));
  nand_5 g12444(.A(new_n14792), .B(new_n14791), .Y(new_n14793));
  nand_5 g12445(.A(new_n14793), .B(new_n14728), .Y(new_n14794));
  nor_5  g12446(.A(pi788), .B(new_n6380), .Y(new_n14795));
  not_8  g12447(.A(new_n14795), .Y(new_n14796));
  nand_5 g12448(.A(pi788), .B(new_n6380), .Y(new_n14797));
  nand_5 g12449(.A(new_n14797), .B(pi148), .Y(new_n14798));
  nand_5 g12450(.A(new_n14798), .B(new_n14796), .Y(new_n14799));
  not_8  g12451(.A(new_n14799), .Y(new_n14800));
  nand_5 g12452(.A(new_n14800), .B(new_n14717), .Y(new_n14801));
  nor_5  g12453(.A(new_n14797), .B(pi148), .Y(new_n14802));
  nand_5 g12454(.A(new_n14802), .B(new_n14723), .Y(new_n14803));
  and_6  g12455(.A(new_n14803), .B(new_n14801), .Y(new_n14804));
  nand_5 g12456(.A(new_n14795), .B(pi148), .Y(new_n14805));
  nor_5  g12457(.A(new_n14805), .B(new_n14717), .Y(new_n14806));
  nor_5  g12458(.A(new_n14800), .B(new_n14723), .Y(new_n14807));
  nor_5  g12459(.A(new_n14807), .B(new_n14806), .Y(new_n14808));
  nand_5 g12460(.A(new_n14808), .B(new_n14804), .Y(new_n14809));
  xor_4  g12461(.A(new_n14809), .B(new_n10630), .Y(new_n14810));
  xnor_4 g12462(.A(new_n14810), .B(new_n14794), .Y(po0133));
  nor_5  g12463(.A(new_n2668), .B(new_n2612), .Y(new_n14812));
  nand_5 g12464(.A(new_n2611), .B(new_n2605), .Y(new_n14813));
  nand_5 g12465(.A(new_n14813), .B(new_n2606), .Y(new_n14814));
  nand_5 g12466(.A(new_n14814), .B(new_n2665), .Y(new_n14815));
  nor_5  g12467(.A(new_n14815), .B(new_n14812), .Y(new_n14816));
  not_8  g12468(.A(new_n14816), .Y(new_n14817));
  nor_5  g12469(.A(new_n6310), .B(pi198), .Y(new_n14818));
  xor_4  g12470(.A(new_n6309), .B(pi198), .Y(new_n14819));
  not_8  g12471(.A(new_n6207), .Y(new_n14820));
  nor_5  g12472(.A(new_n6134), .B(new_n6444), .Y(new_n14821));
  nand_5 g12473(.A(new_n6135), .B(pi284), .Y(new_n14822));
  xor_4  g12474(.A(new_n6133), .B(new_n6444), .Y(new_n14823));
  nor_5  g12475(.A(new_n14823), .B(new_n14822), .Y(new_n14824));
  or_6   g12476(.A(new_n14824), .B(new_n14821), .Y(new_n14825));
  nor_5  g12477(.A(new_n14825), .B(new_n6132), .Y(new_n14826));
  xor_4  g12478(.A(new_n14825), .B(new_n6132), .Y(new_n14827));
  nand_5 g12479(.A(new_n14827), .B(new_n6434), .Y(new_n14828));
  not_8  g12480(.A(new_n14828), .Y(new_n14829));
  nor_5  g12481(.A(new_n14829), .B(new_n14826), .Y(new_n14830));
  nand_5 g12482(.A(new_n14830), .B(new_n6157), .Y(new_n14831));
  xor_4  g12483(.A(new_n14830), .B(new_n6158), .Y(new_n14832));
  or_6   g12484(.A(new_n14832), .B(new_n6432), .Y(new_n14833));
  nand_5 g12485(.A(new_n14833), .B(new_n14831), .Y(new_n14834));
  or_6   g12486(.A(new_n14834), .B(new_n6170), .Y(new_n14835));
  xor_4  g12487(.A(new_n14834), .B(new_n6170), .Y(new_n14836));
  nand_5 g12488(.A(new_n14836), .B(new_n6429), .Y(new_n14837));
  nand_5 g12489(.A(new_n14837), .B(new_n14835), .Y(new_n14838));
  nand_5 g12490(.A(new_n14838), .B(new_n14820), .Y(new_n14839));
  xor_4  g12491(.A(new_n14838), .B(new_n14820), .Y(new_n14840));
  nand_5 g12492(.A(new_n14840), .B(new_n6556), .Y(new_n14841));
  nand_5 g12493(.A(new_n14841), .B(new_n14839), .Y(new_n14842));
  nand_5 g12494(.A(new_n14842), .B(new_n6280), .Y(new_n14843));
  xor_4  g12495(.A(new_n14842), .B(new_n6280), .Y(new_n14844));
  nand_5 g12496(.A(new_n14844), .B(new_n6554), .Y(new_n14845));
  nand_5 g12497(.A(new_n14845), .B(new_n14843), .Y(new_n14846));
  or_6   g12498(.A(new_n14846), .B(new_n6311), .Y(new_n14847));
  nand_5 g12499(.A(new_n14846), .B(new_n6311), .Y(new_n14848));
  nand_5 g12500(.A(new_n14848), .B(pi112), .Y(new_n14849));
  nand_5 g12501(.A(new_n14849), .B(new_n14847), .Y(new_n14850));
  nor_5  g12502(.A(new_n14850), .B(new_n14819), .Y(new_n14851));
  nor_5  g12503(.A(new_n14851), .B(new_n14818), .Y(new_n14852));
  nor_5  g12504(.A(new_n14852), .B(new_n6347), .Y(new_n14853));
  xor_4  g12505(.A(new_n14852), .B(new_n6347), .Y(new_n14854));
  nand_5 g12506(.A(new_n14854), .B(new_n12597), .Y(new_n14855));
  not_8  g12507(.A(new_n14855), .Y(new_n14856));
  nor_5  g12508(.A(new_n14856), .B(new_n14853), .Y(new_n14857));
  nor_5  g12509(.A(new_n14857), .B(new_n6378), .Y(new_n14858));
  xor_4  g12510(.A(new_n14854), .B(pi170), .Y(new_n14859));
  nor_5  g12511(.A(new_n14859), .B(new_n2669), .Y(new_n14860));
  not_8  g12512(.A(new_n2669), .Y(new_n14861));
  xor_4  g12513(.A(new_n14859), .B(new_n14861), .Y(new_n14862));
  xor_4  g12514(.A(new_n14850), .B(new_n14819), .Y(new_n14863));
  or_6   g12515(.A(new_n14863), .B(new_n2826), .Y(new_n14864));
  nand_5 g12516(.A(new_n14848), .B(new_n14847), .Y(new_n14865));
  xor_4  g12517(.A(new_n14865), .B(pi112), .Y(new_n14866));
  nor_5  g12518(.A(new_n14866), .B(new_n2742), .Y(new_n14867));
  xor_4  g12519(.A(new_n14866), .B(new_n2741), .Y(new_n14868));
  xor_4  g12520(.A(new_n14844), .B(pi053), .Y(new_n14869));
  nor_5  g12521(.A(new_n14869), .B(new_n2797), .Y(new_n14870));
  xor_4  g12522(.A(new_n14840), .B(pi154), .Y(new_n14871));
  nor_5  g12523(.A(new_n14871), .B(new_n2788), .Y(new_n14872));
  xor_4  g12524(.A(new_n14871), .B(new_n2789), .Y(new_n14873));
  xor_4  g12525(.A(new_n14836), .B(pi267), .Y(new_n14874));
  nor_5  g12526(.A(new_n14874), .B(new_n2779), .Y(new_n14875));
  not_8  g12527(.A(new_n2779), .Y(new_n14876));
  xor_4  g12528(.A(new_n14874), .B(new_n14876), .Y(new_n14877));
  xor_4  g12529(.A(new_n14832), .B(pi312), .Y(new_n14878));
  and_6  g12530(.A(new_n14878), .B(new_n2770), .Y(new_n14879));
  xor_4  g12531(.A(new_n14878), .B(new_n2771), .Y(new_n14880));
  xor_4  g12532(.A(new_n14827), .B(pi471), .Y(new_n14881));
  nor_5  g12533(.A(new_n14881), .B(new_n2763), .Y(new_n14882));
  nand_5 g12534(.A(new_n2754), .B(new_n2744), .Y(new_n14883));
  nand_5 g12535(.A(new_n14883), .B(new_n14824), .Y(new_n14884));
  or_6   g12536(.A(new_n14823), .B(new_n2745), .Y(new_n14885));
  nor_5  g12537(.A(new_n6135), .B(pi284), .Y(new_n14886));
  nand_5 g12538(.A(new_n14886), .B(new_n2755), .Y(new_n14887));
  or_6   g12539(.A(new_n14822), .B(new_n2755), .Y(new_n14888));
  nand_5 g12540(.A(new_n14888), .B(new_n14887), .Y(new_n14889));
  xor_4  g12541(.A(new_n14823), .B(new_n2745), .Y(new_n14890));
  or_6   g12542(.A(new_n14890), .B(new_n14889), .Y(new_n14891));
  nand_5 g12543(.A(new_n14891), .B(new_n14887), .Y(new_n14892));
  nand_5 g12544(.A(new_n14892), .B(new_n14885), .Y(new_n14893));
  and_6  g12545(.A(new_n14893), .B(new_n14884), .Y(new_n14894));
  xor_4  g12546(.A(new_n14881), .B(new_n2765), .Y(new_n14895));
  nor_5  g12547(.A(new_n14895), .B(new_n14894), .Y(new_n14896));
  nor_5  g12548(.A(new_n14896), .B(new_n14882), .Y(new_n14897));
  nor_5  g12549(.A(new_n14897), .B(new_n14880), .Y(new_n14898));
  nor_5  g12550(.A(new_n14898), .B(new_n14879), .Y(new_n14899));
  nor_5  g12551(.A(new_n14899), .B(new_n14877), .Y(new_n14900));
  nor_5  g12552(.A(new_n14900), .B(new_n14875), .Y(new_n14901));
  nor_5  g12553(.A(new_n14901), .B(new_n14873), .Y(new_n14902));
  nor_5  g12554(.A(new_n14902), .B(new_n14872), .Y(new_n14903));
  xor_4  g12555(.A(new_n14869), .B(new_n2801), .Y(new_n14904));
  nor_5  g12556(.A(new_n14904), .B(new_n14903), .Y(new_n14905));
  or_6   g12557(.A(new_n14905), .B(new_n14870), .Y(new_n14906));
  nor_5  g12558(.A(new_n14906), .B(new_n14868), .Y(new_n14907));
  or_6   g12559(.A(new_n14907), .B(new_n14867), .Y(new_n14908));
  xor_4  g12560(.A(new_n14863), .B(new_n2826), .Y(new_n14909));
  nand_5 g12561(.A(new_n14909), .B(new_n14908), .Y(new_n14910));
  nand_5 g12562(.A(new_n14910), .B(new_n14864), .Y(new_n14911));
  nor_5  g12563(.A(new_n14911), .B(new_n14862), .Y(new_n14912));
  or_6   g12564(.A(new_n14912), .B(new_n14860), .Y(new_n14913));
  nand_5 g12565(.A(new_n14913), .B(new_n14858), .Y(new_n14914));
  nor_5  g12566(.A(new_n14814), .B(new_n2665), .Y(new_n14915));
  nor_5  g12567(.A(new_n2609), .B(new_n2605), .Y(new_n14916));
  nand_5 g12568(.A(new_n14916), .B(new_n2667), .Y(new_n14917));
  not_8  g12569(.A(new_n14917), .Y(new_n14918));
  nor_5  g12570(.A(new_n14918), .B(new_n14915), .Y(new_n14919));
  nand_5 g12571(.A(new_n14857), .B(new_n6378), .Y(new_n14920));
  and_6  g12572(.A(new_n14920), .B(new_n14913), .Y(new_n14921));
  or_6   g12573(.A(new_n14921), .B(new_n14858), .Y(new_n14922));
  nand_5 g12574(.A(new_n14922), .B(new_n14919), .Y(new_n14923));
  nand_5 g12575(.A(new_n14923), .B(new_n14914), .Y(new_n14924));
  nand_5 g12576(.A(new_n14924), .B(new_n14817), .Y(new_n14925));
  not_8  g12577(.A(new_n14914), .Y(new_n14926));
  nor_5  g12578(.A(new_n14920), .B(new_n14913), .Y(new_n14927));
  not_8  g12579(.A(new_n14927), .Y(new_n14928));
  nand_5 g12580(.A(new_n14928), .B(new_n14816), .Y(new_n14929));
  nor_5  g12581(.A(new_n14929), .B(new_n14926), .Y(new_n14930));
  nor_5  g12582(.A(new_n14928), .B(new_n14919), .Y(new_n14931));
  nor_5  g12583(.A(new_n14931), .B(new_n14930), .Y(new_n14932));
  nand_5 g12584(.A(new_n14932), .B(new_n14925), .Y(po0134));
  xor_4  g12585(.A(pi406), .B(new_n9488), .Y(new_n14934));
  nand_5 g12586(.A(pi151), .B(new_n2912), .Y(new_n14935));
  xor_4  g12587(.A(pi151), .B(new_n2912), .Y(new_n14936));
  nand_5 g12588(.A(new_n5287), .B(pi570), .Y(new_n14937));
  xor_4  g12589(.A(pi801), .B(new_n5246), .Y(new_n14938));
  nand_5 g12590(.A(pi144), .B(new_n2920), .Y(new_n14939));
  nand_5 g12591(.A(new_n5354), .B(pi181), .Y(new_n14940));
  nand_5 g12592(.A(new_n14940), .B(new_n14939), .Y(new_n14941));
  nand_5 g12593(.A(new_n14941), .B(new_n14938), .Y(new_n14942));
  nand_5 g12594(.A(new_n14942), .B(new_n14937), .Y(new_n14943));
  nand_5 g12595(.A(new_n14943), .B(new_n14936), .Y(new_n14944));
  nand_5 g12596(.A(new_n14944), .B(new_n14935), .Y(new_n14945));
  xnor_4 g12597(.A(new_n14945), .B(new_n14934), .Y(new_n14946));
  nor_5  g12598(.A(new_n14946), .B(new_n4250), .Y(new_n14947));
  xnor_4 g12599(.A(new_n14946), .B(new_n4250), .Y(new_n14948));
  xnor_4 g12600(.A(new_n14943), .B(new_n14936), .Y(new_n14949));
  nor_5  g12601(.A(new_n14949), .B(new_n4200), .Y(new_n14950));
  xnor_4 g12602(.A(new_n14949), .B(new_n4200), .Y(new_n14951));
  xnor_4 g12603(.A(new_n14941), .B(new_n14938), .Y(new_n14952));
  nor_5  g12604(.A(new_n14952), .B(new_n4221), .Y(new_n14953));
  not_8  g12605(.A(new_n4207), .Y(new_n14954));
  nand_5 g12606(.A(new_n5339), .B(new_n14954), .Y(new_n14955));
  nand_5 g12607(.A(new_n5341), .B(new_n4207), .Y(new_n14956));
  nand_5 g12608(.A(new_n14956), .B(new_n14955), .Y(new_n14957));
  xor_4  g12609(.A(new_n14957), .B(new_n5355), .Y(new_n14958));
  nand_5 g12610(.A(new_n14958), .B(new_n4214), .Y(new_n14959));
  nand_5 g12611(.A(new_n14957), .B(new_n5354), .Y(new_n14960));
  nand_5 g12612(.A(new_n14956), .B(new_n14940), .Y(new_n14961));
  nand_5 g12613(.A(new_n14961), .B(new_n14960), .Y(new_n14962));
  nand_5 g12614(.A(new_n14962), .B(new_n14959), .Y(new_n14963));
  xor_4  g12615(.A(new_n14952), .B(new_n4220), .Y(new_n14964));
  nor_5  g12616(.A(new_n14964), .B(new_n14963), .Y(new_n14965));
  nor_5  g12617(.A(new_n14965), .B(new_n14953), .Y(new_n14966));
  nor_5  g12618(.A(new_n14966), .B(new_n14951), .Y(new_n14967));
  nor_5  g12619(.A(new_n14967), .B(new_n14950), .Y(new_n14968));
  nor_5  g12620(.A(new_n14968), .B(new_n14948), .Y(new_n14969));
  nor_5  g12621(.A(new_n14969), .B(new_n14947), .Y(new_n14970));
  xor_4  g12622(.A(pi177), .B(new_n7263), .Y(new_n14971));
  nand_5 g12623(.A(pi432), .B(new_n3846), .Y(new_n14972));
  not_8  g12624(.A(new_n14972), .Y(new_n14973));
  not_8  g12625(.A(new_n4239), .Y(new_n14974));
  nor_5  g12626(.A(new_n4243), .B(new_n14974), .Y(new_n14975));
  nor_5  g12627(.A(new_n14975), .B(new_n14973), .Y(new_n14976));
  xor_4  g12628(.A(new_n14976), .B(new_n14971), .Y(new_n14977));
  not_8  g12629(.A(new_n14977), .Y(new_n14978));
  nand_5 g12630(.A(new_n4248), .B(new_n4244), .Y(new_n14979));
  or_6   g12631(.A(new_n4249), .B(new_n4238), .Y(new_n14980));
  nand_5 g12632(.A(new_n14980), .B(new_n14979), .Y(new_n14981));
  xor_4  g12633(.A(new_n14981), .B(new_n14978), .Y(new_n14982));
  xor_4  g12634(.A(new_n14982), .B(new_n11182), .Y(new_n14983));
  not_8  g12635(.A(new_n14983), .Y(new_n14984));
  nand_5 g12636(.A(new_n2909), .B(pi172), .Y(new_n14985));
  nand_5 g12637(.A(new_n14945), .B(new_n14934), .Y(new_n14986));
  nand_5 g12638(.A(new_n14986), .B(new_n14985), .Y(new_n14987));
  xor_4  g12639(.A(pi229), .B(pi061), .Y(new_n14988));
  xor_4  g12640(.A(new_n14988), .B(new_n14987), .Y(new_n14989));
  xor_4  g12641(.A(new_n14989), .B(new_n14984), .Y(new_n14990));
  not_8  g12642(.A(new_n14990), .Y(new_n14991));
  xor_4  g12643(.A(new_n14991), .B(new_n14970), .Y(po0135));
  xor_4  g12644(.A(new_n14010), .B(new_n12936), .Y(po0136));
  xor_4  g12645(.A(pi381), .B(new_n13053), .Y(new_n14994));
  nand_5 g12646(.A(new_n7483), .B(pi541), .Y(new_n14995));
  xor_4  g12647(.A(pi607), .B(new_n10966), .Y(new_n14996));
  nand_5 g12648(.A(pi164), .B(new_n7471), .Y(new_n14997));
  xor_4  g12649(.A(pi164), .B(new_n7471), .Y(new_n14998));
  nand_5 g12650(.A(pi484), .B(new_n3710), .Y(new_n14999));
  xor_4  g12651(.A(pi484), .B(new_n3710), .Y(new_n15000));
  nand_5 g12652(.A(pi814), .B(new_n3714), .Y(new_n15001));
  xor_4  g12653(.A(pi814), .B(new_n3714), .Y(new_n15002));
  nand_5 g12654(.A(pi604), .B(new_n3718), .Y(new_n15003));
  nand_5 g12655(.A(new_n4230), .B(new_n4226), .Y(new_n15004));
  nand_5 g12656(.A(new_n15004), .B(new_n15003), .Y(new_n15005));
  nand_5 g12657(.A(new_n15005), .B(new_n15002), .Y(new_n15006));
  nand_5 g12658(.A(new_n15006), .B(new_n15001), .Y(new_n15007));
  nand_5 g12659(.A(new_n15007), .B(new_n15000), .Y(new_n15008));
  nand_5 g12660(.A(new_n15008), .B(new_n14999), .Y(new_n15009));
  nand_5 g12661(.A(new_n15009), .B(new_n14998), .Y(new_n15010));
  nand_5 g12662(.A(new_n15010), .B(new_n14997), .Y(new_n15011));
  nand_5 g12663(.A(new_n15011), .B(new_n14996), .Y(new_n15012));
  nand_5 g12664(.A(new_n15012), .B(new_n14995), .Y(new_n15013));
  xor_4  g12665(.A(new_n15013), .B(new_n14994), .Y(new_n15014));
  xor_4  g12666(.A(new_n15011), .B(new_n14996), .Y(new_n15015));
  xor_4  g12667(.A(new_n15009), .B(new_n14998), .Y(new_n15016));
  xor_4  g12668(.A(new_n15005), .B(new_n15002), .Y(new_n15017));
  not_8  g12669(.A(new_n15017), .Y(new_n15018));
  nand_5 g12670(.A(new_n4250), .B(new_n4232), .Y(new_n15019));
  nand_5 g12671(.A(new_n4251), .B(new_n4225), .Y(new_n15020));
  nand_5 g12672(.A(new_n15020), .B(new_n15019), .Y(new_n15021));
  nor_5  g12673(.A(new_n15021), .B(new_n15018), .Y(new_n15022));
  xor_4  g12674(.A(new_n15021), .B(new_n15017), .Y(new_n15023));
  nor_5  g12675(.A(new_n15023), .B(new_n14983), .Y(new_n15024));
  or_6   g12676(.A(new_n15024), .B(new_n15022), .Y(new_n15025));
  nand_5 g12677(.A(new_n3805), .B(pi120), .Y(new_n15026));
  not_8  g12678(.A(new_n14976), .Y(new_n15027));
  nand_5 g12679(.A(new_n15027), .B(new_n14971), .Y(new_n15028));
  nand_5 g12680(.A(new_n15028), .B(new_n15026), .Y(new_n15029));
  nand_5 g12681(.A(pi146), .B(new_n5941), .Y(new_n15030));
  nand_5 g12682(.A(new_n5940), .B(pi143), .Y(new_n15031));
  and_6  g12683(.A(new_n15031), .B(new_n15030), .Y(new_n15032));
  xor_4  g12684(.A(new_n15032), .B(new_n15029), .Y(new_n15033));
  nand_5 g12685(.A(new_n14981), .B(new_n14977), .Y(new_n15034));
  or_6   g12686(.A(new_n14982), .B(new_n11182), .Y(new_n15035));
  nand_5 g12687(.A(new_n15035), .B(new_n15034), .Y(new_n15036));
  nand_5 g12688(.A(new_n15036), .B(new_n11177), .Y(new_n15037));
  nor_5  g12689(.A(new_n15036), .B(new_n11177), .Y(new_n15038));
  not_8  g12690(.A(new_n15038), .Y(new_n15039));
  nand_5 g12691(.A(new_n15039), .B(new_n15037), .Y(new_n15040));
  xor_4  g12692(.A(new_n15040), .B(new_n15033), .Y(new_n15041));
  not_8  g12693(.A(new_n15041), .Y(new_n15042));
  nand_5 g12694(.A(new_n15042), .B(new_n15025), .Y(new_n15043));
  xor_4  g12695(.A(new_n15007), .B(new_n15000), .Y(new_n15044));
  not_8  g12696(.A(new_n15044), .Y(new_n15045));
  xor_4  g12697(.A(new_n15041), .B(new_n15025), .Y(new_n15046));
  or_6   g12698(.A(new_n15046), .B(new_n15045), .Y(new_n15047));
  nand_5 g12699(.A(new_n15047), .B(new_n15043), .Y(new_n15048));
  nand_5 g12700(.A(new_n15048), .B(new_n15016), .Y(new_n15049));
  xor_4  g12701(.A(pi621), .B(new_n12002), .Y(new_n15050));
  nand_5 g12702(.A(new_n15031), .B(new_n15029), .Y(new_n15051));
  nand_5 g12703(.A(new_n15051), .B(new_n15030), .Y(new_n15052));
  xor_4  g12704(.A(new_n15052), .B(new_n15050), .Y(new_n15053));
  not_8  g12705(.A(new_n15033), .Y(new_n15054));
  nand_5 g12706(.A(new_n15039), .B(new_n15054), .Y(new_n15055));
  nand_5 g12707(.A(new_n15055), .B(new_n15037), .Y(new_n15056));
  xor_4  g12708(.A(new_n15056), .B(new_n15053), .Y(new_n15057));
  xor_4  g12709(.A(new_n15057), .B(new_n11171), .Y(new_n15058));
  xnor_4 g12710(.A(new_n15048), .B(new_n15016), .Y(new_n15059));
  or_6   g12711(.A(new_n15059), .B(new_n15058), .Y(new_n15060));
  nand_5 g12712(.A(new_n15060), .B(new_n15049), .Y(new_n15061));
  nor_5  g12713(.A(new_n15061), .B(new_n15015), .Y(new_n15062));
  xor_4  g12714(.A(new_n15061), .B(new_n15015), .Y(new_n15063));
  xor_4  g12715(.A(pi185), .B(new_n7255), .Y(new_n15064));
  nand_5 g12716(.A(pi621), .B(new_n12002), .Y(new_n15065));
  nand_5 g12717(.A(new_n15052), .B(new_n15050), .Y(new_n15066));
  nand_5 g12718(.A(new_n15066), .B(new_n15065), .Y(new_n15067));
  xor_4  g12719(.A(new_n15067), .B(new_n15064), .Y(new_n15068));
  not_8  g12720(.A(new_n15068), .Y(new_n15069));
  not_8  g12721(.A(new_n15053), .Y(new_n15070));
  nand_5 g12722(.A(new_n15056), .B(new_n15070), .Y(new_n15071));
  not_8  g12723(.A(new_n15071), .Y(new_n15072));
  nor_5  g12724(.A(new_n15057), .B(new_n11171), .Y(new_n15073));
  nor_5  g12725(.A(new_n15073), .B(new_n15072), .Y(new_n15074));
  xor_4  g12726(.A(new_n15074), .B(new_n15069), .Y(new_n15075));
  xor_4  g12727(.A(new_n15075), .B(new_n11168), .Y(new_n15076));
  nand_5 g12728(.A(new_n15076), .B(new_n15063), .Y(new_n15077));
  not_8  g12729(.A(new_n15077), .Y(new_n15078));
  nor_5  g12730(.A(new_n15078), .B(new_n15062), .Y(new_n15079));
  nand_5 g12731(.A(new_n15079), .B(new_n15014), .Y(new_n15080));
  nand_5 g12732(.A(new_n11995), .B(pi092), .Y(new_n15081));
  nand_5 g12733(.A(new_n15067), .B(new_n15064), .Y(new_n15082));
  nand_5 g12734(.A(new_n15082), .B(new_n15081), .Y(new_n15083));
  xor_4  g12735(.A(new_n15083), .B(new_n6092), .Y(new_n15084));
  not_8  g12736(.A(new_n15084), .Y(new_n15085));
  xor_4  g12737(.A(new_n15085), .B(new_n11163), .Y(new_n15086));
  nand_5 g12738(.A(new_n15074), .B(new_n15068), .Y(new_n15087));
  or_6   g12739(.A(new_n15075), .B(new_n11220), .Y(new_n15088));
  nand_5 g12740(.A(new_n15088), .B(new_n15087), .Y(new_n15089));
  xor_4  g12741(.A(new_n15089), .B(new_n15086), .Y(new_n15090));
  xnor_4 g12742(.A(new_n15079), .B(new_n15014), .Y(new_n15091));
  not_8  g12743(.A(new_n15091), .Y(new_n15092));
  nand_5 g12744(.A(new_n15092), .B(new_n15090), .Y(new_n15093));
  nand_5 g12745(.A(new_n15093), .B(new_n15080), .Y(new_n15094));
  nand_5 g12746(.A(new_n7494), .B(pi292), .Y(new_n15095));
  nand_5 g12747(.A(new_n15013), .B(new_n14994), .Y(new_n15096));
  nand_5 g12748(.A(new_n15096), .B(new_n15095), .Y(new_n15097));
  not_8  g12749(.A(new_n15097), .Y(new_n15098));
  xor_4  g12750(.A(new_n15098), .B(new_n15094), .Y(new_n15099));
  nand_5 g12751(.A(new_n11994), .B(pi280), .Y(new_n15100));
  nand_5 g12752(.A(new_n15083), .B(new_n6092), .Y(new_n15101));
  nand_5 g12753(.A(new_n15101), .B(new_n15100), .Y(new_n15102));
  xor_4  g12754(.A(new_n15102), .B(new_n11159), .Y(new_n15103));
  or_6   g12755(.A(new_n15085), .B(new_n11163), .Y(new_n15104));
  nand_5 g12756(.A(new_n15089), .B(new_n15086), .Y(new_n15105));
  nand_5 g12757(.A(new_n15105), .B(new_n15104), .Y(new_n15106));
  xor_4  g12758(.A(new_n15106), .B(new_n15103), .Y(new_n15107));
  xnor_4 g12759(.A(new_n15107), .B(new_n15099), .Y(po0137));
  xor_4  g12760(.A(pi701), .B(new_n2837), .Y(new_n15109));
  nand_5 g12761(.A(pi279), .B(new_n2814), .Y(new_n15110));
  xor_4  g12762(.A(pi279), .B(new_n2814), .Y(new_n15111));
  nand_5 g12763(.A(pi786), .B(new_n2857), .Y(new_n15112));
  xor_4  g12764(.A(pi786), .B(new_n2857), .Y(new_n15113));
  nand_5 g12765(.A(new_n2675), .B(pi187), .Y(new_n15114));
  xor_4  g12766(.A(pi407), .B(new_n10233), .Y(new_n15115));
  nand_5 g12767(.A(pi720), .B(new_n2864), .Y(new_n15116));
  xor_4  g12768(.A(pi720), .B(new_n2864), .Y(new_n15117));
  nand_5 g12769(.A(new_n2867), .B(pi339), .Y(new_n15118));
  not_8  g12770(.A(new_n13748), .Y(new_n15119));
  nand_5 g12771(.A(new_n15119), .B(new_n13738), .Y(new_n15120));
  nand_5 g12772(.A(new_n15120), .B(new_n15118), .Y(new_n15121));
  nand_5 g12773(.A(new_n15121), .B(new_n15117), .Y(new_n15122));
  nand_5 g12774(.A(new_n15122), .B(new_n15116), .Y(new_n15123));
  nand_5 g12775(.A(new_n15123), .B(new_n15115), .Y(new_n15124));
  nand_5 g12776(.A(new_n15124), .B(new_n15114), .Y(new_n15125));
  nand_5 g12777(.A(new_n15125), .B(new_n15113), .Y(new_n15126));
  nand_5 g12778(.A(new_n15126), .B(new_n15112), .Y(new_n15127));
  nand_5 g12779(.A(new_n15127), .B(new_n15111), .Y(new_n15128));
  nand_5 g12780(.A(new_n15128), .B(new_n15110), .Y(new_n15129));
  xor_4  g12781(.A(new_n15129), .B(new_n15109), .Y(new_n15130));
  xor_4  g12782(.A(new_n15127), .B(new_n15111), .Y(new_n15131));
  nand_5 g12783(.A(new_n15131), .B(new_n7318), .Y(new_n15132));
  xor_4  g12784(.A(new_n15131), .B(new_n7318), .Y(new_n15133));
  xor_4  g12785(.A(new_n15125), .B(new_n15113), .Y(new_n15134));
  not_8  g12786(.A(new_n15134), .Y(new_n15135));
  xor_4  g12787(.A(new_n15123), .B(new_n15115), .Y(new_n15136));
  not_8  g12788(.A(new_n15136), .Y(new_n15137));
  xor_4  g12789(.A(new_n15121), .B(new_n15117), .Y(new_n15138));
  not_8  g12790(.A(new_n15138), .Y(new_n15139));
  nand_5 g12791(.A(new_n13749), .B(new_n7338), .Y(new_n15140));
  nand_5 g12792(.A(new_n14042), .B(new_n14030), .Y(new_n15141));
  nand_5 g12793(.A(new_n15141), .B(new_n15140), .Y(new_n15142));
  nand_5 g12794(.A(new_n15142), .B(new_n15139), .Y(new_n15143));
  xor_4  g12795(.A(new_n15142), .B(new_n15138), .Y(new_n15144));
  or_6   g12796(.A(new_n15144), .B(new_n7332), .Y(new_n15145));
  nand_5 g12797(.A(new_n15145), .B(new_n15143), .Y(new_n15146));
  nand_5 g12798(.A(new_n15146), .B(new_n15137), .Y(new_n15147));
  xor_4  g12799(.A(new_n15146), .B(new_n15136), .Y(new_n15148));
  or_6   g12800(.A(new_n15148), .B(new_n7328), .Y(new_n15149));
  nand_5 g12801(.A(new_n15149), .B(new_n15147), .Y(new_n15150));
  nand_5 g12802(.A(new_n15150), .B(new_n15135), .Y(new_n15151));
  not_8  g12803(.A(new_n15151), .Y(new_n15152));
  xor_4  g12804(.A(new_n15150), .B(new_n15134), .Y(new_n15153));
  nor_5  g12805(.A(new_n15153), .B(new_n7324), .Y(new_n15154));
  nor_5  g12806(.A(new_n15154), .B(new_n15152), .Y(new_n15155));
  nand_5 g12807(.A(new_n15155), .B(new_n15133), .Y(new_n15156));
  nand_5 g12808(.A(new_n15156), .B(new_n15132), .Y(new_n15157));
  xnor_4 g12809(.A(new_n15157), .B(new_n15130), .Y(new_n15158));
  xor_4  g12810(.A(new_n15158), .B(new_n7313), .Y(new_n15159));
  xor_4  g12811(.A(pi687), .B(new_n8796), .Y(new_n15160));
  not_8  g12812(.A(new_n15160), .Y(new_n15161));
  nor_5  g12813(.A(pi123), .B(new_n2855), .Y(new_n15162));
  nand_5 g12814(.A(pi811), .B(new_n2859), .Y(new_n15163));
  xor_4  g12815(.A(pi811), .B(new_n2859), .Y(new_n15164));
  nand_5 g12816(.A(pi804), .B(new_n2862), .Y(new_n15165));
  nand_5 g12817(.A(pi573), .B(new_n9488), .Y(new_n15166));
  nand_5 g12818(.A(pi273), .B(new_n2883), .Y(new_n15167));
  nand_5 g12819(.A(new_n14052), .B(new_n14051), .Y(new_n15168));
  nand_5 g12820(.A(new_n15168), .B(new_n15167), .Y(new_n15169));
  xor_4  g12821(.A(pi573), .B(pi172), .Y(new_n15170));
  not_8  g12822(.A(new_n15170), .Y(new_n15171));
  nand_5 g12823(.A(new_n15171), .B(new_n15169), .Y(new_n15172));
  nand_5 g12824(.A(new_n15172), .B(new_n15166), .Y(new_n15173));
  xor_4  g12825(.A(pi804), .B(new_n2862), .Y(new_n15174));
  nand_5 g12826(.A(new_n15174), .B(new_n15173), .Y(new_n15175));
  nand_5 g12827(.A(new_n15175), .B(new_n15165), .Y(new_n15176));
  nand_5 g12828(.A(new_n15176), .B(new_n15164), .Y(new_n15177));
  nand_5 g12829(.A(new_n15177), .B(new_n15163), .Y(new_n15178));
  xor_4  g12830(.A(pi123), .B(pi047), .Y(new_n15179));
  nor_5  g12831(.A(new_n15179), .B(new_n15178), .Y(new_n15180));
  nor_5  g12832(.A(new_n15180), .B(new_n15162), .Y(new_n15181));
  xor_4  g12833(.A(new_n15181), .B(new_n15161), .Y(new_n15182));
  not_8  g12834(.A(new_n15182), .Y(new_n15183));
  xor_4  g12835(.A(new_n15183), .B(new_n15159), .Y(new_n15184));
  not_8  g12836(.A(new_n15184), .Y(new_n15185));
  xor_4  g12837(.A(new_n15155), .B(new_n15133), .Y(new_n15186));
  not_8  g12838(.A(new_n15186), .Y(new_n15187));
  xor_4  g12839(.A(new_n15179), .B(new_n15178), .Y(new_n15188));
  nor_5  g12840(.A(new_n15188), .B(new_n15187), .Y(new_n15189));
  xor_4  g12841(.A(new_n15188), .B(new_n15186), .Y(new_n15190));
  xor_4  g12842(.A(new_n15153), .B(new_n7325), .Y(new_n15191));
  xor_4  g12843(.A(new_n15176), .B(new_n15164), .Y(new_n15192));
  nor_5  g12844(.A(new_n15192), .B(new_n15191), .Y(new_n15193));
  xor_4  g12845(.A(new_n15192), .B(new_n15191), .Y(new_n15194));
  not_8  g12846(.A(new_n15194), .Y(new_n15195));
  xor_4  g12847(.A(new_n15148), .B(new_n7329), .Y(new_n15196));
  not_8  g12848(.A(new_n15196), .Y(new_n15197));
  xnor_4 g12849(.A(new_n15174), .B(new_n15173), .Y(new_n15198));
  nor_5  g12850(.A(new_n15198), .B(new_n15197), .Y(new_n15199));
  xor_4  g12851(.A(new_n15198), .B(new_n15196), .Y(new_n15200));
  xor_4  g12852(.A(new_n15144), .B(new_n7332), .Y(new_n15201));
  xor_4  g12853(.A(new_n15170), .B(new_n15169), .Y(new_n15202));
  nand_5 g12854(.A(new_n15202), .B(new_n15201), .Y(new_n15203));
  or_6   g12855(.A(new_n14053), .B(new_n14043), .Y(new_n15204));
  nand_5 g12856(.A(new_n14074), .B(new_n14054), .Y(new_n15205));
  nand_5 g12857(.A(new_n15205), .B(new_n15204), .Y(new_n15206));
  not_8  g12858(.A(new_n15201), .Y(new_n15207));
  xor_4  g12859(.A(new_n15202), .B(new_n15207), .Y(new_n15208));
  not_8  g12860(.A(new_n15208), .Y(new_n15209));
  nand_5 g12861(.A(new_n15209), .B(new_n15206), .Y(new_n15210));
  nand_5 g12862(.A(new_n15210), .B(new_n15203), .Y(new_n15211));
  nor_5  g12863(.A(new_n15211), .B(new_n15200), .Y(new_n15212));
  or_6   g12864(.A(new_n15212), .B(new_n15199), .Y(new_n15213));
  nor_5  g12865(.A(new_n15213), .B(new_n15195), .Y(new_n15214));
  or_6   g12866(.A(new_n15214), .B(new_n15193), .Y(new_n15215));
  nor_5  g12867(.A(new_n15215), .B(new_n15190), .Y(new_n15216));
  or_6   g12868(.A(new_n15216), .B(new_n15189), .Y(new_n15217));
  xor_4  g12869(.A(new_n15217), .B(new_n15185), .Y(po0138));
  xnor_4 g12870(.A(new_n14602), .B(new_n14601), .Y(po0139));
  nand_5 g12871(.A(new_n11460), .B(new_n11459), .Y(new_n15220));
  xnor_4 g12872(.A(new_n15220), .B(new_n11486), .Y(po0140));
  xnor_4 g12873(.A(new_n2541), .B(new_n2514), .Y(po0141));
  xnor_4 g12874(.A(new_n6704), .B(new_n6703), .Y(po0142));
  xor_4  g12875(.A(new_n11864), .B(new_n9066), .Y(po0143));
  xnor_4 g12876(.A(new_n6047), .B(new_n6046), .Y(po0144));
  xor_4  g12877(.A(new_n9985), .B(new_n2753), .Y(new_n15226));
  xor_4  g12878(.A(new_n15226), .B(new_n9934), .Y(po0145));
  xor_4  g12879(.A(pi343), .B(new_n4763), .Y(new_n15228));
  or_6   g12880(.A(pi599), .B(new_n9229), .Y(new_n15229));
  xor_4  g12881(.A(pi599), .B(new_n9229), .Y(new_n15230));
  nand_5 g12882(.A(pi480), .B(new_n4770), .Y(new_n15231));
  nand_5 g12883(.A(new_n7923), .B(pi000), .Y(new_n15232));
  not_8  g12884(.A(new_n15232), .Y(new_n15233));
  xor_4  g12885(.A(pi480), .B(new_n4770), .Y(new_n15234));
  nand_5 g12886(.A(new_n15234), .B(new_n15233), .Y(new_n15235));
  nand_5 g12887(.A(new_n15235), .B(new_n15231), .Y(new_n15236));
  nand_5 g12888(.A(new_n15236), .B(new_n15230), .Y(new_n15237));
  nand_5 g12889(.A(new_n15237), .B(new_n15229), .Y(new_n15238));
  xor_4  g12890(.A(new_n15238), .B(new_n15228), .Y(new_n15239));
  xor_4  g12891(.A(new_n15239), .B(new_n10802), .Y(new_n15240));
  xor_4  g12892(.A(new_n15236), .B(new_n15230), .Y(new_n15241));
  nor_5  g12893(.A(new_n15241), .B(new_n10803), .Y(new_n15242));
  xnor_4 g12894(.A(new_n15241), .B(new_n10803), .Y(new_n15243));
  xor_4  g12895(.A(new_n15234), .B(new_n15233), .Y(new_n15244));
  xor_4  g12896(.A(pi482), .B(new_n9235), .Y(new_n15245));
  not_8  g12897(.A(new_n15245), .Y(new_n15246));
  nand_5 g12898(.A(new_n15246), .B(new_n5773), .Y(new_n15247));
  nor_5  g12899(.A(new_n15247), .B(new_n15244), .Y(new_n15248));
  not_8  g12900(.A(new_n15244), .Y(new_n15249));
  xor_4  g12901(.A(new_n15247), .B(new_n15249), .Y(new_n15250));
  nor_5  g12902(.A(new_n15250), .B(new_n5772), .Y(new_n15251));
  nor_5  g12903(.A(new_n15251), .B(new_n15248), .Y(new_n15252));
  nor_5  g12904(.A(new_n15252), .B(new_n15243), .Y(new_n15253));
  or_6   g12905(.A(new_n15253), .B(new_n15242), .Y(new_n15254));
  xor_4  g12906(.A(new_n15254), .B(new_n15240), .Y(po0146));
  nor_5  g12907(.A(new_n5162), .B(new_n5137), .Y(new_n15256));
  xor_4  g12908(.A(new_n15256), .B(new_n5157), .Y(po0147));
  nand_5 g12909(.A(pi663), .B(pi582), .Y(new_n15258));
  xor_4  g12910(.A(pi663), .B(pi582), .Y(new_n15259));
  nor_5  g12911(.A(pi835), .B(pi404), .Y(new_n15260));
  nor_5  g12912(.A(new_n2979), .B(new_n2977), .Y(new_n15261));
  nor_5  g12913(.A(new_n15261), .B(new_n15260), .Y(new_n15262));
  nand_5 g12914(.A(new_n15262), .B(new_n15259), .Y(new_n15263));
  nand_5 g12915(.A(new_n15263), .B(new_n15258), .Y(new_n15264));
  not_8  g12916(.A(new_n15264), .Y(new_n15265));
  xor_4  g12917(.A(new_n15262), .B(new_n15259), .Y(new_n15266));
  or_6   g12918(.A(new_n2980), .B(new_n2837), .Y(new_n15267));
  not_8  g12919(.A(new_n2984), .Y(new_n15268));
  nand_5 g12920(.A(new_n13503), .B(new_n2995), .Y(new_n15269));
  nand_5 g12921(.A(new_n13504), .B(new_n2675), .Y(new_n15270));
  nand_5 g12922(.A(new_n15270), .B(new_n15269), .Y(new_n15271));
  or_6   g12923(.A(new_n15271), .B(new_n2990), .Y(new_n15272));
  xor_4  g12924(.A(new_n15271), .B(new_n2990), .Y(new_n15273));
  nand_5 g12925(.A(new_n15273), .B(pi691), .Y(new_n15274));
  nand_5 g12926(.A(new_n15274), .B(new_n15272), .Y(new_n15275));
  nor_5  g12927(.A(new_n15275), .B(new_n15268), .Y(new_n15276));
  xor_4  g12928(.A(new_n15275), .B(new_n15268), .Y(new_n15277));
  nand_5 g12929(.A(new_n15277), .B(new_n2814), .Y(new_n15278));
  not_8  g12930(.A(new_n15278), .Y(new_n15279));
  nor_5  g12931(.A(new_n15279), .B(new_n15276), .Y(new_n15280));
  xor_4  g12932(.A(new_n2980), .B(new_n2837), .Y(new_n15281));
  nand_5 g12933(.A(new_n15281), .B(new_n15280), .Y(new_n15282));
  nand_5 g12934(.A(new_n15282), .B(new_n15267), .Y(new_n15283));
  or_6   g12935(.A(new_n15283), .B(new_n15266), .Y(new_n15284));
  nand_5 g12936(.A(new_n15283), .B(new_n15266), .Y(new_n15285));
  nand_5 g12937(.A(new_n15285), .B(new_n10405), .Y(new_n15286));
  nand_5 g12938(.A(new_n15286), .B(new_n15284), .Y(new_n15287));
  nor_5  g12939(.A(new_n15287), .B(new_n15265), .Y(new_n15288));
  xor_4  g12940(.A(new_n15277), .B(pi233), .Y(new_n15289));
  nor_5  g12941(.A(new_n15289), .B(new_n11566), .Y(new_n15290));
  nand_5 g12942(.A(new_n13505), .B(new_n12180), .Y(new_n15291));
  or_6   g12943(.A(new_n13532), .B(new_n13506), .Y(new_n15292));
  nand_5 g12944(.A(new_n15292), .B(new_n15291), .Y(new_n15293));
  nor_5  g12945(.A(new_n15293), .B(new_n12143), .Y(new_n15294));
  xor_4  g12946(.A(new_n15273), .B(pi691), .Y(new_n15295));
  xor_4  g12947(.A(new_n15293), .B(new_n11579), .Y(new_n15296));
  nor_5  g12948(.A(new_n15296), .B(new_n15295), .Y(new_n15297));
  nor_5  g12949(.A(new_n15297), .B(new_n15294), .Y(new_n15298));
  xor_4  g12950(.A(new_n15289), .B(new_n11565), .Y(new_n15299));
  nor_5  g12951(.A(new_n15299), .B(new_n15298), .Y(new_n15300));
  nor_5  g12952(.A(new_n15300), .B(new_n15290), .Y(new_n15301));
  xor_4  g12953(.A(new_n15281), .B(new_n15280), .Y(new_n15302));
  nand_5 g12954(.A(new_n15302), .B(new_n15301), .Y(new_n15303));
  xnor_4 g12955(.A(new_n15302), .B(new_n15301), .Y(new_n15304));
  or_6   g12956(.A(new_n15304), .B(new_n11587), .Y(new_n15305));
  nand_5 g12957(.A(new_n15305), .B(new_n15303), .Y(new_n15306));
  nand_5 g12958(.A(new_n15284), .B(new_n15285), .Y(new_n15307));
  xor_4  g12959(.A(new_n15307), .B(pi095), .Y(new_n15308));
  not_8  g12960(.A(new_n15308), .Y(new_n15309));
  nand_5 g12961(.A(new_n15309), .B(new_n15306), .Y(new_n15310));
  xor_4  g12962(.A(new_n15308), .B(new_n15306), .Y(new_n15311));
  or_6   g12963(.A(new_n15311), .B(new_n11563), .Y(new_n15312));
  nand_5 g12964(.A(new_n15312), .B(new_n15310), .Y(new_n15313));
  nor_5  g12965(.A(new_n15313), .B(new_n11561), .Y(new_n15314));
  xor_4  g12966(.A(new_n15313), .B(new_n11562), .Y(new_n15315));
  not_8  g12967(.A(new_n15315), .Y(new_n15316));
  xor_4  g12968(.A(new_n15287), .B(new_n15264), .Y(new_n15317));
  nand_5 g12969(.A(new_n15317), .B(new_n15316), .Y(new_n15318));
  xor_4  g12970(.A(new_n15318), .B(new_n11558), .Y(new_n15319));
  nor_5  g12971(.A(new_n15319), .B(new_n15314), .Y(new_n15320));
  xor_4  g12972(.A(new_n15320), .B(new_n15288), .Y(po0148));
  xnor_4 g12973(.A(new_n12186), .B(new_n12142), .Y(po0149));
  xnor_4 g12974(.A(new_n14895), .B(new_n14894), .Y(po0151));
  xnor_4 g12975(.A(new_n11336), .B(new_n11323), .Y(po0152));
  xor_4  g12976(.A(new_n11537), .B(pi286), .Y(new_n15325));
  nand_5 g12977(.A(pi759), .B(new_n8724), .Y(new_n15326));
  xor_4  g12978(.A(pi759), .B(new_n8724), .Y(new_n15327));
  nand_5 g12979(.A(pi815), .B(new_n8727), .Y(new_n15328));
  xor_4  g12980(.A(pi815), .B(new_n8727), .Y(new_n15329));
  nand_5 g12981(.A(new_n9659), .B(pi496), .Y(new_n15330));
  xor_4  g12982(.A(pi535), .B(new_n2651), .Y(new_n15331));
  nand_5 g12983(.A(new_n2590), .B(pi283), .Y(new_n15332));
  xor_4  g12984(.A(new_n2590), .B(pi283), .Y(new_n15333));
  nand_5 g12985(.A(pi502), .B(new_n2638), .Y(new_n15334));
  nand_5 g12986(.A(pi725), .B(new_n2752), .Y(new_n15335));
  not_8  g12987(.A(new_n15335), .Y(new_n15336));
  xor_4  g12988(.A(pi502), .B(new_n2638), .Y(new_n15337));
  nand_5 g12989(.A(new_n15337), .B(new_n15336), .Y(new_n15338));
  nand_5 g12990(.A(new_n15338), .B(new_n15334), .Y(new_n15339));
  nand_5 g12991(.A(new_n15339), .B(new_n15333), .Y(new_n15340));
  nand_5 g12992(.A(new_n15340), .B(new_n15332), .Y(new_n15341));
  nand_5 g12993(.A(new_n15341), .B(new_n15331), .Y(new_n15342));
  nand_5 g12994(.A(new_n15342), .B(new_n15330), .Y(new_n15343));
  nand_5 g12995(.A(new_n15343), .B(new_n15329), .Y(new_n15344));
  nand_5 g12996(.A(new_n15344), .B(new_n15328), .Y(new_n15345));
  nand_5 g12997(.A(new_n15345), .B(new_n15327), .Y(new_n15346));
  nand_5 g12998(.A(new_n15346), .B(new_n15326), .Y(new_n15347));
  xor_4  g12999(.A(new_n15347), .B(new_n15325), .Y(new_n15348));
  nand_5 g13000(.A(pi723), .B(new_n11104), .Y(new_n15349));
  not_8  g13001(.A(new_n9897), .Y(new_n15350));
  nand_5 g13002(.A(pi206), .B(new_n8015), .Y(new_n15351));
  nand_5 g13003(.A(new_n13736), .B(new_n9900), .Y(new_n15352));
  nand_5 g13004(.A(new_n15352), .B(new_n15351), .Y(new_n15353));
  nand_5 g13005(.A(new_n15353), .B(new_n15350), .Y(new_n15354));
  nand_5 g13006(.A(new_n15354), .B(new_n15349), .Y(new_n15355));
  xor_4  g13007(.A(new_n15355), .B(new_n9895), .Y(new_n15356));
  nand_5 g13008(.A(new_n15356), .B(new_n15137), .Y(new_n15357));
  xor_4  g13009(.A(new_n15356), .B(new_n15137), .Y(new_n15358));
  xor_4  g13010(.A(new_n15353), .B(new_n15350), .Y(new_n15359));
  not_8  g13011(.A(new_n15359), .Y(new_n15360));
  nand_5 g13012(.A(new_n15360), .B(new_n15139), .Y(new_n15361));
  or_6   g13013(.A(new_n13749), .B(new_n13737), .Y(new_n15362));
  nand_5 g13014(.A(new_n13778), .B(new_n13750), .Y(new_n15363));
  nand_5 g13015(.A(new_n15363), .B(new_n15362), .Y(new_n15364));
  xor_4  g13016(.A(new_n15359), .B(new_n15139), .Y(new_n15365));
  or_6   g13017(.A(new_n15365), .B(new_n15364), .Y(new_n15366));
  nand_5 g13018(.A(new_n15366), .B(new_n15361), .Y(new_n15367));
  nand_5 g13019(.A(new_n15367), .B(new_n15358), .Y(new_n15368));
  nand_5 g13020(.A(new_n15368), .B(new_n15357), .Y(new_n15369));
  nand_5 g13021(.A(new_n15355), .B(new_n9894), .Y(new_n15370));
  nand_5 g13022(.A(new_n15370), .B(new_n9893), .Y(new_n15371));
  xor_4  g13023(.A(new_n15371), .B(new_n9890), .Y(new_n15372));
  xor_4  g13024(.A(new_n15372), .B(new_n15134), .Y(new_n15373));
  xor_4  g13025(.A(new_n15373), .B(new_n15369), .Y(new_n15374));
  nand_5 g13026(.A(new_n15374), .B(new_n15348), .Y(new_n15375));
  xor_4  g13027(.A(new_n15345), .B(new_n15327), .Y(new_n15376));
  xnor_4 g13028(.A(new_n15367), .B(new_n15358), .Y(new_n15377));
  nor_5  g13029(.A(new_n15377), .B(new_n15376), .Y(new_n15378));
  xor_4  g13030(.A(new_n15377), .B(new_n15376), .Y(new_n15379));
  not_8  g13031(.A(new_n15379), .Y(new_n15380));
  xor_4  g13032(.A(new_n15343), .B(new_n15329), .Y(new_n15381));
  xnor_4 g13033(.A(new_n15365), .B(new_n15364), .Y(new_n15382));
  nand_5 g13034(.A(new_n15382), .B(new_n15381), .Y(new_n15383));
  xor_4  g13035(.A(new_n15341), .B(new_n15331), .Y(new_n15384));
  or_6   g13036(.A(new_n15384), .B(new_n13779), .Y(new_n15385));
  xor_4  g13037(.A(new_n15384), .B(new_n13779), .Y(new_n15386));
  xor_4  g13038(.A(new_n15339), .B(new_n15333), .Y(new_n15387));
  nand_5 g13039(.A(new_n15387), .B(new_n13793), .Y(new_n15388));
  not_8  g13040(.A(new_n15387), .Y(new_n15389));
  xor_4  g13041(.A(new_n15389), .B(new_n13793), .Y(new_n15390));
  xor_4  g13042(.A(new_n15337), .B(new_n15336), .Y(new_n15391));
  not_8  g13043(.A(new_n15391), .Y(new_n15392));
  nor_5  g13044(.A(new_n13799), .B(new_n2753), .Y(new_n15393));
  nor_5  g13045(.A(new_n15393), .B(new_n15392), .Y(new_n15394));
  xor_4  g13046(.A(new_n15393), .B(new_n15391), .Y(new_n15395));
  nor_5  g13047(.A(new_n15395), .B(new_n13808), .Y(new_n15396));
  nor_5  g13048(.A(new_n15396), .B(new_n15394), .Y(new_n15397));
  or_6   g13049(.A(new_n15397), .B(new_n15390), .Y(new_n15398));
  nand_5 g13050(.A(new_n15398), .B(new_n15388), .Y(new_n15399));
  not_8  g13051(.A(new_n15399), .Y(new_n15400));
  nand_5 g13052(.A(new_n15400), .B(new_n15386), .Y(new_n15401));
  nand_5 g13053(.A(new_n15401), .B(new_n15385), .Y(new_n15402));
  not_8  g13054(.A(new_n15381), .Y(new_n15403));
  xor_4  g13055(.A(new_n15382), .B(new_n15403), .Y(new_n15404));
  or_6   g13056(.A(new_n15404), .B(new_n15402), .Y(new_n15405));
  nand_5 g13057(.A(new_n15405), .B(new_n15383), .Y(new_n15406));
  nor_5  g13058(.A(new_n15406), .B(new_n15380), .Y(new_n15407));
  or_6   g13059(.A(new_n15407), .B(new_n15378), .Y(new_n15408));
  xnor_4 g13060(.A(new_n15374), .B(new_n15348), .Y(new_n15409));
  or_6   g13061(.A(new_n15409), .B(new_n15408), .Y(new_n15410));
  nand_5 g13062(.A(new_n15410), .B(new_n15375), .Y(new_n15411));
  not_8  g13063(.A(new_n15411), .Y(new_n15412));
  not_8  g13064(.A(pi551), .Y(new_n15413));
  xor_4  g13065(.A(pi581), .B(new_n15413), .Y(new_n15414));
  nand_5 g13066(.A(new_n11537), .B(pi286), .Y(new_n15415));
  nand_5 g13067(.A(new_n15347), .B(new_n15325), .Y(new_n15416));
  nand_5 g13068(.A(new_n15416), .B(new_n15415), .Y(new_n15417));
  xor_4  g13069(.A(new_n15417), .B(new_n15414), .Y(new_n15418));
  not_8  g13070(.A(new_n15372), .Y(new_n15419));
  nand_5 g13071(.A(new_n15419), .B(new_n15134), .Y(new_n15420));
  or_6   g13072(.A(new_n15373), .B(new_n15369), .Y(new_n15421));
  nand_5 g13073(.A(new_n15421), .B(new_n15420), .Y(new_n15422));
  nor_5  g13074(.A(new_n8008), .B(pi186), .Y(new_n15423));
  nor_5  g13075(.A(new_n15371), .B(new_n9890), .Y(new_n15424));
  nor_5  g13076(.A(new_n15424), .B(new_n15423), .Y(new_n15425));
  xor_4  g13077(.A(new_n15425), .B(new_n10084), .Y(new_n15426));
  not_8  g13078(.A(new_n15426), .Y(new_n15427));
  xor_4  g13079(.A(new_n15427), .B(new_n15131), .Y(new_n15428));
  xnor_4 g13080(.A(new_n15428), .B(new_n15422), .Y(new_n15429));
  xor_4  g13081(.A(new_n15429), .B(new_n15418), .Y(new_n15430));
  xor_4  g13082(.A(new_n15430), .B(new_n15412), .Y(po0153));
  xnor_4 g13083(.A(new_n12374), .B(new_n12373), .Y(po0154));
  not_8  g13084(.A(new_n5042), .Y(new_n15433));
  xor_4  g13085(.A(new_n9575), .B(pi733), .Y(new_n15434));
  nand_5 g13086(.A(new_n14514), .B(pi654), .Y(new_n15435));
  not_8  g13087(.A(new_n5059), .Y(new_n15436));
  xor_4  g13088(.A(new_n8609), .B(new_n5043), .Y(new_n15437));
  nand_5 g13089(.A(new_n15437), .B(new_n15436), .Y(new_n15438));
  nand_5 g13090(.A(new_n15438), .B(new_n15435), .Y(new_n15439));
  nand_5 g13091(.A(new_n15439), .B(new_n15434), .Y(new_n15440));
  xor_4  g13092(.A(new_n15439), .B(new_n15434), .Y(new_n15441));
  nand_5 g13093(.A(new_n15441), .B(new_n5068), .Y(new_n15442));
  nand_5 g13094(.A(new_n15442), .B(new_n15440), .Y(new_n15443));
  nor_5  g13095(.A(new_n15443), .B(new_n15433), .Y(new_n15444));
  xor_4  g13096(.A(new_n15443), .B(new_n5042), .Y(new_n15445));
  nand_5 g13097(.A(new_n9575), .B(pi733), .Y(new_n15446));
  xor_4  g13098(.A(new_n15446), .B(pi127), .Y(new_n15447));
  xor_4  g13099(.A(new_n15447), .B(new_n9573), .Y(new_n15448));
  nor_5  g13100(.A(new_n15448), .B(new_n15445), .Y(new_n15449));
  or_6   g13101(.A(new_n15449), .B(new_n15444), .Y(new_n15450));
  nor_5  g13102(.A(new_n15446), .B(new_n5131), .Y(new_n15451));
  nor_5  g13103(.A(new_n15447), .B(new_n9573), .Y(new_n15452));
  or_6   g13104(.A(new_n15452), .B(new_n15451), .Y(new_n15453));
  xor_4  g13105(.A(new_n9597), .B(new_n5128), .Y(new_n15454));
  xor_4  g13106(.A(new_n15454), .B(new_n15453), .Y(new_n15455));
  nand_5 g13107(.A(new_n15455), .B(new_n15450), .Y(new_n15456));
  xor_4  g13108(.A(pi831), .B(pi414), .Y(new_n15457));
  nor_5  g13109(.A(pi550), .B(pi501), .Y(new_n15458));
  not_8  g13110(.A(new_n5022), .Y(new_n15459));
  nor_5  g13111(.A(new_n5029), .B(new_n15459), .Y(new_n15460));
  nor_5  g13112(.A(new_n15460), .B(new_n15458), .Y(new_n15461));
  xor_4  g13113(.A(new_n15461), .B(new_n15457), .Y(new_n15462));
  not_8  g13114(.A(new_n15462), .Y(new_n15463));
  or_6   g13115(.A(new_n5040), .B(new_n5030), .Y(new_n15464));
  nand_5 g13116(.A(new_n5041), .B(pi276), .Y(new_n15465));
  nand_5 g13117(.A(new_n15465), .B(new_n15464), .Y(new_n15466));
  xor_4  g13118(.A(new_n15466), .B(pi228), .Y(new_n15467));
  xor_4  g13119(.A(new_n15467), .B(new_n15463), .Y(new_n15468));
  xnor_4 g13120(.A(new_n15455), .B(new_n15450), .Y(new_n15469));
  or_6   g13121(.A(new_n15469), .B(new_n15468), .Y(new_n15470));
  nand_5 g13122(.A(new_n15470), .B(new_n15456), .Y(new_n15471));
  xor_4  g13123(.A(pi662), .B(pi171), .Y(new_n15472));
  nand_5 g13124(.A(pi831), .B(pi414), .Y(new_n15473));
  nand_5 g13125(.A(new_n15461), .B(new_n15457), .Y(new_n15474));
  nand_5 g13126(.A(new_n15474), .B(new_n15473), .Y(new_n15475));
  xor_4  g13127(.A(new_n15475), .B(new_n15472), .Y(new_n15476));
  nand_5 g13128(.A(new_n15466), .B(pi228), .Y(new_n15477));
  nand_5 g13129(.A(new_n15467), .B(new_n15463), .Y(new_n15478));
  nand_5 g13130(.A(new_n15478), .B(new_n15477), .Y(new_n15479));
  xor_4  g13131(.A(new_n15479), .B(new_n15476), .Y(new_n15480));
  xor_4  g13132(.A(new_n15480), .B(new_n8591), .Y(new_n15481));
  nand_5 g13133(.A(new_n14509), .B(new_n5128), .Y(new_n15482));
  or_6   g13134(.A(new_n15454), .B(new_n15453), .Y(new_n15483));
  nand_5 g13135(.A(new_n15483), .B(new_n15482), .Y(new_n15484));
  xor_4  g13136(.A(new_n15484), .B(new_n14505), .Y(new_n15485));
  xor_4  g13137(.A(new_n15485), .B(pi653), .Y(new_n15486));
  or_6   g13138(.A(new_n15486), .B(new_n15481), .Y(new_n15487));
  nand_5 g13139(.A(new_n15486), .B(new_n15481), .Y(new_n15488));
  nand_5 g13140(.A(new_n15488), .B(new_n15487), .Y(new_n15489));
  xor_4  g13141(.A(new_n15489), .B(new_n15471), .Y(po0155));
  not_8  g13142(.A(pi101), .Y(new_n15491));
  not_8  g13143(.A(new_n10857), .Y(new_n15492));
  not_8  g13144(.A(new_n10863), .Y(new_n15493));
  nand_5 g13145(.A(new_n15493), .B(pi389), .Y(new_n15494));
  nand_5 g13146(.A(new_n13545), .B(new_n13543), .Y(new_n15495));
  nand_5 g13147(.A(new_n15495), .B(new_n15494), .Y(new_n15496));
  nand_5 g13148(.A(new_n15496), .B(pi693), .Y(new_n15497));
  xor_4  g13149(.A(new_n15496), .B(pi693), .Y(new_n15498));
  nand_5 g13150(.A(new_n15498), .B(new_n10858), .Y(new_n15499));
  nand_5 g13151(.A(new_n15499), .B(new_n15497), .Y(new_n15500));
  or_6   g13152(.A(new_n15500), .B(pi591), .Y(new_n15501));
  xor_4  g13153(.A(new_n15500), .B(pi591), .Y(new_n15502));
  nand_5 g13154(.A(new_n15502), .B(new_n10873), .Y(new_n15503));
  nand_5 g13155(.A(new_n15503), .B(new_n15501), .Y(new_n15504));
  xor_4  g13156(.A(new_n15504), .B(new_n15492), .Y(new_n15505));
  xor_4  g13157(.A(new_n15505), .B(new_n15491), .Y(new_n15506));
  not_8  g13158(.A(new_n15506), .Y(new_n15507));
  xor_4  g13159(.A(new_n15502), .B(new_n10873), .Y(new_n15508));
  not_8  g13160(.A(new_n15508), .Y(new_n15509));
  or_6   g13161(.A(new_n13546), .B(new_n13542), .Y(new_n15510));
  nand_5 g13162(.A(new_n13547), .B(new_n13535), .Y(new_n15511));
  nand_5 g13163(.A(new_n15511), .B(new_n15510), .Y(new_n15512));
  nand_5 g13164(.A(new_n15512), .B(new_n10016), .Y(new_n15513));
  not_8  g13165(.A(new_n15513), .Y(new_n15514));
  nor_5  g13166(.A(new_n15512), .B(new_n10016), .Y(new_n15515));
  xor_4  g13167(.A(new_n15498), .B(new_n10859), .Y(new_n15516));
  not_8  g13168(.A(new_n15516), .Y(new_n15517));
  nor_5  g13169(.A(new_n15517), .B(new_n15515), .Y(new_n15518));
  nor_5  g13170(.A(new_n15518), .B(new_n15514), .Y(new_n15519));
  nor_5  g13171(.A(new_n15519), .B(new_n15509), .Y(new_n15520));
  xor_4  g13172(.A(new_n15519), .B(new_n15508), .Y(new_n15521));
  nor_5  g13173(.A(new_n15521), .B(new_n10023), .Y(new_n15522));
  or_6   g13174(.A(new_n15522), .B(new_n15520), .Y(new_n15523));
  xor_4  g13175(.A(new_n15523), .B(new_n15507), .Y(new_n15524));
  xor_4  g13176(.A(new_n15524), .B(new_n10001), .Y(po0156));
  xor_4  g13177(.A(new_n13528), .B(new_n12153), .Y(po0157));
  nand_5 g13178(.A(new_n10650), .B(new_n8103), .Y(new_n15527));
  nand_5 g13179(.A(new_n10651), .B(new_n11096), .Y(new_n15528));
  nand_5 g13180(.A(new_n15528), .B(new_n15527), .Y(new_n15529));
  nor_5  g13181(.A(new_n15529), .B(new_n10972), .Y(new_n15530));
  nor_5  g13182(.A(new_n15530), .B(pi028), .Y(new_n15531));
  nand_5 g13183(.A(new_n15529), .B(new_n10972), .Y(new_n15532));
  not_8  g13184(.A(new_n15532), .Y(new_n15533));
  nor_5  g13185(.A(new_n15533), .B(new_n15531), .Y(new_n15534));
  nand_5 g13186(.A(new_n15534), .B(pi534), .Y(new_n15535));
  xor_4  g13187(.A(new_n15534), .B(pi534), .Y(new_n15536));
  nand_5 g13188(.A(new_n15536), .B(new_n8049), .Y(new_n15537));
  nand_5 g13189(.A(new_n15537), .B(new_n15535), .Y(new_n15538));
  xor_4  g13190(.A(new_n15538), .B(new_n8047), .Y(new_n15539));
  or_6   g13191(.A(new_n13068), .B(pi292), .Y(new_n15540));
  nand_5 g13192(.A(new_n13073), .B(pi713), .Y(new_n15541));
  not_8  g13193(.A(new_n15541), .Y(new_n15542));
  nand_5 g13194(.A(new_n15542), .B(new_n15540), .Y(new_n15543));
  nand_5 g13195(.A(new_n13068), .B(pi292), .Y(new_n15544));
  not_8  g13196(.A(new_n15544), .Y(new_n15545));
  not_8  g13197(.A(pi713), .Y(new_n15546));
  or_6   g13198(.A(new_n13074), .B(new_n15546), .Y(new_n15547));
  nand_5 g13199(.A(new_n15547), .B(new_n13072), .Y(new_n15548));
  nand_5 g13200(.A(new_n15548), .B(new_n15545), .Y(new_n15549));
  nand_5 g13201(.A(new_n15549), .B(new_n15543), .Y(new_n15550));
  not_8  g13202(.A(new_n15550), .Y(new_n15551));
  nand_5 g13203(.A(new_n13074), .B(new_n15546), .Y(new_n15552));
  not_8  g13204(.A(new_n15552), .Y(new_n15553));
  nand_5 g13205(.A(new_n15553), .B(new_n15544), .Y(new_n15554));
  not_8  g13206(.A(new_n15554), .Y(new_n15555));
  nor_5  g13207(.A(new_n15548), .B(new_n15540), .Y(new_n15556));
  nor_5  g13208(.A(new_n15556), .B(new_n15555), .Y(new_n15557));
  nand_5 g13209(.A(new_n15557), .B(new_n15551), .Y(new_n15558));
  and_6  g13210(.A(new_n15558), .B(new_n15539), .Y(new_n15559));
  xor_4  g13211(.A(new_n15536), .B(new_n8049), .Y(new_n15560));
  not_8  g13212(.A(new_n15560), .Y(new_n15561));
  nand_5 g13213(.A(new_n13081), .B(new_n10710), .Y(new_n15562));
  or_6   g13214(.A(new_n10722), .B(new_n10652), .Y(new_n15563));
  nand_5 g13215(.A(new_n15563), .B(new_n15562), .Y(new_n15564));
  nor_5  g13216(.A(new_n15533), .B(new_n15530), .Y(new_n15565));
  xor_4  g13217(.A(new_n15565), .B(new_n7257), .Y(new_n15566));
  nand_5 g13218(.A(new_n15566), .B(new_n15564), .Y(new_n15567));
  xnor_4 g13219(.A(new_n15566), .B(new_n15564), .Y(new_n15568));
  or_6   g13220(.A(new_n15568), .B(new_n13080), .Y(new_n15569));
  nand_5 g13221(.A(new_n15569), .B(new_n15567), .Y(new_n15570));
  nand_5 g13222(.A(new_n15570), .B(new_n15561), .Y(new_n15571));
  xor_4  g13223(.A(new_n15570), .B(new_n15560), .Y(new_n15572));
  or_6   g13224(.A(new_n15572), .B(new_n13077), .Y(new_n15573));
  nand_5 g13225(.A(new_n15573), .B(new_n15571), .Y(new_n15574));
  xnor_4 g13226(.A(new_n15558), .B(new_n15539), .Y(new_n15575));
  nor_5  g13227(.A(new_n15575), .B(new_n15574), .Y(new_n15576));
  nor_5  g13228(.A(new_n15576), .B(new_n15559), .Y(new_n15577));
  nand_5 g13229(.A(new_n15538), .B(new_n8047), .Y(new_n15578));
  xor_4  g13230(.A(new_n15551), .B(new_n15578), .Y(new_n15579));
  xor_4  g13231(.A(new_n15579), .B(new_n15577), .Y(po0158));
  xor_4  g13232(.A(pi440), .B(new_n10711), .Y(new_n15581));
  nand_5 g13233(.A(pi762), .B(new_n10718), .Y(new_n15582));
  xor_4  g13234(.A(pi762), .B(new_n10718), .Y(new_n15583));
  nand_5 g13235(.A(new_n10701), .B(pi165), .Y(new_n15584));
  not_8  g13236(.A(pi165), .Y(new_n15585));
  xor_4  g13237(.A(pi814), .B(new_n15585), .Y(new_n15586));
  nand_5 g13238(.A(new_n10655), .B(pi101), .Y(new_n15587));
  xor_4  g13239(.A(pi604), .B(new_n15491), .Y(new_n15588));
  nand_5 g13240(.A(pi591), .B(new_n4130), .Y(new_n15589));
  or_6   g13241(.A(new_n13790), .B(new_n13789), .Y(new_n15590));
  nand_5 g13242(.A(new_n15590), .B(new_n15589), .Y(new_n15591));
  nand_5 g13243(.A(new_n15591), .B(new_n15588), .Y(new_n15592));
  nand_5 g13244(.A(new_n15592), .B(new_n15587), .Y(new_n15593));
  nand_5 g13245(.A(new_n15593), .B(new_n15586), .Y(new_n15594));
  nand_5 g13246(.A(new_n15594), .B(new_n15584), .Y(new_n15595));
  nand_5 g13247(.A(new_n15595), .B(new_n15583), .Y(new_n15596));
  nand_5 g13248(.A(new_n15596), .B(new_n15582), .Y(new_n15597));
  xor_4  g13249(.A(new_n15597), .B(new_n15581), .Y(new_n15598));
  not_8  g13250(.A(new_n15598), .Y(new_n15599));
  xor_4  g13251(.A(new_n15599), .B(new_n15429), .Y(new_n15600));
  xor_4  g13252(.A(new_n15595), .B(new_n15583), .Y(new_n15601));
  or_6   g13253(.A(new_n15601), .B(new_n15374), .Y(new_n15602));
  xor_4  g13254(.A(new_n15593), .B(new_n15586), .Y(new_n15603));
  or_6   g13255(.A(new_n15603), .B(new_n15377), .Y(new_n15604));
  xor_4  g13256(.A(new_n15591), .B(new_n15588), .Y(new_n15605));
  or_6   g13257(.A(new_n15605), .B(new_n15382), .Y(new_n15606));
  xor_4  g13258(.A(new_n15605), .B(new_n15382), .Y(new_n15607));
  or_6   g13259(.A(new_n13791), .B(new_n13779), .Y(new_n15608));
  nand_5 g13260(.A(new_n13814), .B(new_n13792), .Y(new_n15609));
  nand_5 g13261(.A(new_n15609), .B(new_n15608), .Y(new_n15610));
  nand_5 g13262(.A(new_n15610), .B(new_n15607), .Y(new_n15611));
  nand_5 g13263(.A(new_n15611), .B(new_n15606), .Y(new_n15612));
  xor_4  g13264(.A(new_n15603), .B(new_n15377), .Y(new_n15613));
  nand_5 g13265(.A(new_n15613), .B(new_n15612), .Y(new_n15614));
  nand_5 g13266(.A(new_n15614), .B(new_n15604), .Y(new_n15615));
  xor_4  g13267(.A(new_n15601), .B(new_n15374), .Y(new_n15616));
  nand_5 g13268(.A(new_n15616), .B(new_n15615), .Y(new_n15617));
  nand_5 g13269(.A(new_n15617), .B(new_n15602), .Y(new_n15618));
  xnor_4 g13270(.A(new_n15618), .B(new_n15600), .Y(po0159));
  nor_5  g13271(.A(new_n12595), .B(pi197), .Y(new_n15620));
  nand_5 g13272(.A(new_n6373), .B(pi170), .Y(new_n15621));
  not_8  g13273(.A(new_n15621), .Y(new_n15622));
  nand_5 g13274(.A(new_n15622), .B(new_n15620), .Y(new_n15623));
  nand_5 g13275(.A(new_n12609), .B(new_n12577), .Y(new_n15624));
  nand_5 g13276(.A(new_n15624), .B(new_n4088), .Y(new_n15625));
  not_8  g13277(.A(new_n15624), .Y(new_n15626));
  nand_5 g13278(.A(new_n4088), .B(pi284), .Y(new_n15627));
  nand_5 g13279(.A(pi307), .B(new_n6442), .Y(new_n15628));
  and_6  g13280(.A(new_n15628), .B(new_n15627), .Y(new_n15629));
  nor_5  g13281(.A(new_n15629), .B(new_n15626), .Y(new_n15630));
  xor_4  g13282(.A(new_n15630), .B(new_n12579), .Y(new_n15631));
  nand_5 g13283(.A(new_n15631), .B(new_n15625), .Y(new_n15632));
  or_6   g13284(.A(new_n15631), .B(new_n4086), .Y(new_n15633));
  nand_5 g13285(.A(new_n15633), .B(new_n15632), .Y(new_n15634));
  nand_5 g13286(.A(new_n15634), .B(new_n12606), .Y(new_n15635));
  xor_4  g13287(.A(new_n15634), .B(new_n12607), .Y(new_n15636));
  or_6   g13288(.A(new_n15636), .B(new_n12096), .Y(new_n15637));
  nand_5 g13289(.A(new_n15637), .B(new_n15635), .Y(new_n15638));
  nand_5 g13290(.A(new_n15638), .B(new_n12605), .Y(new_n15639));
  not_8  g13291(.A(new_n15639), .Y(new_n15640));
  nor_5  g13292(.A(new_n15638), .B(new_n12605), .Y(new_n15641));
  nor_5  g13293(.A(new_n15641), .B(new_n8875), .Y(new_n15642));
  nor_5  g13294(.A(new_n15642), .B(new_n15640), .Y(new_n15643));
  nand_5 g13295(.A(new_n15643), .B(new_n12604), .Y(new_n15644));
  xor_4  g13296(.A(new_n15643), .B(new_n12604), .Y(new_n15645));
  nand_5 g13297(.A(new_n15645), .B(new_n6165), .Y(new_n15646));
  nand_5 g13298(.A(new_n15646), .B(new_n15644), .Y(new_n15647));
  or_6   g13299(.A(new_n15647), .B(new_n12638), .Y(new_n15648));
  nand_5 g13300(.A(new_n15647), .B(new_n12638), .Y(new_n15649));
  nand_5 g13301(.A(new_n15649), .B(pi726), .Y(new_n15650));
  nand_5 g13302(.A(new_n15650), .B(new_n15648), .Y(new_n15651));
  nand_5 g13303(.A(new_n15651), .B(pi578), .Y(new_n15652));
  xor_4  g13304(.A(new_n15651), .B(new_n8868), .Y(new_n15653));
  or_6   g13305(.A(new_n15653), .B(new_n12646), .Y(new_n15654));
  nand_5 g13306(.A(new_n15654), .B(new_n15652), .Y(new_n15655));
  nand_5 g13307(.A(new_n15655), .B(new_n12653), .Y(new_n15656));
  not_8  g13308(.A(new_n15656), .Y(new_n15657));
  nor_5  g13309(.A(new_n15655), .B(new_n12653), .Y(new_n15658));
  nor_5  g13310(.A(new_n15658), .B(new_n8865), .Y(new_n15659));
  nor_5  g13311(.A(new_n15659), .B(new_n15657), .Y(new_n15660));
  not_8  g13312(.A(new_n15660), .Y(new_n15661));
  nand_5 g13313(.A(new_n15661), .B(new_n12659), .Y(new_n15662));
  xor_4  g13314(.A(new_n15660), .B(new_n12659), .Y(new_n15663));
  or_6   g13315(.A(new_n15663), .B(new_n6307), .Y(new_n15664));
  nand_5 g13316(.A(new_n15664), .B(new_n15662), .Y(new_n15665));
  not_8  g13317(.A(new_n15665), .Y(new_n15666));
  nand_5 g13318(.A(new_n15666), .B(new_n12600), .Y(new_n15667));
  nand_5 g13319(.A(pi335), .B(new_n12597), .Y(new_n15668));
  nand_5 g13320(.A(new_n15668), .B(new_n15621), .Y(new_n15669));
  not_8  g13321(.A(new_n15669), .Y(new_n15670));
  xor_4  g13322(.A(new_n15670), .B(new_n12598), .Y(new_n15671));
  not_8  g13323(.A(new_n15671), .Y(new_n15672));
  nor_5  g13324(.A(new_n15666), .B(new_n12600), .Y(new_n15673));
  nor_5  g13325(.A(new_n15673), .B(new_n15672), .Y(new_n15674));
  nand_5 g13326(.A(new_n15674), .B(new_n15667), .Y(new_n15675));
  nand_5 g13327(.A(new_n15675), .B(new_n15623), .Y(new_n15676));
  nor_5  g13328(.A(new_n15676), .B(new_n12600), .Y(new_n15677));
  not_8  g13329(.A(new_n15677), .Y(new_n15678));
  nor_5  g13330(.A(pi581), .B(new_n15413), .Y(new_n15679));
  not_8  g13331(.A(new_n15414), .Y(new_n15680));
  nor_5  g13332(.A(new_n15417), .B(new_n15680), .Y(new_n15681));
  nor_5  g13333(.A(new_n15681), .B(new_n15679), .Y(new_n15682));
  xor_4  g13334(.A(pi592), .B(pi463), .Y(new_n15683));
  xor_4  g13335(.A(new_n15683), .B(new_n15682), .Y(new_n15684));
  not_8  g13336(.A(new_n15684), .Y(new_n15685));
  not_8  g13337(.A(new_n15418), .Y(new_n15686));
  not_8  g13338(.A(new_n15376), .Y(new_n15687));
  not_8  g13339(.A(new_n15384), .Y(new_n15688));
  nand_5 g13340(.A(new_n2753), .B(pi156), .Y(new_n15689));
  or_6   g13341(.A(new_n15689), .B(new_n6440), .Y(new_n15690));
  xor_4  g13342(.A(new_n15689), .B(new_n6440), .Y(new_n15691));
  nand_5 g13343(.A(new_n15691), .B(new_n15391), .Y(new_n15692));
  nand_5 g13344(.A(new_n15692), .B(new_n15690), .Y(new_n15693));
  or_6   g13345(.A(new_n15693), .B(new_n15387), .Y(new_n15694));
  nand_5 g13346(.A(new_n15693), .B(new_n15387), .Y(new_n15695));
  nand_5 g13347(.A(new_n15695), .B(new_n6437), .Y(new_n15696));
  nand_5 g13348(.A(new_n15696), .B(new_n15694), .Y(new_n15697));
  nand_5 g13349(.A(new_n15697), .B(new_n15688), .Y(new_n15698));
  or_6   g13350(.A(new_n15697), .B(new_n15688), .Y(new_n15699));
  nand_5 g13351(.A(new_n15699), .B(new_n12436), .Y(new_n15700));
  nand_5 g13352(.A(new_n15700), .B(new_n15698), .Y(new_n15701));
  nand_5 g13353(.A(new_n15701), .B(new_n15403), .Y(new_n15702));
  or_6   g13354(.A(new_n15701), .B(new_n15403), .Y(new_n15703));
  nand_5 g13355(.A(new_n15703), .B(new_n12444), .Y(new_n15704));
  nand_5 g13356(.A(new_n15704), .B(new_n15702), .Y(new_n15705));
  or_6   g13357(.A(new_n15705), .B(new_n15687), .Y(new_n15706));
  nand_5 g13358(.A(new_n15705), .B(new_n15687), .Y(new_n15707));
  nand_5 g13359(.A(new_n15707), .B(pi030), .Y(new_n15708));
  nand_5 g13360(.A(new_n15708), .B(new_n15706), .Y(new_n15709));
  or_6   g13361(.A(new_n15709), .B(new_n15348), .Y(new_n15710));
  nand_5 g13362(.A(new_n15709), .B(new_n15348), .Y(new_n15711));
  nand_5 g13363(.A(new_n15711), .B(new_n12415), .Y(new_n15712));
  nand_5 g13364(.A(new_n15712), .B(new_n15710), .Y(new_n15713));
  or_6   g13365(.A(new_n15713), .B(new_n15686), .Y(new_n15714));
  nand_5 g13366(.A(new_n15713), .B(new_n15686), .Y(new_n15715));
  nand_5 g13367(.A(new_n15715), .B(pi119), .Y(new_n15716));
  nand_5 g13368(.A(new_n15716), .B(new_n15714), .Y(new_n15717));
  or_6   g13369(.A(new_n15717), .B(new_n15685), .Y(new_n15718));
  nand_5 g13370(.A(new_n15717), .B(new_n15685), .Y(new_n15719));
  nand_5 g13371(.A(new_n15719), .B(new_n12535), .Y(new_n15720));
  nand_5 g13372(.A(new_n15720), .B(new_n15718), .Y(new_n15721));
  nand_5 g13373(.A(pi592), .B(new_n2614), .Y(new_n15722));
  not_8  g13374(.A(new_n15722), .Y(new_n15723));
  nor_5  g13375(.A(new_n15683), .B(new_n15682), .Y(new_n15724));
  nor_5  g13376(.A(new_n15724), .B(new_n15723), .Y(new_n15725));
  not_8  g13377(.A(new_n15725), .Y(new_n15726));
  nand_5 g13378(.A(pi778), .B(new_n2608), .Y(new_n15727));
  nand_5 g13379(.A(new_n2613), .B(pi610), .Y(new_n15728));
  and_6  g13380(.A(new_n15728), .B(new_n15727), .Y(new_n15729));
  xor_4  g13381(.A(new_n15729), .B(new_n15726), .Y(new_n15730));
  or_6   g13382(.A(new_n15730), .B(new_n15721), .Y(new_n15731));
  nand_5 g13383(.A(new_n15730), .B(new_n15721), .Y(new_n15732));
  nand_5 g13384(.A(new_n15732), .B(pi327), .Y(new_n15733));
  nand_5 g13385(.A(new_n15733), .B(new_n15731), .Y(new_n15734));
  nand_5 g13386(.A(new_n15727), .B(new_n15726), .Y(new_n15735));
  nand_5 g13387(.A(new_n15735), .B(new_n15728), .Y(new_n15736));
  nand_5 g13388(.A(new_n15736), .B(new_n15734), .Y(new_n15737));
  nor_5  g13389(.A(new_n15737), .B(new_n15678), .Y(new_n15738));
  and_6  g13390(.A(new_n15737), .B(new_n15678), .Y(new_n15739));
  nor_5  g13391(.A(new_n15739), .B(new_n15738), .Y(new_n15740));
  xor_4  g13392(.A(new_n15736), .B(new_n15734), .Y(new_n15741));
  not_8  g13393(.A(new_n15741), .Y(new_n15742));
  xor_4  g13394(.A(new_n15663), .B(pi247), .Y(new_n15743));
  nand_5 g13395(.A(new_n15718), .B(new_n15719), .Y(new_n15744));
  xor_4  g13396(.A(new_n15744), .B(pi070), .Y(new_n15745));
  not_8  g13397(.A(new_n15745), .Y(new_n15746));
  nand_5 g13398(.A(new_n15746), .B(new_n15743), .Y(new_n15747));
  xor_4  g13399(.A(new_n15745), .B(new_n15743), .Y(new_n15748));
  nand_5 g13400(.A(new_n15715), .B(new_n15714), .Y(new_n15749));
  xor_4  g13401(.A(new_n15749), .B(new_n12518), .Y(new_n15750));
  nor_5  g13402(.A(new_n15658), .B(new_n15657), .Y(new_n15751));
  xor_4  g13403(.A(new_n15751), .B(new_n8865), .Y(new_n15752));
  nor_5  g13404(.A(new_n15752), .B(new_n15750), .Y(new_n15753));
  not_8  g13405(.A(new_n15750), .Y(new_n15754));
  xor_4  g13406(.A(new_n15752), .B(new_n15754), .Y(new_n15755));
  and_6  g13407(.A(new_n15703), .B(new_n15702), .Y(new_n15756));
  xor_4  g13408(.A(new_n15756), .B(pi456), .Y(new_n15757));
  and_6  g13409(.A(new_n15695), .B(new_n15694), .Y(new_n15758));
  xor_4  g13410(.A(new_n15758), .B(pi188), .Y(new_n15759));
  xor_4  g13411(.A(new_n15631), .B(pi356), .Y(new_n15760));
  xor_4  g13412(.A(new_n2753), .B(pi156), .Y(new_n15761));
  xor_4  g13413(.A(new_n15624), .B(new_n4088), .Y(new_n15762));
  nor_5  g13414(.A(new_n15762), .B(new_n15761), .Y(new_n15763));
  not_8  g13415(.A(new_n15763), .Y(new_n15764));
  nand_5 g13416(.A(new_n15764), .B(new_n15760), .Y(new_n15765));
  xor_4  g13417(.A(new_n15763), .B(new_n15760), .Y(new_n15766));
  xor_4  g13418(.A(new_n15691), .B(new_n15392), .Y(new_n15767));
  or_6   g13419(.A(new_n15767), .B(new_n15766), .Y(new_n15768));
  nand_5 g13420(.A(new_n15768), .B(new_n15765), .Y(new_n15769));
  nand_5 g13421(.A(new_n15769), .B(new_n15759), .Y(new_n15770));
  not_8  g13422(.A(new_n15759), .Y(new_n15771));
  xor_4  g13423(.A(new_n15769), .B(new_n15771), .Y(new_n15772));
  xor_4  g13424(.A(new_n15636), .B(new_n12096), .Y(new_n15773));
  or_6   g13425(.A(new_n15773), .B(new_n15772), .Y(new_n15774));
  nand_5 g13426(.A(new_n15774), .B(new_n15770), .Y(new_n15775));
  nor_5  g13427(.A(new_n15641), .B(new_n15640), .Y(new_n15776));
  xor_4  g13428(.A(new_n15776), .B(new_n8875), .Y(new_n15777));
  nand_5 g13429(.A(new_n15777), .B(new_n15775), .Y(new_n15778));
  xnor_4 g13430(.A(new_n15777), .B(new_n15775), .Y(new_n15779));
  nand_5 g13431(.A(new_n15698), .B(new_n15699), .Y(new_n15780));
  xor_4  g13432(.A(new_n15780), .B(pi098), .Y(new_n15781));
  or_6   g13433(.A(new_n15781), .B(new_n15779), .Y(new_n15782));
  nand_5 g13434(.A(new_n15782), .B(new_n15778), .Y(new_n15783));
  nand_5 g13435(.A(new_n15783), .B(new_n15757), .Y(new_n15784));
  xor_4  g13436(.A(new_n15645), .B(pi644), .Y(new_n15785));
  not_8  g13437(.A(new_n15757), .Y(new_n15786));
  xor_4  g13438(.A(new_n15783), .B(new_n15786), .Y(new_n15787));
  or_6   g13439(.A(new_n15787), .B(new_n15785), .Y(new_n15788));
  nand_5 g13440(.A(new_n15788), .B(new_n15784), .Y(new_n15789));
  nand_5 g13441(.A(new_n15649), .B(new_n15648), .Y(new_n15790));
  xor_4  g13442(.A(new_n15790), .B(pi726), .Y(new_n15791));
  or_6   g13443(.A(new_n15791), .B(new_n15789), .Y(new_n15792));
  xor_4  g13444(.A(new_n15791), .B(new_n15789), .Y(new_n15793));
  nand_5 g13445(.A(new_n15707), .B(new_n15706), .Y(new_n15794));
  xor_4  g13446(.A(new_n15794), .B(pi030), .Y(new_n15795));
  nand_5 g13447(.A(new_n15795), .B(new_n15793), .Y(new_n15796));
  nand_5 g13448(.A(new_n15796), .B(new_n15792), .Y(new_n15797));
  xor_4  g13449(.A(new_n15653), .B(new_n12645), .Y(new_n15798));
  not_8  g13450(.A(new_n15798), .Y(new_n15799));
  nor_5  g13451(.A(new_n15799), .B(new_n15797), .Y(new_n15800));
  xor_4  g13452(.A(new_n15798), .B(new_n15797), .Y(new_n15801));
  nand_5 g13453(.A(new_n15711), .B(new_n15710), .Y(new_n15802));
  xor_4  g13454(.A(new_n15802), .B(pi517), .Y(new_n15803));
  nor_5  g13455(.A(new_n15803), .B(new_n15801), .Y(new_n15804));
  or_6   g13456(.A(new_n15804), .B(new_n15800), .Y(new_n15805));
  nor_5  g13457(.A(new_n15805), .B(new_n15755), .Y(new_n15806));
  or_6   g13458(.A(new_n15806), .B(new_n15753), .Y(new_n15807));
  or_6   g13459(.A(new_n15807), .B(new_n15748), .Y(new_n15808));
  nand_5 g13460(.A(new_n15808), .B(new_n15747), .Y(new_n15809));
  nand_5 g13461(.A(new_n15732), .B(new_n15731), .Y(new_n15810));
  xor_4  g13462(.A(new_n15810), .B(pi327), .Y(new_n15811));
  not_8  g13463(.A(new_n15811), .Y(new_n15812));
  nor_5  g13464(.A(new_n15812), .B(new_n15809), .Y(new_n15813));
  xor_4  g13465(.A(new_n15672), .B(new_n15665), .Y(new_n15814));
  xor_4  g13466(.A(new_n15811), .B(new_n15809), .Y(new_n15815));
  nor_5  g13467(.A(new_n15815), .B(new_n15814), .Y(new_n15816));
  or_6   g13468(.A(new_n15816), .B(new_n15813), .Y(new_n15817));
  or_6   g13469(.A(new_n15817), .B(new_n15742), .Y(new_n15818));
  nor_5  g13470(.A(new_n15668), .B(new_n12596), .Y(new_n15819));
  or_6   g13471(.A(new_n15819), .B(new_n15676), .Y(new_n15820));
  xor_4  g13472(.A(new_n15817), .B(new_n15741), .Y(new_n15821));
  or_6   g13473(.A(new_n15821), .B(new_n15820), .Y(new_n15822));
  nand_5 g13474(.A(new_n15822), .B(new_n15818), .Y(new_n15823));
  xor_4  g13475(.A(new_n15823), .B(new_n15740), .Y(po0160));
  xnor_4 g13476(.A(new_n6516), .B(new_n6488), .Y(po0161));
  xor_4  g13477(.A(new_n4637), .B(new_n4628), .Y(po0162));
  xor_4  g13478(.A(new_n12279), .B(new_n12278), .Y(po0163));
  nand_5 g13479(.A(pi219), .B(pi010), .Y(new_n15828));
  nand_5 g13480(.A(new_n5520), .B(new_n3954), .Y(new_n15829));
  nand_5 g13481(.A(pi675), .B(pi528), .Y(new_n15830));
  nand_5 g13482(.A(new_n15830), .B(new_n15829), .Y(new_n15831));
  xor_4  g13483(.A(new_n15831), .B(pi218), .Y(new_n15832));
  xor_4  g13484(.A(new_n15832), .B(new_n15828), .Y(new_n15833));
  xor_4  g13485(.A(pi219), .B(new_n2555), .Y(new_n15834));
  nand_5 g13486(.A(new_n15834), .B(pi656), .Y(new_n15835));
  nand_5 g13487(.A(new_n15835), .B(new_n13889), .Y(new_n15836));
  not_8  g13488(.A(new_n13889), .Y(new_n15837));
  or_6   g13489(.A(new_n15834), .B(pi656), .Y(new_n15838));
  nand_5 g13490(.A(new_n15838), .B(new_n15837), .Y(new_n15839));
  nand_5 g13491(.A(new_n15839), .B(new_n15836), .Y(new_n15840));
  xor_4  g13492(.A(new_n15840), .B(new_n15833), .Y(new_n15841));
  xor_4  g13493(.A(new_n15841), .B(new_n13901), .Y(po0164));
  xnor_4 g13494(.A(new_n10953), .B(new_n10916), .Y(po0165));
  xor_4  g13495(.A(pi770), .B(pi562), .Y(new_n15844));
  nor_5  g13496(.A(pi596), .B(pi387), .Y(new_n15845));
  xor_4  g13497(.A(pi596), .B(pi387), .Y(new_n15846));
  not_8  g13498(.A(new_n15846), .Y(new_n15847));
  nor_5  g13499(.A(pi416), .B(pi051), .Y(new_n15848));
  xor_4  g13500(.A(pi416), .B(new_n4084), .Y(new_n15849));
  nand_5 g13501(.A(pi680), .B(pi564), .Y(new_n15850));
  not_8  g13502(.A(new_n15850), .Y(new_n15851));
  nor_5  g13503(.A(new_n15851), .B(new_n15849), .Y(new_n15852));
  nor_5  g13504(.A(new_n15852), .B(new_n15848), .Y(new_n15853));
  nor_5  g13505(.A(new_n15853), .B(new_n15847), .Y(new_n15854));
  nor_5  g13506(.A(new_n15854), .B(new_n15845), .Y(new_n15855));
  xor_4  g13507(.A(new_n15855), .B(new_n15844), .Y(new_n15856));
  xor_4  g13508(.A(new_n15850), .B(new_n15849), .Y(new_n15857));
  not_8  g13509(.A(new_n15857), .Y(new_n15858));
  xor_4  g13510(.A(pi680), .B(pi564), .Y(new_n15859));
  nand_5 g13511(.A(pi745), .B(pi499), .Y(new_n15860));
  xor_4  g13512(.A(pi745), .B(new_n5785), .Y(new_n15861));
  or_6   g13513(.A(new_n15861), .B(new_n4118), .Y(new_n15862));
  nand_5 g13514(.A(new_n15862), .B(new_n15860), .Y(new_n15863));
  or_6   g13515(.A(new_n15863), .B(new_n15859), .Y(new_n15864));
  nand_5 g13516(.A(new_n15863), .B(new_n15859), .Y(new_n15865));
  nand_5 g13517(.A(new_n15865), .B(new_n6837), .Y(new_n15866));
  nand_5 g13518(.A(new_n15866), .B(new_n15864), .Y(new_n15867));
  nor_5  g13519(.A(new_n15867), .B(new_n15858), .Y(new_n15868));
  xor_4  g13520(.A(new_n15867), .B(new_n15857), .Y(new_n15869));
  nor_5  g13521(.A(new_n15869), .B(new_n4083), .Y(new_n15870));
  or_6   g13522(.A(new_n15870), .B(new_n15868), .Y(new_n15871));
  xor_4  g13523(.A(new_n15853), .B(new_n15847), .Y(new_n15872));
  not_8  g13524(.A(new_n15872), .Y(new_n15873));
  nand_5 g13525(.A(new_n15873), .B(new_n15871), .Y(new_n15874));
  xor_4  g13526(.A(new_n15873), .B(new_n15871), .Y(new_n15875));
  nand_5 g13527(.A(new_n15875), .B(new_n6835), .Y(new_n15876));
  nand_5 g13528(.A(new_n15876), .B(new_n15874), .Y(new_n15877));
  nand_5 g13529(.A(new_n15877), .B(new_n15856), .Y(new_n15878));
  or_6   g13530(.A(new_n15877), .B(new_n15856), .Y(new_n15879));
  nand_5 g13531(.A(new_n15879), .B(new_n6831), .Y(new_n15880));
  nand_5 g13532(.A(new_n15880), .B(new_n15878), .Y(new_n15881));
  xor_4  g13533(.A(new_n15881), .B(new_n6856), .Y(new_n15882));
  xor_4  g13534(.A(pi357), .B(pi347), .Y(new_n15883));
  nand_5 g13535(.A(pi770), .B(pi562), .Y(new_n15884));
  nand_5 g13536(.A(new_n15855), .B(new_n15844), .Y(new_n15885));
  nand_5 g13537(.A(new_n15885), .B(new_n15884), .Y(new_n15886));
  xor_4  g13538(.A(new_n15886), .B(new_n15883), .Y(new_n15887));
  xor_4  g13539(.A(new_n15887), .B(new_n15882), .Y(new_n15888));
  not_8  g13540(.A(new_n6835), .Y(new_n15889));
  xor_4  g13541(.A(new_n15875), .B(new_n15889), .Y(new_n15890));
  not_8  g13542(.A(new_n10511), .Y(new_n15891));
  not_8  g13543(.A(new_n5799), .Y(new_n15892));
  xor_4  g13544(.A(new_n15861), .B(new_n4118), .Y(new_n15893));
  nor_5  g13545(.A(new_n15893), .B(new_n5788), .Y(new_n15894));
  nand_5 g13546(.A(new_n15894), .B(new_n15892), .Y(new_n15895));
  xor_4  g13547(.A(new_n15894), .B(new_n15892), .Y(new_n15896));
  nand_5 g13548(.A(new_n15864), .B(new_n15865), .Y(new_n15897));
  xor_4  g13549(.A(new_n15897), .B(new_n6838), .Y(new_n15898));
  nand_5 g13550(.A(new_n15898), .B(new_n15896), .Y(new_n15899));
  nand_5 g13551(.A(new_n15899), .B(new_n15895), .Y(new_n15900));
  nand_5 g13552(.A(new_n15900), .B(new_n15891), .Y(new_n15901));
  not_8  g13553(.A(new_n15901), .Y(new_n15902));
  xor_4  g13554(.A(new_n15869), .B(new_n4083), .Y(new_n15903));
  xor_4  g13555(.A(new_n15900), .B(new_n10511), .Y(new_n15904));
  nor_5  g13556(.A(new_n15904), .B(new_n15903), .Y(new_n15905));
  nor_5  g13557(.A(new_n15905), .B(new_n15902), .Y(new_n15906));
  not_8  g13558(.A(new_n15906), .Y(new_n15907));
  nor_5  g13559(.A(new_n15907), .B(new_n15890), .Y(new_n15908));
  xor_4  g13560(.A(new_n15906), .B(new_n15890), .Y(new_n15909));
  nor_5  g13561(.A(new_n15909), .B(new_n10520), .Y(new_n15910));
  or_6   g13562(.A(new_n15910), .B(new_n15908), .Y(new_n15911));
  nand_5 g13563(.A(new_n15879), .B(new_n15878), .Y(new_n15912));
  xor_4  g13564(.A(new_n15912), .B(new_n6831), .Y(new_n15913));
  not_8  g13565(.A(new_n15913), .Y(new_n15914));
  nor_5  g13566(.A(new_n15914), .B(new_n15911), .Y(new_n15915));
  xor_4  g13567(.A(new_n15913), .B(new_n15911), .Y(new_n15916));
  nor_5  g13568(.A(new_n15916), .B(new_n10508), .Y(new_n15917));
  or_6   g13569(.A(new_n15917), .B(new_n15915), .Y(new_n15918));
  nand_5 g13570(.A(new_n15918), .B(new_n15888), .Y(new_n15919));
  xor_4  g13571(.A(new_n15918), .B(new_n15888), .Y(new_n15920));
  nand_5 g13572(.A(new_n15920), .B(new_n10507), .Y(new_n15921));
  nand_5 g13573(.A(new_n15921), .B(new_n15919), .Y(new_n15922));
  xor_4  g13574(.A(pi543), .B(pi489), .Y(new_n15923));
  nand_5 g13575(.A(pi357), .B(pi347), .Y(new_n15924));
  nand_5 g13576(.A(new_n15886), .B(new_n15883), .Y(new_n15925));
  nand_5 g13577(.A(new_n15925), .B(new_n15924), .Y(new_n15926));
  xor_4  g13578(.A(new_n15926), .B(new_n15923), .Y(new_n15927));
  not_8  g13579(.A(new_n6856), .Y(new_n15928));
  or_6   g13580(.A(new_n15881), .B(new_n15928), .Y(new_n15929));
  or_6   g13581(.A(new_n15887), .B(new_n15882), .Y(new_n15930));
  nand_5 g13582(.A(new_n15930), .B(new_n15929), .Y(new_n15931));
  xor_4  g13583(.A(new_n15931), .B(new_n15927), .Y(new_n15932));
  xor_4  g13584(.A(new_n15932), .B(new_n6862), .Y(new_n15933));
  xor_4  g13585(.A(new_n15933), .B(new_n10504), .Y(new_n15934));
  xnor_4 g13586(.A(new_n15934), .B(new_n15922), .Y(po0166));
  nor_5  g13587(.A(new_n9173), .B(new_n9171), .Y(new_n15936));
  xor_4  g13588(.A(new_n15936), .B(new_n9186), .Y(new_n15937));
  xor_4  g13589(.A(new_n15937), .B(new_n9184), .Y(po0167));
  not_8  g13590(.A(new_n2835), .Y(new_n15939));
  or_6   g13591(.A(new_n2845), .B(new_n2831), .Y(new_n15940));
  not_8  g13592(.A(new_n15940), .Y(new_n15941));
  nand_5 g13593(.A(new_n10410), .B(new_n2848), .Y(new_n15942));
  nor_5  g13594(.A(new_n15942), .B(new_n15941), .Y(new_n15943));
  nor_5  g13595(.A(new_n15943), .B(new_n15939), .Y(new_n15944));
  nand_5 g13596(.A(new_n10411), .B(new_n2848), .Y(new_n15945));
  nand_5 g13597(.A(new_n10410), .B(new_n2845), .Y(new_n15946));
  nand_5 g13598(.A(new_n15946), .B(new_n15945), .Y(new_n15947));
  nand_5 g13599(.A(new_n15947), .B(new_n15939), .Y(new_n15948));
  nand_5 g13600(.A(new_n15948), .B(new_n2830), .Y(new_n15949));
  nor_5  g13601(.A(new_n15949), .B(new_n15944), .Y(new_n15950));
  nand_5 g13602(.A(new_n2850), .B(new_n15939), .Y(new_n15951));
  nand_5 g13603(.A(new_n15951), .B(new_n2848), .Y(new_n15952));
  nand_5 g13604(.A(new_n15952), .B(new_n10411), .Y(new_n15953));
  nor_5  g13605(.A(new_n15953), .B(new_n2832), .Y(new_n15954));
  nor_5  g13606(.A(new_n15954), .B(new_n15950), .Y(new_n15955));
  nor_5  g13607(.A(new_n15955), .B(new_n14817), .Y(new_n15956));
  nor_5  g13608(.A(new_n15952), .B(new_n10411), .Y(new_n15957));
  xor_4  g13609(.A(new_n15955), .B(new_n14817), .Y(new_n15958));
  nand_5 g13610(.A(new_n14919), .B(new_n14817), .Y(new_n15959));
  not_8  g13611(.A(new_n15959), .Y(new_n15960));
  not_8  g13612(.A(new_n2830), .Y(new_n15961));
  nor_5  g13613(.A(new_n15952), .B(new_n10410), .Y(new_n15962));
  nand_5 g13614(.A(new_n15962), .B(new_n15961), .Y(new_n15963));
  nor_5  g13615(.A(new_n2850), .B(new_n15939), .Y(new_n15964));
  nand_5 g13616(.A(new_n15947), .B(new_n15964), .Y(new_n15965));
  or_6   g13617(.A(new_n2848), .B(new_n15961), .Y(new_n15966));
  nor_5  g13618(.A(new_n15946), .B(new_n2835), .Y(new_n15967));
  nand_5 g13619(.A(new_n15967), .B(new_n15966), .Y(new_n15968));
  nand_5 g13620(.A(new_n15968), .B(new_n15965), .Y(new_n15969));
  nand_5 g13621(.A(new_n15969), .B(new_n2832), .Y(new_n15970));
  and_6  g13622(.A(new_n15970), .B(new_n15963), .Y(new_n15971));
  and_6  g13623(.A(new_n15971), .B(new_n15955), .Y(new_n15972));
  nand_5 g13624(.A(new_n15972), .B(new_n15960), .Y(new_n15973));
  not_8  g13625(.A(new_n15973), .Y(new_n15974));
  nor_5  g13626(.A(new_n15974), .B(new_n15958), .Y(new_n15975));
  nor_5  g13627(.A(new_n15975), .B(new_n15957), .Y(new_n15976));
  nor_5  g13628(.A(new_n15976), .B(new_n15956), .Y(po0168));
  or_6   g13629(.A(pi439), .B(new_n2943), .Y(new_n15978));
  nand_5 g13630(.A(new_n10736), .B(new_n10724), .Y(new_n15979));
  nand_5 g13631(.A(new_n15979), .B(new_n15978), .Y(new_n15980));
  xor_4  g13632(.A(pi380), .B(pi046), .Y(new_n15981));
  xor_4  g13633(.A(new_n15981), .B(new_n15980), .Y(new_n15982));
  not_8  g13634(.A(new_n15982), .Y(new_n15983));
  nor_5  g13635(.A(new_n10761), .B(new_n10737), .Y(new_n15984));
  not_8  g13636(.A(new_n10762), .Y(new_n15985));
  nor_5  g13637(.A(new_n10798), .B(new_n15985), .Y(new_n15986));
  nor_5  g13638(.A(new_n15986), .B(new_n15984), .Y(new_n15987));
  xor_4  g13639(.A(new_n15987), .B(new_n15983), .Y(new_n15988));
  nand_5 g13640(.A(new_n9554), .B(pi473), .Y(new_n15989));
  nand_5 g13641(.A(new_n10760), .B(new_n10738), .Y(new_n15990));
  nand_5 g13642(.A(new_n15990), .B(new_n15989), .Y(new_n15991));
  nand_5 g13643(.A(pi505), .B(new_n14261), .Y(new_n15992));
  nand_5 g13644(.A(new_n8005), .B(pi459), .Y(new_n15993));
  and_6  g13645(.A(new_n15993), .B(new_n15992), .Y(new_n15994));
  xor_4  g13646(.A(new_n15994), .B(new_n15991), .Y(new_n15995));
  xor_4  g13647(.A(new_n15995), .B(new_n15988), .Y(new_n15996));
  nand_5 g13648(.A(new_n10823), .B(new_n10799), .Y(new_n15997));
  not_8  g13649(.A(new_n5569), .Y(new_n15998));
  or_6   g13650(.A(new_n10824), .B(new_n15998), .Y(new_n15999));
  nand_5 g13651(.A(new_n15999), .B(new_n15997), .Y(new_n16000));
  xor_4  g13652(.A(new_n16000), .B(new_n15996), .Y(new_n16001));
  xor_4  g13653(.A(new_n16001), .B(new_n10432), .Y(po0169));
  nand_5 g13654(.A(new_n6022), .B(new_n6023), .Y(new_n16003));
  xor_4  g13655(.A(new_n16003), .B(new_n6029), .Y(po0170));
  xor_4  g13656(.A(pi678), .B(new_n7193), .Y(new_n16005));
  nand_5 g13657(.A(pi408), .B(new_n12811), .Y(new_n16006));
  xor_4  g13658(.A(pi408), .B(new_n12811), .Y(new_n16007));
  nand_5 g13659(.A(pi423), .B(new_n12794), .Y(new_n16008));
  xor_4  g13660(.A(pi423), .B(new_n12794), .Y(new_n16009));
  nand_5 g13661(.A(new_n12776), .B(pi071), .Y(new_n16010));
  xor_4  g13662(.A(pi513), .B(new_n6997), .Y(new_n16011));
  nand_5 g13663(.A(new_n4711), .B(new_n4708), .Y(new_n16012));
  nand_5 g13664(.A(new_n16012), .B(new_n4710), .Y(new_n16013));
  nand_5 g13665(.A(new_n16013), .B(new_n16011), .Y(new_n16014));
  nand_5 g13666(.A(new_n16014), .B(new_n16010), .Y(new_n16015));
  nand_5 g13667(.A(new_n16015), .B(new_n16009), .Y(new_n16016));
  nand_5 g13668(.A(new_n16016), .B(new_n16008), .Y(new_n16017));
  nand_5 g13669(.A(new_n16017), .B(new_n16007), .Y(new_n16018));
  nand_5 g13670(.A(new_n16018), .B(new_n16006), .Y(new_n16019));
  xor_4  g13671(.A(new_n16019), .B(new_n16005), .Y(new_n16020));
  xnor_4 g13672(.A(new_n16017), .B(new_n16007), .Y(new_n16021));
  nor_5  g13673(.A(new_n16021), .B(new_n11491), .Y(new_n16022));
  xnor_4 g13674(.A(new_n16015), .B(new_n16009), .Y(new_n16023));
  nor_5  g13675(.A(new_n4713), .B(new_n4704), .Y(new_n16024));
  nand_5 g13676(.A(new_n4714), .B(new_n4678), .Y(new_n16025));
  not_8  g13677(.A(new_n16025), .Y(new_n16026));
  nor_5  g13678(.A(new_n16026), .B(new_n16024), .Y(new_n16027));
  xor_4  g13679(.A(new_n16013), .B(new_n16011), .Y(new_n16028));
  not_8  g13680(.A(new_n16028), .Y(new_n16029));
  nand_5 g13681(.A(new_n16029), .B(new_n16027), .Y(new_n16030));
  xor_4  g13682(.A(new_n16028), .B(new_n16027), .Y(new_n16031));
  or_6   g13683(.A(new_n16031), .B(new_n11458), .Y(new_n16032));
  nand_5 g13684(.A(new_n16032), .B(new_n16030), .Y(new_n16033));
  nand_5 g13685(.A(new_n16033), .B(new_n16023), .Y(new_n16034));
  xor_4  g13686(.A(new_n16033), .B(new_n16023), .Y(new_n16035));
  nand_5 g13687(.A(new_n16035), .B(new_n11453), .Y(new_n16036));
  nand_5 g13688(.A(new_n16036), .B(new_n16034), .Y(new_n16037));
  xor_4  g13689(.A(new_n16021), .B(new_n11449), .Y(new_n16038));
  nor_5  g13690(.A(new_n16038), .B(new_n16037), .Y(new_n16039));
  or_6   g13691(.A(new_n16039), .B(new_n16022), .Y(new_n16040));
  xor_4  g13692(.A(new_n16040), .B(new_n16020), .Y(new_n16041));
  not_8  g13693(.A(new_n16041), .Y(new_n16042));
  xor_4  g13694(.A(new_n16042), .B(new_n11432), .Y(po0171));
  xor_4  g13695(.A(pi512), .B(pi142), .Y(new_n16044));
  nand_5 g13696(.A(pi721), .B(pi224), .Y(new_n16045));
  xor_4  g13697(.A(pi721), .B(pi224), .Y(new_n16046));
  nand_5 g13698(.A(pi600), .B(pi417), .Y(new_n16047));
  xor_4  g13699(.A(pi600), .B(pi417), .Y(new_n16048));
  nand_5 g13700(.A(pi724), .B(pi348), .Y(new_n16049));
  xor_4  g13701(.A(pi724), .B(pi348), .Y(new_n16050));
  nand_5 g13702(.A(pi756), .B(pi659), .Y(new_n16051));
  xor_4  g13703(.A(pi756), .B(pi659), .Y(new_n16052));
  nand_5 g13704(.A(pi662), .B(pi171), .Y(new_n16053));
  nand_5 g13705(.A(new_n15475), .B(new_n15472), .Y(new_n16054));
  nand_5 g13706(.A(new_n16054), .B(new_n16053), .Y(new_n16055));
  nand_5 g13707(.A(new_n16055), .B(new_n16052), .Y(new_n16056));
  nand_5 g13708(.A(new_n16056), .B(new_n16051), .Y(new_n16057));
  nand_5 g13709(.A(new_n16057), .B(new_n16050), .Y(new_n16058));
  nand_5 g13710(.A(new_n16058), .B(new_n16049), .Y(new_n16059));
  nand_5 g13711(.A(new_n16059), .B(new_n16048), .Y(new_n16060));
  nand_5 g13712(.A(new_n16060), .B(new_n16047), .Y(new_n16061));
  nand_5 g13713(.A(new_n16061), .B(new_n16046), .Y(new_n16062));
  nand_5 g13714(.A(new_n16062), .B(new_n16045), .Y(new_n16063));
  xor_4  g13715(.A(new_n16063), .B(new_n16044), .Y(new_n16064));
  not_8  g13716(.A(new_n16064), .Y(new_n16065));
  not_8  g13717(.A(pi111), .Y(new_n16066));
  xor_4  g13718(.A(new_n16061), .B(new_n16046), .Y(new_n16067));
  not_8  g13719(.A(new_n16067), .Y(new_n16068));
  nand_5 g13720(.A(new_n16068), .B(pi537), .Y(new_n16069));
  not_8  g13721(.A(pi537), .Y(new_n16070));
  xor_4  g13722(.A(new_n16067), .B(new_n16070), .Y(new_n16071));
  xor_4  g13723(.A(new_n16059), .B(new_n16048), .Y(new_n16072));
  xor_4  g13724(.A(new_n16057), .B(new_n16050), .Y(new_n16073));
  not_8  g13725(.A(new_n16073), .Y(new_n16074));
  xor_4  g13726(.A(new_n16055), .B(new_n16052), .Y(new_n16075));
  not_8  g13727(.A(new_n16075), .Y(new_n16076));
  not_8  g13728(.A(new_n15476), .Y(new_n16077));
  nand_5 g13729(.A(new_n15479), .B(new_n16077), .Y(new_n16078));
  or_6   g13730(.A(new_n15480), .B(new_n8591), .Y(new_n16079));
  nand_5 g13731(.A(new_n16079), .B(new_n16078), .Y(new_n16080));
  nand_5 g13732(.A(new_n16080), .B(new_n16076), .Y(new_n16081));
  or_6   g13733(.A(new_n16080), .B(new_n16076), .Y(new_n16082));
  nand_5 g13734(.A(new_n16082), .B(pi026), .Y(new_n16083));
  nand_5 g13735(.A(new_n16083), .B(new_n16081), .Y(new_n16084));
  or_6   g13736(.A(new_n16084), .B(new_n16074), .Y(new_n16085));
  nand_5 g13737(.A(new_n16084), .B(new_n16074), .Y(new_n16086));
  nand_5 g13738(.A(new_n16086), .B(new_n8641), .Y(new_n16087));
  nand_5 g13739(.A(new_n16087), .B(new_n16085), .Y(new_n16088));
  nand_5 g13740(.A(new_n16088), .B(new_n16072), .Y(new_n16089));
  nand_5 g13741(.A(new_n16089), .B(pi671), .Y(new_n16090));
  or_6   g13742(.A(new_n16088), .B(new_n16072), .Y(new_n16091));
  nand_5 g13743(.A(new_n16091), .B(new_n16090), .Y(new_n16092));
  nand_5 g13744(.A(new_n16092), .B(new_n16071), .Y(new_n16093));
  nand_5 g13745(.A(new_n16093), .B(new_n16069), .Y(new_n16094));
  xor_4  g13746(.A(new_n16094), .B(new_n16066), .Y(new_n16095));
  xor_4  g13747(.A(new_n16095), .B(new_n16065), .Y(new_n16096));
  xor_4  g13748(.A(new_n16092), .B(new_n16071), .Y(new_n16097));
  not_8  g13749(.A(new_n16097), .Y(new_n16098));
  and_6  g13750(.A(new_n16082), .B(new_n16081), .Y(new_n16099));
  xor_4  g13751(.A(new_n16099), .B(pi026), .Y(new_n16100));
  not_8  g13752(.A(new_n16100), .Y(new_n16101));
  not_8  g13753(.A(pi268), .Y(new_n16102));
  nor_5  g13754(.A(new_n3235), .B(pi127), .Y(new_n16103));
  nor_5  g13755(.A(new_n5076), .B(new_n5074), .Y(new_n16104));
  nor_5  g13756(.A(new_n16104), .B(new_n16103), .Y(new_n16105));
  xor_4  g13757(.A(pi548), .B(pi074), .Y(new_n16106));
  xor_4  g13758(.A(new_n16106), .B(new_n16105), .Y(new_n16107));
  nand_5 g13759(.A(new_n16107), .B(new_n16102), .Y(new_n16108));
  nand_5 g13760(.A(new_n5078), .B(new_n5072), .Y(new_n16109));
  nand_5 g13761(.A(new_n5077), .B(new_n5073), .Y(new_n16110));
  nand_5 g13762(.A(new_n16110), .B(new_n16109), .Y(new_n16111));
  xor_4  g13763(.A(new_n16107), .B(pi268), .Y(new_n16112));
  not_8  g13764(.A(new_n16112), .Y(new_n16113));
  nand_5 g13765(.A(new_n16113), .B(new_n16111), .Y(new_n16114));
  nand_5 g13766(.A(new_n16114), .B(new_n16108), .Y(new_n16115));
  not_8  g13767(.A(pi296), .Y(new_n16116));
  xor_4  g13768(.A(pi653), .B(new_n3226), .Y(new_n16117));
  nand_5 g13769(.A(new_n5128), .B(pi074), .Y(new_n16118));
  or_6   g13770(.A(new_n16106), .B(new_n16105), .Y(new_n16119));
  nand_5 g13771(.A(new_n16119), .B(new_n16118), .Y(new_n16120));
  xnor_4 g13772(.A(new_n16120), .B(new_n16117), .Y(new_n16121));
  xor_4  g13773(.A(new_n16121), .B(new_n16116), .Y(new_n16122));
  not_8  g13774(.A(new_n16122), .Y(new_n16123));
  xor_4  g13775(.A(new_n16123), .B(new_n16115), .Y(new_n16124));
  xor_4  g13776(.A(new_n16113), .B(new_n16111), .Y(new_n16125));
  not_8  g13777(.A(new_n16125), .Y(new_n16126));
  not_8  g13778(.A(new_n5079), .Y(new_n16127));
  nand_5 g13779(.A(new_n16127), .B(new_n5071), .Y(new_n16128));
  or_6   g13780(.A(new_n5080), .B(new_n5042), .Y(new_n16129));
  nand_5 g13781(.A(new_n16129), .B(new_n16128), .Y(new_n16130));
  nor_5  g13782(.A(new_n16130), .B(new_n16126), .Y(new_n16131));
  xor_4  g13783(.A(new_n16130), .B(new_n16125), .Y(new_n16132));
  nor_5  g13784(.A(new_n16132), .B(new_n15468), .Y(new_n16133));
  or_6   g13785(.A(new_n16133), .B(new_n16131), .Y(new_n16134));
  nand_5 g13786(.A(new_n16134), .B(new_n16124), .Y(new_n16135));
  xnor_4 g13787(.A(new_n16134), .B(new_n16124), .Y(new_n16136));
  or_6   g13788(.A(new_n16136), .B(new_n15481), .Y(new_n16137));
  nand_5 g13789(.A(new_n16137), .B(new_n16135), .Y(new_n16138));
  or_6   g13790(.A(new_n16138), .B(new_n16101), .Y(new_n16139));
  xor_4  g13791(.A(new_n16138), .B(new_n16101), .Y(new_n16140));
  nand_5 g13792(.A(new_n16123), .B(new_n16115), .Y(new_n16141));
  not_8  g13793(.A(new_n16141), .Y(new_n16142));
  nor_5  g13794(.A(new_n16121), .B(pi296), .Y(new_n16143));
  nor_5  g13795(.A(new_n16143), .B(new_n16142), .Y(new_n16144));
  not_8  g13796(.A(pi392), .Y(new_n16145));
  nand_5 g13797(.A(new_n5192), .B(pi584), .Y(new_n16146));
  nand_5 g13798(.A(new_n16120), .B(new_n16117), .Y(new_n16147));
  nand_5 g13799(.A(new_n16147), .B(new_n16146), .Y(new_n16148));
  nand_5 g13800(.A(pi225), .B(new_n5196), .Y(new_n16149));
  nand_5 g13801(.A(new_n3222), .B(pi174), .Y(new_n16150));
  nand_5 g13802(.A(new_n16150), .B(new_n16149), .Y(new_n16151));
  xor_4  g13803(.A(new_n16151), .B(new_n16148), .Y(new_n16152));
  xor_4  g13804(.A(new_n16152), .B(new_n16145), .Y(new_n16153));
  not_8  g13805(.A(new_n16153), .Y(new_n16154));
  xor_4  g13806(.A(new_n16154), .B(new_n16144), .Y(new_n16155));
  nand_5 g13807(.A(new_n16155), .B(new_n16140), .Y(new_n16156));
  nand_5 g13808(.A(new_n16156), .B(new_n16139), .Y(new_n16157));
  nand_5 g13809(.A(new_n16086), .B(new_n16085), .Y(new_n16158));
  xor_4  g13810(.A(new_n16158), .B(pi768), .Y(new_n16159));
  not_8  g13811(.A(new_n16159), .Y(new_n16160));
  nor_5  g13812(.A(new_n16160), .B(new_n16157), .Y(new_n16161));
  xor_4  g13813(.A(new_n16159), .B(new_n16157), .Y(new_n16162));
  nor_5  g13814(.A(new_n16153), .B(new_n16144), .Y(new_n16163));
  nor_5  g13815(.A(new_n16152), .B(pi392), .Y(new_n16164));
  or_6   g13816(.A(new_n16164), .B(new_n16163), .Y(new_n16165));
  not_8  g13817(.A(pi287), .Y(new_n16166));
  not_8  g13818(.A(pi131), .Y(new_n16167));
  xor_4  g13819(.A(pi575), .B(new_n16167), .Y(new_n16168));
  nand_5 g13820(.A(new_n16150), .B(new_n16148), .Y(new_n16169));
  nand_5 g13821(.A(new_n16169), .B(new_n16149), .Y(new_n16170));
  xor_4  g13822(.A(new_n16170), .B(new_n16168), .Y(new_n16171));
  xor_4  g13823(.A(new_n16171), .B(new_n16166), .Y(new_n16172));
  not_8  g13824(.A(new_n16172), .Y(new_n16173));
  xor_4  g13825(.A(new_n16173), .B(new_n16165), .Y(new_n16174));
  nor_5  g13826(.A(new_n16174), .B(new_n16162), .Y(new_n16175));
  or_6   g13827(.A(new_n16175), .B(new_n16161), .Y(new_n16176));
  not_8  g13828(.A(pi671), .Y(new_n16177));
  and_6  g13829(.A(new_n16091), .B(new_n16089), .Y(new_n16178));
  xor_4  g13830(.A(new_n16178), .B(new_n16177), .Y(new_n16179));
  nand_5 g13831(.A(new_n16179), .B(new_n16176), .Y(new_n16180));
  nor_5  g13832(.A(new_n16179), .B(new_n16176), .Y(new_n16181));
  nor_5  g13833(.A(new_n16171), .B(new_n16166), .Y(new_n16182));
  nor_5  g13834(.A(new_n16173), .B(new_n16165), .Y(new_n16183));
  nor_5  g13835(.A(new_n16183), .B(new_n16182), .Y(new_n16184));
  nand_5 g13836(.A(pi575), .B(new_n16167), .Y(new_n16185));
  nand_5 g13837(.A(new_n16170), .B(new_n16168), .Y(new_n16186));
  nand_5 g13838(.A(new_n16186), .B(new_n16185), .Y(new_n16187));
  xor_4  g13839(.A(pi690), .B(pi365), .Y(new_n16188));
  xor_4  g13840(.A(new_n16188), .B(new_n16187), .Y(new_n16189));
  or_6   g13841(.A(new_n16189), .B(pi485), .Y(new_n16190));
  nand_5 g13842(.A(new_n16189), .B(pi485), .Y(new_n16191));
  nand_5 g13843(.A(new_n16191), .B(new_n16190), .Y(new_n16192));
  xor_4  g13844(.A(new_n16192), .B(new_n16184), .Y(new_n16193));
  or_6   g13845(.A(new_n16193), .B(new_n16181), .Y(new_n16194));
  nand_5 g13846(.A(new_n16194), .B(new_n16180), .Y(new_n16195));
  nand_5 g13847(.A(new_n16195), .B(new_n16098), .Y(new_n16196));
  xor_4  g13848(.A(new_n16195), .B(new_n16097), .Y(new_n16197));
  xor_4  g13849(.A(pi715), .B(new_n3213), .Y(new_n16198));
  not_8  g13850(.A(pi365), .Y(new_n16199));
  nor_5  g13851(.A(pi690), .B(new_n16199), .Y(new_n16200));
  nor_5  g13852(.A(new_n16188), .B(new_n16187), .Y(new_n16201));
  nor_5  g13853(.A(new_n16201), .B(new_n16200), .Y(new_n16202));
  xor_4  g13854(.A(new_n16202), .B(new_n16198), .Y(new_n16203));
  not_8  g13855(.A(new_n16203), .Y(new_n16204));
  xor_4  g13856(.A(new_n16204), .B(pi159), .Y(new_n16205));
  not_8  g13857(.A(new_n16205), .Y(new_n16206));
  nand_5 g13858(.A(new_n16191), .B(new_n16184), .Y(new_n16207));
  nand_5 g13859(.A(new_n16207), .B(new_n16190), .Y(new_n16208));
  xor_4  g13860(.A(new_n16208), .B(new_n16206), .Y(new_n16209));
  or_6   g13861(.A(new_n16209), .B(new_n16197), .Y(new_n16210));
  nand_5 g13862(.A(new_n16210), .B(new_n16196), .Y(new_n16211));
  nor_5  g13863(.A(new_n16211), .B(new_n16096), .Y(new_n16212));
  not_8  g13864(.A(new_n16212), .Y(new_n16213));
  nand_5 g13865(.A(new_n16211), .B(new_n16096), .Y(new_n16214));
  nand_5 g13866(.A(new_n16214), .B(new_n16213), .Y(new_n16215));
  not_8  g13867(.A(pi216), .Y(new_n16216));
  nand_5 g13868(.A(new_n16216), .B(pi166), .Y(new_n16217));
  nand_5 g13869(.A(pi216), .B(new_n3208), .Y(new_n16218));
  and_6  g13870(.A(new_n16218), .B(new_n16217), .Y(new_n16219));
  not_8  g13871(.A(pi715), .Y(new_n16220));
  nand_5 g13872(.A(new_n16220), .B(pi509), .Y(new_n16221));
  nand_5 g13873(.A(new_n16202), .B(new_n16198), .Y(new_n16222));
  nand_5 g13874(.A(new_n16222), .B(new_n16221), .Y(new_n16223));
  xor_4  g13875(.A(new_n16223), .B(new_n16219), .Y(new_n16224));
  xor_4  g13876(.A(new_n16224), .B(pi425), .Y(new_n16225));
  nand_5 g13877(.A(new_n16204), .B(pi159), .Y(new_n16226));
  not_8  g13878(.A(new_n16226), .Y(new_n16227));
  nor_5  g13879(.A(new_n16208), .B(new_n16206), .Y(new_n16228));
  nor_5  g13880(.A(new_n16228), .B(new_n16227), .Y(new_n16229));
  not_8  g13881(.A(new_n16229), .Y(new_n16230));
  xor_4  g13882(.A(new_n16230), .B(new_n16225), .Y(new_n16231));
  xor_4  g13883(.A(new_n16231), .B(new_n16215), .Y(po0172));
  nand_5 g13884(.A(new_n9651), .B(new_n9678), .Y(new_n16233));
  nand_5 g13885(.A(new_n7249), .B(new_n7244), .Y(new_n16234));
  nor_5  g13886(.A(new_n16234), .B(new_n16233), .Y(new_n16235));
  nor_5  g13887(.A(new_n9651), .B(new_n9678), .Y(new_n16236));
  and_6  g13888(.A(new_n16236), .B(new_n16234), .Y(new_n16237));
  or_6   g13889(.A(new_n16237), .B(new_n16235), .Y(new_n16238));
  xor_4  g13890(.A(new_n16238), .B(pi529), .Y(new_n16239));
  xor_4  g13891(.A(new_n16239), .B(new_n14668), .Y(new_n16240));
  xor_4  g13892(.A(pi821), .B(new_n9678), .Y(new_n16241));
  nand_5 g13893(.A(new_n16241), .B(new_n14643), .Y(new_n16242));
  nand_5 g13894(.A(pi806), .B(pi448), .Y(new_n16243));
  not_8  g13895(.A(new_n16243), .Y(new_n16244));
  nand_5 g13896(.A(new_n16244), .B(new_n16242), .Y(new_n16245));
  not_8  g13897(.A(new_n16234), .Y(new_n16246));
  nand_5 g13898(.A(new_n16241), .B(new_n16246), .Y(new_n16247));
  nand_5 g13899(.A(new_n16247), .B(new_n16245), .Y(new_n16248));
  nand_5 g13900(.A(new_n16248), .B(pi318), .Y(new_n16249));
  nand_5 g13901(.A(new_n16246), .B(new_n6568), .Y(new_n16250));
  not_8  g13902(.A(new_n16250), .Y(new_n16251));
  or_6   g13903(.A(new_n16251), .B(new_n16241), .Y(new_n16252));
  nand_5 g13904(.A(new_n16252), .B(new_n16247), .Y(new_n16253));
  nand_5 g13905(.A(new_n16253), .B(pi685), .Y(new_n16254));
  nand_5 g13906(.A(new_n16254), .B(new_n16249), .Y(new_n16255));
  nand_5 g13907(.A(new_n16255), .B(new_n16240), .Y(new_n16256));
  not_8  g13908(.A(new_n16240), .Y(new_n16257));
  nand_5 g13909(.A(new_n16257), .B(pi577), .Y(new_n16258));
  nand_5 g13910(.A(new_n16258), .B(new_n16256), .Y(new_n16259));
  nor_5  g13911(.A(new_n16259), .B(pi730), .Y(new_n16260));
  xor_4  g13912(.A(pi478), .B(pi371), .Y(new_n16261));
  nand_5 g13913(.A(new_n16239), .B(new_n11680), .Y(new_n16262));
  not_8  g13914(.A(new_n16262), .Y(new_n16263));
  nand_5 g13915(.A(new_n16263), .B(new_n16235), .Y(new_n16264));
  nor_5  g13916(.A(new_n16238), .B(pi529), .Y(new_n16265));
  nor_5  g13917(.A(new_n16265), .B(new_n16235), .Y(new_n16266));
  nand_5 g13918(.A(new_n16266), .B(new_n16262), .Y(new_n16267));
  nand_5 g13919(.A(new_n16267), .B(new_n16264), .Y(new_n16268));
  xor_4  g13920(.A(new_n16268), .B(new_n16261), .Y(new_n16269));
  xnor_4 g13921(.A(new_n16259), .B(pi730), .Y(new_n16270));
  nor_5  g13922(.A(new_n16270), .B(new_n16269), .Y(new_n16271));
  or_6   g13923(.A(new_n16271), .B(new_n16260), .Y(new_n16272));
  xor_4  g13924(.A(new_n16272), .B(pi060), .Y(new_n16273));
  xor_4  g13925(.A(pi594), .B(pi133), .Y(new_n16274));
  nand_5 g13926(.A(new_n9696), .B(new_n11674), .Y(new_n16275));
  not_8  g13927(.A(new_n16267), .Y(new_n16276));
  nor_5  g13928(.A(new_n16268), .B(new_n16261), .Y(new_n16277));
  nor_5  g13929(.A(new_n16277), .B(new_n16276), .Y(new_n16278));
  xor_4  g13930(.A(new_n16278), .B(new_n16275), .Y(new_n16279));
  xor_4  g13931(.A(new_n16279), .B(new_n16274), .Y(new_n16280));
  xor_4  g13932(.A(new_n16280), .B(new_n16273), .Y(new_n16281));
  nand_5 g13933(.A(new_n16281), .B(new_n6883), .Y(new_n16282));
  xor_4  g13934(.A(new_n16281), .B(new_n6882), .Y(new_n16283));
  xnor_4 g13935(.A(new_n16270), .B(new_n16269), .Y(new_n16284));
  nand_5 g13936(.A(new_n16284), .B(new_n6917), .Y(new_n16285));
  xor_4  g13937(.A(new_n16284), .B(new_n6889), .Y(new_n16286));
  xor_4  g13938(.A(new_n16255), .B(new_n16240), .Y(new_n16287));
  nand_5 g13939(.A(new_n16287), .B(new_n6893), .Y(new_n16288));
  xor_4  g13940(.A(new_n16287), .B(new_n6893), .Y(new_n16289));
  xor_4  g13941(.A(new_n16241), .B(new_n14643), .Y(new_n16290));
  nor_5  g13942(.A(pi448), .B(pi318), .Y(new_n16291));
  xor_4  g13943(.A(new_n6569), .B(new_n7249), .Y(new_n16292));
  nor_5  g13944(.A(new_n16292), .B(new_n16291), .Y(new_n16293));
  nand_5 g13945(.A(new_n16250), .B(new_n16243), .Y(new_n16294));
  nor_5  g13946(.A(new_n16294), .B(new_n6904), .Y(new_n16295));
  nor_5  g13947(.A(new_n16295), .B(new_n16293), .Y(new_n16296));
  nand_5 g13948(.A(new_n16292), .B(new_n6902), .Y(new_n16297));
  nand_5 g13949(.A(new_n16297), .B(new_n16244), .Y(new_n16298));
  nand_5 g13950(.A(new_n16298), .B(new_n16296), .Y(new_n16299));
  xor_4  g13951(.A(new_n16299), .B(new_n6899), .Y(new_n16300));
  xor_4  g13952(.A(new_n16300), .B(new_n16290), .Y(po0483));
  nand_5 g13953(.A(po0483), .B(new_n6900), .Y(new_n16302));
  not_8  g13954(.A(new_n16290), .Y(new_n16303));
  nor_5  g13955(.A(new_n16296), .B(new_n16303), .Y(new_n16304));
  and_6  g13956(.A(new_n16294), .B(new_n16303), .Y(new_n16305));
  and_6  g13957(.A(new_n16305), .B(new_n16298), .Y(new_n16306));
  nor_5  g13958(.A(new_n16306), .B(new_n16304), .Y(new_n16307));
  nand_5 g13959(.A(new_n16307), .B(new_n16302), .Y(new_n16308));
  nand_5 g13960(.A(new_n16308), .B(new_n16289), .Y(new_n16309));
  and_6  g13961(.A(new_n16309), .B(new_n16288), .Y(new_n16310));
  or_6   g13962(.A(new_n16310), .B(new_n16286), .Y(new_n16311));
  nand_5 g13963(.A(new_n16311), .B(new_n16285), .Y(new_n16312));
  or_6   g13964(.A(new_n16312), .B(new_n16283), .Y(new_n16313));
  nand_5 g13965(.A(new_n16313), .B(new_n16282), .Y(new_n16314));
  nor_5  g13966(.A(new_n16314), .B(new_n6878), .Y(new_n16315));
  not_8  g13967(.A(new_n6878), .Y(new_n16316));
  xor_4  g13968(.A(new_n16314), .B(new_n16316), .Y(new_n16317));
  nor_5  g13969(.A(pi594), .B(pi133), .Y(new_n16318));
  nor_5  g13970(.A(new_n16264), .B(new_n16275), .Y(new_n16319));
  nand_5 g13971(.A(new_n16319), .B(new_n16318), .Y(new_n16320));
  not_8  g13972(.A(new_n16279), .Y(new_n16321));
  nand_5 g13973(.A(new_n16321), .B(new_n16274), .Y(new_n16322));
  nor_5  g13974(.A(new_n16319), .B(new_n16318), .Y(new_n16323));
  nand_5 g13975(.A(new_n16323), .B(new_n16322), .Y(new_n16324));
  nand_5 g13976(.A(new_n16324), .B(new_n16320), .Y(new_n16325));
  xor_4  g13977(.A(pi819), .B(new_n11609), .Y(new_n16326));
  xor_4  g13978(.A(new_n16326), .B(new_n16325), .Y(new_n16327));
  not_8  g13979(.A(new_n16327), .Y(new_n16328));
  nor_5  g13980(.A(new_n16272), .B(new_n14638), .Y(new_n16329));
  not_8  g13981(.A(new_n16280), .Y(new_n16330));
  nor_5  g13982(.A(new_n16330), .B(new_n16273), .Y(new_n16331));
  or_6   g13983(.A(new_n16331), .B(new_n16329), .Y(new_n16332));
  nand_5 g13984(.A(new_n16332), .B(pi532), .Y(new_n16333));
  or_6   g13985(.A(new_n16332), .B(pi532), .Y(new_n16334));
  nand_5 g13986(.A(new_n16334), .B(new_n16333), .Y(new_n16335));
  xor_4  g13987(.A(new_n16335), .B(new_n16328), .Y(new_n16336));
  nor_5  g13988(.A(new_n16336), .B(new_n16317), .Y(new_n16337));
  or_6   g13989(.A(new_n16337), .B(new_n16315), .Y(new_n16338));
  xor_4  g13990(.A(new_n16338), .B(new_n6873), .Y(new_n16339));
  nand_5 g13991(.A(new_n16334), .B(new_n16328), .Y(new_n16340));
  nand_5 g13992(.A(new_n16340), .B(new_n16333), .Y(new_n16341));
  xor_4  g13993(.A(new_n16341), .B(new_n14634), .Y(new_n16342));
  xor_4  g13994(.A(pi808), .B(pi113), .Y(new_n16343));
  nand_5 g13995(.A(new_n16328), .B(new_n10987), .Y(new_n16344));
  nand_5 g13996(.A(new_n16324), .B(new_n11609), .Y(new_n16345));
  nor_5  g13997(.A(new_n16345), .B(new_n16344), .Y(new_n16346));
  and_6  g13998(.A(new_n16345), .B(new_n16320), .Y(new_n16347));
  and_6  g13999(.A(new_n16347), .B(new_n16344), .Y(new_n16348));
  nor_5  g14000(.A(new_n16348), .B(new_n16346), .Y(new_n16349));
  xnor_4 g14001(.A(new_n16349), .B(new_n16343), .Y(new_n16350));
  xor_4  g14002(.A(new_n16350), .B(new_n16342), .Y(new_n16351));
  xor_4  g14003(.A(new_n16351), .B(new_n16339), .Y(po0173));
  nand_5 g14004(.A(new_n5792), .B(new_n5789), .Y(new_n16353));
  xor_4  g14005(.A(new_n16353), .B(new_n5786), .Y(po0174));
  nor_5  g14006(.A(new_n5907), .B(pi436), .Y(new_n16355));
  nand_5 g14007(.A(new_n5871), .B(pi510), .Y(new_n16356));
  nand_5 g14008(.A(new_n16356), .B(new_n3441), .Y(new_n16357));
  xor_4  g14009(.A(new_n16356), .B(new_n3441), .Y(new_n16358));
  nand_5 g14010(.A(new_n16358), .B(new_n5875), .Y(new_n16359));
  nand_5 g14011(.A(new_n16359), .B(new_n16357), .Y(new_n16360));
  nand_5 g14012(.A(new_n16360), .B(new_n5870), .Y(new_n16361));
  xor_4  g14013(.A(new_n16360), .B(new_n5870), .Y(new_n16362));
  nand_5 g14014(.A(new_n16362), .B(new_n3438), .Y(new_n16363));
  nand_5 g14015(.A(new_n16363), .B(new_n16361), .Y(new_n16364));
  or_6   g14016(.A(new_n16364), .B(new_n3435), .Y(new_n16365));
  not_8  g14017(.A(new_n5866), .Y(new_n16366));
  xor_4  g14018(.A(new_n16364), .B(new_n3435), .Y(new_n16367));
  nand_5 g14019(.A(new_n16367), .B(new_n16366), .Y(new_n16368));
  nand_5 g14020(.A(new_n16368), .B(new_n16365), .Y(new_n16369));
  or_6   g14021(.A(new_n16369), .B(new_n13626), .Y(new_n16370));
  nand_5 g14022(.A(new_n16370), .B(pi300), .Y(new_n16371));
  nand_5 g14023(.A(new_n16369), .B(new_n13626), .Y(new_n16372));
  nand_5 g14024(.A(new_n16372), .B(new_n16371), .Y(new_n16373));
  nand_5 g14025(.A(new_n16373), .B(new_n5899), .Y(new_n16374));
  xor_4  g14026(.A(new_n16373), .B(new_n5899), .Y(new_n16375));
  nand_5 g14027(.A(new_n16375), .B(pi008), .Y(new_n16376));
  nand_5 g14028(.A(new_n16376), .B(new_n16374), .Y(new_n16377));
  xor_4  g14029(.A(new_n5906), .B(pi436), .Y(new_n16378));
  nor_5  g14030(.A(new_n16378), .B(new_n16377), .Y(new_n16379));
  nor_5  g14031(.A(new_n16379), .B(new_n16355), .Y(new_n16380));
  nand_5 g14032(.A(new_n16380), .B(new_n5925), .Y(new_n16381));
  or_6   g14033(.A(new_n16380), .B(new_n5925), .Y(new_n16382));
  nand_5 g14034(.A(new_n16382), .B(new_n16381), .Y(new_n16383));
  xor_4  g14035(.A(new_n16383), .B(pi227), .Y(new_n16384));
  xor_4  g14036(.A(new_n6009), .B(new_n4922), .Y(new_n16385));
  nor_5  g14037(.A(new_n5965), .B(new_n4879), .Y(new_n16386));
  not_8  g14038(.A(new_n8548), .Y(new_n16387));
  nor_5  g14039(.A(new_n8574), .B(new_n16387), .Y(new_n16388));
  nor_5  g14040(.A(new_n16388), .B(new_n16386), .Y(new_n16389));
  xor_4  g14041(.A(new_n16389), .B(new_n16385), .Y(new_n16390));
  xor_4  g14042(.A(new_n16375), .B(pi008), .Y(new_n16391));
  xor_4  g14043(.A(new_n16367), .B(new_n5866), .Y(new_n16392));
  nor_5  g14044(.A(new_n16392), .B(new_n8599), .Y(new_n16393));
  xor_4  g14045(.A(new_n16362), .B(pi011), .Y(new_n16394));
  nor_5  g14046(.A(new_n16394), .B(new_n8600), .Y(new_n16395));
  xor_4  g14047(.A(new_n16394), .B(new_n8601), .Y(new_n16396));
  nand_5 g14048(.A(new_n6024), .B(pi230), .Y(new_n16397));
  nand_5 g14049(.A(new_n6026), .B(new_n3448), .Y(new_n16398));
  nand_5 g14050(.A(new_n16398), .B(new_n8610), .Y(new_n16399));
  nand_5 g14051(.A(new_n16399), .B(new_n16397), .Y(new_n16400));
  nand_5 g14052(.A(new_n16400), .B(new_n8621), .Y(new_n16401));
  xor_4  g14053(.A(new_n5871), .B(new_n3445), .Y(new_n16402));
  not_8  g14054(.A(new_n8621), .Y(new_n16403));
  xor_4  g14055(.A(new_n16400), .B(new_n16403), .Y(new_n16404));
  or_6   g14056(.A(new_n16404), .B(new_n16402), .Y(new_n16405));
  nand_5 g14057(.A(new_n16405), .B(new_n16401), .Y(new_n16406));
  nand_5 g14058(.A(new_n16406), .B(new_n8604), .Y(new_n16407));
  xor_4  g14059(.A(new_n16406), .B(new_n8605), .Y(new_n16408));
  xor_4  g14060(.A(new_n16358), .B(new_n5875), .Y(new_n16409));
  or_6   g14061(.A(new_n16409), .B(new_n16408), .Y(new_n16410));
  nand_5 g14062(.A(new_n16410), .B(new_n16407), .Y(new_n16411));
  nor_5  g14063(.A(new_n16411), .B(new_n16396), .Y(new_n16412));
  or_6   g14064(.A(new_n16412), .B(new_n16395), .Y(new_n16413));
  xor_4  g14065(.A(new_n16392), .B(new_n8598), .Y(new_n16414));
  nor_5  g14066(.A(new_n16414), .B(new_n16413), .Y(new_n16415));
  or_6   g14067(.A(new_n16415), .B(new_n16393), .Y(new_n16416));
  nand_5 g14068(.A(new_n16372), .B(new_n16370), .Y(new_n16417));
  xor_4  g14069(.A(new_n16417), .B(pi300), .Y(new_n16418));
  not_8  g14070(.A(new_n16418), .Y(new_n16419));
  nor_5  g14071(.A(new_n16419), .B(new_n16416), .Y(new_n16420));
  xor_4  g14072(.A(new_n16418), .B(new_n16416), .Y(new_n16421));
  nor_5  g14073(.A(new_n16421), .B(new_n8635), .Y(new_n16422));
  nor_5  g14074(.A(new_n16422), .B(new_n16420), .Y(new_n16423));
  nand_5 g14075(.A(new_n16423), .B(new_n16391), .Y(new_n16424));
  not_8  g14076(.A(new_n8575), .Y(new_n16425));
  xnor_4 g14077(.A(new_n16423), .B(new_n16391), .Y(new_n16426));
  or_6   g14078(.A(new_n16426), .B(new_n16425), .Y(new_n16427));
  nand_5 g14079(.A(new_n16427), .B(new_n16424), .Y(new_n16428));
  nand_5 g14080(.A(new_n16428), .B(new_n16390), .Y(new_n16429));
  not_8  g14081(.A(new_n16390), .Y(new_n16430));
  xor_4  g14082(.A(new_n16428), .B(new_n16430), .Y(new_n16431));
  xor_4  g14083(.A(new_n16378), .B(new_n16377), .Y(new_n16432));
  or_6   g14084(.A(new_n16432), .B(new_n16431), .Y(new_n16433));
  nand_5 g14085(.A(new_n16433), .B(new_n16429), .Y(new_n16434));
  nand_5 g14086(.A(new_n6009), .B(new_n4922), .Y(new_n16435));
  nand_5 g14087(.A(new_n16389), .B(new_n16385), .Y(new_n16436));
  nand_5 g14088(.A(new_n16436), .B(new_n16435), .Y(new_n16437));
  or_6   g14089(.A(new_n6073), .B(pi093), .Y(new_n16438));
  nand_5 g14090(.A(new_n6073), .B(pi093), .Y(new_n16439));
  and_6  g14091(.A(new_n16439), .B(new_n16438), .Y(new_n16440));
  xor_4  g14092(.A(new_n16440), .B(new_n16437), .Y(new_n16441));
  not_8  g14093(.A(new_n16441), .Y(new_n16442));
  xor_4  g14094(.A(new_n16442), .B(new_n16434), .Y(new_n16443));
  xnor_4 g14095(.A(new_n16443), .B(new_n16384), .Y(po0175));
  and_6  g14096(.A(new_n13233), .B(new_n10400), .Y(new_n16445));
  nor_5  g14097(.A(new_n16445), .B(new_n13230), .Y(new_n16446));
  nand_5 g14098(.A(new_n13224), .B(new_n13218), .Y(new_n16447));
  nand_5 g14099(.A(new_n16447), .B(new_n13219), .Y(new_n16448));
  xor_4  g14100(.A(new_n16448), .B(new_n16446), .Y(new_n16449));
  not_8  g14101(.A(new_n13226), .Y(new_n16450));
  nand_5 g14102(.A(new_n13234), .B(new_n16450), .Y(new_n16451));
  not_8  g14103(.A(new_n13235), .Y(new_n16452));
  nand_5 g14104(.A(new_n13237), .B(new_n16452), .Y(new_n16453));
  nand_5 g14105(.A(new_n16453), .B(new_n16451), .Y(new_n16454));
  xor_4  g14106(.A(new_n16454), .B(new_n16449), .Y(new_n16455));
  not_8  g14107(.A(new_n16455), .Y(new_n16456));
  nand_5 g14108(.A(new_n5404), .B(new_n4160), .Y(new_n16457));
  or_6   g14109(.A(new_n5404), .B(new_n4160), .Y(new_n16458));
  nor_5  g14110(.A(new_n5348), .B(new_n4187), .Y(new_n16459));
  nor_5  g14111(.A(new_n16459), .B(new_n4183), .Y(new_n16460));
  not_8  g14112(.A(new_n4183), .Y(new_n16461));
  xor_4  g14113(.A(new_n16459), .B(new_n16461), .Y(new_n16462));
  nor_5  g14114(.A(new_n16462), .B(new_n5364), .Y(new_n16463));
  or_6   g14115(.A(new_n16463), .B(new_n16460), .Y(new_n16464));
  nand_5 g14116(.A(new_n16464), .B(new_n4176), .Y(new_n16465));
  xor_4  g14117(.A(new_n16464), .B(new_n4175), .Y(new_n16466));
  or_6   g14118(.A(new_n16466), .B(new_n5421), .Y(new_n16467));
  nand_5 g14119(.A(new_n16467), .B(new_n16465), .Y(new_n16468));
  nand_5 g14120(.A(new_n16468), .B(new_n16458), .Y(new_n16469));
  nand_5 g14121(.A(new_n16469), .B(new_n16457), .Y(new_n16470));
  nand_5 g14122(.A(new_n16470), .B(new_n5431), .Y(new_n16471));
  not_8  g14123(.A(new_n16471), .Y(new_n16472));
  nor_5  g14124(.A(new_n16470), .B(new_n5431), .Y(new_n16473));
  nor_5  g14125(.A(new_n16473), .B(new_n4244), .Y(new_n16474));
  nor_5  g14126(.A(new_n16474), .B(new_n16472), .Y(new_n16475));
  nand_5 g14127(.A(new_n16475), .B(new_n14977), .Y(new_n16476));
  xor_4  g14128(.A(new_n16475), .B(new_n14978), .Y(new_n16477));
  or_6   g14129(.A(new_n16477), .B(new_n5435), .Y(new_n16478));
  nand_5 g14130(.A(new_n16478), .B(new_n16476), .Y(new_n16479));
  nor_5  g14131(.A(new_n16479), .B(new_n15054), .Y(new_n16480));
  xor_4  g14132(.A(new_n16479), .B(new_n15033), .Y(new_n16481));
  nor_5  g14133(.A(new_n16481), .B(new_n5444), .Y(new_n16482));
  or_6   g14134(.A(new_n16482), .B(new_n16480), .Y(new_n16483));
  nor_5  g14135(.A(new_n16483), .B(new_n15053), .Y(new_n16484));
  xor_4  g14136(.A(new_n16483), .B(new_n15053), .Y(new_n16485));
  nand_5 g14137(.A(new_n16485), .B(new_n5396), .Y(new_n16486));
  not_8  g14138(.A(new_n16486), .Y(new_n16487));
  nor_5  g14139(.A(new_n16487), .B(new_n16484), .Y(new_n16488));
  nand_5 g14140(.A(new_n16488), .B(new_n5393), .Y(new_n16489));
  xor_4  g14141(.A(new_n16488), .B(new_n5393), .Y(new_n16490));
  nand_5 g14142(.A(new_n16490), .B(new_n15068), .Y(new_n16491));
  nand_5 g14143(.A(new_n16491), .B(new_n16489), .Y(new_n16492));
  nand_5 g14144(.A(new_n16492), .B(new_n15084), .Y(new_n16493));
  xor_4  g14145(.A(new_n16492), .B(new_n15084), .Y(new_n16494));
  nand_5 g14146(.A(new_n16494), .B(new_n13238), .Y(new_n16495));
  nand_5 g14147(.A(new_n16495), .B(new_n16493), .Y(new_n16496));
  xor_4  g14148(.A(new_n16496), .B(new_n16456), .Y(new_n16497));
  xor_4  g14149(.A(new_n16497), .B(new_n15102), .Y(po0176));
  xor_4  g14150(.A(new_n10856), .B(pi762), .Y(new_n16499));
  nor_5  g14151(.A(new_n15504), .B(new_n10857), .Y(new_n16500));
  nor_5  g14152(.A(new_n15505), .B(new_n15491), .Y(new_n16501));
  or_6   g14153(.A(new_n16501), .B(new_n16500), .Y(new_n16502));
  or_6   g14154(.A(new_n16502), .B(new_n10883), .Y(new_n16503));
  nand_5 g14155(.A(new_n16503), .B(pi165), .Y(new_n16504));
  nand_5 g14156(.A(new_n16502), .B(new_n10883), .Y(new_n16505));
  nand_5 g14157(.A(new_n16505), .B(new_n16504), .Y(new_n16506));
  xor_4  g14158(.A(new_n16506), .B(new_n16499), .Y(new_n16507));
  not_8  g14159(.A(new_n16507), .Y(new_n16508));
  nand_5 g14160(.A(new_n15523), .B(new_n15507), .Y(new_n16509));
  nand_5 g14161(.A(new_n15524), .B(new_n10001), .Y(new_n16510));
  nand_5 g14162(.A(new_n16510), .B(new_n16509), .Y(new_n16511));
  nand_5 g14163(.A(new_n16505), .B(new_n16503), .Y(new_n16512));
  xor_4  g14164(.A(new_n16512), .B(pi165), .Y(new_n16513));
  nand_5 g14165(.A(new_n16513), .B(new_n16511), .Y(new_n16514));
  not_8  g14166(.A(new_n10029), .Y(new_n16515));
  xor_4  g14167(.A(new_n16513), .B(new_n16511), .Y(new_n16516));
  nand_5 g14168(.A(new_n16516), .B(new_n16515), .Y(new_n16517));
  nand_5 g14169(.A(new_n16517), .B(new_n16514), .Y(new_n16518));
  xor_4  g14170(.A(new_n16518), .B(new_n16508), .Y(new_n16519));
  xor_4  g14171(.A(new_n16519), .B(new_n10049), .Y(po0177));
  xor_4  g14172(.A(new_n9133), .B(new_n9132), .Y(po0178));
  nand_5 g14173(.A(pi543), .B(pi489), .Y(new_n16522));
  nand_5 g14174(.A(new_n15926), .B(new_n15923), .Y(new_n16523));
  nand_5 g14175(.A(new_n16523), .B(new_n16522), .Y(new_n16524));
  nand_5 g14176(.A(pi668), .B(pi014), .Y(new_n16525));
  not_8  g14177(.A(pi014), .Y(new_n16526));
  nand_5 g14178(.A(new_n10459), .B(new_n16526), .Y(new_n16527));
  nand_5 g14179(.A(new_n16527), .B(new_n16525), .Y(new_n16528));
  xor_4  g14180(.A(new_n16528), .B(new_n16524), .Y(new_n16529));
  or_6   g14181(.A(new_n16529), .B(new_n6827), .Y(new_n16530));
  xor_4  g14182(.A(new_n16529), .B(new_n6827), .Y(new_n16531));
  not_8  g14183(.A(new_n15931), .Y(new_n16532));
  nand_5 g14184(.A(new_n16532), .B(new_n15927), .Y(new_n16533));
  or_6   g14185(.A(new_n15932), .B(new_n6874), .Y(new_n16534));
  nand_5 g14186(.A(new_n16534), .B(new_n16533), .Y(new_n16535));
  nand_5 g14187(.A(new_n16535), .B(new_n16531), .Y(new_n16536));
  nand_5 g14188(.A(new_n16536), .B(new_n16530), .Y(new_n16537));
  xor_4  g14189(.A(pi571), .B(pi137), .Y(new_n16538));
  nand_5 g14190(.A(new_n16527), .B(new_n16524), .Y(new_n16539));
  nand_5 g14191(.A(new_n16539), .B(new_n16525), .Y(new_n16540));
  xor_4  g14192(.A(new_n16540), .B(new_n16538), .Y(new_n16541));
  nand_5 g14193(.A(new_n16541), .B(new_n16537), .Y(new_n16542));
  xor_4  g14194(.A(new_n16541), .B(new_n16537), .Y(new_n16543));
  nand_5 g14195(.A(new_n16543), .B(new_n6944), .Y(new_n16544));
  nand_5 g14196(.A(new_n16544), .B(new_n16542), .Y(new_n16545));
  xor_4  g14197(.A(pi461), .B(pi084), .Y(new_n16546));
  nand_5 g14198(.A(pi571), .B(pi137), .Y(new_n16547));
  nand_5 g14199(.A(new_n16540), .B(new_n16538), .Y(new_n16548));
  nand_5 g14200(.A(new_n16548), .B(new_n16547), .Y(new_n16549));
  xor_4  g14201(.A(new_n16549), .B(new_n16546), .Y(new_n16550));
  nand_5 g14202(.A(new_n16550), .B(new_n16545), .Y(new_n16551));
  xnor_4 g14203(.A(new_n16550), .B(new_n16545), .Y(new_n16552));
  or_6   g14204(.A(new_n16552), .B(new_n12085), .Y(new_n16553));
  nand_5 g14205(.A(new_n16553), .B(new_n16551), .Y(new_n16554));
  xor_4  g14206(.A(new_n16552), .B(new_n12085), .Y(new_n16555));
  not_8  g14207(.A(new_n16555), .Y(new_n16556));
  xor_4  g14208(.A(new_n16543), .B(new_n6943), .Y(new_n16557));
  nand_5 g14209(.A(new_n16557), .B(new_n10501), .Y(new_n16558));
  xor_4  g14210(.A(new_n16557), .B(new_n10501), .Y(new_n16559));
  xor_4  g14211(.A(new_n16535), .B(new_n16531), .Y(new_n16560));
  nor_5  g14212(.A(new_n15933), .B(new_n10505), .Y(new_n16561));
  nor_5  g14213(.A(new_n15934), .B(new_n15922), .Y(new_n16562));
  or_6   g14214(.A(new_n16562), .B(new_n16561), .Y(new_n16563));
  or_6   g14215(.A(new_n16563), .B(new_n16560), .Y(new_n16564));
  xor_4  g14216(.A(new_n16563), .B(new_n16560), .Y(new_n16565));
  nand_5 g14217(.A(new_n16565), .B(new_n10503), .Y(new_n16566));
  nand_5 g14218(.A(new_n16566), .B(new_n16564), .Y(new_n16567));
  nand_5 g14219(.A(new_n16567), .B(new_n16559), .Y(new_n16568));
  nand_5 g14220(.A(new_n16568), .B(new_n16558), .Y(new_n16569));
  nor_5  g14221(.A(new_n16569), .B(new_n16556), .Y(new_n16570));
  xor_4  g14222(.A(new_n16569), .B(new_n16555), .Y(new_n16571));
  nor_5  g14223(.A(new_n16571), .B(new_n10551), .Y(new_n16572));
  or_6   g14224(.A(new_n16572), .B(new_n16570), .Y(new_n16573));
  nand_5 g14225(.A(new_n16573), .B(new_n16554), .Y(new_n16574));
  not_8  g14226(.A(new_n16574), .Y(new_n16575));
  nand_5 g14227(.A(pi461), .B(pi084), .Y(new_n16576));
  nand_5 g14228(.A(new_n16549), .B(new_n16546), .Y(new_n16577));
  nand_5 g14229(.A(new_n16577), .B(new_n16576), .Y(new_n16578));
  or_6   g14230(.A(new_n16578), .B(new_n10563), .Y(new_n16579));
  nand_5 g14231(.A(new_n16578), .B(new_n10563), .Y(new_n16580));
  nand_5 g14232(.A(new_n16580), .B(new_n16579), .Y(new_n16581));
  or_6   g14233(.A(new_n16581), .B(new_n12083), .Y(new_n16582));
  nand_5 g14234(.A(new_n16582), .B(new_n16579), .Y(new_n16583));
  not_8  g14235(.A(new_n16583), .Y(new_n16584));
  nand_5 g14236(.A(new_n16584), .B(new_n16575), .Y(new_n16585));
  nor_5  g14237(.A(new_n16573), .B(new_n16554), .Y(new_n16586));
  not_8  g14238(.A(new_n16586), .Y(new_n16587));
  nor_5  g14239(.A(new_n16580), .B(new_n12082), .Y(new_n16588));
  nand_5 g14240(.A(new_n16588), .B(new_n16587), .Y(new_n16589));
  nand_5 g14241(.A(new_n16589), .B(new_n16585), .Y(po0269));
  or_6   g14242(.A(new_n16579), .B(new_n12083), .Y(new_n16591));
  or_6   g14243(.A(new_n16591), .B(new_n16575), .Y(new_n16592));
  nand_5 g14244(.A(new_n16586), .B(new_n16583), .Y(new_n16593));
  nand_5 g14245(.A(new_n16593), .B(new_n16592), .Y(new_n16594));
  or_6   g14246(.A(new_n16594), .B(po0269), .Y(po0179));
  xnor_4 g14247(.A(new_n3882), .B(new_n3851), .Y(po0180));
  xnor_4 g14248(.A(new_n13639), .B(new_n3482), .Y(po0181));
  nand_5 g14249(.A(new_n4984), .B(new_n4734), .Y(new_n16598));
  not_8  g14250(.A(new_n4988), .Y(new_n16599));
  nand_5 g14251(.A(new_n10980), .B(new_n16599), .Y(new_n16600));
  nand_5 g14252(.A(new_n16600), .B(new_n4987), .Y(new_n16601));
  xnor_4 g14253(.A(new_n16601), .B(new_n16598), .Y(new_n16602));
  nor_5  g14254(.A(pi670), .B(pi455), .Y(new_n16603));
  nor_5  g14255(.A(new_n10979), .B(new_n6026), .Y(new_n16604));
  nor_5  g14256(.A(new_n16604), .B(new_n16603), .Y(new_n16605));
  xor_4  g14257(.A(new_n16605), .B(new_n13253), .Y(new_n16606));
  xor_4  g14258(.A(new_n16606), .B(new_n5855), .Y(new_n16607));
  xnor_4 g14259(.A(new_n16607), .B(new_n16602), .Y(po0182));
  xor_4  g14260(.A(new_n12361), .B(new_n8841), .Y(po0183));
  xor_4  g14261(.A(new_n14958), .B(new_n4214), .Y(po0184));
  not_8  g14262(.A(pi774), .Y(new_n16611));
  nand_5 g14263(.A(pi642), .B(pi622), .Y(new_n16612));
  and_6  g14264(.A(new_n16612), .B(new_n16611), .Y(new_n16613));
  nor_5  g14265(.A(new_n16612), .B(new_n16611), .Y(new_n16614));
  nor_5  g14266(.A(new_n16614), .B(new_n16613), .Y(new_n16615));
  xor_4  g14267(.A(pi255), .B(pi163), .Y(new_n16616));
  not_8  g14268(.A(new_n16616), .Y(new_n16617));
  xor_4  g14269(.A(new_n16617), .B(new_n16615), .Y(new_n16618));
  nand_5 g14270(.A(new_n16618), .B(pi477), .Y(new_n16619));
  not_8  g14271(.A(new_n15761), .Y(new_n16620));
  xor_4  g14272(.A(pi642), .B(pi622), .Y(new_n16621));
  nor_5  g14273(.A(new_n16621), .B(new_n16620), .Y(new_n16622));
  nand_5 g14274(.A(new_n16622), .B(pi477), .Y(new_n16623));
  not_8  g14275(.A(new_n16618), .Y(new_n16624));
  nand_5 g14276(.A(new_n16621), .B(new_n16620), .Y(new_n16625));
  nor_5  g14277(.A(new_n16625), .B(pi477), .Y(new_n16626));
  not_8  g14278(.A(new_n16626), .Y(new_n16627));
  nand_5 g14279(.A(new_n16627), .B(new_n16623), .Y(new_n16628));
  or_6   g14280(.A(new_n16628), .B(new_n16624), .Y(new_n16629));
  nand_5 g14281(.A(new_n16629), .B(new_n16623), .Y(new_n16630));
  nand_5 g14282(.A(new_n16630), .B(new_n16619), .Y(new_n16631));
  xor_4  g14283(.A(new_n16628), .B(new_n16618), .Y(new_n16632));
  or_6   g14284(.A(new_n16632), .B(new_n15767), .Y(new_n16633));
  nand_5 g14285(.A(new_n16633), .B(new_n16631), .Y(new_n16634));
  nand_5 g14286(.A(new_n16624), .B(pi163), .Y(new_n16635));
  nand_5 g14287(.A(new_n16635), .B(new_n16619), .Y(new_n16636));
  not_8  g14288(.A(pi595), .Y(new_n16637));
  xor_4  g14289(.A(pi658), .B(pi017), .Y(new_n16638));
  nor_5  g14290(.A(new_n16614), .B(pi255), .Y(new_n16639));
  nor_5  g14291(.A(new_n16639), .B(new_n16613), .Y(new_n16640));
  xor_4  g14292(.A(new_n16640), .B(new_n16638), .Y(new_n16641));
  or_6   g14293(.A(new_n16641), .B(new_n16637), .Y(new_n16642));
  nand_5 g14294(.A(new_n16641), .B(new_n16637), .Y(new_n16643));
  nand_5 g14295(.A(new_n16643), .B(new_n16642), .Y(new_n16644));
  xor_4  g14296(.A(new_n16644), .B(new_n16636), .Y(new_n16645));
  xor_4  g14297(.A(new_n16645), .B(new_n15759), .Y(new_n16646));
  xor_4  g14298(.A(new_n16646), .B(new_n16634), .Y(po0185));
  xnor_4 g14299(.A(new_n16409), .B(new_n16408), .Y(po0186));
  xor_4  g14300(.A(pi571), .B(new_n6307), .Y(new_n16649));
  nand_5 g14301(.A(new_n8865), .B(pi014), .Y(new_n16650));
  xor_4  g14302(.A(pi205), .B(new_n16526), .Y(new_n16651));
  nand_5 g14303(.A(new_n8868), .B(pi543), .Y(new_n16652));
  xor_4  g14304(.A(new_n8868), .B(pi543), .Y(new_n16653));
  nand_5 g14305(.A(new_n6201), .B(pi347), .Y(new_n16654));
  nand_5 g14306(.A(pi770), .B(new_n6165), .Y(new_n16655));
  nand_5 g14307(.A(pi596), .B(new_n8875), .Y(new_n16656));
  xor_4  g14308(.A(pi596), .B(new_n8875), .Y(new_n16657));
  nand_5 g14309(.A(new_n12096), .B(pi051), .Y(new_n16658));
  nand_5 g14310(.A(new_n4093), .B(new_n4085), .Y(new_n16659));
  nand_5 g14311(.A(new_n16659), .B(new_n16658), .Y(new_n16660));
  nand_5 g14312(.A(new_n16660), .B(new_n16657), .Y(new_n16661));
  nand_5 g14313(.A(new_n16661), .B(new_n16656), .Y(new_n16662));
  xor_4  g14314(.A(pi770), .B(pi644), .Y(new_n16663));
  not_8  g14315(.A(new_n16663), .Y(new_n16664));
  nand_5 g14316(.A(new_n16664), .B(new_n16662), .Y(new_n16665));
  nand_5 g14317(.A(new_n16665), .B(new_n16655), .Y(new_n16666));
  xor_4  g14318(.A(pi726), .B(pi347), .Y(new_n16667));
  not_8  g14319(.A(new_n16667), .Y(new_n16668));
  nand_5 g14320(.A(new_n16668), .B(new_n16666), .Y(new_n16669));
  nand_5 g14321(.A(new_n16669), .B(new_n16654), .Y(new_n16670));
  nand_5 g14322(.A(new_n16670), .B(new_n16653), .Y(new_n16671));
  nand_5 g14323(.A(new_n16671), .B(new_n16652), .Y(new_n16672));
  nand_5 g14324(.A(new_n16672), .B(new_n16651), .Y(new_n16673));
  nand_5 g14325(.A(new_n16673), .B(new_n16650), .Y(new_n16674));
  xor_4  g14326(.A(new_n16674), .B(new_n16649), .Y(new_n16675));
  xor_4  g14327(.A(new_n16667), .B(new_n16666), .Y(new_n16676));
  not_8  g14328(.A(new_n16676), .Y(new_n16677));
  xor_4  g14329(.A(new_n16660), .B(new_n16657), .Y(new_n16678));
  nand_5 g14330(.A(new_n4107), .B(new_n4094), .Y(new_n16679));
  or_6   g14331(.A(new_n4108), .B(new_n4083), .Y(new_n16680));
  nand_5 g14332(.A(new_n16680), .B(new_n16679), .Y(new_n16681));
  nand_5 g14333(.A(new_n16681), .B(new_n16678), .Y(new_n16682));
  xor_4  g14334(.A(new_n16681), .B(new_n16678), .Y(new_n16683));
  nand_5 g14335(.A(new_n16683), .B(new_n6835), .Y(new_n16684));
  nand_5 g14336(.A(new_n16684), .B(new_n16682), .Y(new_n16685));
  xor_4  g14337(.A(new_n16663), .B(new_n16662), .Y(new_n16686));
  not_8  g14338(.A(new_n16686), .Y(new_n16687));
  nand_5 g14339(.A(new_n16687), .B(new_n16685), .Y(new_n16688));
  or_6   g14340(.A(new_n16687), .B(new_n16685), .Y(new_n16689));
  nand_5 g14341(.A(new_n16689), .B(new_n6831), .Y(new_n16690));
  nand_5 g14342(.A(new_n16690), .B(new_n16688), .Y(new_n16691));
  nand_5 g14343(.A(new_n16691), .B(new_n16677), .Y(new_n16692));
  xor_4  g14344(.A(new_n16691), .B(new_n16676), .Y(new_n16693));
  or_6   g14345(.A(new_n16693), .B(new_n6856), .Y(new_n16694));
  nand_5 g14346(.A(new_n16694), .B(new_n16692), .Y(new_n16695));
  nand_5 g14347(.A(new_n16695), .B(new_n6862), .Y(new_n16696));
  xor_4  g14348(.A(new_n16670), .B(new_n16653), .Y(new_n16697));
  xor_4  g14349(.A(new_n16695), .B(new_n6862), .Y(new_n16698));
  nand_5 g14350(.A(new_n16698), .B(new_n16697), .Y(new_n16699));
  nand_5 g14351(.A(new_n16699), .B(new_n16696), .Y(new_n16700));
  nor_5  g14352(.A(new_n16700), .B(new_n6828), .Y(new_n16701));
  xor_4  g14353(.A(new_n16672), .B(new_n16651), .Y(new_n16702));
  xor_4  g14354(.A(new_n16700), .B(new_n6827), .Y(new_n16703));
  nor_5  g14355(.A(new_n16703), .B(new_n16702), .Y(new_n16704));
  or_6   g14356(.A(new_n16704), .B(new_n16701), .Y(new_n16705));
  xor_4  g14357(.A(new_n16705), .B(new_n16675), .Y(new_n16706));
  xor_4  g14358(.A(new_n16706), .B(new_n6944), .Y(new_n16707));
  nor_5  g14359(.A(new_n16707), .B(new_n6329), .Y(new_n16708));
  xor_4  g14360(.A(new_n16707), .B(new_n6301), .Y(new_n16709));
  xor_4  g14361(.A(new_n16698), .B(new_n16697), .Y(new_n16710));
  not_8  g14362(.A(new_n16710), .Y(new_n16711));
  xor_4  g14363(.A(new_n16693), .B(new_n15928), .Y(new_n16712));
  nand_5 g14364(.A(new_n16712), .B(new_n6124), .Y(new_n16713));
  xor_4  g14365(.A(new_n16712), .B(new_n6124), .Y(new_n16714));
  xor_4  g14366(.A(new_n16683), .B(new_n15889), .Y(new_n16715));
  nand_5 g14367(.A(new_n4126), .B(new_n4114), .Y(new_n16716));
  not_8  g14368(.A(new_n16716), .Y(new_n16717));
  nor_5  g14369(.A(new_n4128), .B(new_n4109), .Y(new_n16718));
  nor_5  g14370(.A(new_n16718), .B(new_n16717), .Y(new_n16719));
  not_8  g14371(.A(new_n16719), .Y(new_n16720));
  nor_5  g14372(.A(new_n16720), .B(new_n16715), .Y(new_n16721));
  xor_4  g14373(.A(new_n16719), .B(new_n16715), .Y(new_n16722));
  nor_5  g14374(.A(new_n16722), .B(new_n6178), .Y(new_n16723));
  or_6   g14375(.A(new_n16723), .B(new_n16721), .Y(new_n16724));
  nand_5 g14376(.A(new_n16689), .B(new_n16688), .Y(new_n16725));
  xor_4  g14377(.A(new_n16725), .B(new_n6831), .Y(new_n16726));
  not_8  g14378(.A(new_n16726), .Y(new_n16727));
  nor_5  g14379(.A(new_n16727), .B(new_n16724), .Y(new_n16728));
  xor_4  g14380(.A(new_n16726), .B(new_n16724), .Y(new_n16729));
  nor_5  g14381(.A(new_n16729), .B(new_n6173), .Y(new_n16730));
  or_6   g14382(.A(new_n16730), .B(new_n16728), .Y(new_n16731));
  nand_5 g14383(.A(new_n16731), .B(new_n16714), .Y(new_n16732));
  nand_5 g14384(.A(new_n16732), .B(new_n16713), .Y(new_n16733));
  nor_5  g14385(.A(new_n16733), .B(new_n16711), .Y(new_n16734));
  not_8  g14386(.A(new_n6225), .Y(new_n16735));
  xor_4  g14387(.A(new_n16733), .B(new_n16710), .Y(new_n16736));
  nor_5  g14388(.A(new_n16736), .B(new_n16735), .Y(new_n16737));
  or_6   g14389(.A(new_n16737), .B(new_n16734), .Y(new_n16738));
  not_8  g14390(.A(new_n16702), .Y(new_n16739));
  xor_4  g14391(.A(new_n16703), .B(new_n16739), .Y(new_n16740));
  or_6   g14392(.A(new_n16740), .B(new_n16738), .Y(new_n16741));
  nand_5 g14393(.A(new_n16740), .B(new_n16738), .Y(new_n16742));
  nand_5 g14394(.A(new_n16742), .B(new_n6269), .Y(new_n16743));
  nand_5 g14395(.A(new_n16743), .B(new_n16741), .Y(new_n16744));
  nor_5  g14396(.A(new_n16744), .B(new_n16709), .Y(new_n16745));
  nor_5  g14397(.A(new_n16745), .B(new_n16708), .Y(new_n16746));
  not_8  g14398(.A(pi084), .Y(new_n16747));
  xor_4  g14399(.A(pi335), .B(new_n16747), .Y(new_n16748));
  nand_5 g14400(.A(pi571), .B(new_n6307), .Y(new_n16749));
  nand_5 g14401(.A(new_n16674), .B(new_n16649), .Y(new_n16750));
  nand_5 g14402(.A(new_n16750), .B(new_n16749), .Y(new_n16751));
  xor_4  g14403(.A(new_n16751), .B(new_n16748), .Y(new_n16752));
  not_8  g14404(.A(new_n16675), .Y(new_n16753));
  nor_5  g14405(.A(new_n16705), .B(new_n16753), .Y(new_n16754));
  nor_5  g14406(.A(new_n16706), .B(new_n6943), .Y(new_n16755));
  or_6   g14407(.A(new_n16755), .B(new_n16754), .Y(new_n16756));
  xnor_4 g14408(.A(new_n16756), .B(new_n16752), .Y(new_n16757));
  xor_4  g14409(.A(new_n16757), .B(new_n12086), .Y(new_n16758));
  xor_4  g14410(.A(new_n16758), .B(new_n6338), .Y(new_n16759));
  xor_4  g14411(.A(new_n16759), .B(new_n16746), .Y(po0187));
  xnor_4 g14412(.A(new_n3869), .B(new_n3868), .Y(po0188));
  xor_4  g14413(.A(pi772), .B(new_n8759), .Y(new_n16762));
  nand_5 g14414(.A(new_n10229), .B(pi332), .Y(new_n16763));
  xor_4  g14415(.A(pi811), .B(new_n10647), .Y(new_n16764));
  nand_5 g14416(.A(new_n8767), .B(pi265), .Y(new_n16765));
  xor_4  g14417(.A(pi804), .B(new_n11101), .Y(new_n16766));
  nand_5 g14418(.A(pi635), .B(new_n8770), .Y(new_n16767));
  xor_4  g14419(.A(pi635), .B(new_n8770), .Y(new_n16768));
  nand_5 g14420(.A(pi545), .B(new_n8773), .Y(new_n16769));
  xor_4  g14421(.A(pi545), .B(new_n8773), .Y(new_n16770));
  nand_5 g14422(.A(new_n10239), .B(pi388), .Y(new_n16771));
  not_8  g14423(.A(new_n16771), .Y(new_n16772));
  xor_4  g14424(.A(pi576), .B(pi388), .Y(new_n16773));
  nand_5 g14425(.A(pi401), .B(new_n8511), .Y(new_n16774));
  nand_5 g14426(.A(new_n8778), .B(pi161), .Y(new_n16775));
  nand_5 g14427(.A(new_n8835), .B(pi281), .Y(new_n16776));
  nand_5 g14428(.A(new_n16776), .B(new_n16775), .Y(new_n16777));
  nand_5 g14429(.A(new_n16777), .B(new_n16774), .Y(new_n16778));
  nor_5  g14430(.A(new_n16778), .B(new_n16773), .Y(new_n16779));
  nor_5  g14431(.A(new_n16779), .B(new_n16772), .Y(new_n16780));
  not_8  g14432(.A(new_n16780), .Y(new_n16781));
  nand_5 g14433(.A(new_n16781), .B(new_n16770), .Y(new_n16782));
  nand_5 g14434(.A(new_n16782), .B(new_n16769), .Y(new_n16783));
  nand_5 g14435(.A(new_n16783), .B(new_n16768), .Y(new_n16784));
  nand_5 g14436(.A(new_n16784), .B(new_n16767), .Y(new_n16785));
  nand_5 g14437(.A(new_n16785), .B(new_n16766), .Y(new_n16786));
  nand_5 g14438(.A(new_n16786), .B(new_n16765), .Y(new_n16787));
  nand_5 g14439(.A(new_n16787), .B(new_n16764), .Y(new_n16788));
  nand_5 g14440(.A(new_n16788), .B(new_n16763), .Y(new_n16789));
  xor_4  g14441(.A(new_n16789), .B(new_n16762), .Y(new_n16790));
  not_8  g14442(.A(new_n16790), .Y(new_n16791));
  nand_5 g14443(.A(new_n16791), .B(pi737), .Y(new_n16792));
  nand_5 g14444(.A(new_n16790), .B(new_n5499), .Y(new_n16793));
  and_6  g14445(.A(new_n16793), .B(new_n16792), .Y(new_n16794));
  xor_4  g14446(.A(new_n16783), .B(new_n16768), .Y(new_n16795));
  xor_4  g14447(.A(new_n16780), .B(new_n16770), .Y(new_n16796));
  nor_5  g14448(.A(new_n16796), .B(pi739), .Y(new_n16797));
  nand_5 g14449(.A(new_n16775), .B(new_n16774), .Y(new_n16798));
  xnor_4 g14450(.A(new_n16798), .B(new_n16776), .Y(new_n16799));
  nand_5 g14451(.A(new_n16799), .B(pi675), .Y(new_n16800));
  nor_5  g14452(.A(new_n16800), .B(new_n5517), .Y(new_n16801));
  xor_4  g14453(.A(new_n16778), .B(new_n16773), .Y(new_n16802));
  xor_4  g14454(.A(new_n16800), .B(new_n5517), .Y(new_n16803));
  not_8  g14455(.A(new_n16803), .Y(new_n16804));
  nor_5  g14456(.A(new_n16804), .B(new_n16802), .Y(new_n16805));
  or_6   g14457(.A(new_n16805), .B(new_n16801), .Y(new_n16806));
  xor_4  g14458(.A(new_n16796), .B(new_n5513), .Y(new_n16807));
  nor_5  g14459(.A(new_n16807), .B(new_n16806), .Y(new_n16808));
  or_6   g14460(.A(new_n16808), .B(new_n16797), .Y(new_n16809));
  nor_5  g14461(.A(new_n16809), .B(new_n16795), .Y(new_n16810));
  xnor_4 g14462(.A(new_n16809), .B(new_n16795), .Y(new_n16811));
  nor_5  g14463(.A(new_n16811), .B(new_n5511), .Y(new_n16812));
  nor_5  g14464(.A(new_n16812), .B(new_n16810), .Y(new_n16813));
  nand_5 g14465(.A(new_n16813), .B(new_n5507), .Y(new_n16814));
  xor_4  g14466(.A(new_n16785), .B(new_n16766), .Y(new_n16815));
  not_8  g14467(.A(new_n16815), .Y(new_n16816));
  xor_4  g14468(.A(new_n16813), .B(pi625), .Y(new_n16817));
  or_6   g14469(.A(new_n16817), .B(new_n16816), .Y(new_n16818));
  nand_5 g14470(.A(new_n16818), .B(new_n16814), .Y(new_n16819));
  nand_5 g14471(.A(new_n16819), .B(new_n5503), .Y(new_n16820));
  xor_4  g14472(.A(new_n16787), .B(new_n16764), .Y(new_n16821));
  xor_4  g14473(.A(new_n16819), .B(new_n5503), .Y(new_n16822));
  nand_5 g14474(.A(new_n16822), .B(new_n16821), .Y(new_n16823));
  nand_5 g14475(.A(new_n16823), .B(new_n16820), .Y(new_n16824));
  xor_4  g14476(.A(new_n16824), .B(new_n16794), .Y(new_n16825));
  not_8  g14477(.A(new_n16825), .Y(new_n16826));
  nor_5  g14478(.A(new_n16826), .B(new_n8225), .Y(new_n16827));
  xor_4  g14479(.A(new_n16825), .B(new_n8225), .Y(new_n16828));
  xor_4  g14480(.A(new_n16822), .B(new_n16821), .Y(new_n16829));
  xor_4  g14481(.A(new_n16817), .B(new_n16816), .Y(new_n16830));
  nor_5  g14482(.A(new_n16830), .B(new_n8261), .Y(new_n16831));
  xor_4  g14483(.A(new_n16807), .B(new_n16806), .Y(new_n16832));
  xor_4  g14484(.A(new_n16799), .B(pi675), .Y(new_n16833));
  xor_4  g14485(.A(pi435), .B(new_n7343), .Y(new_n16834));
  or_6   g14486(.A(new_n16834), .B(new_n2555), .Y(new_n16835));
  not_8  g14487(.A(new_n2554), .Y(new_n16836));
  xor_4  g14488(.A(new_n16834), .B(new_n2555), .Y(new_n16837));
  nand_5 g14489(.A(new_n16837), .B(new_n16836), .Y(new_n16838));
  nand_5 g14490(.A(new_n16838), .B(new_n16835), .Y(new_n16839));
  nand_5 g14491(.A(new_n16839), .B(new_n16833), .Y(new_n16840));
  not_8  g14492(.A(new_n8243), .Y(new_n16841));
  xor_4  g14493(.A(new_n16839), .B(new_n16833), .Y(new_n16842));
  nand_5 g14494(.A(new_n16842), .B(new_n16841), .Y(new_n16843));
  nand_5 g14495(.A(new_n16843), .B(new_n16840), .Y(new_n16844));
  and_6  g14496(.A(new_n16844), .B(new_n8236), .Y(new_n16845));
  xor_4  g14497(.A(new_n16804), .B(new_n16802), .Y(new_n16846));
  not_8  g14498(.A(new_n16846), .Y(new_n16847));
  xor_4  g14499(.A(new_n16844), .B(new_n8237), .Y(new_n16848));
  nor_5  g14500(.A(new_n16848), .B(new_n16847), .Y(new_n16849));
  nor_5  g14501(.A(new_n16849), .B(new_n16845), .Y(new_n16850));
  nand_5 g14502(.A(new_n16850), .B(new_n16832), .Y(new_n16851));
  xnor_4 g14503(.A(new_n16850), .B(new_n16832), .Y(new_n16852));
  or_6   g14504(.A(new_n16852), .B(new_n8255), .Y(new_n16853));
  nand_5 g14505(.A(new_n16853), .B(new_n16851), .Y(new_n16854));
  xor_4  g14506(.A(new_n16811), .B(pi128), .Y(new_n16855));
  nor_5  g14507(.A(new_n16855), .B(new_n16854), .Y(new_n16856));
  xor_4  g14508(.A(new_n16855), .B(new_n16854), .Y(new_n16857));
  nand_5 g14509(.A(new_n16857), .B(new_n8232), .Y(new_n16858));
  not_8  g14510(.A(new_n16858), .Y(new_n16859));
  nor_5  g14511(.A(new_n16859), .B(new_n16856), .Y(new_n16860));
  xor_4  g14512(.A(new_n16830), .B(new_n8261), .Y(new_n16861));
  not_8  g14513(.A(new_n16861), .Y(new_n16862));
  nor_5  g14514(.A(new_n16862), .B(new_n16860), .Y(new_n16863));
  nor_5  g14515(.A(new_n16863), .B(new_n16831), .Y(new_n16864));
  and_6  g14516(.A(new_n16864), .B(new_n16829), .Y(new_n16865));
  xnor_4 g14517(.A(new_n16864), .B(new_n16829), .Y(new_n16866));
  nor_5  g14518(.A(new_n16866), .B(new_n8228), .Y(new_n16867));
  nor_5  g14519(.A(new_n16867), .B(new_n16865), .Y(new_n16868));
  nor_5  g14520(.A(new_n16868), .B(new_n16828), .Y(new_n16869));
  or_6   g14521(.A(new_n16869), .B(new_n16827), .Y(new_n16870));
  xor_4  g14522(.A(pi469), .B(new_n7257), .Y(new_n16871));
  nand_5 g14523(.A(new_n11096), .B(pi123), .Y(new_n16872));
  not_8  g14524(.A(new_n16872), .Y(new_n16873));
  not_8  g14525(.A(new_n16762), .Y(new_n16874));
  nor_5  g14526(.A(new_n16789), .B(new_n16874), .Y(new_n16875));
  nor_5  g14527(.A(new_n16875), .B(new_n16873), .Y(new_n16876));
  xor_4  g14528(.A(new_n16876), .B(new_n16871), .Y(new_n16877));
  nand_5 g14529(.A(new_n16824), .B(new_n16792), .Y(new_n16878));
  nand_5 g14530(.A(new_n16878), .B(new_n16793), .Y(new_n16879));
  or_6   g14531(.A(new_n16879), .B(new_n16877), .Y(new_n16880));
  nand_5 g14532(.A(new_n16879), .B(new_n16877), .Y(new_n16881));
  nand_5 g14533(.A(new_n16881), .B(new_n16880), .Y(new_n16882));
  xor_4  g14534(.A(new_n16882), .B(pi827), .Y(new_n16883));
  xnor_4 g14535(.A(new_n16883), .B(new_n16870), .Y(new_n16884));
  xnor_4 g14536(.A(new_n16884), .B(new_n8222), .Y(po0190));
  xor_4  g14537(.A(pi675), .B(pi401), .Y(new_n16886));
  xor_4  g14538(.A(new_n16886), .B(new_n5522), .Y(new_n16887));
  nand_5 g14539(.A(new_n5595), .B(new_n8835), .Y(new_n16888));
  nand_5 g14540(.A(new_n16888), .B(new_n5597), .Y(new_n16889));
  xor_4  g14541(.A(new_n16889), .B(new_n16887), .Y(new_n16890));
  xnor_4 g14542(.A(new_n16890), .B(new_n6598), .Y(new_n16891));
  not_8  g14543(.A(new_n5763), .Y(new_n16892));
  xor_4  g14544(.A(new_n16834), .B(new_n5598), .Y(new_n16893));
  xor_4  g14545(.A(new_n16893), .B(new_n16892), .Y(po1152));
  nand_5 g14546(.A(po1152), .B(new_n6611), .Y(new_n16895));
  xnor_4 g14547(.A(new_n16895), .B(new_n16891), .Y(po0191));
  not_8  g14548(.A(new_n7456), .Y(new_n16897));
  xor_4  g14549(.A(pi829), .B(new_n6716), .Y(new_n16898));
  nand_5 g14550(.A(pi579), .B(new_n5259), .Y(new_n16899));
  nand_5 g14551(.A(new_n2386), .B(pi483), .Y(new_n16900));
  nand_5 g14552(.A(new_n2389), .B(pi264), .Y(new_n16901));
  xor_4  g14553(.A(pi755), .B(pi264), .Y(new_n16902));
  nand_5 g14554(.A(new_n11371), .B(new_n6766), .Y(new_n16903));
  nand_5 g14555(.A(new_n16903), .B(new_n11370), .Y(new_n16904));
  or_6   g14556(.A(new_n16904), .B(new_n16902), .Y(new_n16905));
  nand_5 g14557(.A(new_n16905), .B(new_n16901), .Y(new_n16906));
  xor_4  g14558(.A(pi749), .B(pi483), .Y(new_n16907));
  not_8  g14559(.A(new_n16907), .Y(new_n16908));
  nand_5 g14560(.A(new_n16908), .B(new_n16906), .Y(new_n16909));
  nand_5 g14561(.A(new_n16909), .B(new_n16900), .Y(new_n16910));
  xor_4  g14562(.A(pi579), .B(pi153), .Y(new_n16911));
  not_8  g14563(.A(new_n16911), .Y(new_n16912));
  nand_5 g14564(.A(new_n16912), .B(new_n16910), .Y(new_n16913));
  nand_5 g14565(.A(new_n16913), .B(new_n16899), .Y(new_n16914));
  xor_4  g14566(.A(new_n16914), .B(new_n16898), .Y(new_n16915));
  xor_4  g14567(.A(new_n16915), .B(new_n16897), .Y(new_n16916));
  xor_4  g14568(.A(new_n16911), .B(new_n16910), .Y(new_n16917));
  nand_5 g14569(.A(new_n16917), .B(new_n7451), .Y(new_n16918));
  xor_4  g14570(.A(new_n16907), .B(new_n16906), .Y(new_n16919));
  not_8  g14571(.A(new_n16919), .Y(new_n16920));
  nor_5  g14572(.A(new_n16920), .B(new_n7419), .Y(new_n16921));
  xor_4  g14573(.A(new_n16920), .B(new_n7419), .Y(new_n16922));
  not_8  g14574(.A(new_n16922), .Y(new_n16923));
  not_8  g14575(.A(new_n7442), .Y(new_n16924));
  xor_4  g14576(.A(new_n16904), .B(new_n16902), .Y(new_n16925));
  nand_5 g14577(.A(new_n16925), .B(new_n16924), .Y(new_n16926));
  xor_4  g14578(.A(new_n16925), .B(new_n16924), .Y(new_n16927));
  xor_4  g14579(.A(new_n11369), .B(new_n6766), .Y(new_n16928));
  nand_5 g14580(.A(new_n16928), .B(po0070), .Y(new_n16929));
  or_6   g14581(.A(new_n16928), .B(new_n7425), .Y(new_n16930));
  nand_5 g14582(.A(new_n16930), .B(new_n16929), .Y(new_n16931));
  nand_5 g14583(.A(new_n16931), .B(new_n16927), .Y(new_n16932));
  nand_5 g14584(.A(new_n16932), .B(new_n16926), .Y(new_n16933));
  nor_5  g14585(.A(new_n16933), .B(new_n16923), .Y(new_n16934));
  or_6   g14586(.A(new_n16934), .B(new_n16921), .Y(new_n16935));
  xnor_4 g14587(.A(new_n16917), .B(new_n7451), .Y(new_n16936));
  not_8  g14588(.A(new_n16936), .Y(new_n16937));
  nand_5 g14589(.A(new_n16937), .B(new_n16935), .Y(new_n16938));
  nand_5 g14590(.A(new_n16938), .B(new_n16918), .Y(new_n16939));
  xor_4  g14591(.A(new_n16939), .B(new_n16916), .Y(po0192));
  not_8  g14592(.A(pi068), .Y(new_n16941));
  xor_4  g14593(.A(pi358), .B(new_n16941), .Y(new_n16942));
  nand_5 g14594(.A(pi687), .B(new_n11899), .Y(new_n16943));
  xor_4  g14595(.A(pi687), .B(new_n11899), .Y(new_n16944));
  nand_5 g14596(.A(new_n2897), .B(pi047), .Y(new_n16945));
  xor_4  g14597(.A(pi239), .B(new_n2855), .Y(new_n16946));
  nand_5 g14598(.A(new_n2932), .B(pi410), .Y(new_n16947));
  not_8  g14599(.A(pi229), .Y(new_n16948));
  nand_5 g14600(.A(new_n16948), .B(pi061), .Y(new_n16949));
  not_8  g14601(.A(new_n14988), .Y(new_n16950));
  nand_5 g14602(.A(new_n16950), .B(new_n14987), .Y(new_n16951));
  nand_5 g14603(.A(new_n16951), .B(new_n16949), .Y(new_n16952));
  xor_4  g14604(.A(pi632), .B(new_n2859), .Y(new_n16953));
  nand_5 g14605(.A(new_n16953), .B(new_n16952), .Y(new_n16954));
  nand_5 g14606(.A(new_n16954), .B(new_n16947), .Y(new_n16955));
  nand_5 g14607(.A(new_n16955), .B(new_n16946), .Y(new_n16956));
  nand_5 g14608(.A(new_n16956), .B(new_n16945), .Y(new_n16957));
  nand_5 g14609(.A(new_n16957), .B(new_n16944), .Y(new_n16958));
  nand_5 g14610(.A(new_n16958), .B(new_n16943), .Y(new_n16959));
  xor_4  g14611(.A(new_n16959), .B(new_n16942), .Y(new_n16960));
  xor_4  g14612(.A(new_n16960), .B(new_n15090), .Y(new_n16961));
  not_8  g14613(.A(new_n15076), .Y(new_n16962));
  xor_4  g14614(.A(new_n16957), .B(new_n16944), .Y(new_n16963));
  nand_5 g14615(.A(new_n16963), .B(new_n16962), .Y(new_n16964));
  xor_4  g14616(.A(new_n16963), .B(new_n15076), .Y(new_n16965));
  not_8  g14617(.A(new_n15058), .Y(new_n16966));
  xor_4  g14618(.A(new_n16955), .B(new_n16946), .Y(new_n16967));
  and_6  g14619(.A(new_n16967), .B(new_n16966), .Y(new_n16968));
  xor_4  g14620(.A(new_n16967), .B(new_n15058), .Y(new_n16969));
  xnor_4 g14621(.A(new_n16953), .B(new_n16952), .Y(new_n16970));
  nor_5  g14622(.A(new_n16970), .B(new_n15041), .Y(new_n16971));
  xor_4  g14623(.A(new_n16970), .B(new_n15042), .Y(new_n16972));
  nand_5 g14624(.A(new_n14989), .B(new_n14983), .Y(new_n16973));
  nand_5 g14625(.A(new_n14991), .B(new_n14970), .Y(new_n16974));
  nand_5 g14626(.A(new_n16974), .B(new_n16973), .Y(new_n16975));
  nor_5  g14627(.A(new_n16975), .B(new_n16972), .Y(new_n16976));
  nor_5  g14628(.A(new_n16976), .B(new_n16971), .Y(new_n16977));
  nor_5  g14629(.A(new_n16977), .B(new_n16969), .Y(new_n16978));
  nor_5  g14630(.A(new_n16978), .B(new_n16968), .Y(new_n16979));
  or_6   g14631(.A(new_n16979), .B(new_n16965), .Y(new_n16980));
  nand_5 g14632(.A(new_n16980), .B(new_n16964), .Y(new_n16981));
  not_8  g14633(.A(new_n16981), .Y(new_n16982));
  xor_4  g14634(.A(new_n16982), .B(new_n16961), .Y(po0193));
  xor_4  g14635(.A(pi809), .B(new_n7471), .Y(new_n16984));
  nand_5 g14636(.A(new_n4724), .B(pi064), .Y(new_n16985));
  nand_5 g14637(.A(new_n3742), .B(new_n3711), .Y(new_n16986));
  nand_5 g14638(.A(new_n16986), .B(new_n16985), .Y(new_n16987));
  xor_4  g14639(.A(new_n16987), .B(new_n16984), .Y(new_n16988));
  xor_4  g14640(.A(new_n16988), .B(pi623), .Y(new_n16989));
  not_8  g14641(.A(new_n3743), .Y(new_n16990));
  nor_5  g14642(.A(new_n3771), .B(new_n16990), .Y(new_n16991));
  nor_5  g14643(.A(new_n3772), .B(pi793), .Y(new_n16992));
  or_6   g14644(.A(new_n16992), .B(new_n16991), .Y(new_n16993));
  xor_4  g14645(.A(new_n16993), .B(new_n16989), .Y(new_n16994));
  nand_5 g14646(.A(new_n3891), .B(new_n12022), .Y(new_n16995));
  or_6   g14647(.A(new_n3892), .B(new_n3773), .Y(new_n16996));
  nand_5 g14648(.A(new_n16996), .B(new_n16995), .Y(new_n16997));
  not_8  g14649(.A(new_n16997), .Y(new_n16998));
  nand_5 g14650(.A(new_n16998), .B(new_n16994), .Y(new_n16999));
  xor_4  g14651(.A(new_n16998), .B(new_n16994), .Y(new_n17000));
  nand_5 g14652(.A(new_n17000), .B(new_n12016), .Y(new_n17001));
  nand_5 g14653(.A(new_n17001), .B(new_n16999), .Y(new_n17002));
  xor_4  g14654(.A(pi607), .B(new_n11934), .Y(new_n17003));
  nand_5 g14655(.A(new_n11901), .B(pi021), .Y(new_n17004));
  nand_5 g14656(.A(new_n16987), .B(new_n16984), .Y(new_n17005));
  nand_5 g14657(.A(new_n17005), .B(new_n17004), .Y(new_n17006));
  xor_4  g14658(.A(new_n17006), .B(new_n17003), .Y(new_n17007));
  not_8  g14659(.A(new_n17007), .Y(new_n17008));
  not_8  g14660(.A(new_n16988), .Y(new_n17009));
  nand_5 g14661(.A(new_n17009), .B(pi623), .Y(new_n17010));
  or_6   g14662(.A(new_n16993), .B(new_n16989), .Y(new_n17011));
  nand_5 g14663(.A(new_n17011), .B(new_n17010), .Y(new_n17012));
  nand_5 g14664(.A(new_n17012), .B(new_n17008), .Y(new_n17013));
  or_6   g14665(.A(new_n17012), .B(new_n17008), .Y(new_n17014));
  nand_5 g14666(.A(new_n17014), .B(new_n17013), .Y(new_n17015));
  xor_4  g14667(.A(new_n17015), .B(new_n4838), .Y(new_n17016));
  xor_4  g14668(.A(new_n17016), .B(new_n12014), .Y(new_n17017));
  xor_4  g14669(.A(new_n17017), .B(new_n17002), .Y(po0194));
  xnor_4 g14670(.A(new_n13090), .B(new_n8530), .Y(po0195));
  or_6   g14671(.A(new_n16448), .B(new_n16446), .Y(new_n17020));
  nand_5 g14672(.A(new_n16454), .B(new_n16449), .Y(new_n17021));
  nand_5 g14673(.A(new_n17021), .B(new_n17020), .Y(new_n17022));
  nor_5  g14674(.A(new_n13215), .B(new_n13208), .Y(new_n17023));
  nor_5  g14675(.A(new_n13238), .B(new_n13217), .Y(new_n17024));
  nor_5  g14676(.A(new_n17024), .B(new_n17023), .Y(new_n17025));
  not_8  g14677(.A(new_n17025), .Y(new_n17026));
  nand_5 g14678(.A(new_n13214), .B(new_n13209), .Y(new_n17027));
  nand_5 g14679(.A(new_n17027), .B(new_n13210), .Y(new_n17028));
  nand_5 g14680(.A(new_n17028), .B(new_n16456), .Y(new_n17029));
  nor_5  g14681(.A(new_n17029), .B(new_n17026), .Y(new_n17030));
  nand_5 g14682(.A(new_n17030), .B(new_n17022), .Y(new_n17031));
  nor_5  g14683(.A(new_n17028), .B(new_n16456), .Y(new_n17032));
  nand_5 g14684(.A(new_n17032), .B(new_n17026), .Y(new_n17033));
  or_6   g14685(.A(new_n17033), .B(new_n17022), .Y(new_n17034));
  nand_5 g14686(.A(new_n17034), .B(new_n17031), .Y(po0196));
  not_8  g14687(.A(new_n8699), .Y(new_n17036));
  nor_5  g14688(.A(new_n8716), .B(new_n17036), .Y(new_n17037));
  nor_5  g14689(.A(new_n8717), .B(new_n8648), .Y(new_n17038));
  or_6   g14690(.A(new_n17038), .B(new_n17037), .Y(new_n17039));
  nand_5 g14691(.A(new_n2454), .B(pi242), .Y(new_n17040));
  or_6   g14692(.A(new_n6666), .B(new_n6665), .Y(new_n17041));
  nand_5 g14693(.A(new_n17041), .B(new_n17040), .Y(new_n17042));
  xor_4  g14694(.A(new_n2413), .B(pi539), .Y(new_n17043));
  xor_4  g14695(.A(new_n17043), .B(new_n17042), .Y(new_n17044));
  not_8  g14696(.A(new_n17044), .Y(new_n17045));
  nor_5  g14697(.A(new_n17045), .B(new_n17039), .Y(new_n17046));
  xor_4  g14698(.A(new_n17044), .B(new_n17039), .Y(new_n17047));
  nand_5 g14699(.A(new_n8698), .B(new_n8691), .Y(new_n17048));
  not_8  g14700(.A(new_n17048), .Y(new_n17049));
  nor_5  g14701(.A(new_n8696), .B(new_n8873), .Y(new_n17050));
  nor_5  g14702(.A(new_n17050), .B(new_n17049), .Y(new_n17051));
  xor_4  g14703(.A(pi792), .B(new_n6716), .Y(new_n17052));
  nand_5 g14704(.A(new_n3227), .B(pi579), .Y(new_n17053));
  nand_5 g14705(.A(new_n8695), .B(new_n8692), .Y(new_n17054));
  nand_5 g14706(.A(new_n17054), .B(new_n17053), .Y(new_n17055));
  xor_4  g14707(.A(new_n17055), .B(new_n17052), .Y(new_n17056));
  xor_4  g14708(.A(new_n17056), .B(pi572), .Y(new_n17057));
  xor_4  g14709(.A(new_n17057), .B(new_n17051), .Y(new_n17058));
  nor_5  g14710(.A(new_n17058), .B(new_n17047), .Y(new_n17059));
  or_6   g14711(.A(new_n17059), .B(new_n17046), .Y(new_n17060));
  or_6   g14712(.A(new_n2413), .B(new_n5648), .Y(new_n17061));
  not_8  g14713(.A(new_n17043), .Y(new_n17062));
  nand_5 g14714(.A(new_n17062), .B(new_n17042), .Y(new_n17063));
  nand_5 g14715(.A(new_n17063), .B(new_n17061), .Y(new_n17064));
  nand_5 g14716(.A(new_n17064), .B(new_n2412), .Y(new_n17065));
  not_8  g14717(.A(new_n17065), .Y(new_n17066));
  nor_5  g14718(.A(new_n17064), .B(new_n2412), .Y(new_n17067));
  nor_5  g14719(.A(new_n17067), .B(new_n17066), .Y(new_n17068));
  xor_4  g14720(.A(new_n17068), .B(new_n6829), .Y(new_n17069));
  nand_5 g14721(.A(new_n17069), .B(new_n17060), .Y(new_n17070));
  not_8  g14722(.A(new_n17069), .Y(new_n17071));
  xor_4  g14723(.A(new_n17071), .B(new_n17060), .Y(new_n17072));
  or_6   g14724(.A(new_n17057), .B(new_n17051), .Y(new_n17073));
  not_8  g14725(.A(new_n17073), .Y(new_n17074));
  nor_5  g14726(.A(new_n17056), .B(new_n6802), .Y(new_n17075));
  nor_5  g14727(.A(new_n17075), .B(new_n17074), .Y(new_n17076));
  xor_4  g14728(.A(pi175), .B(new_n6714), .Y(new_n17077));
  nand_5 g14729(.A(new_n3223), .B(pi615), .Y(new_n17078));
  nand_5 g14730(.A(new_n17055), .B(new_n17052), .Y(new_n17079));
  nand_5 g14731(.A(new_n17079), .B(new_n17078), .Y(new_n17080));
  xor_4  g14732(.A(new_n17080), .B(new_n17077), .Y(new_n17081));
  xor_4  g14733(.A(new_n17081), .B(pi033), .Y(new_n17082));
  xor_4  g14734(.A(new_n17082), .B(new_n17076), .Y(new_n17083));
  or_6   g14735(.A(new_n17083), .B(new_n17072), .Y(new_n17084));
  nand_5 g14736(.A(new_n17084), .B(new_n17070), .Y(new_n17085));
  nor_5  g14737(.A(new_n17067), .B(new_n6829), .Y(new_n17086));
  nor_5  g14738(.A(new_n17086), .B(new_n17066), .Y(new_n17087));
  or_6   g14739(.A(new_n17087), .B(new_n7563), .Y(new_n17088));
  nand_5 g14740(.A(new_n17087), .B(new_n7563), .Y(new_n17089));
  nand_5 g14741(.A(new_n17089), .B(new_n17088), .Y(new_n17090));
  xor_4  g14742(.A(new_n17090), .B(pi377), .Y(new_n17091));
  xnor_4 g14743(.A(new_n17091), .B(new_n17085), .Y(new_n17092));
  or_6   g14744(.A(new_n17082), .B(new_n17076), .Y(new_n17093));
  not_8  g14745(.A(new_n17093), .Y(new_n17094));
  nor_5  g14746(.A(new_n17081), .B(new_n6799), .Y(new_n17095));
  nor_5  g14747(.A(new_n17095), .B(new_n17094), .Y(new_n17096));
  xor_4  g14748(.A(pi105), .B(new_n6787), .Y(new_n17097));
  nand_5 g14749(.A(new_n3218), .B(pi022), .Y(new_n17098));
  nand_5 g14750(.A(new_n17080), .B(new_n17077), .Y(new_n17099));
  nand_5 g14751(.A(new_n17099), .B(new_n17098), .Y(new_n17100));
  xor_4  g14752(.A(new_n17100), .B(new_n17097), .Y(new_n17101));
  xor_4  g14753(.A(new_n17101), .B(pi437), .Y(new_n17102));
  xor_4  g14754(.A(new_n17102), .B(new_n17096), .Y(new_n17103));
  xnor_4 g14755(.A(new_n17103), .B(new_n17092), .Y(po0197));
  not_8  g14756(.A(new_n15102), .Y(new_n17105));
  and_6  g14757(.A(new_n17105), .B(new_n13014), .Y(new_n17106));
  nand_5 g14758(.A(new_n15069), .B(new_n12869), .Y(new_n17107));
  xor_4  g14759(.A(new_n15068), .B(new_n12870), .Y(new_n17108));
  or_6   g14760(.A(new_n15053), .B(new_n12871), .Y(new_n17109));
  nand_5 g14761(.A(new_n15053), .B(new_n12871), .Y(new_n17110));
  nand_5 g14762(.A(new_n15054), .B(new_n12872), .Y(new_n17111));
  nand_5 g14763(.A(new_n15033), .B(new_n12873), .Y(new_n17112));
  nand_5 g14764(.A(new_n14977), .B(new_n12905), .Y(new_n17113));
  xor_4  g14765(.A(new_n14977), .B(new_n12905), .Y(new_n17114));
  nand_5 g14766(.A(new_n12874), .B(new_n4244), .Y(new_n17115));
  xor_4  g14767(.A(new_n12874), .B(new_n4244), .Y(new_n17116));
  nor_5  g14768(.A(new_n12876), .B(new_n4160), .Y(new_n17117));
  xnor_4 g14769(.A(new_n12876), .B(new_n4160), .Y(new_n17118));
  nand_5 g14770(.A(new_n12958), .B(new_n4176), .Y(new_n17119));
  nand_5 g14771(.A(new_n12892), .B(new_n4175), .Y(new_n17120));
  nand_5 g14772(.A(new_n4182), .B(new_n4154), .Y(new_n17121));
  nand_5 g14773(.A(new_n4185), .B(new_n4181), .Y(new_n17122));
  nand_5 g14774(.A(new_n17122), .B(new_n17121), .Y(new_n17123));
  nand_5 g14775(.A(new_n12846), .B(new_n4187), .Y(new_n17124));
  nand_5 g14776(.A(new_n12877), .B(new_n4186), .Y(new_n17125));
  nand_5 g14777(.A(new_n17125), .B(new_n17124), .Y(new_n17126));
  xor_4  g14778(.A(new_n17126), .B(new_n16461), .Y(new_n17127));
  xor_4  g14779(.A(new_n17127), .B(new_n12886), .Y(new_n17128));
  nand_5 g14780(.A(new_n4185), .B(new_n4182), .Y(new_n17129));
  nand_5 g14781(.A(new_n17129), .B(new_n17128), .Y(new_n17130));
  nand_5 g14782(.A(new_n17130), .B(new_n17123), .Y(new_n17131));
  nand_5 g14783(.A(new_n4182), .B(pi385), .Y(new_n17132));
  not_8  g14784(.A(new_n17122), .Y(new_n17133));
  nor_5  g14785(.A(new_n17133), .B(new_n12877), .Y(new_n17134));
  nand_5 g14786(.A(new_n17134), .B(new_n17132), .Y(new_n17135));
  nor_5  g14787(.A(new_n12881), .B(new_n12885), .Y(new_n17136));
  nand_5 g14788(.A(new_n17136), .B(new_n17135), .Y(new_n17137));
  nand_5 g14789(.A(new_n17137), .B(new_n17131), .Y(new_n17138));
  nand_5 g14790(.A(new_n17138), .B(new_n17120), .Y(new_n17139));
  nand_5 g14791(.A(new_n17139), .B(new_n17119), .Y(new_n17140));
  nor_5  g14792(.A(new_n17140), .B(new_n17118), .Y(new_n17141));
  nor_5  g14793(.A(new_n17141), .B(new_n17117), .Y(new_n17142));
  not_8  g14794(.A(new_n17142), .Y(new_n17143));
  nand_5 g14795(.A(new_n17143), .B(new_n17116), .Y(new_n17144));
  nand_5 g14796(.A(new_n17144), .B(new_n17115), .Y(new_n17145));
  nand_5 g14797(.A(new_n17145), .B(new_n17114), .Y(new_n17146));
  nand_5 g14798(.A(new_n17146), .B(new_n17113), .Y(new_n17147));
  nand_5 g14799(.A(new_n17147), .B(new_n17112), .Y(new_n17148));
  nand_5 g14800(.A(new_n17148), .B(new_n17111), .Y(new_n17149));
  nand_5 g14801(.A(new_n17149), .B(new_n17110), .Y(new_n17150));
  nand_5 g14802(.A(new_n17150), .B(new_n17109), .Y(new_n17151));
  nand_5 g14803(.A(new_n17151), .B(new_n17108), .Y(new_n17152));
  nand_5 g14804(.A(new_n17152), .B(new_n17107), .Y(new_n17153));
  nand_5 g14805(.A(new_n17153), .B(new_n15085), .Y(new_n17154));
  nand_5 g14806(.A(new_n17154), .B(new_n13016), .Y(new_n17155));
  nor_5  g14807(.A(new_n17153), .B(new_n15085), .Y(new_n17156));
  not_8  g14808(.A(new_n17156), .Y(new_n17157));
  nand_5 g14809(.A(new_n17157), .B(new_n13020), .Y(new_n17158));
  nand_5 g14810(.A(new_n17158), .B(new_n17155), .Y(new_n17159));
  nand_5 g14811(.A(new_n17157), .B(new_n17154), .Y(new_n17160));
  or_6   g14812(.A(new_n17160), .B(new_n15102), .Y(new_n17161));
  nor_5  g14813(.A(new_n17161), .B(new_n17159), .Y(new_n17162));
  nand_5 g14814(.A(new_n17159), .B(new_n15102), .Y(new_n17163));
  nor_5  g14815(.A(new_n17105), .B(new_n13014), .Y(new_n17164));
  nor_5  g14816(.A(new_n17164), .B(new_n17106), .Y(new_n17165));
  not_8  g14817(.A(new_n17165), .Y(new_n17166));
  nor_5  g14818(.A(new_n17166), .B(new_n17154), .Y(new_n17167));
  nor_5  g14819(.A(new_n17165), .B(new_n17157), .Y(new_n17168));
  nor_5  g14820(.A(new_n17168), .B(new_n17167), .Y(new_n17169));
  nand_5 g14821(.A(new_n17169), .B(new_n17163), .Y(new_n17170));
  nor_5  g14822(.A(new_n17170), .B(new_n17162), .Y(new_n17171));
  not_8  g14823(.A(new_n17171), .Y(new_n17172));
  nor_5  g14824(.A(new_n17172), .B(new_n17106), .Y(new_n17173));
  xor_4  g14825(.A(new_n17160), .B(new_n12868), .Y(new_n17174));
  nand_5 g14826(.A(new_n5914), .B(pi013), .Y(new_n17175));
  xor_4  g14827(.A(pi136), .B(new_n4838), .Y(new_n17176));
  nand_5 g14828(.A(new_n5919), .B(pi623), .Y(new_n17177));
  xor_4  g14829(.A(pi823), .B(new_n4843), .Y(new_n17178));
  nand_5 g14830(.A(pi793), .B(new_n5896), .Y(new_n17179));
  xor_4  g14831(.A(pi793), .B(new_n5896), .Y(new_n17180));
  nand_5 g14832(.A(new_n5891), .B(pi103), .Y(new_n17181));
  xor_4  g14833(.A(pi106), .B(new_n4756), .Y(new_n17182));
  nand_5 g14834(.A(pi298), .B(new_n5842), .Y(new_n17183));
  nand_5 g14835(.A(new_n5845), .B(pi157), .Y(new_n17184));
  xor_4  g14836(.A(pi399), .B(new_n3758), .Y(new_n17185));
  nand_5 g14837(.A(new_n5848), .B(pi241), .Y(new_n17186));
  xor_4  g14838(.A(pi261), .B(pi241), .Y(new_n17187));
  nand_5 g14839(.A(pi753), .B(new_n6018), .Y(new_n17188));
  nand_5 g14840(.A(new_n5852), .B(pi488), .Y(new_n17189));
  nand_5 g14841(.A(new_n17189), .B(new_n3860), .Y(new_n17190));
  nand_5 g14842(.A(new_n17190), .B(new_n17188), .Y(new_n17191));
  or_6   g14843(.A(new_n17191), .B(new_n17187), .Y(new_n17192));
  nand_5 g14844(.A(new_n17192), .B(new_n17186), .Y(new_n17193));
  nand_5 g14845(.A(new_n17193), .B(new_n17185), .Y(new_n17194));
  nand_5 g14846(.A(new_n17194), .B(new_n17184), .Y(new_n17195));
  xor_4  g14847(.A(pi298), .B(pi254), .Y(new_n17196));
  not_8  g14848(.A(new_n17196), .Y(new_n17197));
  nand_5 g14849(.A(new_n17197), .B(new_n17195), .Y(new_n17198));
  nand_5 g14850(.A(new_n17198), .B(new_n17183), .Y(new_n17199));
  nand_5 g14851(.A(new_n17199), .B(new_n17182), .Y(new_n17200));
  nand_5 g14852(.A(new_n17200), .B(new_n17181), .Y(new_n17201));
  nand_5 g14853(.A(new_n17201), .B(new_n17180), .Y(new_n17202));
  nand_5 g14854(.A(new_n17202), .B(new_n17179), .Y(new_n17203));
  nand_5 g14855(.A(new_n17203), .B(new_n17178), .Y(new_n17204));
  nand_5 g14856(.A(new_n17204), .B(new_n17177), .Y(new_n17205));
  nand_5 g14857(.A(new_n17205), .B(new_n17176), .Y(new_n17206));
  nand_5 g14858(.A(new_n17206), .B(new_n17175), .Y(new_n17207));
  xor_4  g14859(.A(pi207), .B(new_n4857), .Y(new_n17208));
  xor_4  g14860(.A(new_n17208), .B(new_n17207), .Y(new_n17209));
  or_6   g14861(.A(new_n17209), .B(new_n17174), .Y(new_n17210));
  xor_4  g14862(.A(new_n17209), .B(new_n17174), .Y(new_n17211));
  xor_4  g14863(.A(new_n17151), .B(new_n17108), .Y(new_n17212));
  xnor_4 g14864(.A(new_n17205), .B(new_n17176), .Y(new_n17213));
  nor_5  g14865(.A(new_n17213), .B(new_n17212), .Y(new_n17214));
  nand_5 g14866(.A(new_n17110), .B(new_n17109), .Y(new_n17215));
  xor_4  g14867(.A(new_n17215), .B(new_n17149), .Y(new_n17216));
  not_8  g14868(.A(new_n17216), .Y(new_n17217));
  xnor_4 g14869(.A(new_n17203), .B(new_n17178), .Y(new_n17218));
  nor_5  g14870(.A(new_n17218), .B(new_n17217), .Y(new_n17219));
  xor_4  g14871(.A(new_n17218), .B(new_n17216), .Y(new_n17220));
  nand_5 g14872(.A(new_n17112), .B(new_n17111), .Y(new_n17221));
  xor_4  g14873(.A(new_n17221), .B(new_n17147), .Y(new_n17222));
  xor_4  g14874(.A(new_n17201), .B(new_n17180), .Y(new_n17223));
  or_6   g14875(.A(new_n17223), .B(new_n17222), .Y(new_n17224));
  xor_4  g14876(.A(new_n17223), .B(new_n17222), .Y(new_n17225));
  xor_4  g14877(.A(new_n17145), .B(new_n17114), .Y(new_n17226));
  xnor_4 g14878(.A(new_n17199), .B(new_n17182), .Y(new_n17227));
  nor_5  g14879(.A(new_n17227), .B(new_n17226), .Y(new_n17228));
  not_8  g14880(.A(new_n17226), .Y(new_n17229));
  xor_4  g14881(.A(new_n17227), .B(new_n17229), .Y(new_n17230));
  xor_4  g14882(.A(new_n17142), .B(new_n17116), .Y(new_n17231));
  not_8  g14883(.A(new_n17231), .Y(new_n17232));
  xor_4  g14884(.A(new_n17196), .B(new_n17195), .Y(new_n17233));
  nand_5 g14885(.A(new_n17233), .B(new_n17232), .Y(new_n17234));
  xor_4  g14886(.A(new_n17233), .B(new_n17232), .Y(new_n17235));
  not_8  g14887(.A(new_n17235), .Y(new_n17236));
  xor_4  g14888(.A(new_n17140), .B(new_n17118), .Y(new_n17237));
  xnor_4 g14889(.A(new_n17193), .B(new_n17185), .Y(new_n17238));
  nor_5  g14890(.A(new_n17238), .B(new_n17237), .Y(new_n17239));
  xnor_4 g14891(.A(new_n17238), .B(new_n17237), .Y(new_n17240));
  nand_5 g14892(.A(new_n17119), .B(new_n17120), .Y(new_n17241));
  xor_4  g14893(.A(new_n17241), .B(new_n17138), .Y(new_n17242));
  xor_4  g14894(.A(new_n17191), .B(new_n17187), .Y(new_n17243));
  not_8  g14895(.A(new_n17243), .Y(new_n17244));
  nand_5 g14896(.A(new_n17244), .B(new_n17242), .Y(new_n17245));
  xor_4  g14897(.A(new_n17244), .B(new_n17242), .Y(new_n17246));
  not_8  g14898(.A(new_n17128), .Y(new_n17247));
  nand_5 g14899(.A(new_n17188), .B(new_n17189), .Y(new_n17248));
  xor_4  g14900(.A(pi631), .B(pi455), .Y(new_n17249));
  not_8  g14901(.A(pi455), .Y(new_n17250));
  xor_4  g14902(.A(new_n12878), .B(new_n4187), .Y(new_n17251));
  xor_4  g14903(.A(new_n17251), .B(new_n17250), .Y(new_n17252));
  nand_5 g14904(.A(new_n17252), .B(new_n17249), .Y(new_n17253));
  xor_4  g14905(.A(new_n17253), .B(new_n17248), .Y(new_n17254));
  nor_5  g14906(.A(new_n17254), .B(new_n17247), .Y(new_n17255));
  nand_5 g14907(.A(new_n3860), .B(new_n17250), .Y(new_n17256));
  not_8  g14908(.A(new_n17251), .Y(new_n17257));
  nand_5 g14909(.A(new_n17249), .B(new_n17257), .Y(new_n17258));
  nand_5 g14910(.A(new_n17258), .B(new_n17256), .Y(new_n17259));
  and_6  g14911(.A(new_n17259), .B(new_n17254), .Y(new_n17260));
  nor_5  g14912(.A(new_n17260), .B(new_n17255), .Y(new_n17261));
  nand_5 g14913(.A(new_n17261), .B(new_n17246), .Y(new_n17262));
  nand_5 g14914(.A(new_n17262), .B(new_n17245), .Y(new_n17263));
  nor_5  g14915(.A(new_n17263), .B(new_n17240), .Y(new_n17264));
  or_6   g14916(.A(new_n17264), .B(new_n17239), .Y(new_n17265));
  or_6   g14917(.A(new_n17265), .B(new_n17236), .Y(new_n17266));
  nand_5 g14918(.A(new_n17266), .B(new_n17234), .Y(new_n17267));
  nor_5  g14919(.A(new_n17267), .B(new_n17230), .Y(new_n17268));
  or_6   g14920(.A(new_n17268), .B(new_n17228), .Y(new_n17269));
  not_8  g14921(.A(new_n17269), .Y(new_n17270));
  nand_5 g14922(.A(new_n17270), .B(new_n17225), .Y(new_n17271));
  nand_5 g14923(.A(new_n17271), .B(new_n17224), .Y(new_n17272));
  nor_5  g14924(.A(new_n17272), .B(new_n17220), .Y(new_n17273));
  or_6   g14925(.A(new_n17273), .B(new_n17219), .Y(new_n17274));
  xor_4  g14926(.A(new_n17213), .B(new_n17212), .Y(new_n17275));
  and_6  g14927(.A(new_n17275), .B(new_n17274), .Y(new_n17276));
  nor_5  g14928(.A(new_n17276), .B(new_n17214), .Y(new_n17277));
  nand_5 g14929(.A(new_n17277), .B(new_n17211), .Y(new_n17278));
  nand_5 g14930(.A(new_n17278), .B(new_n17210), .Y(new_n17279));
  nor_5  g14931(.A(new_n17279), .B(new_n17172), .Y(new_n17280));
  nand_5 g14932(.A(new_n5929), .B(pi097), .Y(new_n17281));
  nand_5 g14933(.A(new_n17208), .B(new_n17207), .Y(new_n17282));
  nand_5 g14934(.A(new_n17282), .B(new_n17281), .Y(new_n17283));
  not_8  g14935(.A(new_n17283), .Y(new_n17284));
  xor_4  g14936(.A(new_n17279), .B(new_n17171), .Y(new_n17285));
  nor_5  g14937(.A(new_n17285), .B(new_n17284), .Y(new_n17286));
  nor_5  g14938(.A(new_n17286), .B(new_n17280), .Y(new_n17287));
  nand_5 g14939(.A(new_n17287), .B(new_n17173), .Y(new_n17288));
  nor_5  g14940(.A(new_n17171), .B(new_n17164), .Y(new_n17289));
  nand_5 g14941(.A(new_n17289), .B(new_n17286), .Y(new_n17290));
  nand_5 g14942(.A(new_n17290), .B(new_n17288), .Y(po0198));
  not_8  g14943(.A(new_n7936), .Y(new_n17292));
  nor_5  g14944(.A(new_n13456), .B(new_n7924), .Y(new_n17293));
  nand_5 g14945(.A(new_n17293), .B(new_n7922), .Y(new_n17294));
  xor_4  g14946(.A(new_n17293), .B(new_n7922), .Y(new_n17295));
  nand_5 g14947(.A(new_n17295), .B(new_n13411), .Y(new_n17296));
  nand_5 g14948(.A(new_n17296), .B(new_n17294), .Y(new_n17297));
  nor_5  g14949(.A(new_n17297), .B(new_n17292), .Y(new_n17298));
  xor_4  g14950(.A(new_n17297), .B(new_n7936), .Y(new_n17299));
  nor_5  g14951(.A(new_n17299), .B(new_n13471), .Y(new_n17300));
  or_6   g14952(.A(new_n17300), .B(new_n17298), .Y(new_n17301));
  nand_5 g14953(.A(new_n17301), .B(new_n13450), .Y(new_n17302));
  xor_4  g14954(.A(new_n17301), .B(new_n13451), .Y(new_n17303));
  or_6   g14955(.A(new_n17303), .B(new_n7945), .Y(new_n17304));
  nand_5 g14956(.A(new_n17304), .B(new_n17302), .Y(new_n17305));
  xor_4  g14957(.A(new_n17305), .B(new_n13432), .Y(new_n17306));
  xor_4  g14958(.A(new_n17306), .B(new_n7917), .Y(po0199));
  not_8  g14959(.A(new_n9163), .Y(new_n17308));
  xor_4  g14960(.A(new_n9164), .B(new_n17308), .Y(po0200));
  nand_5 g14961(.A(new_n14420), .B(new_n13540), .Y(new_n17310));
  nand_5 g14962(.A(new_n17310), .B(new_n13538), .Y(new_n17311));
  xor_4  g14963(.A(new_n17311), .B(new_n13545), .Y(new_n17312));
  nor_5  g14964(.A(new_n17312), .B(new_n14419), .Y(new_n17313));
  nor_5  g14965(.A(new_n14420), .B(new_n13539), .Y(new_n17314));
  nor_5  g14966(.A(new_n17314), .B(new_n13546), .Y(new_n17315));
  nor_5  g14967(.A(new_n17315), .B(new_n17313), .Y(new_n17316));
  or_6   g14968(.A(new_n17316), .B(new_n15517), .Y(new_n17317));
  xor_4  g14969(.A(new_n17316), .B(new_n15517), .Y(new_n17318));
  nand_5 g14970(.A(new_n17318), .B(new_n14417), .Y(new_n17319));
  nand_5 g14971(.A(new_n17319), .B(new_n17317), .Y(new_n17320));
  xor_4  g14972(.A(new_n17320), .B(new_n15509), .Y(new_n17321));
  xor_4  g14973(.A(new_n17321), .B(new_n14408), .Y(po0201));
  xnor_4 g14974(.A(new_n12703), .B(new_n12688), .Y(po0202));
  xnor_4 g14975(.A(new_n13010), .B(new_n12929), .Y(po0203));
  xor_4  g14976(.A(new_n6059), .B(new_n6058), .Y(po0204));
  not_8  g14977(.A(new_n12407), .Y(new_n17326));
  nand_5 g14978(.A(new_n8993), .B(new_n8985), .Y(new_n17327));
  nand_5 g14979(.A(new_n8994), .B(new_n8963), .Y(new_n17328));
  nand_5 g14980(.A(new_n17328), .B(new_n17327), .Y(new_n17329));
  xor_4  g14981(.A(new_n17329), .B(new_n17326), .Y(new_n17330));
  nand_5 g14982(.A(new_n8992), .B(new_n8987), .Y(new_n17331));
  nand_5 g14983(.A(new_n17331), .B(new_n8988), .Y(new_n17332));
  xor_4  g14984(.A(new_n17332), .B(new_n12407), .Y(new_n17333));
  nand_5 g14985(.A(new_n17333), .B(new_n17330), .Y(new_n17334));
  xor_4  g14986(.A(new_n17334), .B(new_n12356), .Y(po0205));
  xor_4  g14987(.A(new_n11636), .B(new_n11635), .Y(po0206));
  xnor_4 g14988(.A(new_n11465), .B(new_n4603), .Y(po0207));
  xor_4  g14989(.A(new_n6532), .B(new_n4575), .Y(po0208));
  xor_4  g14990(.A(new_n9109), .B(new_n9030), .Y(po0209));
  xor_4  g14991(.A(new_n16862), .B(new_n16860), .Y(po0210));
  nand_5 g14992(.A(new_n6935), .B(new_n5454), .Y(new_n17341));
  not_8  g14993(.A(new_n6936), .Y(new_n17342));
  nand_5 g14994(.A(new_n6938), .B(new_n17342), .Y(new_n17343));
  nand_5 g14995(.A(new_n17343), .B(new_n17341), .Y(new_n17344));
  nor_5  g14996(.A(new_n17344), .B(new_n5451), .Y(new_n17345));
  xor_4  g14997(.A(new_n17344), .B(new_n5451), .Y(new_n17346));
  not_8  g14998(.A(new_n17346), .Y(new_n17347));
  nor_5  g14999(.A(new_n17347), .B(new_n11530), .Y(new_n17348));
  or_6   g15000(.A(new_n17348), .B(new_n17345), .Y(new_n17349));
  nand_5 g15001(.A(new_n17349), .B(new_n11557), .Y(new_n17350));
  not_8  g15002(.A(new_n17350), .Y(new_n17351));
  xor_4  g15003(.A(new_n17349), .B(new_n11557), .Y(new_n17352));
  not_8  g15004(.A(new_n17352), .Y(new_n17353));
  xor_4  g15005(.A(new_n17347), .B(new_n11530), .Y(new_n17354));
  not_8  g15006(.A(new_n17354), .Y(new_n17355));
  nor_5  g15007(.A(new_n16341), .B(pi260), .Y(new_n17356));
  nor_5  g15008(.A(new_n16350), .B(new_n16342), .Y(new_n17357));
  nor_5  g15009(.A(new_n17357), .B(new_n17356), .Y(new_n17358));
  nand_5 g15010(.A(new_n11580), .B(new_n11071), .Y(new_n17359));
  not_8  g15011(.A(new_n17359), .Y(new_n17360));
  nand_5 g15012(.A(new_n16346), .B(new_n17360), .Y(new_n17361));
  nand_5 g15013(.A(new_n16349), .B(new_n16343), .Y(new_n17362));
  nor_5  g15014(.A(new_n16346), .B(new_n17360), .Y(new_n17363));
  nand_5 g15015(.A(new_n17363), .B(new_n17362), .Y(new_n17364));
  nand_5 g15016(.A(new_n17364), .B(new_n17361), .Y(new_n17365));
  xor_4  g15017(.A(new_n14697), .B(pi179), .Y(new_n17366));
  xor_4  g15018(.A(new_n17366), .B(new_n17365), .Y(new_n17367));
  xnor_4 g15019(.A(new_n17367), .B(new_n17358), .Y(new_n17368));
  nor_5  g15020(.A(new_n17368), .B(new_n6796), .Y(new_n17369));
  nor_5  g15021(.A(new_n16338), .B(new_n6873), .Y(new_n17370));
  nand_5 g15022(.A(new_n16351), .B(new_n16339), .Y(new_n17371));
  not_8  g15023(.A(new_n17371), .Y(new_n17372));
  nor_5  g15024(.A(new_n17372), .B(new_n17370), .Y(new_n17373));
  xor_4  g15025(.A(new_n17368), .B(new_n6796), .Y(new_n17374));
  not_8  g15026(.A(new_n17374), .Y(new_n17375));
  nor_5  g15027(.A(new_n17375), .B(new_n17373), .Y(new_n17376));
  nor_5  g15028(.A(new_n17376), .B(new_n17369), .Y(new_n17377));
  or_6   g15029(.A(new_n17367), .B(new_n17358), .Y(new_n17378));
  nand_5 g15030(.A(new_n17367), .B(new_n14701), .Y(new_n17379));
  nand_5 g15031(.A(new_n17379), .B(new_n17378), .Y(new_n17380));
  xor_4  g15032(.A(new_n17380), .B(pi794), .Y(new_n17381));
  nand_5 g15033(.A(new_n11588), .B(new_n11505), .Y(new_n17382));
  nand_5 g15034(.A(pi525), .B(pi135), .Y(new_n17383));
  nand_5 g15035(.A(new_n17383), .B(new_n17382), .Y(new_n17384));
  nand_5 g15036(.A(new_n11512), .B(new_n11568), .Y(new_n17385));
  not_8  g15037(.A(new_n17385), .Y(new_n17386));
  nor_5  g15038(.A(new_n17386), .B(new_n17364), .Y(new_n17387));
  nor_5  g15039(.A(new_n11512), .B(new_n11568), .Y(new_n17388));
  nand_5 g15040(.A(new_n17388), .B(new_n17361), .Y(new_n17389));
  nor_5  g15041(.A(new_n17385), .B(new_n17361), .Y(new_n17390));
  not_8  g15042(.A(new_n17390), .Y(new_n17391));
  nand_5 g15043(.A(new_n17391), .B(new_n17389), .Y(new_n17392));
  nor_5  g15044(.A(new_n17392), .B(new_n17387), .Y(new_n17393));
  xnor_4 g15045(.A(new_n17393), .B(new_n17384), .Y(new_n17394));
  xor_4  g15046(.A(new_n17394), .B(new_n17381), .Y(new_n17395));
  nand_5 g15047(.A(new_n17395), .B(new_n17377), .Y(new_n17396));
  xnor_4 g15048(.A(new_n17395), .B(new_n17377), .Y(new_n17397));
  or_6   g15049(.A(new_n17397), .B(new_n6939), .Y(new_n17398));
  nand_5 g15050(.A(new_n17398), .B(new_n17396), .Y(new_n17399));
  nand_5 g15051(.A(new_n17399), .B(new_n17355), .Y(new_n17400));
  nor_5  g15052(.A(new_n17380), .B(new_n14708), .Y(new_n17401));
  nor_5  g15053(.A(new_n17394), .B(new_n17381), .Y(new_n17402));
  nor_5  g15054(.A(new_n17402), .B(new_n17401), .Y(new_n17403));
  nor_5  g15055(.A(new_n17391), .B(new_n17382), .Y(new_n17404));
  not_8  g15056(.A(new_n17404), .Y(new_n17405));
  or_6   g15057(.A(new_n17393), .B(new_n17384), .Y(new_n17406));
  nand_5 g15058(.A(new_n17406), .B(new_n17383), .Y(new_n17407));
  nand_5 g15059(.A(new_n17407), .B(new_n17391), .Y(new_n17408));
  nand_5 g15060(.A(new_n17408), .B(new_n17405), .Y(new_n17409));
  xor_4  g15061(.A(new_n17409), .B(pi243), .Y(new_n17410));
  xor_4  g15062(.A(new_n17410), .B(new_n14725), .Y(new_n17411));
  xnor_4 g15063(.A(new_n17411), .B(new_n17403), .Y(new_n17412));
  xor_4  g15064(.A(new_n17399), .B(new_n17354), .Y(new_n17413));
  or_6   g15065(.A(new_n17413), .B(new_n17412), .Y(new_n17414));
  nand_5 g15066(.A(new_n17414), .B(new_n17400), .Y(new_n17415));
  nand_5 g15067(.A(new_n17415), .B(new_n17353), .Y(new_n17416));
  xor_4  g15068(.A(new_n17415), .B(new_n17352), .Y(new_n17417));
  or_6   g15069(.A(new_n17411), .B(new_n17403), .Y(new_n17418));
  nand_5 g15070(.A(new_n17411), .B(pi788), .Y(new_n17419));
  nand_5 g15071(.A(new_n17419), .B(new_n17418), .Y(new_n17420));
  not_8  g15072(.A(new_n17420), .Y(new_n17421));
  nand_5 g15073(.A(new_n11594), .B(new_n11499), .Y(new_n17422));
  not_8  g15074(.A(new_n17422), .Y(new_n17423));
  nand_5 g15075(.A(new_n17423), .B(new_n17404), .Y(new_n17424));
  nor_5  g15076(.A(new_n17423), .B(new_n17408), .Y(new_n17425));
  nand_5 g15077(.A(pi243), .B(pi148), .Y(new_n17426));
  nor_5  g15078(.A(new_n17426), .B(new_n17404), .Y(new_n17427));
  nor_5  g15079(.A(new_n17427), .B(new_n17425), .Y(new_n17428));
  nand_5 g15080(.A(new_n17428), .B(new_n17424), .Y(new_n17429));
  xor_4  g15081(.A(new_n17429), .B(new_n17421), .Y(new_n17430));
  or_6   g15082(.A(new_n17430), .B(new_n17417), .Y(new_n17431));
  nand_5 g15083(.A(new_n17431), .B(new_n17416), .Y(new_n17432));
  nor_5  g15084(.A(new_n17428), .B(new_n17421), .Y(new_n17433));
  nor_5  g15085(.A(new_n17424), .B(new_n17420), .Y(new_n17434));
  nor_5  g15086(.A(new_n17434), .B(new_n17433), .Y(new_n17435));
  xor_4  g15087(.A(new_n17435), .B(new_n17432), .Y(new_n17436));
  nor_5  g15088(.A(new_n17436), .B(new_n17351), .Y(new_n17437));
  not_8  g15089(.A(new_n17435), .Y(new_n17438));
  nand_5 g15090(.A(new_n17438), .B(new_n17432), .Y(new_n17439));
  nor_5  g15091(.A(new_n17439), .B(new_n17404), .Y(new_n17440));
  or_6   g15092(.A(new_n17440), .B(new_n17437), .Y(po0211));
  nand_5 g15093(.A(new_n13488), .B(new_n13480), .Y(new_n17442));
  or_6   g15094(.A(new_n13489), .B(new_n13429), .Y(new_n17443));
  nand_5 g15095(.A(new_n17443), .B(new_n17442), .Y(new_n17444));
  xor_4  g15096(.A(pi768), .B(new_n8332), .Y(new_n17445));
  nand_5 g15097(.A(new_n13486), .B(new_n13483), .Y(new_n17446));
  nand_5 g15098(.A(new_n17446), .B(new_n13484), .Y(new_n17447));
  xor_4  g15099(.A(new_n17447), .B(new_n17445), .Y(new_n17448));
  nand_5 g15100(.A(new_n17448), .B(new_n17444), .Y(new_n17449));
  nand_5 g15101(.A(pi676), .B(new_n3460), .Y(new_n17450));
  not_8  g15102(.A(new_n13394), .Y(new_n17451));
  nand_5 g15103(.A(new_n17451), .B(new_n13393), .Y(new_n17452));
  nand_5 g15104(.A(new_n17452), .B(new_n17450), .Y(new_n17453));
  xor_4  g15105(.A(pi757), .B(pi752), .Y(new_n17454));
  xor_4  g15106(.A(new_n17454), .B(new_n17453), .Y(new_n17455));
  not_8  g15107(.A(new_n17455), .Y(new_n17456));
  xor_4  g15108(.A(new_n17456), .B(new_n7803), .Y(new_n17457));
  or_6   g15109(.A(new_n13396), .B(new_n7859), .Y(new_n17458));
  nand_5 g15110(.A(new_n13428), .B(new_n13397), .Y(new_n17459));
  nand_5 g15111(.A(new_n17459), .B(new_n17458), .Y(new_n17460));
  xor_4  g15112(.A(new_n17460), .B(new_n17457), .Y(new_n17461));
  xnor_4 g15113(.A(new_n17448), .B(new_n17444), .Y(new_n17462));
  or_6   g15114(.A(new_n17462), .B(new_n17461), .Y(new_n17463));
  nand_5 g15115(.A(new_n17463), .B(new_n17449), .Y(new_n17464));
  or_6   g15116(.A(new_n17456), .B(new_n7803), .Y(new_n17465));
  nand_5 g15117(.A(new_n17460), .B(new_n17457), .Y(new_n17466));
  nand_5 g15118(.A(new_n17466), .B(new_n17465), .Y(new_n17467));
  xor_4  g15119(.A(pi553), .B(new_n4922), .Y(new_n17468));
  nand_5 g15120(.A(new_n4725), .B(pi752), .Y(new_n17469));
  not_8  g15121(.A(new_n17454), .Y(new_n17470));
  nand_5 g15122(.A(new_n17470), .B(new_n17453), .Y(new_n17471));
  nand_5 g15123(.A(new_n17471), .B(new_n17469), .Y(new_n17472));
  xor_4  g15124(.A(new_n17472), .B(new_n17468), .Y(new_n17473));
  xor_4  g15125(.A(new_n17473), .B(new_n7798), .Y(new_n17474));
  xor_4  g15126(.A(new_n17474), .B(new_n17467), .Y(new_n17475));
  not_8  g15127(.A(new_n17475), .Y(new_n17476));
  nand_5 g15128(.A(pi768), .B(new_n8332), .Y(new_n17477));
  nand_5 g15129(.A(new_n17447), .B(new_n17445), .Y(new_n17478));
  nand_5 g15130(.A(new_n17478), .B(new_n17477), .Y(new_n17479));
  xor_4  g15131(.A(pi671), .B(pi180), .Y(new_n17480));
  xor_4  g15132(.A(new_n17480), .B(new_n17479), .Y(new_n17481));
  xor_4  g15133(.A(new_n17481), .B(new_n17476), .Y(new_n17482));
  xnor_4 g15134(.A(new_n17482), .B(new_n17464), .Y(po0212));
  not_8  g15135(.A(pi663), .Y(new_n17484));
  xor_4  g15136(.A(pi697), .B(new_n17484), .Y(new_n17485));
  nand_5 g15137(.A(pi835), .B(new_n7533), .Y(new_n17486));
  xor_4  g15138(.A(pi835), .B(new_n7533), .Y(new_n17487));
  nand_5 g15139(.A(pi380), .B(new_n7751), .Y(new_n17488));
  not_8  g15140(.A(new_n15981), .Y(new_n17489));
  nand_5 g15141(.A(new_n17489), .B(new_n15980), .Y(new_n17490));
  nand_5 g15142(.A(new_n17490), .B(new_n17488), .Y(new_n17491));
  nand_5 g15143(.A(new_n17491), .B(new_n17487), .Y(new_n17492));
  nand_5 g15144(.A(new_n17492), .B(new_n17486), .Y(new_n17493));
  xor_4  g15145(.A(new_n17493), .B(new_n17485), .Y(new_n17494));
  not_8  g15146(.A(new_n17494), .Y(new_n17495));
  xnor_4 g15147(.A(new_n17491), .B(new_n17487), .Y(new_n17496));
  nor_5  g15148(.A(new_n9597), .B(new_n9591), .Y(new_n17497));
  not_8  g15149(.A(new_n9598), .Y(new_n17498));
  nor_5  g15150(.A(new_n9603), .B(new_n17498), .Y(new_n17499));
  or_6   g15151(.A(new_n17499), .B(new_n17497), .Y(new_n17500));
  nand_5 g15152(.A(new_n17500), .B(new_n14505), .Y(new_n17501));
  xor_4  g15153(.A(new_n17500), .B(new_n14505), .Y(new_n17502));
  nand_5 g15154(.A(new_n17502), .B(new_n10789), .Y(new_n17503));
  nand_5 g15155(.A(new_n17503), .B(new_n17501), .Y(new_n17504));
  nand_5 g15156(.A(new_n17504), .B(new_n14503), .Y(new_n17505));
  xor_4  g15157(.A(new_n17504), .B(new_n14527), .Y(new_n17506));
  not_8  g15158(.A(new_n17506), .Y(new_n17507));
  nand_5 g15159(.A(new_n17507), .B(new_n10764), .Y(new_n17508));
  nand_5 g15160(.A(new_n17508), .B(new_n17505), .Y(new_n17509));
  nand_5 g15161(.A(new_n17509), .B(new_n14499), .Y(new_n17510));
  xor_4  g15162(.A(new_n17509), .B(new_n14500), .Y(new_n17511));
  not_8  g15163(.A(new_n17511), .Y(new_n17512));
  nand_5 g15164(.A(new_n17512), .B(new_n10737), .Y(new_n17513));
  nand_5 g15165(.A(new_n17513), .B(new_n17510), .Y(new_n17514));
  nor_5  g15166(.A(new_n17514), .B(new_n14497), .Y(new_n17515));
  not_8  g15167(.A(new_n14497), .Y(new_n17516));
  xor_4  g15168(.A(new_n17514), .B(new_n17516), .Y(new_n17517));
  nor_5  g15169(.A(new_n17517), .B(new_n15983), .Y(new_n17518));
  or_6   g15170(.A(new_n17518), .B(new_n17515), .Y(new_n17519));
  nand_5 g15171(.A(new_n17519), .B(new_n17496), .Y(new_n17520));
  xnor_4 g15172(.A(new_n17519), .B(new_n17496), .Y(new_n17521));
  or_6   g15173(.A(new_n17521), .B(new_n14626), .Y(new_n17522));
  nand_5 g15174(.A(new_n17522), .B(new_n17520), .Y(new_n17523));
  nand_5 g15175(.A(new_n4873), .B(pi121), .Y(new_n17524));
  nand_5 g15176(.A(pi124), .B(new_n7700), .Y(new_n17525));
  and_6  g15177(.A(new_n17525), .B(new_n17524), .Y(new_n17526));
  nand_5 g15178(.A(new_n4930), .B(pi066), .Y(new_n17527));
  nand_5 g15179(.A(new_n14625), .B(new_n14622), .Y(new_n17528));
  nand_5 g15180(.A(new_n17528), .B(new_n17527), .Y(new_n17529));
  xor_4  g15181(.A(new_n17529), .B(new_n17526), .Y(new_n17530));
  xor_4  g15182(.A(new_n17530), .B(new_n17523), .Y(new_n17531));
  xor_4  g15183(.A(new_n17531), .B(new_n17495), .Y(new_n17532));
  nand_5 g15184(.A(new_n15546), .B(pi315), .Y(new_n17533));
  nand_5 g15185(.A(pi713), .B(new_n4858), .Y(new_n17534));
  nand_5 g15186(.A(new_n17534), .B(new_n17533), .Y(new_n17535));
  nand_5 g15187(.A(new_n4839), .B(pi341), .Y(new_n17536));
  xor_4  g15188(.A(pi812), .B(new_n9210), .Y(new_n17537));
  nand_5 g15189(.A(new_n4842), .B(pi203), .Y(new_n17538));
  xor_4  g15190(.A(pi547), .B(new_n9213), .Y(new_n17539));
  nand_5 g15191(.A(pi451), .B(new_n4754), .Y(new_n17540));
  xor_4  g15192(.A(pi451), .B(new_n4754), .Y(new_n17541));
  nand_5 g15193(.A(new_n4757), .B(pi363), .Y(new_n17542));
  xor_4  g15194(.A(pi375), .B(new_n9220), .Y(new_n17543));
  nand_5 g15195(.A(new_n4760), .B(pi104), .Y(new_n17544));
  xor_4  g15196(.A(pi427), .B(new_n9223), .Y(new_n17545));
  nand_5 g15197(.A(pi343), .B(new_n4763), .Y(new_n17546));
  nand_5 g15198(.A(new_n15238), .B(new_n15228), .Y(new_n17547));
  nand_5 g15199(.A(new_n17547), .B(new_n17546), .Y(new_n17548));
  nand_5 g15200(.A(new_n17548), .B(new_n17545), .Y(new_n17549));
  nand_5 g15201(.A(new_n17549), .B(new_n17544), .Y(new_n17550));
  nand_5 g15202(.A(new_n17550), .B(new_n17543), .Y(new_n17551));
  nand_5 g15203(.A(new_n17551), .B(new_n17542), .Y(new_n17552));
  nand_5 g15204(.A(new_n17552), .B(new_n17541), .Y(new_n17553));
  nand_5 g15205(.A(new_n17553), .B(new_n17540), .Y(new_n17554));
  nand_5 g15206(.A(new_n17554), .B(new_n17539), .Y(new_n17555));
  nand_5 g15207(.A(new_n17555), .B(new_n17538), .Y(new_n17556));
  nand_5 g15208(.A(new_n17556), .B(new_n17537), .Y(new_n17557));
  nand_5 g15209(.A(new_n17557), .B(new_n17536), .Y(new_n17558));
  xnor_4 g15210(.A(new_n17558), .B(new_n17535), .Y(new_n17559));
  xor_4  g15211(.A(new_n17559), .B(new_n17532), .Y(new_n17560));
  xor_4  g15212(.A(new_n17556), .B(new_n17537), .Y(new_n17561));
  xnor_4 g15213(.A(new_n17521), .B(new_n14626), .Y(new_n17562));
  or_6   g15214(.A(new_n17562), .B(new_n17561), .Y(new_n17563));
  xor_4  g15215(.A(new_n17562), .B(new_n17561), .Y(new_n17564));
  xor_4  g15216(.A(new_n17517), .B(new_n15983), .Y(new_n17565));
  xnor_4 g15217(.A(new_n17554), .B(new_n17539), .Y(new_n17566));
  nand_5 g15218(.A(new_n17566), .B(new_n17565), .Y(new_n17567));
  xor_4  g15219(.A(new_n17566), .B(new_n17565), .Y(new_n17568));
  xor_4  g15220(.A(new_n17552), .B(new_n17541), .Y(new_n17569));
  xor_4  g15221(.A(new_n17511), .B(new_n10737), .Y(new_n17570));
  not_8  g15222(.A(new_n17570), .Y(new_n17571));
  or_6   g15223(.A(new_n17571), .B(new_n17569), .Y(new_n17572));
  xor_4  g15224(.A(new_n17571), .B(new_n17569), .Y(new_n17573));
  xor_4  g15225(.A(new_n17550), .B(new_n17543), .Y(new_n17574));
  not_8  g15226(.A(new_n17574), .Y(new_n17575));
  xor_4  g15227(.A(new_n17506), .B(new_n10764), .Y(new_n17576));
  nand_5 g15228(.A(new_n17576), .B(new_n17575), .Y(new_n17577));
  xor_4  g15229(.A(new_n17576), .B(new_n17575), .Y(new_n17578));
  xor_4  g15230(.A(new_n17548), .B(new_n17545), .Y(new_n17579));
  not_8  g15231(.A(new_n17579), .Y(new_n17580));
  xor_4  g15232(.A(new_n17502), .B(new_n10790), .Y(new_n17581));
  nor_5  g15233(.A(new_n17581), .B(new_n17580), .Y(new_n17582));
  xor_4  g15234(.A(new_n17581), .B(new_n17579), .Y(new_n17583));
  not_8  g15235(.A(new_n15239), .Y(new_n17584));
  nor_5  g15236(.A(new_n17584), .B(new_n9604), .Y(new_n17585));
  or_6   g15237(.A(new_n15241), .B(new_n9620), .Y(new_n17586));
  nor_5  g15238(.A(new_n15245), .B(new_n9629), .Y(new_n17587));
  nand_5 g15239(.A(new_n17587), .B(new_n15249), .Y(new_n17588));
  not_8  g15240(.A(new_n9624), .Y(new_n17589));
  xor_4  g15241(.A(new_n17587), .B(new_n15249), .Y(new_n17590));
  nand_5 g15242(.A(new_n17590), .B(new_n17589), .Y(new_n17591));
  nand_5 g15243(.A(new_n17591), .B(new_n17588), .Y(new_n17592));
  xor_4  g15244(.A(new_n15241), .B(new_n9620), .Y(new_n17593));
  nand_5 g15245(.A(new_n17593), .B(new_n17592), .Y(new_n17594));
  nand_5 g15246(.A(new_n17594), .B(new_n17586), .Y(new_n17595));
  xor_4  g15247(.A(new_n15239), .B(new_n9604), .Y(new_n17596));
  nor_5  g15248(.A(new_n17596), .B(new_n17595), .Y(new_n17597));
  nor_5  g15249(.A(new_n17597), .B(new_n17585), .Y(new_n17598));
  nor_5  g15250(.A(new_n17598), .B(new_n17583), .Y(new_n17599));
  nor_5  g15251(.A(new_n17599), .B(new_n17582), .Y(new_n17600));
  nand_5 g15252(.A(new_n17600), .B(new_n17578), .Y(new_n17601));
  nand_5 g15253(.A(new_n17601), .B(new_n17577), .Y(new_n17602));
  nand_5 g15254(.A(new_n17602), .B(new_n17573), .Y(new_n17603));
  nand_5 g15255(.A(new_n17603), .B(new_n17572), .Y(new_n17604));
  nand_5 g15256(.A(new_n17604), .B(new_n17568), .Y(new_n17605));
  nand_5 g15257(.A(new_n17605), .B(new_n17567), .Y(new_n17606));
  nand_5 g15258(.A(new_n17606), .B(new_n17564), .Y(new_n17607));
  nand_5 g15259(.A(new_n17607), .B(new_n17563), .Y(new_n17608));
  xor_4  g15260(.A(new_n17608), .B(new_n17560), .Y(po0213));
  or_6   g15261(.A(new_n10716), .B(new_n4842), .Y(new_n17610));
  nand_5 g15262(.A(new_n10716), .B(new_n4842), .Y(new_n17611));
  and_6  g15263(.A(new_n17611), .B(new_n17610), .Y(new_n17612));
  nand_5 g15264(.A(new_n13165), .B(pi427), .Y(new_n17613));
  nand_5 g15265(.A(new_n17613), .B(new_n13166), .Y(new_n17614));
  nand_5 g15266(.A(new_n17614), .B(new_n10684), .Y(new_n17615));
  or_6   g15267(.A(new_n17614), .B(new_n10684), .Y(new_n17616));
  nand_5 g15268(.A(new_n17616), .B(pi375), .Y(new_n17617));
  nand_5 g15269(.A(new_n17617), .B(new_n17615), .Y(new_n17618));
  nor_5  g15270(.A(new_n17618), .B(pi236), .Y(new_n17619));
  xor_4  g15271(.A(new_n17618), .B(pi236), .Y(new_n17620));
  not_8  g15272(.A(new_n17620), .Y(new_n17621));
  nor_5  g15273(.A(new_n17621), .B(new_n10700), .Y(new_n17622));
  or_6   g15274(.A(new_n17622), .B(new_n17619), .Y(new_n17623));
  xor_4  g15275(.A(new_n17623), .B(new_n17612), .Y(new_n17624));
  and_6  g15276(.A(new_n17616), .B(new_n17615), .Y(new_n17625));
  xor_4  g15277(.A(new_n17625), .B(new_n4757), .Y(new_n17626));
  nor_5  g15278(.A(new_n8615), .B(new_n6612), .Y(new_n17627));
  or_6   g15279(.A(new_n17627), .B(new_n6608), .Y(new_n17628));
  xor_4  g15280(.A(new_n17627), .B(new_n6607), .Y(new_n17629));
  or_6   g15281(.A(new_n17629), .B(new_n8621), .Y(new_n17630));
  nand_5 g15282(.A(new_n17630), .B(new_n17628), .Y(new_n17631));
  and_6  g15283(.A(new_n17631), .B(new_n8605), .Y(new_n17632));
  xor_4  g15284(.A(new_n17631), .B(new_n8604), .Y(new_n17633));
  nor_5  g15285(.A(new_n17633), .B(new_n6628), .Y(new_n17634));
  nor_5  g15286(.A(new_n17634), .B(new_n17632), .Y(new_n17635));
  nand_5 g15287(.A(new_n17635), .B(new_n6648), .Y(new_n17636));
  or_6   g15288(.A(new_n17635), .B(new_n6648), .Y(new_n17637));
  nand_5 g15289(.A(new_n17637), .B(new_n8600), .Y(new_n17638));
  nand_5 g15290(.A(new_n17638), .B(new_n17636), .Y(new_n17639));
  nor_5  g15291(.A(new_n17639), .B(new_n13169), .Y(new_n17640));
  xor_4  g15292(.A(new_n17639), .B(new_n13168), .Y(new_n17641));
  nor_5  g15293(.A(new_n17641), .B(new_n8598), .Y(new_n17642));
  or_6   g15294(.A(new_n17642), .B(new_n17640), .Y(new_n17643));
  nor_5  g15295(.A(new_n17643), .B(new_n17626), .Y(new_n17644));
  not_8  g15296(.A(new_n17626), .Y(new_n17645));
  xor_4  g15297(.A(new_n17643), .B(new_n17645), .Y(new_n17646));
  nor_5  g15298(.A(new_n17646), .B(new_n8636), .Y(new_n17647));
  or_6   g15299(.A(new_n17647), .B(new_n17644), .Y(new_n17648));
  nand_5 g15300(.A(new_n17648), .B(new_n8575), .Y(new_n17649));
  xor_4  g15301(.A(new_n17621), .B(new_n10700), .Y(new_n17650));
  xor_4  g15302(.A(new_n17648), .B(new_n16425), .Y(new_n17651));
  or_6   g15303(.A(new_n17651), .B(new_n17650), .Y(new_n17652));
  nand_5 g15304(.A(new_n17652), .B(new_n17649), .Y(new_n17653));
  xor_4  g15305(.A(new_n17653), .B(new_n17624), .Y(new_n17654));
  xor_4  g15306(.A(new_n17654), .B(new_n16390), .Y(po0214));
  xnor_4 g15307(.A(new_n10808), .B(new_n10805), .Y(po0215));
  nand_5 g15308(.A(new_n17014), .B(pi013), .Y(new_n17657));
  nand_5 g15309(.A(new_n17657), .B(new_n17013), .Y(new_n17658));
  not_8  g15310(.A(pi323), .Y(new_n17659));
  xor_4  g15311(.A(pi381), .B(new_n17659), .Y(new_n17660));
  nand_5 g15312(.A(pi607), .B(new_n11934), .Y(new_n17661));
  nand_5 g15313(.A(new_n17006), .B(new_n17003), .Y(new_n17662));
  nand_5 g15314(.A(new_n17662), .B(new_n17661), .Y(new_n17663));
  xnor_4 g15315(.A(new_n17663), .B(new_n17660), .Y(new_n17664));
  nand_5 g15316(.A(new_n17664), .B(new_n17658), .Y(new_n17665));
  nor_5  g15317(.A(new_n17664), .B(new_n17658), .Y(new_n17666));
  not_8  g15318(.A(new_n17666), .Y(new_n17667));
  nand_5 g15319(.A(new_n17667), .B(new_n17665), .Y(new_n17668));
  xor_4  g15320(.A(new_n17668), .B(new_n4857), .Y(new_n17669));
  xnor_4 g15321(.A(new_n17669), .B(new_n12011), .Y(new_n17670));
  nand_5 g15322(.A(new_n17016), .B(new_n12014), .Y(new_n17671));
  nand_5 g15323(.A(new_n17017), .B(new_n17002), .Y(new_n17672));
  nand_5 g15324(.A(new_n17672), .B(new_n17671), .Y(new_n17673));
  xnor_4 g15325(.A(new_n17673), .B(new_n17670), .Y(po0216));
  xor_4  g15326(.A(new_n6921), .B(new_n6887), .Y(po0217));
  nand_5 g15327(.A(new_n16606), .B(new_n5855), .Y(new_n17676));
  nor_5  g15328(.A(new_n16605), .B(new_n13253), .Y(new_n17677));
  nor_5  g15329(.A(new_n17677), .B(new_n5857), .Y(new_n17678));
  nand_5 g15330(.A(new_n17678), .B(new_n17676), .Y(new_n17679));
  xor_4  g15331(.A(new_n17679), .B(new_n13262), .Y(new_n17680));
  xor_4  g15332(.A(new_n17680), .B(new_n13553), .Y(new_n17681));
  nand_5 g15333(.A(new_n16601), .B(new_n16598), .Y(new_n17682));
  or_6   g15334(.A(new_n16607), .B(new_n16602), .Y(new_n17683));
  nand_5 g15335(.A(new_n17683), .B(new_n17682), .Y(new_n17684));
  xor_4  g15336(.A(new_n17684), .B(new_n4996), .Y(new_n17685));
  xor_4  g15337(.A(new_n17685), .B(new_n17681), .Y(po0218));
  xor_4  g15338(.A(new_n11283), .B(new_n11282), .Y(po0219));
  xor_4  g15339(.A(new_n13200), .B(new_n3756), .Y(po0220));
  not_8  g15340(.A(new_n10970), .Y(new_n17689));
  not_8  g15341(.A(new_n10907), .Y(new_n17690));
  nand_5 g15342(.A(new_n10856), .B(pi762), .Y(new_n17691));
  nand_5 g15343(.A(new_n16506), .B(new_n16499), .Y(new_n17692));
  nand_5 g15344(.A(new_n17692), .B(new_n17691), .Y(new_n17693));
  nand_5 g15345(.A(new_n17693), .B(new_n10898), .Y(new_n17694));
  or_6   g15346(.A(new_n17693), .B(new_n10898), .Y(new_n17695));
  nand_5 g15347(.A(new_n17695), .B(pi440), .Y(new_n17696));
  nand_5 g15348(.A(new_n17696), .B(new_n17694), .Y(new_n17697));
  or_6   g15349(.A(new_n17697), .B(new_n17690), .Y(new_n17698));
  nand_5 g15350(.A(new_n17698), .B(pi193), .Y(new_n17699));
  nand_5 g15351(.A(new_n17697), .B(new_n17690), .Y(new_n17700));
  nand_5 g15352(.A(new_n17700), .B(new_n17699), .Y(new_n17701));
  nand_5 g15353(.A(new_n17701), .B(new_n17689), .Y(new_n17702));
  not_8  g15354(.A(new_n17702), .Y(new_n17703));
  not_8  g15355(.A(pi057), .Y(new_n17704));
  nor_5  g15356(.A(new_n17701), .B(new_n17689), .Y(new_n17705));
  nor_5  g15357(.A(new_n17705), .B(new_n17704), .Y(new_n17706));
  nor_5  g15358(.A(new_n17706), .B(new_n17703), .Y(new_n17707));
  nand_5 g15359(.A(new_n13053), .B(new_n9207), .Y(new_n17708));
  nand_5 g15360(.A(new_n10969), .B(new_n10964), .Y(new_n17709));
  nand_5 g15361(.A(new_n17709), .B(new_n17708), .Y(new_n17710));
  xor_4  g15362(.A(new_n17710), .B(new_n17707), .Y(new_n17711));
  nand_5 g15363(.A(new_n17700), .B(new_n17698), .Y(new_n17712));
  xor_4  g15364(.A(new_n17712), .B(pi193), .Y(new_n17713));
  not_8  g15365(.A(new_n17713), .Y(new_n17714));
  nand_5 g15366(.A(new_n17714), .B(new_n10134), .Y(new_n17715));
  nand_5 g15367(.A(new_n17713), .B(new_n10133), .Y(new_n17716));
  and_6  g15368(.A(new_n17695), .B(new_n17694), .Y(new_n17717));
  xor_4  g15369(.A(new_n17717), .B(pi440), .Y(new_n17718));
  nand_5 g15370(.A(new_n17718), .B(new_n10089), .Y(new_n17719));
  not_8  g15371(.A(new_n17719), .Y(new_n17720));
  nand_5 g15372(.A(new_n16518), .B(new_n16508), .Y(new_n17721));
  nand_5 g15373(.A(new_n16519), .B(new_n10049), .Y(new_n17722));
  nand_5 g15374(.A(new_n17722), .B(new_n17721), .Y(new_n17723));
  xnor_4 g15375(.A(new_n17718), .B(new_n10089), .Y(new_n17724));
  nor_5  g15376(.A(new_n17724), .B(new_n17723), .Y(new_n17725));
  nor_5  g15377(.A(new_n17725), .B(new_n17720), .Y(new_n17726));
  not_8  g15378(.A(new_n17726), .Y(new_n17727));
  nand_5 g15379(.A(new_n17727), .B(new_n17716), .Y(new_n17728));
  nand_5 g15380(.A(new_n17728), .B(new_n17715), .Y(new_n17729));
  nand_5 g15381(.A(new_n17729), .B(new_n10181), .Y(new_n17730));
  or_6   g15382(.A(new_n17729), .B(new_n10181), .Y(new_n17731));
  or_6   g15383(.A(new_n17705), .B(new_n17703), .Y(new_n17732));
  xor_4  g15384(.A(new_n17732), .B(pi057), .Y(new_n17733));
  not_8  g15385(.A(new_n17733), .Y(new_n17734));
  nand_5 g15386(.A(new_n17734), .B(new_n17731), .Y(new_n17735));
  nand_5 g15387(.A(new_n17735), .B(new_n17730), .Y(new_n17736));
  xor_4  g15388(.A(new_n17736), .B(new_n17711), .Y(new_n17737));
  xnor_4 g15389(.A(new_n17737), .B(new_n10219), .Y(po0221));
  xnor_4 g15390(.A(new_n14968), .B(new_n14948), .Y(po0222));
  nand_5 g15391(.A(new_n17081), .B(pi033), .Y(new_n17740));
  nand_5 g15392(.A(new_n17056), .B(pi572), .Y(new_n17741));
  nand_5 g15393(.A(new_n8696), .B(pi587), .Y(new_n17742));
  not_8  g15394(.A(pi779), .Y(new_n17743));
  nand_5 g15395(.A(new_n8661), .B(new_n17743), .Y(new_n17744));
  nand_5 g15396(.A(new_n8653), .B(pi837), .Y(new_n17745));
  and_6  g15397(.A(new_n8670), .B(new_n8654), .Y(new_n17746));
  nand_5 g15398(.A(new_n17746), .B(new_n17745), .Y(new_n17747));
  nor_5  g15399(.A(new_n8653), .B(pi837), .Y(new_n17748));
  nor_5  g15400(.A(new_n17748), .B(new_n8681), .Y(new_n17749));
  nand_5 g15401(.A(new_n17749), .B(new_n17747), .Y(new_n17750));
  nand_5 g15402(.A(new_n17750), .B(new_n8665), .Y(new_n17751));
  nand_5 g15403(.A(new_n17751), .B(new_n8666), .Y(new_n17752));
  nand_5 g15404(.A(new_n17752), .B(new_n8688), .Y(new_n17753));
  nand_5 g15405(.A(new_n17753), .B(new_n17744), .Y(new_n17754));
  or_6   g15406(.A(new_n17754), .B(new_n8698), .Y(new_n17755));
  nand_5 g15407(.A(new_n17755), .B(new_n17742), .Y(new_n17756));
  nand_5 g15408(.A(new_n17756), .B(new_n17057), .Y(new_n17757));
  nand_5 g15409(.A(new_n17757), .B(new_n17741), .Y(new_n17758));
  nand_5 g15410(.A(new_n17758), .B(new_n17082), .Y(new_n17759));
  nand_5 g15411(.A(new_n17759), .B(new_n17740), .Y(new_n17760));
  xnor_4 g15412(.A(new_n17760), .B(new_n17102), .Y(new_n17761));
  xor_4  g15413(.A(new_n17758), .B(new_n17082), .Y(new_n17762));
  not_8  g15414(.A(new_n17762), .Y(new_n17763));
  xor_4  g15415(.A(new_n17756), .B(new_n17057), .Y(new_n17764));
  or_6   g15416(.A(new_n17764), .B(new_n12292), .Y(new_n17765));
  xor_4  g15417(.A(new_n17764), .B(new_n12292), .Y(new_n17766));
  xor_4  g15418(.A(new_n17754), .B(new_n8698), .Y(new_n17767));
  not_8  g15419(.A(new_n17767), .Y(new_n17768));
  xor_4  g15420(.A(new_n17752), .B(new_n8689), .Y(new_n17769));
  not_8  g15421(.A(new_n12252), .Y(new_n17770));
  nand_5 g15422(.A(new_n12260), .B(new_n8678), .Y(new_n17771));
  nand_5 g15423(.A(new_n12258), .B(pi708), .Y(new_n17772));
  nand_5 g15424(.A(new_n17772), .B(new_n17771), .Y(new_n17773));
  xor_4  g15425(.A(new_n17773), .B(new_n8674), .Y(new_n17774));
  or_6   g15426(.A(new_n17774), .B(new_n17770), .Y(new_n17775));
  or_6   g15427(.A(new_n12258), .B(new_n8703), .Y(new_n17776));
  nand_5 g15428(.A(new_n17776), .B(new_n17774), .Y(new_n17777));
  nand_5 g15429(.A(new_n17777), .B(new_n17775), .Y(new_n17778));
  xor_4  g15430(.A(new_n17750), .B(new_n8667), .Y(new_n17779));
  nand_5 g15431(.A(new_n17779), .B(new_n17778), .Y(new_n17780));
  or_6   g15432(.A(new_n17779), .B(new_n17778), .Y(new_n17781));
  nand_5 g15433(.A(new_n17781), .B(new_n12273), .Y(new_n17782));
  nand_5 g15434(.A(new_n17782), .B(new_n17780), .Y(new_n17783));
  or_6   g15435(.A(new_n17783), .B(new_n17769), .Y(new_n17784));
  xor_4  g15436(.A(new_n17783), .B(new_n17769), .Y(new_n17785));
  nand_5 g15437(.A(new_n17785), .B(new_n12278), .Y(new_n17786));
  nand_5 g15438(.A(new_n17786), .B(new_n17784), .Y(new_n17787));
  nor_5  g15439(.A(new_n17787), .B(new_n17768), .Y(new_n17788));
  xor_4  g15440(.A(new_n17787), .B(new_n17767), .Y(new_n17789));
  nor_5  g15441(.A(new_n17789), .B(new_n12233), .Y(new_n17790));
  or_6   g15442(.A(new_n17790), .B(new_n17788), .Y(new_n17791));
  not_8  g15443(.A(new_n17791), .Y(new_n17792));
  nand_5 g15444(.A(new_n17792), .B(new_n17766), .Y(new_n17793));
  nand_5 g15445(.A(new_n17793), .B(new_n17765), .Y(new_n17794));
  or_6   g15446(.A(new_n17794), .B(new_n17763), .Y(new_n17795));
  nand_5 g15447(.A(new_n17795), .B(new_n12232), .Y(new_n17796));
  nand_5 g15448(.A(new_n17794), .B(new_n17763), .Y(new_n17797));
  nand_5 g15449(.A(new_n17797), .B(new_n17796), .Y(new_n17798));
  xor_4  g15450(.A(new_n5318), .B(pi123), .Y(new_n17799));
  nand_5 g15451(.A(new_n5383), .B(new_n10229), .Y(new_n17800));
  not_8  g15452(.A(new_n17800), .Y(new_n17801));
  not_8  g15453(.A(new_n12205), .Y(new_n17802));
  nor_5  g15454(.A(new_n12230), .B(new_n17802), .Y(new_n17803));
  nor_5  g15455(.A(new_n17803), .B(new_n17801), .Y(new_n17804));
  xor_4  g15456(.A(new_n17804), .B(new_n17799), .Y(new_n17805));
  xor_4  g15457(.A(new_n17805), .B(new_n17798), .Y(new_n17806));
  not_8  g15458(.A(new_n17806), .Y(new_n17807));
  xor_4  g15459(.A(new_n17807), .B(new_n17761), .Y(po0223));
  xor_4  g15460(.A(pi715), .B(new_n3527), .Y(new_n17809));
  nor_5  g15461(.A(pi428), .B(new_n16199), .Y(new_n17810));
  xor_4  g15462(.A(pi428), .B(new_n16199), .Y(new_n17811));
  not_8  g15463(.A(new_n17811), .Y(new_n17812));
  nand_5 g15464(.A(pi196), .B(new_n16167), .Y(new_n17813));
  xor_4  g15465(.A(pi196), .B(new_n16167), .Y(new_n17814));
  nand_5 g15466(.A(new_n5198), .B(new_n5195), .Y(new_n17815));
  nand_5 g15467(.A(new_n17815), .B(new_n5197), .Y(new_n17816));
  nand_5 g15468(.A(new_n17816), .B(new_n17814), .Y(new_n17817));
  nand_5 g15469(.A(new_n17817), .B(new_n17813), .Y(new_n17818));
  nor_5  g15470(.A(new_n17818), .B(new_n17812), .Y(new_n17819));
  nor_5  g15471(.A(new_n17819), .B(new_n17810), .Y(new_n17820));
  xor_4  g15472(.A(new_n17820), .B(new_n17809), .Y(new_n17821));
  not_8  g15473(.A(new_n17821), .Y(new_n17822));
  nor_5  g15474(.A(new_n17822), .B(new_n13340), .Y(new_n17823));
  xor_4  g15475(.A(new_n17821), .B(new_n13340), .Y(new_n17824));
  xor_4  g15476(.A(new_n17818), .B(new_n17811), .Y(new_n17825));
  and_6  g15477(.A(new_n17825), .B(new_n13343), .Y(new_n17826));
  not_8  g15478(.A(new_n13356), .Y(new_n17827));
  xnor_4 g15479(.A(new_n17816), .B(new_n17814), .Y(new_n17828));
  nor_5  g15480(.A(new_n17828), .B(new_n17827), .Y(new_n17829));
  xor_4  g15481(.A(new_n17828), .B(new_n13356), .Y(new_n17830));
  nand_5 g15482(.A(new_n5200), .B(new_n5191), .Y(new_n17831));
  nand_5 g15483(.A(new_n5201), .B(new_n5176), .Y(new_n17832));
  and_6  g15484(.A(new_n17832), .B(new_n17831), .Y(new_n17833));
  nor_5  g15485(.A(new_n17833), .B(new_n17830), .Y(new_n17834));
  nor_5  g15486(.A(new_n17834), .B(new_n17829), .Y(new_n17835));
  xnor_4 g15487(.A(new_n17825), .B(new_n13343), .Y(new_n17836));
  nor_5  g15488(.A(new_n17836), .B(new_n17835), .Y(new_n17837));
  nor_5  g15489(.A(new_n17837), .B(new_n17826), .Y(new_n17838));
  nor_5  g15490(.A(new_n17838), .B(new_n17824), .Y(new_n17839));
  or_6   g15491(.A(new_n17839), .B(new_n17823), .Y(new_n17840));
  xor_4  g15492(.A(pi785), .B(new_n16216), .Y(new_n17841));
  nor_5  g15493(.A(new_n16220), .B(pi331), .Y(new_n17842));
  not_8  g15494(.A(new_n17809), .Y(new_n17843));
  nor_5  g15495(.A(new_n17820), .B(new_n17843), .Y(new_n17844));
  nor_5  g15496(.A(new_n17844), .B(new_n17842), .Y(new_n17845));
  xnor_4 g15497(.A(new_n17845), .B(new_n17841), .Y(new_n17846));
  xor_4  g15498(.A(new_n17846), .B(new_n13336), .Y(new_n17847));
  xnor_4 g15499(.A(new_n17847), .B(new_n17840), .Y(po0224));
  nand_5 g15500(.A(new_n11768), .B(new_n6392), .Y(new_n17849));
  nor_5  g15501(.A(new_n11768), .B(new_n6392), .Y(new_n17850));
  not_8  g15502(.A(new_n17850), .Y(new_n17851));
  nand_5 g15503(.A(new_n17851), .B(new_n17849), .Y(new_n17852));
  not_8  g15504(.A(new_n17852), .Y(new_n17853));
  nand_5 g15505(.A(new_n6255), .B(new_n14080), .Y(new_n17854));
  xor_4  g15506(.A(new_n6255), .B(new_n14080), .Y(new_n17855));
  nand_5 g15507(.A(new_n4065), .B(new_n4060), .Y(new_n17856));
  nand_5 g15508(.A(new_n4071), .B(new_n4066), .Y(new_n17857));
  nand_5 g15509(.A(new_n17857), .B(new_n17856), .Y(new_n17858));
  nand_5 g15510(.A(new_n17858), .B(new_n17855), .Y(new_n17859));
  nand_5 g15511(.A(new_n17859), .B(new_n17854), .Y(new_n17860));
  nand_5 g15512(.A(new_n17860), .B(new_n14078), .Y(new_n17861));
  xor_4  g15513(.A(new_n17860), .B(new_n14078), .Y(new_n17862));
  not_8  g15514(.A(new_n17862), .Y(new_n17863));
  or_6   g15515(.A(new_n17863), .B(new_n6279), .Y(new_n17864));
  nand_5 g15516(.A(new_n17864), .B(new_n17861), .Y(new_n17865));
  nand_5 g15517(.A(new_n17865), .B(new_n14174), .Y(new_n17866));
  not_8  g15518(.A(new_n17866), .Y(new_n17867));
  xor_4  g15519(.A(new_n17865), .B(pi419), .Y(new_n17868));
  nor_5  g15520(.A(new_n17868), .B(new_n6327), .Y(new_n17869));
  nor_5  g15521(.A(new_n17869), .B(new_n17867), .Y(new_n17870));
  not_8  g15522(.A(new_n17870), .Y(new_n17871));
  nand_5 g15523(.A(new_n6361), .B(pi056), .Y(new_n17872));
  nand_5 g15524(.A(new_n6360), .B(new_n6372), .Y(new_n17873));
  nand_5 g15525(.A(new_n17873), .B(new_n17872), .Y(new_n17874));
  xor_4  g15526(.A(new_n17874), .B(new_n17871), .Y(new_n17875));
  nor_5  g15527(.A(new_n17875), .B(new_n11848), .Y(new_n17876));
  xor_4  g15528(.A(new_n17868), .B(new_n6326), .Y(new_n17877));
  or_6   g15529(.A(new_n17877), .B(new_n11784), .Y(new_n17878));
  xor_4  g15530(.A(new_n17863), .B(new_n6279), .Y(new_n17879));
  nand_5 g15531(.A(new_n17879), .B(new_n11793), .Y(new_n17880));
  xor_4  g15532(.A(new_n17858), .B(new_n17855), .Y(new_n17881));
  not_8  g15533(.A(new_n17881), .Y(new_n17882));
  nor_5  g15534(.A(new_n17882), .B(new_n11796), .Y(new_n17883));
  nor_5  g15535(.A(new_n4072), .B(new_n4058), .Y(new_n17884));
  or_6   g15536(.A(new_n4073), .B(new_n4041), .Y(new_n17885));
  not_8  g15537(.A(new_n17885), .Y(new_n17886));
  nor_5  g15538(.A(new_n17886), .B(new_n17884), .Y(new_n17887));
  xor_4  g15539(.A(new_n17881), .B(new_n11796), .Y(new_n17888));
  nor_5  g15540(.A(new_n17888), .B(new_n17887), .Y(new_n17889));
  nor_5  g15541(.A(new_n17889), .B(new_n17883), .Y(new_n17890));
  not_8  g15542(.A(new_n17890), .Y(new_n17891));
  xor_4  g15543(.A(new_n17879), .B(new_n11793), .Y(new_n17892));
  nand_5 g15544(.A(new_n17892), .B(new_n17891), .Y(new_n17893));
  nand_5 g15545(.A(new_n17893), .B(new_n17880), .Y(new_n17894));
  xor_4  g15546(.A(new_n17877), .B(new_n11784), .Y(new_n17895));
  nand_5 g15547(.A(new_n17895), .B(new_n17894), .Y(new_n17896));
  nand_5 g15548(.A(new_n17896), .B(new_n17878), .Y(new_n17897));
  xor_4  g15549(.A(new_n17875), .B(new_n11848), .Y(new_n17898));
  nand_5 g15550(.A(new_n17898), .B(new_n17897), .Y(new_n17899));
  not_8  g15551(.A(new_n17899), .Y(new_n17900));
  nor_5  g15552(.A(new_n17900), .B(new_n17876), .Y(new_n17901));
  nand_5 g15553(.A(new_n17872), .B(new_n17871), .Y(new_n17902));
  nand_5 g15554(.A(new_n17902), .B(new_n17873), .Y(new_n17903));
  xor_4  g15555(.A(new_n17903), .B(new_n17901), .Y(new_n17904));
  xor_4  g15556(.A(new_n17904), .B(new_n17853), .Y(po0225));
  nor_5  g15557(.A(new_n12640), .B(new_n12639), .Y(new_n17906));
  xor_4  g15558(.A(new_n17906), .B(new_n12641), .Y(po0226));
  xnor_4 g15559(.A(new_n6065), .B(new_n6064), .Y(po0227));
  xor_4  g15560(.A(new_n13102), .B(new_n6051), .Y(po0228));
  xnor_4 g15561(.A(new_n14444), .B(new_n14398), .Y(po0229));
  or_6   g15562(.A(pi466), .B(new_n4930), .Y(new_n17911));
  xor_4  g15563(.A(pi466), .B(new_n4930), .Y(new_n17912));
  nand_5 g15564(.A(new_n4721), .B(pi086), .Y(new_n17913));
  nand_5 g15565(.A(new_n17472), .B(new_n17468), .Y(new_n17914));
  nand_5 g15566(.A(new_n17914), .B(new_n17913), .Y(new_n17915));
  nand_5 g15567(.A(new_n17915), .B(new_n17912), .Y(new_n17916));
  nand_5 g15568(.A(new_n17916), .B(new_n17911), .Y(new_n17917));
  not_8  g15569(.A(new_n17917), .Y(new_n17918));
  nand_5 g15570(.A(new_n4873), .B(pi118), .Y(new_n17919));
  not_8  g15571(.A(pi118), .Y(new_n17920));
  nand_5 g15572(.A(pi124), .B(new_n17920), .Y(new_n17921));
  nand_5 g15573(.A(new_n17921), .B(new_n17919), .Y(new_n17922));
  xnor_4 g15574(.A(new_n17915), .B(new_n17912), .Y(new_n17923));
  or_6   g15575(.A(new_n17923), .B(new_n7792), .Y(new_n17924));
  xor_4  g15576(.A(new_n17923), .B(new_n7792), .Y(new_n17925));
  not_8  g15577(.A(new_n17473), .Y(new_n17926));
  nor_5  g15578(.A(new_n17926), .B(new_n7798), .Y(new_n17927));
  nor_5  g15579(.A(new_n17474), .B(new_n17467), .Y(new_n17928));
  or_6   g15580(.A(new_n17928), .B(new_n17927), .Y(new_n17929));
  nand_5 g15581(.A(new_n17929), .B(new_n17925), .Y(new_n17930));
  nand_5 g15582(.A(new_n17930), .B(new_n17924), .Y(new_n17931));
  nand_5 g15583(.A(new_n17931), .B(new_n7870), .Y(new_n17932));
  nor_5  g15584(.A(new_n17931), .B(new_n7870), .Y(new_n17933));
  not_8  g15585(.A(new_n17933), .Y(new_n17934));
  nand_5 g15586(.A(new_n17934), .B(new_n17932), .Y(new_n17935));
  xor_4  g15587(.A(new_n17935), .B(new_n17922), .Y(new_n17936));
  xor_4  g15588(.A(new_n17936), .B(new_n17918), .Y(new_n17937));
  xor_4  g15589(.A(new_n17929), .B(new_n17925), .Y(new_n17938));
  or_6   g15590(.A(new_n17938), .B(new_n7909), .Y(new_n17939));
  nand_5 g15591(.A(new_n17938), .B(new_n7909), .Y(new_n17940));
  nand_5 g15592(.A(new_n17305), .B(new_n13477), .Y(new_n17941));
  or_6   g15593(.A(new_n17306), .B(new_n7918), .Y(new_n17942));
  nand_5 g15594(.A(new_n17942), .B(new_n17941), .Y(new_n17943));
  or_6   g15595(.A(new_n17943), .B(new_n13430), .Y(new_n17944));
  xor_4  g15596(.A(new_n17943), .B(new_n13430), .Y(new_n17945));
  nand_5 g15597(.A(new_n17945), .B(new_n7916), .Y(new_n17946));
  nand_5 g15598(.A(new_n17946), .B(new_n17944), .Y(new_n17947));
  or_6   g15599(.A(new_n17947), .B(new_n17461), .Y(new_n17948));
  nand_5 g15600(.A(new_n17947), .B(new_n17461), .Y(new_n17949));
  nand_5 g15601(.A(new_n17949), .B(new_n7914), .Y(new_n17950));
  nand_5 g15602(.A(new_n17950), .B(new_n17948), .Y(new_n17951));
  nor_5  g15603(.A(new_n17951), .B(new_n17475), .Y(new_n17952));
  xor_4  g15604(.A(new_n17951), .B(new_n17475), .Y(new_n17953));
  not_8  g15605(.A(new_n17953), .Y(new_n17954));
  nor_5  g15606(.A(new_n17954), .B(new_n7913), .Y(new_n17955));
  or_6   g15607(.A(new_n17955), .B(new_n17952), .Y(new_n17956));
  nand_5 g15608(.A(new_n17956), .B(new_n17940), .Y(new_n17957));
  nand_5 g15609(.A(new_n17957), .B(new_n17939), .Y(new_n17958));
  and_6  g15610(.A(new_n17958), .B(new_n17937), .Y(new_n17959));
  not_8  g15611(.A(new_n13819), .Y(new_n17960));
  nor_5  g15612(.A(new_n17958), .B(new_n17937), .Y(new_n17961));
  and_6  g15613(.A(new_n17961), .B(new_n13820), .Y(new_n17962));
  nor_5  g15614(.A(new_n17962), .B(new_n17960), .Y(new_n17963));
  nor_5  g15615(.A(new_n17963), .B(new_n17959), .Y(new_n17964));
  not_8  g15616(.A(new_n17964), .Y(new_n17965));
  nand_5 g15617(.A(new_n17965), .B(new_n13820), .Y(new_n17966));
  nor_5  g15618(.A(new_n17959), .B(new_n7991), .Y(new_n17967));
  nand_5 g15619(.A(new_n17961), .B(new_n13821), .Y(new_n17968));
  not_8  g15620(.A(new_n17921), .Y(new_n17969));
  nand_5 g15621(.A(new_n17932), .B(new_n17918), .Y(new_n17970));
  nand_5 g15622(.A(new_n17970), .B(new_n17969), .Y(new_n17971));
  nand_5 g15623(.A(new_n17919), .B(new_n17917), .Y(new_n17972));
  or_6   g15624(.A(new_n17972), .B(new_n17932), .Y(new_n17973));
  nand_5 g15625(.A(new_n17973), .B(new_n17971), .Y(new_n17974));
  nand_5 g15626(.A(new_n17974), .B(new_n17934), .Y(new_n17975));
  nand_5 g15627(.A(new_n17972), .B(new_n17921), .Y(new_n17976));
  nor_5  g15628(.A(new_n17976), .B(new_n17934), .Y(new_n17977));
  nor_5  g15629(.A(new_n17970), .B(new_n17919), .Y(new_n17978));
  nor_5  g15630(.A(new_n17978), .B(new_n17977), .Y(new_n17979));
  nand_5 g15631(.A(new_n17979), .B(new_n17975), .Y(new_n17980));
  xor_4  g15632(.A(new_n17980), .B(new_n11868), .Y(new_n17981));
  nand_5 g15633(.A(new_n17981), .B(new_n17968), .Y(new_n17982));
  nor_5  g15634(.A(new_n17982), .B(new_n17967), .Y(new_n17983));
  nand_5 g15635(.A(new_n17983), .B(new_n17966), .Y(new_n17984));
  or_6   g15636(.A(new_n17961), .B(new_n17959), .Y(new_n17985));
  nor_5  g15637(.A(new_n17985), .B(new_n7993), .Y(new_n17986));
  nand_5 g15638(.A(new_n17959), .B(new_n13821), .Y(new_n17987));
  nor_5  g15639(.A(new_n17981), .B(new_n17962), .Y(new_n17988));
  nand_5 g15640(.A(new_n17988), .B(new_n17987), .Y(new_n17989));
  or_6   g15641(.A(new_n17989), .B(new_n17986), .Y(new_n17990));
  and_6  g15642(.A(new_n17990), .B(new_n17984), .Y(po0230));
  xor_4  g15643(.A(new_n14466), .B(new_n14454), .Y(po0231));
  xor_4  g15644(.A(pi228), .B(new_n10729), .Y(new_n17993));
  nand_5 g15645(.A(pi514), .B(new_n5021), .Y(new_n17994));
  xor_4  g15646(.A(pi514), .B(new_n5021), .Y(new_n17995));
  nand_5 g15647(.A(new_n5031), .B(pi369), .Y(new_n17996));
  nand_5 g15648(.A(pi438), .B(new_n5058), .Y(new_n17997));
  not_8  g15649(.A(new_n17997), .Y(new_n17998));
  xor_4  g15650(.A(pi617), .B(new_n2360), .Y(new_n17999));
  nand_5 g15651(.A(new_n17999), .B(new_n17998), .Y(new_n18000));
  nand_5 g15652(.A(new_n18000), .B(new_n17996), .Y(new_n18001));
  nand_5 g15653(.A(new_n18001), .B(new_n17995), .Y(new_n18002));
  nand_5 g15654(.A(new_n18002), .B(new_n17994), .Y(new_n18003));
  xnor_4 g15655(.A(new_n18003), .B(new_n17993), .Y(new_n18004));
  xor_4  g15656(.A(new_n18004), .B(new_n3066), .Y(new_n18005));
  xor_4  g15657(.A(new_n18001), .B(new_n17995), .Y(new_n18006));
  or_6   g15658(.A(new_n18006), .B(new_n3071), .Y(new_n18007));
  nand_5 g15659(.A(new_n18006), .B(new_n3071), .Y(new_n18008));
  and_6  g15660(.A(new_n3087), .B(new_n3076), .Y(new_n18009));
  or_6   g15661(.A(new_n18009), .B(new_n18000), .Y(new_n18010));
  nand_5 g15662(.A(new_n2420), .B(pi396), .Y(new_n18011));
  or_6   g15663(.A(new_n18011), .B(new_n3076), .Y(new_n18012));
  nand_5 g15664(.A(new_n17998), .B(new_n3076), .Y(new_n18013));
  nand_5 g15665(.A(new_n18013), .B(new_n18012), .Y(new_n18014));
  xor_4  g15666(.A(new_n18014), .B(new_n17999), .Y(new_n18015));
  nor_5  g15667(.A(new_n18015), .B(new_n3087), .Y(new_n18016));
  nor_5  g15668(.A(new_n18012), .B(new_n17999), .Y(new_n18017));
  nor_5  g15669(.A(new_n18017), .B(new_n18016), .Y(new_n18018));
  nand_5 g15670(.A(new_n18018), .B(new_n18010), .Y(new_n18019));
  nand_5 g15671(.A(new_n18019), .B(new_n18008), .Y(new_n18020));
  nand_5 g15672(.A(new_n18020), .B(new_n18007), .Y(new_n18021));
  xnor_4 g15673(.A(new_n18021), .B(new_n18005), .Y(po0232));
  xor_4  g15674(.A(new_n10812), .B(new_n5582), .Y(po0233));
  nand_5 g15675(.A(new_n6089), .B(new_n6091), .Y(new_n18024));
  or_6   g15676(.A(new_n6096), .B(new_n11994), .Y(new_n18025));
  not_8  g15677(.A(new_n18025), .Y(new_n18026));
  nand_5 g15678(.A(new_n18026), .B(new_n18024), .Y(new_n18027));
  nand_5 g15679(.A(new_n6090), .B(pi280), .Y(new_n18028));
  not_8  g15680(.A(new_n18028), .Y(new_n18029));
  nand_5 g15681(.A(new_n6098), .B(pi661), .Y(new_n18030));
  nand_5 g15682(.A(new_n18030), .B(new_n6096), .Y(new_n18031));
  nand_5 g15683(.A(new_n18031), .B(new_n18029), .Y(new_n18032));
  nand_5 g15684(.A(new_n18032), .B(new_n18027), .Y(new_n18033));
  not_8  g15685(.A(new_n18033), .Y(new_n18034));
  nand_5 g15686(.A(new_n6097), .B(new_n11994), .Y(new_n18035));
  not_8  g15687(.A(new_n18035), .Y(new_n18036));
  nand_5 g15688(.A(new_n18036), .B(new_n18028), .Y(new_n18037));
  not_8  g15689(.A(new_n18037), .Y(new_n18038));
  nor_5  g15690(.A(new_n18031), .B(new_n18024), .Y(new_n18039));
  nor_5  g15691(.A(new_n18039), .B(new_n18038), .Y(new_n18040));
  nand_5 g15692(.A(new_n18040), .B(new_n18034), .Y(new_n18041));
  not_8  g15693(.A(new_n18041), .Y(new_n18042));
  nand_5 g15694(.A(new_n18042), .B(new_n15558), .Y(new_n18043));
  not_8  g15695(.A(new_n18043), .Y(new_n18044));
  xor_4  g15696(.A(new_n18042), .B(new_n15558), .Y(new_n18045));
  not_8  g15697(.A(new_n18045), .Y(new_n18046));
  nand_5 g15698(.A(new_n13122), .B(new_n6101), .Y(new_n18047));
  or_6   g15699(.A(new_n13123), .B(new_n13077), .Y(new_n18048));
  nand_5 g15700(.A(new_n18048), .B(new_n18047), .Y(new_n18049));
  nor_5  g15701(.A(new_n18049), .B(new_n18046), .Y(new_n18050));
  nor_5  g15702(.A(new_n18050), .B(new_n18044), .Y(new_n18051));
  xor_4  g15703(.A(new_n18033), .B(new_n15550), .Y(new_n18052));
  xor_4  g15704(.A(new_n18052), .B(new_n18051), .Y(po0234));
  xor_4  g15705(.A(new_n9807), .B(new_n6139), .Y(po0235));
  xor_4  g15706(.A(new_n5698), .B(new_n5697), .Y(po0236));
  xnor_4 g15707(.A(new_n13906), .B(new_n13884), .Y(po0237));
  nand_5 g15708(.A(new_n16625), .B(pi477), .Y(new_n18057));
  nor_5  g15709(.A(new_n16626), .B(new_n16622), .Y(new_n18058));
  nand_5 g15710(.A(new_n18058), .B(new_n18057), .Y(new_n18059));
  nand_5 g15711(.A(new_n18059), .B(new_n16623), .Y(po0238));
  xor_4  g15712(.A(pi468), .B(new_n6836), .Y(new_n18061));
  nand_5 g15713(.A(pi783), .B(new_n6651), .Y(new_n18062));
  xor_4  g15714(.A(pi783), .B(new_n6651), .Y(new_n18063));
  nand_5 g15715(.A(new_n18063), .B(pi508), .Y(new_n18064));
  nand_5 g15716(.A(new_n18064), .B(new_n18062), .Y(new_n18065));
  xnor_4 g15717(.A(new_n18065), .B(new_n18061), .Y(new_n18066));
  xor_4  g15718(.A(pi223), .B(new_n2487), .Y(new_n18067));
  nor_5  g15719(.A(new_n9104), .B(new_n9083), .Y(new_n18068));
  xor_4  g15720(.A(new_n18068), .B(new_n18067), .Y(new_n18069));
  not_8  g15721(.A(new_n18069), .Y(new_n18070));
  nand_5 g15722(.A(new_n18070), .B(pi393), .Y(new_n18071));
  nand_5 g15723(.A(new_n18071), .B(new_n18064), .Y(new_n18072));
  nand_5 g15724(.A(new_n18069), .B(new_n5693), .Y(new_n18073));
  and_6  g15725(.A(new_n18073), .B(new_n18071), .Y(new_n18074));
  or_6   g15726(.A(new_n18074), .B(pi508), .Y(new_n18075));
  xor_4  g15727(.A(new_n18073), .B(new_n18063), .Y(new_n18076));
  xor_4  g15728(.A(new_n18076), .B(new_n18075), .Y(new_n18077));
  nand_5 g15729(.A(new_n18077), .B(new_n18072), .Y(new_n18078));
  xor_4  g15730(.A(pi839), .B(pi611), .Y(new_n18079));
  xor_4  g15731(.A(new_n18079), .B(new_n5037), .Y(new_n18080));
  nand_5 g15732(.A(new_n2428), .B(new_n5596), .Y(new_n18081));
  nand_5 g15733(.A(new_n18081), .B(new_n5033), .Y(new_n18082));
  nand_5 g15734(.A(pi223), .B(pi214), .Y(new_n18083));
  nand_5 g15735(.A(new_n18083), .B(new_n18082), .Y(new_n18084));
  xor_4  g15736(.A(new_n18084), .B(new_n18080), .Y(new_n18085));
  or_6   g15737(.A(new_n18085), .B(new_n18077), .Y(new_n18086));
  nand_5 g15738(.A(new_n18086), .B(new_n18078), .Y(new_n18087));
  nand_5 g15739(.A(new_n18087), .B(new_n18066), .Y(new_n18088));
  nand_5 g15740(.A(new_n9434), .B(new_n2388), .Y(new_n18089));
  nand_5 g15741(.A(pi836), .B(pi486), .Y(new_n18090));
  nand_5 g15742(.A(new_n18090), .B(new_n18089), .Y(new_n18091));
  nor_5  g15743(.A(new_n18085), .B(new_n5036), .Y(new_n18092));
  xor_4  g15744(.A(new_n18092), .B(new_n18091), .Y(new_n18093));
  nor_5  g15745(.A(pi839), .B(pi611), .Y(new_n18094));
  or_6   g15746(.A(new_n18084), .B(new_n18094), .Y(new_n18095));
  nand_5 g15747(.A(pi839), .B(pi611), .Y(new_n18096));
  nand_5 g15748(.A(new_n18084), .B(new_n18096), .Y(new_n18097));
  nand_5 g15749(.A(new_n18097), .B(new_n18095), .Y(new_n18098));
  xor_4  g15750(.A(new_n18098), .B(new_n18093), .Y(new_n18099));
  xor_4  g15751(.A(new_n18099), .B(new_n5030), .Y(new_n18100));
  xor_4  g15752(.A(new_n18087), .B(new_n18066), .Y(new_n18101));
  nand_5 g15753(.A(new_n18101), .B(new_n18100), .Y(new_n18102));
  nand_5 g15754(.A(new_n18102), .B(new_n18088), .Y(new_n18103));
  xor_4  g15755(.A(pi252), .B(new_n3230), .Y(new_n18104));
  nand_5 g15756(.A(pi468), .B(new_n6836), .Y(new_n18105));
  nand_5 g15757(.A(new_n18065), .B(new_n18061), .Y(new_n18106));
  nand_5 g15758(.A(new_n18106), .B(new_n18105), .Y(new_n18107));
  xnor_4 g15759(.A(new_n18107), .B(new_n18104), .Y(new_n18108));
  or_6   g15760(.A(new_n18108), .B(new_n18103), .Y(new_n18109));
  xor_4  g15761(.A(new_n18108), .B(new_n18103), .Y(new_n18110));
  not_8  g15762(.A(new_n5030), .Y(new_n18111));
  or_6   g15763(.A(new_n18099), .B(new_n18111), .Y(new_n18112));
  nor_5  g15764(.A(new_n18079), .B(new_n5036), .Y(new_n18113));
  nor_5  g15765(.A(new_n18084), .B(new_n18080), .Y(new_n18114));
  or_6   g15766(.A(new_n18114), .B(new_n18113), .Y(new_n18115));
  nand_5 g15767(.A(new_n18115), .B(new_n18099), .Y(new_n18116));
  nand_5 g15768(.A(new_n18116), .B(new_n18112), .Y(new_n18117));
  xor_4  g15769(.A(pi289), .B(pi200), .Y(new_n18118));
  nand_5 g15770(.A(new_n18090), .B(new_n18096), .Y(new_n18119));
  nand_5 g15771(.A(new_n18119), .B(new_n18089), .Y(new_n18120));
  xor_4  g15772(.A(new_n18120), .B(new_n18118), .Y(new_n18121));
  xor_4  g15773(.A(new_n18121), .B(new_n15462), .Y(new_n18122));
  xor_4  g15774(.A(new_n18122), .B(new_n18117), .Y(new_n18123));
  nand_5 g15775(.A(new_n18123), .B(new_n18110), .Y(new_n18124));
  nand_5 g15776(.A(new_n18124), .B(new_n18109), .Y(new_n18125));
  nand_5 g15777(.A(new_n5654), .B(pi074), .Y(new_n18126));
  nand_5 g15778(.A(new_n18107), .B(new_n18104), .Y(new_n18127));
  nand_5 g15779(.A(new_n18127), .B(new_n18126), .Y(new_n18128));
  xor_4  g15780(.A(pi584), .B(new_n5651), .Y(new_n18129));
  xor_4  g15781(.A(new_n18129), .B(new_n18128), .Y(new_n18130));
  or_6   g15782(.A(new_n18130), .B(new_n18125), .Y(new_n18131));
  nand_5 g15783(.A(new_n18130), .B(new_n18125), .Y(new_n18132));
  nand_5 g15784(.A(new_n2385), .B(new_n5515), .Y(new_n18133));
  nand_5 g15785(.A(new_n18120), .B(new_n18118), .Y(new_n18134));
  nand_5 g15786(.A(new_n18134), .B(new_n18133), .Y(new_n18135));
  nand_5 g15787(.A(new_n9526), .B(new_n2405), .Y(new_n18136));
  nand_5 g15788(.A(pi492), .B(pi055), .Y(new_n18137));
  nand_5 g15789(.A(new_n18137), .B(new_n18136), .Y(new_n18138));
  xor_4  g15790(.A(new_n18138), .B(new_n18135), .Y(new_n18139));
  xor_4  g15791(.A(new_n18139), .B(new_n15476), .Y(new_n18140));
  not_8  g15792(.A(new_n18140), .Y(new_n18141));
  nor_5  g15793(.A(new_n18121), .B(new_n15462), .Y(new_n18142));
  not_8  g15794(.A(new_n18122), .Y(new_n18143));
  nor_5  g15795(.A(new_n18143), .B(new_n18117), .Y(new_n18144));
  nor_5  g15796(.A(new_n18144), .B(new_n18142), .Y(new_n18145));
  xor_4  g15797(.A(new_n18145), .B(new_n18141), .Y(new_n18146));
  not_8  g15798(.A(new_n18146), .Y(new_n18147));
  nand_5 g15799(.A(new_n18147), .B(new_n18132), .Y(new_n18148));
  nand_5 g15800(.A(new_n18148), .B(new_n18131), .Y(new_n18149));
  nand_5 g15801(.A(pi584), .B(new_n5651), .Y(new_n18150));
  nand_5 g15802(.A(new_n18129), .B(new_n18128), .Y(new_n18151));
  nand_5 g15803(.A(new_n18151), .B(new_n18150), .Y(new_n18152));
  nand_5 g15804(.A(new_n5648), .B(pi225), .Y(new_n18153));
  nand_5 g15805(.A(pi539), .B(new_n3222), .Y(new_n18154));
  nand_5 g15806(.A(new_n18154), .B(new_n18153), .Y(new_n18155));
  xor_4  g15807(.A(new_n18155), .B(new_n18152), .Y(new_n18156));
  xor_4  g15808(.A(new_n18156), .B(new_n18149), .Y(new_n18157));
  xor_4  g15809(.A(pi699), .B(pi373), .Y(new_n18158));
  nand_5 g15810(.A(new_n18137), .B(new_n18135), .Y(new_n18159));
  nand_5 g15811(.A(new_n18159), .B(new_n18136), .Y(new_n18160));
  xor_4  g15812(.A(new_n18160), .B(new_n18158), .Y(new_n18161));
  xor_4  g15813(.A(new_n18161), .B(new_n16075), .Y(new_n18162));
  or_6   g15814(.A(new_n18139), .B(new_n16077), .Y(new_n18163));
  nand_5 g15815(.A(new_n18145), .B(new_n18141), .Y(new_n18164));
  nand_5 g15816(.A(new_n18164), .B(new_n18163), .Y(new_n18165));
  xor_4  g15817(.A(new_n18165), .B(new_n18162), .Y(new_n18166));
  xor_4  g15818(.A(new_n18166), .B(new_n18157), .Y(po0239));
  xor_4  g15819(.A(new_n14180), .B(new_n14178), .Y(po0240));
  xnor_4 g15820(.A(new_n15781), .B(new_n15779), .Y(po0241));
  not_8  g15821(.A(new_n17710), .Y(new_n18170));
  nand_5 g15822(.A(new_n9253), .B(pi542), .Y(new_n18171));
  nand_5 g15823(.A(new_n9254), .B(new_n15546), .Y(new_n18172));
  nand_5 g15824(.A(new_n18172), .B(new_n18171), .Y(new_n18173));
  nor_5  g15825(.A(new_n18173), .B(new_n18170), .Y(new_n18174));
  xor_4  g15826(.A(new_n18173), .B(new_n17710), .Y(new_n18175));
  nor_5  g15827(.A(new_n18175), .B(new_n8048), .Y(new_n18176));
  nor_5  g15828(.A(new_n18176), .B(new_n18174), .Y(new_n18177));
  not_8  g15829(.A(new_n10961), .Y(new_n18178));
  nor_5  g15830(.A(new_n10974), .B(new_n17689), .Y(new_n18179));
  nand_5 g15831(.A(new_n18179), .B(new_n18178), .Y(new_n18180));
  nor_5  g15832(.A(new_n18179), .B(new_n18178), .Y(new_n18181));
  nand_5 g15833(.A(new_n10974), .B(new_n17689), .Y(new_n18182));
  nand_5 g15834(.A(new_n18182), .B(new_n10962), .Y(new_n18183));
  nor_5  g15835(.A(new_n18183), .B(new_n18181), .Y(new_n18184));
  nand_5 g15836(.A(new_n18184), .B(new_n10958), .Y(new_n18185));
  nand_5 g15837(.A(new_n18185), .B(new_n18180), .Y(new_n18186));
  not_8  g15838(.A(new_n18186), .Y(new_n18187));
  nor_5  g15839(.A(new_n18187), .B(new_n18177), .Y(new_n18188));
  nor_5  g15840(.A(new_n18182), .B(new_n10962), .Y(new_n18189));
  nand_5 g15841(.A(new_n18183), .B(new_n18181), .Y(new_n18190));
  nor_5  g15842(.A(new_n18190), .B(new_n10958), .Y(new_n18191));
  or_6   g15843(.A(new_n18191), .B(new_n18189), .Y(new_n18192));
  nand_5 g15844(.A(new_n18174), .B(new_n8047), .Y(new_n18193));
  nor_5  g15845(.A(new_n18193), .B(new_n18192), .Y(new_n18194));
  nor_5  g15846(.A(new_n18194), .B(new_n18188), .Y(po0242));
  xnor_4 g15847(.A(new_n16404), .B(new_n16402), .Y(po0243));
  xor_4  g15848(.A(new_n17270), .B(new_n17225), .Y(po0244));
  xnor_4 g15849(.A(new_n17430), .B(new_n17417), .Y(po0245));
  xnor_4 g15850(.A(new_n16414), .B(new_n16413), .Y(po0246));
  xor_4  g15851(.A(new_n9449), .B(new_n9456), .Y(po0247));
  xor_4  g15852(.A(pi704), .B(new_n8086), .Y(new_n18201));
  nand_5 g15853(.A(new_n8062), .B(pi065), .Y(new_n18202));
  xor_4  g15854(.A(new_n8062), .B(pi065), .Y(new_n18203));
  nand_5 g15855(.A(new_n8075), .B(pi195), .Y(new_n18204));
  xor_4  g15856(.A(new_n8075), .B(pi195), .Y(new_n18205));
  nand_5 g15857(.A(new_n8063), .B(pi379), .Y(new_n18206));
  not_8  g15858(.A(new_n9983), .Y(new_n18207));
  xor_4  g15859(.A(pi474), .B(new_n9978), .Y(new_n18208));
  nand_5 g15860(.A(new_n18208), .B(new_n18207), .Y(new_n18209));
  nand_5 g15861(.A(new_n18209), .B(new_n18206), .Y(new_n18210));
  nand_5 g15862(.A(new_n18210), .B(new_n18205), .Y(new_n18211));
  nand_5 g15863(.A(new_n18211), .B(new_n18204), .Y(new_n18212));
  nand_5 g15864(.A(new_n18212), .B(new_n18203), .Y(new_n18213));
  nand_5 g15865(.A(new_n18213), .B(new_n18202), .Y(new_n18214));
  xor_4  g15866(.A(new_n18214), .B(new_n18201), .Y(new_n18215));
  xor_4  g15867(.A(new_n18215), .B(new_n15381), .Y(new_n18216));
  xnor_4 g15868(.A(new_n18212), .B(new_n18203), .Y(new_n18217));
  nor_5  g15869(.A(new_n18217), .B(new_n15688), .Y(new_n18218));
  xor_4  g15870(.A(new_n18217), .B(new_n15688), .Y(new_n18219));
  not_8  g15871(.A(new_n18219), .Y(new_n18220));
  xnor_4 g15872(.A(new_n18210), .B(new_n18205), .Y(new_n18221));
  or_6   g15873(.A(new_n18221), .B(new_n15389), .Y(new_n18222));
  nand_5 g15874(.A(new_n18208), .B(new_n15391), .Y(new_n18223));
  or_6   g15875(.A(new_n9984), .B(new_n2753), .Y(new_n18224));
  nand_5 g15876(.A(new_n18207), .B(new_n2753), .Y(new_n18225));
  nand_5 g15877(.A(new_n18225), .B(new_n18224), .Y(new_n18226));
  xor_4  g15878(.A(new_n18208), .B(new_n15392), .Y(new_n18227));
  not_8  g15879(.A(new_n18227), .Y(new_n18228));
  or_6   g15880(.A(new_n18228), .B(new_n18226), .Y(new_n18229));
  nand_5 g15881(.A(new_n18229), .B(new_n18224), .Y(new_n18230));
  nand_5 g15882(.A(new_n18230), .B(new_n18223), .Y(new_n18231));
  and_6  g15883(.A(new_n15337), .B(new_n2753), .Y(new_n18232));
  or_6   g15884(.A(new_n18232), .B(new_n18209), .Y(new_n18233));
  nand_5 g15885(.A(new_n18233), .B(new_n18231), .Y(new_n18234));
  nand_5 g15886(.A(new_n18234), .B(new_n18222), .Y(new_n18235));
  nand_5 g15887(.A(new_n18221), .B(new_n15389), .Y(new_n18236));
  nand_5 g15888(.A(new_n18236), .B(new_n18235), .Y(new_n18237));
  nor_5  g15889(.A(new_n18237), .B(new_n18220), .Y(new_n18238));
  nor_5  g15890(.A(new_n18238), .B(new_n18218), .Y(new_n18239));
  xor_4  g15891(.A(new_n18239), .B(new_n18216), .Y(new_n18240));
  xor_4  g15892(.A(new_n18227), .B(new_n18226), .Y(new_n18241));
  not_8  g15893(.A(new_n18241), .Y(new_n18242));
  not_8  g15894(.A(new_n15226), .Y(new_n18243));
  nor_5  g15895(.A(new_n18243), .B(new_n9933), .Y(new_n18244));
  nor_5  g15896(.A(new_n15226), .B(new_n9931), .Y(new_n18245));
  or_6   g15897(.A(new_n18245), .B(new_n18244), .Y(new_n18246));
  xor_4  g15898(.A(new_n18246), .B(new_n9927), .Y(new_n18247));
  or_6   g15899(.A(new_n18247), .B(new_n18242), .Y(new_n18248));
  or_6   g15900(.A(new_n18246), .B(new_n9927), .Y(new_n18249));
  not_8  g15901(.A(new_n13733), .Y(new_n18250));
  nor_5  g15902(.A(new_n18244), .B(new_n18250), .Y(new_n18251));
  nand_5 g15903(.A(new_n18251), .B(new_n18249), .Y(new_n18252));
  nand_5 g15904(.A(new_n18252), .B(new_n18248), .Y(new_n18253));
  nand_5 g15905(.A(new_n18253), .B(new_n13752), .Y(new_n18254));
  not_8  g15906(.A(new_n18254), .Y(new_n18255));
  xor_4  g15907(.A(new_n18253), .B(new_n13751), .Y(new_n18256));
  nand_5 g15908(.A(new_n18236), .B(new_n18222), .Y(new_n18257));
  xor_4  g15909(.A(new_n18257), .B(new_n18234), .Y(new_n18258));
  not_8  g15910(.A(new_n18258), .Y(new_n18259));
  nor_5  g15911(.A(new_n18259), .B(new_n18256), .Y(new_n18260));
  nor_5  g15912(.A(new_n18260), .B(new_n18255), .Y(new_n18261));
  xor_4  g15913(.A(new_n18237), .B(new_n18219), .Y(new_n18262));
  nand_5 g15914(.A(new_n18262), .B(new_n18261), .Y(new_n18263));
  not_8  g15915(.A(new_n18262), .Y(new_n18264));
  xor_4  g15916(.A(new_n18264), .B(new_n18261), .Y(new_n18265));
  not_8  g15917(.A(new_n18265), .Y(new_n18266));
  nand_5 g15918(.A(new_n18266), .B(new_n13737), .Y(new_n18267));
  nand_5 g15919(.A(new_n18267), .B(new_n18263), .Y(new_n18268));
  nand_5 g15920(.A(new_n18268), .B(new_n18240), .Y(new_n18269));
  xor_4  g15921(.A(new_n18268), .B(new_n18240), .Y(new_n18270));
  nand_5 g15922(.A(new_n18270), .B(new_n15360), .Y(new_n18271));
  nand_5 g15923(.A(new_n18271), .B(new_n18269), .Y(new_n18272));
  nand_5 g15924(.A(pi704), .B(new_n8086), .Y(new_n18273));
  nand_5 g15925(.A(new_n18214), .B(new_n18201), .Y(new_n18274));
  nand_5 g15926(.A(new_n18274), .B(new_n18273), .Y(new_n18275));
  nand_5 g15927(.A(new_n8091), .B(pi222), .Y(new_n18276));
  or_6   g15928(.A(new_n8091), .B(pi222), .Y(new_n18277));
  nand_5 g15929(.A(new_n18277), .B(new_n18276), .Y(new_n18278));
  xor_4  g15930(.A(new_n18278), .B(new_n18275), .Y(new_n18279));
  xor_4  g15931(.A(new_n18279), .B(new_n15687), .Y(new_n18280));
  or_6   g15932(.A(new_n18215), .B(new_n15381), .Y(new_n18281));
  nand_5 g15933(.A(new_n18239), .B(new_n18216), .Y(new_n18282));
  nand_5 g15934(.A(new_n18282), .B(new_n18281), .Y(new_n18283));
  xor_4  g15935(.A(new_n18283), .B(new_n18280), .Y(new_n18284));
  not_8  g15936(.A(new_n18284), .Y(new_n18285));
  xor_4  g15937(.A(new_n18285), .B(new_n18272), .Y(new_n18286));
  xnor_4 g15938(.A(new_n18286), .B(new_n15356), .Y(po0248));
  nand_5 g15939(.A(new_n17716), .B(new_n17715), .Y(new_n18288));
  xor_4  g15940(.A(new_n18288), .B(new_n17727), .Y(po0249));
  xor_4  g15941(.A(new_n7553), .B(new_n10554), .Y(new_n18290));
  nand_5 g15942(.A(new_n17089), .B(pi377), .Y(new_n18291));
  nand_5 g15943(.A(new_n18291), .B(new_n17088), .Y(new_n18292));
  nor_5  g15944(.A(new_n18292), .B(new_n7557), .Y(new_n18293));
  nor_5  g15945(.A(new_n18293), .B(new_n10470), .Y(new_n18294));
  nand_5 g15946(.A(new_n18292), .B(new_n7557), .Y(new_n18295));
  not_8  g15947(.A(new_n18295), .Y(new_n18296));
  nor_5  g15948(.A(new_n18296), .B(new_n18294), .Y(new_n18297));
  not_8  g15949(.A(new_n18297), .Y(new_n18298));
  or_6   g15950(.A(new_n18298), .B(new_n18290), .Y(new_n18299));
  nor_5  g15951(.A(new_n7553), .B(pi735), .Y(new_n18300));
  nor_5  g15952(.A(new_n18300), .B(new_n7528), .Y(new_n18301));
  nand_5 g15953(.A(new_n18301), .B(new_n18299), .Y(new_n18302));
  nand_5 g15954(.A(new_n7528), .B(new_n10554), .Y(new_n18303));
  nor_5  g15955(.A(new_n18303), .B(new_n18298), .Y(new_n18304));
  nand_5 g15956(.A(new_n18298), .B(pi735), .Y(new_n18305));
  not_8  g15957(.A(new_n7526), .Y(new_n18306));
  nor_5  g15958(.A(new_n18306), .B(new_n7514), .Y(new_n18307));
  nand_5 g15959(.A(new_n18307), .B(new_n18305), .Y(new_n18308));
  not_8  g15960(.A(new_n18308), .Y(new_n18309));
  nor_5  g15961(.A(new_n18309), .B(new_n18304), .Y(new_n18310));
  nand_5 g15962(.A(new_n18310), .B(new_n18302), .Y(new_n18311));
  nand_5 g15963(.A(pi728), .B(new_n3212), .Y(new_n18312));
  xor_4  g15964(.A(pi728), .B(new_n3212), .Y(new_n18313));
  nand_5 g15965(.A(new_n5205), .B(pi073), .Y(new_n18314));
  nand_5 g15966(.A(new_n17100), .B(new_n17097), .Y(new_n18315));
  nand_5 g15967(.A(new_n18315), .B(new_n18314), .Y(new_n18316));
  nand_5 g15968(.A(new_n18316), .B(new_n18313), .Y(new_n18317));
  nand_5 g15969(.A(new_n18317), .B(new_n18312), .Y(new_n18318));
  nand_5 g15970(.A(new_n18318), .B(pi096), .Y(new_n18319));
  nand_5 g15971(.A(pi800), .B(pi244), .Y(new_n18320));
  xor_4  g15972(.A(new_n18316), .B(new_n18313), .Y(new_n18321));
  nor_5  g15973(.A(new_n18321), .B(new_n12073), .Y(new_n18322));
  or_6   g15974(.A(new_n17102), .B(new_n17096), .Y(new_n18323));
  not_8  g15975(.A(new_n18323), .Y(new_n18324));
  nor_5  g15976(.A(new_n17101), .B(new_n6824), .Y(new_n18325));
  nor_5  g15977(.A(new_n18325), .B(new_n18324), .Y(new_n18326));
  xor_4  g15978(.A(new_n18321), .B(pi666), .Y(new_n18327));
  nor_5  g15979(.A(new_n18327), .B(new_n18326), .Y(new_n18328));
  nor_5  g15980(.A(new_n18328), .B(new_n18322), .Y(new_n18329));
  not_8  g15981(.A(new_n18329), .Y(new_n18330));
  nand_5 g15982(.A(new_n8986), .B(new_n3209), .Y(new_n18331));
  nand_5 g15983(.A(new_n18331), .B(new_n18330), .Y(new_n18332));
  nand_5 g15984(.A(new_n18332), .B(new_n18320), .Y(new_n18333));
  or_6   g15985(.A(new_n18333), .B(new_n18319), .Y(new_n18334));
  nor_5  g15986(.A(new_n18318), .B(pi096), .Y(new_n18335));
  nor_5  g15987(.A(new_n18335), .B(new_n18331), .Y(new_n18336));
  nand_5 g15988(.A(new_n18336), .B(new_n18329), .Y(new_n18337));
  nand_5 g15989(.A(new_n18337), .B(new_n18334), .Y(new_n18338));
  not_8  g15990(.A(new_n18319), .Y(new_n18339));
  nor_5  g15991(.A(new_n18320), .B(new_n18339), .Y(new_n18340));
  nand_5 g15992(.A(new_n18340), .B(new_n18330), .Y(new_n18341));
  nand_5 g15993(.A(new_n18335), .B(new_n18333), .Y(new_n18342));
  nand_5 g15994(.A(new_n18342), .B(new_n18341), .Y(new_n18343));
  nor_5  g15995(.A(new_n18343), .B(new_n18338), .Y(new_n18344));
  xor_4  g15996(.A(new_n18344), .B(new_n18311), .Y(new_n18345));
  xor_4  g15997(.A(new_n18297), .B(new_n18290), .Y(new_n18346));
  nor_5  g15998(.A(new_n18335), .B(new_n18339), .Y(new_n18347));
  and_6  g15999(.A(new_n18331), .B(new_n18320), .Y(new_n18348));
  xor_4  g16000(.A(new_n18348), .B(new_n18347), .Y(new_n18349));
  not_8  g16001(.A(new_n18349), .Y(new_n18350));
  xor_4  g16002(.A(new_n18350), .B(new_n18329), .Y(new_n18351));
  nor_5  g16003(.A(new_n18351), .B(new_n18346), .Y(new_n18352));
  nor_5  g16004(.A(new_n18296), .B(new_n18293), .Y(new_n18353));
  xor_4  g16005(.A(new_n18353), .B(pi533), .Y(new_n18354));
  xor_4  g16006(.A(new_n18327), .B(new_n18326), .Y(new_n18355));
  or_6   g16007(.A(new_n18355), .B(new_n18354), .Y(new_n18356));
  nand_5 g16008(.A(new_n18355), .B(new_n18354), .Y(new_n18357));
  nand_5 g16009(.A(new_n17091), .B(new_n17085), .Y(new_n18358));
  or_6   g16010(.A(new_n17103), .B(new_n17092), .Y(new_n18359));
  nand_5 g16011(.A(new_n18359), .B(new_n18358), .Y(new_n18360));
  nand_5 g16012(.A(new_n18360), .B(new_n18357), .Y(new_n18361));
  nand_5 g16013(.A(new_n18361), .B(new_n18356), .Y(new_n18362));
  xor_4  g16014(.A(new_n18351), .B(new_n18346), .Y(new_n18363));
  nand_5 g16015(.A(new_n18363), .B(new_n18362), .Y(new_n18364));
  not_8  g16016(.A(new_n18364), .Y(new_n18365));
  nor_5  g16017(.A(new_n18365), .B(new_n18352), .Y(new_n18366));
  nand_5 g16018(.A(new_n18366), .B(new_n18345), .Y(new_n18367));
  nor_5  g16019(.A(new_n18335), .B(pi244), .Y(new_n18368));
  nor_5  g16020(.A(new_n18368), .B(new_n18339), .Y(new_n18369));
  nor_5  g16021(.A(new_n18369), .B(new_n18338), .Y(new_n18370));
  xor_4  g16022(.A(new_n18370), .B(new_n18302), .Y(new_n18371));
  nor_5  g16023(.A(new_n18371), .B(new_n18367), .Y(new_n18372));
  not_8  g16024(.A(new_n18367), .Y(new_n18373));
  or_6   g16025(.A(new_n18344), .B(new_n18311), .Y(new_n18374));
  nand_5 g16026(.A(new_n18371), .B(new_n18374), .Y(new_n18375));
  nor_5  g16027(.A(new_n18375), .B(new_n18373), .Y(new_n18376));
  or_6   g16028(.A(new_n18376), .B(new_n18372), .Y(po0250));
  nand_5 g16029(.A(new_n9169), .B(new_n16941), .Y(new_n18378));
  not_8  g16030(.A(new_n18378), .Y(new_n18379));
  xor_4  g16031(.A(pi512), .B(pi068), .Y(new_n18380));
  not_8  g16032(.A(new_n18380), .Y(new_n18381));
  nand_5 g16033(.A(new_n11899), .B(new_n9154), .Y(new_n18382));
  not_8  g16034(.A(new_n18382), .Y(new_n18383));
  not_8  g16035(.A(new_n2896), .Y(new_n18384));
  nor_5  g16036(.A(new_n2937), .B(new_n18384), .Y(new_n18385));
  nor_5  g16037(.A(new_n18385), .B(new_n18383), .Y(new_n18386));
  nor_5  g16038(.A(new_n18386), .B(new_n18381), .Y(new_n18387));
  nor_5  g16039(.A(new_n18387), .B(new_n18379), .Y(new_n18388));
  not_8  g16040(.A(new_n15266), .Y(new_n18389));
  xor_4  g16041(.A(new_n18386), .B(new_n18380), .Y(new_n18390));
  nand_5 g16042(.A(new_n18390), .B(new_n18389), .Y(new_n18391));
  not_8  g16043(.A(new_n18390), .Y(new_n18392));
  xor_4  g16044(.A(new_n18392), .B(new_n15266), .Y(new_n18393));
  nand_5 g16045(.A(new_n2980), .B(new_n2938), .Y(new_n18394));
  nand_5 g16046(.A(new_n3044), .B(new_n2981), .Y(new_n18395));
  nand_5 g16047(.A(new_n18395), .B(new_n18394), .Y(new_n18396));
  nand_5 g16048(.A(new_n18396), .B(new_n18393), .Y(new_n18397));
  nand_5 g16049(.A(new_n18397), .B(new_n18391), .Y(new_n18398));
  nand_5 g16050(.A(new_n18398), .B(new_n18388), .Y(new_n18399));
  nand_5 g16051(.A(new_n18399), .B(new_n15264), .Y(new_n18400));
  nor_5  g16052(.A(new_n18398), .B(new_n18388), .Y(new_n18401));
  not_8  g16053(.A(new_n18401), .Y(new_n18402));
  nand_5 g16054(.A(new_n18402), .B(new_n18400), .Y(new_n18403));
  nor_5  g16055(.A(new_n18399), .B(new_n15264), .Y(new_n18404));
  not_8  g16056(.A(new_n18404), .Y(new_n18405));
  nand_5 g16057(.A(new_n18401), .B(new_n15264), .Y(new_n18406));
  nand_5 g16058(.A(new_n18406), .B(new_n18405), .Y(new_n18407));
  not_8  g16059(.A(new_n18407), .Y(new_n18408));
  nand_5 g16060(.A(new_n18408), .B(new_n18403), .Y(new_n18409));
  nand_5 g16061(.A(pi358), .B(new_n10405), .Y(new_n18410));
  xor_4  g16062(.A(pi358), .B(new_n10405), .Y(new_n18411));
  nand_5 g16063(.A(pi687), .B(new_n2837), .Y(new_n18412));
  nand_5 g16064(.A(new_n2894), .B(new_n2853), .Y(new_n18413));
  nand_5 g16065(.A(new_n18413), .B(new_n18412), .Y(new_n18414));
  nand_5 g16066(.A(new_n18414), .B(new_n18411), .Y(new_n18415));
  nand_5 g16067(.A(new_n18415), .B(new_n18410), .Y(new_n18416));
  nand_5 g16068(.A(new_n18409), .B(new_n18405), .Y(new_n18417));
  xor_4  g16069(.A(new_n18417), .B(new_n18416), .Y(new_n18418));
  not_8  g16070(.A(new_n18418), .Y(new_n18419));
  nor_5  g16071(.A(new_n18419), .B(new_n18400), .Y(new_n18420));
  and_6  g16072(.A(new_n18416), .B(new_n18405), .Y(new_n18421));
  nor_5  g16073(.A(new_n18416), .B(new_n18401), .Y(new_n18422));
  or_6   g16074(.A(new_n18422), .B(new_n18421), .Y(new_n18423));
  xor_4  g16075(.A(new_n18414), .B(new_n18411), .Y(new_n18424));
  xor_4  g16076(.A(new_n18396), .B(new_n18393), .Y(new_n18425));
  nand_5 g16077(.A(new_n18425), .B(new_n18424), .Y(new_n18426));
  xor_4  g16078(.A(new_n18425), .B(new_n18424), .Y(new_n18427));
  nand_5 g16079(.A(new_n3045), .B(new_n2895), .Y(new_n18428));
  nand_5 g16080(.A(new_n3104), .B(new_n3046), .Y(new_n18429));
  nand_5 g16081(.A(new_n18429), .B(new_n18428), .Y(new_n18430));
  nand_5 g16082(.A(new_n18430), .B(new_n18427), .Y(new_n18431));
  nand_5 g16083(.A(new_n18431), .B(new_n18426), .Y(new_n18432));
  not_8  g16084(.A(new_n18432), .Y(new_n18433));
  nand_5 g16085(.A(new_n18433), .B(new_n18419), .Y(new_n18434));
  nand_5 g16086(.A(new_n18434), .B(new_n18423), .Y(new_n18435));
  nor_5  g16087(.A(new_n18435), .B(new_n18420), .Y(new_n18436));
  nor_5  g16088(.A(new_n18434), .B(new_n18423), .Y(new_n18437));
  nor_5  g16089(.A(new_n18437), .B(new_n18436), .Y(po0411));
  or_6   g16090(.A(po0411), .B(new_n18409), .Y(new_n18439));
  not_8  g16091(.A(new_n18434), .Y(new_n18440));
  nand_5 g16092(.A(new_n18440), .B(new_n18422), .Y(new_n18441));
  nand_5 g16093(.A(new_n18441), .B(new_n18439), .Y(po0251));
  nand_5 g16094(.A(new_n3026), .B(pi369), .Y(new_n18443));
  nor_5  g16095(.A(new_n18443), .B(new_n2358), .Y(new_n18444));
  xor_4  g16096(.A(new_n18443), .B(pi514), .Y(new_n18445));
  nor_5  g16097(.A(new_n18445), .B(new_n3011), .Y(new_n18446));
  or_6   g16098(.A(new_n18446), .B(new_n18444), .Y(new_n18447));
  xor_4  g16099(.A(new_n18447), .B(new_n3006), .Y(new_n18448));
  xor_4  g16100(.A(new_n18448), .B(new_n10729), .Y(new_n18449));
  nor_5  g16101(.A(new_n18449), .B(new_n6889), .Y(new_n18450));
  xor_4  g16102(.A(new_n18449), .B(new_n6917), .Y(new_n18451));
  xor_4  g16103(.A(new_n18445), .B(new_n3011), .Y(new_n18452));
  xor_4  g16104(.A(new_n3025), .B(pi369), .Y(new_n18453));
  nand_5 g16105(.A(new_n3022), .B(pi438), .Y(new_n18454));
  nand_5 g16106(.A(new_n3021), .B(new_n2420), .Y(new_n18455));
  nand_5 g16107(.A(new_n18455), .B(new_n6902), .Y(new_n18456));
  nand_5 g16108(.A(new_n18456), .B(new_n18454), .Y(new_n18457));
  not_8  g16109(.A(new_n18457), .Y(new_n18458));
  nor_5  g16110(.A(new_n18458), .B(new_n18453), .Y(new_n18459));
  xor_4  g16111(.A(new_n18457), .B(new_n18453), .Y(new_n18460));
  nor_5  g16112(.A(new_n18460), .B(new_n6899), .Y(new_n18461));
  or_6   g16113(.A(new_n18461), .B(new_n18459), .Y(new_n18462));
  and_6  g16114(.A(new_n18462), .B(new_n18452), .Y(new_n18463));
  xnor_4 g16115(.A(new_n18462), .B(new_n18452), .Y(new_n18464));
  nor_5  g16116(.A(new_n18464), .B(new_n6897), .Y(new_n18465));
  nor_5  g16117(.A(new_n18465), .B(new_n18463), .Y(new_n18466));
  nor_5  g16118(.A(new_n18466), .B(new_n18451), .Y(new_n18467));
  or_6   g16119(.A(new_n18467), .B(new_n18450), .Y(new_n18468));
  nand_5 g16120(.A(new_n18447), .B(new_n3006), .Y(new_n18469));
  nand_5 g16121(.A(new_n18448), .B(pi117), .Y(new_n18470));
  nand_5 g16122(.A(new_n18470), .B(new_n18469), .Y(new_n18471));
  nand_5 g16123(.A(new_n18471), .B(new_n3000), .Y(new_n18472));
  or_6   g16124(.A(new_n18471), .B(new_n3000), .Y(new_n18473));
  and_6  g16125(.A(new_n18473), .B(new_n18472), .Y(new_n18474));
  xor_4  g16126(.A(new_n18474), .B(new_n7758), .Y(new_n18475));
  xor_4  g16127(.A(new_n18475), .B(new_n18468), .Y(new_n18476));
  xor_4  g16128(.A(new_n18476), .B(new_n6882), .Y(po0252));
  xnor_4 g16129(.A(new_n3672), .B(new_n3671), .Y(po0253));
  xor_4  g16130(.A(new_n5810), .B(new_n3861), .Y(po0254));
  xor_4  g16131(.A(new_n12714), .B(new_n12682), .Y(po0255));
  nand_5 g16132(.A(pi612), .B(new_n7019), .Y(new_n18481));
  nand_5 g16133(.A(new_n3552), .B(pi337), .Y(new_n18482));
  and_6  g16134(.A(new_n18482), .B(new_n18481), .Y(new_n18483));
  xor_4  g16135(.A(pi617), .B(pi270), .Y(new_n18484));
  xor_4  g16136(.A(new_n18484), .B(new_n2363), .Y(new_n18485));
  nand_5 g16137(.A(pi396), .B(pi367), .Y(new_n18486));
  nand_5 g16138(.A(new_n5058), .B(new_n6975), .Y(new_n18487));
  nand_5 g16139(.A(new_n18487), .B(new_n2365), .Y(new_n18488));
  nand_5 g16140(.A(new_n18488), .B(new_n18486), .Y(new_n18489));
  nor_5  g16141(.A(new_n18489), .B(new_n2427), .Y(new_n18490));
  nor_5  g16142(.A(new_n18486), .B(new_n2421), .Y(new_n18491));
  nor_5  g16143(.A(new_n18491), .B(new_n18490), .Y(new_n18492));
  xor_4  g16144(.A(new_n18492), .B(new_n18485), .Y(new_n18493));
  nand_5 g16145(.A(new_n7138), .B(new_n6976), .Y(new_n18494));
  nand_5 g16146(.A(new_n18011), .B(new_n17997), .Y(new_n18495));
  xor_4  g16147(.A(new_n18495), .B(new_n18494), .Y(new_n18496));
  nand_5 g16148(.A(new_n18496), .B(new_n7059), .Y(new_n18497));
  not_8  g16149(.A(new_n18496), .Y(new_n18498));
  nand_5 g16150(.A(new_n18498), .B(new_n7056), .Y(new_n18499));
  nand_5 g16151(.A(new_n18499), .B(new_n18497), .Y(new_n18500));
  xor_4  g16152(.A(new_n18500), .B(new_n18493), .Y(new_n18501));
  xor_4  g16153(.A(new_n18501), .B(new_n18483), .Y(po0256));
  xnor_4 g16154(.A(new_n13891), .B(new_n2561), .Y(po0257));
  xor_4  g16155(.A(new_n15046), .B(new_n15044), .Y(po0258));
  xor_4  g16156(.A(new_n16411), .B(new_n16396), .Y(po0259));
  nand_5 g16157(.A(new_n14527), .B(pi174), .Y(new_n18506));
  xor_4  g16158(.A(new_n14503), .B(new_n5196), .Y(new_n18507));
  or_6   g16159(.A(new_n15484), .B(new_n14505), .Y(new_n18508));
  nand_5 g16160(.A(new_n15485), .B(pi653), .Y(new_n18509));
  nand_5 g16161(.A(new_n18509), .B(new_n18508), .Y(new_n18510));
  nand_5 g16162(.A(new_n18510), .B(new_n18507), .Y(new_n18511));
  nand_5 g16163(.A(new_n18511), .B(new_n18506), .Y(new_n18512));
  nand_5 g16164(.A(new_n18512), .B(new_n14500), .Y(new_n18513));
  xor_4  g16165(.A(new_n18512), .B(new_n14499), .Y(new_n18514));
  or_6   g16166(.A(new_n18514), .B(new_n16167), .Y(new_n18515));
  nand_5 g16167(.A(new_n18515), .B(new_n18513), .Y(new_n18516));
  nand_5 g16168(.A(new_n18516), .B(new_n17516), .Y(new_n18517));
  xor_4  g16169(.A(new_n18516), .B(new_n14497), .Y(new_n18518));
  or_6   g16170(.A(new_n18518), .B(new_n16199), .Y(new_n18519));
  nand_5 g16171(.A(new_n18519), .B(new_n18517), .Y(new_n18520));
  nand_5 g16172(.A(new_n18520), .B(pi715), .Y(new_n18521));
  xor_4  g16173(.A(new_n18520), .B(new_n16220), .Y(new_n18522));
  or_6   g16174(.A(new_n18522), .B(new_n14626), .Y(new_n18523));
  nand_5 g16175(.A(new_n18523), .B(new_n18521), .Y(new_n18524));
  xor_4  g16176(.A(new_n18524), .B(new_n17530), .Y(new_n18525));
  xor_4  g16177(.A(new_n18525), .B(new_n16216), .Y(new_n18526));
  xor_4  g16178(.A(new_n18518), .B(new_n16199), .Y(new_n18527));
  xor_4  g16179(.A(new_n18510), .B(new_n18507), .Y(new_n18528));
  not_8  g16180(.A(new_n18528), .Y(new_n18529));
  nand_5 g16181(.A(new_n15488), .B(new_n15471), .Y(new_n18530));
  nand_5 g16182(.A(new_n18530), .B(new_n15487), .Y(new_n18531));
  nand_5 g16183(.A(new_n18531), .B(new_n18529), .Y(new_n18532));
  xor_4  g16184(.A(new_n18531), .B(new_n18528), .Y(new_n18533));
  or_6   g16185(.A(new_n18533), .B(new_n16100), .Y(new_n18534));
  nand_5 g16186(.A(new_n18534), .B(new_n18532), .Y(new_n18535));
  or_6   g16187(.A(new_n18535), .B(new_n16159), .Y(new_n18536));
  xor_4  g16188(.A(new_n18535), .B(new_n16159), .Y(new_n18537));
  xor_4  g16189(.A(new_n18514), .B(new_n16167), .Y(new_n18538));
  nand_5 g16190(.A(new_n18538), .B(new_n18537), .Y(new_n18539));
  nand_5 g16191(.A(new_n18539), .B(new_n18536), .Y(new_n18540));
  nand_5 g16192(.A(new_n18540), .B(new_n18527), .Y(new_n18541));
  not_8  g16193(.A(new_n16179), .Y(new_n18542));
  xor_4  g16194(.A(new_n18540), .B(new_n18527), .Y(new_n18543));
  nand_5 g16195(.A(new_n18543), .B(new_n18542), .Y(new_n18544));
  nand_5 g16196(.A(new_n18544), .B(new_n18541), .Y(new_n18545));
  xor_4  g16197(.A(new_n18522), .B(new_n14626), .Y(new_n18546));
  or_6   g16198(.A(new_n18546), .B(new_n18545), .Y(new_n18547));
  nand_5 g16199(.A(new_n18546), .B(new_n18545), .Y(new_n18548));
  nand_5 g16200(.A(new_n18548), .B(new_n16098), .Y(new_n18549));
  nand_5 g16201(.A(new_n18549), .B(new_n18547), .Y(new_n18550));
  xnor_4 g16202(.A(new_n18550), .B(new_n16096), .Y(new_n18551));
  xnor_4 g16203(.A(new_n18551), .B(new_n18526), .Y(po0260));
  not_8  g16204(.A(new_n4325), .Y(new_n18553));
  nor_5  g16205(.A(new_n4524), .B(new_n18553), .Y(new_n18554));
  nor_5  g16206(.A(new_n4530), .B(new_n4325), .Y(new_n18555));
  or_6   g16207(.A(new_n18555), .B(new_n18554), .Y(po0261));
  nand_5 g16208(.A(new_n11389), .B(new_n11387), .Y(new_n18557));
  nand_5 g16209(.A(new_n18557), .B(new_n11388), .Y(new_n18558));
  not_8  g16210(.A(new_n18558), .Y(new_n18559));
  xor_4  g16211(.A(new_n18559), .B(new_n7242), .Y(new_n18560));
  or_6   g16212(.A(new_n11392), .B(new_n7211), .Y(new_n18561));
  not_8  g16213(.A(new_n7113), .Y(new_n18562));
  nor_5  g16214(.A(new_n11410), .B(new_n18562), .Y(new_n18563));
  nor_5  g16215(.A(new_n12716), .B(new_n12679), .Y(new_n18564));
  or_6   g16216(.A(new_n18564), .B(new_n18563), .Y(new_n18565));
  xor_4  g16217(.A(new_n11392), .B(new_n7211), .Y(new_n18566));
  nand_5 g16218(.A(new_n18566), .B(new_n18565), .Y(new_n18567));
  nand_5 g16219(.A(new_n18567), .B(new_n18561), .Y(new_n18568));
  not_8  g16220(.A(new_n18568), .Y(new_n18569));
  xor_4  g16221(.A(new_n18569), .B(new_n18560), .Y(po0262));
  xor_4  g16222(.A(new_n6631), .B(new_n6628), .Y(po0263));
  xnor_4 g16223(.A(new_n17272), .B(new_n17220), .Y(po0264));
  xor_4  g16224(.A(pi253), .B(new_n6714), .Y(new_n18573));
  nand_5 g16225(.A(new_n3264), .B(pi615), .Y(new_n18574));
  nand_5 g16226(.A(new_n16914), .B(new_n16898), .Y(new_n18575));
  nand_5 g16227(.A(new_n18575), .B(new_n18574), .Y(new_n18576));
  xnor_4 g16228(.A(new_n18576), .B(new_n18573), .Y(new_n18577));
  nor_5  g16229(.A(new_n18577), .B(new_n7396), .Y(new_n18578));
  xor_4  g16230(.A(new_n18577), .B(new_n7397), .Y(new_n18579));
  or_6   g16231(.A(new_n16915), .B(new_n16897), .Y(new_n18580));
  nand_5 g16232(.A(new_n16939), .B(new_n16916), .Y(new_n18581));
  nand_5 g16233(.A(new_n18581), .B(new_n18580), .Y(new_n18582));
  nor_5  g16234(.A(new_n18582), .B(new_n18579), .Y(new_n18583));
  or_6   g16235(.A(new_n18583), .B(new_n18578), .Y(new_n18584));
  nand_5 g16236(.A(new_n3333), .B(pi022), .Y(new_n18585));
  nand_5 g16237(.A(new_n18576), .B(new_n18573), .Y(new_n18586));
  nand_5 g16238(.A(new_n18586), .B(new_n18585), .Y(new_n18587));
  nand_5 g16239(.A(new_n3303), .B(pi073), .Y(new_n18588));
  nand_5 g16240(.A(pi637), .B(new_n6787), .Y(new_n18589));
  nand_5 g16241(.A(new_n18589), .B(new_n18588), .Y(new_n18590));
  xor_4  g16242(.A(new_n18590), .B(new_n18587), .Y(new_n18591));
  xor_4  g16243(.A(new_n18591), .B(new_n7395), .Y(new_n18592));
  xnor_4 g16244(.A(new_n18592), .B(new_n18584), .Y(po0265));
  nand_5 g16245(.A(new_n7250), .B(pi622), .Y(new_n18594));
  or_6   g16246(.A(new_n18594), .B(new_n16611), .Y(new_n18595));
  xor_4  g16247(.A(new_n18594), .B(new_n16611), .Y(new_n18596));
  nand_5 g16248(.A(new_n18596), .B(new_n8833), .Y(new_n18597));
  nand_5 g16249(.A(new_n18597), .B(new_n18595), .Y(new_n18598));
  nand_5 g16250(.A(new_n18598), .B(new_n8825), .Y(new_n18599));
  or_6   g16251(.A(new_n18598), .B(new_n8825), .Y(new_n18600));
  nand_5 g16252(.A(new_n18600), .B(pi017), .Y(new_n18601));
  nand_5 g16253(.A(new_n18601), .B(new_n18599), .Y(new_n18602));
  nand_5 g16254(.A(new_n18602), .B(new_n8820), .Y(new_n18603));
  or_6   g16255(.A(new_n18602), .B(new_n8820), .Y(new_n18604));
  nand_5 g16256(.A(new_n18604), .B(pi129), .Y(new_n18605));
  nand_5 g16257(.A(new_n18605), .B(new_n18603), .Y(new_n18606));
  nand_5 g16258(.A(new_n18606), .B(new_n8815), .Y(new_n18607));
  or_6   g16259(.A(new_n18606), .B(new_n8815), .Y(new_n18608));
  nand_5 g16260(.A(new_n18608), .B(new_n18607), .Y(new_n18609));
  xor_4  g16261(.A(new_n18609), .B(pi210), .Y(new_n18610));
  and_6  g16262(.A(new_n18604), .B(new_n18603), .Y(new_n18611));
  xor_4  g16263(.A(new_n18611), .B(pi129), .Y(new_n18612));
  not_8  g16264(.A(new_n18612), .Y(new_n18613));
  nand_5 g16265(.A(new_n4104), .B(new_n4075), .Y(new_n18614));
  nor_5  g16266(.A(new_n4099), .B(pi708), .Y(new_n18615));
  nand_5 g16267(.A(new_n4096), .B(pi837), .Y(new_n18616));
  nand_5 g16268(.A(new_n18616), .B(new_n18615), .Y(new_n18617));
  nand_5 g16269(.A(new_n18617), .B(new_n18614), .Y(new_n18618));
  nand_5 g16270(.A(new_n18618), .B(new_n4095), .Y(new_n18619));
  or_6   g16271(.A(new_n18618), .B(new_n4095), .Y(new_n18620));
  nand_5 g16272(.A(new_n18620), .B(new_n6809), .Y(new_n18621));
  nand_5 g16273(.A(new_n18621), .B(new_n18619), .Y(new_n18622));
  xor_4  g16274(.A(new_n18622), .B(new_n16678), .Y(new_n18623));
  xor_4  g16275(.A(new_n18623), .B(new_n17743), .Y(new_n18624));
  nor_5  g16276(.A(new_n18624), .B(new_n18613), .Y(new_n18625));
  xor_4  g16277(.A(new_n18624), .B(new_n18612), .Y(new_n18626));
  nand_5 g16278(.A(new_n18600), .B(new_n18599), .Y(new_n18627));
  xor_4  g16279(.A(new_n18627), .B(pi017), .Y(new_n18628));
  nand_5 g16280(.A(new_n18619), .B(new_n18620), .Y(new_n18629));
  xor_4  g16281(.A(new_n18629), .B(pi760), .Y(new_n18630));
  not_8  g16282(.A(new_n18630), .Y(new_n18631));
  nor_5  g16283(.A(new_n18631), .B(new_n18628), .Y(new_n18632));
  xor_4  g16284(.A(new_n18596), .B(new_n8833), .Y(new_n18633));
  nand_5 g16285(.A(new_n18614), .B(new_n18616), .Y(new_n18634));
  not_8  g16286(.A(new_n18615), .Y(new_n18635));
  nand_5 g16287(.A(new_n8996), .B(new_n18635), .Y(new_n18636));
  nand_5 g16288(.A(new_n4099), .B(pi708), .Y(new_n18637));
  not_8  g16289(.A(new_n8996), .Y(new_n18638));
  nand_5 g16290(.A(new_n18638), .B(new_n18637), .Y(new_n18639));
  nand_5 g16291(.A(new_n18639), .B(new_n18636), .Y(new_n18640));
  xnor_4 g16292(.A(new_n18640), .B(new_n18634), .Y(new_n18641));
  and_6  g16293(.A(new_n18641), .B(new_n18633), .Y(new_n18642));
  and_6  g16294(.A(new_n18637), .B(new_n18635), .Y(new_n18643));
  nor_5  g16295(.A(new_n8996), .B(new_n18643), .Y(new_n18644));
  nor_5  g16296(.A(new_n18644), .B(new_n18641), .Y(new_n18645));
  nor_5  g16297(.A(new_n18645), .B(new_n18642), .Y(new_n18646));
  xor_4  g16298(.A(new_n18630), .B(new_n18628), .Y(new_n18647));
  nor_5  g16299(.A(new_n18647), .B(new_n18646), .Y(new_n18648));
  nor_5  g16300(.A(new_n18648), .B(new_n18632), .Y(new_n18649));
  nor_5  g16301(.A(new_n18649), .B(new_n18626), .Y(new_n18650));
  or_6   g16302(.A(new_n18650), .B(new_n18625), .Y(new_n18651));
  not_8  g16303(.A(new_n16678), .Y(new_n18652));
  nor_5  g16304(.A(new_n18622), .B(new_n18652), .Y(new_n18653));
  nor_5  g16305(.A(new_n18623), .B(new_n17743), .Y(new_n18654));
  or_6   g16306(.A(new_n18654), .B(new_n18653), .Y(new_n18655));
  nand_5 g16307(.A(new_n18655), .B(new_n16687), .Y(new_n18656));
  or_6   g16308(.A(new_n18655), .B(new_n16687), .Y(new_n18657));
  nand_5 g16309(.A(new_n18657), .B(new_n18656), .Y(new_n18658));
  xor_4  g16310(.A(new_n18658), .B(pi587), .Y(new_n18659));
  xnor_4 g16311(.A(new_n18659), .B(new_n18651), .Y(new_n18660));
  xnor_4 g16312(.A(new_n18660), .B(new_n18610), .Y(po0266));
  nor_5  g16313(.A(new_n18559), .B(new_n7239), .Y(new_n18662));
  xor_4  g16314(.A(new_n18559), .B(new_n7239), .Y(new_n18663));
  not_8  g16315(.A(new_n18663), .Y(new_n18664));
  not_8  g16316(.A(new_n7242), .Y(new_n18665));
  nand_5 g16317(.A(new_n18558), .B(new_n18665), .Y(new_n18666));
  nand_5 g16318(.A(new_n18569), .B(new_n18560), .Y(new_n18667));
  nand_5 g16319(.A(new_n18667), .B(new_n18666), .Y(new_n18668));
  nor_5  g16320(.A(new_n18668), .B(new_n18664), .Y(new_n18669));
  or_6   g16321(.A(new_n18669), .B(new_n18662), .Y(po0267));
  not_8  g16322(.A(new_n5544), .Y(new_n18671));
  nand_5 g16323(.A(new_n5497), .B(new_n9174), .Y(new_n18672));
  not_8  g16324(.A(new_n18672), .Y(new_n18673));
  nand_5 g16325(.A(pi811), .B(pi692), .Y(new_n18674));
  nand_5 g16326(.A(pi804), .B(pi625), .Y(new_n18675));
  nand_5 g16327(.A(new_n8770), .B(new_n5511), .Y(new_n18676));
  not_8  g16328(.A(new_n18676), .Y(new_n18677));
  nor_5  g16329(.A(pi739), .B(pi273), .Y(new_n18678));
  nor_5  g16330(.A(pi576), .B(pi067), .Y(new_n18679));
  nand_5 g16331(.A(pi675), .B(pi401), .Y(new_n18680));
  not_8  g16332(.A(new_n18680), .Y(new_n18681));
  xor_4  g16333(.A(pi576), .B(new_n5517), .Y(new_n18682));
  nor_5  g16334(.A(new_n18682), .B(new_n18681), .Y(new_n18683));
  nor_5  g16335(.A(new_n18683), .B(new_n18679), .Y(new_n18684));
  xor_4  g16336(.A(pi739), .B(new_n8773), .Y(new_n18685));
  nor_5  g16337(.A(new_n18685), .B(new_n18684), .Y(new_n18686));
  nor_5  g16338(.A(new_n18686), .B(new_n18678), .Y(new_n18687));
  xor_4  g16339(.A(pi573), .B(new_n5511), .Y(new_n18688));
  nor_5  g16340(.A(new_n18688), .B(new_n18687), .Y(new_n18689));
  nor_5  g16341(.A(new_n18689), .B(new_n18677), .Y(new_n18690));
  not_8  g16342(.A(new_n18690), .Y(new_n18691));
  xor_4  g16343(.A(pi804), .B(new_n5507), .Y(new_n18692));
  or_6   g16344(.A(new_n18692), .B(new_n18691), .Y(new_n18693));
  nand_5 g16345(.A(new_n18693), .B(new_n18675), .Y(new_n18694));
  xor_4  g16346(.A(pi811), .B(pi692), .Y(new_n18695));
  nand_5 g16347(.A(new_n18695), .B(new_n18694), .Y(new_n18696));
  nand_5 g16348(.A(new_n18696), .B(new_n18674), .Y(new_n18697));
  nand_5 g16349(.A(new_n5499), .B(new_n8759), .Y(new_n18698));
  nand_5 g16350(.A(pi737), .B(pi123), .Y(new_n18699));
  nand_5 g16351(.A(new_n18699), .B(new_n18698), .Y(new_n18700));
  xnor_4 g16352(.A(new_n18700), .B(new_n18697), .Y(new_n18701));
  nand_5 g16353(.A(new_n18701), .B(pi342), .Y(new_n18702));
  xor_4  g16354(.A(new_n18701), .B(pi342), .Y(new_n18703));
  xnor_4 g16355(.A(new_n18695), .B(new_n18694), .Y(new_n18704));
  or_6   g16356(.A(new_n18704), .B(new_n5505), .Y(new_n18705));
  xor_4  g16357(.A(new_n18692), .B(new_n18690), .Y(new_n18706));
  nor_5  g16358(.A(new_n18706), .B(new_n5509), .Y(new_n18707));
  xor_4  g16359(.A(new_n18706), .B(pi373), .Y(new_n18708));
  xor_4  g16360(.A(new_n18688), .B(new_n18687), .Y(new_n18709));
  nor_5  g16361(.A(new_n18709), .B(new_n9526), .Y(new_n18710));
  xor_4  g16362(.A(new_n18685), .B(new_n18684), .Y(new_n18711));
  nor_5  g16363(.A(new_n18711), .B(new_n5515), .Y(new_n18712));
  xor_4  g16364(.A(new_n18682), .B(new_n18680), .Y(new_n18713));
  nor_5  g16365(.A(new_n18713), .B(pi836), .Y(new_n18714));
  xor_4  g16366(.A(new_n18713), .B(pi836), .Y(new_n18715));
  not_8  g16367(.A(new_n18715), .Y(new_n18716));
  nand_5 g16368(.A(new_n16886), .B(pi839), .Y(new_n18717));
  or_6   g16369(.A(new_n16889), .B(new_n16887), .Y(new_n18718));
  nand_5 g16370(.A(new_n18718), .B(new_n18717), .Y(new_n18719));
  nor_5  g16371(.A(new_n18719), .B(new_n18716), .Y(new_n18720));
  or_6   g16372(.A(new_n18720), .B(new_n18714), .Y(new_n18721));
  xor_4  g16373(.A(new_n18711), .B(pi200), .Y(new_n18722));
  nor_5  g16374(.A(new_n18722), .B(new_n18721), .Y(new_n18723));
  nor_5  g16375(.A(new_n18723), .B(new_n18712), .Y(new_n18724));
  xor_4  g16376(.A(new_n18709), .B(pi492), .Y(new_n18725));
  nor_5  g16377(.A(new_n18725), .B(new_n18724), .Y(new_n18726));
  or_6   g16378(.A(new_n18726), .B(new_n18710), .Y(new_n18727));
  not_8  g16379(.A(new_n18727), .Y(new_n18728));
  nor_5  g16380(.A(new_n18728), .B(new_n18708), .Y(new_n18729));
  or_6   g16381(.A(new_n18729), .B(new_n18707), .Y(new_n18730));
  xor_4  g16382(.A(new_n18704), .B(pi549), .Y(new_n18731));
  not_8  g16383(.A(new_n18731), .Y(new_n18732));
  nand_5 g16384(.A(new_n18732), .B(new_n18730), .Y(new_n18733));
  nand_5 g16385(.A(new_n18733), .B(new_n18705), .Y(new_n18734));
  nand_5 g16386(.A(new_n18734), .B(new_n18703), .Y(new_n18735));
  nand_5 g16387(.A(new_n18735), .B(new_n18702), .Y(new_n18736));
  nand_5 g16388(.A(new_n18698), .B(new_n18697), .Y(new_n18737));
  nand_5 g16389(.A(new_n18737), .B(new_n18699), .Y(new_n18738));
  nand_5 g16390(.A(new_n18738), .B(pi469), .Y(new_n18739));
  or_6   g16391(.A(new_n18738), .B(pi469), .Y(new_n18740));
  nand_5 g16392(.A(new_n18740), .B(new_n18739), .Y(new_n18741));
  xor_4  g16393(.A(new_n18741), .B(new_n5540), .Y(new_n18742));
  nor_5  g16394(.A(new_n18742), .B(new_n18736), .Y(new_n18743));
  nor_5  g16395(.A(new_n18743), .B(new_n18673), .Y(new_n18744));
  or_6   g16396(.A(new_n18741), .B(new_n5540), .Y(new_n18745));
  nand_5 g16397(.A(new_n18745), .B(new_n18739), .Y(new_n18746));
  nand_5 g16398(.A(new_n18746), .B(new_n18744), .Y(new_n18747));
  not_8  g16399(.A(new_n18747), .Y(new_n18748));
  nand_5 g16400(.A(new_n18748), .B(new_n18671), .Y(new_n18749));
  not_8  g16401(.A(new_n18749), .Y(new_n18750));
  nand_5 g16402(.A(new_n18743), .B(new_n18673), .Y(new_n18751));
  and_6  g16403(.A(new_n18751), .B(new_n18740), .Y(new_n18752));
  or_6   g16404(.A(new_n18752), .B(new_n18744), .Y(new_n18753));
  nor_5  g16405(.A(new_n18748), .B(new_n18671), .Y(new_n18754));
  nand_5 g16406(.A(new_n5547), .B(pi397), .Y(new_n18755));
  nor_5  g16407(.A(new_n18755), .B(new_n18754), .Y(new_n18756));
  and_6  g16408(.A(new_n18756), .B(new_n18753), .Y(new_n18757));
  nor_5  g16409(.A(new_n18757), .B(new_n18750), .Y(new_n18758));
  nand_5 g16410(.A(new_n14252), .B(pi716), .Y(new_n18759));
  nand_5 g16411(.A(pi769), .B(new_n4511), .Y(new_n18760));
  nand_5 g16412(.A(new_n18760), .B(new_n18759), .Y(new_n18761));
  xor_4  g16413(.A(new_n18761), .B(new_n11091), .Y(new_n18762));
  nand_5 g16414(.A(new_n4374), .B(new_n14258), .Y(new_n18763));
  nand_5 g16415(.A(new_n13155), .B(new_n13149), .Y(new_n18764));
  nand_5 g16416(.A(new_n13156), .B(pi125), .Y(new_n18765));
  nand_5 g16417(.A(new_n18765), .B(new_n18764), .Y(new_n18766));
  nor_5  g16418(.A(new_n13153), .B(pi635), .Y(new_n18767));
  nand_5 g16419(.A(new_n13153), .B(pi635), .Y(new_n18768));
  nand_5 g16420(.A(new_n18768), .B(new_n10742), .Y(new_n18769));
  not_8  g16421(.A(new_n18769), .Y(new_n18770));
  nor_5  g16422(.A(new_n18770), .B(new_n18767), .Y(new_n18771));
  nand_5 g16423(.A(pi712), .B(pi265), .Y(new_n18772));
  nand_5 g16424(.A(new_n9512), .B(new_n11101), .Y(new_n18773));
  nand_5 g16425(.A(new_n18773), .B(new_n18772), .Y(new_n18774));
  xor_4  g16426(.A(new_n18774), .B(new_n18771), .Y(new_n18775));
  not_8  g16427(.A(new_n18775), .Y(new_n18776));
  nand_5 g16428(.A(new_n18776), .B(new_n18766), .Y(new_n18777));
  xor_4  g16429(.A(new_n18775), .B(new_n18766), .Y(new_n18778));
  or_6   g16430(.A(new_n18778), .B(new_n10740), .Y(new_n18779));
  nand_5 g16431(.A(new_n18779), .B(new_n18777), .Y(new_n18780));
  nand_5 g16432(.A(new_n9554), .B(new_n10647), .Y(new_n18781));
  nand_5 g16433(.A(pi530), .B(pi332), .Y(new_n18782));
  nand_5 g16434(.A(new_n18782), .B(new_n18781), .Y(new_n18783));
  not_8  g16435(.A(new_n18771), .Y(new_n18784));
  nand_5 g16436(.A(new_n18772), .B(new_n18784), .Y(new_n18785));
  nand_5 g16437(.A(new_n18785), .B(new_n18773), .Y(new_n18786));
  xor_4  g16438(.A(new_n18786), .B(new_n18783), .Y(new_n18787));
  nand_5 g16439(.A(new_n18787), .B(new_n18780), .Y(new_n18788));
  or_6   g16440(.A(new_n18787), .B(new_n18780), .Y(new_n18789));
  nand_5 g16441(.A(new_n18789), .B(pi473), .Y(new_n18790));
  nand_5 g16442(.A(new_n18790), .B(new_n18788), .Y(new_n18791));
  nand_5 g16443(.A(new_n18786), .B(new_n18782), .Y(new_n18792));
  nand_5 g16444(.A(new_n18792), .B(new_n18781), .Y(new_n18793));
  nand_5 g16445(.A(pi772), .B(pi459), .Y(new_n18794));
  nand_5 g16446(.A(new_n11096), .B(new_n14261), .Y(new_n18795));
  nand_5 g16447(.A(new_n18795), .B(new_n18794), .Y(new_n18796));
  xor_4  g16448(.A(new_n18796), .B(new_n18793), .Y(new_n18797));
  or_6   g16449(.A(new_n18797), .B(new_n18791), .Y(new_n18798));
  nand_5 g16450(.A(new_n18798), .B(pi505), .Y(new_n18799));
  nand_5 g16451(.A(new_n18797), .B(new_n18791), .Y(new_n18800));
  nand_5 g16452(.A(new_n18800), .B(new_n18799), .Y(new_n18801));
  nand_5 g16453(.A(pi368), .B(pi275), .Y(new_n18802));
  nand_5 g16454(.A(new_n18802), .B(new_n18763), .Y(new_n18803));
  nand_5 g16455(.A(new_n18794), .B(new_n18793), .Y(new_n18804));
  nand_5 g16456(.A(new_n18804), .B(new_n18795), .Y(new_n18805));
  nor_5  g16457(.A(new_n18805), .B(new_n7257), .Y(new_n18806));
  nand_5 g16458(.A(new_n18805), .B(new_n7257), .Y(new_n18807));
  not_8  g16459(.A(new_n18807), .Y(new_n18808));
  nor_5  g16460(.A(new_n18808), .B(new_n18806), .Y(new_n18809));
  xor_4  g16461(.A(new_n18809), .B(new_n18803), .Y(new_n18810));
  nor_5  g16462(.A(new_n18810), .B(new_n18801), .Y(new_n18811));
  not_8  g16463(.A(new_n18811), .Y(new_n18812));
  nand_5 g16464(.A(new_n18812), .B(new_n18763), .Y(new_n18813));
  not_8  g16465(.A(new_n18813), .Y(new_n18814));
  nor_5  g16466(.A(new_n18812), .B(new_n18763), .Y(new_n18815));
  nor_5  g16467(.A(new_n18815), .B(new_n18808), .Y(new_n18816));
  nor_5  g16468(.A(new_n18816), .B(new_n18814), .Y(new_n18817));
  nand_5 g16469(.A(new_n18814), .B(new_n18806), .Y(new_n18818));
  nor_5  g16470(.A(new_n18808), .B(new_n18802), .Y(new_n18819));
  nand_5 g16471(.A(new_n18819), .B(new_n18812), .Y(new_n18820));
  nand_5 g16472(.A(new_n18820), .B(new_n18818), .Y(new_n18821));
  nor_5  g16473(.A(new_n18821), .B(new_n18817), .Y(new_n18822));
  nand_5 g16474(.A(new_n18822), .B(new_n18762), .Y(new_n18823));
  not_8  g16475(.A(new_n18823), .Y(new_n18824));
  nand_5 g16476(.A(new_n18761), .B(new_n11091), .Y(new_n18825));
  nand_5 g16477(.A(new_n14252), .B(new_n4511), .Y(new_n18826));
  nand_5 g16478(.A(new_n18826), .B(new_n18825), .Y(new_n18827));
  or_6   g16479(.A(new_n18827), .B(new_n18817), .Y(new_n18828));
  nor_5  g16480(.A(new_n18828), .B(new_n18824), .Y(new_n18829));
  xor_4  g16481(.A(new_n18829), .B(new_n18758), .Y(new_n18830));
  not_8  g16482(.A(new_n18830), .Y(new_n18831));
  or_6   g16483(.A(new_n18826), .B(pi534), .Y(new_n18832));
  or_6   g16484(.A(new_n18832), .B(new_n18821), .Y(new_n18833));
  nand_5 g16485(.A(new_n18827), .B(new_n18817), .Y(new_n18834));
  nand_5 g16486(.A(new_n18834), .B(new_n18833), .Y(new_n18835));
  or_6   g16487(.A(new_n18835), .B(new_n18829), .Y(new_n18836));
  nor_5  g16488(.A(new_n5547), .B(pi397), .Y(new_n18837));
  nand_5 g16489(.A(new_n18837), .B(new_n18747), .Y(new_n18838));
  not_8  g16490(.A(new_n18838), .Y(new_n18839));
  nand_5 g16491(.A(new_n18755), .B(new_n5544), .Y(new_n18840));
  nor_5  g16492(.A(new_n18840), .B(new_n18753), .Y(new_n18841));
  nor_5  g16493(.A(new_n18841), .B(new_n18839), .Y(new_n18842));
  nand_5 g16494(.A(new_n18842), .B(new_n18758), .Y(new_n18843));
  not_8  g16495(.A(new_n18843), .Y(new_n18844));
  and_6  g16496(.A(new_n18844), .B(new_n18836), .Y(new_n18845));
  xor_4  g16497(.A(new_n18844), .B(new_n18836), .Y(new_n18846));
  not_8  g16498(.A(new_n18846), .Y(new_n18847));
  xnor_4 g16499(.A(new_n18810), .B(new_n18801), .Y(new_n18848));
  xor_4  g16500(.A(new_n18742), .B(new_n18736), .Y(new_n18849));
  or_6   g16501(.A(new_n18849), .B(new_n18848), .Y(new_n18850));
  xnor_4 g16502(.A(new_n18734), .B(new_n18703), .Y(new_n18851));
  and_6  g16503(.A(new_n18800), .B(new_n18798), .Y(new_n18852));
  xor_4  g16504(.A(new_n18852), .B(new_n8005), .Y(new_n18853));
  not_8  g16505(.A(new_n18853), .Y(new_n18854));
  nor_5  g16506(.A(new_n18854), .B(new_n18851), .Y(new_n18855));
  nand_5 g16507(.A(new_n18789), .B(new_n18788), .Y(new_n18856));
  xor_4  g16508(.A(new_n18856), .B(pi473), .Y(new_n18857));
  xor_4  g16509(.A(new_n18731), .B(new_n18730), .Y(new_n18858));
  not_8  g16510(.A(new_n18858), .Y(new_n18859));
  nor_5  g16511(.A(new_n18859), .B(new_n18857), .Y(new_n18860));
  xor_4  g16512(.A(new_n18858), .B(new_n18857), .Y(new_n18861));
  xor_4  g16513(.A(new_n18728), .B(new_n18708), .Y(new_n18862));
  xor_4  g16514(.A(new_n18778), .B(pi248), .Y(new_n18863));
  nand_5 g16515(.A(new_n18863), .B(new_n18862), .Y(new_n18864));
  xor_4  g16516(.A(new_n18725), .B(new_n18724), .Y(new_n18865));
  nor_5  g16517(.A(new_n18865), .B(new_n13157), .Y(new_n18866));
  xnor_4 g16518(.A(new_n18865), .B(new_n13157), .Y(new_n18867));
  xnor_4 g16519(.A(new_n18722), .B(new_n18721), .Y(new_n18868));
  or_6   g16520(.A(new_n18868), .B(new_n6596), .Y(new_n18869));
  xor_4  g16521(.A(new_n18719), .B(new_n18716), .Y(new_n18870));
  nand_5 g16522(.A(new_n18870), .B(new_n6597), .Y(new_n18871));
  xor_4  g16523(.A(new_n18870), .B(new_n6630), .Y(new_n18872));
  nor_5  g16524(.A(new_n16890), .B(new_n6598), .Y(new_n18873));
  nor_5  g16525(.A(new_n16895), .B(new_n16891), .Y(new_n18874));
  nor_5  g16526(.A(new_n18874), .B(new_n18873), .Y(new_n18875));
  or_6   g16527(.A(new_n18875), .B(new_n18872), .Y(new_n18876));
  nand_5 g16528(.A(new_n18876), .B(new_n18871), .Y(new_n18877));
  not_8  g16529(.A(new_n18877), .Y(new_n18878));
  xor_4  g16530(.A(new_n18868), .B(new_n6596), .Y(new_n18879));
  nand_5 g16531(.A(new_n18879), .B(new_n18878), .Y(new_n18880));
  nand_5 g16532(.A(new_n18880), .B(new_n18869), .Y(new_n18881));
  nor_5  g16533(.A(new_n18881), .B(new_n18867), .Y(new_n18882));
  or_6   g16534(.A(new_n18882), .B(new_n18866), .Y(new_n18883));
  xnor_4 g16535(.A(new_n18863), .B(new_n18862), .Y(new_n18884));
  or_6   g16536(.A(new_n18884), .B(new_n18883), .Y(new_n18885));
  nand_5 g16537(.A(new_n18885), .B(new_n18864), .Y(new_n18886));
  nor_5  g16538(.A(new_n18886), .B(new_n18861), .Y(new_n18887));
  or_6   g16539(.A(new_n18887), .B(new_n18860), .Y(new_n18888));
  xor_4  g16540(.A(new_n18853), .B(new_n18851), .Y(new_n18889));
  nor_5  g16541(.A(new_n18889), .B(new_n18888), .Y(new_n18890));
  or_6   g16542(.A(new_n18890), .B(new_n18855), .Y(new_n18891));
  xor_4  g16543(.A(new_n18849), .B(new_n18848), .Y(new_n18892));
  nand_5 g16544(.A(new_n18892), .B(new_n18891), .Y(new_n18893));
  nand_5 g16545(.A(new_n18893), .B(new_n18850), .Y(new_n18894));
  nand_5 g16546(.A(new_n18753), .B(new_n18747), .Y(new_n18895));
  xor_4  g16547(.A(new_n18895), .B(pi397), .Y(new_n18896));
  xor_4  g16548(.A(new_n18896), .B(new_n5549), .Y(new_n18897));
  not_8  g16549(.A(new_n18897), .Y(new_n18898));
  nor_5  g16550(.A(new_n18898), .B(new_n18894), .Y(new_n18899));
  xor_4  g16551(.A(new_n18897), .B(new_n18894), .Y(new_n18900));
  xor_4  g16552(.A(new_n18822), .B(new_n18762), .Y(new_n18901));
  nor_5  g16553(.A(new_n18901), .B(new_n18900), .Y(new_n18902));
  or_6   g16554(.A(new_n18902), .B(new_n18899), .Y(new_n18903));
  nor_5  g16555(.A(new_n18903), .B(new_n18847), .Y(new_n18904));
  nor_5  g16556(.A(new_n18904), .B(new_n18845), .Y(new_n18905));
  xor_4  g16557(.A(new_n18905), .B(new_n18831), .Y(po0268));
  not_8  g16558(.A(new_n11993), .Y(new_n18907));
  nor_5  g16559(.A(new_n12011), .B(new_n18907), .Y(new_n18908));
  nor_5  g16560(.A(new_n12068), .B(new_n12012), .Y(new_n18909));
  or_6   g16561(.A(new_n18909), .B(new_n18908), .Y(new_n18910));
  nor_5  g16562(.A(new_n12008), .B(new_n7381), .Y(new_n18911));
  nor_5  g16563(.A(new_n7308), .B(new_n7294), .Y(new_n18912));
  and_6  g16564(.A(new_n18912), .B(new_n12009), .Y(new_n18913));
  nor_5  g16565(.A(new_n7307), .B(new_n7296), .Y(new_n18914));
  nand_5 g16566(.A(new_n18914), .B(new_n12008), .Y(new_n18915));
  or_6   g16567(.A(new_n12009), .B(new_n7380), .Y(new_n18916));
  nand_5 g16568(.A(new_n18916), .B(new_n18915), .Y(new_n18917));
  nor_5  g16569(.A(new_n18917), .B(new_n18913), .Y(new_n18918));
  not_8  g16570(.A(new_n18918), .Y(new_n18919));
  nor_5  g16571(.A(new_n18919), .B(new_n18911), .Y(new_n18920));
  nand_5 g16572(.A(pi323), .B(pi072), .Y(new_n18921));
  nand_5 g16573(.A(new_n17659), .B(new_n7187), .Y(new_n18922));
  nand_5 g16574(.A(new_n18922), .B(new_n16941), .Y(new_n18923));
  nand_5 g16575(.A(new_n18923), .B(new_n18921), .Y(new_n18924));
  or_6   g16576(.A(new_n18924), .B(new_n11987), .Y(new_n18925));
  nor_5  g16577(.A(new_n18922), .B(new_n16941), .Y(new_n18926));
  nand_5 g16578(.A(new_n18926), .B(new_n11990), .Y(new_n18927));
  nand_5 g16579(.A(new_n18927), .B(new_n18925), .Y(new_n18928));
  nor_5  g16580(.A(new_n18921), .B(pi068), .Y(new_n18929));
  nand_5 g16581(.A(new_n18929), .B(new_n11987), .Y(new_n18930));
  not_8  g16582(.A(new_n11990), .Y(new_n18931));
  nand_5 g16583(.A(new_n18924), .B(new_n18931), .Y(new_n18932));
  nand_5 g16584(.A(new_n18932), .B(new_n18930), .Y(new_n18933));
  or_6   g16585(.A(new_n18933), .B(new_n18928), .Y(new_n18934));
  xor_4  g16586(.A(new_n18934), .B(new_n18920), .Y(new_n18935));
  nand_5 g16587(.A(new_n18935), .B(new_n18910), .Y(new_n18936));
  not_8  g16588(.A(new_n18936), .Y(new_n18937));
  nand_5 g16589(.A(new_n18918), .B(new_n7381), .Y(new_n18938));
  not_8  g16590(.A(new_n18938), .Y(new_n18939));
  xor_4  g16591(.A(new_n18939), .B(new_n18928), .Y(new_n18940));
  nand_5 g16592(.A(new_n18940), .B(new_n18937), .Y(new_n18941));
  nor_5  g16593(.A(new_n18934), .B(new_n18920), .Y(new_n18942));
  nor_5  g16594(.A(new_n18940), .B(new_n18942), .Y(new_n18943));
  nand_5 g16595(.A(new_n18943), .B(new_n18936), .Y(new_n18944));
  nand_5 g16596(.A(new_n18944), .B(new_n18941), .Y(po0270));
  nand_5 g16597(.A(new_n17667), .B(pi097), .Y(new_n18946));
  nand_5 g16598(.A(new_n18946), .B(new_n17665), .Y(new_n18947));
  nand_5 g16599(.A(pi381), .B(new_n17659), .Y(new_n18948));
  nand_5 g16600(.A(new_n17663), .B(new_n17660), .Y(new_n18949));
  nand_5 g16601(.A(new_n18949), .B(new_n18948), .Y(new_n18950));
  xor_4  g16602(.A(new_n18950), .B(new_n18947), .Y(new_n18951));
  nand_5 g16603(.A(new_n18951), .B(new_n18920), .Y(new_n18952));
  nor_5  g16604(.A(new_n17669), .B(new_n12011), .Y(new_n18953));
  nor_5  g16605(.A(new_n17673), .B(new_n17670), .Y(new_n18954));
  nor_5  g16606(.A(new_n18954), .B(new_n18953), .Y(new_n18955));
  xor_4  g16607(.A(new_n18951), .B(new_n18920), .Y(new_n18956));
  nand_5 g16608(.A(new_n18956), .B(new_n18955), .Y(new_n18957));
  nand_5 g16609(.A(new_n18957), .B(new_n18952), .Y(new_n18958));
  nand_5 g16610(.A(new_n18950), .B(new_n18947), .Y(new_n18959));
  xor_4  g16611(.A(new_n18959), .B(new_n18939), .Y(new_n18960));
  not_8  g16612(.A(new_n18960), .Y(new_n18961));
  xor_4  g16613(.A(new_n18961), .B(new_n18958), .Y(po0271));
  xor_4  g16614(.A(new_n15795), .B(new_n15793), .Y(po0272));
  nand_5 g16615(.A(new_n14809), .B(new_n10630), .Y(new_n18964));
  nand_5 g16616(.A(new_n14810), .B(new_n14794), .Y(new_n18965));
  and_6  g16617(.A(new_n18965), .B(new_n18964), .Y(new_n18966));
  not_8  g16618(.A(new_n10469), .Y(new_n18967));
  nand_5 g16619(.A(new_n14804), .B(new_n18967), .Y(new_n18968));
  nor_5  g16620(.A(new_n18968), .B(new_n18966), .Y(po0273));
  xor_4  g16621(.A(new_n12378), .B(new_n8910), .Y(po0274));
  xnor_4 g16622(.A(new_n8432), .B(new_n8395), .Y(po0275));
  xor_4  g16623(.A(new_n18366), .B(new_n18345), .Y(po0276));
  nand_5 g16624(.A(new_n13939), .B(new_n4751), .Y(new_n18973));
  nor_5  g16625(.A(new_n13939), .B(new_n4751), .Y(new_n18974));
  not_8  g16626(.A(new_n18974), .Y(new_n18975));
  nand_5 g16627(.A(new_n18975), .B(new_n18973), .Y(new_n18976));
  xor_4  g16628(.A(new_n18976), .B(new_n13718), .Y(new_n18977));
  or_6   g16629(.A(new_n13277), .B(new_n5870), .Y(new_n18978));
  xor_4  g16630(.A(new_n13277), .B(new_n5870), .Y(new_n18979));
  not_8  g16631(.A(new_n13262), .Y(new_n18980));
  nor_5  g16632(.A(new_n17679), .B(new_n18980), .Y(new_n18981));
  nor_5  g16633(.A(new_n17680), .B(new_n5875), .Y(new_n18982));
  or_6   g16634(.A(new_n18982), .B(new_n18981), .Y(new_n18983));
  nand_5 g16635(.A(new_n18983), .B(new_n18979), .Y(new_n18984));
  nand_5 g16636(.A(new_n18984), .B(new_n18978), .Y(new_n18985));
  nor_5  g16637(.A(new_n18985), .B(new_n16366), .Y(new_n18986));
  xor_4  g16638(.A(new_n18985), .B(new_n5866), .Y(new_n18987));
  nor_5  g16639(.A(new_n18987), .B(new_n13950), .Y(new_n18988));
  or_6   g16640(.A(new_n18988), .B(new_n18986), .Y(new_n18989));
  nor_5  g16641(.A(new_n18989), .B(new_n13959), .Y(new_n18990));
  xnor_4 g16642(.A(new_n18989), .B(new_n13959), .Y(new_n18991));
  nor_5  g16643(.A(new_n18991), .B(new_n5865), .Y(new_n18992));
  or_6   g16644(.A(new_n18992), .B(new_n18990), .Y(new_n18993));
  nand_5 g16645(.A(new_n18993), .B(new_n13949), .Y(new_n18994));
  xor_4  g16646(.A(new_n18993), .B(new_n13948), .Y(new_n18995));
  or_6   g16647(.A(new_n18995), .B(new_n5900), .Y(new_n18996));
  nand_5 g16648(.A(new_n18996), .B(new_n18994), .Y(new_n18997));
  nor_5  g16649(.A(new_n18997), .B(new_n5907), .Y(new_n18998));
  xor_4  g16650(.A(new_n18997), .B(new_n5906), .Y(new_n18999));
  nor_5  g16651(.A(new_n18999), .B(new_n13944), .Y(new_n19000));
  or_6   g16652(.A(new_n19000), .B(new_n18998), .Y(new_n19001));
  nor_5  g16653(.A(new_n19001), .B(new_n13943), .Y(new_n19002));
  xor_4  g16654(.A(new_n19001), .B(new_n13942), .Y(new_n19003));
  nor_5  g16655(.A(new_n19003), .B(new_n5924), .Y(new_n19004));
  nor_5  g16656(.A(new_n19004), .B(new_n19002), .Y(new_n19005));
  nand_5 g16657(.A(new_n19005), .B(new_n13941), .Y(new_n19006));
  xor_4  g16658(.A(new_n19005), .B(new_n13940), .Y(new_n19007));
  or_6   g16659(.A(new_n19007), .B(new_n13710), .Y(new_n19008));
  nand_5 g16660(.A(new_n19008), .B(new_n19006), .Y(new_n19009));
  xor_4  g16661(.A(new_n19007), .B(new_n13710), .Y(new_n19010));
  not_8  g16662(.A(new_n19010), .Y(new_n19011));
  xor_4  g16663(.A(new_n18999), .B(new_n13945), .Y(new_n19012));
  nand_5 g16664(.A(new_n19012), .B(new_n4953), .Y(new_n19013));
  xor_4  g16665(.A(new_n19012), .B(new_n4954), .Y(new_n19014));
  xor_4  g16666(.A(new_n18995), .B(new_n5899), .Y(new_n19015));
  nor_5  g16667(.A(new_n19015), .B(new_n4960), .Y(new_n19016));
  not_8  g16668(.A(new_n4960), .Y(new_n19017));
  xor_4  g16669(.A(new_n19015), .B(new_n19017), .Y(new_n19018));
  xor_4  g16670(.A(new_n18991), .B(new_n5865), .Y(new_n19019));
  xor_4  g16671(.A(new_n18987), .B(new_n13950), .Y(new_n19020));
  not_8  g16672(.A(new_n19020), .Y(new_n19021));
  or_6   g16673(.A(new_n17684), .B(new_n4996), .Y(new_n19022));
  nand_5 g16674(.A(new_n17685), .B(new_n17681), .Y(new_n19023));
  nand_5 g16675(.A(new_n19023), .B(new_n19022), .Y(new_n19024));
  nor_5  g16676(.A(new_n19024), .B(new_n4976), .Y(new_n19025));
  xnor_4 g16677(.A(new_n18983), .B(new_n18979), .Y(new_n19026));
  xor_4  g16678(.A(new_n19024), .B(new_n4975), .Y(new_n19027));
  nor_5  g16679(.A(new_n19027), .B(new_n19026), .Y(new_n19028));
  or_6   g16680(.A(new_n19028), .B(new_n19025), .Y(new_n19029));
  nand_5 g16681(.A(new_n19029), .B(new_n19021), .Y(new_n19030));
  xor_4  g16682(.A(new_n19029), .B(new_n19020), .Y(new_n19031));
  or_6   g16683(.A(new_n19031), .B(new_n4969), .Y(new_n19032));
  nand_5 g16684(.A(new_n19032), .B(new_n19030), .Y(new_n19033));
  and_6  g16685(.A(new_n19033), .B(new_n19019), .Y(new_n19034));
  nor_5  g16686(.A(new_n19033), .B(new_n19019), .Y(new_n19035));
  nor_5  g16687(.A(new_n19035), .B(new_n4966), .Y(new_n19036));
  nor_5  g16688(.A(new_n19036), .B(new_n19034), .Y(new_n19037));
  nor_5  g16689(.A(new_n19037), .B(new_n19018), .Y(new_n19038));
  nor_5  g16690(.A(new_n19038), .B(new_n19016), .Y(new_n19039));
  or_6   g16691(.A(new_n19039), .B(new_n19014), .Y(new_n19040));
  nand_5 g16692(.A(new_n19040), .B(new_n19013), .Y(new_n19041));
  nand_5 g16693(.A(new_n19041), .B(new_n4948), .Y(new_n19042));
  xor_4  g16694(.A(new_n19003), .B(new_n5925), .Y(new_n19043));
  xor_4  g16695(.A(new_n19041), .B(new_n4947), .Y(new_n19044));
  or_6   g16696(.A(new_n19044), .B(new_n19043), .Y(new_n19045));
  nand_5 g16697(.A(new_n19045), .B(new_n19042), .Y(new_n19046));
  nand_5 g16698(.A(new_n19046), .B(new_n19011), .Y(new_n19047));
  not_8  g16699(.A(new_n19047), .Y(new_n19048));
  xor_4  g16700(.A(new_n19046), .B(new_n19010), .Y(new_n19049));
  nor_5  g16701(.A(new_n19049), .B(new_n4944), .Y(new_n19050));
  nor_5  g16702(.A(new_n19050), .B(new_n19048), .Y(new_n19051));
  xor_4  g16703(.A(new_n19051), .B(new_n19009), .Y(new_n19052));
  not_8  g16704(.A(new_n19052), .Y(new_n19053));
  nor_5  g16705(.A(new_n19053), .B(new_n18977), .Y(new_n19054));
  nand_5 g16706(.A(new_n19051), .B(new_n19009), .Y(new_n19055));
  or_6   g16707(.A(new_n18976), .B(new_n13718), .Y(new_n19056));
  nand_5 g16708(.A(new_n19056), .B(new_n18975), .Y(new_n19057));
  nand_5 g16709(.A(new_n19057), .B(new_n19055), .Y(new_n19058));
  nor_5  g16710(.A(new_n19058), .B(new_n19054), .Y(po1287));
  nor_5  g16711(.A(new_n19051), .B(new_n19009), .Y(new_n19060));
  or_6   g16712(.A(new_n18973), .B(new_n13719), .Y(new_n19061));
  nor_5  g16713(.A(new_n19061), .B(new_n19060), .Y(new_n19062));
  nor_5  g16714(.A(new_n19057), .B(new_n19055), .Y(new_n19063));
  or_6   g16715(.A(new_n19063), .B(new_n19062), .Y(new_n19064));
  or_6   g16716(.A(new_n19064), .B(po1287), .Y(po0277));
  xnor_4 g16717(.A(new_n6914), .B(new_n6898), .Y(po0278));
  not_8  g16718(.A(new_n14399), .Y(new_n19067));
  nor_5  g16719(.A(new_n17320), .B(new_n15508), .Y(new_n19068));
  nor_5  g16720(.A(new_n17321), .B(new_n14409), .Y(new_n19069));
  or_6   g16721(.A(new_n19069), .B(new_n19068), .Y(new_n19070));
  or_6   g16722(.A(new_n19070), .B(new_n15506), .Y(new_n19071));
  not_8  g16723(.A(new_n14403), .Y(new_n19072));
  xor_4  g16724(.A(new_n19070), .B(new_n15506), .Y(new_n19073));
  nand_5 g16725(.A(new_n19073), .B(new_n19072), .Y(new_n19074));
  nand_5 g16726(.A(new_n19074), .B(new_n19071), .Y(new_n19075));
  nor_5  g16727(.A(new_n19075), .B(new_n19067), .Y(new_n19076));
  xor_4  g16728(.A(new_n19075), .B(new_n14399), .Y(new_n19077));
  nor_5  g16729(.A(new_n19077), .B(new_n16513), .Y(new_n19078));
  or_6   g16730(.A(new_n19078), .B(new_n19076), .Y(new_n19079));
  nand_5 g16731(.A(new_n19079), .B(new_n14394), .Y(new_n19080));
  xor_4  g16732(.A(new_n19079), .B(new_n14395), .Y(new_n19081));
  or_6   g16733(.A(new_n19081), .B(new_n16508), .Y(new_n19082));
  nand_5 g16734(.A(new_n19082), .B(new_n19080), .Y(new_n19083));
  xor_4  g16735(.A(new_n17718), .B(new_n14390), .Y(new_n19084));
  xor_4  g16736(.A(new_n19084), .B(new_n19083), .Y(po0279));
  nand_5 g16737(.A(new_n8641), .B(pi439), .Y(new_n19086));
  nand_5 g16738(.A(pi822), .B(new_n13485), .Y(new_n19087));
  xor_4  g16739(.A(pi822), .B(new_n13485), .Y(new_n19088));
  nand_5 g16740(.A(new_n8591), .B(pi100), .Y(new_n19089));
  xor_4  g16741(.A(pi557), .B(new_n7758), .Y(new_n19090));
  nand_5 g16742(.A(new_n8576), .B(pi117), .Y(new_n19091));
  nand_5 g16743(.A(new_n18003), .B(new_n17993), .Y(new_n19092));
  nand_5 g16744(.A(new_n19092), .B(new_n19091), .Y(new_n19093));
  nand_5 g16745(.A(new_n19093), .B(new_n19090), .Y(new_n19094));
  nand_5 g16746(.A(new_n19094), .B(new_n19089), .Y(new_n19095));
  nand_5 g16747(.A(new_n19095), .B(new_n19088), .Y(new_n19096));
  nand_5 g16748(.A(new_n19096), .B(new_n19087), .Y(new_n19097));
  xor_4  g16749(.A(pi768), .B(pi439), .Y(new_n19098));
  not_8  g16750(.A(new_n19098), .Y(new_n19099));
  nand_5 g16751(.A(new_n19099), .B(new_n19097), .Y(new_n19100));
  nand_5 g16752(.A(new_n19100), .B(new_n19086), .Y(new_n19101));
  nand_5 g16753(.A(new_n16177), .B(pi046), .Y(new_n19102));
  nand_5 g16754(.A(pi671), .B(new_n7751), .Y(new_n19103));
  nand_5 g16755(.A(new_n19103), .B(new_n19102), .Y(new_n19104));
  xor_4  g16756(.A(new_n19104), .B(new_n19101), .Y(new_n19105));
  nor_5  g16757(.A(new_n19105), .B(new_n3047), .Y(new_n19106));
  xor_4  g16758(.A(new_n19105), .B(new_n3048), .Y(new_n19107));
  xor_4  g16759(.A(new_n19098), .B(new_n19097), .Y(new_n19108));
  nand_5 g16760(.A(new_n19108), .B(new_n3053), .Y(new_n19109));
  xor_4  g16761(.A(new_n19095), .B(new_n19088), .Y(new_n19110));
  or_6   g16762(.A(new_n19110), .B(new_n3058), .Y(new_n19111));
  xor_4  g16763(.A(new_n19110), .B(new_n3058), .Y(new_n19112));
  xor_4  g16764(.A(new_n19093), .B(new_n19090), .Y(new_n19113));
  nand_5 g16765(.A(new_n19113), .B(new_n3063), .Y(new_n19114));
  not_8  g16766(.A(new_n19114), .Y(new_n19115));
  xnor_4 g16767(.A(new_n19113), .B(new_n3063), .Y(new_n19116));
  not_8  g16768(.A(new_n3066), .Y(new_n19117));
  nor_5  g16769(.A(new_n18004), .B(new_n19117), .Y(new_n19118));
  nor_5  g16770(.A(new_n18021), .B(new_n18005), .Y(new_n19119));
  nor_5  g16771(.A(new_n19119), .B(new_n19118), .Y(new_n19120));
  nor_5  g16772(.A(new_n19120), .B(new_n19116), .Y(new_n19121));
  nor_5  g16773(.A(new_n19121), .B(new_n19115), .Y(new_n19122));
  nand_5 g16774(.A(new_n19122), .B(new_n19112), .Y(new_n19123));
  nand_5 g16775(.A(new_n19123), .B(new_n19111), .Y(new_n19124));
  xor_4  g16776(.A(new_n19108), .B(new_n3053), .Y(new_n19125));
  nand_5 g16777(.A(new_n19125), .B(new_n19124), .Y(new_n19126));
  nand_5 g16778(.A(new_n19126), .B(new_n19109), .Y(new_n19127));
  nor_5  g16779(.A(new_n19127), .B(new_n19107), .Y(new_n19128));
  nor_5  g16780(.A(new_n19128), .B(new_n19106), .Y(new_n19129));
  xor_4  g16781(.A(pi537), .B(pi452), .Y(new_n19130));
  not_8  g16782(.A(new_n19130), .Y(new_n19131));
  nand_5 g16783(.A(new_n19103), .B(new_n19101), .Y(new_n19132));
  nand_5 g16784(.A(new_n19132), .B(new_n19102), .Y(new_n19133));
  xor_4  g16785(.A(new_n19133), .B(new_n19131), .Y(new_n19134));
  xor_4  g16786(.A(new_n19134), .B(new_n3045), .Y(new_n19135));
  xnor_4 g16787(.A(new_n19135), .B(new_n19129), .Y(po0280));
  xnor_4 g16788(.A(new_n13530), .B(new_n13509), .Y(po0281));
  nand_5 g16789(.A(new_n3327), .B(pi096), .Y(new_n19138));
  nand_5 g16790(.A(pi728), .B(new_n3262), .Y(new_n19139));
  xor_4  g16791(.A(pi728), .B(new_n3262), .Y(new_n19140));
  nand_5 g16792(.A(new_n18589), .B(new_n18587), .Y(new_n19141));
  nand_5 g16793(.A(new_n19141), .B(new_n18588), .Y(new_n19142));
  nand_5 g16794(.A(new_n19142), .B(new_n19140), .Y(new_n19143));
  nand_5 g16795(.A(new_n19143), .B(new_n19139), .Y(new_n19144));
  nand_5 g16796(.A(pi114), .B(new_n7590), .Y(new_n19145));
  nand_5 g16797(.A(new_n19145), .B(new_n19144), .Y(new_n19146));
  nand_5 g16798(.A(new_n19146), .B(new_n19138), .Y(new_n19147));
  not_8  g16799(.A(new_n7394), .Y(new_n19148));
  xor_4  g16800(.A(new_n19142), .B(new_n19140), .Y(new_n19149));
  not_8  g16801(.A(new_n19149), .Y(new_n19150));
  nand_5 g16802(.A(new_n19150), .B(new_n7489), .Y(new_n19151));
  not_8  g16803(.A(new_n19151), .Y(new_n19152));
  xor_4  g16804(.A(new_n19150), .B(new_n7489), .Y(new_n19153));
  not_8  g16805(.A(new_n19153), .Y(new_n19154));
  or_6   g16806(.A(new_n18591), .B(new_n7395), .Y(new_n19155));
  nand_5 g16807(.A(new_n18592), .B(new_n18584), .Y(new_n19156));
  nand_5 g16808(.A(new_n19156), .B(new_n19155), .Y(new_n19157));
  nor_5  g16809(.A(new_n19157), .B(new_n19154), .Y(new_n19158));
  nor_5  g16810(.A(new_n19158), .B(new_n19152), .Y(new_n19159));
  nand_5 g16811(.A(new_n19159), .B(new_n19148), .Y(new_n19160));
  not_8  g16812(.A(new_n19160), .Y(new_n19161));
  nand_5 g16813(.A(new_n19161), .B(new_n19147), .Y(new_n19162));
  nor_5  g16814(.A(new_n19159), .B(new_n19148), .Y(new_n19163));
  not_8  g16815(.A(new_n19163), .Y(new_n19164));
  not_8  g16816(.A(new_n19144), .Y(new_n19165));
  nor_5  g16817(.A(new_n19165), .B(new_n19138), .Y(new_n19166));
  nand_5 g16818(.A(new_n19166), .B(new_n19164), .Y(new_n19167));
  nand_5 g16819(.A(new_n19167), .B(new_n19162), .Y(new_n19168));
  nand_5 g16820(.A(new_n7388), .B(new_n7384), .Y(new_n19169));
  not_8  g16821(.A(new_n19169), .Y(new_n19170));
  nand_5 g16822(.A(new_n19170), .B(new_n19168), .Y(new_n19171));
  nor_5  g16823(.A(new_n19164), .B(new_n19147), .Y(new_n19172));
  nor_5  g16824(.A(new_n19145), .B(new_n19144), .Y(new_n19173));
  nand_5 g16825(.A(new_n19173), .B(new_n19160), .Y(new_n19174));
  not_8  g16826(.A(new_n19174), .Y(new_n19175));
  nor_5  g16827(.A(new_n19175), .B(new_n19172), .Y(new_n19176));
  not_8  g16828(.A(new_n19176), .Y(new_n19177));
  nor_5  g16829(.A(new_n19177), .B(new_n7389), .Y(new_n19178));
  and_6  g16830(.A(new_n19178), .B(new_n19171), .Y(new_n19179));
  nand_5 g16831(.A(new_n19168), .B(new_n7390), .Y(new_n19180));
  nand_5 g16832(.A(new_n7391), .B(new_n7384), .Y(new_n19181));
  or_6   g16833(.A(new_n19181), .B(new_n19176), .Y(new_n19182));
  nand_5 g16834(.A(new_n19182), .B(new_n19180), .Y(new_n19183));
  nor_5  g16835(.A(new_n19183), .B(new_n19179), .Y(po0282));
  xor_4  g16836(.A(new_n10966), .B(pi193), .Y(new_n19185));
  nand_5 g16837(.A(pi440), .B(new_n10711), .Y(new_n19186));
  nand_5 g16838(.A(new_n15597), .B(new_n15581), .Y(new_n19187));
  nand_5 g16839(.A(new_n19187), .B(new_n19186), .Y(new_n19188));
  xor_4  g16840(.A(new_n19188), .B(new_n19185), .Y(new_n19189));
  not_8  g16841(.A(new_n19189), .Y(new_n19190));
  or_6   g16842(.A(new_n15601), .B(new_n15191), .Y(new_n19191));
  xor_4  g16843(.A(new_n15601), .B(new_n15191), .Y(new_n19192));
  nor_5  g16844(.A(new_n14061), .B(new_n13800), .Y(new_n19193));
  nand_5 g16845(.A(new_n19193), .B(new_n13803), .Y(new_n19194));
  xor_4  g16846(.A(new_n19193), .B(new_n13809), .Y(new_n19195));
  or_6   g16847(.A(new_n19195), .B(new_n14062), .Y(new_n19196));
  nand_5 g16848(.A(new_n19196), .B(new_n19194), .Y(new_n19197));
  or_6   g16849(.A(new_n19197), .B(new_n13794), .Y(new_n19198));
  nand_5 g16850(.A(new_n19197), .B(new_n13794), .Y(new_n19199));
  nand_5 g16851(.A(new_n19199), .B(new_n14056), .Y(new_n19200));
  nand_5 g16852(.A(new_n19200), .B(new_n19198), .Y(new_n19201));
  nor_5  g16853(.A(new_n19201), .B(new_n14043), .Y(new_n19202));
  xnor_4 g16854(.A(new_n19201), .B(new_n14043), .Y(new_n19203));
  nor_5  g16855(.A(new_n19203), .B(new_n13791), .Y(new_n19204));
  nor_5  g16856(.A(new_n19204), .B(new_n19202), .Y(new_n19205));
  nand_5 g16857(.A(new_n19205), .B(new_n15605), .Y(new_n19206));
  xnor_4 g16858(.A(new_n19205), .B(new_n15605), .Y(new_n19207));
  or_6   g16859(.A(new_n19207), .B(new_n15201), .Y(new_n19208));
  nand_5 g16860(.A(new_n19208), .B(new_n19206), .Y(new_n19209));
  and_6  g16861(.A(new_n19209), .B(new_n15603), .Y(new_n19210));
  xnor_4 g16862(.A(new_n19209), .B(new_n15603), .Y(new_n19211));
  nor_5  g16863(.A(new_n19211), .B(new_n15197), .Y(new_n19212));
  nor_5  g16864(.A(new_n19212), .B(new_n19210), .Y(new_n19213));
  nand_5 g16865(.A(new_n19213), .B(new_n19192), .Y(new_n19214));
  nand_5 g16866(.A(new_n19214), .B(new_n19191), .Y(new_n19215));
  nand_5 g16867(.A(new_n19215), .B(new_n15599), .Y(new_n19216));
  xor_4  g16868(.A(new_n19215), .B(new_n15599), .Y(new_n19217));
  nand_5 g16869(.A(new_n19217), .B(new_n15187), .Y(new_n19218));
  nand_5 g16870(.A(new_n19218), .B(new_n19216), .Y(new_n19219));
  xor_4  g16871(.A(new_n19219), .B(new_n19190), .Y(new_n19220));
  xnor_4 g16872(.A(new_n19220), .B(new_n15159), .Y(po0283));
  xnor_4 g16873(.A(new_n14890), .B(new_n14889), .Y(po0284));
  xor_4  g16874(.A(new_n15904), .B(new_n15903), .Y(po0285));
  xnor_4 g16875(.A(new_n10627), .B(new_n10572), .Y(po0286));
  nand_5 g16876(.A(new_n5031), .B(new_n6972), .Y(new_n19225));
  nand_5 g16877(.A(new_n18486), .B(new_n18484), .Y(new_n19226));
  and_6  g16878(.A(new_n19226), .B(new_n19225), .Y(new_n19227));
  xor_4  g16879(.A(pi731), .B(new_n5021), .Y(new_n19228));
  xor_4  g16880(.A(new_n19228), .B(new_n19227), .Y(new_n19229));
  xor_4  g16881(.A(new_n19229), .B(new_n2414), .Y(new_n19230));
  nand_5 g16882(.A(new_n18498), .B(new_n18493), .Y(new_n19231));
  and_6  g16883(.A(new_n18490), .B(new_n2363), .Y(new_n19232));
  nor_5  g16884(.A(new_n19232), .B(new_n19226), .Y(new_n19233));
  nor_5  g16885(.A(new_n18484), .B(new_n2363), .Y(new_n19234));
  nand_5 g16886(.A(new_n18489), .B(new_n19234), .Y(new_n19235));
  nand_5 g16887(.A(new_n19235), .B(new_n2423), .Y(new_n19236));
  nor_5  g16888(.A(new_n19236), .B(new_n19233), .Y(new_n19237));
  nand_5 g16889(.A(new_n19237), .B(new_n19231), .Y(new_n19238));
  xor_4  g16890(.A(new_n19238), .B(new_n19230), .Y(new_n19239));
  xor_4  g16891(.A(pi294), .B(pi204), .Y(new_n19240));
  nand_5 g16892(.A(new_n18481), .B(new_n3641), .Y(new_n19241));
  nand_5 g16893(.A(new_n19241), .B(new_n18482), .Y(new_n19242));
  xor_4  g16894(.A(new_n19242), .B(new_n19240), .Y(new_n19243));
  xor_4  g16895(.A(new_n19243), .B(new_n19239), .Y(new_n19244));
  or_6   g16896(.A(new_n18483), .B(new_n7059), .Y(new_n19245));
  and_6  g16897(.A(new_n19245), .B(new_n19231), .Y(new_n19246));
  not_8  g16898(.A(new_n18493), .Y(new_n19247));
  not_8  g16899(.A(new_n18500), .Y(new_n19248));
  nand_5 g16900(.A(new_n19248), .B(new_n19247), .Y(new_n19249));
  nand_5 g16901(.A(new_n18483), .B(pi238), .Y(new_n19250));
  nand_5 g16902(.A(new_n19250), .B(new_n19249), .Y(new_n19251));
  nor_5  g16903(.A(new_n19251), .B(new_n19246), .Y(new_n19252));
  nor_5  g16904(.A(new_n19248), .B(new_n18493), .Y(new_n19253));
  nand_5 g16905(.A(new_n18483), .B(new_n3641), .Y(new_n19254));
  nor_5  g16906(.A(new_n19254), .B(new_n19253), .Y(new_n19255));
  nor_5  g16907(.A(new_n19255), .B(new_n19252), .Y(new_n19256));
  xnor_4 g16908(.A(new_n19256), .B(new_n19244), .Y(po0287));
  xor_4  g16909(.A(new_n13812), .B(new_n13797), .Y(po0288));
  xor_4  g16910(.A(new_n12647), .B(new_n12646), .Y(po0289));
  xnor_4 g16911(.A(new_n2802), .B(new_n2800), .Y(po0290));
  nor_5  g16912(.A(pi731), .B(pi276), .Y(new_n19261));
  nor_5  g16913(.A(new_n19228), .B(new_n19227), .Y(new_n19262));
  nor_5  g16914(.A(new_n19262), .B(new_n19261), .Y(new_n19263));
  xor_4  g16915(.A(pi454), .B(new_n8576), .Y(new_n19264));
  xor_4  g16916(.A(new_n19264), .B(new_n19263), .Y(new_n19265));
  or_6   g16917(.A(new_n19265), .B(new_n2448), .Y(new_n19266));
  xor_4  g16918(.A(new_n19265), .B(new_n2448), .Y(new_n19267));
  or_6   g16919(.A(new_n19229), .B(new_n2414), .Y(new_n19268));
  nand_5 g16920(.A(new_n19238), .B(new_n19230), .Y(new_n19269));
  nand_5 g16921(.A(new_n19269), .B(new_n19268), .Y(new_n19270));
  nand_5 g16922(.A(new_n19270), .B(new_n19267), .Y(new_n19271));
  nand_5 g16923(.A(new_n19271), .B(new_n19266), .Y(new_n19272));
  nor_5  g16924(.A(pi454), .B(pi228), .Y(new_n19273));
  nor_5  g16925(.A(new_n19264), .B(new_n19263), .Y(new_n19274));
  nor_5  g16926(.A(new_n19274), .B(new_n19273), .Y(new_n19275));
  not_8  g16927(.A(new_n19275), .Y(new_n19276));
  nand_5 g16928(.A(new_n8591), .B(new_n6963), .Y(new_n19277));
  nand_5 g16929(.A(pi557), .B(pi145), .Y(new_n19278));
  nand_5 g16930(.A(new_n19278), .B(new_n19277), .Y(new_n19279));
  xor_4  g16931(.A(new_n19279), .B(new_n19276), .Y(new_n19280));
  xor_4  g16932(.A(new_n19280), .B(new_n2456), .Y(new_n19281));
  xor_4  g16933(.A(new_n19281), .B(new_n19272), .Y(new_n19282));
  xor_4  g16934(.A(pi590), .B(new_n2909), .Y(new_n19283));
  nand_5 g16935(.A(pi328), .B(new_n2912), .Y(new_n19284));
  xor_4  g16936(.A(pi328), .B(new_n2912), .Y(new_n19285));
  nand_5 g16937(.A(new_n5287), .B(pi277), .Y(new_n19286));
  xor_4  g16938(.A(pi801), .B(new_n2960), .Y(new_n19287));
  nand_5 g16939(.A(pi313), .B(new_n2920), .Y(new_n19288));
  xor_4  g16940(.A(pi313), .B(new_n2920), .Y(new_n19289));
  nand_5 g16941(.A(pi832), .B(new_n5340), .Y(new_n19290));
  not_8  g16942(.A(new_n19290), .Y(new_n19291));
  nand_5 g16943(.A(new_n19291), .B(new_n19289), .Y(new_n19292));
  nand_5 g16944(.A(new_n19292), .B(new_n19288), .Y(new_n19293));
  nand_5 g16945(.A(new_n19293), .B(new_n19287), .Y(new_n19294));
  nand_5 g16946(.A(new_n19294), .B(new_n19286), .Y(new_n19295));
  nand_5 g16947(.A(new_n19295), .B(new_n19285), .Y(new_n19296));
  nand_5 g16948(.A(new_n19296), .B(new_n19284), .Y(new_n19297));
  xor_4  g16949(.A(new_n19297), .B(new_n19283), .Y(new_n19298));
  or_6   g16950(.A(new_n19298), .B(new_n19282), .Y(new_n19299));
  xor_4  g16951(.A(new_n19270), .B(new_n19267), .Y(new_n19300));
  xor_4  g16952(.A(new_n19295), .B(new_n19285), .Y(new_n19301));
  not_8  g16953(.A(new_n19301), .Y(new_n19302));
  nand_5 g16954(.A(new_n19302), .B(new_n19300), .Y(new_n19303));
  xor_4  g16955(.A(new_n19302), .B(new_n19300), .Y(new_n19304));
  xor_4  g16956(.A(new_n19293), .B(new_n19287), .Y(new_n19305));
  not_8  g16957(.A(new_n19305), .Y(new_n19306));
  nand_5 g16958(.A(new_n19306), .B(new_n19239), .Y(new_n19307));
  not_8  g16959(.A(new_n19292), .Y(new_n19308));
  nand_5 g16960(.A(new_n19308), .B(new_n19231), .Y(new_n19309));
  not_8  g16961(.A(new_n19289), .Y(new_n19310));
  nand_5 g16962(.A(new_n19291), .B(new_n18498), .Y(new_n19311));
  not_8  g16963(.A(new_n19311), .Y(new_n19312));
  nand_5 g16964(.A(new_n3815), .B(pi038), .Y(new_n19313));
  nor_5  g16965(.A(new_n19313), .B(new_n18498), .Y(new_n19314));
  nor_5  g16966(.A(new_n19314), .B(new_n19312), .Y(new_n19315));
  xor_4  g16967(.A(new_n19315), .B(new_n19247), .Y(new_n19316));
  nor_5  g16968(.A(new_n19316), .B(new_n19310), .Y(new_n19317));
  nand_5 g16969(.A(new_n19315), .B(new_n18493), .Y(new_n19318));
  nand_5 g16970(.A(new_n19318), .B(new_n19311), .Y(new_n19319));
  or_6   g16971(.A(new_n19319), .B(new_n19317), .Y(new_n19320));
  nand_5 g16972(.A(new_n19320), .B(new_n19309), .Y(new_n19321));
  xor_4  g16973(.A(new_n19306), .B(new_n19239), .Y(new_n19322));
  nand_5 g16974(.A(new_n19322), .B(new_n19321), .Y(new_n19323));
  nand_5 g16975(.A(new_n19323), .B(new_n19307), .Y(new_n19324));
  nand_5 g16976(.A(new_n19324), .B(new_n19304), .Y(new_n19325));
  nand_5 g16977(.A(new_n19325), .B(new_n19303), .Y(new_n19326));
  xor_4  g16978(.A(new_n19298), .B(new_n19282), .Y(new_n19327));
  nand_5 g16979(.A(new_n19327), .B(new_n19326), .Y(new_n19328));
  nand_5 g16980(.A(new_n19328), .B(new_n19299), .Y(new_n19329));
  nor_5  g16981(.A(new_n19280), .B(new_n2506), .Y(new_n19330));
  nor_5  g16982(.A(new_n19281), .B(new_n19272), .Y(new_n19331));
  nor_5  g16983(.A(new_n19331), .B(new_n19330), .Y(new_n19332));
  xor_4  g16984(.A(pi566), .B(new_n13485), .Y(new_n19333));
  nand_5 g16985(.A(new_n19278), .B(new_n19276), .Y(new_n19334));
  nand_5 g16986(.A(new_n19334), .B(new_n19277), .Y(new_n19335));
  xor_4  g16987(.A(new_n19335), .B(new_n19333), .Y(new_n19336));
  xor_4  g16988(.A(new_n19336), .B(new_n2461), .Y(new_n19337));
  xor_4  g16989(.A(new_n19337), .B(new_n19332), .Y(new_n19338));
  nand_5 g16990(.A(pi590), .B(new_n2909), .Y(new_n19339));
  nand_5 g16991(.A(new_n19297), .B(new_n19283), .Y(new_n19340));
  nand_5 g16992(.A(new_n19340), .B(new_n19339), .Y(new_n19341));
  nand_5 g16993(.A(pi709), .B(new_n16948), .Y(new_n19342));
  nand_5 g16994(.A(new_n11143), .B(pi229), .Y(new_n19343));
  nand_5 g16995(.A(new_n19343), .B(new_n19342), .Y(new_n19344));
  xnor_4 g16996(.A(new_n19344), .B(new_n19341), .Y(new_n19345));
  xor_4  g16997(.A(new_n19345), .B(new_n19338), .Y(new_n19346));
  xor_4  g16998(.A(new_n19346), .B(new_n19329), .Y(po0291));
  xor_4  g16999(.A(new_n12635), .B(new_n12634), .Y(po0292));
  xnor_4 g17000(.A(new_n19120), .B(new_n19116), .Y(po0293));
  xor_4  g17001(.A(new_n13131), .B(new_n4210), .Y(po0294));
  xor_4  g17002(.A(new_n19203), .B(new_n13791), .Y(po0295));
  nand_5 g17003(.A(new_n18608), .B(pi210), .Y(new_n19352));
  nand_5 g17004(.A(new_n19352), .B(new_n18607), .Y(new_n19353));
  nand_5 g17005(.A(new_n19353), .B(new_n8812), .Y(new_n19354));
  or_6   g17006(.A(new_n19353), .B(new_n8812), .Y(new_n19355));
  and_6  g17007(.A(new_n19355), .B(new_n19354), .Y(new_n19356));
  xor_4  g17008(.A(new_n19356), .B(pi826), .Y(new_n19357));
  not_8  g17009(.A(new_n19357), .Y(new_n19358));
  nand_5 g17010(.A(new_n18657), .B(pi587), .Y(new_n19359));
  nand_5 g17011(.A(new_n19359), .B(new_n18656), .Y(new_n19360));
  nand_5 g17012(.A(new_n19360), .B(new_n16677), .Y(new_n19361));
  or_6   g17013(.A(new_n19360), .B(new_n16677), .Y(new_n19362));
  nand_5 g17014(.A(new_n19362), .B(new_n19361), .Y(new_n19363));
  xor_4  g17015(.A(new_n19363), .B(pi572), .Y(new_n19364));
  xor_4  g17016(.A(new_n19364), .B(new_n19358), .Y(new_n19365));
  nand_5 g17017(.A(new_n18659), .B(new_n18651), .Y(new_n19366));
  or_6   g17018(.A(new_n18660), .B(new_n18610), .Y(new_n19367));
  nand_5 g17019(.A(new_n19367), .B(new_n19366), .Y(new_n19368));
  xor_4  g17020(.A(new_n19368), .B(new_n19365), .Y(po0296));
  xor_4  g17021(.A(pi724), .B(new_n2943), .Y(new_n19370));
  nand_5 g17022(.A(pi756), .B(new_n4341), .Y(new_n19371));
  xor_4  g17023(.A(pi756), .B(new_n4341), .Y(new_n19372));
  nand_5 g17024(.A(new_n2966), .B(pi171), .Y(new_n19373));
  xor_4  g17025(.A(pi263), .B(new_n2908), .Y(new_n19374));
  nand_5 g17026(.A(new_n2949), .B(pi414), .Y(new_n19375));
  xor_4  g17027(.A(pi766), .B(new_n2913), .Y(new_n19376));
  nand_5 g17028(.A(pi550), .B(new_n4347), .Y(new_n19377));
  xor_4  g17029(.A(pi550), .B(pi504), .Y(new_n19378));
  nand_5 g17030(.A(pi309), .B(new_n5026), .Y(new_n19379));
  nand_5 g17031(.A(new_n2956), .B(pi209), .Y(new_n19380));
  nand_5 g17032(.A(new_n19380), .B(new_n9081), .Y(new_n19381));
  nand_5 g17033(.A(new_n19381), .B(new_n19379), .Y(new_n19382));
  or_6   g17034(.A(new_n19382), .B(new_n19378), .Y(new_n19383));
  nand_5 g17035(.A(new_n19383), .B(new_n19377), .Y(new_n19384));
  nand_5 g17036(.A(new_n19384), .B(new_n19376), .Y(new_n19385));
  nand_5 g17037(.A(new_n19385), .B(new_n19375), .Y(new_n19386));
  nand_5 g17038(.A(new_n19386), .B(new_n19374), .Y(new_n19387));
  nand_5 g17039(.A(new_n19387), .B(new_n19373), .Y(new_n19388));
  nand_5 g17040(.A(new_n19388), .B(new_n19372), .Y(new_n19389));
  nand_5 g17041(.A(new_n19389), .B(new_n19371), .Y(new_n19390));
  xor_4  g17042(.A(new_n19390), .B(new_n19370), .Y(new_n19391));
  nor_5  g17043(.A(new_n19391), .B(new_n10339), .Y(new_n19392));
  not_8  g17044(.A(new_n10342), .Y(new_n19393));
  xor_4  g17045(.A(new_n19388), .B(new_n19372), .Y(new_n19394));
  nand_5 g17046(.A(new_n19394), .B(new_n19393), .Y(new_n19395));
  xor_4  g17047(.A(new_n19394), .B(new_n19393), .Y(new_n19396));
  not_8  g17048(.A(new_n19396), .Y(new_n19397));
  xor_4  g17049(.A(new_n19386), .B(new_n19374), .Y(new_n19398));
  not_8  g17050(.A(new_n19398), .Y(new_n19399));
  nand_5 g17051(.A(new_n19399), .B(new_n10344), .Y(new_n19400));
  xor_4  g17052(.A(new_n19384), .B(new_n19376), .Y(new_n19401));
  nand_5 g17053(.A(new_n19401), .B(new_n10349), .Y(new_n19402));
  xnor_4 g17054(.A(new_n19401), .B(new_n10349), .Y(new_n19403));
  xor_4  g17055(.A(new_n19382), .B(new_n19378), .Y(new_n19404));
  nor_5  g17056(.A(new_n19404), .B(new_n10354), .Y(new_n19405));
  xnor_4 g17057(.A(new_n19404), .B(new_n10354), .Y(new_n19406));
  and_6  g17058(.A(new_n19379), .B(new_n19380), .Y(new_n19407));
  xor_4  g17059(.A(new_n19407), .B(new_n10357), .Y(new_n19408));
  nand_5 g17060(.A(new_n9081), .B(pi062), .Y(new_n19409));
  nand_5 g17061(.A(new_n19409), .B(new_n10359), .Y(new_n19410));
  nand_5 g17062(.A(pi491), .B(new_n3020), .Y(new_n19411));
  nand_5 g17063(.A(new_n19411), .B(new_n10363), .Y(new_n19412));
  nand_5 g17064(.A(new_n19412), .B(new_n19410), .Y(new_n19413));
  nor_5  g17065(.A(new_n19413), .B(new_n19408), .Y(new_n19414));
  or_6   g17066(.A(new_n19407), .B(new_n10358), .Y(new_n19415));
  nand_5 g17067(.A(new_n19415), .B(pi491), .Y(new_n19416));
  nor_5  g17068(.A(new_n19416), .B(new_n19414), .Y(new_n19417));
  nand_5 g17069(.A(new_n10361), .B(pi062), .Y(new_n19418));
  nand_5 g17070(.A(new_n19413), .B(new_n19408), .Y(new_n19419));
  nor_5  g17071(.A(new_n19407), .B(pi491), .Y(new_n19420));
  nand_5 g17072(.A(new_n19420), .B(new_n19419), .Y(new_n19421));
  nand_5 g17073(.A(new_n19421), .B(new_n19418), .Y(new_n19422));
  nor_5  g17074(.A(new_n19422), .B(new_n19417), .Y(new_n19423));
  nor_5  g17075(.A(new_n19423), .B(new_n19406), .Y(new_n19424));
  or_6   g17076(.A(new_n19424), .B(new_n19405), .Y(new_n19425));
  or_6   g17077(.A(new_n19425), .B(new_n19403), .Y(new_n19426));
  nand_5 g17078(.A(new_n19426), .B(new_n19402), .Y(new_n19427));
  xor_4  g17079(.A(new_n19398), .B(new_n10344), .Y(new_n19428));
  or_6   g17080(.A(new_n19428), .B(new_n19427), .Y(new_n19429));
  nand_5 g17081(.A(new_n19429), .B(new_n19400), .Y(new_n19430));
  or_6   g17082(.A(new_n19430), .B(new_n19397), .Y(new_n19431));
  nand_5 g17083(.A(new_n19431), .B(new_n19395), .Y(new_n19432));
  xnor_4 g17084(.A(new_n19391), .B(new_n10339), .Y(new_n19433));
  nor_5  g17085(.A(new_n19433), .B(new_n19432), .Y(new_n19434));
  or_6   g17086(.A(new_n19434), .B(new_n19392), .Y(new_n19435));
  xor_4  g17087(.A(pi600), .B(new_n2939), .Y(new_n19436));
  nand_5 g17088(.A(pi724), .B(new_n2943), .Y(new_n19437));
  nand_5 g17089(.A(new_n19390), .B(new_n19370), .Y(new_n19438));
  nand_5 g17090(.A(new_n19438), .B(new_n19437), .Y(new_n19439));
  xnor_4 g17091(.A(new_n19439), .B(new_n19436), .Y(new_n19440));
  or_6   g17092(.A(new_n19440), .B(new_n10333), .Y(new_n19441));
  nand_5 g17093(.A(new_n19441), .B(new_n19435), .Y(new_n19442));
  nand_5 g17094(.A(new_n19440), .B(new_n10333), .Y(new_n19443));
  and_6  g17095(.A(new_n19443), .B(new_n19442), .Y(new_n19444));
  xor_4  g17096(.A(pi835), .B(new_n9154), .Y(new_n19445));
  nand_5 g17097(.A(pi600), .B(new_n2939), .Y(new_n19446));
  nand_5 g17098(.A(new_n19439), .B(new_n19436), .Y(new_n19447));
  nand_5 g17099(.A(new_n19447), .B(new_n19446), .Y(new_n19448));
  xnor_4 g17100(.A(new_n19448), .B(new_n19445), .Y(new_n19449));
  xor_4  g17101(.A(new_n19449), .B(new_n10329), .Y(new_n19450));
  xor_4  g17102(.A(new_n19450), .B(new_n19444), .Y(po0297));
  xor_4  g17103(.A(new_n12041), .B(new_n3864), .Y(po0298));
  xnor_4 g17104(.A(new_n10050), .B(new_n10048), .Y(po0299));
  xor_4  g17105(.A(new_n14442), .B(new_n14441), .Y(po0300));
  or_6   g17106(.A(new_n16171), .B(pi287), .Y(new_n19455));
  nand_5 g17107(.A(new_n16152), .B(new_n16145), .Y(new_n19456));
  nor_5  g17108(.A(new_n16121), .B(new_n16116), .Y(new_n19457));
  nor_5  g17109(.A(new_n16107), .B(pi268), .Y(new_n19458));
  nor_5  g17110(.A(new_n5077), .B(pi355), .Y(new_n19459));
  nand_5 g17111(.A(new_n5061), .B(new_n5051), .Y(new_n19460));
  nand_5 g17112(.A(new_n19460), .B(new_n5052), .Y(new_n19461));
  nor_5  g17113(.A(new_n19461), .B(new_n5078), .Y(new_n19462));
  nor_5  g17114(.A(new_n19462), .B(new_n19459), .Y(new_n19463));
  nor_5  g17115(.A(new_n19463), .B(new_n16113), .Y(new_n19464));
  or_6   g17116(.A(new_n19464), .B(new_n19458), .Y(new_n19465));
  nor_5  g17117(.A(new_n19465), .B(new_n16123), .Y(new_n19466));
  nor_5  g17118(.A(new_n19466), .B(new_n19457), .Y(new_n19467));
  nand_5 g17119(.A(new_n19467), .B(new_n16153), .Y(new_n19468));
  nand_5 g17120(.A(new_n19468), .B(new_n19456), .Y(new_n19469));
  nand_5 g17121(.A(new_n19469), .B(new_n16173), .Y(new_n19470));
  nand_5 g17122(.A(new_n19470), .B(new_n19455), .Y(new_n19471));
  xor_4  g17123(.A(new_n19471), .B(new_n16192), .Y(new_n19472));
  nand_5 g17124(.A(new_n19472), .B(new_n3263), .Y(new_n19473));
  not_8  g17125(.A(new_n3297), .Y(new_n19474));
  xor_4  g17126(.A(new_n19469), .B(new_n16172), .Y(new_n19475));
  or_6   g17127(.A(new_n19475), .B(new_n19474), .Y(new_n19476));
  xor_4  g17128(.A(new_n19467), .B(new_n16154), .Y(new_n19477));
  nor_5  g17129(.A(new_n19477), .B(new_n3265), .Y(new_n19478));
  xnor_4 g17130(.A(new_n19477), .B(new_n3265), .Y(new_n19479));
  xor_4  g17131(.A(new_n19465), .B(new_n16122), .Y(new_n19480));
  or_6   g17132(.A(new_n19480), .B(new_n3290), .Y(new_n19481));
  xor_4  g17133(.A(new_n19463), .B(new_n16113), .Y(new_n19482));
  or_6   g17134(.A(new_n19482), .B(new_n3284), .Y(new_n19483));
  xor_4  g17135(.A(new_n19482), .B(new_n3284), .Y(new_n19484));
  xnor_4 g17136(.A(new_n19461), .B(new_n5078), .Y(new_n19485));
  nor_5  g17137(.A(new_n19485), .B(new_n3276), .Y(new_n19486));
  xor_4  g17138(.A(new_n19485), .B(new_n3276), .Y(new_n19487));
  nand_5 g17139(.A(new_n5060), .B(new_n3269), .Y(new_n19488));
  or_6   g17140(.A(new_n5062), .B(new_n3269), .Y(new_n19489));
  and_6  g17141(.A(new_n19489), .B(new_n19488), .Y(new_n19490));
  xor_4  g17142(.A(new_n19490), .B(new_n3273), .Y(new_n19491));
  xor_4  g17143(.A(new_n19491), .B(new_n5053), .Y(po0679));
  nand_5 g17144(.A(po0679), .B(new_n3273), .Y(new_n19493));
  nor_5  g17145(.A(new_n19488), .B(new_n5054), .Y(new_n19494));
  nor_5  g17146(.A(new_n5060), .B(new_n5053), .Y(new_n19495));
  and_6  g17147(.A(new_n19495), .B(new_n19490), .Y(new_n19496));
  nor_5  g17148(.A(new_n19496), .B(new_n19494), .Y(new_n19497));
  nand_5 g17149(.A(new_n19497), .B(new_n19493), .Y(new_n19498));
  and_6  g17150(.A(new_n19498), .B(new_n19487), .Y(new_n19499));
  nor_5  g17151(.A(new_n19499), .B(new_n19486), .Y(new_n19500));
  nand_5 g17152(.A(new_n19500), .B(new_n19484), .Y(new_n19501));
  nand_5 g17153(.A(new_n19501), .B(new_n19483), .Y(new_n19502));
  xor_4  g17154(.A(new_n19480), .B(new_n3290), .Y(new_n19503));
  nand_5 g17155(.A(new_n19503), .B(new_n19502), .Y(new_n19504));
  nand_5 g17156(.A(new_n19504), .B(new_n19481), .Y(new_n19505));
  nor_5  g17157(.A(new_n19505), .B(new_n19479), .Y(new_n19506));
  or_6   g17158(.A(new_n19506), .B(new_n19478), .Y(new_n19507));
  xor_4  g17159(.A(new_n19475), .B(new_n19474), .Y(new_n19508));
  nand_5 g17160(.A(new_n19508), .B(new_n19507), .Y(new_n19509));
  nand_5 g17161(.A(new_n19509), .B(new_n19476), .Y(new_n19510));
  xor_4  g17162(.A(new_n19472), .B(new_n3263), .Y(new_n19511));
  nand_5 g17163(.A(new_n19511), .B(new_n19510), .Y(new_n19512));
  nand_5 g17164(.A(new_n19512), .B(new_n19473), .Y(new_n19513));
  not_8  g17165(.A(new_n16192), .Y(new_n19514));
  nor_5  g17166(.A(new_n19471), .B(new_n19514), .Y(new_n19515));
  not_8  g17167(.A(pi485), .Y(new_n19516));
  nor_5  g17168(.A(new_n16189), .B(new_n19516), .Y(new_n19517));
  nor_5  g17169(.A(new_n19517), .B(new_n19515), .Y(new_n19518));
  xor_4  g17170(.A(new_n19518), .B(new_n16205), .Y(new_n19519));
  xor_4  g17171(.A(new_n19519), .B(new_n3309), .Y(new_n19520));
  xnor_4 g17172(.A(new_n19520), .B(new_n19513), .Y(po0301));
  xor_4  g17173(.A(new_n11342), .B(new_n11317), .Y(po0302));
  nand_5 g17174(.A(new_n14272), .B(pi121), .Y(new_n19523));
  xor_4  g17175(.A(new_n14272), .B(pi121), .Y(new_n19524));
  not_8  g17176(.A(new_n14282), .Y(new_n19525));
  nand_5 g17177(.A(new_n19525), .B(pi162), .Y(new_n19526));
  xor_4  g17178(.A(new_n14282), .B(new_n6005), .Y(new_n19527));
  nand_5 g17179(.A(new_n9561), .B(pi352), .Y(new_n19528));
  nand_5 g17180(.A(new_n19528), .B(new_n9562), .Y(new_n19529));
  nand_5 g17181(.A(new_n19529), .B(new_n19527), .Y(new_n19530));
  nand_5 g17182(.A(new_n19530), .B(new_n19526), .Y(new_n19531));
  nand_5 g17183(.A(new_n19531), .B(new_n14279), .Y(new_n19532));
  xor_4  g17184(.A(new_n19531), .B(new_n14277), .Y(new_n19533));
  or_6   g17185(.A(new_n19533), .B(new_n7703), .Y(new_n19534));
  nand_5 g17186(.A(new_n19534), .B(new_n19532), .Y(new_n19535));
  nand_5 g17187(.A(new_n19535), .B(new_n19524), .Y(new_n19536));
  nand_5 g17188(.A(new_n19536), .B(new_n19523), .Y(new_n19537));
  nand_5 g17189(.A(new_n19537), .B(new_n14270), .Y(new_n19538));
  not_8  g17190(.A(new_n19538), .Y(new_n19539));
  nand_5 g17191(.A(new_n9547), .B(pi724), .Y(new_n19540));
  nand_5 g17192(.A(new_n19540), .B(new_n9546), .Y(new_n19541));
  and_6  g17193(.A(new_n19541), .B(new_n10281), .Y(new_n19542));
  nor_5  g17194(.A(new_n19541), .B(new_n10281), .Y(new_n19543));
  nor_5  g17195(.A(new_n19543), .B(new_n2898), .Y(new_n19544));
  nor_5  g17196(.A(new_n19544), .B(new_n19542), .Y(new_n19545));
  nand_5 g17197(.A(new_n19545), .B(new_n10319), .Y(new_n19546));
  xor_4  g17198(.A(new_n19545), .B(new_n10319), .Y(new_n19547));
  nand_5 g17199(.A(new_n19547), .B(new_n9154), .Y(new_n19548));
  nand_5 g17200(.A(new_n19548), .B(new_n19546), .Y(new_n19549));
  or_6   g17201(.A(new_n19549), .B(new_n10278), .Y(new_n19550));
  xor_4  g17202(.A(new_n19549), .B(new_n10278), .Y(new_n19551));
  nand_5 g17203(.A(new_n19551), .B(pi512), .Y(new_n19552));
  nand_5 g17204(.A(new_n19552), .B(new_n19550), .Y(new_n19553));
  nand_5 g17205(.A(new_n19553), .B(new_n10404), .Y(new_n19554));
  xor_4  g17206(.A(new_n19554), .B(new_n19539), .Y(new_n19555));
  not_8  g17207(.A(new_n19555), .Y(new_n19556));
  nor_5  g17208(.A(new_n19537), .B(new_n14270), .Y(new_n19557));
  nor_5  g17209(.A(new_n19557), .B(new_n19539), .Y(new_n19558));
  xor_4  g17210(.A(new_n19553), .B(new_n10403), .Y(new_n19559));
  nand_5 g17211(.A(new_n19559), .B(new_n19558), .Y(new_n19560));
  xor_4  g17212(.A(new_n19533), .B(new_n7703), .Y(new_n19561));
  not_8  g17213(.A(new_n19561), .Y(new_n19562));
  xor_4  g17214(.A(new_n19547), .B(pi224), .Y(new_n19563));
  nor_5  g17215(.A(new_n19563), .B(new_n19562), .Y(new_n19564));
  xor_4  g17216(.A(new_n19563), .B(new_n19562), .Y(new_n19565));
  not_8  g17217(.A(new_n19565), .Y(new_n19566));
  xor_4  g17218(.A(new_n19529), .B(new_n19527), .Y(new_n19567));
  nor_5  g17219(.A(new_n19543), .B(new_n19542), .Y(new_n19568));
  xor_4  g17220(.A(new_n19568), .B(new_n2898), .Y(new_n19569));
  or_6   g17221(.A(new_n19569), .B(new_n19567), .Y(new_n19570));
  not_8  g17222(.A(new_n9564), .Y(new_n19571));
  nor_5  g17223(.A(new_n19571), .B(new_n9549), .Y(new_n19572));
  nor_5  g17224(.A(new_n9565), .B(new_n9537), .Y(new_n19573));
  or_6   g17225(.A(new_n19573), .B(new_n19572), .Y(new_n19574));
  xor_4  g17226(.A(new_n19569), .B(new_n19567), .Y(new_n19575));
  nand_5 g17227(.A(new_n19575), .B(new_n19574), .Y(new_n19576));
  nand_5 g17228(.A(new_n19576), .B(new_n19570), .Y(new_n19577));
  nor_5  g17229(.A(new_n19577), .B(new_n19566), .Y(new_n19578));
  or_6   g17230(.A(new_n19578), .B(new_n19564), .Y(new_n19579));
  xor_4  g17231(.A(new_n19551), .B(new_n9169), .Y(new_n19580));
  nand_5 g17232(.A(new_n19580), .B(new_n19579), .Y(new_n19581));
  xor_4  g17233(.A(new_n19535), .B(new_n19524), .Y(new_n19582));
  xor_4  g17234(.A(new_n19580), .B(new_n19579), .Y(new_n19583));
  nand_5 g17235(.A(new_n19583), .B(new_n19582), .Y(new_n19584));
  nand_5 g17236(.A(new_n19584), .B(new_n19581), .Y(new_n19585));
  xor_4  g17237(.A(new_n19559), .B(new_n19558), .Y(new_n19586));
  nand_5 g17238(.A(new_n19586), .B(new_n19585), .Y(new_n19587));
  nand_5 g17239(.A(new_n19587), .B(new_n19560), .Y(new_n19588));
  xor_4  g17240(.A(new_n19588), .B(new_n19556), .Y(po0303));
  xor_4  g17241(.A(new_n19211), .B(new_n15196), .Y(po0304));
  nand_5 g17242(.A(new_n16883), .B(new_n16870), .Y(new_n19591));
  or_6   g17243(.A(new_n16884), .B(new_n8222), .Y(new_n19592));
  nand_5 g17244(.A(new_n19592), .B(new_n19591), .Y(new_n19593));
  xor_4  g17245(.A(new_n19593), .B(new_n8283), .Y(new_n19594));
  not_8  g17246(.A(new_n19594), .Y(new_n19595));
  xor_4  g17247(.A(pi534), .B(new_n8981), .Y(new_n19596));
  nand_5 g17248(.A(pi469), .B(new_n7257), .Y(new_n19597));
  not_8  g17249(.A(new_n19597), .Y(new_n19598));
  not_8  g17250(.A(new_n16871), .Y(new_n19599));
  nor_5  g17251(.A(new_n16876), .B(new_n19599), .Y(new_n19600));
  nor_5  g17252(.A(new_n19600), .B(new_n19598), .Y(new_n19601));
  xor_4  g17253(.A(new_n19601), .B(new_n19596), .Y(new_n19602));
  not_8  g17254(.A(new_n19602), .Y(new_n19603));
  nand_5 g17255(.A(new_n16881), .B(pi827), .Y(new_n19604));
  nand_5 g17256(.A(new_n19604), .B(new_n16880), .Y(new_n19605));
  nand_5 g17257(.A(new_n19605), .B(new_n19603), .Y(new_n19606));
  or_6   g17258(.A(new_n19605), .B(new_n19603), .Y(new_n19607));
  nand_5 g17259(.A(new_n19607), .B(new_n19606), .Y(new_n19608));
  xor_4  g17260(.A(new_n19608), .B(pi405), .Y(new_n19609));
  xor_4  g17261(.A(new_n19609), .B(new_n19595), .Y(po0305));
  not_8  g17262(.A(new_n4527), .Y(new_n19611));
  nand_5 g17263(.A(new_n15546), .B(pi141), .Y(new_n19612));
  nor_5  g17264(.A(new_n9253), .B(pi542), .Y(new_n19613));
  nand_5 g17265(.A(new_n19613), .B(new_n19612), .Y(new_n19614));
  or_6   g17266(.A(new_n19614), .B(new_n9308), .Y(new_n19615));
  nor_5  g17267(.A(new_n9308), .B(new_n9255), .Y(new_n19616));
  nor_5  g17268(.A(new_n19616), .B(new_n19613), .Y(new_n19617));
  or_6   g17269(.A(new_n9254), .B(new_n9209), .Y(new_n19618));
  nand_5 g17270(.A(new_n19618), .B(new_n19612), .Y(new_n19619));
  xor_4  g17271(.A(new_n19619), .B(new_n19617), .Y(new_n19620));
  nand_5 g17272(.A(new_n19620), .B(new_n19615), .Y(new_n19621));
  nor_5  g17273(.A(new_n19621), .B(new_n19611), .Y(new_n19622));
  xor_4  g17274(.A(new_n19621), .B(new_n19611), .Y(new_n19623));
  or_6   g17275(.A(new_n9309), .B(new_n4432), .Y(new_n19624));
  nand_5 g17276(.A(new_n9373), .B(new_n9310), .Y(new_n19625));
  nand_5 g17277(.A(new_n19625), .B(new_n19624), .Y(new_n19626));
  nand_5 g17278(.A(new_n19626), .B(new_n19623), .Y(new_n19627));
  not_8  g17279(.A(new_n19627), .Y(new_n19628));
  nor_5  g17280(.A(new_n19628), .B(new_n19622), .Y(new_n19629));
  nor_5  g17281(.A(new_n19621), .B(new_n18173), .Y(new_n19630));
  nand_5 g17282(.A(new_n19630), .B(new_n4522), .Y(new_n19631));
  and_6  g17283(.A(new_n19631), .B(new_n19629), .Y(new_n19632));
  nor_5  g17284(.A(new_n19630), .B(new_n4522), .Y(new_n19633));
  nor_5  g17285(.A(new_n19633), .B(new_n19629), .Y(new_n19634));
  nor_5  g17286(.A(new_n19634), .B(new_n19632), .Y(po0306));
  xor_4  g17287(.A(pi671), .B(pi555), .Y(new_n19636));
  nand_5 g17288(.A(new_n8641), .B(new_n6957), .Y(new_n19637));
  nand_5 g17289(.A(new_n6960), .B(new_n13485), .Y(new_n19638));
  not_8  g17290(.A(new_n19333), .Y(new_n19639));
  nand_5 g17291(.A(new_n19335), .B(new_n19639), .Y(new_n19640));
  nand_5 g17292(.A(new_n19640), .B(new_n19638), .Y(new_n19641));
  not_8  g17293(.A(new_n19641), .Y(new_n19642));
  xor_4  g17294(.A(pi768), .B(new_n6957), .Y(new_n19643));
  or_6   g17295(.A(new_n19643), .B(new_n19642), .Y(new_n19644));
  nand_5 g17296(.A(new_n19644), .B(new_n19637), .Y(new_n19645));
  xor_4  g17297(.A(new_n19645), .B(new_n19636), .Y(new_n19646));
  not_8  g17298(.A(new_n19646), .Y(new_n19647));
  xor_4  g17299(.A(new_n19647), .B(new_n7564), .Y(new_n19648));
  xor_4  g17300(.A(new_n19643), .B(new_n19641), .Y(new_n19649));
  nor_5  g17301(.A(new_n19649), .B(new_n2380), .Y(new_n19650));
  xor_4  g17302(.A(new_n19649), .B(new_n2380), .Y(new_n19651));
  nor_5  g17303(.A(new_n19336), .B(new_n2462), .Y(new_n19652));
  nor_5  g17304(.A(new_n19337), .B(new_n19332), .Y(new_n19653));
  or_6   g17305(.A(new_n19653), .B(new_n19652), .Y(new_n19654));
  and_6  g17306(.A(new_n19654), .B(new_n19651), .Y(new_n19655));
  nor_5  g17307(.A(new_n19655), .B(new_n19650), .Y(new_n19656));
  xor_4  g17308(.A(new_n19656), .B(new_n19648), .Y(new_n19657));
  xor_4  g17309(.A(pi527), .B(new_n2897), .Y(new_n19658));
  nand_5 g17310(.A(pi816), .B(new_n2932), .Y(new_n19659));
  xor_4  g17311(.A(pi816), .B(new_n2932), .Y(new_n19660));
  nand_5 g17312(.A(new_n19343), .B(new_n19341), .Y(new_n19661));
  nand_5 g17313(.A(new_n19661), .B(new_n19342), .Y(new_n19662));
  nand_5 g17314(.A(new_n19662), .B(new_n19660), .Y(new_n19663));
  nand_5 g17315(.A(new_n19663), .B(new_n19659), .Y(new_n19664));
  xor_4  g17316(.A(new_n19664), .B(new_n19658), .Y(new_n19665));
  xor_4  g17317(.A(new_n19665), .B(new_n19657), .Y(new_n19666));
  xor_4  g17318(.A(new_n19654), .B(new_n19651), .Y(new_n19667));
  not_8  g17319(.A(new_n19667), .Y(new_n19668));
  xnor_4 g17320(.A(new_n19662), .B(new_n19660), .Y(new_n19669));
  nor_5  g17321(.A(new_n19669), .B(new_n19668), .Y(new_n19670));
  xor_4  g17322(.A(new_n19669), .B(new_n19667), .Y(new_n19671));
  or_6   g17323(.A(new_n19345), .B(new_n19338), .Y(new_n19672));
  nand_5 g17324(.A(new_n19346), .B(new_n19329), .Y(new_n19673));
  nand_5 g17325(.A(new_n19673), .B(new_n19672), .Y(new_n19674));
  nor_5  g17326(.A(new_n19674), .B(new_n19671), .Y(new_n19675));
  nor_5  g17327(.A(new_n19675), .B(new_n19670), .Y(new_n19676));
  xnor_4 g17328(.A(new_n19676), .B(new_n19666), .Y(po0307));
  xor_4  g17329(.A(new_n19413), .B(new_n19408), .Y(po0308));
  xor_4  g17330(.A(new_n19425), .B(new_n19403), .Y(po0309));
  xor_4  g17331(.A(pi705), .B(new_n8055), .Y(new_n19680));
  nand_5 g17332(.A(pi798), .B(new_n8762), .Y(new_n19681));
  nand_5 g17333(.A(new_n18277), .B(new_n18275), .Y(new_n19682));
  nand_5 g17334(.A(new_n19682), .B(new_n18276), .Y(new_n19683));
  nand_5 g17335(.A(new_n19683), .B(new_n10037), .Y(new_n19684));
  nand_5 g17336(.A(new_n19684), .B(new_n19681), .Y(new_n19685));
  xor_4  g17337(.A(new_n19685), .B(new_n19680), .Y(new_n19686));
  or_6   g17338(.A(new_n19686), .B(new_n15418), .Y(new_n19687));
  xor_4  g17339(.A(new_n19686), .B(new_n15418), .Y(new_n19688));
  xor_4  g17340(.A(new_n19683), .B(new_n10037), .Y(new_n19689));
  or_6   g17341(.A(new_n19689), .B(new_n15348), .Y(new_n19690));
  xor_4  g17342(.A(new_n19689), .B(new_n15348), .Y(new_n19691));
  nor_5  g17343(.A(new_n18279), .B(new_n15687), .Y(new_n19692));
  not_8  g17344(.A(new_n18280), .Y(new_n19693));
  nor_5  g17345(.A(new_n18283), .B(new_n19693), .Y(new_n19694));
  nor_5  g17346(.A(new_n19694), .B(new_n19692), .Y(new_n19695));
  nand_5 g17347(.A(new_n19695), .B(new_n19691), .Y(new_n19696));
  nand_5 g17348(.A(new_n19696), .B(new_n19690), .Y(new_n19697));
  nand_5 g17349(.A(new_n19697), .B(new_n19688), .Y(new_n19698));
  nand_5 g17350(.A(new_n19698), .B(new_n19687), .Y(new_n19699));
  nand_5 g17351(.A(pi705), .B(new_n8055), .Y(new_n19700));
  nand_5 g17352(.A(new_n19685), .B(new_n19680), .Y(new_n19701));
  nand_5 g17353(.A(new_n19701), .B(new_n19700), .Y(new_n19702));
  xor_4  g17354(.A(new_n19702), .B(new_n10095), .Y(new_n19703));
  xor_4  g17355(.A(new_n19703), .B(new_n15685), .Y(new_n19704));
  xor_4  g17356(.A(new_n19704), .B(new_n19699), .Y(new_n19705));
  not_8  g17357(.A(new_n10112), .Y(new_n19706));
  nor_5  g17358(.A(new_n15425), .B(new_n10083), .Y(new_n19707));
  nor_5  g17359(.A(new_n19707), .B(new_n10081), .Y(new_n19708));
  xor_4  g17360(.A(new_n19708), .B(new_n19706), .Y(new_n19709));
  xor_4  g17361(.A(new_n19709), .B(new_n19705), .Y(new_n19710));
  xor_4  g17362(.A(new_n19697), .B(new_n19688), .Y(new_n19711));
  not_8  g17363(.A(new_n19711), .Y(new_n19712));
  xor_4  g17364(.A(new_n19695), .B(new_n19691), .Y(new_n19713));
  not_8  g17365(.A(new_n19713), .Y(new_n19714));
  nor_5  g17366(.A(new_n18284), .B(new_n18272), .Y(new_n19715));
  nor_5  g17367(.A(new_n18286), .B(new_n15356), .Y(new_n19716));
  or_6   g17368(.A(new_n19716), .B(new_n19715), .Y(new_n19717));
  nand_5 g17369(.A(new_n19717), .B(new_n19714), .Y(new_n19718));
  xor_4  g17370(.A(new_n19717), .B(new_n19713), .Y(new_n19719));
  or_6   g17371(.A(new_n19719), .B(new_n15372), .Y(new_n19720));
  nand_5 g17372(.A(new_n19720), .B(new_n19718), .Y(new_n19721));
  or_6   g17373(.A(new_n19721), .B(new_n19712), .Y(new_n19722));
  nand_5 g17374(.A(new_n19721), .B(new_n19712), .Y(new_n19723));
  nand_5 g17375(.A(new_n19723), .B(new_n15427), .Y(new_n19724));
  nand_5 g17376(.A(new_n19724), .B(new_n19722), .Y(new_n19725));
  xor_4  g17377(.A(new_n19725), .B(new_n19710), .Y(po0310));
  xor_4  g17378(.A(pi462), .B(new_n9217), .Y(new_n19727));
  nand_5 g17379(.A(new_n9220), .B(pi099), .Y(new_n19728));
  xor_4  g17380(.A(pi363), .B(new_n9322), .Y(new_n19729));
  nand_5 g17381(.A(new_n9223), .B(pi083), .Y(new_n19730));
  xor_4  g17382(.A(pi104), .B(new_n9285), .Y(new_n19731));
  nand_5 g17383(.A(new_n9226), .B(pi087), .Y(new_n19732));
  not_8  g17384(.A(new_n14247), .Y(new_n19733));
  nand_5 g17385(.A(new_n19733), .B(new_n14246), .Y(new_n19734));
  nand_5 g17386(.A(new_n19734), .B(new_n19732), .Y(new_n19735));
  nand_5 g17387(.A(new_n19735), .B(new_n19731), .Y(new_n19736));
  nand_5 g17388(.A(new_n19736), .B(new_n19730), .Y(new_n19737));
  nand_5 g17389(.A(new_n19737), .B(new_n19729), .Y(new_n19738));
  nand_5 g17390(.A(new_n19738), .B(new_n19728), .Y(new_n19739));
  xor_4  g17391(.A(new_n19739), .B(new_n19727), .Y(new_n19740));
  xnor_4 g17392(.A(new_n19737), .B(new_n19729), .Y(new_n19741));
  not_8  g17393(.A(new_n9099), .Y(new_n19742));
  not_8  g17394(.A(new_n14243), .Y(new_n19743));
  nand_5 g17395(.A(new_n14248), .B(new_n19743), .Y(new_n19744));
  nand_5 g17396(.A(new_n14250), .B(new_n9123), .Y(new_n19745));
  nand_5 g17397(.A(new_n19745), .B(new_n19744), .Y(new_n19746));
  nand_5 g17398(.A(new_n19746), .B(new_n19742), .Y(new_n19747));
  xnor_4 g17399(.A(new_n19735), .B(new_n19731), .Y(new_n19748));
  xor_4  g17400(.A(new_n19746), .B(new_n9099), .Y(new_n19749));
  not_8  g17401(.A(new_n19749), .Y(new_n19750));
  nand_5 g17402(.A(new_n19750), .B(new_n19748), .Y(new_n19751));
  nand_5 g17403(.A(new_n19751), .B(new_n19747), .Y(new_n19752));
  nand_5 g17404(.A(new_n19752), .B(new_n19741), .Y(new_n19753));
  xor_4  g17405(.A(new_n19752), .B(new_n19741), .Y(new_n19754));
  nand_5 g17406(.A(new_n19754), .B(new_n9132), .Y(new_n19755));
  nand_5 g17407(.A(new_n19755), .B(new_n19753), .Y(new_n19756));
  xor_4  g17408(.A(new_n19756), .B(new_n19740), .Y(new_n19757));
  xor_4  g17409(.A(new_n19757), .B(new_n9137), .Y(po0311));
  xor_4  g17410(.A(pi609), .B(new_n6434), .Y(new_n19759));
  nand_5 g17411(.A(pi640), .B(new_n4086), .Y(new_n19760));
  not_8  g17412(.A(new_n15627), .Y(new_n19761));
  xor_4  g17413(.A(pi640), .B(new_n4086), .Y(new_n19762));
  nand_5 g17414(.A(new_n19762), .B(new_n19761), .Y(new_n19763));
  nand_5 g17415(.A(new_n19763), .B(new_n19760), .Y(new_n19764));
  xor_4  g17416(.A(new_n19764), .B(new_n19759), .Y(new_n19765));
  xor_4  g17417(.A(new_n19765), .B(new_n18258), .Y(new_n19766));
  nor_5  g17418(.A(new_n15627), .B(new_n18243), .Y(new_n19767));
  nand_5 g17419(.A(new_n19762), .B(new_n18241), .Y(new_n19768));
  nor_5  g17420(.A(new_n19768), .B(new_n19767), .Y(new_n19769));
  or_6   g17421(.A(new_n15628), .B(new_n18243), .Y(new_n19770));
  nand_5 g17422(.A(new_n19761), .B(new_n18243), .Y(new_n19771));
  nand_5 g17423(.A(new_n19771), .B(new_n19770), .Y(new_n19772));
  xor_4  g17424(.A(new_n19762), .B(new_n18241), .Y(new_n19773));
  nor_5  g17425(.A(new_n19773), .B(new_n19772), .Y(new_n19774));
  nand_5 g17426(.A(new_n19770), .B(new_n19763), .Y(new_n19775));
  nor_5  g17427(.A(new_n19775), .B(new_n19774), .Y(new_n19776));
  nor_5  g17428(.A(new_n19776), .B(new_n19769), .Y(new_n19777));
  xor_4  g17429(.A(new_n19777), .B(new_n19766), .Y(po0312));
  xnor_4 g17430(.A(new_n14241), .B(new_n9116), .Y(po0313));
  xnor_4 g17431(.A(new_n18935), .B(new_n18910), .Y(po0314));
  nand_5 g17432(.A(new_n10356), .B(new_n10355), .Y(new_n19781));
  xnor_4 g17433(.A(new_n19781), .B(new_n10372), .Y(po0315));
  nand_5 g17434(.A(new_n17484), .B(pi512), .Y(new_n19783));
  nand_5 g17435(.A(pi663), .B(new_n9169), .Y(new_n19784));
  nand_5 g17436(.A(new_n19784), .B(new_n19783), .Y(new_n19785));
  nand_5 g17437(.A(new_n4335), .B(pi224), .Y(new_n19786));
  nand_5 g17438(.A(new_n19448), .B(new_n19445), .Y(new_n19787));
  nand_5 g17439(.A(new_n19787), .B(new_n19786), .Y(new_n19788));
  xnor_4 g17440(.A(new_n19788), .B(new_n19785), .Y(new_n19789));
  not_8  g17441(.A(new_n19789), .Y(new_n19790));
  xor_4  g17442(.A(new_n19790), .B(new_n10324), .Y(new_n19791));
  or_6   g17443(.A(new_n19449), .B(new_n10329), .Y(new_n19792));
  nand_5 g17444(.A(new_n19450), .B(new_n19444), .Y(new_n19793));
  nand_5 g17445(.A(new_n19793), .B(new_n19792), .Y(new_n19794));
  xnor_4 g17446(.A(new_n19794), .B(new_n19791), .Y(po0316));
  xor_4  g17447(.A(new_n15059), .B(new_n16966), .Y(po0317));
  not_8  g17448(.A(pi722), .Y(new_n19797));
  nand_5 g17449(.A(new_n19797), .B(pi278), .Y(new_n19798));
  nand_5 g17450(.A(new_n19708), .B(new_n19706), .Y(new_n19799));
  nand_5 g17451(.A(new_n19799), .B(new_n19798), .Y(new_n19800));
  nand_5 g17452(.A(pi465), .B(new_n10165), .Y(new_n19801));
  nand_5 g17453(.A(new_n19801), .B(new_n19800), .Y(new_n19802));
  nand_5 g17454(.A(new_n10166), .B(pi431), .Y(new_n19803));
  nand_5 g17455(.A(new_n19803), .B(new_n19802), .Y(new_n19804));
  nand_5 g17456(.A(pi443), .B(new_n10405), .Y(new_n19805));
  xor_4  g17457(.A(pi443), .B(new_n10405), .Y(new_n19806));
  nand_5 g17458(.A(pi701), .B(new_n2837), .Y(new_n19807));
  nand_5 g17459(.A(new_n15129), .B(new_n15109), .Y(new_n19808));
  nand_5 g17460(.A(new_n19808), .B(new_n19807), .Y(new_n19809));
  nand_5 g17461(.A(new_n19809), .B(new_n19806), .Y(new_n19810));
  nand_5 g17462(.A(new_n19810), .B(new_n19805), .Y(new_n19811));
  xor_4  g17463(.A(new_n19811), .B(new_n19804), .Y(new_n19812));
  xor_4  g17464(.A(new_n19800), .B(new_n10169), .Y(new_n19813));
  xor_4  g17465(.A(new_n19809), .B(new_n19806), .Y(new_n19814));
  nand_5 g17466(.A(new_n19814), .B(new_n19813), .Y(new_n19815));
  not_8  g17467(.A(new_n19813), .Y(new_n19816));
  not_8  g17468(.A(new_n19814), .Y(new_n19817));
  nand_5 g17469(.A(new_n19817), .B(new_n19816), .Y(new_n19818));
  nand_5 g17470(.A(new_n19709), .B(new_n15130), .Y(new_n19819));
  xor_4  g17471(.A(new_n19709), .B(new_n15130), .Y(new_n19820));
  nor_5  g17472(.A(new_n15426), .B(new_n15131), .Y(new_n19821));
  nor_5  g17473(.A(new_n15428), .B(new_n15422), .Y(new_n19822));
  nor_5  g17474(.A(new_n19822), .B(new_n19821), .Y(new_n19823));
  nand_5 g17475(.A(new_n19823), .B(new_n19820), .Y(new_n19824));
  nand_5 g17476(.A(new_n19824), .B(new_n19819), .Y(new_n19825));
  nand_5 g17477(.A(new_n19825), .B(new_n19818), .Y(new_n19826));
  nand_5 g17478(.A(new_n19826), .B(new_n19815), .Y(new_n19827));
  xor_4  g17479(.A(new_n19827), .B(new_n19812), .Y(new_n19828));
  nand_5 g17480(.A(new_n13053), .B(pi057), .Y(new_n19829));
  nand_5 g17481(.A(new_n10966), .B(pi193), .Y(new_n19830));
  nand_5 g17482(.A(new_n19188), .B(new_n19185), .Y(new_n19831));
  nand_5 g17483(.A(new_n19831), .B(new_n19830), .Y(new_n19832));
  nand_5 g17484(.A(pi292), .B(new_n17704), .Y(new_n19833));
  nand_5 g17485(.A(new_n19833), .B(new_n19829), .Y(new_n19834));
  not_8  g17486(.A(new_n19834), .Y(new_n19835));
  nand_5 g17487(.A(new_n19835), .B(new_n19832), .Y(new_n19836));
  nand_5 g17488(.A(new_n19836), .B(new_n19829), .Y(new_n19837));
  nand_5 g17489(.A(new_n19818), .B(new_n19815), .Y(new_n19838));
  xor_4  g17490(.A(new_n19838), .B(new_n19825), .Y(new_n19839));
  not_8  g17491(.A(new_n19839), .Y(new_n19840));
  xnor_4 g17492(.A(new_n19823), .B(new_n19820), .Y(new_n19841));
  nor_5  g17493(.A(new_n19841), .B(new_n19190), .Y(new_n19842));
  and_6  g17494(.A(new_n15598), .B(new_n15429), .Y(new_n19843));
  nor_5  g17495(.A(new_n15618), .B(new_n15600), .Y(new_n19844));
  nor_5  g17496(.A(new_n19844), .B(new_n19843), .Y(new_n19845));
  xor_4  g17497(.A(new_n19841), .B(new_n19189), .Y(new_n19846));
  nor_5  g17498(.A(new_n19846), .B(new_n19845), .Y(new_n19847));
  nor_5  g17499(.A(new_n19847), .B(new_n19842), .Y(new_n19848));
  not_8  g17500(.A(new_n19848), .Y(new_n19849));
  nand_5 g17501(.A(new_n19849), .B(new_n19840), .Y(new_n19850));
  and_6  g17502(.A(new_n19850), .B(new_n19837), .Y(new_n19851));
  not_8  g17503(.A(new_n19832), .Y(new_n19852));
  nor_5  g17504(.A(new_n19852), .B(new_n19829), .Y(new_n19853));
  nand_5 g17505(.A(new_n19848), .B(new_n19839), .Y(new_n19854));
  nand_5 g17506(.A(new_n19854), .B(new_n19853), .Y(new_n19855));
  nand_5 g17507(.A(new_n19855), .B(new_n19851), .Y(new_n19856));
  nand_5 g17508(.A(new_n19856), .B(new_n19828), .Y(new_n19857));
  nor_5  g17509(.A(new_n19833), .B(new_n19832), .Y(new_n19858));
  nand_5 g17510(.A(new_n19858), .B(new_n19850), .Y(new_n19859));
  not_8  g17511(.A(new_n19837), .Y(new_n19860));
  and_6  g17512(.A(new_n19854), .B(new_n19860), .Y(new_n19861));
  nand_5 g17513(.A(new_n19861), .B(new_n19859), .Y(new_n19862));
  nand_5 g17514(.A(new_n19862), .B(new_n19857), .Y(new_n19863));
  nand_5 g17515(.A(new_n19811), .B(new_n19804), .Y(new_n19864));
  nand_5 g17516(.A(new_n19827), .B(new_n19812), .Y(new_n19865));
  nand_5 g17517(.A(new_n19865), .B(new_n19864), .Y(new_n19866));
  xor_4  g17518(.A(new_n19866), .B(new_n19837), .Y(new_n19867));
  xnor_4 g17519(.A(new_n19867), .B(new_n19863), .Y(po0318));
  xor_4  g17520(.A(new_n18879), .B(new_n18878), .Y(po0319));
  xnor_4 g17521(.A(new_n16979), .B(new_n16965), .Y(po0320));
  xor_4  g17522(.A(new_n16731), .B(new_n16714), .Y(po0321));
  nand_5 g17523(.A(new_n5936), .B(new_n4857), .Y(new_n19872));
  nand_5 g17524(.A(new_n19872), .B(new_n5937), .Y(new_n19873));
  nor_5  g17525(.A(new_n19873), .B(new_n13718), .Y(new_n19874));
  nand_5 g17526(.A(new_n19874), .B(new_n18034), .Y(new_n19875));
  nand_5 g17527(.A(new_n6101), .B(new_n6086), .Y(new_n19876));
  nand_5 g17528(.A(new_n6102), .B(new_n5939), .Y(new_n19877));
  nand_5 g17529(.A(new_n19877), .B(new_n19876), .Y(new_n19878));
  xor_4  g17530(.A(new_n19873), .B(new_n13719), .Y(new_n19879));
  not_8  g17531(.A(new_n19879), .Y(new_n19880));
  nand_5 g17532(.A(new_n19880), .B(new_n19878), .Y(new_n19881));
  xor_4  g17533(.A(new_n19879), .B(new_n19878), .Y(new_n19882));
  or_6   g17534(.A(new_n19882), .B(new_n18042), .Y(new_n19883));
  nand_5 g17535(.A(new_n19883), .B(new_n19881), .Y(new_n19884));
  xor_4  g17536(.A(new_n19874), .B(new_n18034), .Y(new_n19885));
  nand_5 g17537(.A(new_n19885), .B(new_n19884), .Y(new_n19886));
  nand_5 g17538(.A(new_n19886), .B(new_n19875), .Y(po0322));
  xor_4  g17539(.A(new_n8637), .B(new_n8636), .Y(po0323));
  xor_4  g17540(.A(new_n14157), .B(new_n14156), .Y(po0324));
  nand_5 g17541(.A(pi234), .B(new_n3327), .Y(new_n19890));
  not_8  g17542(.A(new_n19890), .Y(new_n19891));
  xor_4  g17543(.A(pi234), .B(new_n3327), .Y(new_n19892));
  not_8  g17544(.A(new_n19892), .Y(new_n19893));
  nand_5 g17545(.A(pi325), .B(new_n13221), .Y(new_n19894));
  nand_5 g17546(.A(new_n3262), .B(pi189), .Y(new_n19895));
  nand_5 g17547(.A(pi637), .B(new_n5272), .Y(new_n19896));
  xor_4  g17548(.A(pi637), .B(new_n5272), .Y(new_n19897));
  nand_5 g17549(.A(pi253), .B(new_n5275), .Y(new_n19898));
  nand_5 g17550(.A(new_n3333), .B(pi018), .Y(new_n19899));
  not_8  g17551(.A(pi217), .Y(new_n19900));
  nand_5 g17552(.A(pi829), .B(new_n19900), .Y(new_n19901));
  nor_5  g17553(.A(pi829), .B(new_n19900), .Y(new_n19902));
  not_8  g17554(.A(pi107), .Y(new_n19903));
  nand_5 g17555(.A(pi153), .B(new_n19903), .Y(new_n19904));
  not_8  g17556(.A(new_n19904), .Y(new_n19905));
  xor_4  g17557(.A(pi153), .B(new_n19903), .Y(new_n19906));
  not_8  g17558(.A(new_n19906), .Y(new_n19907));
  nand_5 g17559(.A(pi749), .B(new_n5283), .Y(new_n19908));
  not_8  g17560(.A(new_n19908), .Y(new_n19909));
  xor_4  g17561(.A(pi749), .B(new_n5283), .Y(new_n19910));
  not_8  g17562(.A(new_n19910), .Y(new_n19911));
  nand_5 g17563(.A(new_n2389), .B(pi076), .Y(new_n19912));
  nand_5 g17564(.A(pi755), .B(new_n5286), .Y(new_n19913));
  nand_5 g17565(.A(new_n5351), .B(new_n5343), .Y(new_n19914));
  nand_5 g17566(.A(new_n19914), .B(new_n5350), .Y(new_n19915));
  nand_5 g17567(.A(new_n19915), .B(new_n19913), .Y(new_n19916));
  nand_5 g17568(.A(new_n19916), .B(new_n19912), .Y(new_n19917));
  nor_5  g17569(.A(new_n19917), .B(new_n19911), .Y(new_n19918));
  nor_5  g17570(.A(new_n19918), .B(new_n19909), .Y(new_n19919));
  nor_5  g17571(.A(new_n19919), .B(new_n19907), .Y(new_n19920));
  nor_5  g17572(.A(new_n19920), .B(new_n19905), .Y(new_n19921));
  or_6   g17573(.A(new_n19921), .B(new_n19902), .Y(new_n19922));
  nand_5 g17574(.A(new_n19922), .B(new_n19901), .Y(new_n19923));
  nand_5 g17575(.A(new_n19923), .B(new_n19899), .Y(new_n19924));
  nand_5 g17576(.A(new_n19924), .B(new_n19898), .Y(new_n19925));
  nand_5 g17577(.A(new_n19925), .B(new_n19897), .Y(new_n19926));
  nand_5 g17578(.A(new_n19926), .B(new_n19896), .Y(new_n19927));
  nand_5 g17579(.A(new_n19927), .B(new_n19895), .Y(new_n19928));
  nand_5 g17580(.A(new_n19928), .B(new_n19894), .Y(new_n19929));
  nor_5  g17581(.A(new_n19929), .B(new_n19893), .Y(new_n19930));
  nor_5  g17582(.A(new_n19930), .B(new_n19891), .Y(new_n19931));
  or_6   g17583(.A(new_n19931), .B(new_n17171), .Y(new_n19932));
  xor_4  g17584(.A(new_n19931), .B(new_n17171), .Y(new_n19933));
  not_8  g17585(.A(new_n17212), .Y(new_n19934));
  nand_5 g17586(.A(new_n17257), .B(new_n5343), .Y(new_n19935));
  nand_5 g17587(.A(new_n17251), .B(new_n5344), .Y(new_n19936));
  nand_5 g17588(.A(new_n19936), .B(new_n19935), .Y(new_n19937));
  xor_4  g17589(.A(new_n19937), .B(new_n5352), .Y(new_n19938));
  or_6   g17590(.A(new_n19938), .B(new_n17247), .Y(new_n19939));
  nand_5 g17591(.A(new_n17251), .B(new_n5345), .Y(new_n19940));
  nand_5 g17592(.A(new_n19940), .B(new_n19938), .Y(new_n19941));
  nand_5 g17593(.A(new_n19941), .B(new_n19939), .Y(new_n19942));
  and_6  g17594(.A(new_n19913), .B(new_n19912), .Y(new_n19943));
  xor_4  g17595(.A(new_n19943), .B(new_n19915), .Y(new_n19944));
  not_8  g17596(.A(new_n19944), .Y(new_n19945));
  nand_5 g17597(.A(new_n19945), .B(new_n19942), .Y(new_n19946));
  xor_4  g17598(.A(new_n19944), .B(new_n19942), .Y(new_n19947));
  or_6   g17599(.A(new_n19947), .B(new_n17242), .Y(new_n19948));
  nand_5 g17600(.A(new_n19948), .B(new_n19946), .Y(new_n19949));
  xor_4  g17601(.A(new_n19917), .B(new_n19910), .Y(new_n19950));
  not_8  g17602(.A(new_n19950), .Y(new_n19951));
  nand_5 g17603(.A(new_n19951), .B(new_n19949), .Y(new_n19952));
  xor_4  g17604(.A(new_n19950), .B(new_n19949), .Y(new_n19953));
  or_6   g17605(.A(new_n19953), .B(new_n17237), .Y(new_n19954));
  nand_5 g17606(.A(new_n19954), .B(new_n19952), .Y(new_n19955));
  xor_4  g17607(.A(new_n19919), .B(new_n19906), .Y(new_n19956));
  not_8  g17608(.A(new_n19956), .Y(new_n19957));
  nand_5 g17609(.A(new_n19957), .B(new_n19955), .Y(new_n19958));
  xor_4  g17610(.A(new_n19956), .B(new_n19955), .Y(new_n19959));
  or_6   g17611(.A(new_n19959), .B(new_n17232), .Y(new_n19960));
  nand_5 g17612(.A(new_n19960), .B(new_n19958), .Y(new_n19961));
  xor_4  g17613(.A(pi829), .B(new_n19900), .Y(new_n19962));
  xor_4  g17614(.A(new_n19962), .B(new_n19921), .Y(new_n19963));
  not_8  g17615(.A(new_n19963), .Y(new_n19964));
  nand_5 g17616(.A(new_n19964), .B(new_n19961), .Y(new_n19965));
  xor_4  g17617(.A(new_n19963), .B(new_n19961), .Y(new_n19966));
  or_6   g17618(.A(new_n19966), .B(new_n17226), .Y(new_n19967));
  nand_5 g17619(.A(new_n19967), .B(new_n19965), .Y(new_n19968));
  nand_5 g17620(.A(new_n19899), .B(new_n19898), .Y(new_n19969));
  xnor_4 g17621(.A(new_n19969), .B(new_n19923), .Y(new_n19970));
  nand_5 g17622(.A(new_n19970), .B(new_n19968), .Y(new_n19971));
  not_8  g17623(.A(new_n17222), .Y(new_n19972));
  xnor_4 g17624(.A(new_n19970), .B(new_n19968), .Y(new_n19973));
  or_6   g17625(.A(new_n19973), .B(new_n19972), .Y(new_n19974));
  nand_5 g17626(.A(new_n19974), .B(new_n19971), .Y(new_n19975));
  xor_4  g17627(.A(new_n19925), .B(new_n19897), .Y(new_n19976));
  nand_5 g17628(.A(new_n19976), .B(new_n19975), .Y(new_n19977));
  xnor_4 g17629(.A(new_n19976), .B(new_n19975), .Y(new_n19978));
  or_6   g17630(.A(new_n19978), .B(new_n17217), .Y(new_n19979));
  nand_5 g17631(.A(new_n19979), .B(new_n19977), .Y(new_n19980));
  nand_5 g17632(.A(new_n19980), .B(new_n19934), .Y(new_n19981));
  xor_4  g17633(.A(new_n19980), .B(new_n17212), .Y(new_n19982));
  nand_5 g17634(.A(new_n19895), .B(new_n19894), .Y(new_n19983));
  xor_4  g17635(.A(new_n19983), .B(new_n19927), .Y(new_n19984));
  or_6   g17636(.A(new_n19984), .B(new_n19982), .Y(new_n19985));
  nand_5 g17637(.A(new_n19985), .B(new_n19981), .Y(new_n19986));
  nor_5  g17638(.A(new_n19986), .B(new_n17174), .Y(new_n19987));
  xor_4  g17639(.A(new_n19986), .B(new_n17174), .Y(new_n19988));
  xor_4  g17640(.A(new_n19929), .B(new_n19892), .Y(new_n19989));
  not_8  g17641(.A(new_n19989), .Y(new_n19990));
  nand_5 g17642(.A(new_n19990), .B(new_n19988), .Y(new_n19991));
  not_8  g17643(.A(new_n19991), .Y(new_n19992));
  nor_5  g17644(.A(new_n19992), .B(new_n19987), .Y(new_n19993));
  not_8  g17645(.A(new_n19993), .Y(new_n19994));
  nand_5 g17646(.A(new_n19994), .B(new_n19933), .Y(new_n19995));
  nand_5 g17647(.A(new_n19995), .B(new_n19932), .Y(new_n19996));
  not_8  g17648(.A(new_n19996), .Y(new_n19997));
  nand_5 g17649(.A(new_n19997), .B(new_n17289), .Y(new_n19998));
  not_8  g17650(.A(new_n19995), .Y(new_n19999));
  nand_5 g17651(.A(new_n19999), .B(new_n17173), .Y(new_n20000));
  nand_5 g17652(.A(new_n20000), .B(new_n19998), .Y(po0325));
  nor_5  g17653(.A(new_n19035), .B(new_n19034), .Y(new_n20002));
  xor_4  g17654(.A(new_n20002), .B(new_n4966), .Y(po0326));
  xnor_4 g17655(.A(new_n14611), .B(new_n14610), .Y(po0327));
  xor_4  g17656(.A(new_n16403), .B(new_n8619), .Y(po0328));
  xor_4  g17657(.A(new_n16565), .B(new_n10503), .Y(po0329));
  xor_4  g17658(.A(new_n4124), .B(new_n4123), .Y(po0330));
  xor_4  g17659(.A(new_n12391), .B(new_n8864), .Y(po0331));
  not_8  g17660(.A(new_n8445), .Y(new_n20009));
  nand_5 g17661(.A(new_n17529), .B(new_n17525), .Y(new_n20010));
  nand_5 g17662(.A(new_n20010), .B(new_n17524), .Y(new_n20011));
  xor_4  g17663(.A(new_n20011), .B(new_n20009), .Y(new_n20012));
  not_8  g17664(.A(new_n20012), .Y(new_n20013));
  not_8  g17665(.A(new_n17530), .Y(new_n20014));
  nor_5  g17666(.A(new_n20014), .B(new_n3702), .Y(new_n20015));
  xor_4  g17667(.A(new_n20014), .B(new_n3702), .Y(new_n20016));
  not_8  g17668(.A(new_n20016), .Y(new_n20017));
  or_6   g17669(.A(new_n14626), .B(new_n3576), .Y(new_n20018));
  nand_5 g17670(.A(new_n14630), .B(new_n14627), .Y(new_n20019));
  nand_5 g17671(.A(new_n20019), .B(new_n20018), .Y(new_n20020));
  nor_5  g17672(.A(new_n20020), .B(new_n20017), .Y(new_n20021));
  nor_5  g17673(.A(new_n20021), .B(new_n20015), .Y(new_n20022));
  nor_5  g17674(.A(new_n20022), .B(new_n20013), .Y(new_n20023));
  not_8  g17675(.A(new_n20023), .Y(new_n20024));
  nand_5 g17676(.A(new_n20022), .B(new_n20013), .Y(new_n20025));
  nand_5 g17677(.A(new_n20025), .B(new_n20024), .Y(new_n20026));
  not_8  g17678(.A(new_n20026), .Y(new_n20027));
  xor_4  g17679(.A(new_n20020), .B(new_n20017), .Y(new_n20028));
  nand_5 g17680(.A(pi650), .B(new_n3426), .Y(new_n20029));
  nand_5 g17681(.A(new_n14620), .B(new_n14617), .Y(new_n20030));
  nand_5 g17682(.A(new_n20030), .B(new_n20029), .Y(new_n20031));
  nand_5 g17683(.A(new_n3423), .B(pi089), .Y(new_n20032));
  nand_5 g17684(.A(pi303), .B(new_n3424), .Y(new_n20033));
  nand_5 g17685(.A(new_n20033), .B(new_n20032), .Y(new_n20034));
  xnor_4 g17686(.A(new_n20034), .B(new_n20031), .Y(new_n20035));
  nand_5 g17687(.A(new_n20035), .B(new_n20028), .Y(new_n20036));
  not_8  g17688(.A(new_n14621), .Y(new_n20037));
  nor_5  g17689(.A(new_n14631), .B(new_n20037), .Y(new_n20038));
  or_6   g17690(.A(new_n14632), .B(new_n14616), .Y(new_n20039));
  not_8  g17691(.A(new_n20039), .Y(new_n20040));
  nor_5  g17692(.A(new_n20040), .B(new_n20038), .Y(new_n20041));
  not_8  g17693(.A(new_n20028), .Y(new_n20042));
  xor_4  g17694(.A(new_n20035), .B(new_n20042), .Y(new_n20043));
  or_6   g17695(.A(new_n20043), .B(new_n20041), .Y(new_n20044));
  nand_5 g17696(.A(new_n20044), .B(new_n20036), .Y(new_n20045));
  xor_4  g17697(.A(new_n20045), .B(new_n20027), .Y(new_n20046));
  nand_5 g17698(.A(new_n20032), .B(new_n20031), .Y(new_n20047));
  nand_5 g17699(.A(new_n20047), .B(new_n20033), .Y(new_n20048));
  xor_4  g17700(.A(new_n20048), .B(new_n20046), .Y(po0332));
  xor_4  g17701(.A(new_n11627), .B(new_n11625), .Y(po0333));
  xor_4  g17702(.A(new_n18538), .B(new_n18537), .Y(po0334));
  xor_4  g17703(.A(new_n9557), .B(new_n9542), .Y(new_n20052));
  nor_5  g17704(.A(new_n9530), .B(new_n9516), .Y(new_n20053));
  xor_4  g17705(.A(new_n9530), .B(new_n9516), .Y(new_n20054));
  not_8  g17706(.A(new_n20054), .Y(new_n20055));
  or_6   g17707(.A(new_n9490), .B(new_n9480), .Y(new_n20056));
  nor_5  g17708(.A(new_n9493), .B(new_n9389), .Y(new_n20057));
  xor_4  g17709(.A(new_n9493), .B(new_n9389), .Y(new_n20058));
  not_8  g17710(.A(new_n20058), .Y(new_n20059));
  or_6   g17711(.A(new_n9427), .B(new_n9403), .Y(new_n20060));
  xor_4  g17712(.A(new_n9427), .B(new_n9403), .Y(new_n20061));
  not_8  g17713(.A(new_n9381), .Y(new_n20062));
  nand_5 g17714(.A(new_n9394), .B(new_n20062), .Y(new_n20063));
  not_8  g17715(.A(new_n20063), .Y(new_n20064));
  nand_5 g17716(.A(new_n9447), .B(new_n9395), .Y(new_n20065));
  nand_5 g17717(.A(new_n20065), .B(new_n9383), .Y(new_n20066));
  nor_5  g17718(.A(new_n20066), .B(new_n20064), .Y(new_n20067));
  nor_5  g17719(.A(new_n20065), .B(new_n20062), .Y(new_n20068));
  nor_5  g17720(.A(new_n20068), .B(new_n20067), .Y(new_n20069));
  nand_5 g17721(.A(new_n20069), .B(new_n9414), .Y(new_n20070));
  not_8  g17722(.A(new_n20070), .Y(new_n20071));
  nor_5  g17723(.A(new_n20071), .B(new_n20067), .Y(new_n20072));
  nand_5 g17724(.A(new_n20072), .B(new_n20061), .Y(new_n20073));
  nand_5 g17725(.A(new_n20073), .B(new_n20060), .Y(new_n20074));
  nor_5  g17726(.A(new_n20074), .B(new_n20059), .Y(new_n20075));
  or_6   g17727(.A(new_n20075), .B(new_n20057), .Y(new_n20076));
  xor_4  g17728(.A(new_n9491), .B(new_n9480), .Y(new_n20077));
  not_8  g17729(.A(new_n20077), .Y(new_n20078));
  nand_5 g17730(.A(new_n20078), .B(new_n20076), .Y(new_n20079));
  nand_5 g17731(.A(new_n20079), .B(new_n20056), .Y(new_n20080));
  nor_5  g17732(.A(new_n20080), .B(new_n20055), .Y(new_n20081));
  nor_5  g17733(.A(new_n20081), .B(new_n20053), .Y(new_n20082));
  xnor_4 g17734(.A(new_n20082), .B(new_n20052), .Y(new_n20083));
  or_6   g17735(.A(new_n20083), .B(new_n16821), .Y(new_n20084));
  xor_4  g17736(.A(new_n20083), .B(new_n16821), .Y(new_n20085));
  xor_4  g17737(.A(new_n9416), .B(new_n9396), .Y(new_n20086));
  nor_5  g17738(.A(new_n20086), .B(new_n16834), .Y(new_n20087));
  nor_5  g17739(.A(new_n20087), .B(new_n16799), .Y(new_n20088));
  xnor_4 g17740(.A(new_n20087), .B(new_n16799), .Y(new_n20089));
  xor_4  g17741(.A(new_n20069), .B(new_n9414), .Y(new_n20090));
  nor_5  g17742(.A(new_n20090), .B(new_n20089), .Y(new_n20091));
  or_6   g17743(.A(new_n20091), .B(new_n20088), .Y(new_n20092));
  or_6   g17744(.A(new_n20092), .B(new_n16802), .Y(new_n20093));
  xor_4  g17745(.A(new_n20092), .B(new_n16802), .Y(new_n20094));
  xnor_4 g17746(.A(new_n20072), .B(new_n20061), .Y(new_n20095));
  nand_5 g17747(.A(new_n20095), .B(new_n20094), .Y(new_n20096));
  nand_5 g17748(.A(new_n20096), .B(new_n20093), .Y(new_n20097));
  xor_4  g17749(.A(new_n20074), .B(new_n20059), .Y(new_n20098));
  nand_5 g17750(.A(new_n20098), .B(new_n20097), .Y(new_n20099));
  xor_4  g17751(.A(new_n20098), .B(new_n20097), .Y(new_n20100));
  nand_5 g17752(.A(new_n20100), .B(new_n16796), .Y(new_n20101));
  nand_5 g17753(.A(new_n20101), .B(new_n20099), .Y(new_n20102));
  xor_4  g17754(.A(new_n20077), .B(new_n20076), .Y(new_n20103));
  not_8  g17755(.A(new_n20103), .Y(new_n20104));
  nand_5 g17756(.A(new_n20104), .B(new_n20102), .Y(new_n20105));
  xor_4  g17757(.A(new_n20103), .B(new_n20102), .Y(new_n20106));
  or_6   g17758(.A(new_n20106), .B(new_n16795), .Y(new_n20107));
  nand_5 g17759(.A(new_n20107), .B(new_n20105), .Y(new_n20108));
  xor_4  g17760(.A(new_n20080), .B(new_n20054), .Y(new_n20109));
  nor_5  g17761(.A(new_n20109), .B(new_n20108), .Y(new_n20110));
  xnor_4 g17762(.A(new_n20109), .B(new_n20108), .Y(new_n20111));
  nor_5  g17763(.A(new_n20111), .B(new_n16816), .Y(new_n20112));
  nor_5  g17764(.A(new_n20112), .B(new_n20110), .Y(new_n20113));
  nand_5 g17765(.A(new_n20113), .B(new_n20085), .Y(new_n20114));
  nand_5 g17766(.A(new_n20114), .B(new_n20084), .Y(new_n20115));
  nor_5  g17767(.A(new_n20115), .B(new_n16791), .Y(new_n20116));
  xor_4  g17768(.A(new_n20115), .B(new_n16790), .Y(new_n20117));
  nand_5 g17769(.A(new_n9558), .B(new_n10311), .Y(new_n20118));
  nand_5 g17770(.A(new_n20082), .B(new_n20052), .Y(new_n20119));
  nand_5 g17771(.A(new_n20119), .B(new_n20118), .Y(new_n20120));
  xor_4  g17772(.A(new_n19525), .B(new_n10280), .Y(new_n20121));
  xor_4  g17773(.A(new_n20121), .B(new_n20120), .Y(new_n20122));
  nor_5  g17774(.A(new_n20122), .B(new_n20117), .Y(new_n20123));
  or_6   g17775(.A(new_n20123), .B(new_n20116), .Y(new_n20124));
  xnor_4 g17776(.A(new_n20124), .B(new_n16877), .Y(new_n20125));
  nand_5 g17777(.A(new_n14282), .B(new_n10281), .Y(new_n20126));
  nand_5 g17778(.A(new_n20121), .B(new_n20120), .Y(new_n20127));
  nand_5 g17779(.A(new_n20127), .B(new_n20126), .Y(new_n20128));
  xor_4  g17780(.A(new_n14277), .B(new_n10319), .Y(new_n20129));
  not_8  g17781(.A(new_n20129), .Y(new_n20130));
  xor_4  g17782(.A(new_n20130), .B(new_n20128), .Y(new_n20131));
  xnor_4 g17783(.A(new_n20131), .B(new_n20125), .Y(po0335));
  not_8  g17784(.A(new_n11597), .Y(new_n20133));
  nand_5 g17785(.A(new_n20133), .B(new_n11559), .Y(new_n20134));
  not_8  g17786(.A(new_n20134), .Y(new_n20135));
  nor_5  g17787(.A(new_n20133), .B(new_n11558), .Y(new_n20136));
  nor_5  g17788(.A(new_n20136), .B(new_n20135), .Y(new_n20137));
  nor_5  g17789(.A(new_n11598), .B(new_n11524), .Y(new_n20138));
  nor_5  g17790(.A(new_n11638), .B(new_n11600), .Y(new_n20139));
  nor_5  g17791(.A(new_n20139), .B(new_n20138), .Y(new_n20140));
  xnor_4 g17792(.A(new_n20140), .B(new_n20137), .Y(po0336));
  xnor_4 g17793(.A(new_n15469), .B(new_n15468), .Y(po0337));
  xor_4  g17794(.A(new_n18015), .B(new_n3087), .Y(po0338));
  nand_5 g17795(.A(new_n6133), .B(pi528), .Y(new_n20144));
  xor_4  g17796(.A(new_n6133), .B(new_n3954), .Y(new_n20145));
  not_8  g17797(.A(new_n20145), .Y(new_n20146));
  nand_5 g17798(.A(new_n20146), .B(new_n6137), .Y(new_n20147));
  nand_5 g17799(.A(new_n20147), .B(new_n20144), .Y(new_n20148));
  or_6   g17800(.A(new_n20148), .B(new_n6132), .Y(new_n20149));
  xor_4  g17801(.A(new_n20148), .B(new_n6132), .Y(new_n20150));
  nand_5 g17802(.A(new_n20150), .B(new_n3946), .Y(new_n20151));
  nand_5 g17803(.A(new_n20151), .B(new_n20149), .Y(new_n20152));
  xor_4  g17804(.A(new_n20152), .B(new_n6158), .Y(new_n20153));
  xor_4  g17805(.A(new_n20153), .B(pi338), .Y(new_n20154));
  xor_4  g17806(.A(new_n20150), .B(pi362), .Y(new_n20155));
  nor_5  g17807(.A(new_n20155), .B(new_n9802), .Y(new_n20156));
  nor_5  g17808(.A(new_n9808), .B(new_n9803), .Y(new_n20157));
  nor_5  g17809(.A(new_n20157), .B(new_n20147), .Y(new_n20158));
  nand_5 g17810(.A(new_n20146), .B(new_n11004), .Y(new_n20159));
  nand_5 g17811(.A(new_n9808), .B(new_n6138), .Y(new_n20160));
  nand_5 g17812(.A(new_n9807), .B(new_n6137), .Y(new_n20161));
  nand_5 g17813(.A(new_n20161), .B(new_n20160), .Y(new_n20162));
  xor_4  g17814(.A(new_n20145), .B(new_n9803), .Y(new_n20163));
  or_6   g17815(.A(new_n20163), .B(new_n20162), .Y(new_n20164));
  nand_5 g17816(.A(new_n20164), .B(new_n20160), .Y(new_n20165));
  and_6  g17817(.A(new_n20165), .B(new_n20159), .Y(new_n20166));
  nor_5  g17818(.A(new_n20166), .B(new_n20158), .Y(new_n20167));
  xor_4  g17819(.A(new_n20155), .B(new_n9801), .Y(new_n20168));
  nor_5  g17820(.A(new_n20168), .B(new_n20167), .Y(new_n20169));
  or_6   g17821(.A(new_n20169), .B(new_n20156), .Y(new_n20170));
  xor_4  g17822(.A(new_n20170), .B(new_n20154), .Y(new_n20171));
  xor_4  g17823(.A(new_n20171), .B(new_n9823), .Y(po0339));
  nand_5 g17824(.A(new_n13850), .B(new_n4050), .Y(new_n20173));
  or_6   g17825(.A(new_n13851), .B(pi274), .Y(new_n20174));
  nand_5 g17826(.A(new_n20174), .B(new_n20173), .Y(new_n20175));
  nand_5 g17827(.A(new_n20175), .B(new_n11643), .Y(new_n20176));
  xor_4  g17828(.A(new_n20175), .B(new_n4304), .Y(new_n20177));
  or_6   g17829(.A(new_n20177), .B(pi031), .Y(new_n20178));
  nand_5 g17830(.A(new_n20178), .B(new_n20176), .Y(new_n20179));
  nand_5 g17831(.A(new_n20179), .B(new_n4441), .Y(new_n20180));
  xor_4  g17832(.A(new_n20179), .B(new_n4312), .Y(new_n20181));
  or_6   g17833(.A(new_n20181), .B(pi310), .Y(new_n20182));
  nand_5 g17834(.A(new_n20182), .B(new_n20180), .Y(new_n20183));
  nor_5  g17835(.A(new_n20183), .B(new_n4436), .Y(new_n20184));
  nand_5 g17836(.A(new_n20183), .B(new_n4436), .Y(new_n20185));
  nand_5 g17837(.A(new_n20185), .B(pi586), .Y(new_n20186));
  not_8  g17838(.A(new_n20186), .Y(new_n20187));
  nor_5  g17839(.A(new_n20187), .B(new_n20184), .Y(new_n20188));
  xor_4  g17840(.A(new_n20188), .B(new_n11640), .Y(new_n20189));
  xor_4  g17841(.A(new_n20189), .B(pi041), .Y(new_n20190));
  not_8  g17842(.A(new_n8150), .Y(new_n20191));
  nand_5 g17843(.A(new_n13869), .B(new_n10740), .Y(new_n20192));
  nand_5 g17844(.A(new_n20192), .B(new_n13868), .Y(new_n20193));
  nand_5 g17845(.A(new_n20193), .B(new_n8193), .Y(new_n20194));
  or_6   g17846(.A(new_n20193), .B(new_n8193), .Y(new_n20195));
  nand_5 g17847(.A(new_n20195), .B(new_n4382), .Y(new_n20196));
  nand_5 g17848(.A(new_n20196), .B(new_n20194), .Y(new_n20197));
  or_6   g17849(.A(new_n20197), .B(new_n8198), .Y(new_n20198));
  xor_4  g17850(.A(new_n20197), .B(new_n8198), .Y(new_n20199));
  nand_5 g17851(.A(new_n20199), .B(pi505), .Y(new_n20200));
  nand_5 g17852(.A(new_n20200), .B(new_n20198), .Y(new_n20201));
  or_6   g17853(.A(new_n20201), .B(new_n8204), .Y(new_n20202));
  nand_5 g17854(.A(new_n20202), .B(pi368), .Y(new_n20203));
  nand_5 g17855(.A(new_n20201), .B(new_n8204), .Y(new_n20204));
  nand_5 g17856(.A(new_n20204), .B(new_n20203), .Y(new_n20205));
  nand_5 g17857(.A(new_n20205), .B(new_n20191), .Y(new_n20206));
  not_8  g17858(.A(new_n20206), .Y(new_n20207));
  nor_5  g17859(.A(new_n20205), .B(new_n20191), .Y(new_n20208));
  nor_5  g17860(.A(new_n20208), .B(new_n20207), .Y(new_n20209));
  xor_4  g17861(.A(new_n20209), .B(new_n4511), .Y(new_n20210));
  xnor_4 g17862(.A(new_n20210), .B(new_n20190), .Y(new_n20211));
  nand_5 g17863(.A(new_n20204), .B(new_n20202), .Y(new_n20212));
  xor_4  g17864(.A(new_n20212), .B(new_n4374), .Y(new_n20213));
  xor_4  g17865(.A(new_n20183), .B(new_n4317), .Y(new_n20214));
  xor_4  g17866(.A(new_n20214), .B(pi586), .Y(new_n20215));
  nand_5 g17867(.A(new_n20215), .B(new_n20213), .Y(new_n20216));
  xor_4  g17868(.A(new_n20215), .B(new_n20213), .Y(new_n20217));
  xor_4  g17869(.A(new_n20199), .B(pi505), .Y(new_n20218));
  not_8  g17870(.A(new_n20218), .Y(new_n20219));
  xor_4  g17871(.A(new_n20181), .B(new_n8152), .Y(new_n20220));
  nor_5  g17872(.A(new_n20220), .B(new_n20219), .Y(new_n20221));
  xor_4  g17873(.A(new_n20220), .B(new_n20218), .Y(new_n20222));
  xor_4  g17874(.A(new_n20177), .B(new_n10039), .Y(new_n20223));
  nand_5 g17875(.A(new_n20195), .B(new_n20194), .Y(new_n20224));
  xor_4  g17876(.A(new_n20224), .B(pi473), .Y(new_n20225));
  nand_5 g17877(.A(new_n20225), .B(new_n20223), .Y(new_n20226));
  xnor_4 g17878(.A(new_n20225), .B(new_n20223), .Y(new_n20227));
  and_6  g17879(.A(new_n13871), .B(new_n13852), .Y(new_n20228));
  nor_5  g17880(.A(new_n13910), .B(new_n13872), .Y(new_n20229));
  nor_5  g17881(.A(new_n20229), .B(new_n20228), .Y(new_n20230));
  or_6   g17882(.A(new_n20230), .B(new_n20227), .Y(new_n20231));
  nand_5 g17883(.A(new_n20231), .B(new_n20226), .Y(new_n20232));
  nor_5  g17884(.A(new_n20232), .B(new_n20222), .Y(new_n20233));
  or_6   g17885(.A(new_n20233), .B(new_n20221), .Y(new_n20234));
  nand_5 g17886(.A(new_n20234), .B(new_n20217), .Y(new_n20235));
  nand_5 g17887(.A(new_n20235), .B(new_n20216), .Y(new_n20236));
  xnor_4 g17888(.A(new_n20236), .B(new_n20211), .Y(po0340));
  xor_4  g17889(.A(new_n19938), .B(new_n17128), .Y(po0341));
  not_8  g17890(.A(new_n18901), .Y(new_n20239));
  xor_4  g17891(.A(new_n20239), .B(new_n18900), .Y(po0342));
  nand_5 g17892(.A(new_n9229), .B(new_n9235), .Y(new_n20241));
  nor_5  g17893(.A(new_n20241), .B(pi480), .Y(new_n20242));
  nand_5 g17894(.A(new_n20242), .B(new_n9226), .Y(new_n20243));
  not_8  g17895(.A(new_n20243), .Y(new_n20244));
  nand_5 g17896(.A(new_n20244), .B(new_n9223), .Y(new_n20245));
  nor_5  g17897(.A(new_n20245), .B(pi363), .Y(new_n20246));
  nand_5 g17898(.A(new_n20246), .B(new_n9217), .Y(new_n20247));
  nor_5  g17899(.A(new_n20247), .B(pi203), .Y(new_n20248));
  nand_5 g17900(.A(new_n20248), .B(new_n9210), .Y(new_n20249));
  xor_4  g17901(.A(new_n20249), .B(pi713), .Y(new_n20250));
  xor_4  g17902(.A(new_n20250), .B(new_n17689), .Y(new_n20251));
  xor_4  g17903(.A(new_n20246), .B(pi451), .Y(new_n20252));
  nor_5  g17904(.A(new_n20252), .B(new_n10856), .Y(new_n20253));
  xor_4  g17905(.A(new_n20245), .B(pi363), .Y(new_n20254));
  and_6  g17906(.A(new_n20254), .B(new_n10882), .Y(new_n20255));
  xor_4  g17907(.A(new_n20254), .B(new_n10882), .Y(new_n20256));
  not_8  g17908(.A(new_n20256), .Y(new_n20257));
  nand_5 g17909(.A(new_n10929), .B(new_n9235), .Y(new_n20258));
  not_8  g17910(.A(new_n20258), .Y(new_n20259));
  nand_5 g17911(.A(new_n10863), .B(new_n9232), .Y(new_n20260));
  nand_5 g17912(.A(new_n20260), .B(new_n20259), .Y(new_n20261));
  nand_5 g17913(.A(new_n15493), .B(pi480), .Y(new_n20262));
  nand_5 g17914(.A(new_n20262), .B(new_n20258), .Y(new_n20263));
  nand_5 g17915(.A(new_n20263), .B(new_n20261), .Y(new_n20264));
  xor_4  g17916(.A(new_n20264), .B(pi090), .Y(new_n20265));
  xor_4  g17917(.A(new_n20265), .B(new_n10858), .Y(new_n20266));
  nand_5 g17918(.A(new_n9232), .B(pi090), .Y(new_n20267));
  nor_5  g17919(.A(new_n20267), .B(new_n20266), .Y(new_n20268));
  nand_5 g17920(.A(new_n10863), .B(new_n10929), .Y(new_n20269));
  nand_5 g17921(.A(new_n20269), .B(new_n20265), .Y(new_n20270));
  nand_5 g17922(.A(new_n20270), .B(new_n10859), .Y(new_n20271));
  nor_5  g17923(.A(new_n20242), .B(pi090), .Y(new_n20272));
  nand_5 g17924(.A(new_n20272), .B(new_n20264), .Y(new_n20273));
  nand_5 g17925(.A(new_n20273), .B(new_n20271), .Y(new_n20274));
  nor_5  g17926(.A(new_n20274), .B(new_n20268), .Y(new_n20275));
  nor_5  g17927(.A(new_n20275), .B(new_n10872), .Y(new_n20276));
  not_8  g17928(.A(new_n20276), .Y(new_n20277));
  xor_4  g17929(.A(new_n20242), .B(pi343), .Y(new_n20278));
  xor_4  g17930(.A(new_n20275), .B(new_n10873), .Y(new_n20279));
  or_6   g17931(.A(new_n20279), .B(new_n20278), .Y(new_n20280));
  nand_5 g17932(.A(new_n20280), .B(new_n20277), .Y(new_n20281));
  nor_5  g17933(.A(new_n20281), .B(new_n20244), .Y(new_n20282));
  nand_5 g17934(.A(new_n20276), .B(new_n9226), .Y(new_n20283));
  xor_4  g17935(.A(new_n10857), .B(pi104), .Y(new_n20284));
  not_8  g17936(.A(new_n20284), .Y(new_n20285));
  nand_5 g17937(.A(new_n20285), .B(new_n20283), .Y(new_n20286));
  nor_5  g17938(.A(new_n20286), .B(new_n20282), .Y(new_n20287));
  nand_5 g17939(.A(new_n20284), .B(new_n20243), .Y(new_n20288));
  nand_5 g17940(.A(new_n20285), .B(new_n20242), .Y(new_n20289));
  nand_5 g17941(.A(new_n20289), .B(new_n20288), .Y(new_n20290));
  nor_5  g17942(.A(new_n20290), .B(new_n20277), .Y(new_n20291));
  nor_5  g17943(.A(new_n20291), .B(new_n20287), .Y(new_n20292));
  nand_5 g17944(.A(new_n20292), .B(new_n15492), .Y(new_n20293));
  nand_5 g17945(.A(new_n20284), .B(new_n20282), .Y(new_n20294));
  nand_5 g17946(.A(new_n20294), .B(new_n20292), .Y(new_n20295));
  and_6  g17947(.A(new_n20295), .B(new_n10857), .Y(new_n20296));
  or_6   g17948(.A(new_n20296), .B(new_n20281), .Y(new_n20297));
  nand_5 g17949(.A(new_n20297), .B(new_n20293), .Y(new_n20298));
  nor_5  g17950(.A(new_n20298), .B(new_n20257), .Y(new_n20299));
  nor_5  g17951(.A(new_n20299), .B(new_n20255), .Y(new_n20300));
  xor_4  g17952(.A(new_n20252), .B(new_n10855), .Y(new_n20301));
  nor_5  g17953(.A(new_n20301), .B(new_n20300), .Y(new_n20302));
  nor_5  g17954(.A(new_n20302), .B(new_n20253), .Y(new_n20303));
  nor_5  g17955(.A(new_n20303), .B(new_n10898), .Y(new_n20304));
  xor_4  g17956(.A(new_n20247), .B(new_n9213), .Y(new_n20305));
  xor_4  g17957(.A(new_n20303), .B(new_n10897), .Y(new_n20306));
  nor_5  g17958(.A(new_n20306), .B(new_n20305), .Y(new_n20307));
  or_6   g17959(.A(new_n20307), .B(new_n20304), .Y(new_n20308));
  xor_4  g17960(.A(new_n20308), .B(new_n10907), .Y(new_n20309));
  nor_5  g17961(.A(new_n20248), .B(new_n9210), .Y(new_n20310));
  nand_5 g17962(.A(new_n20310), .B(new_n20309), .Y(new_n20311));
  nand_5 g17963(.A(new_n20304), .B(new_n10907), .Y(new_n20312));
  or_6   g17964(.A(new_n20308), .B(new_n10907), .Y(new_n20313));
  nand_5 g17965(.A(new_n20313), .B(new_n20249), .Y(new_n20314));
  nand_5 g17966(.A(new_n20314), .B(new_n20312), .Y(new_n20315));
  nand_5 g17967(.A(new_n20315), .B(new_n20311), .Y(new_n20316));
  nor_5  g17968(.A(new_n20316), .B(new_n20251), .Y(new_n20317));
  nand_5 g17969(.A(new_n20249), .B(pi713), .Y(new_n20318));
  nand_5 g17970(.A(new_n20250), .B(new_n17689), .Y(new_n20319));
  nand_5 g17971(.A(new_n20319), .B(new_n20318), .Y(new_n20320));
  xor_4  g17972(.A(new_n20320), .B(new_n17710), .Y(new_n20321));
  xor_4  g17973(.A(new_n20321), .B(new_n20317), .Y(new_n20322));
  not_8  g17974(.A(new_n19582), .Y(new_n20323));
  xor_4  g17975(.A(new_n20301), .B(new_n20300), .Y(new_n20324));
  nor_5  g17976(.A(new_n10929), .B(new_n9235), .Y(new_n20325));
  or_6   g17977(.A(new_n20325), .B(new_n20259), .Y(new_n20326));
  nor_5  g17978(.A(new_n20326), .B(new_n9456), .Y(new_n20327));
  nor_5  g17979(.A(new_n20327), .B(new_n20325), .Y(new_n20328));
  nand_5 g17980(.A(new_n20262), .B(new_n20260), .Y(new_n20329));
  xor_4  g17981(.A(new_n20329), .B(new_n9444), .Y(new_n20330));
  nor_5  g17982(.A(new_n20330), .B(new_n20328), .Y(new_n20331));
  or_6   g17983(.A(new_n20329), .B(new_n9445), .Y(new_n20332));
  nand_5 g17984(.A(new_n20329), .B(new_n20259), .Y(new_n20333));
  nand_5 g17985(.A(new_n20333), .B(new_n20332), .Y(new_n20334));
  nor_5  g17986(.A(new_n20334), .B(new_n20331), .Y(new_n20335));
  nor_5  g17987(.A(new_n20335), .B(new_n9443), .Y(new_n20336));
  and_6  g17988(.A(new_n20335), .B(new_n9443), .Y(new_n20337));
  nor_5  g17989(.A(new_n20337), .B(new_n20266), .Y(new_n20338));
  nor_5  g17990(.A(new_n20338), .B(new_n20336), .Y(new_n20339));
  nand_5 g17991(.A(new_n20339), .B(new_n9409), .Y(new_n20340));
  xor_4  g17992(.A(new_n20279), .B(new_n20278), .Y(new_n20341));
  xor_4  g17993(.A(new_n20339), .B(new_n9409), .Y(new_n20342));
  nand_5 g17994(.A(new_n20342), .B(new_n20341), .Y(new_n20343));
  nand_5 g17995(.A(new_n20343), .B(new_n20340), .Y(new_n20344));
  not_8  g17996(.A(new_n20344), .Y(new_n20345));
  nand_5 g17997(.A(new_n20345), .B(new_n20295), .Y(new_n20346));
  xor_4  g17998(.A(new_n20344), .B(new_n20295), .Y(new_n20347));
  or_6   g17999(.A(new_n20347), .B(new_n9482), .Y(new_n20348));
  nand_5 g18000(.A(new_n20348), .B(new_n20346), .Y(new_n20349));
  nor_5  g18001(.A(new_n20349), .B(new_n9520), .Y(new_n20350));
  xor_4  g18002(.A(new_n20349), .B(new_n9520), .Y(new_n20351));
  not_8  g18003(.A(new_n20351), .Y(new_n20352));
  xor_4  g18004(.A(new_n20298), .B(new_n20256), .Y(new_n20353));
  nor_5  g18005(.A(new_n20353), .B(new_n20352), .Y(new_n20354));
  or_6   g18006(.A(new_n20354), .B(new_n20350), .Y(new_n20355));
  nand_5 g18007(.A(new_n20355), .B(new_n20324), .Y(new_n20356));
  xor_4  g18008(.A(new_n20355), .B(new_n20324), .Y(new_n20357));
  nand_5 g18009(.A(new_n20357), .B(new_n19571), .Y(new_n20358));
  nand_5 g18010(.A(new_n20358), .B(new_n20356), .Y(new_n20359));
  nor_5  g18011(.A(new_n20359), .B(new_n19567), .Y(new_n20360));
  not_8  g18012(.A(new_n19567), .Y(new_n20361));
  xor_4  g18013(.A(new_n20359), .B(new_n20361), .Y(new_n20362));
  xor_4  g18014(.A(new_n20306), .B(new_n20305), .Y(new_n20363));
  nor_5  g18015(.A(new_n20363), .B(new_n20362), .Y(new_n20364));
  or_6   g18016(.A(new_n20364), .B(new_n20360), .Y(new_n20365));
  nor_5  g18017(.A(new_n20365), .B(new_n19562), .Y(new_n20366));
  xor_4  g18018(.A(new_n20248), .B(new_n9210), .Y(new_n20367));
  xor_4  g18019(.A(new_n20367), .B(new_n20309), .Y(new_n20368));
  xor_4  g18020(.A(new_n20365), .B(new_n19562), .Y(new_n20369));
  and_6  g18021(.A(new_n20369), .B(new_n20368), .Y(new_n20370));
  nor_5  g18022(.A(new_n20370), .B(new_n20366), .Y(new_n20371));
  nand_5 g18023(.A(new_n20371), .B(new_n20323), .Y(new_n20372));
  not_8  g18024(.A(new_n20372), .Y(new_n20373));
  nor_5  g18025(.A(new_n20371), .B(new_n20323), .Y(new_n20374));
  xor_4  g18026(.A(new_n20316), .B(new_n20251), .Y(new_n20375));
  nor_5  g18027(.A(new_n20375), .B(new_n20374), .Y(new_n20376));
  nor_5  g18028(.A(new_n20376), .B(new_n20373), .Y(new_n20377));
  nand_5 g18029(.A(new_n20377), .B(new_n20322), .Y(new_n20378));
  nor_5  g18030(.A(new_n20378), .B(new_n19538), .Y(new_n20379));
  not_8  g18031(.A(new_n19558), .Y(new_n20380));
  xor_4  g18032(.A(new_n20377), .B(new_n20322), .Y(new_n20381));
  nor_5  g18033(.A(new_n20381), .B(new_n20380), .Y(new_n20382));
  or_6   g18034(.A(new_n20382), .B(new_n19557), .Y(new_n20383));
  and_6  g18035(.A(new_n20383), .B(new_n20378), .Y(new_n20384));
  nor_5  g18036(.A(new_n20384), .B(new_n20379), .Y(new_n20385));
  nand_5 g18037(.A(new_n20320), .B(new_n18170), .Y(new_n20386));
  nor_5  g18038(.A(new_n20386), .B(new_n20317), .Y(new_n20387));
  nor_5  g18039(.A(new_n20320), .B(new_n18170), .Y(new_n20388));
  nand_5 g18040(.A(new_n20388), .B(new_n20317), .Y(new_n20389));
  not_8  g18041(.A(new_n20389), .Y(new_n20390));
  nor_5  g18042(.A(new_n20390), .B(new_n20387), .Y(new_n20391));
  xor_4  g18043(.A(new_n20391), .B(new_n20385), .Y(po0343));
  xnor_4 g18044(.A(new_n2775), .B(new_n2774), .Y(po0344));
  xor_4  g18045(.A(pi507), .B(new_n8328), .Y(new_n20394));
  nand_5 g18046(.A(new_n8332), .B(pi324), .Y(new_n20395));
  xor_4  g18047(.A(pi738), .B(new_n2468), .Y(new_n20396));
  nand_5 g18048(.A(pi790), .B(new_n8336), .Y(new_n20397));
  nand_5 g18049(.A(new_n7010), .B(pi316), .Y(new_n20398));
  nand_5 g18050(.A(pi102), .B(new_n7013), .Y(new_n20399));
  xor_4  g18051(.A(pi102), .B(new_n7013), .Y(new_n20400));
  nand_5 g18052(.A(new_n7016), .B(pi204), .Y(new_n20401));
  or_6   g18053(.A(new_n19242), .B(new_n19240), .Y(new_n20402));
  nand_5 g18054(.A(new_n20402), .B(new_n20401), .Y(new_n20403));
  nand_5 g18055(.A(new_n20403), .B(new_n20400), .Y(new_n20404));
  nand_5 g18056(.A(new_n20404), .B(new_n20399), .Y(new_n20405));
  xor_4  g18057(.A(pi747), .B(new_n2474), .Y(new_n20406));
  nand_5 g18058(.A(new_n20406), .B(new_n20405), .Y(new_n20407));
  nand_5 g18059(.A(new_n20407), .B(new_n20398), .Y(new_n20408));
  xor_4  g18060(.A(pi790), .B(new_n8336), .Y(new_n20409));
  nand_5 g18061(.A(new_n20409), .B(new_n20408), .Y(new_n20410));
  nand_5 g18062(.A(new_n20410), .B(new_n20397), .Y(new_n20411));
  nand_5 g18063(.A(new_n20411), .B(new_n20396), .Y(new_n20412));
  nand_5 g18064(.A(new_n20412), .B(new_n20395), .Y(new_n20413));
  xor_4  g18065(.A(new_n20413), .B(new_n20394), .Y(new_n20414));
  not_8  g18066(.A(new_n20414), .Y(new_n20415));
  nor_5  g18067(.A(new_n20415), .B(new_n19657), .Y(new_n20416));
  xor_4  g18068(.A(new_n20414), .B(new_n19657), .Y(new_n20417));
  xor_4  g18069(.A(new_n20411), .B(new_n20396), .Y(new_n20418));
  or_6   g18070(.A(new_n20418), .B(new_n19667), .Y(new_n20419));
  not_8  g18071(.A(new_n19338), .Y(new_n20420));
  xnor_4 g18072(.A(new_n20409), .B(new_n20408), .Y(new_n20421));
  nand_5 g18073(.A(new_n20421), .B(new_n20420), .Y(new_n20422));
  or_6   g18074(.A(new_n20421), .B(new_n20420), .Y(new_n20423));
  xor_4  g18075(.A(new_n20406), .B(new_n20405), .Y(new_n20424));
  or_6   g18076(.A(new_n20424), .B(new_n19282), .Y(new_n20425));
  xor_4  g18077(.A(new_n20424), .B(new_n19282), .Y(new_n20426));
  xor_4  g18078(.A(new_n20403), .B(new_n20400), .Y(new_n20427));
  not_8  g18079(.A(new_n20427), .Y(new_n20428));
  or_6   g18080(.A(new_n20428), .B(new_n19300), .Y(new_n20429));
  not_8  g18081(.A(new_n19243), .Y(new_n20430));
  nor_5  g18082(.A(new_n20430), .B(new_n19239), .Y(new_n20431));
  nor_5  g18083(.A(new_n19256), .B(new_n19244), .Y(new_n20432));
  or_6   g18084(.A(new_n20432), .B(new_n20431), .Y(new_n20433));
  xor_4  g18085(.A(new_n20428), .B(new_n19300), .Y(new_n20434));
  nand_5 g18086(.A(new_n20434), .B(new_n20433), .Y(new_n20435));
  nand_5 g18087(.A(new_n20435), .B(new_n20429), .Y(new_n20436));
  not_8  g18088(.A(new_n20436), .Y(new_n20437));
  nand_5 g18089(.A(new_n20437), .B(new_n20426), .Y(new_n20438));
  nand_5 g18090(.A(new_n20438), .B(new_n20425), .Y(new_n20439));
  nand_5 g18091(.A(new_n20439), .B(new_n20423), .Y(new_n20440));
  nand_5 g18092(.A(new_n20440), .B(new_n20422), .Y(new_n20441));
  xor_4  g18093(.A(new_n20418), .B(new_n19667), .Y(new_n20442));
  nand_5 g18094(.A(new_n20442), .B(new_n20441), .Y(new_n20443));
  nand_5 g18095(.A(new_n20443), .B(new_n20419), .Y(new_n20444));
  nor_5  g18096(.A(new_n20444), .B(new_n20417), .Y(new_n20445));
  or_6   g18097(.A(new_n20445), .B(new_n20416), .Y(new_n20446));
  xor_4  g18098(.A(pi775), .B(pi537), .Y(new_n20447));
  nand_5 g18099(.A(new_n16177), .B(new_n6953), .Y(new_n20448));
  nand_5 g18100(.A(new_n19645), .B(new_n19636), .Y(new_n20449));
  nand_5 g18101(.A(new_n20449), .B(new_n20448), .Y(new_n20450));
  xor_4  g18102(.A(new_n20450), .B(new_n20447), .Y(new_n20451));
  not_8  g18103(.A(new_n20451), .Y(new_n20452));
  xor_4  g18104(.A(new_n20452), .B(new_n7560), .Y(new_n20453));
  nor_5  g18105(.A(new_n19647), .B(new_n7564), .Y(new_n20454));
  not_8  g18106(.A(new_n19648), .Y(new_n20455));
  nor_5  g18107(.A(new_n19656), .B(new_n20455), .Y(new_n20456));
  or_6   g18108(.A(new_n20456), .B(new_n20454), .Y(new_n20457));
  xnor_4 g18109(.A(new_n20457), .B(new_n20453), .Y(new_n20458));
  nand_5 g18110(.A(pi507), .B(new_n8328), .Y(new_n20459));
  nand_5 g18111(.A(new_n20413), .B(new_n20394), .Y(new_n20460));
  nand_5 g18112(.A(new_n20460), .B(new_n20459), .Y(new_n20461));
  not_8  g18113(.A(pi009), .Y(new_n20462));
  nand_5 g18114(.A(pi446), .B(new_n20462), .Y(new_n20463));
  nand_5 g18115(.A(new_n3525), .B(pi009), .Y(new_n20464));
  nand_5 g18116(.A(new_n20464), .B(new_n20463), .Y(new_n20465));
  xor_4  g18117(.A(new_n20465), .B(new_n20461), .Y(new_n20466));
  xor_4  g18118(.A(new_n20466), .B(new_n20458), .Y(new_n20467));
  xnor_4 g18119(.A(new_n20467), .B(new_n20446), .Y(po0345));
  xnor_4 g18120(.A(new_n6527), .B(new_n4579), .Y(po0346));
  xnor_4 g18121(.A(new_n12706), .B(new_n12705), .Y(po0347));
  xnor_4 g18122(.A(new_n12177), .B(new_n12176), .Y(po0348));
  xnor_4 g18123(.A(new_n9469), .B(new_n9468), .Y(po0349));
  xor_4  g18124(.A(new_n13621), .B(new_n13611), .Y(new_n20473));
  xor_4  g18125(.A(new_n20473), .B(new_n3487), .Y(po0350));
  nand_5 g18126(.A(new_n20140), .B(new_n20137), .Y(new_n20475));
  nand_5 g18127(.A(new_n20475), .B(new_n20134), .Y(po0351));
  xor_4  g18128(.A(new_n16729), .B(new_n6173), .Y(po0352));
  xnor_4 g18129(.A(new_n12410), .B(new_n12409), .Y(po0353));
  nand_5 g18130(.A(pi827), .B(pi472), .Y(new_n20479));
  not_8  g18131(.A(new_n20479), .Y(new_n20480));
  nand_5 g18132(.A(new_n5497), .B(new_n5636), .Y(new_n20481));
  nand_5 g18133(.A(new_n20481), .B(new_n20479), .Y(new_n20482));
  nor_5  g18134(.A(new_n20482), .B(pi419), .Y(new_n20483));
  nor_5  g18135(.A(new_n20483), .B(new_n20480), .Y(new_n20484));
  nand_5 g18136(.A(new_n5640), .B(new_n5499), .Y(new_n20485));
  nand_5 g18137(.A(pi834), .B(pi737), .Y(new_n20486));
  nand_5 g18138(.A(new_n20486), .B(new_n20485), .Y(new_n20487));
  nand_5 g18139(.A(pi692), .B(pi297), .Y(new_n20488));
  not_8  g18140(.A(new_n20488), .Y(new_n20489));
  nor_5  g18141(.A(pi692), .B(pi297), .Y(new_n20490));
  nor_5  g18142(.A(new_n5507), .B(new_n5646), .Y(new_n20491));
  nor_5  g18143(.A(new_n3991), .B(new_n5511), .Y(new_n20492));
  nor_5  g18144(.A(new_n5513), .B(new_n3993), .Y(new_n20493));
  xor_4  g18145(.A(pi739), .B(new_n3993), .Y(new_n20494));
  nand_5 g18146(.A(new_n3946), .B(new_n5517), .Y(new_n20495));
  nand_5 g18147(.A(pi362), .B(pi067), .Y(new_n20496));
  nand_5 g18148(.A(new_n15830), .B(new_n15828), .Y(new_n20497));
  nand_5 g18149(.A(new_n20497), .B(new_n15829), .Y(new_n20498));
  nand_5 g18150(.A(new_n20498), .B(new_n20496), .Y(new_n20499));
  nand_5 g18151(.A(new_n20499), .B(new_n20495), .Y(new_n20500));
  nor_5  g18152(.A(new_n20500), .B(new_n20494), .Y(new_n20501));
  nor_5  g18153(.A(new_n20501), .B(new_n20493), .Y(new_n20502));
  xor_4  g18154(.A(pi250), .B(new_n5511), .Y(new_n20503));
  nor_5  g18155(.A(new_n20503), .B(new_n20502), .Y(new_n20504));
  nor_5  g18156(.A(new_n20504), .B(new_n20492), .Y(new_n20505));
  xor_4  g18157(.A(pi625), .B(new_n5646), .Y(new_n20506));
  nor_5  g18158(.A(new_n20506), .B(new_n20505), .Y(new_n20507));
  nor_5  g18159(.A(new_n20507), .B(new_n20491), .Y(new_n20508));
  nor_5  g18160(.A(new_n20508), .B(new_n20490), .Y(new_n20509));
  nor_5  g18161(.A(new_n20509), .B(new_n20489), .Y(new_n20510));
  xor_4  g18162(.A(new_n20510), .B(new_n20487), .Y(new_n20511));
  nand_5 g18163(.A(new_n20511), .B(new_n14078), .Y(new_n20512));
  not_8  g18164(.A(new_n20512), .Y(new_n20513));
  xor_4  g18165(.A(new_n20511), .B(new_n14078), .Y(new_n20514));
  not_8  g18166(.A(new_n20514), .Y(new_n20515));
  nor_5  g18167(.A(new_n20490), .B(new_n20489), .Y(new_n20516));
  xor_4  g18168(.A(new_n20516), .B(new_n20508), .Y(new_n20517));
  or_6   g18169(.A(new_n20517), .B(pi647), .Y(new_n20518));
  not_8  g18170(.A(new_n20518), .Y(new_n20519));
  xor_4  g18171(.A(new_n20517), .B(pi647), .Y(new_n20520));
  not_8  g18172(.A(new_n20520), .Y(new_n20521));
  xor_4  g18173(.A(new_n20506), .B(new_n20505), .Y(new_n20522));
  or_6   g18174(.A(new_n20522), .B(new_n4060), .Y(new_n20523));
  xor_4  g18175(.A(new_n20522), .B(new_n4060), .Y(new_n20524));
  xnor_4 g18176(.A(new_n20503), .B(new_n20502), .Y(new_n20525));
  nor_5  g18177(.A(new_n20525), .B(pi602), .Y(new_n20526));
  xor_4  g18178(.A(new_n20525), .B(pi602), .Y(new_n20527));
  xor_4  g18179(.A(new_n20500), .B(new_n20494), .Y(new_n20528));
  nor_5  g18180(.A(new_n20528), .B(new_n3962), .Y(new_n20529));
  nand_5 g18181(.A(new_n20496), .B(new_n20495), .Y(new_n20530));
  xnor_4 g18182(.A(new_n20530), .B(new_n20498), .Y(new_n20531));
  nand_5 g18183(.A(new_n20531), .B(pi271), .Y(new_n20532));
  xor_4  g18184(.A(new_n20531), .B(pi271), .Y(new_n20533));
  and_6  g18185(.A(new_n15833), .B(pi218), .Y(new_n20534));
  nor_5  g18186(.A(new_n15835), .B(new_n15833), .Y(new_n20535));
  or_6   g18187(.A(new_n20535), .B(new_n20534), .Y(new_n20536));
  nand_5 g18188(.A(new_n20536), .B(new_n20533), .Y(new_n20537));
  nand_5 g18189(.A(new_n20537), .B(new_n20532), .Y(new_n20538));
  xor_4  g18190(.A(new_n20528), .B(pi614), .Y(new_n20539));
  not_8  g18191(.A(new_n20539), .Y(new_n20540));
  nand_5 g18192(.A(new_n20540), .B(new_n20538), .Y(new_n20541));
  not_8  g18193(.A(new_n20541), .Y(new_n20542));
  nor_5  g18194(.A(new_n20542), .B(new_n20529), .Y(new_n20543));
  and_6  g18195(.A(new_n20543), .B(new_n20527), .Y(new_n20544));
  nor_5  g18196(.A(new_n20544), .B(new_n20526), .Y(new_n20545));
  nand_5 g18197(.A(new_n20545), .B(new_n20524), .Y(new_n20546));
  nand_5 g18198(.A(new_n20546), .B(new_n20523), .Y(new_n20547));
  nor_5  g18199(.A(new_n20547), .B(new_n20521), .Y(new_n20548));
  nor_5  g18200(.A(new_n20548), .B(new_n20519), .Y(new_n20549));
  nor_5  g18201(.A(new_n20549), .B(new_n20515), .Y(new_n20550));
  nor_5  g18202(.A(new_n20550), .B(new_n20513), .Y(new_n20551));
  not_8  g18203(.A(new_n20551), .Y(new_n20552));
  not_8  g18204(.A(new_n20486), .Y(new_n20553));
  not_8  g18205(.A(new_n20485), .Y(new_n20554));
  nor_5  g18206(.A(new_n20510), .B(new_n20554), .Y(new_n20555));
  nor_5  g18207(.A(new_n20555), .B(new_n20553), .Y(new_n20556));
  not_8  g18208(.A(new_n20556), .Y(new_n20557));
  nand_5 g18209(.A(new_n20557), .B(new_n20552), .Y(new_n20558));
  or_6   g18210(.A(new_n20558), .B(new_n20484), .Y(new_n20559));
  not_8  g18211(.A(new_n20559), .Y(new_n20560));
  nand_5 g18212(.A(new_n20556), .B(new_n20551), .Y(new_n20561));
  not_8  g18213(.A(new_n20561), .Y(new_n20562));
  nand_5 g18214(.A(new_n20480), .B(new_n14174), .Y(new_n20563));
  nor_5  g18215(.A(new_n20563), .B(new_n20562), .Y(new_n20564));
  nor_5  g18216(.A(new_n20564), .B(new_n20560), .Y(new_n20565));
  not_8  g18217(.A(new_n20565), .Y(new_n20566));
  nand_5 g18218(.A(new_n20562), .B(new_n20484), .Y(new_n20567));
  nor_5  g18219(.A(new_n20481), .B(new_n14174), .Y(new_n20568));
  nand_5 g18220(.A(new_n20568), .B(new_n20558), .Y(new_n20569));
  nand_5 g18221(.A(new_n20569), .B(new_n20567), .Y(new_n20570));
  nor_5  g18222(.A(new_n20570), .B(new_n20566), .Y(new_n20571));
  xor_4  g18223(.A(pi405), .B(pi056), .Y(new_n20572));
  xor_4  g18224(.A(new_n20572), .B(pi282), .Y(new_n20573));
  xor_4  g18225(.A(new_n20573), .B(new_n20571), .Y(new_n20574));
  nand_5 g18226(.A(new_n20574), .B(new_n20190), .Y(new_n20575));
  xnor_4 g18227(.A(new_n20574), .B(new_n20190), .Y(new_n20576));
  nand_5 g18228(.A(new_n20561), .B(new_n20558), .Y(new_n20577));
  xor_4  g18229(.A(new_n20482), .B(new_n14174), .Y(new_n20578));
  xor_4  g18230(.A(new_n20578), .B(new_n20577), .Y(new_n20579));
  nand_5 g18231(.A(new_n20579), .B(new_n20215), .Y(new_n20580));
  xor_4  g18232(.A(new_n20579), .B(new_n20215), .Y(new_n20581));
  xor_4  g18233(.A(new_n20549), .B(new_n20514), .Y(new_n20582));
  nand_5 g18234(.A(new_n20582), .B(new_n20220), .Y(new_n20583));
  not_8  g18235(.A(new_n20583), .Y(new_n20584));
  xnor_4 g18236(.A(new_n20582), .B(new_n20220), .Y(new_n20585));
  xor_4  g18237(.A(new_n20547), .B(new_n20520), .Y(new_n20586));
  and_6  g18238(.A(new_n20586), .B(new_n20223), .Y(new_n20587));
  xor_4  g18239(.A(new_n20545), .B(new_n20524), .Y(new_n20588));
  and_6  g18240(.A(new_n20588), .B(new_n13852), .Y(new_n20589));
  xnor_4 g18241(.A(new_n20588), .B(new_n13852), .Y(new_n20590));
  not_8  g18242(.A(new_n20527), .Y(new_n20591));
  xor_4  g18243(.A(new_n20543), .B(new_n20591), .Y(new_n20592));
  not_8  g18244(.A(new_n20592), .Y(new_n20593));
  nor_5  g18245(.A(new_n20593), .B(new_n13874), .Y(new_n20594));
  xor_4  g18246(.A(new_n20539), .B(new_n20538), .Y(new_n20595));
  not_8  g18247(.A(new_n20595), .Y(new_n20596));
  or_6   g18248(.A(new_n20596), .B(new_n13880), .Y(new_n20597));
  nor_5  g18249(.A(new_n20535), .B(new_n20534), .Y(new_n20598));
  xor_4  g18250(.A(new_n20598), .B(new_n20533), .Y(new_n20599));
  not_8  g18251(.A(new_n20599), .Y(new_n20600));
  nor_5  g18252(.A(new_n20600), .B(new_n13885), .Y(new_n20601));
  nor_5  g18253(.A(new_n15841), .B(new_n13901), .Y(new_n20602));
  nand_5 g18254(.A(new_n15838), .B(new_n15835), .Y(new_n20603));
  and_6  g18255(.A(new_n20603), .B(new_n15837), .Y(new_n20604));
  and_6  g18256(.A(new_n20604), .B(new_n15841), .Y(new_n20605));
  nor_5  g18257(.A(new_n20605), .B(new_n20602), .Y(new_n20606));
  xor_4  g18258(.A(new_n20599), .B(new_n13885), .Y(new_n20607));
  nor_5  g18259(.A(new_n20607), .B(new_n20606), .Y(new_n20608));
  or_6   g18260(.A(new_n20608), .B(new_n20601), .Y(new_n20609));
  xor_4  g18261(.A(new_n20595), .B(new_n13880), .Y(new_n20610));
  not_8  g18262(.A(new_n20610), .Y(new_n20611));
  nand_5 g18263(.A(new_n20611), .B(new_n20609), .Y(new_n20612));
  nand_5 g18264(.A(new_n20612), .B(new_n20597), .Y(new_n20613));
  xor_4  g18265(.A(new_n20592), .B(new_n13874), .Y(new_n20614));
  nor_5  g18266(.A(new_n20614), .B(new_n20613), .Y(new_n20615));
  nor_5  g18267(.A(new_n20615), .B(new_n20594), .Y(new_n20616));
  nor_5  g18268(.A(new_n20616), .B(new_n20590), .Y(new_n20617));
  nor_5  g18269(.A(new_n20617), .B(new_n20589), .Y(new_n20618));
  xnor_4 g18270(.A(new_n20586), .B(new_n20223), .Y(new_n20619));
  nor_5  g18271(.A(new_n20619), .B(new_n20618), .Y(new_n20620));
  nor_5  g18272(.A(new_n20620), .B(new_n20587), .Y(new_n20621));
  nor_5  g18273(.A(new_n20621), .B(new_n20585), .Y(new_n20622));
  nor_5  g18274(.A(new_n20622), .B(new_n20584), .Y(new_n20623));
  nand_5 g18275(.A(new_n20623), .B(new_n20581), .Y(new_n20624));
  nand_5 g18276(.A(new_n20624), .B(new_n20580), .Y(new_n20625));
  or_6   g18277(.A(new_n20625), .B(new_n20576), .Y(new_n20626));
  nand_5 g18278(.A(new_n20626), .B(new_n20575), .Y(new_n20627));
  nand_5 g18279(.A(new_n20188), .B(new_n11640), .Y(new_n20628));
  nand_5 g18280(.A(new_n20189), .B(new_n8209), .Y(new_n20629));
  nand_5 g18281(.A(new_n20629), .B(new_n20628), .Y(new_n20630));
  xor_4  g18282(.A(new_n20630), .B(new_n4278), .Y(new_n20631));
  not_8  g18283(.A(new_n20631), .Y(new_n20632));
  nand_5 g18284(.A(pi405), .B(pi282), .Y(new_n20633));
  nand_5 g18285(.A(new_n5546), .B(new_n5634), .Y(new_n20634));
  nand_5 g18286(.A(new_n20634), .B(new_n6372), .Y(new_n20635));
  nand_5 g18287(.A(new_n20635), .B(new_n20633), .Y(new_n20636));
  not_8  g18288(.A(new_n20636), .Y(new_n20637));
  nand_5 g18289(.A(new_n20637), .B(new_n20570), .Y(new_n20638));
  nor_5  g18290(.A(new_n20634), .B(new_n6372), .Y(new_n20639));
  nand_5 g18291(.A(new_n20639), .B(new_n20565), .Y(new_n20640));
  nand_5 g18292(.A(new_n20640), .B(new_n20638), .Y(new_n20641));
  not_8  g18293(.A(new_n20641), .Y(new_n20642));
  or_6   g18294(.A(new_n20633), .B(pi056), .Y(new_n20643));
  nor_5  g18295(.A(new_n20643), .B(new_n20570), .Y(new_n20644));
  nor_5  g18296(.A(new_n20637), .B(new_n20565), .Y(new_n20645));
  nor_5  g18297(.A(new_n20645), .B(new_n20644), .Y(new_n20646));
  nand_5 g18298(.A(new_n20646), .B(new_n20642), .Y(new_n20647));
  xor_4  g18299(.A(new_n20647), .B(new_n20632), .Y(new_n20648));
  xnor_4 g18300(.A(new_n20648), .B(new_n20627), .Y(po0354));
  xor_4  g18301(.A(new_n17249), .B(new_n12969), .Y(po0355));
  xor_4  g18302(.A(pi430), .B(pi403), .Y(new_n20651));
  not_8  g18303(.A(new_n20651), .Y(new_n20652));
  nor_5  g18304(.A(new_n5454), .B(new_n9174), .Y(new_n20653));
  nor_5  g18305(.A(new_n5501), .B(new_n5457), .Y(new_n20654));
  xor_4  g18306(.A(pi342), .B(pi319), .Y(new_n20655));
  not_8  g18307(.A(new_n20655), .Y(new_n20656));
  nor_5  g18308(.A(new_n5505), .B(new_n5460), .Y(new_n20657));
  xor_4  g18309(.A(pi549), .B(pi429), .Y(new_n20658));
  not_8  g18310(.A(new_n20658), .Y(new_n20659));
  nor_5  g18311(.A(new_n5463), .B(new_n5509), .Y(new_n20660));
  not_8  g18312(.A(new_n18158), .Y(new_n20661));
  nor_5  g18313(.A(new_n18160), .B(new_n20661), .Y(new_n20662));
  nor_5  g18314(.A(new_n20662), .B(new_n20660), .Y(new_n20663));
  nor_5  g18315(.A(new_n20663), .B(new_n20659), .Y(new_n20664));
  nor_5  g18316(.A(new_n20664), .B(new_n20657), .Y(new_n20665));
  nor_5  g18317(.A(new_n20665), .B(new_n20656), .Y(new_n20666));
  nor_5  g18318(.A(new_n20666), .B(new_n20654), .Y(new_n20667));
  xor_4  g18319(.A(pi777), .B(pi334), .Y(new_n20668));
  not_8  g18320(.A(new_n20668), .Y(new_n20669));
  nor_5  g18321(.A(new_n20669), .B(new_n20667), .Y(new_n20670));
  nor_5  g18322(.A(new_n20670), .B(new_n20653), .Y(new_n20671));
  xor_4  g18323(.A(new_n20671), .B(new_n20652), .Y(new_n20672));
  xor_4  g18324(.A(new_n20672), .B(new_n16065), .Y(new_n20673));
  not_8  g18325(.A(new_n20673), .Y(new_n20674));
  xor_4  g18326(.A(new_n20668), .B(new_n20667), .Y(new_n20675));
  nand_5 g18327(.A(new_n20675), .B(new_n16067), .Y(new_n20676));
  xor_4  g18328(.A(new_n20665), .B(new_n20655), .Y(new_n20677));
  nor_5  g18329(.A(new_n20677), .B(new_n16072), .Y(new_n20678));
  xor_4  g18330(.A(new_n20663), .B(new_n20658), .Y(new_n20679));
  or_6   g18331(.A(new_n20679), .B(new_n16073), .Y(new_n20680));
  xor_4  g18332(.A(new_n20679), .B(new_n16073), .Y(new_n20681));
  or_6   g18333(.A(new_n18161), .B(new_n16075), .Y(new_n20682));
  not_8  g18334(.A(new_n18165), .Y(new_n20683));
  nand_5 g18335(.A(new_n20683), .B(new_n18162), .Y(new_n20684));
  nand_5 g18336(.A(new_n20684), .B(new_n20682), .Y(new_n20685));
  nand_5 g18337(.A(new_n20685), .B(new_n20681), .Y(new_n20686));
  nand_5 g18338(.A(new_n20686), .B(new_n20680), .Y(new_n20687));
  not_8  g18339(.A(new_n20687), .Y(new_n20688));
  xnor_4 g18340(.A(new_n20677), .B(new_n16072), .Y(new_n20689));
  nor_5  g18341(.A(new_n20689), .B(new_n20688), .Y(new_n20690));
  or_6   g18342(.A(new_n20690), .B(new_n20678), .Y(new_n20691));
  xor_4  g18343(.A(new_n20675), .B(new_n16068), .Y(new_n20692));
  or_6   g18344(.A(new_n20692), .B(new_n20691), .Y(new_n20693));
  nand_5 g18345(.A(new_n20693), .B(new_n20676), .Y(new_n20694));
  xor_4  g18346(.A(new_n20694), .B(new_n20674), .Y(new_n20695));
  not_8  g18347(.A(new_n20695), .Y(new_n20696));
  xor_4  g18348(.A(pi690), .B(new_n5642), .Y(new_n20697));
  nand_5 g18349(.A(new_n6829), .B(pi575), .Y(new_n20698));
  xor_4  g18350(.A(pi714), .B(new_n3219), .Y(new_n20699));
  nand_5 g18351(.A(new_n18154), .B(new_n18152), .Y(new_n20700));
  nand_5 g18352(.A(new_n20700), .B(new_n18153), .Y(new_n20701));
  nand_5 g18353(.A(new_n20701), .B(new_n20699), .Y(new_n20702));
  nand_5 g18354(.A(new_n20702), .B(new_n20698), .Y(new_n20703));
  xor_4  g18355(.A(new_n20703), .B(new_n20697), .Y(new_n20704));
  not_8  g18356(.A(new_n20704), .Y(new_n20705));
  or_6   g18357(.A(new_n18156), .B(new_n18149), .Y(new_n20706));
  nand_5 g18358(.A(new_n18166), .B(new_n18157), .Y(new_n20707));
  nand_5 g18359(.A(new_n20707), .B(new_n20706), .Y(new_n20708));
  xor_4  g18360(.A(new_n20685), .B(new_n20681), .Y(new_n20709));
  not_8  g18361(.A(new_n20709), .Y(new_n20710));
  or_6   g18362(.A(new_n20710), .B(new_n20708), .Y(new_n20711));
  nand_5 g18363(.A(new_n20710), .B(new_n20708), .Y(new_n20712));
  xnor_4 g18364(.A(new_n20701), .B(new_n20699), .Y(new_n20713));
  nand_5 g18365(.A(new_n20713), .B(new_n20712), .Y(new_n20714));
  nand_5 g18366(.A(new_n20714), .B(new_n20711), .Y(new_n20715));
  nand_5 g18367(.A(new_n20715), .B(new_n20705), .Y(new_n20716));
  xor_4  g18368(.A(new_n20715), .B(new_n20704), .Y(new_n20717));
  xor_4  g18369(.A(new_n20689), .B(new_n20687), .Y(new_n20718));
  or_6   g18370(.A(new_n20718), .B(new_n20717), .Y(new_n20719));
  nand_5 g18371(.A(new_n20719), .B(new_n20716), .Y(new_n20720));
  nand_5 g18372(.A(pi533), .B(new_n3213), .Y(new_n20721));
  nand_5 g18373(.A(new_n10470), .B(pi509), .Y(new_n20722));
  and_6  g18374(.A(new_n20722), .B(new_n20721), .Y(new_n20723));
  nand_5 g18375(.A(pi690), .B(new_n5642), .Y(new_n20724));
  nand_5 g18376(.A(new_n20703), .B(new_n20697), .Y(new_n20725));
  nand_5 g18377(.A(new_n20725), .B(new_n20724), .Y(new_n20726));
  xor_4  g18378(.A(new_n20726), .B(new_n20723), .Y(new_n20727));
  not_8  g18379(.A(new_n20727), .Y(new_n20728));
  nor_5  g18380(.A(new_n20728), .B(new_n20720), .Y(new_n20729));
  xor_4  g18381(.A(new_n20692), .B(new_n20691), .Y(new_n20730));
  xor_4  g18382(.A(new_n20727), .B(new_n20720), .Y(new_n20731));
  not_8  g18383(.A(new_n20731), .Y(new_n20732));
  nand_5 g18384(.A(new_n20732), .B(new_n20730), .Y(new_n20733));
  not_8  g18385(.A(new_n20733), .Y(new_n20734));
  nor_5  g18386(.A(new_n20734), .B(new_n20729), .Y(new_n20735));
  xor_4  g18387(.A(pi735), .B(new_n3208), .Y(new_n20736));
  not_8  g18388(.A(new_n20736), .Y(new_n20737));
  nand_5 g18389(.A(new_n20726), .B(new_n20721), .Y(new_n20738));
  nand_5 g18390(.A(new_n20738), .B(new_n20722), .Y(new_n20739));
  xor_4  g18391(.A(new_n20739), .B(new_n20737), .Y(new_n20740));
  xor_4  g18392(.A(new_n20740), .B(new_n20735), .Y(new_n20741));
  xor_4  g18393(.A(new_n20741), .B(new_n20696), .Y(po0356));
  xor_4  g18394(.A(new_n3649), .B(new_n3648), .Y(po0357));
  xor_4  g18395(.A(new_n16421), .B(new_n8635), .Y(po0358));
  xnor_4 g18396(.A(new_n10025), .B(new_n10002), .Y(po0359));
  not_8  g18397(.A(new_n18388), .Y(new_n20746));
  not_8  g18398(.A(new_n2938), .Y(new_n20747));
  nand_5 g18399(.A(new_n3016), .B(new_n2872), .Y(new_n20748));
  nand_5 g18400(.A(new_n3017), .B(pi144), .Y(new_n20749));
  nand_5 g18401(.A(new_n20749), .B(new_n5780), .Y(new_n20750));
  nand_5 g18402(.A(new_n20750), .B(new_n20748), .Y(new_n20751));
  nor_5  g18403(.A(new_n20751), .B(new_n5246), .Y(new_n20752));
  xor_4  g18404(.A(new_n20751), .B(pi570), .Y(new_n20753));
  nor_5  g18405(.A(new_n20753), .B(new_n3013), .Y(new_n20754));
  or_6   g18406(.A(new_n20754), .B(new_n20752), .Y(new_n20755));
  nand_5 g18407(.A(new_n20755), .B(new_n3008), .Y(new_n20756));
  or_6   g18408(.A(new_n20755), .B(new_n3008), .Y(new_n20757));
  nand_5 g18409(.A(new_n20757), .B(pi151), .Y(new_n20758));
  nand_5 g18410(.A(new_n20758), .B(new_n20756), .Y(new_n20759));
  nand_5 g18411(.A(new_n20759), .B(new_n2999), .Y(new_n20760));
  or_6   g18412(.A(new_n20759), .B(new_n2999), .Y(new_n20761));
  nand_5 g18413(.A(new_n20761), .B(pi172), .Y(new_n20762));
  nand_5 g18414(.A(new_n20762), .B(new_n20760), .Y(new_n20763));
  nand_5 g18415(.A(new_n20763), .B(new_n2993), .Y(new_n20764));
  or_6   g18416(.A(new_n20763), .B(new_n2993), .Y(new_n20765));
  nand_5 g18417(.A(new_n20765), .B(pi061), .Y(new_n20766));
  nand_5 g18418(.A(new_n20766), .B(new_n20764), .Y(new_n20767));
  nand_5 g18419(.A(new_n20767), .B(new_n2988), .Y(new_n20768));
  or_6   g18420(.A(new_n20767), .B(new_n2988), .Y(new_n20769));
  nand_5 g18421(.A(new_n20769), .B(pi410), .Y(new_n20770));
  nand_5 g18422(.A(new_n20770), .B(new_n20768), .Y(new_n20771));
  or_6   g18423(.A(new_n20771), .B(new_n2982), .Y(new_n20772));
  xor_4  g18424(.A(new_n20771), .B(new_n2982), .Y(new_n20773));
  nand_5 g18425(.A(new_n20773), .B(new_n2855), .Y(new_n20774));
  nand_5 g18426(.A(new_n20774), .B(new_n20772), .Y(new_n20775));
  or_6   g18427(.A(new_n20775), .B(new_n20747), .Y(new_n20776));
  nand_5 g18428(.A(new_n20775), .B(new_n20747), .Y(new_n20777));
  nand_5 g18429(.A(new_n20777), .B(pi687), .Y(new_n20778));
  nand_5 g18430(.A(new_n20778), .B(new_n20776), .Y(new_n20779));
  nor_5  g18431(.A(new_n20779), .B(new_n18390), .Y(new_n20780));
  xor_4  g18432(.A(new_n20779), .B(new_n18392), .Y(new_n20781));
  nor_5  g18433(.A(new_n20781), .B(pi358), .Y(new_n20782));
  nor_5  g18434(.A(new_n20782), .B(new_n20780), .Y(new_n20783));
  xor_4  g18435(.A(new_n20783), .B(new_n20746), .Y(new_n20784));
  nor_5  g18436(.A(new_n20784), .B(new_n18042), .Y(new_n20785));
  xor_4  g18437(.A(new_n20784), .B(new_n18042), .Y(new_n20786));
  not_8  g18438(.A(new_n20786), .Y(new_n20787));
  xor_4  g18439(.A(new_n20773), .B(pi047), .Y(new_n20788));
  nand_5 g18440(.A(new_n20788), .B(new_n6063), .Y(new_n20789));
  nand_5 g18441(.A(new_n20757), .B(new_n20756), .Y(new_n20790));
  xor_4  g18442(.A(new_n20790), .B(pi151), .Y(new_n20791));
  xor_4  g18443(.A(new_n20753), .B(new_n3010), .Y(new_n20792));
  or_6   g18444(.A(new_n20792), .B(new_n6016), .Y(new_n20793));
  xor_4  g18445(.A(new_n20792), .B(new_n6016), .Y(new_n20794));
  nand_5 g18446(.A(new_n20748), .B(new_n20749), .Y(new_n20795));
  nand_5 g18447(.A(new_n5780), .B(new_n5779), .Y(new_n20796));
  nand_5 g18448(.A(new_n5781), .B(new_n13084), .Y(new_n20797));
  nand_5 g18449(.A(new_n20797), .B(new_n20796), .Y(new_n20798));
  xor_4  g18450(.A(new_n20798), .B(new_n20795), .Y(new_n20799));
  nor_5  g18451(.A(new_n20799), .B(new_n6020), .Y(new_n20800));
  and_6  g18452(.A(new_n5782), .B(new_n13084), .Y(new_n20801));
  and_6  g18453(.A(new_n20799), .B(new_n20801), .Y(new_n20802));
  nor_5  g18454(.A(new_n20802), .B(new_n20800), .Y(new_n20803));
  nand_5 g18455(.A(new_n20803), .B(new_n20794), .Y(new_n20804));
  nand_5 g18456(.A(new_n20804), .B(new_n20793), .Y(new_n20805));
  not_8  g18457(.A(new_n20805), .Y(new_n20806));
  nor_5  g18458(.A(new_n20806), .B(new_n20791), .Y(new_n20807));
  xor_4  g18459(.A(new_n20805), .B(new_n20791), .Y(new_n20808));
  nor_5  g18460(.A(new_n20808), .B(new_n6014), .Y(new_n20809));
  nor_5  g18461(.A(new_n20809), .B(new_n20807), .Y(new_n20810));
  nand_5 g18462(.A(new_n20761), .B(new_n20760), .Y(new_n20811));
  xor_4  g18463(.A(new_n20811), .B(pi172), .Y(new_n20812));
  nand_5 g18464(.A(new_n20812), .B(new_n20810), .Y(new_n20813));
  xnor_4 g18465(.A(new_n20812), .B(new_n20810), .Y(new_n20814));
  or_6   g18466(.A(new_n20814), .B(new_n6044), .Y(new_n20815));
  nand_5 g18467(.A(new_n20815), .B(new_n20813), .Y(new_n20816));
  nand_5 g18468(.A(new_n20764), .B(new_n20765), .Y(new_n20817));
  xor_4  g18469(.A(new_n20817), .B(pi061), .Y(new_n20818));
  nand_5 g18470(.A(new_n20818), .B(new_n20816), .Y(new_n20819));
  xnor_4 g18471(.A(new_n20818), .B(new_n20816), .Y(new_n20820));
  or_6   g18472(.A(new_n20820), .B(new_n13102), .Y(new_n20821));
  nand_5 g18473(.A(new_n20821), .B(new_n20819), .Y(new_n20822));
  nand_5 g18474(.A(new_n20769), .B(new_n20768), .Y(new_n20823));
  xor_4  g18475(.A(new_n20823), .B(pi410), .Y(new_n20824));
  or_6   g18476(.A(new_n20824), .B(new_n20822), .Y(new_n20825));
  xor_4  g18477(.A(new_n20824), .B(new_n20822), .Y(new_n20826));
  nand_5 g18478(.A(new_n20826), .B(new_n6055), .Y(new_n20827));
  nand_5 g18479(.A(new_n20827), .B(new_n20825), .Y(new_n20828));
  xor_4  g18480(.A(new_n20788), .B(new_n6063), .Y(new_n20829));
  nand_5 g18481(.A(new_n20829), .B(new_n20828), .Y(new_n20830));
  nand_5 g18482(.A(new_n20830), .B(new_n20789), .Y(new_n20831));
  or_6   g18483(.A(new_n20831), .B(new_n6081), .Y(new_n20832));
  nand_5 g18484(.A(new_n20831), .B(new_n6081), .Y(new_n20833));
  nand_5 g18485(.A(new_n20777), .B(new_n20776), .Y(new_n20834));
  xor_4  g18486(.A(new_n20834), .B(pi687), .Y(new_n20835));
  nand_5 g18487(.A(new_n20835), .B(new_n20833), .Y(new_n20836));
  nand_5 g18488(.A(new_n20836), .B(new_n20832), .Y(new_n20837));
  nand_5 g18489(.A(new_n20837), .B(new_n13078), .Y(new_n20838));
  xor_4  g18490(.A(new_n20781), .B(new_n10400), .Y(new_n20839));
  xor_4  g18491(.A(new_n20837), .B(new_n6101), .Y(new_n20840));
  or_6   g18492(.A(new_n20840), .B(new_n20839), .Y(new_n20841));
  nand_5 g18493(.A(new_n20841), .B(new_n20838), .Y(new_n20842));
  nor_5  g18494(.A(new_n20842), .B(new_n20787), .Y(new_n20843));
  nor_5  g18495(.A(new_n20843), .B(new_n20785), .Y(new_n20844));
  nand_5 g18496(.A(new_n20783), .B(new_n18388), .Y(new_n20845));
  xor_4  g18497(.A(new_n20845), .B(new_n18034), .Y(new_n20846));
  xor_4  g18498(.A(new_n20846), .B(new_n20844), .Y(po0360));
  nand_5 g18499(.A(new_n13141), .B(new_n11256), .Y(new_n20848));
  nand_5 g18500(.A(new_n13142), .B(new_n4232), .Y(new_n20849));
  nand_5 g18501(.A(new_n20849), .B(new_n20848), .Y(new_n20850));
  nor_5  g18502(.A(new_n20850), .B(new_n15018), .Y(new_n20851));
  xor_4  g18503(.A(new_n20850), .B(new_n15017), .Y(new_n20852));
  nor_5  g18504(.A(new_n20852), .B(new_n11261), .Y(new_n20853));
  nor_5  g18505(.A(new_n20853), .B(new_n20851), .Y(new_n20854));
  xor_4  g18506(.A(new_n20854), .B(new_n15044), .Y(new_n20855));
  xor_4  g18507(.A(new_n20855), .B(new_n11266), .Y(po0361));
  nor_5  g18508(.A(pi773), .B(new_n11393), .Y(new_n20857));
  nand_5 g18509(.A(new_n11407), .B(new_n11394), .Y(new_n20858));
  not_8  g18510(.A(new_n20858), .Y(new_n20859));
  nor_5  g18511(.A(new_n20859), .B(new_n20857), .Y(new_n20860));
  not_8  g18512(.A(new_n20860), .Y(new_n20861));
  nand_5 g18513(.A(new_n20861), .B(new_n18558), .Y(new_n20862));
  xor_4  g18514(.A(new_n20860), .B(new_n18559), .Y(new_n20863));
  or_6   g18515(.A(new_n11408), .B(new_n11392), .Y(new_n20864));
  nand_5 g18516(.A(new_n11431), .B(new_n11409), .Y(new_n20865));
  nand_5 g18517(.A(new_n20865), .B(new_n20864), .Y(new_n20866));
  nand_5 g18518(.A(new_n20866), .B(new_n20863), .Y(new_n20867));
  nand_5 g18519(.A(new_n20867), .B(new_n20862), .Y(new_n20868));
  nor_5  g18520(.A(new_n16040), .B(new_n16020), .Y(new_n20869));
  nor_5  g18521(.A(new_n16042), .B(new_n11432), .Y(new_n20870));
  or_6   g18522(.A(new_n20870), .B(new_n20869), .Y(new_n20871));
  xor_4  g18523(.A(new_n20866), .B(new_n20863), .Y(new_n20872));
  nand_5 g18524(.A(new_n13031), .B(pi272), .Y(new_n20873));
  nand_5 g18525(.A(new_n16019), .B(new_n16005), .Y(new_n20874));
  nand_5 g18526(.A(new_n20874), .B(new_n20873), .Y(new_n20875));
  nand_5 g18527(.A(new_n20875), .B(new_n20872), .Y(new_n20876));
  nor_5  g18528(.A(new_n20876), .B(new_n20871), .Y(new_n20877));
  nor_5  g18529(.A(new_n20877), .B(new_n20868), .Y(new_n20878));
  nor_5  g18530(.A(new_n20875), .B(new_n20872), .Y(new_n20879));
  nand_5 g18531(.A(new_n20879), .B(new_n20871), .Y(new_n20880));
  and_6  g18532(.A(new_n20880), .B(new_n20868), .Y(new_n20881));
  nor_5  g18533(.A(new_n20881), .B(new_n20878), .Y(po0362));
  nand_5 g18534(.A(new_n6083), .B(new_n6082), .Y(new_n20883));
  xor_4  g18535(.A(new_n20883), .B(new_n6084), .Y(po0363));
  nand_5 g18536(.A(new_n17949), .B(new_n17948), .Y(new_n20885));
  xor_4  g18537(.A(new_n20885), .B(new_n7914), .Y(po0364));
  xor_4  g18538(.A(new_n7467), .B(new_n7465), .Y(po0365));
  xor_4  g18539(.A(new_n14614), .B(new_n14563), .Y(po0366));
  xnor_4 g18540(.A(new_n20090), .B(new_n20089), .Y(po0367));
  nand_5 g18541(.A(new_n15098), .B(new_n11228), .Y(new_n20890));
  nand_5 g18542(.A(new_n15097), .B(new_n11227), .Y(new_n20891));
  nand_5 g18543(.A(new_n20891), .B(new_n20890), .Y(new_n20892));
  nand_5 g18544(.A(new_n20854), .B(new_n15045), .Y(new_n20893));
  or_6   g18545(.A(new_n20855), .B(new_n11266), .Y(new_n20894));
  nand_5 g18546(.A(new_n20894), .B(new_n20893), .Y(new_n20895));
  or_6   g18547(.A(new_n20895), .B(new_n11231), .Y(new_n20896));
  xor_4  g18548(.A(new_n20895), .B(new_n11231), .Y(new_n20897));
  nand_5 g18549(.A(new_n20897), .B(new_n15016), .Y(new_n20898));
  nand_5 g18550(.A(new_n20898), .B(new_n20896), .Y(new_n20899));
  nand_5 g18551(.A(new_n20899), .B(new_n15015), .Y(new_n20900));
  xor_4  g18552(.A(new_n20899), .B(new_n15015), .Y(new_n20901));
  nand_5 g18553(.A(new_n20901), .B(new_n11275), .Y(new_n20902));
  nand_5 g18554(.A(new_n20902), .B(new_n20900), .Y(new_n20903));
  nand_5 g18555(.A(new_n20903), .B(new_n15014), .Y(new_n20904));
  not_8  g18556(.A(new_n11283), .Y(new_n20905));
  xor_4  g18557(.A(new_n20903), .B(new_n15014), .Y(new_n20906));
  nand_5 g18558(.A(new_n20906), .B(new_n20905), .Y(new_n20907));
  nand_5 g18559(.A(new_n20907), .B(new_n20904), .Y(new_n20908));
  xor_4  g18560(.A(new_n20908), .B(new_n20892), .Y(po0368));
  xor_4  g18561(.A(new_n14909), .B(new_n14908), .Y(po0369));
  xor_4  g18562(.A(new_n11204), .B(new_n8928), .Y(po0370));
  xor_4  g18563(.A(new_n19978), .B(new_n17216), .Y(po0371));
  xor_4  g18564(.A(new_n17774), .B(new_n12252), .Y(po0372));
  xnor_4 g18565(.A(new_n7433), .B(new_n7425), .Y(po0373));
  xor_4  g18566(.A(new_n15972), .B(new_n15960), .Y(po0374));
  xor_4  g18567(.A(new_n8623), .B(new_n8608), .Y(po0375));
  xor_4  g18568(.A(new_n19207), .B(new_n15207), .Y(po0376));
  nand_5 g18569(.A(new_n13359), .B(new_n13357), .Y(new_n20918));
  xnor_4 g18570(.A(new_n20918), .B(new_n13354), .Y(po0377));
  xor_4  g18571(.A(new_n16292), .B(new_n6904), .Y(po0378));
  nand_5 g18572(.A(new_n11091), .B(pi397), .Y(new_n20921));
  not_8  g18573(.A(new_n20921), .Y(new_n20922));
  not_8  g18574(.A(new_n19596), .Y(new_n20923));
  nor_5  g18575(.A(new_n19601), .B(new_n20923), .Y(new_n20924));
  nor_5  g18576(.A(new_n20924), .B(new_n20922), .Y(new_n20925));
  nand_5 g18577(.A(new_n20925), .B(new_n14271), .Y(new_n20926));
  not_8  g18578(.A(new_n20925), .Y(new_n20927));
  xor_4  g18579(.A(new_n20927), .B(new_n14270), .Y(new_n20928));
  nand_5 g18580(.A(new_n20928), .B(new_n10404), .Y(new_n20929));
  nand_5 g18581(.A(new_n20929), .B(new_n20926), .Y(new_n20930));
  nand_5 g18582(.A(new_n19602), .B(new_n10278), .Y(new_n20931));
  xor_4  g18583(.A(new_n19603), .B(new_n10278), .Y(new_n20932));
  or_6   g18584(.A(new_n20932), .B(new_n14273), .Y(new_n20933));
  nand_5 g18585(.A(new_n20933), .B(new_n20931), .Y(new_n20934));
  xor_4  g18586(.A(new_n20928), .B(new_n10403), .Y(new_n20935));
  or_6   g18587(.A(new_n20935), .B(new_n20934), .Y(new_n20936));
  xor_4  g18588(.A(new_n20932), .B(new_n14273), .Y(new_n20937));
  nor_5  g18589(.A(new_n14279), .B(new_n10319), .Y(new_n20938));
  nand_5 g18590(.A(new_n20130), .B(new_n20128), .Y(new_n20939));
  not_8  g18591(.A(new_n20939), .Y(new_n20940));
  nor_5  g18592(.A(new_n20940), .B(new_n20938), .Y(new_n20941));
  nor_5  g18593(.A(new_n20941), .B(new_n20937), .Y(new_n20942));
  nand_5 g18594(.A(new_n20124), .B(new_n16877), .Y(new_n20943));
  or_6   g18595(.A(new_n20131), .B(new_n20125), .Y(new_n20944));
  nand_5 g18596(.A(new_n20944), .B(new_n20943), .Y(new_n20945));
  and_6  g18597(.A(new_n20941), .B(new_n20937), .Y(new_n20946));
  nor_5  g18598(.A(new_n20946), .B(new_n20945), .Y(new_n20947));
  or_6   g18599(.A(new_n20947), .B(new_n20942), .Y(new_n20948));
  nand_5 g18600(.A(new_n20935), .B(new_n20934), .Y(new_n20949));
  nand_5 g18601(.A(new_n20949), .B(new_n20948), .Y(new_n20950));
  nand_5 g18602(.A(new_n20950), .B(new_n20936), .Y(new_n20951));
  xnor_4 g18603(.A(new_n20951), .B(new_n20930), .Y(po0379));
  not_8  g18604(.A(new_n19804), .Y(new_n20953));
  or_6   g18605(.A(new_n19709), .B(new_n19705), .Y(new_n20954));
  nand_5 g18606(.A(new_n19725), .B(new_n19710), .Y(new_n20955));
  nand_5 g18607(.A(new_n20955), .B(new_n20954), .Y(new_n20956));
  nor_5  g18608(.A(new_n19703), .B(new_n15684), .Y(new_n20957));
  nor_5  g18609(.A(new_n19704), .B(new_n19699), .Y(new_n20958));
  nor_5  g18610(.A(new_n20958), .B(new_n20957), .Y(new_n20959));
  not_8  g18611(.A(new_n15730), .Y(new_n20960));
  nand_5 g18612(.A(new_n19702), .B(new_n10093), .Y(new_n20961));
  nand_5 g18613(.A(new_n20961), .B(new_n10094), .Y(new_n20962));
  nand_5 g18614(.A(new_n20962), .B(new_n20960), .Y(new_n20963));
  nor_5  g18615(.A(new_n20962), .B(new_n20960), .Y(new_n20964));
  not_8  g18616(.A(new_n20964), .Y(new_n20965));
  nand_5 g18617(.A(new_n20965), .B(new_n20963), .Y(new_n20966));
  xor_4  g18618(.A(new_n20966), .B(new_n10141), .Y(new_n20967));
  xor_4  g18619(.A(new_n20967), .B(new_n20959), .Y(new_n20968));
  nor_5  g18620(.A(new_n20968), .B(new_n20956), .Y(new_n20969));
  not_8  g18621(.A(new_n20968), .Y(new_n20970));
  xor_4  g18622(.A(new_n20970), .B(new_n20956), .Y(new_n20971));
  nor_5  g18623(.A(new_n20971), .B(new_n19816), .Y(new_n20972));
  or_6   g18624(.A(new_n20972), .B(new_n20969), .Y(new_n20973));
  xor_4  g18625(.A(new_n20973), .B(new_n20953), .Y(new_n20974));
  nand_5 g18626(.A(new_n8052), .B(pi079), .Y(new_n20975));
  nand_5 g18627(.A(new_n20975), .B(new_n20959), .Y(new_n20976));
  nand_5 g18628(.A(pi700), .B(new_n10138), .Y(new_n20977));
  not_8  g18629(.A(new_n20977), .Y(new_n20978));
  nor_5  g18630(.A(new_n20978), .B(new_n20963), .Y(new_n20979));
  nand_5 g18631(.A(new_n20979), .B(new_n20976), .Y(new_n20980));
  or_6   g18632(.A(new_n20975), .B(new_n20964), .Y(new_n20981));
  or_6   g18633(.A(new_n20981), .B(new_n20959), .Y(new_n20982));
  nand_5 g18634(.A(new_n20982), .B(new_n20980), .Y(new_n20983));
  nand_5 g18635(.A(new_n20983), .B(new_n15736), .Y(new_n20984));
  not_8  g18636(.A(new_n15736), .Y(new_n20985));
  nand_5 g18637(.A(new_n20978), .B(new_n20964), .Y(new_n20986));
  nand_5 g18638(.A(new_n20977), .B(new_n20965), .Y(new_n20987));
  nand_5 g18639(.A(new_n20987), .B(new_n20963), .Y(new_n20988));
  or_6   g18640(.A(new_n20988), .B(new_n20976), .Y(new_n20989));
  nand_5 g18641(.A(new_n20989), .B(new_n20986), .Y(new_n20990));
  nand_5 g18642(.A(new_n20990), .B(new_n20985), .Y(new_n20991));
  nor_5  g18643(.A(new_n20990), .B(new_n20985), .Y(new_n20992));
  nor_5  g18644(.A(new_n20992), .B(new_n20983), .Y(new_n20993));
  nand_5 g18645(.A(new_n20993), .B(new_n20991), .Y(new_n20994));
  nand_5 g18646(.A(new_n20994), .B(new_n20984), .Y(new_n20995));
  xor_4  g18647(.A(new_n20995), .B(new_n20974), .Y(po0380));
  nand_5 g18648(.A(new_n11025), .B(new_n11077), .Y(new_n20997));
  xor_4  g18649(.A(new_n20997), .B(pi069), .Y(new_n20998));
  nand_5 g18650(.A(new_n11072), .B(new_n11077), .Y(new_n20999));
  not_8  g18651(.A(pi320), .Y(new_n21000));
  nand_5 g18652(.A(new_n10999), .B(new_n21000), .Y(new_n21001));
  xor_4  g18653(.A(new_n10999), .B(new_n21000), .Y(new_n21002));
  not_8  g18654(.A(pi042), .Y(new_n21003));
  nand_5 g18655(.A(new_n7245), .B(new_n10996), .Y(new_n21004));
  nand_5 g18656(.A(new_n21004), .B(pi366), .Y(new_n21005));
  nor_5  g18657(.A(new_n21005), .B(new_n9650), .Y(new_n21006));
  or_6   g18658(.A(new_n21004), .B(pi366), .Y(new_n21007));
  nor_5  g18659(.A(new_n21007), .B(pi255), .Y(new_n21008));
  or_6   g18660(.A(new_n21008), .B(new_n21006), .Y(new_n21009));
  xor_4  g18661(.A(pi658), .B(new_n10995), .Y(new_n21010));
  xor_4  g18662(.A(new_n21010), .B(new_n21009), .Y(new_n21011));
  nor_5  g18663(.A(pi658), .B(pi169), .Y(new_n21012));
  nor_5  g18664(.A(new_n21012), .B(new_n21008), .Y(new_n21013));
  nand_5 g18665(.A(new_n21013), .B(new_n21011), .Y(new_n21014));
  nand_5 g18666(.A(new_n21010), .B(new_n21009), .Y(new_n21015));
  nor_5  g18667(.A(new_n9648), .B(pi366), .Y(new_n21016));
  nor_5  g18668(.A(new_n21016), .B(new_n21015), .Y(new_n21017));
  nor_5  g18669(.A(new_n21017), .B(pi651), .Y(new_n21018));
  nand_5 g18670(.A(new_n21018), .B(new_n21014), .Y(new_n21019));
  not_8  g18671(.A(new_n21011), .Y(new_n21020));
  nand_5 g18672(.A(new_n21020), .B(new_n9648), .Y(new_n21021));
  nand_5 g18673(.A(new_n10992), .B(new_n10995), .Y(new_n21022));
  nand_5 g18674(.A(new_n21022), .B(pi651), .Y(new_n21023));
  nand_5 g18675(.A(new_n21023), .B(new_n10994), .Y(new_n21024));
  or_6   g18676(.A(new_n21024), .B(new_n21021), .Y(new_n21025));
  nand_5 g18677(.A(new_n21025), .B(new_n21019), .Y(new_n21026));
  nand_5 g18678(.A(pi366), .B(pi169), .Y(new_n21027));
  nor_5  g18679(.A(new_n21027), .B(new_n10993), .Y(new_n21028));
  nand_5 g18680(.A(new_n21028), .B(new_n21021), .Y(new_n21029));
  nor_5  g18681(.A(new_n21023), .B(new_n9648), .Y(new_n21030));
  nand_5 g18682(.A(new_n21030), .B(new_n21011), .Y(new_n21031));
  nand_5 g18683(.A(new_n21031), .B(new_n21029), .Y(new_n21032));
  nor_5  g18684(.A(new_n21032), .B(new_n21026), .Y(new_n21033));
  nand_5 g18685(.A(new_n21033), .B(new_n21003), .Y(new_n21034));
  nand_5 g18686(.A(new_n21026), .B(new_n11015), .Y(new_n21035));
  nand_5 g18687(.A(new_n21035), .B(new_n21034), .Y(new_n21036));
  nand_5 g18688(.A(new_n21036), .B(new_n21002), .Y(new_n21037));
  nand_5 g18689(.A(new_n21037), .B(new_n21001), .Y(new_n21038));
  nand_5 g18690(.A(new_n21038), .B(new_n10986), .Y(new_n21039));
  nand_5 g18691(.A(new_n21039), .B(new_n11026), .Y(new_n21040));
  nand_5 g18692(.A(new_n11024), .B(pi643), .Y(new_n21041));
  or_6   g18693(.A(new_n21041), .B(new_n21038), .Y(new_n21042));
  nand_5 g18694(.A(new_n21042), .B(new_n21040), .Y(new_n21043));
  nand_5 g18695(.A(new_n21043), .B(new_n20999), .Y(new_n21044));
  nor_5  g18696(.A(new_n21039), .B(new_n11024), .Y(new_n21045));
  nand_5 g18697(.A(pi627), .B(pi015), .Y(new_n21046));
  nor_5  g18698(.A(new_n21046), .B(new_n21045), .Y(new_n21047));
  not_8  g18699(.A(new_n21045), .Y(new_n21048));
  nor_5  g18700(.A(new_n21048), .B(new_n20999), .Y(new_n21049));
  nor_5  g18701(.A(new_n21049), .B(new_n21047), .Y(new_n21050));
  nand_5 g18702(.A(new_n21050), .B(new_n21044), .Y(new_n21051));
  xor_4  g18703(.A(new_n21051), .B(pi069), .Y(new_n21052));
  not_8  g18704(.A(new_n21052), .Y(new_n21053));
  nand_5 g18705(.A(new_n21053), .B(new_n20998), .Y(new_n21054));
  nand_5 g18706(.A(new_n21052), .B(new_n11511), .Y(new_n21055));
  nand_5 g18707(.A(new_n21055), .B(new_n21054), .Y(new_n21056));
  nand_5 g18708(.A(new_n21056), .B(new_n11506), .Y(new_n21057));
  not_8  g18709(.A(pi736), .Y(new_n21058));
  or_6   g18710(.A(new_n20997), .B(pi069), .Y(new_n21059));
  nor_5  g18711(.A(new_n21059), .B(pi415), .Y(new_n21060));
  nand_5 g18712(.A(new_n21060), .B(new_n21058), .Y(new_n21061));
  not_8  g18713(.A(new_n21061), .Y(new_n21062));
  nand_5 g18714(.A(new_n21062), .B(new_n11500), .Y(new_n21063));
  nor_5  g18715(.A(new_n21063), .B(new_n21057), .Y(new_n21064));
  xor_4  g18716(.A(new_n21059), .B(pi415), .Y(new_n21065));
  or_6   g18717(.A(new_n21065), .B(new_n21056), .Y(new_n21066));
  nand_5 g18718(.A(new_n21065), .B(new_n21056), .Y(new_n21067));
  nand_5 g18719(.A(new_n21067), .B(pi561), .Y(new_n21068));
  nand_5 g18720(.A(new_n21068), .B(new_n21066), .Y(new_n21069));
  or_6   g18721(.A(new_n21060), .B(new_n21058), .Y(new_n21070));
  nand_5 g18722(.A(new_n21070), .B(new_n21061), .Y(new_n21071));
  xor_4  g18723(.A(new_n21071), .B(new_n11500), .Y(new_n21072));
  xor_4  g18724(.A(new_n21072), .B(new_n21069), .Y(new_n21073));
  nand_5 g18725(.A(new_n21058), .B(new_n11500), .Y(new_n21074));
  and_6  g18726(.A(new_n21074), .B(new_n21057), .Y(new_n21075));
  nand_5 g18727(.A(new_n21075), .B(new_n21073), .Y(new_n21076));
  nor_5  g18728(.A(new_n21070), .B(new_n11500), .Y(new_n21077));
  nor_5  g18729(.A(new_n21077), .B(new_n21064), .Y(new_n21078));
  nand_5 g18730(.A(new_n21078), .B(new_n21076), .Y(new_n21079));
  nand_5 g18731(.A(new_n21079), .B(new_n15959), .Y(new_n21080));
  not_8  g18732(.A(pi321), .Y(new_n21081));
  nor_5  g18733(.A(new_n14861), .B(new_n21081), .Y(new_n21082));
  xor_4  g18734(.A(new_n2669), .B(pi321), .Y(new_n21083));
  not_8  g18735(.A(new_n21083), .Y(new_n21084));
  nor_5  g18736(.A(new_n21084), .B(new_n21073), .Y(new_n21085));
  nor_5  g18737(.A(new_n21085), .B(new_n21082), .Y(new_n21086));
  xor_4  g18738(.A(pi561), .B(pi194), .Y(new_n21087));
  nand_5 g18739(.A(new_n21066), .B(new_n21067), .Y(new_n21088));
  xor_4  g18740(.A(new_n21088), .B(new_n21087), .Y(new_n21089));
  not_8  g18741(.A(new_n21089), .Y(new_n21090));
  nor_5  g18742(.A(new_n21090), .B(pi194), .Y(new_n21091));
  xor_4  g18743(.A(new_n21052), .B(pi199), .Y(new_n21092));
  nand_5 g18744(.A(new_n21020), .B(pi595), .Y(new_n21093));
  xor_4  g18745(.A(new_n21011), .B(pi595), .Y(new_n21094));
  xor_4  g18746(.A(pi642), .B(pi481), .Y(new_n21095));
  not_8  g18747(.A(new_n21095), .Y(new_n21096));
  nand_5 g18748(.A(new_n21096), .B(pi477), .Y(new_n21097));
  not_8  g18749(.A(new_n21097), .Y(new_n21098));
  nand_5 g18750(.A(new_n21007), .B(new_n21005), .Y(new_n21099));
  xor_4  g18751(.A(new_n21099), .B(new_n16616), .Y(new_n21100));
  nand_5 g18752(.A(new_n21100), .B(new_n21098), .Y(new_n21101));
  not_8  g18753(.A(new_n21100), .Y(new_n21102));
  nand_5 g18754(.A(new_n21102), .B(pi163), .Y(new_n21103));
  nand_5 g18755(.A(new_n21103), .B(new_n21101), .Y(new_n21104));
  not_8  g18756(.A(new_n21104), .Y(new_n21105));
  or_6   g18757(.A(new_n21105), .B(new_n21094), .Y(new_n21106));
  nand_5 g18758(.A(new_n21106), .B(new_n21093), .Y(new_n21107));
  nand_5 g18759(.A(new_n21107), .B(pi746), .Y(new_n21108));
  xor_4  g18760(.A(new_n21033), .B(new_n21003), .Y(new_n21109));
  xnor_4 g18761(.A(new_n21107), .B(pi746), .Y(new_n21110));
  or_6   g18762(.A(new_n21110), .B(new_n21109), .Y(new_n21111));
  nand_5 g18763(.A(new_n21111), .B(new_n21108), .Y(new_n21112));
  nand_5 g18764(.A(new_n21112), .B(pi269), .Y(new_n21113));
  xor_4  g18765(.A(new_n21036), .B(new_n21002), .Y(new_n21114));
  not_8  g18766(.A(pi269), .Y(new_n21115));
  xor_4  g18767(.A(new_n21112), .B(new_n21115), .Y(new_n21116));
  or_6   g18768(.A(new_n21116), .B(new_n21114), .Y(new_n21117));
  nand_5 g18769(.A(new_n21117), .B(new_n21113), .Y(new_n21118));
  xor_4  g18770(.A(new_n11027), .B(pi643), .Y(new_n21119));
  xor_4  g18771(.A(new_n21119), .B(new_n21038), .Y(new_n21120));
  nand_5 g18772(.A(new_n21120), .B(new_n21118), .Y(new_n21121));
  xor_4  g18773(.A(new_n21120), .B(new_n21118), .Y(new_n21122));
  nand_5 g18774(.A(new_n21122), .B(pi538), .Y(new_n21123));
  nand_5 g18775(.A(new_n21123), .B(new_n21121), .Y(new_n21124));
  nand_5 g18776(.A(new_n11027), .B(new_n10986), .Y(new_n21125));
  not_8  g18777(.A(new_n21119), .Y(new_n21126));
  nand_5 g18778(.A(new_n21126), .B(new_n21038), .Y(new_n21127));
  nand_5 g18779(.A(new_n21127), .B(new_n21125), .Y(new_n21128));
  xor_4  g18780(.A(new_n11078), .B(new_n11072), .Y(new_n21129));
  xor_4  g18781(.A(new_n21129), .B(new_n21128), .Y(new_n21130));
  nand_5 g18782(.A(new_n21130), .B(new_n21124), .Y(new_n21131));
  xor_4  g18783(.A(new_n21130), .B(new_n21124), .Y(new_n21132));
  nand_5 g18784(.A(new_n21132), .B(pi063), .Y(new_n21133));
  nand_5 g18785(.A(new_n21133), .B(new_n21131), .Y(new_n21134));
  or_6   g18786(.A(new_n21134), .B(new_n21092), .Y(new_n21135));
  nand_5 g18787(.A(new_n21135), .B(pi202), .Y(new_n21136));
  nand_5 g18788(.A(new_n21134), .B(new_n21092), .Y(new_n21137));
  nand_5 g18789(.A(new_n21137), .B(new_n21136), .Y(new_n21138));
  nor_5  g18790(.A(new_n21138), .B(new_n21089), .Y(new_n21139));
  nor_5  g18791(.A(new_n21139), .B(new_n21091), .Y(new_n21140));
  not_8  g18792(.A(new_n21140), .Y(new_n21141));
  xor_4  g18793(.A(new_n21138), .B(new_n21090), .Y(new_n21142));
  nor_5  g18794(.A(new_n21142), .B(new_n2670), .Y(new_n21143));
  xor_4  g18795(.A(new_n21142), .B(new_n2826), .Y(new_n21144));
  xnor_4 g18796(.A(new_n21132), .B(pi063), .Y(new_n21145));
  nor_5  g18797(.A(new_n21145), .B(new_n2801), .Y(new_n21146));
  xor_4  g18798(.A(new_n21145), .B(new_n2797), .Y(new_n21147));
  xor_4  g18799(.A(new_n21104), .B(new_n21094), .Y(new_n21148));
  nand_5 g18800(.A(new_n21148), .B(new_n2765), .Y(new_n21149));
  nand_5 g18801(.A(new_n21100), .B(new_n2744), .Y(new_n21150));
  or_6   g18802(.A(new_n21096), .B(pi477), .Y(new_n21151));
  nor_5  g18803(.A(new_n21151), .B(new_n2754), .Y(new_n21152));
  nor_5  g18804(.A(new_n21097), .B(new_n2755), .Y(new_n21153));
  or_6   g18805(.A(new_n21153), .B(new_n21152), .Y(new_n21154));
  xor_4  g18806(.A(new_n21100), .B(new_n2744), .Y(new_n21155));
  nor_5  g18807(.A(new_n21155), .B(new_n21154), .Y(new_n21156));
  or_6   g18808(.A(new_n21156), .B(new_n21152), .Y(new_n21157));
  nand_5 g18809(.A(new_n21157), .B(new_n21150), .Y(new_n21158));
  not_8  g18810(.A(new_n21101), .Y(new_n21159));
  nand_5 g18811(.A(new_n21159), .B(new_n14883), .Y(new_n21160));
  nand_5 g18812(.A(new_n21160), .B(new_n21158), .Y(new_n21161));
  or_6   g18813(.A(new_n21148), .B(new_n2765), .Y(new_n21162));
  nand_5 g18814(.A(new_n21162), .B(new_n21161), .Y(new_n21163));
  nand_5 g18815(.A(new_n21163), .B(new_n21149), .Y(new_n21164));
  nand_5 g18816(.A(new_n21164), .B(new_n2770), .Y(new_n21165));
  xor_4  g18817(.A(new_n21164), .B(new_n2770), .Y(new_n21166));
  not_8  g18818(.A(new_n21166), .Y(new_n21167));
  xor_4  g18819(.A(new_n21110), .B(new_n21109), .Y(new_n21168));
  or_6   g18820(.A(new_n21168), .B(new_n21167), .Y(new_n21169));
  nand_5 g18821(.A(new_n21169), .B(new_n21165), .Y(new_n21170));
  nor_5  g18822(.A(new_n21170), .B(new_n14876), .Y(new_n21171));
  xnor_4 g18823(.A(new_n21116), .B(new_n21114), .Y(new_n21172));
  xor_4  g18824(.A(new_n21170), .B(new_n2779), .Y(new_n21173));
  nor_5  g18825(.A(new_n21173), .B(new_n21172), .Y(new_n21174));
  or_6   g18826(.A(new_n21174), .B(new_n21171), .Y(new_n21175));
  xor_4  g18827(.A(new_n21122), .B(pi538), .Y(new_n21176));
  or_6   g18828(.A(new_n21176), .B(new_n21175), .Y(new_n21177));
  xor_4  g18829(.A(new_n21176), .B(new_n21175), .Y(new_n21178));
  nand_5 g18830(.A(new_n21178), .B(new_n2789), .Y(new_n21179));
  nand_5 g18831(.A(new_n21179), .B(new_n21177), .Y(new_n21180));
  nor_5  g18832(.A(new_n21180), .B(new_n21147), .Y(new_n21181));
  or_6   g18833(.A(new_n21181), .B(new_n21146), .Y(new_n21182));
  not_8  g18834(.A(pi202), .Y(new_n21183));
  nand_5 g18835(.A(new_n21137), .B(new_n21135), .Y(new_n21184));
  xor_4  g18836(.A(new_n21184), .B(new_n21183), .Y(new_n21185));
  nand_5 g18837(.A(new_n21185), .B(new_n21182), .Y(new_n21186));
  or_6   g18838(.A(new_n21185), .B(new_n21182), .Y(new_n21187));
  nand_5 g18839(.A(new_n21187), .B(new_n2741), .Y(new_n21188));
  nand_5 g18840(.A(new_n21188), .B(new_n21186), .Y(new_n21189));
  nor_5  g18841(.A(new_n21189), .B(new_n21144), .Y(new_n21190));
  or_6   g18842(.A(new_n21190), .B(new_n21143), .Y(new_n21191));
  nand_5 g18843(.A(new_n21191), .B(new_n21141), .Y(new_n21192));
  xor_4  g18844(.A(new_n21084), .B(new_n21073), .Y(new_n21193));
  xor_4  g18845(.A(new_n21191), .B(new_n21140), .Y(new_n21194));
  or_6   g18846(.A(new_n21194), .B(new_n21193), .Y(new_n21195));
  nand_5 g18847(.A(new_n21195), .B(new_n21192), .Y(new_n21196));
  nor_5  g18848(.A(new_n21196), .B(new_n21086), .Y(new_n21197));
  nand_5 g18849(.A(new_n21197), .B(new_n21080), .Y(new_n21198));
  or_6   g18850(.A(new_n21079), .B(new_n15959), .Y(new_n21199));
  nand_5 g18851(.A(new_n21199), .B(new_n21080), .Y(new_n21200));
  nand_5 g18852(.A(new_n21196), .B(new_n21086), .Y(new_n21201));
  nor_5  g18853(.A(new_n21201), .B(new_n21200), .Y(new_n21202));
  not_8  g18854(.A(new_n21197), .Y(new_n21203));
  nand_5 g18855(.A(new_n21199), .B(new_n21203), .Y(new_n21204));
  or_6   g18856(.A(new_n21204), .B(new_n21202), .Y(new_n21205));
  nand_5 g18857(.A(new_n21205), .B(new_n21198), .Y(new_n21206));
  xor_4  g18858(.A(new_n21206), .B(new_n21064), .Y(new_n21207));
  xor_4  g18859(.A(new_n21207), .B(new_n14816), .Y(po0381));
  xor_4  g18860(.A(new_n13523), .B(new_n9688), .Y(po0382));
  xor_4  g18861(.A(new_n5718), .B(new_n5717), .Y(po0383));
  xor_4  g18862(.A(new_n19577), .B(new_n19565), .Y(po0384));
  nand_5 g18863(.A(new_n19811), .B(new_n7377), .Y(new_n21212));
  nor_5  g18864(.A(new_n15157), .B(new_n15130), .Y(new_n21213));
  nor_5  g18865(.A(new_n15158), .B(new_n7312), .Y(new_n21214));
  or_6   g18866(.A(new_n21214), .B(new_n21213), .Y(new_n21215));
  nand_5 g18867(.A(new_n21215), .B(new_n19817), .Y(new_n21216));
  xor_4  g18868(.A(new_n21215), .B(new_n19814), .Y(new_n21217));
  or_6   g18869(.A(new_n21217), .B(new_n7293), .Y(new_n21218));
  nand_5 g18870(.A(new_n21218), .B(new_n21216), .Y(new_n21219));
  or_6   g18871(.A(new_n21219), .B(new_n21212), .Y(new_n21220));
  nand_5 g18872(.A(new_n21219), .B(new_n21212), .Y(new_n21221));
  nor_5  g18873(.A(new_n19811), .B(new_n7377), .Y(new_n21222));
  not_8  g18874(.A(new_n21222), .Y(new_n21223));
  nand_5 g18875(.A(new_n21223), .B(new_n21221), .Y(new_n21224));
  nand_5 g18876(.A(new_n21222), .B(new_n21219), .Y(new_n21225));
  nand_5 g18877(.A(new_n21225), .B(new_n21224), .Y(new_n21226));
  nand_5 g18878(.A(new_n21226), .B(new_n21220), .Y(new_n21227));
  or_6   g18879(.A(new_n19219), .B(new_n19190), .Y(new_n21228));
  nand_5 g18880(.A(new_n19220), .B(new_n15159), .Y(new_n21229));
  nand_5 g18881(.A(new_n21229), .B(new_n21228), .Y(new_n21230));
  xor_4  g18882(.A(new_n21217), .B(new_n7293), .Y(new_n21231));
  not_8  g18883(.A(new_n21231), .Y(new_n21232));
  nand_5 g18884(.A(new_n21232), .B(new_n21230), .Y(new_n21233));
  xor_4  g18885(.A(new_n19835), .B(new_n19832), .Y(new_n21234));
  xor_4  g18886(.A(new_n21232), .B(new_n21230), .Y(new_n21235));
  nand_5 g18887(.A(new_n21235), .B(new_n21234), .Y(new_n21236));
  nand_5 g18888(.A(new_n21236), .B(new_n21233), .Y(new_n21237));
  xor_4  g18889(.A(new_n21237), .B(new_n21227), .Y(new_n21238));
  xor_4  g18890(.A(new_n21238), .B(new_n19837), .Y(po0385));
  xnor_4 g18891(.A(new_n3665), .B(new_n3664), .Y(po0386));
  nand_5 g18892(.A(new_n14202), .B(new_n14191), .Y(new_n21241));
  nand_5 g18893(.A(new_n14205), .B(new_n14209), .Y(new_n21242));
  nand_5 g18894(.A(new_n21242), .B(new_n21241), .Y(new_n21243));
  xor_4  g18895(.A(new_n21243), .B(new_n20861), .Y(new_n21244));
  not_8  g18896(.A(new_n21244), .Y(new_n21245));
  xor_4  g18897(.A(new_n14207), .B(new_n14191), .Y(new_n21246));
  nand_5 g18898(.A(new_n21246), .B(new_n20860), .Y(new_n21247));
  xor_4  g18899(.A(new_n21246), .B(new_n20861), .Y(new_n21248));
  nand_5 g18900(.A(new_n14155), .B(new_n11412), .Y(new_n21249));
  nand_5 g18901(.A(new_n14156), .B(new_n11411), .Y(new_n21250));
  nand_5 g18902(.A(new_n6565), .B(new_n6545), .Y(new_n21251));
  nand_5 g18903(.A(new_n6566), .B(new_n6539), .Y(new_n21252));
  nand_5 g18904(.A(new_n21252), .B(new_n21251), .Y(new_n21253));
  nand_5 g18905(.A(new_n21253), .B(new_n14117), .Y(new_n21254));
  xor_4  g18906(.A(new_n21253), .B(new_n14117), .Y(new_n21255));
  not_8  g18907(.A(new_n21255), .Y(new_n21256));
  or_6   g18908(.A(new_n21256), .B(new_n11416), .Y(new_n21257));
  nand_5 g18909(.A(new_n21257), .B(new_n21254), .Y(new_n21258));
  nand_5 g18910(.A(new_n21258), .B(new_n21250), .Y(new_n21259));
  nand_5 g18911(.A(new_n21259), .B(new_n21249), .Y(new_n21260));
  nand_5 g18912(.A(new_n21260), .B(new_n11408), .Y(new_n21261));
  xor_4  g18913(.A(new_n21260), .B(new_n11408), .Y(new_n21262));
  nand_5 g18914(.A(new_n21262), .B(new_n14179), .Y(new_n21263));
  nand_5 g18915(.A(new_n21263), .B(new_n21261), .Y(new_n21264));
  or_6   g18916(.A(new_n21264), .B(new_n21248), .Y(new_n21265));
  nand_5 g18917(.A(new_n21265), .B(new_n21247), .Y(new_n21266));
  xor_4  g18918(.A(new_n21266), .B(new_n21245), .Y(po0387));
  xor_4  g18919(.A(new_n21194), .B(new_n21193), .Y(po0388));
  nand_5 g18920(.A(new_n19790), .B(new_n10325), .Y(new_n21269));
  or_6   g18921(.A(new_n19794), .B(new_n19791), .Y(new_n21270));
  nand_5 g18922(.A(new_n21270), .B(new_n21269), .Y(new_n21271));
  nand_5 g18923(.A(new_n19788), .B(new_n19784), .Y(new_n21272));
  nand_5 g18924(.A(new_n21272), .B(new_n19783), .Y(new_n21273));
  not_8  g18925(.A(new_n21273), .Y(new_n21274));
  and_6  g18926(.A(new_n21274), .B(new_n21271), .Y(new_n21275));
  nor_5  g18927(.A(new_n21274), .B(new_n21271), .Y(new_n21276));
  nor_5  g18928(.A(new_n21276), .B(new_n21275), .Y(new_n21277));
  xor_4  g18929(.A(new_n21277), .B(new_n10425), .Y(po0389));
  xor_4  g18930(.A(new_n9125), .B(new_n9123), .Y(po0390));
  xnor_4 g18931(.A(new_n9371), .B(new_n9314), .Y(po0391));
  xor_4  g18932(.A(new_n20111), .B(new_n16815), .Y(po0392));
  nand_5 g18933(.A(new_n18034), .B(new_n15550), .Y(new_n21282));
  not_8  g18934(.A(new_n18052), .Y(new_n21283));
  nand_5 g18935(.A(new_n21283), .B(new_n18051), .Y(new_n21284));
  nand_5 g18936(.A(new_n21284), .B(new_n21282), .Y(po0393));
  xor_4  g18937(.A(new_n5167), .B(new_n5158), .Y(po0394));
  xor_4  g18938(.A(new_n8948), .B(new_n8947), .Y(po0395));
  or_6   g18939(.A(new_n6946), .B(new_n6944), .Y(new_n21288));
  nand_5 g18940(.A(new_n6947), .B(pi533), .Y(new_n21289));
  nand_5 g18941(.A(new_n21289), .B(new_n21288), .Y(new_n21290));
  xor_4  g18942(.A(new_n21290), .B(new_n12085), .Y(new_n21291));
  xor_4  g18943(.A(new_n21291), .B(pi735), .Y(new_n21292));
  nor_5  g18944(.A(new_n21292), .B(new_n17355), .Y(new_n21293));
  not_8  g18945(.A(new_n6939), .Y(new_n21294));
  nand_5 g18946(.A(new_n6948), .B(new_n21294), .Y(new_n21295));
  or_6   g18947(.A(new_n6949), .B(new_n6930), .Y(new_n21296));
  nand_5 g18948(.A(new_n21296), .B(new_n21295), .Y(new_n21297));
  xor_4  g18949(.A(new_n21292), .B(new_n17354), .Y(new_n21298));
  nor_5  g18950(.A(new_n21298), .B(new_n21297), .Y(new_n21299));
  or_6   g18951(.A(new_n21299), .B(new_n21293), .Y(new_n21300));
  or_6   g18952(.A(new_n21290), .B(new_n12085), .Y(new_n21301));
  nand_5 g18953(.A(new_n21291), .B(new_n10554), .Y(new_n21302));
  nand_5 g18954(.A(new_n21302), .B(new_n21301), .Y(new_n21303));
  xor_4  g18955(.A(new_n21303), .B(new_n12083), .Y(new_n21304));
  xor_4  g18956(.A(new_n21304), .B(new_n17353), .Y(new_n21305));
  xnor_4 g18957(.A(new_n21305), .B(new_n21300), .Y(po0396));
  xnor_4 g18958(.A(new_n10948), .B(new_n10921), .Y(po0397));
  nor_5  g18959(.A(new_n12168), .B(new_n12166), .Y(po0398));
  or_6   g18960(.A(new_n20152), .B(new_n6158), .Y(new_n21309));
  nand_5 g18961(.A(new_n20153), .B(pi338), .Y(new_n21310));
  nand_5 g18962(.A(new_n21310), .B(new_n21309), .Y(new_n21311));
  xor_4  g18963(.A(new_n6169), .B(new_n3991), .Y(new_n21312));
  not_8  g18964(.A(new_n21312), .Y(new_n21313));
  xor_4  g18965(.A(new_n21313), .B(new_n21311), .Y(new_n21314));
  not_8  g18966(.A(new_n20154), .Y(new_n21315));
  nor_5  g18967(.A(new_n20170), .B(new_n21315), .Y(new_n21316));
  nor_5  g18968(.A(new_n20171), .B(new_n9823), .Y(new_n21317));
  or_6   g18969(.A(new_n21317), .B(new_n21316), .Y(new_n21318));
  xor_4  g18970(.A(new_n21318), .B(new_n21314), .Y(new_n21319));
  xor_4  g18971(.A(new_n21319), .B(new_n9830), .Y(po0399));
  xor_4  g18972(.A(new_n21065), .B(new_n9763), .Y(new_n21321));
  not_8  g18973(.A(new_n21321), .Y(new_n21322));
  or_6   g18974(.A(new_n20998), .B(new_n9796), .Y(new_n21323));
  xor_4  g18975(.A(new_n20998), .B(new_n9796), .Y(new_n21324));
  nor_5  g18976(.A(new_n11078), .B(new_n9843), .Y(new_n21325));
  nor_5  g18977(.A(new_n11083), .B(new_n11080), .Y(new_n21326));
  nor_5  g18978(.A(new_n21326), .B(new_n21325), .Y(new_n21327));
  nand_5 g18979(.A(new_n21327), .B(new_n21324), .Y(new_n21328));
  nand_5 g18980(.A(new_n21328), .B(new_n21323), .Y(new_n21329));
  xor_4  g18981(.A(new_n21329), .B(new_n21322), .Y(new_n21330));
  not_8  g18982(.A(new_n21330), .Y(new_n21331));
  xor_4  g18983(.A(new_n21331), .B(new_n11623), .Y(new_n21332));
  not_8  g18984(.A(new_n21332), .Y(new_n21333));
  xor_4  g18985(.A(new_n21327), .B(new_n21324), .Y(new_n21334));
  nand_5 g18986(.A(new_n21334), .B(new_n11602), .Y(new_n21335));
  xor_4  g18987(.A(new_n21334), .B(new_n11602), .Y(new_n21336));
  or_6   g18988(.A(new_n11084), .B(new_n11076), .Y(new_n21337));
  not_8  g18989(.A(new_n11067), .Y(new_n21338));
  nand_5 g18990(.A(new_n11085), .B(new_n21338), .Y(new_n21339));
  nand_5 g18991(.A(new_n21339), .B(new_n21337), .Y(new_n21340));
  nand_5 g18992(.A(new_n21340), .B(new_n21336), .Y(new_n21341));
  nand_5 g18993(.A(new_n21341), .B(new_n21335), .Y(new_n21342));
  xor_4  g18994(.A(new_n21342), .B(new_n21333), .Y(po0400));
  or_6   g18995(.A(new_n20709), .B(new_n7802), .Y(new_n21344));
  not_8  g18996(.A(new_n18085), .Y(new_n21345));
  nand_5 g18997(.A(new_n18070), .B(new_n7820), .Y(new_n21346));
  nand_5 g18998(.A(new_n18069), .B(new_n7818), .Y(new_n21347));
  nand_5 g18999(.A(new_n21347), .B(new_n21346), .Y(new_n21348));
  xor_4  g19000(.A(new_n21348), .B(new_n7725), .Y(new_n21349));
  nand_5 g19001(.A(new_n21349), .B(new_n21345), .Y(new_n21350));
  not_8  g19002(.A(new_n21349), .Y(new_n21351));
  nand_5 g19003(.A(new_n18069), .B(new_n7821), .Y(new_n21352));
  nand_5 g19004(.A(new_n21352), .B(new_n21351), .Y(new_n21353));
  nand_5 g19005(.A(new_n21353), .B(new_n21350), .Y(new_n21354));
  nand_5 g19006(.A(new_n21354), .B(new_n7814), .Y(new_n21355));
  xor_4  g19007(.A(new_n21354), .B(new_n7814), .Y(new_n21356));
  nand_5 g19008(.A(new_n21356), .B(new_n18100), .Y(new_n21357));
  nand_5 g19009(.A(new_n21357), .B(new_n21355), .Y(new_n21358));
  or_6   g19010(.A(new_n21358), .B(new_n7812), .Y(new_n21359));
  xor_4  g19011(.A(new_n21358), .B(new_n7813), .Y(new_n21360));
  not_8  g19012(.A(new_n21360), .Y(new_n21361));
  nand_5 g19013(.A(new_n21361), .B(new_n18123), .Y(new_n21362));
  nand_5 g19014(.A(new_n21362), .B(new_n21359), .Y(new_n21363));
  nor_5  g19015(.A(new_n21363), .B(new_n18146), .Y(new_n21364));
  xor_4  g19016(.A(new_n21363), .B(new_n18147), .Y(new_n21365));
  nor_5  g19017(.A(new_n21365), .B(new_n7810), .Y(new_n21366));
  or_6   g19018(.A(new_n21366), .B(new_n21364), .Y(new_n21367));
  or_6   g19019(.A(new_n21367), .B(new_n7806), .Y(new_n21368));
  xor_4  g19020(.A(new_n21367), .B(new_n7806), .Y(new_n21369));
  nand_5 g19021(.A(new_n21369), .B(new_n18166), .Y(new_n21370));
  nand_5 g19022(.A(new_n21370), .B(new_n21368), .Y(new_n21371));
  xor_4  g19023(.A(new_n20709), .B(new_n7802), .Y(new_n21372));
  nand_5 g19024(.A(new_n21372), .B(new_n21371), .Y(new_n21373));
  nand_5 g19025(.A(new_n21373), .B(new_n21344), .Y(new_n21374));
  nand_5 g19026(.A(new_n21374), .B(new_n7797), .Y(new_n21375));
  xor_4  g19027(.A(new_n21374), .B(new_n7797), .Y(new_n21376));
  nand_5 g19028(.A(new_n21376), .B(new_n20718), .Y(new_n21377));
  nand_5 g19029(.A(new_n21377), .B(new_n21375), .Y(new_n21378));
  nor_5  g19030(.A(new_n21378), .B(new_n7791), .Y(new_n21379));
  xor_4  g19031(.A(new_n21378), .B(new_n7790), .Y(new_n21380));
  nor_5  g19032(.A(new_n21380), .B(new_n20730), .Y(new_n21381));
  nor_5  g19033(.A(new_n21381), .B(new_n21379), .Y(new_n21382));
  xor_4  g19034(.A(new_n21382), .B(new_n7788), .Y(new_n21383));
  xor_4  g19035(.A(new_n21383), .B(new_n20695), .Y(po0401));
  xor_4  g19036(.A(pi721), .B(new_n16220), .Y(new_n21385));
  nand_5 g19037(.A(pi417), .B(new_n16199), .Y(new_n21386));
  xor_4  g19038(.A(pi417), .B(new_n16199), .Y(new_n21387));
  nand_5 g19039(.A(pi348), .B(new_n16167), .Y(new_n21388));
  xor_4  g19040(.A(pi348), .B(new_n16167), .Y(new_n21389));
  nand_5 g19041(.A(pi659), .B(new_n5196), .Y(new_n21390));
  xor_4  g19042(.A(pi659), .B(new_n5196), .Y(new_n21391));
  nand_5 g19043(.A(pi662), .B(new_n5192), .Y(new_n21392));
  nand_5 g19044(.A(pi831), .B(new_n5128), .Y(new_n21393));
  xor_4  g19045(.A(pi831), .B(new_n5128), .Y(new_n21394));
  nand_5 g19046(.A(pi501), .B(new_n5131), .Y(new_n21395));
  xor_4  g19047(.A(pi501), .B(new_n5131), .Y(new_n21396));
  nand_5 g19048(.A(new_n5046), .B(pi589), .Y(new_n21397));
  xor_4  g19049(.A(pi733), .B(new_n2484), .Y(new_n21398));
  nand_5 g19050(.A(new_n5043), .B(pi077), .Y(new_n21399));
  not_8  g19051(.A(new_n21399), .Y(new_n21400));
  nand_5 g19052(.A(new_n21400), .B(new_n21398), .Y(new_n21401));
  nand_5 g19053(.A(new_n21401), .B(new_n21397), .Y(new_n21402));
  nand_5 g19054(.A(new_n21402), .B(new_n21396), .Y(new_n21403));
  nand_5 g19055(.A(new_n21403), .B(new_n21395), .Y(new_n21404));
  nand_5 g19056(.A(new_n21404), .B(new_n21394), .Y(new_n21405));
  nand_5 g19057(.A(new_n21405), .B(new_n21393), .Y(new_n21406));
  xor_4  g19058(.A(pi662), .B(new_n5192), .Y(new_n21407));
  nand_5 g19059(.A(new_n21407), .B(new_n21406), .Y(new_n21408));
  nand_5 g19060(.A(new_n21408), .B(new_n21392), .Y(new_n21409));
  nand_5 g19061(.A(new_n21409), .B(new_n21391), .Y(new_n21410));
  nand_5 g19062(.A(new_n21410), .B(new_n21390), .Y(new_n21411));
  nand_5 g19063(.A(new_n21411), .B(new_n21389), .Y(new_n21412));
  nand_5 g19064(.A(new_n21412), .B(new_n21388), .Y(new_n21413));
  nand_5 g19065(.A(new_n21413), .B(new_n21387), .Y(new_n21414));
  nand_5 g19066(.A(new_n21414), .B(new_n21386), .Y(new_n21415));
  xor_4  g19067(.A(new_n21415), .B(new_n21385), .Y(new_n21416));
  xor_4  g19068(.A(new_n21416), .B(new_n14631), .Y(new_n21417));
  xnor_4 g19069(.A(new_n21413), .B(new_n21387), .Y(new_n21418));
  nor_5  g19070(.A(new_n21418), .B(new_n14534), .Y(new_n21419));
  xor_4  g19071(.A(new_n21418), .B(new_n14535), .Y(new_n21420));
  xor_4  g19072(.A(new_n21411), .B(new_n21389), .Y(new_n21421));
  not_8  g19073(.A(new_n21421), .Y(new_n21422));
  nand_5 g19074(.A(new_n21422), .B(new_n14564), .Y(new_n21423));
  xor_4  g19075(.A(new_n21409), .B(new_n21391), .Y(new_n21424));
  or_6   g19076(.A(new_n21424), .B(new_n14568), .Y(new_n21425));
  xor_4  g19077(.A(new_n21424), .B(new_n14568), .Y(new_n21426));
  xor_4  g19078(.A(new_n21407), .B(new_n21406), .Y(new_n21427));
  or_6   g19079(.A(new_n21427), .B(new_n14571), .Y(new_n21428));
  xor_4  g19080(.A(new_n21427), .B(new_n14571), .Y(new_n21429));
  xnor_4 g19081(.A(new_n21404), .B(new_n21394), .Y(new_n21430));
  or_6   g19082(.A(new_n21430), .B(new_n14575), .Y(new_n21431));
  xor_4  g19083(.A(new_n21402), .B(new_n21396), .Y(new_n21432));
  nor_5  g19084(.A(new_n21432), .B(new_n14579), .Y(new_n21433));
  xor_4  g19085(.A(new_n21432), .B(new_n14579), .Y(new_n21434));
  nor_5  g19086(.A(new_n21399), .B(new_n14583), .Y(new_n21435));
  nand_5 g19087(.A(new_n21398), .B(new_n14586), .Y(new_n21436));
  nor_5  g19088(.A(new_n21436), .B(new_n21435), .Y(new_n21437));
  nand_5 g19089(.A(pi654), .B(new_n2487), .Y(new_n21438));
  nor_5  g19090(.A(new_n21438), .B(new_n14583), .Y(new_n21439));
  not_8  g19091(.A(new_n21439), .Y(new_n21440));
  nand_5 g19092(.A(new_n21400), .B(new_n14583), .Y(new_n21441));
  nand_5 g19093(.A(new_n21441), .B(new_n21440), .Y(new_n21442));
  xor_4  g19094(.A(new_n21398), .B(new_n14593), .Y(new_n21443));
  not_8  g19095(.A(new_n21443), .Y(new_n21444));
  nor_5  g19096(.A(new_n21444), .B(new_n21442), .Y(new_n21445));
  nand_5 g19097(.A(new_n21440), .B(new_n21401), .Y(new_n21446));
  nor_5  g19098(.A(new_n21446), .B(new_n21445), .Y(new_n21447));
  nor_5  g19099(.A(new_n21447), .B(new_n21437), .Y(new_n21448));
  and_6  g19100(.A(new_n21448), .B(new_n21434), .Y(new_n21449));
  nor_5  g19101(.A(new_n21449), .B(new_n21433), .Y(new_n21450));
  xor_4  g19102(.A(new_n21430), .B(new_n14575), .Y(new_n21451));
  nand_5 g19103(.A(new_n21451), .B(new_n21450), .Y(new_n21452));
  nand_5 g19104(.A(new_n21452), .B(new_n21431), .Y(new_n21453));
  not_8  g19105(.A(new_n21453), .Y(new_n21454));
  nand_5 g19106(.A(new_n21454), .B(new_n21429), .Y(new_n21455));
  nand_5 g19107(.A(new_n21455), .B(new_n21428), .Y(new_n21456));
  nand_5 g19108(.A(new_n21456), .B(new_n21426), .Y(new_n21457));
  nand_5 g19109(.A(new_n21457), .B(new_n21425), .Y(new_n21458));
  xor_4  g19110(.A(new_n21421), .B(new_n14564), .Y(new_n21459));
  not_8  g19111(.A(new_n21459), .Y(new_n21460));
  nand_5 g19112(.A(new_n21460), .B(new_n21458), .Y(new_n21461));
  nand_5 g19113(.A(new_n21461), .B(new_n21423), .Y(new_n21462));
  nor_5  g19114(.A(new_n21462), .B(new_n21420), .Y(new_n21463));
  nor_5  g19115(.A(new_n21463), .B(new_n21419), .Y(new_n21464));
  xnor_4 g19116(.A(new_n21464), .B(new_n21417), .Y(po0402));
  xor_4  g19117(.A(new_n18049), .B(new_n18046), .Y(po0403));
  xnor_4 g19118(.A(new_n5006), .B(new_n4974), .Y(po0404));
  xor_4  g19119(.A(new_n3362), .B(new_n3360), .Y(po0405));
  nand_5 g19120(.A(pi321), .B(new_n6379), .Y(new_n21469));
  nand_5 g19121(.A(new_n21081), .B(pi197), .Y(new_n21470));
  nand_5 g19122(.A(new_n21470), .B(new_n11500), .Y(new_n21471));
  and_6  g19123(.A(new_n21471), .B(new_n21469), .Y(new_n21472));
  nor_5  g19124(.A(new_n11506), .B(pi194), .Y(new_n21473));
  nor_5  g19125(.A(new_n21087), .B(new_n6294), .Y(new_n21474));
  nor_5  g19126(.A(new_n21474), .B(new_n21473), .Y(new_n21475));
  xor_4  g19127(.A(new_n21087), .B(new_n6294), .Y(new_n21476));
  nand_5 g19128(.A(pi782), .B(pi199), .Y(new_n21477));
  xor_4  g19129(.A(pi782), .B(pi199), .Y(new_n21478));
  nand_5 g19130(.A(pi627), .B(pi150), .Y(new_n21479));
  nand_5 g19131(.A(pi826), .B(pi643), .Y(new_n21480));
  xor_4  g19132(.A(pi826), .B(pi643), .Y(new_n21481));
  nand_5 g19133(.A(pi320), .B(pi210), .Y(new_n21482));
  nand_5 g19134(.A(new_n21000), .B(new_n6106), .Y(new_n21483));
  nand_5 g19135(.A(pi129), .B(pi042), .Y(new_n21484));
  xor_4  g19136(.A(pi129), .B(pi042), .Y(new_n21485));
  nand_5 g19137(.A(pi658), .B(pi017), .Y(new_n21486));
  nand_5 g19138(.A(new_n16640), .B(new_n16638), .Y(new_n21487));
  nand_5 g19139(.A(new_n21487), .B(new_n21486), .Y(new_n21488));
  nand_5 g19140(.A(new_n21488), .B(new_n21485), .Y(new_n21489));
  nand_5 g19141(.A(new_n21489), .B(new_n21484), .Y(new_n21490));
  nand_5 g19142(.A(new_n21490), .B(new_n21483), .Y(new_n21491));
  nand_5 g19143(.A(new_n21491), .B(new_n21482), .Y(new_n21492));
  nand_5 g19144(.A(new_n21492), .B(new_n21481), .Y(new_n21493));
  nand_5 g19145(.A(new_n21493), .B(new_n21480), .Y(new_n21494));
  xor_4  g19146(.A(pi627), .B(pi150), .Y(new_n21495));
  nand_5 g19147(.A(new_n21495), .B(new_n21494), .Y(new_n21496));
  nand_5 g19148(.A(new_n21496), .B(new_n21479), .Y(new_n21497));
  nand_5 g19149(.A(new_n21497), .B(new_n21478), .Y(new_n21498));
  nand_5 g19150(.A(new_n21498), .B(new_n21477), .Y(new_n21499));
  and_6  g19151(.A(new_n21499), .B(new_n21476), .Y(new_n21500));
  xnor_4 g19152(.A(new_n21497), .B(new_n21478), .Y(new_n21501));
  nor_5  g19153(.A(new_n21501), .B(pi202), .Y(new_n21502));
  xnor_4 g19154(.A(new_n21495), .B(new_n21494), .Y(new_n21503));
  nand_5 g19155(.A(new_n21503), .B(pi063), .Y(new_n21504));
  xor_4  g19156(.A(new_n21503), .B(pi063), .Y(new_n21505));
  not_8  g19157(.A(pi538), .Y(new_n21506));
  xor_4  g19158(.A(new_n21492), .B(new_n21481), .Y(new_n21507));
  or_6   g19159(.A(new_n21507), .B(new_n21506), .Y(new_n21508));
  nand_5 g19160(.A(new_n21483), .B(new_n21482), .Y(new_n21509));
  xnor_4 g19161(.A(new_n21509), .B(new_n21490), .Y(new_n21510));
  or_6   g19162(.A(new_n21510), .B(new_n21115), .Y(new_n21511));
  nand_5 g19163(.A(new_n21510), .B(new_n21115), .Y(new_n21512));
  xnor_4 g19164(.A(new_n21488), .B(new_n21485), .Y(new_n21513));
  nand_5 g19165(.A(new_n21513), .B(pi746), .Y(new_n21514));
  xor_4  g19166(.A(new_n21513), .B(pi746), .Y(new_n21515));
  nand_5 g19167(.A(new_n16643), .B(new_n16636), .Y(new_n21516));
  nand_5 g19168(.A(new_n21516), .B(new_n16642), .Y(new_n21517));
  nand_5 g19169(.A(new_n21517), .B(new_n21515), .Y(new_n21518));
  nand_5 g19170(.A(new_n21518), .B(new_n21514), .Y(new_n21519));
  nand_5 g19171(.A(new_n21519), .B(new_n21512), .Y(new_n21520));
  nand_5 g19172(.A(new_n21520), .B(new_n21511), .Y(new_n21521));
  xor_4  g19173(.A(new_n21507), .B(new_n21506), .Y(new_n21522));
  nand_5 g19174(.A(new_n21522), .B(new_n21521), .Y(new_n21523));
  nand_5 g19175(.A(new_n21523), .B(new_n21508), .Y(new_n21524));
  nand_5 g19176(.A(new_n21524), .B(new_n21505), .Y(new_n21525));
  nand_5 g19177(.A(new_n21525), .B(new_n21504), .Y(new_n21526));
  xor_4  g19178(.A(new_n21501), .B(new_n21183), .Y(new_n21527));
  nor_5  g19179(.A(new_n21527), .B(new_n21526), .Y(new_n21528));
  nor_5  g19180(.A(new_n21528), .B(new_n21502), .Y(new_n21529));
  xor_4  g19181(.A(new_n21499), .B(new_n21476), .Y(new_n21530));
  not_8  g19182(.A(new_n21530), .Y(new_n21531));
  nor_5  g19183(.A(new_n21531), .B(new_n21529), .Y(new_n21532));
  nor_5  g19184(.A(new_n21532), .B(new_n21500), .Y(new_n21533));
  nand_5 g19185(.A(new_n21533), .B(new_n21475), .Y(new_n21534));
  or_6   g19186(.A(new_n21534), .B(new_n21472), .Y(new_n21535));
  nor_5  g19187(.A(new_n21533), .B(new_n21475), .Y(new_n21536));
  not_8  g19188(.A(new_n21536), .Y(new_n21537));
  nor_5  g19189(.A(new_n21469), .B(pi340), .Y(new_n21538));
  nand_5 g19190(.A(new_n21538), .B(new_n21537), .Y(new_n21539));
  nand_5 g19191(.A(new_n21539), .B(new_n21535), .Y(new_n21540));
  xnor_4 g19192(.A(new_n21540), .B(new_n15737), .Y(new_n21541));
  xor_4  g19193(.A(new_n21530), .B(new_n21529), .Y(new_n21542));
  nand_5 g19194(.A(new_n21542), .B(new_n15746), .Y(new_n21543));
  xor_4  g19195(.A(new_n21527), .B(new_n21526), .Y(new_n21544));
  nor_5  g19196(.A(new_n21544), .B(new_n15754), .Y(new_n21545));
  xor_4  g19197(.A(new_n21524), .B(new_n21505), .Y(new_n21546));
  not_8  g19198(.A(new_n21546), .Y(new_n21547));
  nor_5  g19199(.A(new_n21547), .B(new_n15803), .Y(new_n21548));
  xor_4  g19200(.A(new_n21546), .B(new_n15803), .Y(new_n21549));
  not_8  g19201(.A(new_n15795), .Y(new_n21550));
  xor_4  g19202(.A(new_n21522), .B(new_n21521), .Y(new_n21551));
  nor_5  g19203(.A(new_n21551), .B(new_n21550), .Y(new_n21552));
  nand_5 g19204(.A(new_n21512), .B(new_n21511), .Y(new_n21553));
  xor_4  g19205(.A(new_n21553), .B(new_n21519), .Y(new_n21554));
  nor_5  g19206(.A(new_n21554), .B(new_n15786), .Y(new_n21555));
  xor_4  g19207(.A(new_n21517), .B(new_n21515), .Y(new_n21556));
  not_8  g19208(.A(new_n21556), .Y(new_n21557));
  nor_5  g19209(.A(new_n21557), .B(new_n15781), .Y(new_n21558));
  xor_4  g19210(.A(new_n21556), .B(new_n15781), .Y(new_n21559));
  nand_5 g19211(.A(new_n16645), .B(new_n15771), .Y(new_n21560));
  or_6   g19212(.A(new_n16646), .B(new_n16634), .Y(new_n21561));
  nand_5 g19213(.A(new_n21561), .B(new_n21560), .Y(new_n21562));
  nor_5  g19214(.A(new_n21562), .B(new_n21559), .Y(new_n21563));
  nor_5  g19215(.A(new_n21563), .B(new_n21558), .Y(new_n21564));
  xor_4  g19216(.A(new_n21554), .B(new_n15757), .Y(new_n21565));
  nor_5  g19217(.A(new_n21565), .B(new_n21564), .Y(new_n21566));
  or_6   g19218(.A(new_n21566), .B(new_n21555), .Y(new_n21567));
  xor_4  g19219(.A(new_n21551), .B(new_n15795), .Y(new_n21568));
  nor_5  g19220(.A(new_n21568), .B(new_n21567), .Y(new_n21569));
  or_6   g19221(.A(new_n21569), .B(new_n21552), .Y(new_n21570));
  nor_5  g19222(.A(new_n21570), .B(new_n21549), .Y(new_n21571));
  nor_5  g19223(.A(new_n21571), .B(new_n21548), .Y(new_n21572));
  xor_4  g19224(.A(new_n21544), .B(new_n15750), .Y(new_n21573));
  nor_5  g19225(.A(new_n21573), .B(new_n21572), .Y(new_n21574));
  nor_5  g19226(.A(new_n21574), .B(new_n21545), .Y(new_n21575));
  xor_4  g19227(.A(new_n21542), .B(new_n15745), .Y(new_n21576));
  or_6   g19228(.A(new_n21576), .B(new_n21575), .Y(new_n21577));
  nand_5 g19229(.A(new_n21577), .B(new_n21543), .Y(new_n21578));
  or_6   g19230(.A(new_n21578), .B(new_n15812), .Y(new_n21579));
  xor_4  g19231(.A(new_n21578), .B(new_n15812), .Y(new_n21580));
  nand_5 g19232(.A(new_n21537), .B(new_n21534), .Y(new_n21581));
  xor_4  g19233(.A(new_n21581), .B(pi340), .Y(new_n21582));
  nand_5 g19234(.A(new_n21470), .B(new_n21469), .Y(new_n21583));
  xor_4  g19235(.A(new_n21583), .B(new_n21582), .Y(new_n21584));
  nand_5 g19236(.A(new_n21584), .B(new_n21580), .Y(new_n21585));
  nand_5 g19237(.A(new_n21585), .B(new_n21579), .Y(new_n21586));
  nor_5  g19238(.A(new_n21470), .B(new_n11500), .Y(new_n21587));
  nand_5 g19239(.A(new_n21587), .B(new_n21534), .Y(new_n21588));
  nand_5 g19240(.A(new_n21536), .B(new_n21472), .Y(new_n21589));
  nand_5 g19241(.A(new_n21589), .B(new_n21588), .Y(new_n21590));
  or_6   g19242(.A(new_n21590), .B(new_n21540), .Y(new_n21591));
  xor_4  g19243(.A(new_n21591), .B(new_n15741), .Y(new_n21592));
  nor_5  g19244(.A(new_n21592), .B(new_n21586), .Y(new_n21593));
  nand_5 g19245(.A(new_n21593), .B(new_n21541), .Y(new_n21594));
  not_8  g19246(.A(new_n21593), .Y(new_n21595));
  nor_5  g19247(.A(new_n21591), .B(new_n15742), .Y(new_n21596));
  nor_5  g19248(.A(new_n21596), .B(new_n21541), .Y(new_n21597));
  nand_5 g19249(.A(new_n21597), .B(new_n21595), .Y(new_n21598));
  nand_5 g19250(.A(new_n21598), .B(new_n21594), .Y(po0406));
  or_6   g19251(.A(new_n18959), .B(new_n18938), .Y(new_n21600));
  nand_5 g19252(.A(new_n18961), .B(new_n18958), .Y(new_n21601));
  nand_5 g19253(.A(new_n21601), .B(new_n21600), .Y(po0407));
  xor_4  g19254(.A(new_n12281), .B(new_n12250), .Y(po0408));
  xor_4  g19255(.A(new_n10030), .B(new_n10029), .Y(po0409));
  xor_4  g19256(.A(new_n20353), .B(new_n20352), .Y(po0410));
  xor_4  g19257(.A(new_n19583), .B(new_n20323), .Y(po0412));
  nand_5 g19258(.A(new_n16439), .B(new_n16437), .Y(new_n21607));
  nand_5 g19259(.A(new_n21607), .B(new_n16438), .Y(new_n21608));
  xor_4  g19260(.A(pi661), .B(pi124), .Y(new_n21609));
  not_8  g19261(.A(new_n21609), .Y(new_n21610));
  xor_4  g19262(.A(new_n21610), .B(new_n6099), .Y(new_n21611));
  not_8  g19263(.A(new_n21611), .Y(new_n21612));
  xor_4  g19264(.A(new_n21612), .B(new_n21608), .Y(new_n21613));
  not_8  g19265(.A(new_n21613), .Y(new_n21614));
  not_8  g19266(.A(new_n2982), .Y(new_n21615));
  nand_5 g19267(.A(new_n2987), .B(new_n8641), .Y(new_n21616));
  not_8  g19268(.A(new_n8645), .Y(new_n21617));
  nand_5 g19269(.A(new_n21617), .B(new_n8642), .Y(new_n21618));
  nand_5 g19270(.A(new_n21618), .B(new_n21616), .Y(new_n21619));
  or_6   g19271(.A(new_n21619), .B(new_n21615), .Y(new_n21620));
  nand_5 g19272(.A(new_n21619), .B(new_n21615), .Y(new_n21621));
  nand_5 g19273(.A(new_n21621), .B(pi671), .Y(new_n21622));
  nand_5 g19274(.A(new_n21622), .B(new_n21620), .Y(new_n21623));
  or_6   g19275(.A(new_n21623), .B(new_n2938), .Y(new_n21624));
  nand_5 g19276(.A(new_n21623), .B(new_n2938), .Y(new_n21625));
  nand_5 g19277(.A(new_n21625), .B(new_n21624), .Y(new_n21626));
  xor_4  g19278(.A(new_n21626), .B(new_n16070), .Y(new_n21627));
  not_8  g19279(.A(new_n21627), .Y(new_n21628));
  nand_5 g19280(.A(new_n8639), .B(new_n8575), .Y(new_n21629));
  nand_5 g19281(.A(new_n8646), .B(new_n8640), .Y(new_n21630));
  nand_5 g19282(.A(new_n21630), .B(new_n21629), .Y(new_n21631));
  not_8  g19283(.A(new_n21631), .Y(new_n21632));
  nand_5 g19284(.A(new_n21621), .B(new_n21620), .Y(new_n21633));
  xor_4  g19285(.A(new_n21633), .B(pi671), .Y(new_n21634));
  nand_5 g19286(.A(new_n21634), .B(new_n21632), .Y(new_n21635));
  xor_4  g19287(.A(new_n21634), .B(new_n21632), .Y(new_n21636));
  nand_5 g19288(.A(new_n21636), .B(new_n16430), .Y(new_n21637));
  nand_5 g19289(.A(new_n21637), .B(new_n21635), .Y(new_n21638));
  nand_5 g19290(.A(new_n21638), .B(new_n21628), .Y(new_n21639));
  xor_4  g19291(.A(new_n21638), .B(new_n21628), .Y(new_n21640));
  nand_5 g19292(.A(new_n21640), .B(new_n16442), .Y(new_n21641));
  nand_5 g19293(.A(new_n21641), .B(new_n21639), .Y(new_n21642));
  xor_4  g19294(.A(new_n18390), .B(new_n16066), .Y(new_n21643));
  nand_5 g19295(.A(new_n21624), .B(pi537), .Y(new_n21644));
  nand_5 g19296(.A(new_n21644), .B(new_n21625), .Y(new_n21645));
  xor_4  g19297(.A(new_n21645), .B(new_n21643), .Y(new_n21646));
  xor_4  g19298(.A(new_n21646), .B(new_n21642), .Y(new_n21647));
  xor_4  g19299(.A(new_n21647), .B(new_n21614), .Y(po0413));
  xor_4  g19300(.A(new_n2612), .B(pi565), .Y(new_n21649));
  nand_5 g19301(.A(new_n2616), .B(new_n11526), .Y(new_n21650));
  not_8  g19302(.A(new_n21650), .Y(new_n21651));
  not_8  g19303(.A(new_n9726), .Y(new_n21652));
  nor_5  g19304(.A(new_n9762), .B(new_n21652), .Y(new_n21653));
  nor_5  g19305(.A(new_n21653), .B(new_n21651), .Y(new_n21654));
  xor_4  g19306(.A(new_n21654), .B(new_n21649), .Y(new_n21655));
  nor_5  g19307(.A(new_n2820), .B(pi835), .Y(new_n21656));
  nor_5  g19308(.A(new_n9792), .B(new_n9791), .Y(new_n21657));
  nor_5  g19309(.A(new_n21657), .B(new_n21656), .Y(new_n21658));
  xor_4  g19310(.A(new_n2844), .B(new_n17484), .Y(new_n21659));
  xor_4  g19311(.A(new_n21659), .B(new_n21658), .Y(new_n21660));
  or_6   g19312(.A(new_n21660), .B(new_n21655), .Y(new_n21661));
  nor_5  g19313(.A(new_n9793), .B(new_n9763), .Y(new_n21662));
  nor_5  g19314(.A(new_n9851), .B(new_n9794), .Y(new_n21663));
  or_6   g19315(.A(new_n21663), .B(new_n21662), .Y(new_n21664));
  xor_4  g19316(.A(new_n21660), .B(new_n21655), .Y(new_n21665));
  nand_5 g19317(.A(new_n21665), .B(new_n21664), .Y(new_n21666));
  nand_5 g19318(.A(new_n21666), .B(new_n21661), .Y(new_n21667));
  nand_5 g19319(.A(new_n2847), .B(new_n17484), .Y(new_n21668));
  not_8  g19320(.A(new_n21668), .Y(new_n21669));
  nor_5  g19321(.A(new_n21659), .B(new_n21658), .Y(new_n21670));
  nor_5  g19322(.A(new_n21670), .B(new_n21669), .Y(new_n21671));
  nand_5 g19323(.A(new_n21671), .B(new_n10410), .Y(new_n21672));
  not_8  g19324(.A(new_n21672), .Y(new_n21673));
  nor_5  g19325(.A(new_n21671), .B(new_n10410), .Y(new_n21674));
  nor_5  g19326(.A(new_n21674), .B(new_n21673), .Y(new_n21675));
  not_8  g19327(.A(new_n14814), .Y(new_n21676));
  nor_5  g19328(.A(new_n2612), .B(pi565), .Y(new_n21677));
  not_8  g19329(.A(new_n21649), .Y(new_n21678));
  nor_5  g19330(.A(new_n21654), .B(new_n21678), .Y(new_n21679));
  or_6   g19331(.A(new_n21679), .B(new_n21677), .Y(new_n21680));
  nand_5 g19332(.A(new_n21680), .B(new_n21676), .Y(new_n21681));
  nor_5  g19333(.A(new_n21680), .B(new_n21676), .Y(new_n21682));
  not_8  g19334(.A(new_n21682), .Y(new_n21683));
  nand_5 g19335(.A(new_n21683), .B(new_n21681), .Y(new_n21684));
  xor_4  g19336(.A(new_n21684), .B(new_n21675), .Y(new_n21685));
  not_8  g19337(.A(new_n21685), .Y(new_n21686));
  xor_4  g19338(.A(new_n21686), .B(new_n21667), .Y(po0414));
  xor_4  g19339(.A(new_n17633), .B(new_n6628), .Y(po0415));
  xor_4  g19340(.A(new_n17593), .B(new_n17592), .Y(po0416));
  xor_4  g19341(.A(new_n21376), .B(new_n20718), .Y(po0417));
  xor_4  g19342(.A(new_n11060), .B(new_n11038), .Y(po0418));
  xor_4  g19343(.A(new_n3088), .B(new_n3087), .Y(po0419));
  xor_4  g19344(.A(new_n3102), .B(new_n3051), .Y(po0420));
  xnor_4 g19345(.A(new_n9840), .B(new_n9838), .Y(po0421));
  xor_4  g19346(.A(new_n19828), .B(new_n15736), .Y(new_n21695));
  not_8  g19347(.A(new_n21695), .Y(new_n21696));
  nand_5 g19348(.A(new_n19839), .B(new_n15730), .Y(new_n21697));
  not_8  g19349(.A(new_n21697), .Y(new_n21698));
  xor_4  g19350(.A(new_n19839), .B(new_n15730), .Y(new_n21699));
  not_8  g19351(.A(new_n21699), .Y(new_n21700));
  nor_5  g19352(.A(new_n19841), .B(new_n15684), .Y(new_n21701));
  xor_4  g19353(.A(new_n19841), .B(new_n15685), .Y(new_n21702));
  or_6   g19354(.A(new_n15429), .B(new_n15418), .Y(new_n21703));
  nand_5 g19355(.A(new_n15430), .B(new_n15412), .Y(new_n21704));
  nand_5 g19356(.A(new_n21704), .B(new_n21703), .Y(new_n21705));
  nor_5  g19357(.A(new_n21705), .B(new_n21702), .Y(new_n21706));
  or_6   g19358(.A(new_n21706), .B(new_n21701), .Y(new_n21707));
  nor_5  g19359(.A(new_n21707), .B(new_n21700), .Y(new_n21708));
  nor_5  g19360(.A(new_n21708), .B(new_n21698), .Y(new_n21709));
  xor_4  g19361(.A(new_n21709), .B(new_n21696), .Y(po0422));
  xor_4  g19362(.A(new_n17641), .B(new_n8598), .Y(po0423));
  xnor_4 g19363(.A(new_n18641), .B(new_n18633), .Y(po0424));
  nand_5 g19364(.A(new_n13161), .B(new_n13157), .Y(new_n21713));
  or_6   g19365(.A(new_n13168), .B(new_n13162), .Y(new_n21714));
  nand_5 g19366(.A(new_n21714), .B(new_n21713), .Y(new_n21715));
  nand_5 g19367(.A(new_n21715), .B(new_n18863), .Y(new_n21716));
  xnor_4 g19368(.A(new_n21715), .B(new_n18863), .Y(new_n21717));
  or_6   g19369(.A(new_n21717), .B(new_n17626), .Y(new_n21718));
  nand_5 g19370(.A(new_n21718), .B(new_n21716), .Y(new_n21719));
  or_6   g19371(.A(new_n21719), .B(new_n18857), .Y(new_n21720));
  xor_4  g19372(.A(new_n21719), .B(new_n18857), .Y(new_n21721));
  nand_5 g19373(.A(new_n21721), .B(new_n17650), .Y(new_n21722));
  nand_5 g19374(.A(new_n21722), .B(new_n21720), .Y(new_n21723));
  nor_5  g19375(.A(new_n21723), .B(new_n18854), .Y(new_n21724));
  xor_4  g19376(.A(new_n21723), .B(new_n18853), .Y(new_n21725));
  nor_5  g19377(.A(new_n21725), .B(new_n17624), .Y(new_n21726));
  or_6   g19378(.A(new_n21726), .B(new_n21724), .Y(new_n21727));
  not_8  g19379(.A(new_n13059), .Y(new_n21728));
  nand_5 g19380(.A(new_n17623), .B(new_n17610), .Y(new_n21729));
  nand_5 g19381(.A(new_n21729), .B(new_n17611), .Y(new_n21730));
  nor_5  g19382(.A(new_n21730), .B(new_n21728), .Y(new_n21731));
  nand_5 g19383(.A(new_n21730), .B(new_n21728), .Y(new_n21732));
  not_8  g19384(.A(new_n21732), .Y(new_n21733));
  nor_5  g19385(.A(new_n21733), .B(new_n21731), .Y(new_n21734));
  xor_4  g19386(.A(new_n21734), .B(new_n4839), .Y(new_n21735));
  not_8  g19387(.A(new_n21735), .Y(new_n21736));
  or_6   g19388(.A(new_n21736), .B(new_n21727), .Y(new_n21737));
  xor_4  g19389(.A(new_n21736), .B(new_n21727), .Y(new_n21738));
  nand_5 g19390(.A(new_n21738), .B(new_n18848), .Y(new_n21739));
  nand_5 g19391(.A(new_n21739), .B(new_n21737), .Y(new_n21740));
  nor_5  g19392(.A(new_n21731), .B(pi812), .Y(new_n21741));
  nor_5  g19393(.A(new_n21741), .B(new_n21733), .Y(new_n21742));
  not_8  g19394(.A(new_n21742), .Y(new_n21743));
  xor_4  g19395(.A(new_n17535), .B(new_n13075), .Y(new_n21744));
  xor_4  g19396(.A(new_n21744), .B(new_n21743), .Y(new_n21745));
  not_8  g19397(.A(new_n21745), .Y(new_n21746));
  xor_4  g19398(.A(new_n21746), .B(new_n21740), .Y(new_n21747));
  xor_4  g19399(.A(new_n21747), .B(new_n18901), .Y(po0425));
  xor_4  g19400(.A(new_n18266), .B(new_n13737), .Y(po0426));
  not_8  g19401(.A(new_n21314), .Y(new_n21750));
  nand_5 g19402(.A(new_n21318), .B(new_n21750), .Y(new_n21751));
  or_6   g19403(.A(new_n21319), .B(new_n9830), .Y(new_n21752));
  nand_5 g19404(.A(new_n21752), .B(new_n21751), .Y(new_n21753));
  nor_5  g19405(.A(new_n21753), .B(new_n9836), .Y(new_n21754));
  nand_5 g19406(.A(new_n6169), .B(new_n3991), .Y(new_n21755));
  or_6   g19407(.A(new_n21313), .B(new_n21311), .Y(new_n21756));
  nand_5 g19408(.A(new_n21756), .B(new_n21755), .Y(new_n21757));
  xor_4  g19409(.A(new_n21757), .B(pi613), .Y(new_n21758));
  xor_4  g19410(.A(new_n21758), .B(new_n14820), .Y(new_n21759));
  xor_4  g19411(.A(new_n21753), .B(new_n9835), .Y(new_n21760));
  nor_5  g19412(.A(new_n21760), .B(new_n21759), .Y(new_n21761));
  or_6   g19413(.A(new_n21761), .B(new_n21754), .Y(new_n21762));
  nand_5 g19414(.A(new_n21757), .B(new_n5646), .Y(new_n21763));
  or_6   g19415(.A(new_n21758), .B(new_n6207), .Y(new_n21764));
  nand_5 g19416(.A(new_n21764), .B(new_n21763), .Y(new_n21765));
  nand_5 g19417(.A(new_n21765), .B(new_n6280), .Y(new_n21766));
  or_6   g19418(.A(new_n21765), .B(new_n6280), .Y(new_n21767));
  nand_5 g19419(.A(new_n21767), .B(new_n21766), .Y(new_n21768));
  xor_4  g19420(.A(new_n21768), .B(pi297), .Y(new_n21769));
  or_6   g19421(.A(new_n21769), .B(new_n21762), .Y(new_n21770));
  xor_4  g19422(.A(new_n21769), .B(new_n21762), .Y(new_n21771));
  nand_5 g19423(.A(new_n21771), .B(new_n9843), .Y(new_n21772));
  nand_5 g19424(.A(new_n21772), .B(new_n21770), .Y(new_n21773));
  nand_5 g19425(.A(new_n21766), .B(pi297), .Y(new_n21774));
  nand_5 g19426(.A(new_n21774), .B(new_n21767), .Y(new_n21775));
  nor_5  g19427(.A(new_n21775), .B(new_n6289), .Y(new_n21776));
  and_6  g19428(.A(new_n21775), .B(new_n6289), .Y(new_n21777));
  nor_5  g19429(.A(new_n21777), .B(new_n21776), .Y(new_n21778));
  xor_4  g19430(.A(new_n21778), .B(new_n5640), .Y(new_n21779));
  not_8  g19431(.A(new_n21779), .Y(new_n21780));
  nor_5  g19432(.A(new_n21780), .B(new_n21773), .Y(new_n21781));
  xor_4  g19433(.A(new_n21779), .B(new_n21773), .Y(new_n21782));
  nor_5  g19434(.A(new_n21782), .B(new_n9797), .Y(new_n21783));
  or_6   g19435(.A(new_n21783), .B(new_n21781), .Y(new_n21784));
  nor_5  g19436(.A(new_n21776), .B(new_n5640), .Y(new_n21785));
  nor_5  g19437(.A(new_n21785), .B(new_n21777), .Y(new_n21786));
  nand_5 g19438(.A(new_n21786), .B(new_n6309), .Y(new_n21787));
  or_6   g19439(.A(new_n21786), .B(new_n6309), .Y(new_n21788));
  nand_5 g19440(.A(new_n21788), .B(new_n21787), .Y(new_n21789));
  xor_4  g19441(.A(new_n21789), .B(pi472), .Y(new_n21790));
  nand_5 g19442(.A(new_n21790), .B(new_n21784), .Y(new_n21791));
  xnor_4 g19443(.A(new_n21790), .B(new_n21784), .Y(new_n21792));
  or_6   g19444(.A(new_n21792), .B(new_n9764), .Y(new_n21793));
  nand_5 g19445(.A(new_n21793), .B(new_n21791), .Y(new_n21794));
  nand_5 g19446(.A(new_n21787), .B(pi472), .Y(new_n21795));
  nand_5 g19447(.A(new_n21795), .B(new_n21788), .Y(new_n21796));
  nor_5  g19448(.A(new_n21796), .B(new_n6347), .Y(new_n21797));
  nand_5 g19449(.A(new_n21796), .B(new_n6347), .Y(new_n21798));
  not_8  g19450(.A(new_n21798), .Y(new_n21799));
  nor_5  g19451(.A(new_n21799), .B(new_n21797), .Y(new_n21800));
  xor_4  g19452(.A(new_n21800), .B(new_n5634), .Y(new_n21801));
  nand_5 g19453(.A(new_n21801), .B(new_n21794), .Y(new_n21802));
  not_8  g19454(.A(new_n21655), .Y(new_n21803));
  xnor_4 g19455(.A(new_n21801), .B(new_n21794), .Y(new_n21804));
  or_6   g19456(.A(new_n21804), .B(new_n21803), .Y(new_n21805));
  nand_5 g19457(.A(new_n21805), .B(new_n21802), .Y(new_n21806));
  xor_4  g19458(.A(new_n21806), .B(new_n21684), .Y(new_n21807));
  nor_5  g19459(.A(new_n21797), .B(new_n5634), .Y(new_n21808));
  nor_5  g19460(.A(new_n21808), .B(new_n21799), .Y(new_n21809));
  xor_4  g19461(.A(new_n21809), .B(new_n12552), .Y(new_n21810));
  nor_5  g19462(.A(new_n21810), .B(new_n21807), .Y(new_n21811));
  not_8  g19463(.A(new_n21684), .Y(new_n21812));
  nand_5 g19464(.A(new_n21806), .B(new_n21812), .Y(new_n21813));
  nand_5 g19465(.A(new_n21813), .B(new_n21683), .Y(new_n21814));
  or_6   g19466(.A(new_n21814), .B(new_n21811), .Y(new_n21815));
  nor_5  g19467(.A(new_n21809), .B(new_n12552), .Y(new_n21816));
  nand_5 g19468(.A(new_n21811), .B(new_n21682), .Y(new_n21817));
  nand_5 g19469(.A(new_n21817), .B(new_n21816), .Y(new_n21818));
  and_6  g19470(.A(new_n21818), .B(new_n21815), .Y(po0427));
  nand_5 g19471(.A(new_n7530), .B(pi663), .Y(new_n21820));
  nand_5 g19472(.A(new_n17493), .B(new_n17485), .Y(new_n21821));
  nand_5 g19473(.A(new_n21821), .B(new_n21820), .Y(new_n21822));
  nand_5 g19474(.A(new_n21822), .B(new_n20011), .Y(new_n21823));
  not_8  g19475(.A(new_n21823), .Y(new_n21824));
  xor_4  g19476(.A(new_n21822), .B(new_n20011), .Y(new_n21825));
  not_8  g19477(.A(new_n21825), .Y(new_n21826));
  nand_5 g19478(.A(new_n20014), .B(new_n17523), .Y(new_n21827));
  or_6   g19479(.A(new_n17531), .B(new_n17494), .Y(new_n21828));
  nand_5 g19480(.A(new_n21828), .B(new_n21827), .Y(new_n21829));
  nor_5  g19481(.A(new_n21829), .B(new_n21826), .Y(new_n21830));
  nor_5  g19482(.A(new_n21830), .B(new_n21824), .Y(new_n21831));
  not_8  g19483(.A(new_n21831), .Y(new_n21832));
  nand_5 g19484(.A(new_n17558), .B(new_n17533), .Y(new_n21833));
  nand_5 g19485(.A(new_n21833), .B(new_n17534), .Y(new_n21834));
  nor_5  g19486(.A(new_n21834), .B(new_n21832), .Y(new_n21835));
  xor_4  g19487(.A(new_n21834), .B(new_n21831), .Y(new_n21836));
  xor_4  g19488(.A(new_n21829), .B(new_n21826), .Y(new_n21837));
  not_8  g19489(.A(new_n21837), .Y(new_n21838));
  nand_5 g19490(.A(new_n21838), .B(new_n21834), .Y(new_n21839));
  not_8  g19491(.A(new_n21834), .Y(new_n21840));
  xor_4  g19492(.A(new_n21837), .B(new_n21840), .Y(new_n21841));
  or_6   g19493(.A(new_n17559), .B(new_n17532), .Y(new_n21842));
  nand_5 g19494(.A(new_n17608), .B(new_n17560), .Y(new_n21843));
  nand_5 g19495(.A(new_n21843), .B(new_n21842), .Y(new_n21844));
  nand_5 g19496(.A(new_n21844), .B(new_n21841), .Y(new_n21845));
  nand_5 g19497(.A(new_n21845), .B(new_n21839), .Y(new_n21846));
  not_8  g19498(.A(new_n21846), .Y(new_n21847));
  nor_5  g19499(.A(new_n21847), .B(new_n21836), .Y(new_n21848));
  nor_5  g19500(.A(new_n21848), .B(new_n21835), .Y(po0428));
  nand_5 g19501(.A(new_n10210), .B(new_n10193), .Y(new_n21850));
  nand_5 g19502(.A(new_n10222), .B(new_n10221), .Y(new_n21851));
  nand_5 g19503(.A(new_n21851), .B(new_n21850), .Y(po0429));
  nand_5 g19504(.A(new_n9210), .B(pi108), .Y(new_n21853));
  xor_4  g19505(.A(pi341), .B(new_n10965), .Y(new_n21854));
  nand_5 g19506(.A(pi442), .B(new_n9213), .Y(new_n21855));
  xor_4  g19507(.A(pi442), .B(new_n9213), .Y(new_n21856));
  nand_5 g19508(.A(pi462), .B(new_n9217), .Y(new_n21857));
  nand_5 g19509(.A(new_n19739), .B(new_n19727), .Y(new_n21858));
  nand_5 g19510(.A(new_n21858), .B(new_n21857), .Y(new_n21859));
  nand_5 g19511(.A(new_n21859), .B(new_n21856), .Y(new_n21860));
  nand_5 g19512(.A(new_n21860), .B(new_n21855), .Y(new_n21861));
  nand_5 g19513(.A(new_n21861), .B(new_n21854), .Y(new_n21862));
  nand_5 g19514(.A(new_n21862), .B(new_n21853), .Y(new_n21863));
  xor_4  g19515(.A(new_n21863), .B(new_n9208), .Y(new_n21864));
  xnor_4 g19516(.A(new_n21861), .B(new_n21854), .Y(new_n21865));
  nor_5  g19517(.A(new_n21865), .B(new_n9163), .Y(new_n21866));
  xor_4  g19518(.A(new_n21865), .B(new_n17308), .Y(new_n21867));
  xnor_4 g19519(.A(new_n21859), .B(new_n21856), .Y(new_n21868));
  nand_5 g19520(.A(new_n21868), .B(new_n9150), .Y(new_n21869));
  or_6   g19521(.A(new_n21868), .B(new_n9150), .Y(new_n21870));
  not_8  g19522(.A(new_n19740), .Y(new_n21871));
  nor_5  g19523(.A(new_n19756), .B(new_n21871), .Y(new_n21872));
  nor_5  g19524(.A(new_n19757), .B(new_n9138), .Y(new_n21873));
  nor_5  g19525(.A(new_n21873), .B(new_n21872), .Y(new_n21874));
  nand_5 g19526(.A(new_n21874), .B(new_n21870), .Y(new_n21875));
  nand_5 g19527(.A(new_n21875), .B(new_n21869), .Y(new_n21876));
  nor_5  g19528(.A(new_n21876), .B(new_n21867), .Y(new_n21877));
  or_6   g19529(.A(new_n21877), .B(new_n21866), .Y(new_n21878));
  nand_5 g19530(.A(new_n21878), .B(new_n21864), .Y(new_n21879));
  xnor_4 g19531(.A(new_n21878), .B(new_n21864), .Y(new_n21880));
  or_6   g19532(.A(new_n21880), .B(new_n9069), .Y(new_n21881));
  nand_5 g19533(.A(new_n21881), .B(new_n21879), .Y(new_n21882));
  nand_5 g19534(.A(new_n21882), .B(new_n9068), .Y(new_n21883));
  or_6   g19535(.A(new_n21882), .B(new_n9068), .Y(new_n21884));
  nand_5 g19536(.A(new_n21884), .B(new_n21883), .Y(new_n21885));
  nand_5 g19537(.A(new_n21863), .B(new_n9208), .Y(new_n21886));
  nand_5 g19538(.A(new_n21886), .B(new_n19612), .Y(new_n21887));
  not_8  g19539(.A(new_n21887), .Y(new_n21888));
  xor_4  g19540(.A(new_n21888), .B(new_n21885), .Y(po0430));
  xor_4  g19541(.A(new_n19081), .B(new_n16507), .Y(po0431));
  nor_5  g19542(.A(new_n19554), .B(new_n19539), .Y(new_n21891));
  nor_5  g19543(.A(new_n19588), .B(new_n19556), .Y(new_n21892));
  nor_5  g19544(.A(new_n21892), .B(new_n21891), .Y(po0432));
  xor_4  g19545(.A(new_n17000), .B(new_n12016), .Y(po0433));
  not_8  g19546(.A(pi142), .Y(new_n21895));
  nand_5 g19547(.A(pi293), .B(new_n21895), .Y(new_n21896));
  nand_5 g19548(.A(new_n3697), .B(pi142), .Y(new_n21897));
  nand_5 g19549(.A(new_n11349), .B(pi446), .Y(new_n21898));
  xor_4  g19550(.A(pi721), .B(new_n3525), .Y(new_n21899));
  nand_5 g19551(.A(pi507), .B(new_n11345), .Y(new_n21900));
  xor_4  g19552(.A(pi507), .B(new_n11345), .Y(new_n21901));
  nand_5 g19553(.A(new_n11294), .B(pi324), .Y(new_n21902));
  nand_5 g19554(.A(new_n2500), .B(new_n2469), .Y(new_n21903));
  nand_5 g19555(.A(new_n21903), .B(new_n21902), .Y(new_n21904));
  nand_5 g19556(.A(new_n21904), .B(new_n21901), .Y(new_n21905));
  nand_5 g19557(.A(new_n21905), .B(new_n21900), .Y(new_n21906));
  nand_5 g19558(.A(new_n21906), .B(new_n21899), .Y(new_n21907));
  nand_5 g19559(.A(new_n21907), .B(new_n21898), .Y(new_n21908));
  nand_5 g19560(.A(new_n21908), .B(new_n21897), .Y(new_n21909));
  nand_5 g19561(.A(new_n21909), .B(new_n21896), .Y(new_n21910));
  not_8  g19562(.A(new_n21910), .Y(new_n21911));
  xor_4  g19563(.A(new_n21911), .B(new_n7587), .Y(new_n21912));
  and_6  g19564(.A(new_n21912), .B(new_n7581), .Y(new_n21913));
  nor_5  g19565(.A(new_n21911), .B(new_n7587), .Y(new_n21914));
  nor_5  g19566(.A(new_n21914), .B(new_n7581), .Y(new_n21915));
  nor_5  g19567(.A(new_n21911), .B(new_n7580), .Y(new_n21916));
  nor_5  g19568(.A(new_n21916), .B(new_n21915), .Y(new_n21917));
  nand_5 g19569(.A(new_n21897), .B(new_n21896), .Y(new_n21918));
  xnor_4 g19570(.A(new_n21918), .B(new_n21908), .Y(new_n21919));
  or_6   g19571(.A(new_n21919), .B(new_n7588), .Y(new_n21920));
  xor_4  g19572(.A(new_n21919), .B(new_n7588), .Y(new_n21921));
  xor_4  g19573(.A(new_n21906), .B(new_n21899), .Y(new_n21922));
  or_6   g19574(.A(new_n21922), .B(new_n7630), .Y(new_n21923));
  xor_4  g19575(.A(new_n21922), .B(new_n7630), .Y(new_n21924));
  xor_4  g19576(.A(new_n21904), .B(new_n21901), .Y(new_n21925));
  or_6   g19577(.A(new_n21925), .B(new_n7633), .Y(new_n21926));
  xor_4  g19578(.A(new_n21925), .B(new_n7633), .Y(new_n21927));
  or_6   g19579(.A(new_n2501), .B(new_n2467), .Y(new_n21928));
  nand_5 g19580(.A(new_n2550), .B(new_n2502), .Y(new_n21929));
  nand_5 g19581(.A(new_n21929), .B(new_n21928), .Y(new_n21930));
  nand_5 g19582(.A(new_n21930), .B(new_n21927), .Y(new_n21931));
  nand_5 g19583(.A(new_n21931), .B(new_n21926), .Y(new_n21932));
  nand_5 g19584(.A(new_n21932), .B(new_n21924), .Y(new_n21933));
  nand_5 g19585(.A(new_n21933), .B(new_n21923), .Y(new_n21934));
  nand_5 g19586(.A(new_n21934), .B(new_n21921), .Y(new_n21935));
  nand_5 g19587(.A(new_n21935), .B(new_n21920), .Y(new_n21936));
  nor_5  g19588(.A(new_n21936), .B(new_n21917), .Y(new_n21937));
  nand_5 g19589(.A(new_n21911), .B(new_n7585), .Y(new_n21938));
  nand_5 g19590(.A(new_n21938), .B(new_n21936), .Y(new_n21939));
  nor_5  g19591(.A(new_n21939), .B(new_n21916), .Y(new_n21940));
  nor_5  g19592(.A(new_n21940), .B(new_n21937), .Y(new_n21941));
  nor_5  g19593(.A(new_n21941), .B(new_n21913), .Y(po0434));
  xor_4  g19594(.A(new_n7658), .B(new_n2527), .Y(po0435));
  not_8  g19595(.A(new_n2990), .Y(new_n21944));
  nand_5 g19596(.A(new_n2994), .B(pi822), .Y(new_n21945));
  xor_4  g19597(.A(new_n2994), .B(pi822), .Y(new_n21946));
  nand_5 g19598(.A(new_n18473), .B(pi100), .Y(new_n21947));
  nand_5 g19599(.A(new_n21947), .B(new_n18472), .Y(new_n21948));
  nand_5 g19600(.A(new_n21948), .B(new_n21946), .Y(new_n21949));
  nand_5 g19601(.A(new_n21949), .B(new_n21945), .Y(new_n21950));
  xor_4  g19602(.A(new_n21950), .B(new_n21944), .Y(new_n21951));
  xor_4  g19603(.A(new_n21951), .B(pi439), .Y(new_n21952));
  xor_4  g19604(.A(new_n21948), .B(new_n21946), .Y(new_n21953));
  not_8  g19605(.A(new_n18475), .Y(new_n21954));
  nor_5  g19606(.A(new_n21954), .B(new_n18468), .Y(new_n21955));
  or_6   g19607(.A(new_n18476), .B(new_n6882), .Y(new_n21956));
  not_8  g19608(.A(new_n21956), .Y(new_n21957));
  nor_5  g19609(.A(new_n21957), .B(new_n21955), .Y(new_n21958));
  or_6   g19610(.A(new_n21958), .B(new_n21953), .Y(new_n21959));
  not_8  g19611(.A(new_n21953), .Y(new_n21960));
  xor_4  g19612(.A(new_n21958), .B(new_n21960), .Y(new_n21961));
  or_6   g19613(.A(new_n21961), .B(new_n16316), .Y(new_n21962));
  nand_5 g19614(.A(new_n21962), .B(new_n21959), .Y(new_n21963));
  xor_4  g19615(.A(new_n21963), .B(new_n21952), .Y(new_n21964));
  xor_4  g19616(.A(new_n21964), .B(new_n6873), .Y(po0436));
  xor_4  g19617(.A(new_n17789), .B(new_n12234), .Y(po0437));
  xnor_4 g19618(.A(new_n3880), .B(new_n3879), .Y(po0438));
  xor_4  g19619(.A(new_n11814), .B(new_n11819), .Y(po0439));
  xor_4  g19620(.A(new_n15023), .B(new_n14984), .Y(po0440));
  xnor_4 g19621(.A(new_n19077), .B(new_n16513), .Y(po0441));
  xnor_4 g19622(.A(new_n20163), .B(new_n20162), .Y(po0442));
  nand_5 g19623(.A(new_n2980), .B(new_n7533), .Y(new_n21972));
  xor_4  g19624(.A(new_n2980), .B(new_n7533), .Y(new_n21973));
  nand_5 g19625(.A(new_n21950), .B(new_n21944), .Y(new_n21974));
  nand_5 g19626(.A(new_n21951), .B(pi439), .Y(new_n21975));
  nand_5 g19627(.A(new_n21975), .B(new_n21974), .Y(new_n21976));
  or_6   g19628(.A(new_n21976), .B(new_n15268), .Y(new_n21977));
  xor_4  g19629(.A(new_n21976), .B(new_n15268), .Y(new_n21978));
  nand_5 g19630(.A(new_n21978), .B(new_n7751), .Y(new_n21979));
  nand_5 g19631(.A(new_n21979), .B(new_n21977), .Y(new_n21980));
  nand_5 g19632(.A(new_n21980), .B(new_n21973), .Y(new_n21981));
  nand_5 g19633(.A(new_n21981), .B(new_n21972), .Y(new_n21982));
  nand_5 g19634(.A(new_n21982), .B(new_n18389), .Y(new_n21983));
  not_8  g19635(.A(new_n21983), .Y(new_n21984));
  nor_5  g19636(.A(new_n21982), .B(new_n18389), .Y(new_n21985));
  nor_5  g19637(.A(new_n21985), .B(pi697), .Y(new_n21986));
  nor_5  g19638(.A(new_n21986), .B(new_n21984), .Y(new_n21987));
  not_8  g19639(.A(new_n21987), .Y(new_n21988));
  nor_5  g19640(.A(new_n21985), .B(new_n21984), .Y(new_n21989));
  xor_4  g19641(.A(new_n21989), .B(new_n7530), .Y(new_n21990));
  xor_4  g19642(.A(new_n21980), .B(new_n21973), .Y(new_n21991));
  xor_4  g19643(.A(new_n21978), .B(new_n7751), .Y(new_n21992));
  nand_5 g19644(.A(new_n21992), .B(new_n6797), .Y(new_n21993));
  not_8  g19645(.A(new_n21963), .Y(new_n21994));
  nor_5  g19646(.A(new_n21994), .B(new_n21952), .Y(new_n21995));
  or_6   g19647(.A(new_n21964), .B(new_n6873), .Y(new_n21996));
  not_8  g19648(.A(new_n21996), .Y(new_n21997));
  nor_5  g19649(.A(new_n21997), .B(new_n21995), .Y(new_n21998));
  xor_4  g19650(.A(new_n21992), .B(new_n6796), .Y(new_n21999));
  or_6   g19651(.A(new_n21999), .B(new_n21998), .Y(new_n22000));
  nand_5 g19652(.A(new_n22000), .B(new_n21993), .Y(new_n22001));
  nand_5 g19653(.A(new_n22001), .B(new_n21991), .Y(new_n22002));
  xor_4  g19654(.A(new_n22001), .B(new_n21991), .Y(new_n22003));
  nand_5 g19655(.A(new_n22003), .B(new_n6939), .Y(new_n22004));
  nand_5 g19656(.A(new_n22004), .B(new_n22002), .Y(new_n22005));
  nor_5  g19657(.A(new_n22005), .B(new_n21990), .Y(new_n22006));
  xnor_4 g19658(.A(new_n22005), .B(new_n21990), .Y(new_n22007));
  nor_5  g19659(.A(new_n22007), .B(new_n17354), .Y(new_n22008));
  nor_5  g19660(.A(new_n22008), .B(new_n22006), .Y(new_n22009));
  nor_5  g19661(.A(new_n22009), .B(new_n21988), .Y(new_n22010));
  nand_5 g19662(.A(new_n22010), .B(new_n15264), .Y(new_n22011));
  nor_5  g19663(.A(new_n21988), .B(new_n15265), .Y(new_n22012));
  nand_5 g19664(.A(new_n22012), .B(new_n17352), .Y(new_n22013));
  not_8  g19665(.A(new_n22009), .Y(new_n22014));
  nand_5 g19666(.A(new_n21988), .B(new_n15265), .Y(new_n22015));
  nor_5  g19667(.A(new_n22015), .B(new_n22014), .Y(new_n22016));
  nor_5  g19668(.A(new_n22016), .B(new_n17350), .Y(new_n22017));
  nand_5 g19669(.A(new_n22017), .B(new_n22011), .Y(new_n22018));
  or_6   g19670(.A(new_n22010), .B(new_n17352), .Y(new_n22019));
  or_6   g19671(.A(new_n22019), .B(new_n22016), .Y(new_n22020));
  xor_4  g19672(.A(new_n21987), .B(new_n15265), .Y(new_n22021));
  nor_5  g19673(.A(new_n22021), .B(new_n22009), .Y(new_n22022));
  nor_5  g19674(.A(new_n22022), .B(new_n17351), .Y(new_n22023));
  nand_5 g19675(.A(new_n22023), .B(new_n22020), .Y(new_n22024));
  nand_5 g19676(.A(new_n22024), .B(new_n22018), .Y(new_n22025));
  nand_5 g19677(.A(new_n22025), .B(new_n22013), .Y(po1400));
  nand_5 g19678(.A(po1400), .B(new_n17350), .Y(new_n22027));
  nand_5 g19679(.A(new_n22027), .B(new_n22011), .Y(po0443));
  xor_4  g19680(.A(pi569), .B(pi390), .Y(new_n22029));
  xor_4  g19681(.A(new_n22029), .B(new_n7427), .Y(po0444));
  xor_4  g19682(.A(new_n7966), .B(new_n7965), .Y(po0445));
  xor_4  g19683(.A(new_n12630), .B(new_n12629), .Y(po0446));
  xnor_4 g19684(.A(new_n16571), .B(new_n10551), .Y(po0447));
  xnor_4 g19685(.A(new_n9151), .B(new_n9150), .Y(po0448));
  xor_4  g19686(.A(new_n9806), .B(new_n9449), .Y(po0449));
  xor_4  g19687(.A(new_n14582), .B(new_n3636), .Y(po0450));
  xor_4  g19688(.A(new_n13098), .B(new_n6043), .Y(po0451));
  nand_5 g19689(.A(new_n10424), .B(new_n10419), .Y(new_n22038));
  not_8  g19690(.A(new_n22038), .Y(new_n22039));
  nand_5 g19691(.A(new_n22039), .B(new_n10397), .Y(new_n22040));
  not_8  g19692(.A(new_n10421), .Y(new_n22041));
  nand_5 g19693(.A(new_n22041), .B(new_n10398), .Y(new_n22042));
  nand_5 g19694(.A(new_n22042), .B(new_n22040), .Y(po0452));
  xor_4  g19695(.A(new_n20603), .B(new_n15837), .Y(po0453));
  xor_4  g19696(.A(new_n16736), .B(new_n6225), .Y(po0454));
  xor_4  g19697(.A(new_n21934), .B(new_n21921), .Y(po0455));
  nand_5 g19698(.A(new_n19854), .B(new_n19850), .Y(new_n22047));
  not_8  g19699(.A(new_n22047), .Y(new_n22048));
  nor_5  g19700(.A(new_n19861), .B(new_n19851), .Y(new_n22049));
  nor_5  g19701(.A(new_n22049), .B(new_n22048), .Y(new_n22050));
  not_8  g19702(.A(new_n19828), .Y(new_n22051));
  nor_5  g19703(.A(new_n19858), .B(new_n19853), .Y(new_n22052));
  nand_5 g19704(.A(new_n22052), .B(new_n22048), .Y(new_n22053));
  nand_5 g19705(.A(new_n22053), .B(new_n22051), .Y(new_n22054));
  nor_5  g19706(.A(new_n22054), .B(new_n22050), .Y(new_n22055));
  and_6  g19707(.A(new_n19855), .B(new_n19828), .Y(new_n22056));
  nand_5 g19708(.A(new_n22056), .B(new_n19859), .Y(new_n22057));
  nor_5  g19709(.A(new_n22057), .B(new_n22049), .Y(new_n22058));
  nor_5  g19710(.A(new_n22058), .B(new_n22055), .Y(po0456));
  xor_4  g19711(.A(new_n12258), .B(new_n8703), .Y(po0457));
  nor_5  g19712(.A(new_n9812), .B(new_n9811), .Y(new_n22061));
  xor_4  g19713(.A(new_n22061), .B(new_n9813), .Y(po0458));
  xor_4  g19714(.A(new_n19575), .B(new_n19574), .Y(po0459));
  xor_4  g19715(.A(new_n20803), .B(new_n20794), .Y(po0460));
  xor_4  g19716(.A(new_n13517), .B(new_n9682), .Y(po0461));
  xnor_4 g19717(.A(new_n6918), .B(new_n6916), .Y(po0462));
  xor_4  g19718(.A(new_n2566), .B(pi702), .Y(new_n22067));
  xor_4  g19719(.A(new_n22067), .B(new_n4468), .Y(po0463));
  xor_4  g19720(.A(new_n7490), .B(new_n7489), .Y(po0464));
  xor_4  g19721(.A(new_n17375), .B(new_n17373), .Y(po0465));
  xor_4  g19722(.A(new_n19122), .B(new_n19112), .Y(po0466));
  xnor_4 g19723(.A(new_n7961), .B(new_n7960), .Y(po0467));
  not_8  g19724(.A(new_n17624), .Y(new_n22073));
  nor_5  g19725(.A(new_n17653), .B(new_n22073), .Y(new_n22074));
  nor_5  g19726(.A(new_n17654), .B(new_n16390), .Y(new_n22075));
  or_6   g19727(.A(new_n22075), .B(new_n22074), .Y(new_n22076));
  nor_5  g19728(.A(new_n22076), .B(new_n21735), .Y(new_n22077));
  xor_4  g19729(.A(new_n22076), .B(new_n21736), .Y(new_n22078));
  nor_5  g19730(.A(new_n22078), .B(new_n16442), .Y(new_n22079));
  or_6   g19731(.A(new_n22079), .B(new_n22077), .Y(new_n22080));
  nor_5  g19732(.A(new_n22080), .B(new_n21746), .Y(new_n22081));
  xor_4  g19733(.A(new_n22080), .B(new_n21745), .Y(new_n22082));
  nor_5  g19734(.A(new_n22082), .B(new_n21614), .Y(new_n22083));
  or_6   g19735(.A(new_n22083), .B(new_n22081), .Y(new_n22084));
  nor_5  g19736(.A(new_n21612), .B(new_n21608), .Y(new_n22085));
  nand_5 g19737(.A(new_n22085), .B(new_n18031), .Y(new_n22086));
  nand_5 g19738(.A(new_n18026), .B(pi124), .Y(new_n22087));
  nand_5 g19739(.A(new_n22087), .B(new_n22086), .Y(new_n22088));
  nand_5 g19740(.A(new_n18036), .B(new_n4873), .Y(new_n22089));
  nor_5  g19741(.A(new_n18036), .B(new_n4873), .Y(new_n22090));
  nor_5  g19742(.A(new_n22090), .B(new_n18031), .Y(new_n22091));
  nand_5 g19743(.A(new_n22091), .B(new_n21608), .Y(new_n22092));
  nand_5 g19744(.A(new_n22092), .B(new_n22089), .Y(new_n22093));
  nor_5  g19745(.A(new_n22093), .B(new_n22088), .Y(new_n22094));
  nand_5 g19746(.A(new_n21743), .B(new_n4858), .Y(new_n22095));
  nand_5 g19747(.A(new_n22095), .B(new_n15542), .Y(new_n22096));
  nand_5 g19748(.A(new_n21742), .B(pi315), .Y(new_n22097));
  not_8  g19749(.A(new_n22097), .Y(new_n22098));
  nand_5 g19750(.A(new_n22098), .B(new_n15548), .Y(new_n22099));
  nand_5 g19751(.A(new_n22099), .B(new_n22096), .Y(new_n22100));
  nand_5 g19752(.A(new_n22097), .B(new_n15553), .Y(new_n22101));
  not_8  g19753(.A(new_n22101), .Y(new_n22102));
  nor_5  g19754(.A(new_n22095), .B(new_n15548), .Y(new_n22103));
  nor_5  g19755(.A(new_n22103), .B(new_n22102), .Y(new_n22104));
  not_8  g19756(.A(new_n22104), .Y(new_n22105));
  nor_5  g19757(.A(new_n22105), .B(new_n22100), .Y(new_n22106));
  xor_4  g19758(.A(new_n22106), .B(new_n22094), .Y(new_n22107));
  xnor_4 g19759(.A(new_n22107), .B(new_n22084), .Y(po0468));
  nand_5 g19760(.A(pi430), .B(pi403), .Y(new_n22109));
  not_8  g19761(.A(new_n22109), .Y(new_n22110));
  nor_5  g19762(.A(new_n20671), .B(new_n20652), .Y(new_n22111));
  nor_5  g19763(.A(new_n22111), .B(new_n22110), .Y(new_n22112));
  nand_5 g19764(.A(pi512), .B(pi142), .Y(new_n22113));
  nand_5 g19765(.A(new_n16063), .B(new_n16044), .Y(new_n22114));
  nand_5 g19766(.A(new_n22114), .B(new_n22113), .Y(new_n22115));
  xor_4  g19767(.A(new_n22115), .B(new_n22112), .Y(new_n22116));
  not_8  g19768(.A(new_n22116), .Y(new_n22117));
  nand_5 g19769(.A(new_n20672), .B(new_n16065), .Y(new_n22118));
  or_6   g19770(.A(new_n20694), .B(new_n20674), .Y(new_n22119));
  nand_5 g19771(.A(new_n22119), .B(new_n22118), .Y(new_n22120));
  xor_4  g19772(.A(new_n22120), .B(new_n22117), .Y(new_n22121));
  nand_5 g19773(.A(new_n21382), .B(new_n7789), .Y(new_n22122));
  or_6   g19774(.A(new_n21383), .B(new_n20695), .Y(new_n22123));
  nand_5 g19775(.A(new_n22123), .B(new_n22122), .Y(new_n22124));
  xor_4  g19776(.A(new_n22124), .B(new_n22121), .Y(new_n22125));
  xor_4  g19777(.A(new_n22125), .B(new_n7745), .Y(po0469));
  nand_5 g19778(.A(new_n18392), .B(new_n16066), .Y(new_n22127));
  or_6   g19779(.A(new_n21645), .B(new_n21643), .Y(new_n22128));
  nand_5 g19780(.A(new_n22128), .B(new_n22127), .Y(new_n22129));
  xor_4  g19781(.A(new_n22129), .B(new_n18388), .Y(new_n22130));
  nand_5 g19782(.A(new_n22130), .B(new_n22094), .Y(new_n22131));
  nand_5 g19783(.A(new_n21646), .B(new_n21642), .Y(new_n22132));
  nand_5 g19784(.A(new_n21647), .B(new_n21613), .Y(new_n22133));
  nand_5 g19785(.A(new_n22133), .B(new_n22132), .Y(new_n22134));
  xor_4  g19786(.A(new_n22130), .B(new_n22094), .Y(new_n22135));
  nand_5 g19787(.A(new_n22135), .B(new_n22134), .Y(new_n22136));
  nand_5 g19788(.A(new_n22136), .B(new_n22131), .Y(new_n22137));
  not_8  g19789(.A(new_n22088), .Y(new_n22138));
  nor_5  g19790(.A(new_n22129), .B(new_n20746), .Y(new_n22139));
  xor_4  g19791(.A(new_n22139), .B(new_n22138), .Y(new_n22140));
  xnor_4 g19792(.A(new_n22140), .B(new_n22137), .Y(po0470));
  xnor_4 g19793(.A(new_n15773), .B(new_n15772), .Y(po0471));
  xor_4  g19794(.A(new_n17945), .B(new_n7916), .Y(po0472));
  xor_4  g19795(.A(new_n14000), .B(new_n12995), .Y(po0473));
  xor_4  g19796(.A(pi111), .B(pi072), .Y(new_n22145));
  nand_5 g19797(.A(new_n7181), .B(new_n16070), .Y(new_n22146));
  nand_5 g19798(.A(new_n20450), .B(new_n20447), .Y(new_n22147));
  nand_5 g19799(.A(new_n22147), .B(new_n22146), .Y(new_n22148));
  xor_4  g19800(.A(new_n22148), .B(new_n22145), .Y(new_n22149));
  xor_4  g19801(.A(new_n22149), .B(new_n7551), .Y(new_n22150));
  or_6   g19802(.A(new_n20452), .B(new_n7560), .Y(new_n22151));
  nand_5 g19803(.A(new_n20457), .B(new_n20453), .Y(new_n22152));
  nand_5 g19804(.A(new_n22152), .B(new_n22151), .Y(new_n22153));
  xor_4  g19805(.A(new_n22153), .B(new_n22150), .Y(new_n22154));
  xor_4  g19806(.A(pi689), .B(new_n3697), .Y(new_n22155));
  nand_5 g19807(.A(new_n20464), .B(new_n20461), .Y(new_n22156));
  nand_5 g19808(.A(new_n22156), .B(new_n20463), .Y(new_n22157));
  xor_4  g19809(.A(new_n22157), .B(new_n22155), .Y(new_n22158));
  xor_4  g19810(.A(new_n22158), .B(new_n22154), .Y(new_n22159));
  or_6   g19811(.A(new_n20466), .B(new_n20458), .Y(new_n22160));
  nand_5 g19812(.A(new_n20467), .B(new_n20446), .Y(new_n22161));
  nand_5 g19813(.A(new_n22161), .B(new_n22160), .Y(new_n22162));
  not_8  g19814(.A(new_n22162), .Y(new_n22163));
  xor_4  g19815(.A(new_n22163), .B(new_n22159), .Y(po0474));
  xor_4  g19816(.A(new_n13904), .B(new_n13903), .Y(po0475));
  nand_5 g19817(.A(new_n19313), .B(new_n19290), .Y(new_n22166));
  xor_4  g19818(.A(new_n22166), .B(new_n18496), .Y(po0476));
  xor_4  g19819(.A(new_n11845), .B(new_n11843), .Y(po0477));
  xnor_4 g19820(.A(new_n11285), .B(new_n11230), .Y(po0478));
  xor_4  g19821(.A(new_n21804), .B(new_n21655), .Y(po0479));
  xnor_4 g19822(.A(new_n5424), .B(new_n5405), .Y(po0480));
  xor_4  g19823(.A(new_n14605), .B(new_n14574), .Y(po0481));
  nand_5 g19824(.A(new_n20648), .B(new_n20627), .Y(new_n22173));
  not_8  g19825(.A(new_n22173), .Y(new_n22174));
  nor_5  g19826(.A(new_n20630), .B(new_n4278), .Y(new_n22175));
  xor_4  g19827(.A(new_n20641), .B(new_n22175), .Y(new_n22176));
  nand_5 g19828(.A(new_n22176), .B(new_n22174), .Y(new_n22177));
  nor_5  g19829(.A(new_n20647), .B(new_n20632), .Y(new_n22178));
  nor_5  g19830(.A(new_n22176), .B(new_n22178), .Y(new_n22179));
  nand_5 g19831(.A(new_n22179), .B(new_n22173), .Y(new_n22180));
  nand_5 g19832(.A(new_n22180), .B(new_n22177), .Y(po0482));
  xor_4  g19833(.A(new_n17602), .B(new_n17573), .Y(po0484));
  xnor_4 g19834(.A(new_n8286), .B(new_n8285), .Y(po0485));
  xor_4  g19835(.A(new_n15441), .B(new_n5068), .Y(po0486));
  nand_5 g19836(.A(new_n20991), .B(new_n20984), .Y(new_n22185));
  xor_4  g19837(.A(new_n22185), .B(new_n19804), .Y(new_n22186));
  nor_5  g19838(.A(new_n20973), .B(new_n20953), .Y(new_n22187));
  nand_5 g19839(.A(new_n20995), .B(new_n20974), .Y(new_n22188));
  not_8  g19840(.A(new_n22188), .Y(new_n22189));
  nor_5  g19841(.A(new_n22189), .B(new_n22187), .Y(new_n22190));
  xnor_4 g19842(.A(new_n22190), .B(new_n22186), .Y(po0487));
  xnor_4 g19843(.A(new_n19511), .B(new_n19510), .Y(po0488));
  xor_4  g19844(.A(new_n8703), .B(new_n6669), .Y(po0489));
  nand_5 g19845(.A(new_n12984), .B(new_n12978), .Y(new_n22194));
  xor_4  g19846(.A(new_n22194), .B(new_n12982), .Y(po0490));
  xor_4  g19847(.A(new_n18432), .B(new_n18419), .Y(po0491));
  xor_4  g19848(.A(new_n7162), .B(new_n7161), .Y(po0492));
  xor_4  g19849(.A(new_n11853), .B(new_n11852), .Y(po0493));
  xor_4  g19850(.A(new_n16485), .B(new_n5396), .Y(po0494));
  xnor_4 g19851(.A(new_n19498), .B(new_n19487), .Y(po0495));
  nand_5 g19852(.A(new_n16070), .B(pi452), .Y(new_n22201));
  nand_5 g19853(.A(new_n19133), .B(new_n19131), .Y(new_n22202));
  nand_5 g19854(.A(new_n22202), .B(new_n22201), .Y(new_n22203));
  xor_4  g19855(.A(pi697), .B(pi111), .Y(new_n22204));
  xor_4  g19856(.A(new_n22204), .B(new_n22203), .Y(new_n22205));
  and_6  g19857(.A(new_n22205), .B(new_n18425), .Y(new_n22206));
  xor_4  g19858(.A(new_n22205), .B(new_n18425), .Y(new_n22207));
  not_8  g19859(.A(new_n22207), .Y(new_n22208));
  not_8  g19860(.A(new_n19134), .Y(new_n22209));
  nor_5  g19861(.A(new_n22209), .B(new_n3045), .Y(new_n22210));
  nor_5  g19862(.A(new_n19135), .B(new_n19129), .Y(new_n22211));
  or_6   g19863(.A(new_n22211), .B(new_n22210), .Y(new_n22212));
  nor_5  g19864(.A(new_n22212), .B(new_n22208), .Y(new_n22213));
  nor_5  g19865(.A(new_n22213), .B(new_n22206), .Y(new_n22214));
  nand_5 g19866(.A(pi697), .B(new_n16066), .Y(new_n22215));
  not_8  g19867(.A(new_n22204), .Y(new_n22216));
  nand_5 g19868(.A(new_n22216), .B(new_n22203), .Y(new_n22217));
  nand_5 g19869(.A(new_n22217), .B(new_n22215), .Y(new_n22218));
  nand_5 g19870(.A(new_n22218), .B(new_n22214), .Y(new_n22219));
  nor_5  g19871(.A(new_n22218), .B(new_n22214), .Y(new_n22220));
  not_8  g19872(.A(new_n22220), .Y(new_n22221));
  and_6  g19873(.A(new_n22221), .B(new_n22219), .Y(new_n22222));
  xnor_4 g19874(.A(new_n22222), .B(new_n18417), .Y(po0496));
  xnor_4 g19875(.A(new_n14435), .B(new_n14418), .Y(po0497));
  xor_4  g19876(.A(new_n19017), .B(new_n4958), .Y(new_n22225));
  xor_4  g19877(.A(new_n22225), .B(new_n5010), .Y(po0498));
  xor_4  g19878(.A(new_n3659), .B(new_n3655), .Y(po0499));
  or_6   g19879(.A(new_n22221), .B(new_n18409), .Y(new_n22228));
  not_8  g19880(.A(new_n18403), .Y(new_n22229));
  nor_5  g19881(.A(new_n22219), .B(new_n18407), .Y(new_n22230));
  nand_5 g19882(.A(new_n22230), .B(new_n22229), .Y(new_n22231));
  nand_5 g19883(.A(new_n22231), .B(new_n22228), .Y(po0500));
  nor_5  g19884(.A(new_n10364), .B(new_n10246), .Y(new_n22233));
  xor_4  g19885(.A(new_n22233), .B(new_n10359), .Y(po0501));
  xor_4  g19886(.A(new_n21847), .B(new_n21836), .Y(po0502));
  xnor_4 g19887(.A(new_n12992), .B(new_n12951), .Y(po0503));
  xnor_4 g19888(.A(new_n21573), .B(new_n21572), .Y(po0504));
  xor_4  g19889(.A(new_n19125), .B(new_n19124), .Y(po0505));
  not_8  g19890(.A(new_n18761), .Y(new_n22239));
  nand_5 g19891(.A(new_n15993), .B(new_n15991), .Y(new_n22240));
  nand_5 g19892(.A(new_n22240), .B(new_n15992), .Y(new_n22241));
  nand_5 g19893(.A(new_n4374), .B(pi275), .Y(new_n22242));
  nand_5 g19894(.A(new_n22242), .B(new_n22241), .Y(new_n22243));
  nand_5 g19895(.A(pi368), .B(new_n14258), .Y(new_n22244));
  nand_5 g19896(.A(new_n22244), .B(new_n22243), .Y(new_n22245));
  xor_4  g19897(.A(new_n22245), .B(new_n22239), .Y(new_n22246));
  not_8  g19898(.A(new_n18803), .Y(new_n22247));
  xor_4  g19899(.A(new_n22241), .B(new_n22247), .Y(new_n22248));
  or_6   g19900(.A(new_n22248), .B(new_n17496), .Y(new_n22249));
  xor_4  g19901(.A(new_n22248), .B(new_n17496), .Y(new_n22250));
  nor_5  g19902(.A(new_n15987), .B(new_n15983), .Y(new_n22251));
  not_8  g19903(.A(new_n15995), .Y(new_n22252));
  nand_5 g19904(.A(new_n22252), .B(new_n15988), .Y(new_n22253));
  not_8  g19905(.A(new_n22253), .Y(new_n22254));
  nor_5  g19906(.A(new_n22254), .B(new_n22251), .Y(new_n22255));
  nand_5 g19907(.A(new_n22255), .B(new_n22250), .Y(new_n22256));
  nand_5 g19908(.A(new_n22256), .B(new_n22249), .Y(new_n22257));
  xor_4  g19909(.A(new_n22257), .B(new_n22246), .Y(new_n22258));
  xor_4  g19910(.A(new_n22258), .B(new_n17494), .Y(new_n22259));
  xor_4  g19911(.A(new_n22259), .B(new_n17559), .Y(new_n22260));
  xor_4  g19912(.A(new_n22255), .B(new_n22250), .Y(new_n22261));
  or_6   g19913(.A(new_n22261), .B(new_n17561), .Y(new_n22262));
  xor_4  g19914(.A(new_n22261), .B(new_n17561), .Y(new_n22263));
  not_8  g19915(.A(new_n15996), .Y(new_n22264));
  nor_5  g19916(.A(new_n17566), .B(new_n22264), .Y(new_n22265));
  xor_4  g19917(.A(new_n17566), .B(new_n15996), .Y(new_n22266));
  nand_5 g19918(.A(new_n17569), .B(new_n10799), .Y(new_n22267));
  not_8  g19919(.A(new_n10820), .Y(new_n22268));
  nand_5 g19920(.A(new_n17574), .B(new_n22268), .Y(new_n22269));
  nand_5 g19921(.A(new_n17580), .B(new_n10800), .Y(new_n22270));
  xor_4  g19922(.A(new_n17580), .B(new_n10800), .Y(new_n22271));
  or_6   g19923(.A(new_n15239), .B(new_n10802), .Y(new_n22272));
  nand_5 g19924(.A(new_n15254), .B(new_n15240), .Y(new_n22273));
  nand_5 g19925(.A(new_n22273), .B(new_n22272), .Y(new_n22274));
  nand_5 g19926(.A(new_n22274), .B(new_n22271), .Y(new_n22275));
  nand_5 g19927(.A(new_n22275), .B(new_n22270), .Y(new_n22276));
  xor_4  g19928(.A(new_n17574), .B(new_n10820), .Y(new_n22277));
  or_6   g19929(.A(new_n22277), .B(new_n22276), .Y(new_n22278));
  nand_5 g19930(.A(new_n22278), .B(new_n22269), .Y(new_n22279));
  xor_4  g19931(.A(new_n17569), .B(new_n10799), .Y(new_n22280));
  nand_5 g19932(.A(new_n22280), .B(new_n22279), .Y(new_n22281));
  and_6  g19933(.A(new_n22281), .B(new_n22267), .Y(new_n22282));
  nor_5  g19934(.A(new_n22282), .B(new_n22266), .Y(new_n22283));
  nor_5  g19935(.A(new_n22283), .B(new_n22265), .Y(new_n22284));
  nand_5 g19936(.A(new_n22284), .B(new_n22263), .Y(new_n22285));
  nand_5 g19937(.A(new_n22285), .B(new_n22262), .Y(new_n22286));
  xor_4  g19938(.A(new_n22286), .B(new_n22260), .Y(po0506));
  xor_4  g19939(.A(new_n16426), .B(new_n8575), .Y(po0507));
  not_8  g19940(.A(new_n19665), .Y(new_n22289));
  nor_5  g19941(.A(new_n22289), .B(new_n19657), .Y(new_n22290));
  nor_5  g19942(.A(new_n19676), .B(new_n19666), .Y(new_n22291));
  or_6   g19943(.A(new_n22291), .B(new_n22290), .Y(new_n22292));
  xor_4  g19944(.A(pi404), .B(new_n11899), .Y(new_n22293));
  not_8  g19945(.A(new_n22293), .Y(new_n22294));
  nand_5 g19946(.A(new_n2940), .B(pi239), .Y(new_n22295));
  not_8  g19947(.A(new_n22295), .Y(new_n22296));
  not_8  g19948(.A(new_n19658), .Y(new_n22297));
  nor_5  g19949(.A(new_n19664), .B(new_n22297), .Y(new_n22298));
  nor_5  g19950(.A(new_n22298), .B(new_n22296), .Y(new_n22299));
  xor_4  g19951(.A(new_n22299), .B(new_n22294), .Y(new_n22300));
  xor_4  g19952(.A(new_n22300), .B(new_n20458), .Y(new_n22301));
  xnor_4 g19953(.A(new_n22301), .B(new_n22292), .Y(po0508));
  nand_5 g19954(.A(new_n8981), .B(pi358), .Y(new_n22303));
  not_8  g19955(.A(new_n22303), .Y(new_n22304));
  nand_5 g19956(.A(pi397), .B(new_n10400), .Y(new_n22305));
  nand_5 g19957(.A(new_n22305), .B(new_n22303), .Y(new_n22306));
  nor_5  g19958(.A(new_n10266), .B(pi469), .Y(new_n22307));
  nor_5  g19959(.A(new_n15181), .B(new_n15161), .Y(new_n22308));
  nor_5  g19960(.A(new_n22308), .B(new_n22307), .Y(new_n22309));
  nor_5  g19961(.A(new_n22309), .B(new_n22306), .Y(new_n22310));
  nor_5  g19962(.A(new_n22310), .B(new_n22304), .Y(new_n22311));
  xor_4  g19963(.A(new_n22309), .B(new_n22306), .Y(new_n22312));
  nor_5  g19964(.A(new_n22312), .B(new_n21231), .Y(new_n22313));
  nor_5  g19965(.A(new_n15183), .B(new_n15159), .Y(new_n22314));
  nor_5  g19966(.A(new_n15217), .B(new_n15185), .Y(new_n22315));
  or_6   g19967(.A(new_n22315), .B(new_n22314), .Y(new_n22316));
  xor_4  g19968(.A(new_n22312), .B(new_n21232), .Y(new_n22317));
  nor_5  g19969(.A(new_n22317), .B(new_n22316), .Y(new_n22318));
  nor_5  g19970(.A(new_n22318), .B(new_n22313), .Y(new_n22319));
  not_8  g19971(.A(new_n22319), .Y(new_n22320));
  or_6   g19972(.A(new_n22320), .B(new_n22311), .Y(new_n22321));
  nand_5 g19973(.A(new_n22320), .B(new_n22311), .Y(new_n22322));
  and_6  g19974(.A(new_n22322), .B(new_n22321), .Y(new_n22323));
  xor_4  g19975(.A(new_n22323), .B(new_n21227), .Y(po0509));
  xnor_4 g19976(.A(new_n15409), .B(new_n15408), .Y(po0510));
  xor_4  g19977(.A(new_n12940), .B(new_n13988), .Y(new_n22326));
  xor_4  g19978(.A(new_n22326), .B(new_n12998), .Y(po0511));
  not_8  g19979(.A(new_n4463), .Y(new_n22328));
  xor_4  g19980(.A(new_n4472), .B(new_n22328), .Y(po0512));
  xor_4  g19981(.A(new_n11235), .B(new_n7250), .Y(po0513));
  nand_5 g19982(.A(new_n21438), .B(new_n21399), .Y(new_n22331));
  xor_4  g19983(.A(new_n22331), .B(new_n14582), .Y(po0514));
  xnor_4 g19984(.A(new_n8631), .B(new_n8630), .Y(po0515));
  xor_4  g19985(.A(new_n16937), .B(new_n16935), .Y(po0516));
  xor_4  g19986(.A(new_n4480), .B(new_n4456), .Y(po0517));
  nand_5 g19987(.A(new_n22245), .B(new_n22239), .Y(new_n22336));
  nand_5 g19988(.A(new_n22336), .B(new_n18759), .Y(new_n22337));
  nand_5 g19989(.A(new_n22337), .B(new_n21822), .Y(new_n22338));
  or_6   g19990(.A(new_n22337), .B(new_n21822), .Y(new_n22339));
  or_6   g19991(.A(new_n22257), .B(new_n22246), .Y(new_n22340));
  nand_5 g19992(.A(new_n22258), .B(new_n17495), .Y(new_n22341));
  nand_5 g19993(.A(new_n22341), .B(new_n22340), .Y(new_n22342));
  not_8  g19994(.A(new_n22342), .Y(new_n22343));
  nand_5 g19995(.A(new_n22343), .B(new_n22339), .Y(new_n22344));
  nand_5 g19996(.A(new_n22344), .B(new_n22338), .Y(new_n22345));
  nor_5  g19997(.A(new_n22345), .B(new_n5495), .Y(new_n22346));
  xor_4  g19998(.A(new_n22345), .B(new_n5495), .Y(new_n22347));
  not_8  g19999(.A(new_n22347), .Y(new_n22348));
  nand_5 g20000(.A(new_n22338), .B(new_n22339), .Y(new_n22349));
  xor_4  g20001(.A(new_n22349), .B(new_n22343), .Y(new_n22350));
  not_8  g20002(.A(new_n22350), .Y(new_n22351));
  or_6   g20003(.A(new_n16000), .B(new_n15996), .Y(new_n22352));
  nand_5 g20004(.A(new_n16001), .B(new_n10432), .Y(new_n22353));
  nand_5 g20005(.A(new_n22353), .B(new_n22352), .Y(new_n22354));
  nor_5  g20006(.A(new_n22354), .B(new_n10429), .Y(new_n22355));
  not_8  g20007(.A(new_n22261), .Y(new_n22356));
  xor_4  g20008(.A(new_n22354), .B(new_n5560), .Y(new_n22357));
  nor_5  g20009(.A(new_n22357), .B(new_n22356), .Y(new_n22358));
  or_6   g20010(.A(new_n22358), .B(new_n22355), .Y(new_n22359));
  nor_5  g20011(.A(new_n22359), .B(new_n22259), .Y(new_n22360));
  xor_4  g20012(.A(new_n22359), .B(new_n22259), .Y(new_n22361));
  nand_5 g20013(.A(new_n22361), .B(new_n10428), .Y(new_n22362));
  not_8  g20014(.A(new_n22362), .Y(new_n22363));
  nor_5  g20015(.A(new_n22363), .B(new_n22360), .Y(new_n22364));
  nand_5 g20016(.A(new_n22364), .B(new_n22351), .Y(new_n22365));
  xor_4  g20017(.A(new_n22364), .B(new_n22351), .Y(new_n22366));
  nand_5 g20018(.A(new_n22366), .B(new_n5496), .Y(new_n22367));
  nand_5 g20019(.A(new_n22367), .B(new_n22365), .Y(new_n22368));
  nor_5  g20020(.A(new_n22368), .B(new_n22348), .Y(new_n22369));
  nor_5  g20021(.A(new_n22369), .B(new_n22346), .Y(po0518));
  xor_4  g20022(.A(new_n19882), .B(new_n18041), .Y(po0519));
  xor_4  g20023(.A(new_n4988), .B(new_n4986), .Y(po0520));
  xnor_4 g20024(.A(new_n10946), .B(new_n10924), .Y(po0521));
  xnor_4 g20025(.A(new_n7679), .B(new_n7678), .Y(po0522));
  nand_5 g20026(.A(new_n16496), .B(new_n16456), .Y(new_n22375));
  nand_5 g20027(.A(new_n16497), .B(new_n17105), .Y(new_n22376));
  nand_5 g20028(.A(new_n22376), .B(new_n22375), .Y(new_n22377));
  xor_4  g20029(.A(new_n17022), .B(new_n17105), .Y(new_n22378));
  xnor_4 g20030(.A(new_n22378), .B(new_n22377), .Y(po0523));
  xor_4  g20031(.A(new_n13540), .B(new_n10007), .Y(po0524));
  xor_4  g20032(.A(new_n3371), .B(new_n3369), .Y(po0525));
  xnor_4 g20033(.A(new_n10089), .B(new_n10070), .Y(po0526));
  xor_4  g20034(.A(new_n13901), .B(new_n13899), .Y(po0527));
  xor_4  g20035(.A(new_n14061), .B(new_n13800), .Y(po0528));
  xor_4  g20036(.A(new_n21930), .B(new_n21927), .Y(po0529));
  xnor_4 g20037(.A(new_n16136), .B(new_n15481), .Y(po0530));
  xnor_4 g20038(.A(new_n6699), .B(new_n6698), .Y(po0531));
  nor_5  g20039(.A(new_n3329), .B(new_n3210), .Y(new_n22388));
  not_8  g20040(.A(new_n22388), .Y(new_n22389));
  not_8  g20041(.A(new_n18354), .Y(new_n22390));
  nand_5 g20042(.A(new_n6689), .B(new_n2472), .Y(new_n22391));
  nand_5 g20043(.A(new_n22391), .B(new_n6688), .Y(new_n22392));
  nand_5 g20044(.A(new_n22392), .B(new_n17045), .Y(new_n22393));
  or_6   g20045(.A(new_n22392), .B(new_n17045), .Y(new_n22394));
  nand_5 g20046(.A(new_n22394), .B(new_n2470), .Y(new_n22395));
  nand_5 g20047(.A(new_n22395), .B(new_n22393), .Y(new_n22396));
  or_6   g20048(.A(new_n22396), .B(new_n17071), .Y(new_n22397));
  xor_4  g20049(.A(new_n22396), .B(new_n17071), .Y(new_n22398));
  nand_5 g20050(.A(new_n22398), .B(pi348), .Y(new_n22399));
  nand_5 g20051(.A(new_n22399), .B(new_n22397), .Y(new_n22400));
  or_6   g20052(.A(new_n22400), .B(new_n17091), .Y(new_n22401));
  nand_5 g20053(.A(new_n22401), .B(pi417), .Y(new_n22402));
  nand_5 g20054(.A(new_n22400), .B(new_n17091), .Y(new_n22403));
  nand_5 g20055(.A(new_n22403), .B(new_n22402), .Y(new_n22404));
  or_6   g20056(.A(new_n22404), .B(new_n22390), .Y(new_n22405));
  xor_4  g20057(.A(new_n22404), .B(new_n22390), .Y(new_n22406));
  nand_5 g20058(.A(new_n22406), .B(new_n11349), .Y(new_n22407));
  nand_5 g20059(.A(new_n22407), .B(new_n22405), .Y(new_n22408));
  nand_5 g20060(.A(new_n22408), .B(new_n18346), .Y(new_n22409));
  nor_5  g20061(.A(new_n22408), .B(new_n18346), .Y(new_n22410));
  not_8  g20062(.A(new_n22410), .Y(new_n22411));
  nand_5 g20063(.A(new_n22411), .B(new_n22409), .Y(new_n22412));
  xor_4  g20064(.A(new_n22412), .B(new_n21895), .Y(new_n22413));
  xor_4  g20065(.A(new_n22406), .B(pi721), .Y(new_n22414));
  nor_5  g20066(.A(new_n6711), .B(new_n6691), .Y(new_n22415));
  nor_5  g20067(.A(new_n6712), .B(new_n3338), .Y(new_n22416));
  or_6   g20068(.A(new_n22416), .B(new_n22415), .Y(new_n22417));
  and_6  g20069(.A(new_n22394), .B(new_n22393), .Y(new_n22418));
  xor_4  g20070(.A(new_n22418), .B(new_n2470), .Y(new_n22419));
  not_8  g20071(.A(new_n22419), .Y(new_n22420));
  nor_5  g20072(.A(new_n22420), .B(new_n22417), .Y(new_n22421));
  xor_4  g20073(.A(new_n22419), .B(new_n22417), .Y(new_n22422));
  nor_5  g20074(.A(new_n22422), .B(new_n3336), .Y(new_n22423));
  or_6   g20075(.A(new_n22423), .B(new_n22421), .Y(new_n22424));
  xor_4  g20076(.A(new_n22398), .B(new_n11294), .Y(new_n22425));
  or_6   g20077(.A(new_n22425), .B(new_n22424), .Y(new_n22426));
  nand_5 g20078(.A(new_n22426), .B(new_n3389), .Y(new_n22427));
  nand_5 g20079(.A(new_n22425), .B(new_n22424), .Y(new_n22428));
  nand_5 g20080(.A(new_n22428), .B(new_n22427), .Y(new_n22429));
  nand_5 g20081(.A(new_n22403), .B(new_n22401), .Y(new_n22430));
  xor_4  g20082(.A(new_n22430), .B(pi417), .Y(new_n22431));
  nor_5  g20083(.A(new_n22431), .B(new_n22429), .Y(new_n22432));
  xnor_4 g20084(.A(new_n22431), .B(new_n22429), .Y(new_n22433));
  nor_5  g20085(.A(new_n22433), .B(new_n3393), .Y(new_n22434));
  or_6   g20086(.A(new_n22434), .B(new_n22432), .Y(new_n22435));
  nand_5 g20087(.A(new_n22435), .B(new_n22414), .Y(new_n22436));
  or_6   g20088(.A(new_n22435), .B(new_n22414), .Y(new_n22437));
  nand_5 g20089(.A(new_n22437), .B(new_n3406), .Y(new_n22438));
  nand_5 g20090(.A(new_n22438), .B(new_n22436), .Y(new_n22439));
  nor_5  g20091(.A(new_n22439), .B(new_n22413), .Y(new_n22440));
  nor_5  g20092(.A(new_n22440), .B(new_n22389), .Y(new_n22441));
  not_8  g20093(.A(new_n3260), .Y(new_n22442));
  nand_5 g20094(.A(new_n22439), .B(new_n22413), .Y(new_n22443));
  nor_5  g20095(.A(new_n22443), .B(new_n22442), .Y(new_n22444));
  nor_5  g20096(.A(new_n22444), .B(new_n22441), .Y(new_n22445));
  nor_5  g20097(.A(new_n3258), .B(new_n3211), .Y(new_n22446));
  or_6   g20098(.A(new_n22446), .B(new_n22440), .Y(new_n22447));
  not_8  g20099(.A(new_n22443), .Y(new_n22448));
  nor_5  g20100(.A(new_n22448), .B(new_n3260), .Y(new_n22449));
  nand_5 g20101(.A(new_n22449), .B(new_n22447), .Y(new_n22450));
  nand_5 g20102(.A(new_n22411), .B(new_n21895), .Y(new_n22451));
  nand_5 g20103(.A(new_n22451), .B(new_n22409), .Y(new_n22452));
  not_8  g20104(.A(new_n22452), .Y(new_n22453));
  xor_4  g20105(.A(new_n22453), .B(new_n18311), .Y(new_n22454));
  nand_5 g20106(.A(new_n22454), .B(new_n22450), .Y(new_n22455));
  nand_5 g20107(.A(new_n22455), .B(new_n22445), .Y(new_n22456));
  nor_5  g20108(.A(new_n22456), .B(new_n18302), .Y(new_n22457));
  nand_5 g20109(.A(new_n22452), .B(new_n18302), .Y(new_n22458));
  nand_5 g20110(.A(new_n22453), .B(new_n18310), .Y(new_n22459));
  nand_5 g20111(.A(new_n22459), .B(new_n22458), .Y(new_n22460));
  nand_5 g20112(.A(new_n22456), .B(new_n18302), .Y(new_n22461));
  nand_5 g20113(.A(new_n22461), .B(new_n22460), .Y(new_n22462));
  nor_5  g20114(.A(new_n22462), .B(new_n22457), .Y(po0532));
  nor_5  g20115(.A(new_n18321), .B(pi666), .Y(new_n22464));
  not_8  g20116(.A(new_n18327), .Y(new_n22465));
  nand_5 g20117(.A(new_n17101), .B(pi437), .Y(new_n22466));
  nand_5 g20118(.A(new_n17760), .B(new_n17102), .Y(new_n22467));
  nand_5 g20119(.A(new_n22467), .B(new_n22466), .Y(new_n22468));
  nor_5  g20120(.A(new_n22468), .B(new_n22465), .Y(new_n22469));
  nor_5  g20121(.A(new_n22469), .B(new_n22464), .Y(new_n22470));
  xor_4  g20122(.A(new_n22470), .B(new_n18349), .Y(new_n22471));
  xor_4  g20123(.A(new_n22306), .B(new_n13233), .Y(new_n22472));
  nand_5 g20124(.A(new_n5269), .B(new_n8796), .Y(new_n22473));
  xor_4  g20125(.A(new_n5269), .B(new_n8796), .Y(new_n22474));
  or_6   g20126(.A(new_n5318), .B(pi123), .Y(new_n22475));
  not_8  g20127(.A(new_n17804), .Y(new_n22476));
  nand_5 g20128(.A(new_n22476), .B(new_n17799), .Y(new_n22477));
  nand_5 g20129(.A(new_n22477), .B(new_n22475), .Y(new_n22478));
  nand_5 g20130(.A(new_n22478), .B(new_n22474), .Y(new_n22479));
  nand_5 g20131(.A(new_n22479), .B(new_n22473), .Y(new_n22480));
  xor_4  g20132(.A(new_n22480), .B(new_n22472), .Y(new_n22481));
  not_8  g20133(.A(new_n22481), .Y(new_n22482));
  or_6   g20134(.A(new_n22482), .B(new_n22471), .Y(new_n22483));
  nand_5 g20135(.A(new_n22482), .B(new_n22471), .Y(new_n22484));
  not_8  g20136(.A(new_n17805), .Y(new_n22485));
  nand_5 g20137(.A(new_n22485), .B(new_n17798), .Y(new_n22486));
  nand_5 g20138(.A(new_n17807), .B(new_n17761), .Y(new_n22487));
  nand_5 g20139(.A(new_n22487), .B(new_n22486), .Y(new_n22488));
  xor_4  g20140(.A(new_n22478), .B(new_n22474), .Y(new_n22489));
  nor_5  g20141(.A(new_n22489), .B(new_n22488), .Y(new_n22490));
  not_8  g20142(.A(new_n22489), .Y(new_n22491));
  xor_4  g20143(.A(new_n22491), .B(new_n22488), .Y(new_n22492));
  xor_4  g20144(.A(new_n22468), .B(new_n22465), .Y(new_n22493));
  nor_5  g20145(.A(new_n22493), .B(new_n22492), .Y(new_n22494));
  nor_5  g20146(.A(new_n22494), .B(new_n22490), .Y(new_n22495));
  not_8  g20147(.A(new_n22495), .Y(new_n22496));
  nand_5 g20148(.A(new_n22496), .B(new_n22484), .Y(new_n22497));
  nand_5 g20149(.A(new_n22497), .B(new_n22483), .Y(new_n22498));
  not_8  g20150(.A(new_n22498), .Y(new_n22499));
  nand_5 g20151(.A(new_n22470), .B(new_n18350), .Y(new_n22500));
  nor_5  g20152(.A(new_n22500), .B(new_n18369), .Y(new_n22501));
  nand_5 g20153(.A(new_n18335), .B(pi244), .Y(new_n22502));
  nand_5 g20154(.A(new_n18369), .B(new_n8986), .Y(new_n22503));
  and_6  g20155(.A(new_n22503), .B(new_n22502), .Y(new_n22504));
  or_6   g20156(.A(new_n22504), .B(new_n22470), .Y(new_n22505));
  nand_5 g20157(.A(new_n18339), .B(pi800), .Y(new_n22506));
  nand_5 g20158(.A(new_n22506), .B(new_n22502), .Y(new_n22507));
  nand_5 g20159(.A(new_n22507), .B(new_n18320), .Y(new_n22508));
  nand_5 g20160(.A(new_n22508), .B(new_n22505), .Y(new_n22509));
  nor_5  g20161(.A(new_n22509), .B(new_n22501), .Y(new_n22510));
  nor_5  g20162(.A(new_n22510), .B(new_n22499), .Y(new_n22511));
  nand_5 g20163(.A(new_n22510), .B(new_n18369), .Y(new_n22512));
  not_8  g20164(.A(new_n22512), .Y(new_n22513));
  nor_5  g20165(.A(new_n22513), .B(new_n22511), .Y(new_n22514));
  not_8  g20166(.A(new_n22305), .Y(new_n22515));
  nand_5 g20167(.A(new_n22515), .B(new_n13230), .Y(new_n22516));
  or_6   g20168(.A(new_n22306), .B(new_n13233), .Y(new_n22517));
  nand_5 g20169(.A(new_n22517), .B(new_n22305), .Y(new_n22518));
  nor_5  g20170(.A(new_n22480), .B(new_n13232), .Y(new_n22519));
  nand_5 g20171(.A(new_n22519), .B(new_n22518), .Y(new_n22520));
  nand_5 g20172(.A(new_n22520), .B(new_n22516), .Y(new_n22521));
  not_8  g20173(.A(new_n22521), .Y(new_n22522));
  nor_5  g20174(.A(new_n22522), .B(new_n22514), .Y(new_n22523));
  xor_4  g20175(.A(new_n22510), .B(new_n22499), .Y(new_n22524));
  nand_5 g20176(.A(new_n22304), .B(new_n13232), .Y(new_n22525));
  not_8  g20177(.A(new_n22525), .Y(new_n22526));
  not_8  g20178(.A(new_n16446), .Y(new_n22527));
  not_8  g20179(.A(new_n22472), .Y(new_n22528));
  nand_5 g20180(.A(new_n22480), .B(new_n22528), .Y(new_n22529));
  nor_5  g20181(.A(new_n22529), .B(new_n22527), .Y(new_n22530));
  nor_5  g20182(.A(new_n22530), .B(new_n22526), .Y(new_n22531));
  nand_5 g20183(.A(new_n22531), .B(new_n22522), .Y(new_n22532));
  nor_5  g20184(.A(new_n22532), .B(new_n22524), .Y(new_n22533));
  nand_5 g20185(.A(new_n22531), .B(new_n22513), .Y(new_n22534));
  nor_5  g20186(.A(new_n22534), .B(new_n22533), .Y(new_n22535));
  nor_5  g20187(.A(new_n22535), .B(new_n22521), .Y(new_n22536));
  nor_5  g20188(.A(new_n22536), .B(new_n22523), .Y(po0533));
  xnor_4 g20189(.A(new_n20043), .B(new_n20041), .Y(po0534));
  not_8  g20190(.A(new_n8113), .Y(new_n22539));
  nor_5  g20191(.A(new_n19593), .B(new_n8283), .Y(new_n22540));
  nor_5  g20192(.A(new_n19609), .B(new_n19595), .Y(new_n22541));
  nor_5  g20193(.A(new_n22541), .B(new_n22540), .Y(new_n22542));
  nand_5 g20194(.A(new_n19606), .B(new_n5546), .Y(new_n22543));
  nand_5 g20195(.A(new_n22543), .B(new_n19607), .Y(new_n22544));
  xor_4  g20196(.A(new_n22544), .B(new_n20927), .Y(new_n22545));
  xor_4  g20197(.A(new_n22545), .B(new_n8114), .Y(new_n22546));
  nor_5  g20198(.A(new_n22546), .B(new_n22542), .Y(new_n22547));
  not_8  g20199(.A(new_n22545), .Y(new_n22548));
  or_6   g20200(.A(new_n22548), .B(new_n8114), .Y(new_n22549));
  nor_5  g20201(.A(new_n22544), .B(new_n20927), .Y(new_n22550));
  xor_4  g20202(.A(new_n22550), .B(new_n8113), .Y(new_n22551));
  nand_5 g20203(.A(new_n22551), .B(new_n22549), .Y(new_n22552));
  nor_5  g20204(.A(new_n22552), .B(new_n22547), .Y(new_n22553));
  nor_5  g20205(.A(new_n22553), .B(new_n22539), .Y(po0535));
  xnor_4 g20206(.A(new_n18363), .B(new_n18362), .Y(po0536));
  nand_5 g20207(.A(new_n21250), .B(new_n21249), .Y(new_n22556));
  xnor_4 g20208(.A(new_n22556), .B(new_n21258), .Y(po0537));
  xor_4  g20209(.A(new_n18543), .B(new_n18542), .Y(po0538));
  xor_4  g20210(.A(new_n21345), .B(new_n18077), .Y(po0539));
  xor_4  g20211(.A(pi185), .B(pi093), .Y(new_n22560));
  nand_5 g20212(.A(new_n12002), .B(new_n4922), .Y(new_n22561));
  not_8  g20213(.A(new_n22561), .Y(new_n22562));
  nand_5 g20214(.A(pi752), .B(pi143), .Y(new_n22563));
  xor_4  g20215(.A(pi752), .B(pi143), .Y(new_n22564));
  nand_5 g20216(.A(pi676), .B(pi177), .Y(new_n22565));
  xor_4  g20217(.A(pi676), .B(pi177), .Y(new_n22566));
  not_8  g20218(.A(new_n22566), .Y(new_n22567));
  nand_5 g20219(.A(new_n4908), .B(new_n3846), .Y(new_n22568));
  nand_5 g20220(.A(new_n13183), .B(new_n13175), .Y(new_n22569));
  nand_5 g20221(.A(new_n22569), .B(new_n22568), .Y(new_n22570));
  or_6   g20222(.A(new_n22570), .B(new_n22567), .Y(new_n22571));
  nand_5 g20223(.A(new_n22571), .B(new_n22565), .Y(new_n22572));
  nand_5 g20224(.A(new_n22572), .B(new_n22564), .Y(new_n22573));
  nand_5 g20225(.A(new_n22573), .B(new_n22563), .Y(new_n22574));
  xor_4  g20226(.A(pi382), .B(new_n4922), .Y(new_n22575));
  nor_5  g20227(.A(new_n22575), .B(new_n22574), .Y(new_n22576));
  nor_5  g20228(.A(new_n22576), .B(new_n22562), .Y(new_n22577));
  not_8  g20229(.A(new_n22577), .Y(new_n22578));
  xor_4  g20230(.A(new_n22578), .B(new_n22560), .Y(new_n22579));
  xor_4  g20231(.A(new_n22579), .B(new_n4849), .Y(new_n22580));
  xor_4  g20232(.A(new_n22575), .B(new_n22574), .Y(new_n22581));
  nor_5  g20233(.A(new_n22581), .B(new_n4791), .Y(new_n22582));
  xor_4  g20234(.A(new_n22581), .B(new_n4790), .Y(new_n22583));
  xnor_4 g20235(.A(new_n22572), .B(new_n22564), .Y(new_n22584));
  nor_5  g20236(.A(new_n22584), .B(new_n4792), .Y(new_n22585));
  xor_4  g20237(.A(new_n22584), .B(new_n4792), .Y(new_n22586));
  not_8  g20238(.A(new_n22586), .Y(new_n22587));
  xor_4  g20239(.A(new_n22570), .B(new_n22566), .Y(new_n22588));
  nor_5  g20240(.A(new_n22588), .B(new_n4794), .Y(new_n22589));
  nand_5 g20241(.A(new_n13184), .B(new_n13174), .Y(new_n22590));
  nand_5 g20242(.A(new_n13192), .B(new_n13185), .Y(new_n22591));
  nand_5 g20243(.A(new_n22591), .B(new_n22590), .Y(new_n22592));
  xor_4  g20244(.A(new_n22588), .B(new_n4793), .Y(new_n22593));
  nor_5  g20245(.A(new_n22593), .B(new_n22592), .Y(new_n22594));
  nor_5  g20246(.A(new_n22594), .B(new_n22589), .Y(new_n22595));
  nor_5  g20247(.A(new_n22595), .B(new_n22587), .Y(new_n22596));
  nor_5  g20248(.A(new_n22596), .B(new_n22585), .Y(new_n22597));
  nor_5  g20249(.A(new_n22597), .B(new_n22583), .Y(new_n22598));
  nor_5  g20250(.A(new_n22598), .B(new_n22582), .Y(new_n22599));
  xor_4  g20251(.A(new_n22599), .B(new_n22580), .Y(new_n22600));
  not_8  g20252(.A(new_n22600), .Y(new_n22601));
  xor_4  g20253(.A(new_n22597), .B(new_n22583), .Y(new_n22602));
  not_8  g20254(.A(new_n13193), .Y(new_n22603));
  nor_5  g20255(.A(new_n13202), .B(new_n22603), .Y(new_n22604));
  nor_5  g20256(.A(new_n13203), .B(new_n3745), .Y(new_n22605));
  or_6   g20257(.A(new_n22605), .B(new_n22604), .Y(new_n22606));
  xnor_4 g20258(.A(new_n22593), .B(new_n22592), .Y(new_n22607));
  or_6   g20259(.A(new_n22607), .B(new_n22606), .Y(new_n22608));
  xor_4  g20260(.A(new_n22607), .B(new_n22606), .Y(new_n22609));
  nand_5 g20261(.A(new_n22609), .B(new_n3767), .Y(new_n22610));
  nand_5 g20262(.A(new_n22610), .B(new_n22608), .Y(new_n22611));
  xor_4  g20263(.A(new_n22595), .B(new_n22587), .Y(new_n22612));
  nor_5  g20264(.A(new_n22612), .B(new_n22611), .Y(new_n22613));
  nand_5 g20265(.A(new_n22612), .B(new_n22611), .Y(new_n22614));
  nand_5 g20266(.A(new_n22614), .B(new_n3743), .Y(new_n22615));
  not_8  g20267(.A(new_n22615), .Y(new_n22616));
  nor_5  g20268(.A(new_n22616), .B(new_n22613), .Y(new_n22617));
  nand_5 g20269(.A(new_n22617), .B(new_n22602), .Y(new_n22618));
  xor_4  g20270(.A(new_n22617), .B(new_n22602), .Y(new_n22619));
  nand_5 g20271(.A(new_n22619), .B(new_n17009), .Y(new_n22620));
  nand_5 g20272(.A(new_n22620), .B(new_n22618), .Y(new_n22621));
  nand_5 g20273(.A(new_n22621), .B(new_n22601), .Y(new_n22622));
  xor_4  g20274(.A(new_n22621), .B(new_n22600), .Y(new_n22623));
  or_6   g20275(.A(new_n22623), .B(new_n17007), .Y(new_n22624));
  nand_5 g20276(.A(new_n22624), .B(new_n22622), .Y(new_n22625));
  nand_5 g20277(.A(new_n11995), .B(new_n4930), .Y(new_n22626));
  nand_5 g20278(.A(new_n22578), .B(new_n22560), .Y(new_n22627));
  nand_5 g20279(.A(new_n22627), .B(new_n22626), .Y(new_n22628));
  xor_4  g20280(.A(new_n22628), .B(new_n21610), .Y(new_n22629));
  xor_4  g20281(.A(new_n22629), .B(new_n4863), .Y(new_n22630));
  nand_5 g20282(.A(new_n22579), .B(new_n4849), .Y(new_n22631));
  nand_5 g20283(.A(new_n22599), .B(new_n22580), .Y(new_n22632));
  nand_5 g20284(.A(new_n22632), .B(new_n22631), .Y(new_n22633));
  xor_4  g20285(.A(new_n22633), .B(new_n22630), .Y(new_n22634));
  not_8  g20286(.A(new_n22634), .Y(new_n22635));
  xor_4  g20287(.A(new_n22635), .B(new_n22625), .Y(new_n22636));
  xor_4  g20288(.A(new_n22636), .B(new_n17664), .Y(po0540));
  nand_5 g20289(.A(new_n20868), .B(new_n14199), .Y(new_n22638));
  nand_5 g20290(.A(new_n11447), .B(new_n11432), .Y(new_n22639));
  nand_5 g20291(.A(new_n11494), .B(new_n11448), .Y(new_n22640));
  nand_5 g20292(.A(new_n22640), .B(new_n22639), .Y(new_n22641));
  nand_5 g20293(.A(new_n22641), .B(new_n14200), .Y(new_n22642));
  xor_4  g20294(.A(new_n22641), .B(new_n14200), .Y(new_n22643));
  nand_5 g20295(.A(new_n22643), .B(new_n20872), .Y(new_n22644));
  nand_5 g20296(.A(new_n22644), .B(new_n22642), .Y(new_n22645));
  xor_4  g20297(.A(new_n20868), .B(new_n14199), .Y(new_n22646));
  nand_5 g20298(.A(new_n22646), .B(new_n22645), .Y(new_n22647));
  nand_5 g20299(.A(new_n22647), .B(new_n22638), .Y(po0541));
  xnor_4 g20300(.A(new_n21665), .B(new_n21664), .Y(po0542));
  nand_5 g20301(.A(new_n15102), .B(new_n11159), .Y(new_n22650));
  nand_5 g20302(.A(new_n15106), .B(new_n15103), .Y(new_n22651));
  nand_5 g20303(.A(new_n22651), .B(new_n22650), .Y(new_n22652));
  nand_5 g20304(.A(new_n22652), .B(new_n15097), .Y(new_n22653));
  nand_5 g20305(.A(new_n15098), .B(new_n15094), .Y(new_n22654));
  nand_5 g20306(.A(new_n15107), .B(new_n15099), .Y(new_n22655));
  nand_5 g20307(.A(new_n22655), .B(new_n22654), .Y(new_n22656));
  xor_4  g20308(.A(new_n22652), .B(new_n15097), .Y(new_n22657));
  nand_5 g20309(.A(new_n22657), .B(new_n22656), .Y(new_n22658));
  nand_5 g20310(.A(new_n22658), .B(new_n22653), .Y(po0543));
  nor_5  g20311(.A(new_n14927), .B(new_n14922), .Y(new_n22660));
  nor_5  g20312(.A(new_n22660), .B(new_n14926), .Y(new_n22661));
  xor_4  g20313(.A(new_n22661), .B(new_n15959), .Y(po0544));
  xor_4  g20314(.A(new_n9715), .B(new_n9714), .Y(po0545));
  xor_4  g20315(.A(new_n10821), .B(new_n22268), .Y(po0546));
  xor_4  g20316(.A(new_n4499), .B(new_n4446), .Y(po0547));
  nand_5 g20317(.A(new_n9169), .B(pi111), .Y(new_n22666));
  not_8  g20318(.A(new_n22666), .Y(new_n22667));
  xor_4  g20319(.A(pi512), .B(new_n16066), .Y(new_n22668));
  not_8  g20320(.A(new_n22668), .Y(new_n22669));
  nand_5 g20321(.A(pi537), .B(new_n9154), .Y(new_n22670));
  not_8  g20322(.A(new_n22670), .Y(new_n22671));
  xor_4  g20323(.A(pi537), .B(new_n9154), .Y(new_n22672));
  not_8  g20324(.A(new_n22672), .Y(new_n22673));
  nand_5 g20325(.A(pi671), .B(new_n2898), .Y(new_n22674));
  not_8  g20326(.A(new_n22674), .Y(new_n22675));
  xor_4  g20327(.A(pi671), .B(new_n2898), .Y(new_n22676));
  not_8  g20328(.A(new_n22676), .Y(new_n22677));
  nand_5 g20329(.A(new_n8641), .B(pi724), .Y(new_n22678));
  xor_4  g20330(.A(pi768), .B(new_n9143), .Y(new_n22679));
  nand_5 g20331(.A(pi756), .B(new_n13485), .Y(new_n22680));
  xor_4  g20332(.A(pi756), .B(new_n13485), .Y(new_n22681));
  nand_5 g20333(.A(new_n8591), .B(pi171), .Y(new_n22682));
  xor_4  g20334(.A(pi557), .B(new_n2908), .Y(new_n22683));
  nand_5 g20335(.A(pi414), .B(new_n8576), .Y(new_n22684));
  not_8  g20336(.A(new_n9616), .Y(new_n22685));
  nand_5 g20337(.A(new_n22685), .B(new_n9605), .Y(new_n22686));
  nand_5 g20338(.A(new_n22686), .B(new_n22684), .Y(new_n22687));
  nand_5 g20339(.A(new_n22687), .B(new_n22683), .Y(new_n22688));
  nand_5 g20340(.A(new_n22688), .B(new_n22682), .Y(new_n22689));
  nand_5 g20341(.A(new_n22689), .B(new_n22681), .Y(new_n22690));
  nand_5 g20342(.A(new_n22690), .B(new_n22680), .Y(new_n22691));
  nand_5 g20343(.A(new_n22691), .B(new_n22679), .Y(new_n22692));
  nand_5 g20344(.A(new_n22692), .B(new_n22678), .Y(new_n22693));
  nor_5  g20345(.A(new_n22693), .B(new_n22677), .Y(new_n22694));
  nor_5  g20346(.A(new_n22694), .B(new_n22675), .Y(new_n22695));
  nor_5  g20347(.A(new_n22695), .B(new_n22673), .Y(new_n22696));
  nor_5  g20348(.A(new_n22696), .B(new_n22671), .Y(new_n22697));
  nor_5  g20349(.A(new_n22697), .B(new_n22669), .Y(new_n22698));
  nor_5  g20350(.A(new_n22698), .B(new_n22667), .Y(new_n22699));
  or_6   g20351(.A(new_n22699), .B(new_n21837), .Y(new_n22700));
  xor_4  g20352(.A(new_n22695), .B(new_n22672), .Y(new_n22701));
  nand_5 g20353(.A(new_n22701), .B(new_n17562), .Y(new_n22702));
  xnor_4 g20354(.A(new_n22701), .B(new_n17562), .Y(new_n22703));
  xor_4  g20355(.A(new_n22693), .B(new_n22677), .Y(new_n22704));
  nand_5 g20356(.A(new_n22704), .B(new_n17565), .Y(new_n22705));
  xnor_4 g20357(.A(new_n22691), .B(new_n22679), .Y(new_n22706));
  nor_5  g20358(.A(new_n22706), .B(new_n17570), .Y(new_n22707));
  xor_4  g20359(.A(new_n22706), .B(new_n17571), .Y(new_n22708));
  not_8  g20360(.A(new_n17576), .Y(new_n22709));
  xor_4  g20361(.A(new_n22689), .B(new_n22681), .Y(new_n22710));
  nor_5  g20362(.A(new_n22710), .B(new_n22709), .Y(new_n22711));
  xor_4  g20363(.A(new_n22687), .B(new_n22683), .Y(new_n22712));
  not_8  g20364(.A(new_n22712), .Y(new_n22713));
  nor_5  g20365(.A(new_n22713), .B(new_n17581), .Y(new_n22714));
  xor_4  g20366(.A(new_n22712), .B(new_n17581), .Y(new_n22715));
  nor_5  g20367(.A(new_n9617), .B(new_n9604), .Y(new_n22716));
  nor_5  g20368(.A(new_n9640), .B(new_n9618), .Y(new_n22717));
  nor_5  g20369(.A(new_n22717), .B(new_n22716), .Y(new_n22718));
  nor_5  g20370(.A(new_n22718), .B(new_n22715), .Y(new_n22719));
  or_6   g20371(.A(new_n22719), .B(new_n22714), .Y(new_n22720));
  xor_4  g20372(.A(new_n22710), .B(new_n17576), .Y(new_n22721));
  nor_5  g20373(.A(new_n22721), .B(new_n22720), .Y(new_n22722));
  or_6   g20374(.A(new_n22722), .B(new_n22711), .Y(new_n22723));
  nor_5  g20375(.A(new_n22723), .B(new_n22708), .Y(new_n22724));
  or_6   g20376(.A(new_n22724), .B(new_n22707), .Y(new_n22725));
  xnor_4 g20377(.A(new_n22704), .B(new_n17565), .Y(new_n22726));
  or_6   g20378(.A(new_n22726), .B(new_n22725), .Y(new_n22727));
  nand_5 g20379(.A(new_n22727), .B(new_n22705), .Y(new_n22728));
  or_6   g20380(.A(new_n22728), .B(new_n22703), .Y(new_n22729));
  nand_5 g20381(.A(new_n22729), .B(new_n22702), .Y(new_n22730));
  xor_4  g20382(.A(new_n22697), .B(new_n22668), .Y(new_n22731));
  or_6   g20383(.A(new_n22731), .B(new_n17532), .Y(new_n22732));
  nand_5 g20384(.A(new_n22732), .B(new_n22730), .Y(new_n22733));
  nand_5 g20385(.A(new_n22731), .B(new_n17532), .Y(new_n22734));
  nand_5 g20386(.A(new_n22734), .B(new_n22733), .Y(new_n22735));
  nor_5  g20387(.A(new_n22735), .B(new_n22700), .Y(new_n22736));
  not_8  g20388(.A(new_n22735), .Y(new_n22737));
  nand_5 g20389(.A(new_n22699), .B(new_n21837), .Y(new_n22738));
  nor_5  g20390(.A(new_n22738), .B(new_n22737), .Y(new_n22739));
  nor_5  g20391(.A(new_n22739), .B(new_n22736), .Y(new_n22740));
  xor_4  g20392(.A(new_n22740), .B(new_n21831), .Y(po0548));
  xnor_4 g20393(.A(new_n13254), .B(new_n13249), .Y(po0549));
  xnor_4 g20394(.A(new_n14776), .B(new_n14737), .Y(po0550));
  xnor_4 g20395(.A(new_n6291), .B(new_n6272), .Y(po0551));
  xnor_4 g20396(.A(new_n18466), .B(new_n18451), .Y(po0552));
  xnor_4 g20397(.A(new_n16038), .B(new_n16037), .Y(po0553));
  xor_4  g20398(.A(new_n17249), .B(new_n17251), .Y(po0554));
  not_8  g20399(.A(new_n22094), .Y(new_n22748));
  nand_5 g20400(.A(new_n22106), .B(new_n22748), .Y(new_n22749));
  not_8  g20401(.A(new_n22749), .Y(new_n22750));
  nor_5  g20402(.A(new_n22107), .B(new_n22084), .Y(new_n22751));
  nor_5  g20403(.A(new_n22751), .B(new_n22750), .Y(new_n22752));
  not_8  g20404(.A(new_n22752), .Y(new_n22753));
  xor_4  g20405(.A(new_n22100), .B(new_n22088), .Y(new_n22754));
  xor_4  g20406(.A(new_n22754), .B(new_n22753), .Y(po0555));
  xor_4  g20407(.A(new_n15209), .B(new_n15206), .Y(po0556));
  xor_4  g20408(.A(new_n14778), .B(new_n14733), .Y(po0557));
  xnor_4 g20409(.A(new_n2767), .B(new_n2766), .Y(po0558));
  xor_4  g20410(.A(new_n20875), .B(new_n20872), .Y(new_n22759));
  xnor_4 g20411(.A(new_n22759), .B(new_n20871), .Y(po0559));
  xor_4  g20412(.A(new_n21584), .B(new_n21580), .Y(po0560));
  xor_4  g20413(.A(new_n17254), .B(new_n17128), .Y(po0561));
  nand_5 g20414(.A(new_n19538), .B(new_n4871), .Y(new_n22763));
  nand_5 g20415(.A(new_n20380), .B(new_n4872), .Y(new_n22764));
  not_8  g20416(.A(new_n22764), .Y(new_n22765));
  nor_5  g20417(.A(new_n9521), .B(new_n4916), .Y(new_n22766));
  xor_4  g20418(.A(new_n9520), .B(new_n4916), .Y(new_n22767));
  or_6   g20419(.A(new_n9481), .B(new_n4906), .Y(new_n22768));
  xor_4  g20420(.A(new_n9481), .B(new_n4906), .Y(new_n22769));
  nand_5 g20421(.A(new_n9409), .B(new_n4899), .Y(new_n22770));
  xor_4  g20422(.A(new_n9409), .B(new_n4899), .Y(new_n22771));
  nand_5 g20423(.A(new_n9446), .B(new_n4887), .Y(new_n22772));
  nor_5  g20424(.A(new_n22772), .B(new_n9445), .Y(new_n22773));
  xor_4  g20425(.A(new_n22772), .B(new_n9444), .Y(new_n22774));
  nor_5  g20426(.A(new_n22774), .B(new_n4882), .Y(new_n22775));
  nor_5  g20427(.A(new_n22775), .B(new_n22773), .Y(new_n22776));
  nand_5 g20428(.A(new_n22776), .B(new_n4893), .Y(new_n22777));
  not_8  g20429(.A(new_n9443), .Y(new_n22778));
  xnor_4 g20430(.A(new_n22776), .B(new_n4893), .Y(new_n22779));
  or_6   g20431(.A(new_n22779), .B(new_n22778), .Y(new_n22780));
  nand_5 g20432(.A(new_n22780), .B(new_n22777), .Y(new_n22781));
  nand_5 g20433(.A(new_n22781), .B(new_n22771), .Y(new_n22782));
  nand_5 g20434(.A(new_n22782), .B(new_n22770), .Y(new_n22783));
  nand_5 g20435(.A(new_n22783), .B(new_n22769), .Y(new_n22784));
  nand_5 g20436(.A(new_n22784), .B(new_n22768), .Y(new_n22785));
  nor_5  g20437(.A(new_n22785), .B(new_n22767), .Y(new_n22786));
  or_6   g20438(.A(new_n22786), .B(new_n22766), .Y(new_n22787));
  or_6   g20439(.A(new_n22787), .B(new_n9564), .Y(new_n22788));
  xor_4  g20440(.A(new_n22787), .B(new_n9564), .Y(new_n22789));
  nand_5 g20441(.A(new_n22789), .B(new_n4877), .Y(new_n22790));
  nand_5 g20442(.A(new_n22790), .B(new_n22788), .Y(new_n22791));
  nor_5  g20443(.A(new_n22791), .B(new_n19567), .Y(new_n22792));
  xor_4  g20444(.A(new_n22791), .B(new_n20361), .Y(new_n22793));
  nor_5  g20445(.A(new_n22793), .B(new_n4875), .Y(new_n22794));
  or_6   g20446(.A(new_n22794), .B(new_n22792), .Y(new_n22795));
  nand_5 g20447(.A(new_n22795), .B(new_n19562), .Y(new_n22796));
  xor_4  g20448(.A(new_n22795), .B(new_n19561), .Y(new_n22797));
  or_6   g20449(.A(new_n22797), .B(new_n4927), .Y(new_n22798));
  nand_5 g20450(.A(new_n22798), .B(new_n22796), .Y(new_n22799));
  or_6   g20451(.A(new_n22799), .B(new_n20323), .Y(new_n22800));
  xor_4  g20452(.A(new_n22799), .B(new_n20323), .Y(new_n22801));
  nand_5 g20453(.A(new_n22801), .B(new_n4935), .Y(new_n22802));
  nand_5 g20454(.A(new_n22802), .B(new_n22800), .Y(new_n22803));
  xor_4  g20455(.A(new_n19558), .B(new_n4872), .Y(new_n22804));
  nor_5  g20456(.A(new_n22804), .B(new_n22803), .Y(new_n22805));
  nor_5  g20457(.A(new_n22805), .B(new_n22765), .Y(new_n22806));
  xor_4  g20458(.A(new_n19539), .B(new_n4871), .Y(new_n22807));
  or_6   g20459(.A(new_n22807), .B(new_n22806), .Y(new_n22808));
  nand_5 g20460(.A(new_n22808), .B(new_n22763), .Y(po0562));
  xor_4  g20461(.A(new_n20106), .B(new_n16795), .Y(po0563));
  not_8  g20462(.A(new_n20391), .Y(new_n22811));
  nor_5  g20463(.A(new_n22811), .B(new_n20385), .Y(new_n22812));
  nor_5  g20464(.A(new_n22812), .B(new_n20387), .Y(new_n22813));
  nor_5  g20465(.A(new_n22813), .B(new_n20379), .Y(po0564));
  xnor_4 g20466(.A(new_n20614), .B(new_n20613), .Y(po0565));
  xor_4  g20467(.A(new_n15805), .B(new_n15755), .Y(po0566));
  xor_4  g20468(.A(new_n9635), .B(new_n9626), .Y(po0567));
  xnor_4 g20469(.A(new_n16132), .B(new_n15468), .Y(po0568));
  nand_5 g20470(.A(new_n16398), .B(new_n16397), .Y(new_n22819));
  xor_4  g20471(.A(new_n22819), .B(new_n8610), .Y(po0569));
  nand_5 g20472(.A(new_n18454), .B(new_n18455), .Y(new_n22821));
  xor_4  g20473(.A(new_n22821), .B(new_n6902), .Y(po0570));
  not_8  g20474(.A(new_n11631), .Y(new_n22823));
  and_6  g20475(.A(new_n21065), .B(new_n9763), .Y(new_n22824));
  nor_5  g20476(.A(new_n21329), .B(new_n21322), .Y(new_n22825));
  nor_5  g20477(.A(new_n22825), .B(new_n22824), .Y(new_n22826));
  xor_4  g20478(.A(new_n21655), .B(new_n21071), .Y(new_n22827));
  xnor_4 g20479(.A(new_n22827), .B(new_n22826), .Y(new_n22828));
  xor_4  g20480(.A(new_n22828), .B(new_n22823), .Y(new_n22829));
  nor_5  g20481(.A(new_n21331), .B(new_n11623), .Y(new_n22830));
  nor_5  g20482(.A(new_n21342), .B(new_n21333), .Y(new_n22831));
  nor_5  g20483(.A(new_n22831), .B(new_n22830), .Y(new_n22832));
  xnor_4 g20484(.A(new_n22832), .B(new_n22829), .Y(po0571));
  xor_4  g20485(.A(new_n11480), .B(new_n4620), .Y(po0572));
  xnor_4 g20486(.A(new_n13598), .B(new_n13596), .Y(po0573));
  nand_5 g20487(.A(new_n17781), .B(new_n17780), .Y(new_n22836));
  xor_4  g20488(.A(new_n22836), .B(new_n12273), .Y(po0574));
  xnor_4 g20489(.A(new_n16336), .B(new_n16317), .Y(po0575));
  xor_4  g20490(.A(new_n15815), .B(new_n15814), .Y(po0576));
  xor_4  g20491(.A(new_n10009), .B(new_n10007), .Y(po0577));
  xor_4  g20492(.A(new_n10011), .B(new_n10010), .Y(po0578));
  xnor_4 g20493(.A(new_n21451), .B(new_n21450), .Y(po0579));
  xor_4  g20494(.A(new_n12668), .B(new_n12667), .Y(po0580));
  nand_5 g20495(.A(new_n16892), .B(new_n5692), .Y(new_n22844));
  nand_5 g20496(.A(new_n22844), .B(new_n5770), .Y(new_n22845));
  xor_4  g20497(.A(new_n22844), .B(new_n10769), .Y(new_n22846));
  not_8  g20498(.A(new_n22846), .Y(new_n22847));
  nand_5 g20499(.A(new_n22847), .B(new_n5698), .Y(new_n22848));
  nand_5 g20500(.A(new_n22848), .B(new_n22845), .Y(new_n22849));
  nand_5 g20501(.A(new_n22849), .B(new_n10768), .Y(new_n22850));
  xor_4  g20502(.A(new_n22849), .B(new_n10774), .Y(new_n22851));
  or_6   g20503(.A(new_n22851), .B(new_n5707), .Y(new_n22852));
  nand_5 g20504(.A(new_n22852), .B(new_n22850), .Y(new_n22853));
  nor_5  g20505(.A(new_n22853), .B(new_n5712), .Y(new_n22854));
  nand_5 g20506(.A(new_n22854), .B(new_n13150), .Y(new_n22855));
  nand_5 g20507(.A(new_n22853), .B(new_n5712), .Y(new_n22856));
  nand_5 g20508(.A(new_n22856), .B(new_n10778), .Y(new_n22857));
  nand_5 g20509(.A(new_n22857), .B(new_n22855), .Y(new_n22858));
  nand_5 g20510(.A(new_n22858), .B(new_n10791), .Y(new_n22859));
  not_8  g20511(.A(new_n22859), .Y(new_n22860));
  nand_5 g20512(.A(new_n22856), .B(new_n10747), .Y(new_n22861));
  nand_5 g20513(.A(new_n22854), .B(pi618), .Y(new_n22862));
  and_6  g20514(.A(new_n22862), .B(new_n22861), .Y(new_n22863));
  nand_5 g20515(.A(new_n10754), .B(new_n10745), .Y(new_n22864));
  nor_5  g20516(.A(new_n22864), .B(new_n22863), .Y(new_n22865));
  nor_5  g20517(.A(new_n22865), .B(new_n22860), .Y(new_n22866));
  xor_4  g20518(.A(new_n22853), .B(new_n5713), .Y(new_n22867));
  or_6   g20519(.A(new_n22867), .B(new_n10780), .Y(new_n22868));
  nand_5 g20520(.A(new_n22868), .B(new_n22856), .Y(new_n22869));
  nand_5 g20521(.A(new_n22869), .B(new_n10767), .Y(new_n22870));
  and_6  g20522(.A(new_n22870), .B(new_n22866), .Y(new_n22871));
  xor_4  g20523(.A(new_n22871), .B(new_n5718), .Y(po0581));
  nor_5  g20524(.A(new_n8445), .B(new_n8443), .Y(new_n22873));
  not_8  g20525(.A(new_n22873), .Y(new_n22874));
  nor_5  g20526(.A(new_n3470), .B(new_n3423), .Y(new_n22875));
  nor_5  g20527(.A(new_n3522), .B(new_n3472), .Y(new_n22876));
  nor_5  g20528(.A(new_n22876), .B(new_n22875), .Y(new_n22877));
  nor_5  g20529(.A(new_n22877), .B(new_n13551), .Y(new_n22878));
  and_6  g20530(.A(new_n22878), .B(new_n22874), .Y(new_n22879));
  nor_5  g20531(.A(new_n22878), .B(new_n22874), .Y(new_n22880));
  nor_5  g20532(.A(new_n22880), .B(new_n22879), .Y(new_n22881));
  xor_4  g20533(.A(new_n22877), .B(new_n13551), .Y(new_n22882));
  or_6   g20534(.A(new_n22882), .B(new_n8447), .Y(new_n22883));
  nor_5  g20535(.A(new_n3706), .B(new_n3691), .Y(new_n22884));
  nor_5  g20536(.A(new_n3707), .B(new_n3523), .Y(new_n22885));
  nor_5  g20537(.A(new_n22885), .B(new_n22884), .Y(new_n22886));
  xor_4  g20538(.A(new_n22882), .B(new_n8446), .Y(new_n22887));
  or_6   g20539(.A(new_n22887), .B(new_n22886), .Y(new_n22888));
  nand_5 g20540(.A(new_n22888), .B(new_n22883), .Y(new_n22889));
  not_8  g20541(.A(new_n22889), .Y(new_n22890));
  xor_4  g20542(.A(new_n22890), .B(new_n22881), .Y(po0582));
  xor_4  g20543(.A(new_n18068), .B(new_n9022), .Y(po0583));
  xor_4  g20544(.A(new_n5342), .B(new_n14954), .Y(po0584));
  xnor_4 g20545(.A(new_n20444), .B(new_n20417), .Y(po0585));
  xnor_4 g20546(.A(new_n6040), .B(new_n6039), .Y(po0586));
  not_8  g20547(.A(pi425), .Y(new_n22896));
  not_8  g20548(.A(new_n16224), .Y(new_n22897));
  nand_5 g20549(.A(new_n22897), .B(new_n22896), .Y(new_n22898));
  nand_5 g20550(.A(new_n16203), .B(pi159), .Y(new_n22899));
  not_8  g20551(.A(new_n22899), .Y(new_n22900));
  nor_5  g20552(.A(new_n19518), .B(new_n16205), .Y(new_n22901));
  nor_5  g20553(.A(new_n22901), .B(new_n22900), .Y(new_n22902));
  nand_5 g20554(.A(new_n22902), .B(new_n16225), .Y(new_n22903));
  nand_5 g20555(.A(new_n22903), .B(new_n22898), .Y(new_n22904));
  nand_5 g20556(.A(new_n16223), .B(new_n16218), .Y(new_n22905));
  nand_5 g20557(.A(new_n22905), .B(new_n16217), .Y(new_n22906));
  nor_5  g20558(.A(new_n22906), .B(new_n22904), .Y(new_n22907));
  and_6  g20559(.A(new_n22906), .B(new_n22904), .Y(new_n22908));
  nor_5  g20560(.A(new_n22908), .B(new_n22907), .Y(new_n22909));
  xor_4  g20561(.A(new_n22909), .B(new_n3324), .Y(new_n22910));
  xor_4  g20562(.A(new_n22902), .B(new_n16225), .Y(new_n22911));
  or_6   g20563(.A(new_n22911), .B(new_n3315), .Y(new_n22912));
  xor_4  g20564(.A(new_n22911), .B(new_n3315), .Y(new_n22913));
  nor_5  g20565(.A(new_n19519), .B(new_n3309), .Y(new_n22914));
  and_6  g20566(.A(new_n19520), .B(new_n19513), .Y(new_n22915));
  nor_5  g20567(.A(new_n22915), .B(new_n22914), .Y(new_n22916));
  nand_5 g20568(.A(new_n22916), .B(new_n22913), .Y(new_n22917));
  nand_5 g20569(.A(new_n22917), .B(new_n22912), .Y(new_n22918));
  not_8  g20570(.A(new_n22918), .Y(new_n22919));
  nor_5  g20571(.A(new_n22919), .B(new_n22910), .Y(new_n22920));
  nor_5  g20572(.A(new_n22907), .B(new_n3323), .Y(new_n22921));
  nor_5  g20573(.A(new_n22907), .B(new_n3207), .Y(new_n22922));
  nor_5  g20574(.A(new_n22908), .B(new_n3416), .Y(new_n22923));
  nor_5  g20575(.A(new_n22923), .B(new_n22922), .Y(new_n22924));
  nor_5  g20576(.A(new_n22924), .B(new_n22921), .Y(new_n22925));
  xor_4  g20577(.A(new_n22925), .B(new_n22920), .Y(po0587));
  xnor_4 g20578(.A(new_n21356), .B(new_n18100), .Y(po0588));
  nand_5 g20579(.A(new_n8997), .B(pi642), .Y(new_n22928));
  nand_5 g20580(.A(new_n8998), .B(new_n7245), .Y(new_n22929));
  nand_5 g20581(.A(new_n22929), .B(new_n22928), .Y(new_n22930));
  nand_5 g20582(.A(pi694), .B(pi680), .Y(new_n22931));
  or_6   g20583(.A(pi694), .B(pi680), .Y(new_n22932));
  nand_5 g20584(.A(new_n22932), .B(new_n22931), .Y(new_n22933));
  xor_4  g20585(.A(new_n22933), .B(new_n9650), .Y(new_n22934));
  xor_4  g20586(.A(new_n22934), .B(new_n22930), .Y(new_n22935));
  nand_5 g20587(.A(new_n8999), .B(pi642), .Y(new_n22936));
  or_6   g20588(.A(new_n22936), .B(new_n9650), .Y(new_n22937));
  nand_5 g20589(.A(new_n22937), .B(new_n22935), .Y(new_n22938));
  nand_5 g20590(.A(new_n22936), .B(new_n9650), .Y(new_n22939));
  nand_5 g20591(.A(new_n22939), .B(new_n22938), .Y(new_n22940));
  xor_4  g20592(.A(new_n22940), .B(pi658), .Y(new_n22941));
  nand_5 g20593(.A(pi529), .B(pi051), .Y(new_n22942));
  nand_5 g20594(.A(new_n9690), .B(new_n4084), .Y(new_n22943));
  nand_5 g20595(.A(new_n22943), .B(new_n22942), .Y(new_n22944));
  nand_5 g20596(.A(new_n22931), .B(new_n8998), .Y(new_n22945));
  nand_5 g20597(.A(new_n22945), .B(new_n22932), .Y(new_n22946));
  xor_4  g20598(.A(new_n22946), .B(new_n22944), .Y(new_n22947));
  xnor_4 g20599(.A(new_n22947), .B(new_n22941), .Y(new_n22948));
  nor_5  g20600(.A(new_n9000), .B(new_n8996), .Y(new_n22949));
  not_8  g20601(.A(new_n22949), .Y(new_n22950));
  nor_5  g20602(.A(new_n22935), .B(new_n22950), .Y(new_n22951));
  xor_4  g20603(.A(new_n22935), .B(new_n22949), .Y(new_n22952));
  nor_5  g20604(.A(new_n22952), .B(new_n18633), .Y(new_n22953));
  nor_5  g20605(.A(new_n22953), .B(new_n22951), .Y(new_n22954));
  xor_4  g20606(.A(new_n22954), .B(new_n22948), .Y(new_n22955));
  xnor_4 g20607(.A(new_n22955), .B(new_n18628), .Y(po0589));
  nand_5 g20608(.A(new_n22115), .B(new_n22112), .Y(new_n22957));
  not_8  g20609(.A(new_n22957), .Y(new_n22958));
  nor_5  g20610(.A(new_n22120), .B(new_n22117), .Y(new_n22959));
  nor_5  g20611(.A(new_n22959), .B(new_n22958), .Y(new_n22960));
  nand_5 g20612(.A(new_n22960), .B(new_n7745), .Y(new_n22961));
  nand_5 g20613(.A(new_n22124), .B(new_n22121), .Y(new_n22962));
  nand_5 g20614(.A(new_n22125), .B(new_n7745), .Y(new_n22963));
  and_6  g20615(.A(new_n22963), .B(new_n22962), .Y(new_n22964));
  xor_4  g20616(.A(new_n22960), .B(new_n9002), .Y(new_n22965));
  not_8  g20617(.A(new_n22965), .Y(new_n22966));
  nand_5 g20618(.A(new_n22966), .B(new_n22964), .Y(new_n22967));
  nand_5 g20619(.A(new_n22967), .B(new_n22961), .Y(po0590));
  xor_4  g20620(.A(new_n22368), .B(new_n22348), .Y(po0591));
  xnor_4 g20621(.A(new_n21876), .B(new_n21867), .Y(po0592));
  or_6   g20622(.A(new_n22546), .B(new_n22542), .Y(new_n22971));
  nor_5  g20623(.A(new_n22551), .B(new_n22971), .Y(new_n22972));
  or_6   g20624(.A(new_n22972), .B(new_n22553), .Y(po0593));
  not_8  g20625(.A(new_n11290), .Y(new_n22974));
  nand_5 g20626(.A(new_n22974), .B(new_n11089), .Y(new_n22975));
  nand_5 g20627(.A(new_n11291), .B(new_n11287), .Y(new_n22976));
  nand_5 g20628(.A(new_n22976), .B(new_n22975), .Y(po0594));
  xnor_4 g20629(.A(new_n12063), .B(new_n12021), .Y(po0595));
  xor_4  g20630(.A(new_n13103), .B(new_n10679), .Y(po0596));
  xor_4  g20631(.A(new_n21640), .B(new_n16441), .Y(po0597));
  nand_5 g20632(.A(new_n12300), .B(new_n6714), .Y(new_n22981));
  nand_5 g20633(.A(new_n22981), .B(new_n12299), .Y(new_n22982));
  nor_5  g20634(.A(new_n22982), .B(new_n7319), .Y(new_n22983));
  xor_4  g20635(.A(new_n22982), .B(new_n7318), .Y(new_n22984));
  nor_5  g20636(.A(new_n22984), .B(new_n6787), .Y(new_n22985));
  or_6   g20637(.A(new_n22985), .B(new_n22983), .Y(new_n22986));
  nand_5 g20638(.A(new_n22986), .B(new_n7312), .Y(new_n22987));
  not_8  g20639(.A(new_n22987), .Y(new_n22988));
  nor_5  g20640(.A(new_n22986), .B(new_n7312), .Y(new_n22989));
  nor_5  g20641(.A(new_n22989), .B(new_n7592), .Y(new_n22990));
  nor_5  g20642(.A(new_n22990), .B(new_n22988), .Y(new_n22991));
  xor_4  g20643(.A(new_n22991), .B(new_n7293), .Y(new_n22992));
  xor_4  g20644(.A(new_n22992), .B(new_n7590), .Y(new_n22993));
  nor_5  g20645(.A(new_n22993), .B(new_n22481), .Y(new_n22994));
  xor_4  g20646(.A(new_n22993), .B(new_n22482), .Y(new_n22995));
  xor_4  g20647(.A(new_n22984), .B(new_n6787), .Y(new_n22996));
  not_8  g20648(.A(new_n22996), .Y(new_n22997));
  or_6   g20649(.A(new_n12302), .B(new_n12296), .Y(new_n22998));
  nand_5 g20650(.A(new_n12303), .B(new_n12232), .Y(new_n22999));
  nand_5 g20651(.A(new_n22999), .B(new_n22998), .Y(new_n23000));
  nor_5  g20652(.A(new_n23000), .B(new_n22997), .Y(new_n23001));
  xor_4  g20653(.A(new_n23000), .B(new_n22996), .Y(new_n23002));
  nor_5  g20654(.A(new_n23002), .B(new_n22485), .Y(new_n23003));
  or_6   g20655(.A(new_n23003), .B(new_n23001), .Y(new_n23004));
  nand_5 g20656(.A(new_n23004), .B(new_n22491), .Y(new_n23005));
  nor_5  g20657(.A(new_n22989), .B(new_n22988), .Y(new_n23006));
  xor_4  g20658(.A(new_n23006), .B(new_n7592), .Y(new_n23007));
  xor_4  g20659(.A(new_n23004), .B(new_n22489), .Y(new_n23008));
  or_6   g20660(.A(new_n23008), .B(new_n23007), .Y(new_n23009));
  nand_5 g20661(.A(new_n23009), .B(new_n23005), .Y(new_n23010));
  nor_5  g20662(.A(new_n23010), .B(new_n22995), .Y(new_n23011));
  or_6   g20663(.A(new_n23011), .B(new_n22994), .Y(new_n23012));
  nor_5  g20664(.A(new_n23012), .B(new_n22532), .Y(new_n23013));
  xor_4  g20665(.A(new_n23012), .B(new_n22532), .Y(new_n23014));
  or_6   g20666(.A(new_n23014), .B(new_n7378), .Y(new_n23015));
  not_8  g20667(.A(new_n7293), .Y(new_n23016));
  nand_5 g20668(.A(new_n22991), .B(new_n23016), .Y(new_n23017));
  or_6   g20669(.A(new_n22992), .B(pi096), .Y(new_n23018));
  nand_5 g20670(.A(new_n23018), .B(new_n23017), .Y(new_n23019));
  xor_4  g20671(.A(new_n23014), .B(new_n7378), .Y(new_n23020));
  nand_5 g20672(.A(new_n23020), .B(new_n23019), .Y(new_n23021));
  nand_5 g20673(.A(new_n23021), .B(new_n23015), .Y(new_n23022));
  nor_5  g20674(.A(new_n23022), .B(new_n23013), .Y(new_n23023));
  and_6  g20675(.A(new_n23022), .B(new_n22522), .Y(new_n23024));
  nor_5  g20676(.A(new_n23024), .B(new_n23023), .Y(po0598));
  nand_5 g20677(.A(new_n19355), .B(pi826), .Y(new_n23026));
  nand_5 g20678(.A(new_n23026), .B(new_n19354), .Y(new_n23027));
  nand_5 g20679(.A(new_n23027), .B(new_n8808), .Y(new_n23028));
  or_6   g20680(.A(new_n23027), .B(new_n8808), .Y(new_n23029));
  nand_5 g20681(.A(new_n23029), .B(pi150), .Y(new_n23030));
  nand_5 g20682(.A(new_n23030), .B(new_n23028), .Y(new_n23031));
  nand_5 g20683(.A(new_n23031), .B(new_n8804), .Y(new_n23032));
  or_6   g20684(.A(new_n23031), .B(new_n8804), .Y(new_n23033));
  nand_5 g20685(.A(new_n23033), .B(new_n23032), .Y(new_n23034));
  xor_4  g20686(.A(new_n23034), .B(pi782), .Y(new_n23035));
  nand_5 g20687(.A(new_n19362), .B(pi572), .Y(new_n23036));
  nand_5 g20688(.A(new_n23036), .B(new_n19361), .Y(new_n23037));
  nor_5  g20689(.A(new_n23037), .B(pi033), .Y(new_n23038));
  xor_4  g20690(.A(new_n23037), .B(new_n6799), .Y(new_n23039));
  nor_5  g20691(.A(new_n23039), .B(new_n16697), .Y(new_n23040));
  or_6   g20692(.A(new_n23040), .B(new_n23038), .Y(new_n23041));
  xor_4  g20693(.A(new_n23041), .B(new_n16702), .Y(new_n23042));
  xor_4  g20694(.A(new_n23042), .B(new_n6824), .Y(new_n23043));
  nor_5  g20695(.A(new_n23043), .B(new_n23035), .Y(new_n23044));
  not_8  g20696(.A(new_n23035), .Y(new_n23045));
  xor_4  g20697(.A(new_n23043), .B(new_n23045), .Y(new_n23046));
  and_6  g20698(.A(new_n23029), .B(new_n23028), .Y(new_n23047));
  xor_4  g20699(.A(new_n23047), .B(new_n6220), .Y(new_n23048));
  xnor_4 g20700(.A(new_n23039), .B(new_n16697), .Y(new_n23049));
  nor_5  g20701(.A(new_n23049), .B(new_n23048), .Y(new_n23050));
  nor_5  g20702(.A(new_n19364), .B(new_n19357), .Y(new_n23051));
  nor_5  g20703(.A(new_n19368), .B(new_n19365), .Y(new_n23052));
  or_6   g20704(.A(new_n23052), .B(new_n23051), .Y(new_n23053));
  not_8  g20705(.A(new_n23048), .Y(new_n23054));
  xor_4  g20706(.A(new_n23049), .B(new_n23054), .Y(new_n23055));
  nor_5  g20707(.A(new_n23055), .B(new_n23053), .Y(new_n23056));
  nor_5  g20708(.A(new_n23056), .B(new_n23050), .Y(new_n23057));
  nor_5  g20709(.A(new_n23057), .B(new_n23046), .Y(new_n23058));
  or_6   g20710(.A(new_n23058), .B(new_n23044), .Y(new_n23059));
  nand_5 g20711(.A(new_n23032), .B(new_n6260), .Y(new_n23060));
  nand_5 g20712(.A(new_n23060), .B(new_n23033), .Y(new_n23061));
  or_6   g20713(.A(new_n23061), .B(new_n8756), .Y(new_n23062));
  nand_5 g20714(.A(new_n23061), .B(new_n8756), .Y(new_n23063));
  and_6  g20715(.A(new_n23063), .B(new_n23062), .Y(new_n23064));
  xor_4  g20716(.A(new_n23064), .B(new_n6294), .Y(new_n23065));
  xor_4  g20717(.A(new_n16675), .B(pi666), .Y(new_n23066));
  nand_5 g20718(.A(new_n23041), .B(new_n16739), .Y(new_n23067));
  or_6   g20719(.A(new_n23042), .B(pi437), .Y(new_n23068));
  nand_5 g20720(.A(new_n23068), .B(new_n23067), .Y(new_n23069));
  xor_4  g20721(.A(new_n23069), .B(new_n23066), .Y(new_n23070));
  xor_4  g20722(.A(new_n23070), .B(new_n23065), .Y(new_n23071));
  xor_4  g20723(.A(new_n23071), .B(new_n23059), .Y(po0599));
  xor_4  g20724(.A(new_n20611), .B(new_n20609), .Y(po0600));
  xor_4  g20725(.A(new_n21361), .B(new_n18123), .Y(po0601));
  xor_4  g20726(.A(new_n14002), .B(new_n13988), .Y(new_n23075));
  xor_4  g20727(.A(new_n23075), .B(new_n14006), .Y(po0602));
  xor_4  g20728(.A(new_n22721), .B(new_n22720), .Y(po0603));
  xor_4  g20729(.A(new_n21444), .B(new_n21442), .Y(po0604));
  xor_4  g20730(.A(new_n6537), .B(new_n4695), .Y(po0605));
  nand_5 g20731(.A(new_n4999), .B(new_n4993), .Y(new_n23080));
  xor_4  g20732(.A(new_n23080), .B(new_n16598), .Y(po0606));
  xnor_4 g20733(.A(new_n15211), .B(new_n15200), .Y(po0607));
  xor_4  g20734(.A(new_n11278), .B(new_n8755), .Y(po0608));
  xor_4  g20735(.A(new_n3644), .B(new_n3633), .Y(po0609));
  xnor_4 g20736(.A(new_n10613), .B(new_n10612), .Y(po0610));
  xnor_4 g20737(.A(new_n14026), .B(new_n14025), .Y(po0611));
  xor_4  g20738(.A(new_n22106), .B(new_n18836), .Y(new_n23087));
  nor_5  g20739(.A(new_n21745), .B(new_n21740), .Y(new_n23088));
  nor_5  g20740(.A(new_n21747), .B(new_n20239), .Y(new_n23089));
  nor_5  g20741(.A(new_n23089), .B(new_n23088), .Y(new_n23090));
  xor_4  g20742(.A(new_n23090), .B(new_n23087), .Y(po0612));
  xnor_4 g20743(.A(new_n8714), .B(new_n8702), .Y(po0613));
  xnor_4 g20744(.A(new_n23057), .B(new_n23046), .Y(po0614));
  nand_5 g20745(.A(new_n13726), .B(new_n13723), .Y(po0615));
  xor_4  g20746(.A(new_n9458), .B(new_n9444), .Y(new_n23095));
  xor_4  g20747(.A(new_n23095), .B(new_n9419), .Y(po0616));
  xor_4  g20748(.A(new_n17028), .B(new_n16456), .Y(new_n23097));
  xor_4  g20749(.A(new_n23097), .B(new_n17025), .Y(po0617));
  xor_4  g20750(.A(new_n14069), .B(new_n14062), .Y(po0618));
  xnor_4 g20751(.A(new_n17267), .B(new_n17230), .Y(po0619));
  xor_4  g20752(.A(new_n11262), .B(new_n8812), .Y(po0620));
  xor_4  g20753(.A(new_n22779), .B(new_n22778), .Y(po0621));
  xor_4  g20754(.A(new_n15299), .B(new_n15298), .Y(po0622));
  nand_5 g20755(.A(pi689), .B(new_n16066), .Y(new_n23104));
  not_8  g20756(.A(new_n23104), .Y(new_n23105));
  nand_5 g20757(.A(new_n8383), .B(pi111), .Y(new_n23106));
  not_8  g20758(.A(new_n23106), .Y(new_n23107));
  nand_5 g20759(.A(new_n16070), .B(pi009), .Y(new_n23108));
  not_8  g20760(.A(new_n23108), .Y(new_n23109));
  nand_5 g20761(.A(pi537), .B(new_n20462), .Y(new_n23110));
  not_8  g20762(.A(new_n23110), .Y(new_n23111));
  nand_5 g20763(.A(new_n16177), .B(pi180), .Y(new_n23112));
  not_8  g20764(.A(new_n23112), .Y(new_n23113));
  nor_5  g20765(.A(new_n17480), .B(new_n17479), .Y(new_n23114));
  nor_5  g20766(.A(new_n23114), .B(new_n23113), .Y(new_n23115));
  nor_5  g20767(.A(new_n23115), .B(new_n23111), .Y(new_n23116));
  nor_5  g20768(.A(new_n23116), .B(new_n23109), .Y(new_n23117));
  nor_5  g20769(.A(new_n23117), .B(new_n23107), .Y(new_n23118));
  nor_5  g20770(.A(new_n23118), .B(new_n23105), .Y(new_n23119));
  or_6   g20771(.A(new_n23119), .B(new_n17981), .Y(new_n23120));
  or_6   g20772(.A(new_n17481), .B(new_n17476), .Y(new_n23121));
  nand_5 g20773(.A(new_n17482), .B(new_n17464), .Y(new_n23122));
  nand_5 g20774(.A(new_n23122), .B(new_n23121), .Y(new_n23123));
  nand_5 g20775(.A(new_n23110), .B(new_n23108), .Y(new_n23124));
  xor_4  g20776(.A(new_n23124), .B(new_n23115), .Y(new_n23125));
  not_8  g20777(.A(new_n23125), .Y(new_n23126));
  nor_5  g20778(.A(new_n23126), .B(new_n23123), .Y(new_n23127));
  xor_4  g20779(.A(new_n23125), .B(new_n23123), .Y(new_n23128));
  nor_5  g20780(.A(new_n23128), .B(new_n17938), .Y(new_n23129));
  or_6   g20781(.A(new_n23129), .B(new_n23127), .Y(new_n23130));
  nand_5 g20782(.A(new_n23106), .B(new_n23104), .Y(new_n23131));
  xor_4  g20783(.A(new_n23131), .B(new_n23117), .Y(new_n23132));
  nor_5  g20784(.A(new_n23132), .B(new_n23130), .Y(new_n23133));
  nand_5 g20785(.A(new_n23132), .B(new_n23130), .Y(new_n23134));
  not_8  g20786(.A(new_n23134), .Y(new_n23135));
  nor_5  g20787(.A(new_n23135), .B(new_n17937), .Y(new_n23136));
  nor_5  g20788(.A(new_n23136), .B(new_n23133), .Y(new_n23137));
  not_8  g20789(.A(new_n23137), .Y(new_n23138));
  nor_5  g20790(.A(new_n23138), .B(new_n23120), .Y(new_n23139));
  nand_5 g20791(.A(new_n23119), .B(new_n17981), .Y(new_n23140));
  nor_5  g20792(.A(new_n23140), .B(new_n23137), .Y(new_n23141));
  nor_5  g20793(.A(new_n23141), .B(new_n23139), .Y(new_n23142));
  nand_5 g20794(.A(new_n17975), .B(new_n11868), .Y(new_n23143));
  nand_5 g20795(.A(new_n17979), .B(new_n7786), .Y(new_n23144));
  nand_5 g20796(.A(new_n23144), .B(new_n23143), .Y(new_n23145));
  xor_4  g20797(.A(new_n23145), .B(new_n23142), .Y(po0623));
  xor_4  g20798(.A(new_n12695), .B(new_n12693), .Y(po0624));
  nand_5 g20799(.A(new_n16758), .B(new_n6338), .Y(new_n23148));
  nand_5 g20800(.A(new_n16759), .B(new_n16746), .Y(new_n23149));
  nand_5 g20801(.A(new_n23149), .B(new_n23148), .Y(new_n23150));
  nand_5 g20802(.A(new_n6373), .B(pi084), .Y(new_n23151));
  nand_5 g20803(.A(new_n16751), .B(new_n16748), .Y(new_n23152));
  nand_5 g20804(.A(new_n23152), .B(new_n23151), .Y(new_n23153));
  xor_4  g20805(.A(new_n23153), .B(new_n6385), .Y(new_n23154));
  xor_4  g20806(.A(new_n23154), .B(new_n12083), .Y(new_n23155));
  nand_5 g20807(.A(new_n16756), .B(new_n16752), .Y(new_n23156));
  or_6   g20808(.A(new_n16757), .B(new_n12085), .Y(new_n23157));
  nand_5 g20809(.A(new_n23157), .B(new_n23156), .Y(new_n23158));
  xor_4  g20810(.A(new_n23158), .B(new_n23155), .Y(new_n23159));
  not_8  g20811(.A(new_n23159), .Y(new_n23160));
  xor_4  g20812(.A(new_n23160), .B(new_n23150), .Y(po0625));
  xor_4  g20813(.A(new_n19500), .B(new_n19484), .Y(po0626));
  xor_4  g20814(.A(new_n21707), .B(new_n21700), .Y(po0627));
  xor_4  g20815(.A(pi574), .B(pi367), .Y(new_n23164));
  xor_4  g20816(.A(new_n23164), .B(new_n12969), .Y(po0628));
  xor_4  g20817(.A(new_n12366), .B(new_n8922), .Y(po0629));
  xor_4  g20818(.A(new_n19324), .B(new_n19304), .Y(po0630));
  nand_5 g20819(.A(new_n23063), .B(pi126), .Y(new_n23168));
  nand_5 g20820(.A(new_n23168), .B(new_n23062), .Y(new_n23169));
  xor_4  g20821(.A(new_n23169), .B(new_n8970), .Y(new_n23170));
  xor_4  g20822(.A(new_n23170), .B(pi197), .Y(new_n23171));
  nor_5  g20823(.A(pi571), .B(new_n11506), .Y(new_n23172));
  not_8  g20824(.A(new_n23172), .Y(new_n23173));
  nand_5 g20825(.A(pi571), .B(new_n11506), .Y(new_n23174));
  nand_5 g20826(.A(new_n23174), .B(new_n23173), .Y(new_n23175));
  xor_4  g20827(.A(new_n23175), .B(pi525), .Y(new_n23176));
  nor_5  g20828(.A(new_n22940), .B(new_n9648), .Y(new_n23177));
  nor_5  g20829(.A(new_n22947), .B(new_n22941), .Y(new_n23178));
  or_6   g20830(.A(new_n23178), .B(new_n23177), .Y(new_n23179));
  nand_5 g20831(.A(new_n22946), .B(new_n22942), .Y(new_n23180));
  nand_5 g20832(.A(new_n23180), .B(new_n22943), .Y(new_n23181));
  or_6   g20833(.A(pi596), .B(pi478), .Y(new_n23182));
  nand_5 g20834(.A(pi596), .B(pi478), .Y(new_n23183));
  nand_5 g20835(.A(new_n23183), .B(new_n23182), .Y(new_n23184));
  xnor_4 g20836(.A(new_n23184), .B(new_n23181), .Y(new_n23185));
  or_6   g20837(.A(new_n23185), .B(new_n23179), .Y(new_n23186));
  xor_4  g20838(.A(new_n23185), .B(new_n23179), .Y(new_n23187));
  nand_5 g20839(.A(new_n23187), .B(new_n21003), .Y(new_n23188));
  nand_5 g20840(.A(new_n23188), .B(new_n23186), .Y(new_n23189));
  xnor_4 g20841(.A(pi770), .B(pi594), .Y(new_n23190));
  nand_5 g20842(.A(new_n23183), .B(new_n23181), .Y(new_n23191));
  nand_5 g20843(.A(new_n23191), .B(new_n23182), .Y(new_n23192));
  xor_4  g20844(.A(new_n23192), .B(new_n23190), .Y(new_n23193));
  or_6   g20845(.A(new_n23193), .B(new_n23189), .Y(new_n23194));
  xor_4  g20846(.A(new_n23193), .B(new_n23189), .Y(new_n23195));
  nand_5 g20847(.A(new_n23195), .B(pi320), .Y(new_n23196));
  nand_5 g20848(.A(new_n23196), .B(new_n23194), .Y(new_n23197));
  nand_5 g20849(.A(new_n23197), .B(pi643), .Y(new_n23198));
  and_6  g20850(.A(pi770), .B(pi594), .Y(new_n23199));
  nor_5  g20851(.A(new_n23192), .B(new_n23190), .Y(new_n23200));
  nor_5  g20852(.A(new_n23200), .B(new_n23199), .Y(new_n23201));
  not_8  g20853(.A(pi347), .Y(new_n23202));
  xor_4  g20854(.A(pi817), .B(new_n23202), .Y(new_n23203));
  xor_4  g20855(.A(new_n23203), .B(new_n23201), .Y(new_n23204));
  xor_4  g20856(.A(new_n23197), .B(new_n10986), .Y(new_n23205));
  or_6   g20857(.A(new_n23205), .B(new_n23204), .Y(new_n23206));
  nand_5 g20858(.A(new_n23206), .B(new_n23198), .Y(new_n23207));
  xor_4  g20859(.A(pi808), .B(pi543), .Y(new_n23208));
  nor_5  g20860(.A(new_n11609), .B(new_n23202), .Y(new_n23209));
  nor_5  g20861(.A(new_n23203), .B(new_n23201), .Y(new_n23210));
  nor_5  g20862(.A(new_n23210), .B(new_n23209), .Y(new_n23211));
  xor_4  g20863(.A(new_n23211), .B(new_n23208), .Y(new_n23212));
  or_6   g20864(.A(new_n23212), .B(new_n23207), .Y(new_n23213));
  nand_5 g20865(.A(new_n23213), .B(pi627), .Y(new_n23214));
  nand_5 g20866(.A(new_n23212), .B(new_n23207), .Y(new_n23215));
  nand_5 g20867(.A(new_n23215), .B(new_n23214), .Y(new_n23216));
  xor_4  g20868(.A(pi179), .B(pi014), .Y(new_n23217));
  nand_5 g20869(.A(pi808), .B(pi543), .Y(new_n23218));
  not_8  g20870(.A(new_n23218), .Y(new_n23219));
  not_8  g20871(.A(new_n23208), .Y(new_n23220));
  nor_5  g20872(.A(new_n23211), .B(new_n23220), .Y(new_n23221));
  nor_5  g20873(.A(new_n23221), .B(new_n23219), .Y(new_n23222));
  xor_4  g20874(.A(new_n23222), .B(new_n23217), .Y(new_n23223));
  or_6   g20875(.A(new_n23223), .B(new_n23216), .Y(new_n23224));
  nand_5 g20876(.A(new_n23224), .B(pi199), .Y(new_n23225));
  nand_5 g20877(.A(new_n23223), .B(new_n23216), .Y(new_n23226));
  nand_5 g20878(.A(new_n23226), .B(new_n23225), .Y(new_n23227));
  nand_5 g20879(.A(pi179), .B(pi014), .Y(new_n23228));
  not_8  g20880(.A(new_n23228), .Y(new_n23229));
  not_8  g20881(.A(new_n23217), .Y(new_n23230));
  nor_5  g20882(.A(new_n23222), .B(new_n23230), .Y(new_n23231));
  nor_5  g20883(.A(new_n23231), .B(new_n23229), .Y(new_n23232));
  nor_5  g20884(.A(new_n23232), .B(new_n23227), .Y(new_n23233));
  not_8  g20885(.A(new_n23233), .Y(new_n23234));
  nand_5 g20886(.A(new_n23232), .B(new_n23227), .Y(new_n23235));
  nand_5 g20887(.A(new_n23235), .B(new_n23234), .Y(new_n23236));
  xor_4  g20888(.A(new_n23236), .B(new_n23176), .Y(new_n23237));
  not_8  g20889(.A(new_n23237), .Y(new_n23238));
  xor_4  g20890(.A(new_n23195), .B(pi320), .Y(new_n23239));
  xor_4  g20891(.A(new_n23187), .B(pi042), .Y(new_n23240));
  nor_5  g20892(.A(new_n23240), .B(new_n18612), .Y(new_n23241));
  xor_4  g20893(.A(new_n23240), .B(new_n18613), .Y(new_n23242));
  not_8  g20894(.A(new_n22954), .Y(new_n23243));
  nor_5  g20895(.A(new_n23243), .B(new_n22948), .Y(new_n23244));
  nor_5  g20896(.A(new_n22955), .B(new_n18628), .Y(new_n23245));
  or_6   g20897(.A(new_n23245), .B(new_n23244), .Y(new_n23246));
  nor_5  g20898(.A(new_n23246), .B(new_n23242), .Y(new_n23247));
  nor_5  g20899(.A(new_n23247), .B(new_n23241), .Y(new_n23248));
  nand_5 g20900(.A(new_n23248), .B(new_n23239), .Y(new_n23249));
  xnor_4 g20901(.A(new_n23248), .B(new_n23239), .Y(new_n23250));
  or_6   g20902(.A(new_n23250), .B(new_n18610), .Y(new_n23251));
  nand_5 g20903(.A(new_n23251), .B(new_n23249), .Y(new_n23252));
  xor_4  g20904(.A(new_n23205), .B(new_n23204), .Y(new_n23253));
  nand_5 g20905(.A(new_n23253), .B(new_n23252), .Y(new_n23254));
  xnor_4 g20906(.A(new_n23253), .B(new_n23252), .Y(new_n23255));
  or_6   g20907(.A(new_n23255), .B(new_n19358), .Y(new_n23256));
  nand_5 g20908(.A(new_n23256), .B(new_n23254), .Y(new_n23257));
  and_6  g20909(.A(new_n23215), .B(new_n23213), .Y(new_n23258));
  xor_4  g20910(.A(new_n23258), .B(new_n11072), .Y(new_n23259));
  not_8  g20911(.A(new_n23259), .Y(new_n23260));
  nand_5 g20912(.A(new_n23260), .B(new_n23257), .Y(new_n23261));
  xor_4  g20913(.A(new_n23259), .B(new_n23257), .Y(new_n23262));
  or_6   g20914(.A(new_n23262), .B(new_n23048), .Y(new_n23263));
  nand_5 g20915(.A(new_n23263), .B(new_n23261), .Y(new_n23264));
  and_6  g20916(.A(new_n23226), .B(new_n23224), .Y(new_n23265));
  xor_4  g20917(.A(new_n23265), .B(new_n11511), .Y(new_n23266));
  not_8  g20918(.A(new_n23266), .Y(new_n23267));
  nand_5 g20919(.A(new_n23267), .B(new_n23264), .Y(new_n23268));
  xor_4  g20920(.A(new_n23266), .B(new_n23264), .Y(new_n23269));
  or_6   g20921(.A(new_n23269), .B(new_n23035), .Y(new_n23270));
  nand_5 g20922(.A(new_n23270), .B(new_n23268), .Y(new_n23271));
  nand_5 g20923(.A(new_n23271), .B(new_n23238), .Y(new_n23272));
  xor_4  g20924(.A(new_n23271), .B(new_n23237), .Y(new_n23273));
  or_6   g20925(.A(new_n23273), .B(new_n23065), .Y(new_n23274));
  nand_5 g20926(.A(new_n23274), .B(new_n23272), .Y(new_n23275));
  or_6   g20927(.A(new_n23275), .B(new_n23171), .Y(new_n23276));
  xor_4  g20928(.A(new_n23275), .B(new_n23171), .Y(new_n23277));
  or_6   g20929(.A(new_n23236), .B(new_n23176), .Y(new_n23278));
  nand_5 g20930(.A(new_n23278), .B(new_n23234), .Y(new_n23279));
  nand_5 g20931(.A(new_n23173), .B(pi525), .Y(new_n23280));
  nand_5 g20932(.A(new_n23280), .B(new_n23174), .Y(new_n23281));
  nand_5 g20933(.A(new_n23281), .B(new_n23279), .Y(new_n23282));
  nor_5  g20934(.A(new_n23281), .B(new_n23235), .Y(new_n23283));
  nand_5 g20935(.A(new_n23172), .B(new_n11588), .Y(new_n23284));
  nor_5  g20936(.A(new_n23284), .B(new_n23233), .Y(new_n23285));
  nor_5  g20937(.A(new_n23285), .B(new_n23283), .Y(new_n23286));
  nand_5 g20938(.A(new_n23286), .B(new_n23282), .Y(new_n23287));
  xor_4  g20939(.A(new_n23287), .B(pi243), .Y(new_n23288));
  nand_5 g20940(.A(new_n11500), .B(pi084), .Y(new_n23289));
  nand_5 g20941(.A(pi340), .B(new_n16747), .Y(new_n23290));
  nand_5 g20942(.A(new_n23290), .B(new_n23289), .Y(new_n23291));
  xor_4  g20943(.A(new_n23291), .B(new_n23288), .Y(new_n23292));
  nand_5 g20944(.A(new_n23292), .B(new_n23277), .Y(new_n23293));
  nand_5 g20945(.A(new_n23293), .B(new_n23276), .Y(new_n23294));
  nand_5 g20946(.A(new_n23169), .B(new_n8970), .Y(new_n23295));
  nand_5 g20947(.A(new_n23170), .B(pi197), .Y(new_n23296));
  nand_5 g20948(.A(new_n23296), .B(new_n23295), .Y(new_n23297));
  xor_4  g20949(.A(new_n23297), .B(new_n11090), .Y(new_n23298));
  not_8  g20950(.A(new_n23298), .Y(new_n23299));
  not_8  g20951(.A(new_n23286), .Y(new_n23300));
  nand_5 g20952(.A(new_n23289), .B(new_n11594), .Y(new_n23301));
  nand_5 g20953(.A(new_n23301), .B(new_n23290), .Y(new_n23302));
  nand_5 g20954(.A(new_n23302), .B(new_n23300), .Y(new_n23303));
  nor_5  g20955(.A(new_n23290), .B(pi243), .Y(new_n23304));
  nand_5 g20956(.A(new_n23304), .B(new_n23282), .Y(new_n23305));
  nand_5 g20957(.A(new_n23305), .B(new_n23303), .Y(new_n23306));
  nor_5  g20958(.A(new_n23289), .B(new_n11594), .Y(new_n23307));
  nand_5 g20959(.A(new_n23307), .B(new_n23286), .Y(new_n23308));
  or_6   g20960(.A(new_n23302), .B(new_n23282), .Y(new_n23309));
  nand_5 g20961(.A(new_n23309), .B(new_n23308), .Y(new_n23310));
  nor_5  g20962(.A(new_n23310), .B(new_n23306), .Y(new_n23311));
  xor_4  g20963(.A(new_n23311), .B(new_n23299), .Y(new_n23312));
  xnor_4 g20964(.A(new_n23312), .B(new_n23294), .Y(po0631));
  xnor_4 g20965(.A(new_n20619), .B(new_n20618), .Y(po0632));
  xor_4  g20966(.A(new_n15616), .B(new_n15615), .Y(po0633));
  or_6   g20967(.A(new_n19177), .B(new_n19168), .Y(new_n23316));
  xor_4  g20968(.A(new_n23316), .B(new_n7393), .Y(po0634));
  xnor_4 g20969(.A(new_n20363), .B(new_n20362), .Y(po0635));
  not_8  g20970(.A(new_n22248), .Y(new_n23319));
  xor_4  g20971(.A(new_n23319), .B(new_n5679), .Y(new_n23320));
  or_6   g20972(.A(new_n15995), .B(new_n5682), .Y(new_n23321));
  or_6   g20973(.A(new_n10761), .B(new_n5728), .Y(new_n23322));
  nand_5 g20974(.A(new_n10795), .B(new_n5724), .Y(new_n23323));
  xor_4  g20975(.A(new_n10765), .B(new_n5723), .Y(new_n23324));
  nand_5 g20976(.A(new_n22871), .B(new_n5718), .Y(new_n23325));
  nand_5 g20977(.A(new_n23325), .B(new_n22866), .Y(new_n23326));
  nand_5 g20978(.A(new_n23326), .B(new_n23324), .Y(new_n23327));
  nand_5 g20979(.A(new_n23327), .B(new_n23323), .Y(new_n23328));
  xor_4  g20980(.A(new_n10761), .B(new_n5728), .Y(new_n23329));
  nand_5 g20981(.A(new_n23329), .B(new_n23328), .Y(new_n23330));
  nand_5 g20982(.A(new_n23330), .B(new_n23322), .Y(new_n23331));
  xor_4  g20983(.A(new_n15995), .B(new_n5682), .Y(new_n23332));
  nand_5 g20984(.A(new_n23332), .B(new_n23331), .Y(new_n23333));
  nand_5 g20985(.A(new_n23333), .B(new_n23321), .Y(new_n23334));
  xor_4  g20986(.A(new_n23334), .B(new_n23320), .Y(po0636));
  xnor_4 g20987(.A(new_n21380), .B(new_n20730), .Y(po0637));
  xor_4  g20988(.A(new_n18956), .B(new_n18955), .Y(po0638));
  nand_5 g20989(.A(new_n19199), .B(new_n19198), .Y(new_n23338));
  xor_4  g20990(.A(new_n23338), .B(new_n14056), .Y(po0639));
  nand_5 g20991(.A(new_n16066), .B(new_n7187), .Y(new_n23340));
  nand_5 g20992(.A(new_n22148), .B(new_n22145), .Y(new_n23341));
  nand_5 g20993(.A(new_n23341), .B(new_n23340), .Y(new_n23342));
  xor_4  g20994(.A(new_n23342), .B(new_n7545), .Y(new_n23343));
  or_6   g20995(.A(new_n22149), .B(new_n7551), .Y(new_n23344));
  not_8  g20996(.A(new_n23344), .Y(new_n23345));
  not_8  g20997(.A(new_n22150), .Y(new_n23346));
  nor_5  g20998(.A(new_n22153), .B(new_n23346), .Y(new_n23347));
  nor_5  g20999(.A(new_n23347), .B(new_n23345), .Y(new_n23348));
  xor_4  g21000(.A(new_n23348), .B(new_n23343), .Y(new_n23349));
  nand_5 g21001(.A(new_n8383), .B(pi293), .Y(new_n23350));
  nand_5 g21002(.A(new_n22157), .B(new_n22155), .Y(new_n23351));
  nand_5 g21003(.A(new_n23351), .B(new_n23350), .Y(new_n23352));
  nor_5  g21004(.A(new_n23352), .B(new_n23349), .Y(new_n23353));
  or_6   g21005(.A(new_n22158), .B(new_n22154), .Y(new_n23354));
  nand_5 g21006(.A(new_n22163), .B(new_n22159), .Y(new_n23355));
  nand_5 g21007(.A(new_n23355), .B(new_n23354), .Y(new_n23356));
  and_6  g21008(.A(new_n23356), .B(new_n23353), .Y(new_n23357));
  nand_5 g21009(.A(new_n23352), .B(new_n23349), .Y(new_n23358));
  nor_5  g21010(.A(new_n23358), .B(new_n23356), .Y(new_n23359));
  or_6   g21011(.A(new_n23359), .B(new_n23357), .Y(new_n23360));
  nand_5 g21012(.A(new_n23342), .B(new_n7545), .Y(new_n23361));
  nand_5 g21013(.A(new_n23348), .B(new_n23343), .Y(new_n23362));
  nand_5 g21014(.A(new_n23362), .B(new_n23361), .Y(new_n23363));
  xor_4  g21015(.A(new_n23363), .B(new_n23360), .Y(po0640));
  nand_5 g21016(.A(new_n8452), .B(new_n22874), .Y(new_n23365));
  or_6   g21017(.A(new_n8458), .B(new_n8447), .Y(new_n23366));
  nand_5 g21018(.A(new_n8459), .B(new_n8440), .Y(new_n23367));
  nand_5 g21019(.A(new_n23367), .B(new_n23366), .Y(new_n23368));
  nor_5  g21020(.A(new_n23368), .B(new_n23365), .Y(po0641));
  xnor_4 g21021(.A(new_n18886), .B(new_n18861), .Y(po0642));
  xor_4  g21022(.A(new_n23128), .B(new_n17938), .Y(po0643));
  xor_4  g21023(.A(new_n19866), .B(new_n15736), .Y(new_n23372));
  nand_5 g21024(.A(new_n22051), .B(new_n20985), .Y(new_n23373));
  not_8  g21025(.A(new_n23373), .Y(new_n23374));
  nor_5  g21026(.A(new_n21709), .B(new_n21696), .Y(new_n23375));
  nor_5  g21027(.A(new_n23375), .B(new_n23374), .Y(new_n23376));
  xor_4  g21028(.A(new_n23376), .B(new_n23372), .Y(po0644));
  xor_4  g21029(.A(new_n22366), .B(new_n5495), .Y(po0645));
  xor_4  g21030(.A(new_n14016), .B(new_n13005), .Y(po0646));
  xor_4  g21031(.A(new_n22007), .B(new_n17355), .Y(po0647));
  xor_4  g21032(.A(new_n18247), .B(new_n18241), .Y(po0648));
  xnor_4 g21033(.A(new_n18495), .B(new_n3076), .Y(po0649));
  xnor_4 g21034(.A(new_n8426), .B(new_n8405), .Y(po0650));
  xnor_4 g21035(.A(new_n19044), .B(new_n19043), .Y(po0651));
  xnor_4 g21036(.A(new_n22851), .B(new_n5707), .Y(po0652));
  nand_5 g21037(.A(new_n16382), .B(pi227), .Y(new_n23386));
  nand_5 g21038(.A(new_n23386), .B(new_n16381), .Y(new_n23387));
  or_6   g21039(.A(new_n23387), .B(new_n13710), .Y(new_n23388));
  nand_5 g21040(.A(new_n23387), .B(new_n13710), .Y(new_n23389));
  nand_5 g21041(.A(new_n23389), .B(new_n23388), .Y(new_n23390));
  xor_4  g21042(.A(new_n23390), .B(pi089), .Y(new_n23391));
  nor_5  g21043(.A(new_n23391), .B(new_n21613), .Y(new_n23392));
  nand_5 g21044(.A(new_n16441), .B(new_n16434), .Y(new_n23393));
  or_6   g21045(.A(new_n16443), .B(new_n16384), .Y(new_n23394));
  nand_5 g21046(.A(new_n23394), .B(new_n23393), .Y(new_n23395));
  xor_4  g21047(.A(new_n23391), .B(new_n21613), .Y(new_n23396));
  nand_5 g21048(.A(new_n23396), .B(new_n23395), .Y(new_n23397));
  not_8  g21049(.A(new_n23397), .Y(new_n23398));
  nor_5  g21050(.A(new_n23398), .B(new_n23392), .Y(new_n23399));
  nand_5 g21051(.A(new_n23388), .B(pi089), .Y(new_n23400));
  nand_5 g21052(.A(new_n23400), .B(new_n23389), .Y(new_n23401));
  nand_5 g21053(.A(new_n23401), .B(new_n13719), .Y(new_n23402));
  or_6   g21054(.A(new_n23401), .B(new_n13719), .Y(new_n23403));
  nand_5 g21055(.A(new_n23403), .B(new_n23402), .Y(new_n23404));
  xor_4  g21056(.A(new_n23404), .B(new_n22094), .Y(new_n23405));
  xor_4  g21057(.A(new_n23405), .B(new_n23399), .Y(po0653));
  xor_4  g21058(.A(new_n15916), .B(new_n10508), .Y(po0654));
  xnor_4 g21059(.A(new_n18649), .B(new_n18626), .Y(po0655));
  xnor_4 g21060(.A(new_n11471), .B(new_n4648), .Y(po0656));
  xor_4  g21061(.A(new_n18533), .B(new_n16101), .Y(po0657));
  xor_4  g21062(.A(new_n16516), .B(new_n16515), .Y(po0658));
  xnor_4 g21063(.A(new_n17058), .B(new_n17047), .Y(po0659));
  xnor_4 g21064(.A(new_n17598), .B(new_n17583), .Y(po0660));
  xor_4  g21065(.A(new_n10815), .B(new_n10814), .Y(po0661));
  xor_4  g21066(.A(new_n16490), .B(new_n15069), .Y(po0662));
  xor_4  g21067(.A(new_n16722), .B(new_n6177), .Y(po0663));
  xor_4  g21068(.A(new_n10387), .B(new_n10331), .Y(po0664));
  nand_5 g21069(.A(new_n22436), .B(new_n22437), .Y(new_n23418));
  xor_4  g21070(.A(new_n23418), .B(new_n3406), .Y(po0665));
  xor_4  g21071(.A(new_n6330), .B(new_n6328), .Y(po0666));
  xor_4  g21072(.A(new_n22781), .B(new_n22771), .Y(po0667));
  xor_4  g21073(.A(new_n10333), .B(new_n10332), .Y(new_n23422));
  xor_4  g21074(.A(new_n23422), .B(new_n10385), .Y(po0668));
  xor_4  g21075(.A(new_n22867), .B(new_n10782), .Y(po0669));
  xor_4  g21076(.A(new_n13511), .B(new_n7251), .Y(po0670));
  xor_4  g21077(.A(new_n9128), .B(new_n9127), .Y(po0671));
  xor_4  g21078(.A(new_n16866), .B(new_n8268), .Y(po0672));
  nand_5 g21079(.A(new_n6201), .B(pi154), .Y(new_n23428));
  nand_5 g21080(.A(new_n6165), .B(pi267), .Y(new_n23429));
  xor_4  g21081(.A(pi644), .B(new_n6429), .Y(new_n23430));
  nand_5 g21082(.A(pi312), .B(new_n8875), .Y(new_n23431));
  xor_4  g21083(.A(pi312), .B(new_n8875), .Y(new_n23432));
  nand_5 g21084(.A(new_n12096), .B(pi471), .Y(new_n23433));
  nand_5 g21085(.A(new_n19764), .B(new_n19759), .Y(new_n23434));
  nand_5 g21086(.A(new_n23434), .B(new_n23433), .Y(new_n23435));
  nand_5 g21087(.A(new_n23435), .B(new_n23432), .Y(new_n23436));
  nand_5 g21088(.A(new_n23436), .B(new_n23431), .Y(new_n23437));
  nand_5 g21089(.A(new_n23437), .B(new_n23430), .Y(new_n23438));
  nand_5 g21090(.A(new_n23438), .B(new_n23429), .Y(new_n23439));
  xor_4  g21091(.A(pi726), .B(new_n6556), .Y(new_n23440));
  nand_5 g21092(.A(new_n23440), .B(new_n23439), .Y(new_n23441));
  nand_5 g21093(.A(new_n23441), .B(new_n23428), .Y(new_n23442));
  nand_5 g21094(.A(new_n8868), .B(pi053), .Y(new_n23443));
  nand_5 g21095(.A(pi578), .B(new_n6554), .Y(new_n23444));
  nand_5 g21096(.A(new_n23444), .B(new_n23443), .Y(new_n23445));
  xor_4  g21097(.A(new_n23445), .B(new_n23442), .Y(new_n23446));
  xor_4  g21098(.A(new_n23446), .B(new_n19714), .Y(new_n23447));
  xor_4  g21099(.A(new_n23440), .B(new_n23439), .Y(new_n23448));
  or_6   g21100(.A(new_n23448), .B(new_n18285), .Y(new_n23449));
  not_8  g21101(.A(new_n18240), .Y(new_n23450));
  xor_4  g21102(.A(new_n23437), .B(new_n23430), .Y(new_n23451));
  or_6   g21103(.A(new_n23451), .B(new_n23450), .Y(new_n23452));
  xor_4  g21104(.A(new_n23451), .B(new_n23450), .Y(new_n23453));
  xnor_4 g21105(.A(new_n23435), .B(new_n23432), .Y(new_n23454));
  nor_5  g21106(.A(new_n23454), .B(new_n18262), .Y(new_n23455));
  or_6   g21107(.A(new_n19765), .B(new_n18258), .Y(new_n23456));
  nand_5 g21108(.A(new_n19777), .B(new_n19766), .Y(new_n23457));
  nand_5 g21109(.A(new_n23457), .B(new_n23456), .Y(new_n23458));
  xor_4  g21110(.A(new_n23454), .B(new_n18264), .Y(new_n23459));
  nor_5  g21111(.A(new_n23459), .B(new_n23458), .Y(new_n23460));
  or_6   g21112(.A(new_n23460), .B(new_n23455), .Y(new_n23461));
  not_8  g21113(.A(new_n23461), .Y(new_n23462));
  nand_5 g21114(.A(new_n23462), .B(new_n23453), .Y(new_n23463));
  nand_5 g21115(.A(new_n23463), .B(new_n23452), .Y(new_n23464));
  xor_4  g21116(.A(new_n23448), .B(new_n18285), .Y(new_n23465));
  nand_5 g21117(.A(new_n23465), .B(new_n23464), .Y(new_n23466));
  nand_5 g21118(.A(new_n23466), .B(new_n23449), .Y(new_n23467));
  xnor_4 g21119(.A(new_n23467), .B(new_n23447), .Y(po0673));
  xnor_4 g21120(.A(new_n21705), .B(new_n21702), .Y(po0674));
  xor_4  g21121(.A(new_n10616), .B(new_n10615), .Y(po0675));
  nor_5  g21122(.A(new_n8711), .B(new_n8710), .Y(new_n23471));
  xor_4  g21123(.A(new_n23471), .B(new_n8712), .Y(po0676));
  nand_5 g21124(.A(new_n5735), .B(new_n5734), .Y(new_n23473));
  xnor_4 g21125(.A(new_n23473), .B(new_n5737), .Y(po0677));
  xnor_4 g21126(.A(new_n7669), .B(new_n7645), .Y(po0678));
  nor_5  g21127(.A(new_n5553), .B(new_n5496), .Y(new_n23476));
  nand_5 g21128(.A(new_n23476), .B(new_n5630), .Y(new_n23477));
  not_8  g21129(.A(new_n22337), .Y(new_n23478));
  not_8  g21130(.A(new_n5743), .Y(new_n23479));
  or_6   g21131(.A(new_n23319), .B(new_n5679), .Y(new_n23480));
  nand_5 g21132(.A(new_n23334), .B(new_n23320), .Y(new_n23481));
  nand_5 g21133(.A(new_n23481), .B(new_n23480), .Y(new_n23482));
  not_8  g21134(.A(new_n23482), .Y(new_n23483));
  nand_5 g21135(.A(new_n23483), .B(new_n23479), .Y(new_n23484));
  nor_5  g21136(.A(new_n23484), .B(new_n23478), .Y(new_n23485));
  nor_5  g21137(.A(new_n23483), .B(new_n23479), .Y(new_n23486));
  not_8  g21138(.A(new_n22245), .Y(new_n23487));
  or_6   g21139(.A(new_n23487), .B(new_n18759), .Y(new_n23488));
  nor_5  g21140(.A(new_n23488), .B(new_n23486), .Y(new_n23489));
  nor_5  g21141(.A(new_n23489), .B(new_n23485), .Y(new_n23490));
  and_6  g21142(.A(new_n23490), .B(new_n9886), .Y(new_n23491));
  nand_5 g21143(.A(new_n23486), .B(new_n23478), .Y(new_n23492));
  nor_5  g21144(.A(new_n22245), .B(new_n18760), .Y(new_n23493));
  nand_5 g21145(.A(new_n23493), .B(new_n23484), .Y(new_n23494));
  nand_5 g21146(.A(new_n23494), .B(new_n23492), .Y(new_n23495));
  nor_5  g21147(.A(new_n23495), .B(new_n23491), .Y(new_n23496));
  nand_5 g21148(.A(new_n23496), .B(new_n5633), .Y(new_n23497));
  nand_5 g21149(.A(new_n23497), .B(new_n23477), .Y(po0680));
  xor_4  g21150(.A(new_n8612), .B(new_n8615), .Y(po0681));
  xor_4  g21151(.A(new_n17261), .B(new_n17246), .Y(po0682));
  nor_5  g21152(.A(new_n19866), .B(new_n20985), .Y(new_n23501));
  nor_5  g21153(.A(new_n23376), .B(new_n23372), .Y(new_n23502));
  nor_5  g21154(.A(new_n23502), .B(new_n23501), .Y(po0683));
  xnor_4 g21155(.A(new_n21462), .B(new_n21420), .Y(po0684));
  nor_5  g21156(.A(new_n21303), .B(new_n12083), .Y(new_n23505));
  nand_5 g21157(.A(new_n21305), .B(new_n21300), .Y(new_n23506));
  or_6   g21158(.A(new_n23506), .B(new_n17350), .Y(new_n23507));
  nand_5 g21159(.A(new_n23507), .B(new_n23505), .Y(new_n23508));
  nor_5  g21160(.A(new_n21304), .B(new_n17353), .Y(new_n23509));
  nor_5  g21161(.A(new_n23509), .B(new_n17351), .Y(new_n23510));
  nand_5 g21162(.A(new_n23510), .B(new_n23506), .Y(new_n23511));
  and_6  g21163(.A(new_n23511), .B(new_n23508), .Y(po0685));
  xnor_4 g21164(.A(new_n22460), .B(new_n22456), .Y(po0686));
  nor_5  g21165(.A(new_n16094), .B(pi111), .Y(new_n23514));
  nor_5  g21166(.A(new_n16095), .B(new_n16065), .Y(new_n23515));
  or_6   g21167(.A(new_n23515), .B(new_n23514), .Y(new_n23516));
  nor_5  g21168(.A(new_n23516), .B(new_n22115), .Y(new_n23517));
  not_8  g21169(.A(new_n23517), .Y(new_n23518));
  nand_5 g21170(.A(new_n23516), .B(new_n22115), .Y(new_n23519));
  nand_5 g21171(.A(new_n23519), .B(new_n23518), .Y(new_n23520));
  not_8  g21172(.A(new_n23520), .Y(new_n23521));
  not_8  g21173(.A(new_n22906), .Y(new_n23522));
  nand_5 g21174(.A(new_n16230), .B(new_n22897), .Y(new_n23523));
  nand_5 g21175(.A(new_n23523), .B(new_n23522), .Y(new_n23524));
  nand_5 g21176(.A(new_n16229), .B(new_n16224), .Y(new_n23525));
  nand_5 g21177(.A(new_n23525), .B(new_n22906), .Y(new_n23526));
  nand_5 g21178(.A(new_n23526), .B(new_n23524), .Y(new_n23527));
  nand_5 g21179(.A(new_n16214), .B(pi425), .Y(new_n23528));
  nand_5 g21180(.A(new_n23528), .B(new_n16213), .Y(new_n23529));
  nor_5  g21181(.A(new_n23529), .B(new_n23527), .Y(new_n23530));
  nand_5 g21182(.A(new_n23525), .B(pi425), .Y(new_n23531));
  or_6   g21183(.A(new_n23531), .B(new_n16213), .Y(new_n23532));
  nand_5 g21184(.A(new_n23523), .B(new_n22896), .Y(new_n23533));
  or_6   g21185(.A(new_n23533), .B(new_n16214), .Y(new_n23534));
  nand_5 g21186(.A(new_n23534), .B(new_n23532), .Y(new_n23535));
  and_6  g21187(.A(new_n23535), .B(new_n22906), .Y(new_n23536));
  nor_5  g21188(.A(new_n23536), .B(new_n23530), .Y(new_n23537));
  nand_5 g21189(.A(new_n23525), .B(new_n23523), .Y(new_n23538));
  or_6   g21190(.A(new_n23538), .B(new_n22906), .Y(new_n23539));
  nor_5  g21191(.A(new_n23539), .B(new_n23535), .Y(new_n23540));
  and_6  g21192(.A(new_n23538), .B(new_n23527), .Y(new_n23541));
  and_6  g21193(.A(new_n23541), .B(new_n23529), .Y(new_n23542));
  nor_5  g21194(.A(new_n23542), .B(new_n23540), .Y(new_n23543));
  nand_5 g21195(.A(new_n23543), .B(new_n23537), .Y(new_n23544));
  nand_5 g21196(.A(new_n23544), .B(new_n23521), .Y(new_n23545));
  nand_5 g21197(.A(new_n23545), .B(new_n23518), .Y(new_n23546));
  not_8  g21198(.A(new_n23546), .Y(new_n23547));
  nand_5 g21199(.A(new_n23537), .B(new_n23524), .Y(new_n23548));
  nand_5 g21200(.A(new_n23548), .B(new_n23532), .Y(new_n23549));
  xor_4  g21201(.A(new_n23549), .B(new_n23547), .Y(po0687));
  xor_4  g21202(.A(new_n11065), .B(new_n11032), .Y(po0688));
  not_8  g21203(.A(new_n15668), .Y(new_n23552));
  nand_5 g21204(.A(pi247), .B(new_n12560), .Y(new_n23553));
  not_8  g21205(.A(new_n23553), .Y(new_n23554));
  xor_4  g21206(.A(pi247), .B(new_n12560), .Y(new_n23555));
  not_8  g21207(.A(new_n23555), .Y(new_n23556));
  nand_5 g21208(.A(new_n8865), .B(pi112), .Y(new_n23557));
  xor_4  g21209(.A(pi205), .B(new_n12563), .Y(new_n23558));
  nand_5 g21210(.A(new_n23444), .B(new_n23442), .Y(new_n23559));
  nand_5 g21211(.A(new_n23559), .B(new_n23443), .Y(new_n23560));
  nand_5 g21212(.A(new_n23560), .B(new_n23558), .Y(new_n23561));
  nand_5 g21213(.A(new_n23561), .B(new_n23557), .Y(new_n23562));
  nor_5  g21214(.A(new_n23562), .B(new_n23556), .Y(new_n23563));
  nor_5  g21215(.A(new_n23563), .B(new_n23554), .Y(new_n23564));
  nor_5  g21216(.A(new_n23564), .B(new_n15622), .Y(new_n23565));
  nor_5  g21217(.A(new_n23565), .B(new_n23552), .Y(new_n23566));
  not_8  g21218(.A(new_n20995), .Y(new_n23567));
  xor_4  g21219(.A(new_n23564), .B(new_n15670), .Y(new_n23568));
  nand_5 g21220(.A(new_n23568), .B(new_n20970), .Y(new_n23569));
  xnor_4 g21221(.A(new_n23560), .B(new_n23558), .Y(new_n23570));
  nor_5  g21222(.A(new_n23570), .B(new_n19711), .Y(new_n23571));
  nor_5  g21223(.A(new_n23446), .B(new_n19713), .Y(new_n23572));
  nor_5  g21224(.A(new_n23467), .B(new_n23447), .Y(new_n23573));
  nor_5  g21225(.A(new_n23573), .B(new_n23572), .Y(new_n23574));
  xor_4  g21226(.A(new_n23570), .B(new_n19712), .Y(new_n23575));
  nor_5  g21227(.A(new_n23575), .B(new_n23574), .Y(new_n23576));
  or_6   g21228(.A(new_n23576), .B(new_n23571), .Y(new_n23577));
  not_8  g21229(.A(new_n19705), .Y(new_n23578));
  xor_4  g21230(.A(new_n23562), .B(new_n23556), .Y(new_n23579));
  nand_5 g21231(.A(new_n23579), .B(new_n23578), .Y(new_n23580));
  nand_5 g21232(.A(new_n23580), .B(new_n23577), .Y(new_n23581));
  or_6   g21233(.A(new_n23579), .B(new_n23578), .Y(new_n23582));
  nand_5 g21234(.A(new_n23582), .B(new_n23581), .Y(new_n23583));
  xor_4  g21235(.A(new_n23568), .B(new_n20970), .Y(new_n23584));
  nand_5 g21236(.A(new_n23584), .B(new_n23583), .Y(new_n23585));
  nand_5 g21237(.A(new_n23585), .B(new_n23569), .Y(new_n23586));
  nand_5 g21238(.A(new_n23586), .B(new_n23567), .Y(new_n23587));
  nand_5 g21239(.A(new_n23587), .B(new_n23566), .Y(new_n23588));
  not_8  g21240(.A(new_n23566), .Y(new_n23589));
  or_6   g21241(.A(new_n23586), .B(new_n23567), .Y(new_n23590));
  nand_5 g21242(.A(new_n23590), .B(new_n23589), .Y(new_n23591));
  nand_5 g21243(.A(new_n23591), .B(new_n23588), .Y(new_n23592));
  xnor_4 g21244(.A(new_n23592), .B(new_n22185), .Y(po0689));
  xor_4  g21245(.A(new_n7443), .B(new_n16924), .Y(po0690));
  xnor_4 g21246(.A(new_n11829), .B(new_n11828), .Y(po0691));
  xnor_4 g21247(.A(new_n20616), .B(new_n20590), .Y(po0692));
  xnor_4 g21248(.A(new_n8257), .B(new_n8233), .Y(po0693));
  xnor_4 g21249(.A(new_n13474), .B(new_n13454), .Y(po0694));
  xnor_4 g21250(.A(new_n6393), .B(new_n6371), .Y(po0695));
  xnor_4 g21251(.A(new_n10219), .B(new_n10203), .Y(po0696));
  xnor_4 g21252(.A(new_n3679), .B(new_n3677), .Y(po0697));
  xor_4  g21253(.A(new_n18460), .B(new_n6900), .Y(po0698));
  xor_4  g21254(.A(new_n15629), .B(new_n18243), .Y(po0699));
  xor_4  g21255(.A(new_n17303), .B(new_n7944), .Y(po0700));
  xor_4  g21256(.A(pi832), .B(pi569), .Y(new_n23605));
  xor_4  g21257(.A(new_n23605), .B(new_n2522), .Y(po0701));
  xnor_4 g21258(.A(new_n7151), .B(new_n7149), .Y(po0702));
  xnor_4 g21259(.A(new_n16209), .B(new_n16197), .Y(po0703));
  xor_4  g21260(.A(new_n9832), .B(new_n9830), .Y(po0704));
  or_6   g21261(.A(new_n20946), .B(new_n20942), .Y(new_n23610));
  xor_4  g21262(.A(new_n23610), .B(new_n20945), .Y(po0705));
  nand_5 g21263(.A(new_n21151), .B(new_n21097), .Y(new_n23612));
  xor_4  g21264(.A(new_n23612), .B(new_n2755), .Y(po0706));
  xor_4  g21265(.A(new_n9348), .B(new_n22328), .Y(po0707));
  xor_4  g21266(.A(new_n7177), .B(new_n7115), .Y(po0708));
  nand_5 g21267(.A(new_n23590), .B(new_n23587), .Y(new_n23616));
  xor_4  g21268(.A(new_n23616), .B(new_n23589), .Y(po0709));
  xor_4  g21269(.A(new_n17888), .B(new_n17887), .Y(po0710));
  xnor_4 g21270(.A(new_n16432), .B(new_n16431), .Y(po0711));
  nor_5  g21271(.A(new_n18524), .B(new_n20014), .Y(new_n23620));
  nor_5  g21272(.A(new_n18525), .B(pi216), .Y(new_n23621));
  nor_5  g21273(.A(new_n23621), .B(new_n23620), .Y(new_n23622));
  nand_5 g21274(.A(new_n23622), .B(new_n20011), .Y(new_n23623));
  nor_5  g21275(.A(new_n23622), .B(new_n20011), .Y(new_n23624));
  not_8  g21276(.A(new_n23624), .Y(new_n23625));
  nand_5 g21277(.A(new_n18550), .B(new_n16096), .Y(new_n23626));
  or_6   g21278(.A(new_n18551), .B(new_n18526), .Y(new_n23627));
  nand_5 g21279(.A(new_n23627), .B(new_n23626), .Y(new_n23628));
  not_8  g21280(.A(new_n23628), .Y(new_n23629));
  nand_5 g21281(.A(new_n23629), .B(new_n23625), .Y(new_n23630));
  nand_5 g21282(.A(new_n23630), .B(new_n23623), .Y(new_n23631));
  or_6   g21283(.A(new_n23631), .B(new_n23519), .Y(new_n23632));
  not_8  g21284(.A(new_n23632), .Y(new_n23633));
  nand_5 g21285(.A(new_n23628), .B(new_n23624), .Y(new_n23634));
  nand_5 g21286(.A(new_n23634), .B(new_n23518), .Y(new_n23635));
  nor_5  g21287(.A(new_n23635), .B(new_n23633), .Y(po0712));
  xnor_4 g21288(.A(new_n21235), .B(new_n21234), .Y(po0713));
  nand_5 g21289(.A(new_n22635), .B(new_n22625), .Y(new_n23638));
  nand_5 g21290(.A(new_n22636), .B(new_n17664), .Y(new_n23639));
  nand_5 g21291(.A(new_n23639), .B(new_n23638), .Y(new_n23640));
  nor_5  g21292(.A(new_n22629), .B(new_n4863), .Y(new_n23641));
  and_6  g21293(.A(new_n22633), .B(new_n22630), .Y(new_n23642));
  nor_5  g21294(.A(new_n23642), .B(new_n23641), .Y(new_n23643));
  nand_5 g21295(.A(new_n23643), .B(new_n23640), .Y(new_n23644));
  not_8  g21296(.A(new_n4868), .Y(new_n23645));
  nor_5  g21297(.A(new_n23643), .B(new_n23640), .Y(new_n23646));
  nor_5  g21298(.A(new_n23646), .B(new_n23645), .Y(new_n23647));
  nand_5 g21299(.A(pi661), .B(pi124), .Y(new_n23648));
  or_6   g21300(.A(new_n22628), .B(new_n21610), .Y(new_n23649));
  nand_5 g21301(.A(new_n23649), .B(new_n23648), .Y(new_n23650));
  or_6   g21302(.A(new_n23650), .B(new_n18950), .Y(new_n23651));
  nor_5  g21303(.A(new_n23651), .B(new_n23647), .Y(new_n23652));
  not_8  g21304(.A(new_n23646), .Y(new_n23653));
  nand_5 g21305(.A(new_n23650), .B(new_n18950), .Y(new_n23654));
  nand_5 g21306(.A(new_n23654), .B(new_n23645), .Y(new_n23655));
  nor_5  g21307(.A(new_n23655), .B(new_n23653), .Y(new_n23656));
  or_6   g21308(.A(new_n23656), .B(new_n23652), .Y(new_n23657));
  and_6  g21309(.A(new_n23657), .B(new_n23644), .Y(po0714));
  xor_4  g21310(.A(new_n13104), .B(new_n13102), .Y(po0715));
  xnor_4 g21311(.A(new_n21173), .B(new_n21172), .Y(po0716));
  not_8  g21312(.A(new_n18829), .Y(new_n23661));
  nand_5 g21313(.A(new_n22100), .B(new_n23661), .Y(new_n23662));
  nor_5  g21314(.A(new_n22106), .B(new_n18836), .Y(new_n23663));
  nand_5 g21315(.A(new_n23090), .B(new_n23087), .Y(new_n23664));
  not_8  g21316(.A(new_n23664), .Y(new_n23665));
  nor_5  g21317(.A(new_n23665), .B(new_n23663), .Y(new_n23666));
  xor_4  g21318(.A(new_n22100), .B(new_n18829), .Y(new_n23667));
  not_8  g21319(.A(new_n23667), .Y(new_n23668));
  nand_5 g21320(.A(new_n23668), .B(new_n23666), .Y(new_n23669));
  nand_5 g21321(.A(new_n23669), .B(new_n23662), .Y(po0717));
  xnor_4 g21322(.A(new_n10620), .B(new_n10585), .Y(po0718));
  xor_4  g21323(.A(new_n11334), .B(new_n11326), .Y(po0719));
  xnor_4 g21324(.A(new_n5819), .B(new_n5818), .Y(po0720));
  xor_4  g21325(.A(new_n13456), .B(new_n7924), .Y(po0721));
  xor_4  g21326(.A(new_n6513), .B(new_n4598), .Y(po0722));
  xor_4  g21327(.A(new_n14781), .B(new_n14780), .Y(po0723));
  nand_5 g21328(.A(pi358), .B(new_n16941), .Y(new_n23677));
  nand_5 g21329(.A(new_n16959), .B(new_n16942), .Y(new_n23678));
  nand_5 g21330(.A(new_n23678), .B(new_n23677), .Y(new_n23679));
  xor_4  g21331(.A(new_n23679), .B(new_n15107), .Y(new_n23680));
  or_6   g21332(.A(new_n16960), .B(new_n15090), .Y(new_n23681));
  nand_5 g21333(.A(new_n16982), .B(new_n16961), .Y(new_n23682));
  nand_5 g21334(.A(new_n23682), .B(new_n23681), .Y(new_n23683));
  xnor_4 g21335(.A(new_n23683), .B(new_n23680), .Y(po0724));
  xor_4  g21336(.A(pi216), .B(new_n21895), .Y(new_n23685));
  nand_5 g21337(.A(pi721), .B(new_n16220), .Y(new_n23686));
  nand_5 g21338(.A(new_n21415), .B(new_n21385), .Y(new_n23687));
  nand_5 g21339(.A(new_n23687), .B(new_n23686), .Y(new_n23688));
  xnor_4 g21340(.A(new_n23688), .B(new_n23685), .Y(new_n23689));
  or_6   g21341(.A(new_n23689), .B(new_n20042), .Y(new_n23690));
  not_8  g21342(.A(new_n21416), .Y(new_n23691));
  nor_5  g21343(.A(new_n23691), .B(new_n14631), .Y(new_n23692));
  nor_5  g21344(.A(new_n21464), .B(new_n21417), .Y(new_n23693));
  or_6   g21345(.A(new_n23693), .B(new_n23692), .Y(new_n23694));
  xor_4  g21346(.A(new_n23689), .B(new_n20042), .Y(new_n23695));
  nand_5 g21347(.A(new_n23695), .B(new_n23694), .Y(new_n23696));
  nand_5 g21348(.A(new_n23696), .B(new_n23690), .Y(new_n23697));
  or_6   g21349(.A(new_n23697), .B(new_n20027), .Y(new_n23698));
  nand_5 g21350(.A(new_n23697), .B(new_n20027), .Y(new_n23699));
  nand_5 g21351(.A(new_n23699), .B(new_n23698), .Y(new_n23700));
  nand_5 g21352(.A(new_n16216), .B(pi142), .Y(new_n23701));
  nand_5 g21353(.A(new_n23688), .B(new_n23685), .Y(new_n23702));
  nand_5 g21354(.A(new_n23702), .B(new_n23701), .Y(new_n23703));
  not_8  g21355(.A(new_n23703), .Y(new_n23704));
  xor_4  g21356(.A(new_n23704), .B(new_n23700), .Y(po0725));
  xor_4  g21357(.A(new_n20086), .B(new_n16834), .Y(po0726));
  xor_4  g21358(.A(new_n17985), .B(new_n13818), .Y(po0727));
  xor_4  g21359(.A(new_n15568), .B(new_n13119), .Y(po0728));
  xnor_4 g21360(.A(new_n18101), .B(new_n18100), .Y(po0729));
  xor_4  g21361(.A(new_n7159), .B(new_n7127), .Y(po0730));
  xor_4  g21362(.A(new_n18123), .B(new_n18110), .Y(po0731));
  xnor_4 g21363(.A(new_n20122), .B(new_n20117), .Y(po0732));
  xnor_4 g21364(.A(new_n6187), .B(new_n6186), .Y(po0733));
  xnor_4 g21365(.A(new_n19947), .B(new_n17242), .Y(po0734));
  xor_4  g21366(.A(new_n20623), .B(new_n20581), .Y(po0735));
  xor_4  g21367(.A(new_n21369), .B(new_n18166), .Y(po0736));
  xor_4  g21368(.A(new_n14774), .B(new_n14741), .Y(po0737));
  xnor_4 g21369(.A(new_n14897), .B(new_n14880), .Y(po0738));
  xnor_4 g21370(.A(new_n10376), .B(new_n10346), .Y(po0739));
  xor_4  g21371(.A(new_n19754), .B(new_n9132), .Y(po0740));
  xnor_4 g21372(.A(new_n13363), .B(new_n13342), .Y(po0741));
  nor_5  g21373(.A(new_n22448), .B(new_n22440), .Y(new_n23722));
  xnor_4 g21374(.A(new_n23722), .B(new_n3331), .Y(po0742));
  xor_4  g21375(.A(new_n21792), .B(new_n9763), .Y(po0743));
  xor_4  g21376(.A(new_n7951), .B(new_n7950), .Y(po0744));
  xor_4  g21377(.A(new_n16462), .B(new_n5363), .Y(po0745));
  xor_4  g21378(.A(new_n5437), .B(new_n5436), .Y(po0746));
  nor_5  g21379(.A(new_n22827), .B(new_n22826), .Y(new_n23728));
  nor_5  g21380(.A(new_n21803), .B(new_n21071), .Y(new_n23729));
  nor_5  g21381(.A(new_n23729), .B(new_n21062), .Y(new_n23730));
  not_8  g21382(.A(new_n23730), .Y(new_n23731));
  nor_5  g21383(.A(new_n23731), .B(new_n23728), .Y(new_n23732));
  not_8  g21384(.A(new_n23732), .Y(new_n23733));
  nor_5  g21385(.A(new_n23733), .B(new_n21681), .Y(new_n23734));
  nor_5  g21386(.A(new_n23732), .B(new_n21683), .Y(new_n23735));
  nor_5  g21387(.A(new_n23735), .B(new_n23734), .Y(new_n23736));
  not_8  g21388(.A(new_n11524), .Y(new_n23737));
  xor_4  g21389(.A(new_n23732), .B(new_n21812), .Y(new_n23738));
  or_6   g21390(.A(new_n23738), .B(new_n23737), .Y(new_n23739));
  nand_5 g21391(.A(new_n23738), .B(new_n23737), .Y(new_n23740));
  nand_5 g21392(.A(new_n22828), .B(new_n22823), .Y(new_n23741));
  nand_5 g21393(.A(new_n22832), .B(new_n22829), .Y(new_n23742));
  nand_5 g21394(.A(new_n23742), .B(new_n23741), .Y(new_n23743));
  nand_5 g21395(.A(new_n23743), .B(new_n23740), .Y(new_n23744));
  nand_5 g21396(.A(new_n23744), .B(new_n23739), .Y(new_n23745));
  and_6  g21397(.A(new_n23745), .B(new_n23736), .Y(new_n23746));
  or_6   g21398(.A(new_n23746), .B(new_n23734), .Y(po0747));
  xnor_4 g21399(.A(new_n12325), .B(new_n6522), .Y(po0748));
  xnor_4 g21400(.A(new_n12711), .B(new_n12684), .Y(po0749));
  xor_4  g21401(.A(new_n20826), .B(new_n6055), .Y(po0750));
  xor_4  g21402(.A(new_n22350), .B(new_n21834), .Y(new_n23751));
  or_6   g21403(.A(new_n22259), .B(new_n17559), .Y(new_n23752));
  nand_5 g21404(.A(new_n22286), .B(new_n22260), .Y(new_n23753));
  nand_5 g21405(.A(new_n23753), .B(new_n23752), .Y(new_n23754));
  xor_4  g21406(.A(new_n23754), .B(new_n23751), .Y(po0751));
  xor_4  g21407(.A(new_n5172), .B(new_n5150), .Y(po0752));
  xnor_4 g21408(.A(new_n4478), .B(new_n4462), .Y(po0753));
  xor_4  g21409(.A(new_n6197), .B(new_n6175), .Y(po0754));
  xnor_4 g21410(.A(new_n6034), .B(new_n6033), .Y(po0755));
  xor_4  g21411(.A(new_n23262), .B(new_n23054), .Y(po0756));
  xor_4  g21412(.A(new_n5004), .B(new_n5002), .Y(po0757));
  nand_5 g21413(.A(new_n17636), .B(new_n17637), .Y(new_n23762));
  xor_4  g21414(.A(new_n23762), .B(new_n8600), .Y(po0758));
  xor_4  g21415(.A(new_n8249), .B(new_n8248), .Y(po0759));
  xor_4  g21416(.A(new_n20369), .B(new_n20368), .Y(po0760));
  xor_4  g21417(.A(new_n19959), .B(new_n17231), .Y(po0761));
  xnor_4 g21418(.A(new_n2793), .B(new_n2792), .Y(po0763));
  xor_4  g21419(.A(new_n14595), .B(new_n14592), .Y(po0764));
  xor_4  g21420(.A(new_n17646), .B(new_n8635), .Y(po0765));
  xor_4  g21421(.A(new_n16035), .B(new_n11453), .Y(po0766));
  xor_4  g21422(.A(new_n18069), .B(new_n7821), .Y(po0767));
  nand_5 g21423(.A(new_n19723), .B(new_n19722), .Y(new_n23772));
  xor_4  g21424(.A(new_n23772), .B(new_n15426), .Y(po0768));
  xnor_4 g21425(.A(new_n11833), .B(new_n11806), .Y(po0769));
  xnor_4 g21426(.A(new_n12066), .B(new_n12065), .Y(po0770));
  xor_4  g21427(.A(new_n21880), .B(new_n9070), .Y(po0771));
  xnor_4 g21428(.A(new_n17462), .B(new_n17461), .Y(po0772));
  xor_4  g21429(.A(new_n19157), .B(new_n19154), .Y(po0773));
  xor_4  g21430(.A(new_n6693), .B(new_n3342), .Y(po0774));
  xnor_4 g21431(.A(new_n8951), .B(new_n8950), .Y(po0775));
  xor_4  g21432(.A(new_n12260), .B(new_n11358), .Y(po0776));
  xor_4  g21433(.A(new_n19973), .B(new_n17222), .Y(po0777));
  not_8  g21434(.A(new_n22652), .Y(new_n23783));
  nand_5 g21435(.A(new_n23679), .B(new_n15107), .Y(new_n23784));
  nor_5  g21436(.A(new_n23683), .B(new_n23784), .Y(new_n23785));
  nor_5  g21437(.A(new_n23679), .B(new_n15107), .Y(new_n23786));
  nand_5 g21438(.A(new_n23683), .B(new_n23786), .Y(new_n23787));
  not_8  g21439(.A(new_n23787), .Y(new_n23788));
  nor_5  g21440(.A(new_n23788), .B(new_n23785), .Y(new_n23789));
  xor_4  g21441(.A(new_n23789), .B(new_n23783), .Y(po0778));
  xnor_4 g21442(.A(new_n21592), .B(new_n21586), .Y(po0779));
  nand_5 g21443(.A(new_n16742), .B(new_n16741), .Y(new_n23792));
  xor_4  g21444(.A(new_n23792), .B(new_n6271), .Y(po0780));
  xor_4  g21445(.A(new_n5431), .B(new_n5429), .Y(po0781));
  xnor_4 g21446(.A(new_n16931), .B(new_n16927), .Y(po0782));
  xor_4  g21447(.A(new_n13705), .B(new_n13703), .Y(po0783));
  xnor_4 g21448(.A(new_n5707), .B(new_n5705), .Y(po0784));
  xor_4  g21449(.A(new_n9466), .B(new_n9465), .Y(po0785));
  xnor_4 g21450(.A(new_n8422), .B(new_n8412), .Y(po0786));
  xor_4  g21451(.A(new_n23292), .B(new_n23277), .Y(po0787));
  xor_4  g21452(.A(new_n23326), .B(new_n23324), .Y(po0788));
  xnor_4 g21453(.A(new_n12656), .B(new_n12654), .Y(po0789));
  xnor_4 g21454(.A(new_n18647), .B(new_n18646), .Y(po0790));
  nor_5  g21455(.A(new_n21888), .B(new_n21883), .Y(new_n23804));
  nor_5  g21456(.A(new_n21887), .B(new_n21884), .Y(new_n23805));
  nor_5  g21457(.A(new_n23805), .B(new_n23804), .Y(new_n23806));
  nor_5  g21458(.A(new_n23806), .B(new_n11860), .Y(po0791));
  xor_4  g21459(.A(new_n22357), .B(new_n22261), .Y(po0792));
  xnor_4 g21460(.A(new_n22793), .B(new_n4875), .Y(po0793));
  not_8  g21461(.A(new_n17903), .Y(new_n23810));
  nand_5 g21462(.A(new_n23810), .B(new_n17901), .Y(new_n23811));
  nand_5 g21463(.A(new_n17904), .B(new_n17853), .Y(new_n23812));
  nand_5 g21464(.A(new_n23812), .B(new_n17849), .Y(new_n23813));
  nand_5 g21465(.A(new_n23813), .B(new_n23811), .Y(new_n23814));
  not_8  g21466(.A(new_n23814), .Y(new_n23815));
  nor_5  g21467(.A(new_n23811), .B(new_n17851), .Y(new_n23816));
  nor_5  g21468(.A(new_n23816), .B(new_n23815), .Y(new_n23817));
  xor_4  g21469(.A(new_n23817), .B(new_n11660), .Y(po0794));
  xor_4  g21470(.A(new_n15762), .B(new_n15761), .Y(po0795));
  xnor_4 g21471(.A(new_n5008), .B(new_n4968), .Y(po0796));
  xnor_4 g21472(.A(new_n11063), .B(new_n11062), .Y(po0797));
  nand_5 g21473(.A(new_n20011), .B(new_n20009), .Y(new_n23822));
  nand_5 g21474(.A(new_n20024), .B(new_n23822), .Y(new_n23823));
  not_8  g21475(.A(new_n23823), .Y(new_n23824));
  nand_5 g21476(.A(new_n23704), .B(new_n23698), .Y(new_n23825));
  nand_5 g21477(.A(new_n23703), .B(new_n23699), .Y(new_n23826));
  nand_5 g21478(.A(new_n23826), .B(new_n23825), .Y(new_n23827));
  xor_4  g21479(.A(new_n23827), .B(new_n23824), .Y(po0798));
  not_8  g21480(.A(new_n12610), .Y(new_n23829));
  nand_5 g21481(.A(new_n12617), .B(new_n23829), .Y(new_n23830));
  nand_5 g21482(.A(new_n12615), .B(new_n12613), .Y(new_n23831));
  xnor_4 g21483(.A(new_n23831), .B(new_n23830), .Y(po0799));
  or_6   g21484(.A(new_n22139), .B(new_n22138), .Y(new_n23833));
  nand_5 g21485(.A(new_n22140), .B(new_n22137), .Y(new_n23834));
  nand_5 g21486(.A(new_n23834), .B(new_n23833), .Y(po0800));
  xor_4  g21487(.A(new_n11239), .B(new_n13128), .Y(po0801));
  xnor_4 g21488(.A(new_n12990), .B(new_n12957), .Y(po0802));
  nand_5 g21489(.A(new_n9502), .B(new_n9500), .Y(new_n23838));
  xor_4  g21490(.A(new_n23838), .B(new_n9471), .Y(po0803));
  xor_4  g21491(.A(new_n23465), .B(new_n23464), .Y(po0804));
  xor_4  g21492(.A(new_n12371), .B(new_n8917), .Y(po0805));
  xor_4  g21493(.A(new_n12680), .B(new_n7173), .Y(po0806));
  xor_4  g21494(.A(new_n9807), .B(new_n9805), .Y(po0807));
  xnor_4 g21495(.A(new_n23008), .B(new_n23007), .Y(po0808));
  xor_4  g21496(.A(new_n22361), .B(new_n10428), .Y(po0809));
  xnor_4 g21497(.A(new_n21936), .B(new_n21912), .Y(po0810));
  xor_4  g21498(.A(new_n14906), .B(new_n14868), .Y(po0811));
  xnor_4 g21499(.A(new_n21298), .B(new_n21297), .Y(po0812));
  xor_4  g21500(.A(new_n17629), .B(new_n8621), .Y(po0813));
  nand_5 g21501(.A(new_n21207), .B(new_n14817), .Y(new_n23850));
  nor_5  g21502(.A(new_n21206), .B(new_n21064), .Y(new_n23851));
  nand_5 g21503(.A(new_n23851), .B(new_n21197), .Y(new_n23852));
  nand_5 g21504(.A(new_n23852), .B(new_n23850), .Y(po0814));
  xor_4  g21505(.A(new_n6476), .B(new_n4628), .Y(po0815));
  nand_5 g21506(.A(new_n23816), .B(new_n11660), .Y(new_n23855));
  nand_5 g21507(.A(new_n23815), .B(new_n11661), .Y(new_n23856));
  nand_5 g21508(.A(new_n23856), .B(new_n23855), .Y(po0816));
  xor_4  g21509(.A(new_n8996), .B(new_n18643), .Y(po0817));
  xnor_4 g21510(.A(new_n13000), .B(new_n12937), .Y(po0818));
  xor_4  g21511(.A(new_n10941), .B(new_n10940), .Y(po0819));
  xor_4  g21512(.A(new_n22846), .B(new_n5698), .Y(po0820));
  xor_4  g21513(.A(new_n9139), .B(new_n9138), .Y(po0821));
  xor_4  g21514(.A(new_n22916), .B(new_n22913), .Y(po0822));
  nor_5  g21515(.A(new_n15550), .B(new_n15578), .Y(new_n23864));
  nor_5  g21516(.A(new_n15579), .B(new_n15577), .Y(new_n23865));
  nor_5  g21517(.A(new_n23865), .B(new_n23864), .Y(po0823));
  xor_4  g21518(.A(new_n18074), .B(new_n3339), .Y(po0824));
  nand_5 g21519(.A(new_n12163), .B(new_n12091), .Y(new_n23868));
  xor_4  g21520(.A(new_n23868), .B(new_n7251), .Y(po0825));
  xnor_4 g21521(.A(new_n19885), .B(new_n19884), .Y(po0826));
  nor_5  g21522(.A(new_n8254), .B(new_n8253), .Y(new_n23871));
  xor_4  g21523(.A(new_n23871), .B(new_n8255), .Y(po0827));
  xnor_4 g21524(.A(new_n11880), .B(new_n11879), .Y(po0828));
  xor_4  g21525(.A(new_n23667), .B(new_n23666), .Y(po0829));
  xor_4  g21526(.A(new_n19053), .B(new_n18977), .Y(po0830));
  not_8  g21527(.A(new_n17030), .Y(new_n23876));
  nand_5 g21528(.A(new_n17033), .B(new_n23876), .Y(new_n23877));
  xnor_4 g21529(.A(new_n23877), .B(new_n17022), .Y(po0831));
  xor_4  g21530(.A(new_n15091), .B(new_n15090), .Y(po0832));
  xor_4  g21531(.A(new_n15437), .B(new_n15436), .Y(po0833));
  xor_4  g21532(.A(new_n20607), .B(new_n20606), .Y(po0834));
  xnor_4 g21533(.A(new_n16494), .B(new_n13238), .Y(po0835));
  xor_4  g21534(.A(new_n5347), .B(new_n4186), .Y(po0836));
  xor_4  g21535(.A(new_n17295), .B(new_n13411), .Y(po0837));
  xor_4  g21536(.A(new_n9847), .B(new_n9846), .Y(po0838));
  xor_4  g21537(.A(new_n14127), .B(new_n14126), .Y(po0839));
  nand_5 g21538(.A(new_n23405), .B(new_n23399), .Y(new_n23887));
  xor_4  g21539(.A(new_n23887), .B(new_n22088), .Y(new_n23888));
  nand_5 g21540(.A(new_n23888), .B(new_n22748), .Y(new_n23889));
  nor_5  g21541(.A(new_n23889), .B(new_n23402), .Y(new_n23890));
  and_6  g21542(.A(new_n23888), .B(new_n23403), .Y(new_n23891));
  nand_5 g21543(.A(new_n23889), .B(new_n23402), .Y(new_n23892));
  nor_5  g21544(.A(new_n23892), .B(new_n23891), .Y(new_n23893));
  nor_5  g21545(.A(new_n23893), .B(new_n23890), .Y(po0840));
  nor_5  g21546(.A(new_n20374), .B(new_n20373), .Y(new_n23895));
  xor_4  g21547(.A(new_n23895), .B(new_n20375), .Y(po0841));
  nor_5  g21548(.A(new_n20337), .B(new_n20336), .Y(new_n23897));
  xor_4  g21549(.A(new_n23897), .B(new_n20266), .Y(po0842));
  nand_5 g21550(.A(new_n12963), .B(new_n12962), .Y(new_n23899));
  xnor_4 g21551(.A(new_n23899), .B(new_n12988), .Y(po0843));
  xnor_4 g21552(.A(new_n23496), .B(new_n5633), .Y(po0844));
  nand_5 g21553(.A(new_n23653), .B(new_n23644), .Y(new_n23902));
  nand_5 g21554(.A(new_n23654), .B(new_n23651), .Y(new_n23903));
  not_8  g21555(.A(new_n23903), .Y(new_n23904));
  nand_5 g21556(.A(new_n23904), .B(new_n23902), .Y(new_n23905));
  nand_5 g21557(.A(new_n23905), .B(new_n23654), .Y(new_n23906));
  nand_5 g21558(.A(new_n23906), .B(new_n23647), .Y(new_n23907));
  nor_5  g21559(.A(new_n23654), .B(new_n23644), .Y(new_n23908));
  nor_5  g21560(.A(new_n23908), .B(po0714), .Y(new_n23909));
  nand_5 g21561(.A(new_n23909), .B(new_n23907), .Y(po0845));
  xnor_4 g21562(.A(new_n9362), .B(new_n9361), .Y(po0846));
  xor_4  g21563(.A(new_n13799), .B(new_n2753), .Y(po0847));
  nor_5  g21564(.A(new_n23312), .B(new_n23294), .Y(new_n23913));
  nand_5 g21565(.A(new_n23913), .B(new_n23306), .Y(new_n23914));
  nand_5 g21566(.A(new_n23297), .B(new_n11090), .Y(new_n23915));
  not_8  g21567(.A(new_n23915), .Y(new_n23916));
  nor_5  g21568(.A(new_n23913), .B(new_n23306), .Y(new_n23917));
  nand_5 g21569(.A(new_n23917), .B(new_n23916), .Y(new_n23918));
  nand_5 g21570(.A(new_n23918), .B(new_n23914), .Y(po0848));
  nand_5 g21571(.A(new_n22889), .B(new_n22880), .Y(new_n23920));
  nand_5 g21572(.A(new_n22890), .B(new_n22879), .Y(new_n23921));
  nand_5 g21573(.A(new_n23921), .B(new_n23920), .Y(po0849));
  xor_4  g21574(.A(new_n23269), .B(new_n23045), .Y(po0850));
  xor_4  g21575(.A(new_n8610), .B(new_n6612), .Y(po0851));
  xor_4  g21576(.A(new_n13817), .B(new_n7990), .Y(po0852));
  xnor_4 g21577(.A(new_n14911), .B(new_n14862), .Y(po0853));
  nand_5 g21578(.A(new_n23582), .B(new_n23580), .Y(new_n23927));
  xor_4  g21579(.A(new_n23927), .B(new_n23577), .Y(po0854));
  xor_4  g21580(.A(new_n15296), .B(new_n15295), .Y(po0855));
  xor_4  g21581(.A(new_n12294), .B(new_n12292), .Y(po0856));
  nand_5 g21582(.A(new_n19164), .B(new_n19160), .Y(new_n23931));
  nand_5 g21583(.A(new_n19145), .B(new_n19138), .Y(new_n23932));
  xor_4  g21584(.A(new_n23932), .B(new_n19165), .Y(new_n23933));
  xor_4  g21585(.A(new_n23933), .B(new_n23931), .Y(po0857));
  xor_4  g21586(.A(new_n21738), .B(new_n18848), .Y(po0858));
  nor_5  g21587(.A(new_n22100), .B(new_n22138), .Y(new_n23936));
  nor_5  g21588(.A(new_n22754), .B(new_n22753), .Y(new_n23937));
  nor_5  g21589(.A(new_n23937), .B(new_n23936), .Y(po0859));
  not_8  g21590(.A(new_n22960), .Y(new_n23939));
  nand_5 g21591(.A(pi735), .B(new_n3208), .Y(new_n23940));
  not_8  g21592(.A(new_n23940), .Y(new_n23941));
  nor_5  g21593(.A(new_n20739), .B(new_n20737), .Y(new_n23942));
  nor_5  g21594(.A(new_n23942), .B(new_n23941), .Y(new_n23943));
  nor_5  g21595(.A(new_n20740), .B(new_n20735), .Y(new_n23944));
  nand_5 g21596(.A(new_n20741), .B(new_n20696), .Y(new_n23945));
  not_8  g21597(.A(new_n23945), .Y(new_n23946));
  nor_5  g21598(.A(new_n23946), .B(new_n23944), .Y(new_n23947));
  not_8  g21599(.A(new_n23947), .Y(new_n23948));
  or_6   g21600(.A(new_n23948), .B(new_n23943), .Y(new_n23949));
  nor_5  g21601(.A(new_n23949), .B(new_n22121), .Y(new_n23950));
  nand_5 g21602(.A(new_n23950), .B(new_n23939), .Y(new_n23951));
  not_8  g21603(.A(new_n22121), .Y(new_n23952));
  nand_5 g21604(.A(new_n23948), .B(new_n23943), .Y(new_n23953));
  nor_5  g21605(.A(new_n23953), .B(new_n23952), .Y(new_n23954));
  nand_5 g21606(.A(new_n23954), .B(new_n22957), .Y(new_n23955));
  nand_5 g21607(.A(new_n23955), .B(new_n23951), .Y(po0860));
  xor_4  g21608(.A(new_n12674), .B(new_n12673), .Y(po0861));
  xnor_4 g21609(.A(new_n11849), .B(new_n11847), .Y(po0862));
  xor_4  g21610(.A(new_n21932), .B(new_n21924), .Y(po0863));
  nand_5 g21611(.A(new_n22484), .B(new_n22483), .Y(new_n23960));
  xor_4  g21612(.A(new_n23960), .B(new_n22496), .Y(po0864));
  xor_4  g21613(.A(new_n9535), .B(new_n9524), .Y(po0865));
  xor_4  g21614(.A(new_n23020), .B(new_n23019), .Y(po0866));
  xor_4  g21615(.A(new_n3382), .B(new_n3381), .Y(po0867));
  xor_4  g21616(.A(new_n14789), .B(new_n10574), .Y(po0868));
  xor_4  g21617(.A(new_n19073), .B(new_n19072), .Y(po0869));
  xor_4  g21618(.A(new_n7925), .B(new_n7924), .Y(po0870));
  xor_4  g21619(.A(new_n22783), .B(new_n22769), .Y(po0871));
  xnor_4 g21620(.A(new_n12662), .B(new_n12661), .Y(po0872));
  xnor_4 g21621(.A(new_n8420), .B(new_n8415), .Y(po0873));
  xor_4  g21622(.A(new_n12174), .B(new_n12156), .Y(po0874));
  xor_4  g21623(.A(new_n9710), .B(new_n9709), .Y(po0875));
  xnor_4 g21624(.A(new_n8497), .B(new_n8481), .Y(po0876));
  nor_5  g21625(.A(new_n20208), .B(new_n4511), .Y(new_n23974));
  nor_5  g21626(.A(new_n23974), .B(new_n20207), .Y(new_n23975));
  or_6   g21627(.A(new_n23975), .B(new_n8218), .Y(new_n23976));
  not_8  g21628(.A(new_n23976), .Y(new_n23977));
  xor_4  g21629(.A(new_n23977), .B(new_n22175), .Y(new_n23978));
  xor_4  g21630(.A(new_n23975), .B(new_n8217), .Y(new_n23979));
  nand_5 g21631(.A(new_n23979), .B(new_n20631), .Y(new_n23980));
  nand_5 g21632(.A(new_n20210), .B(new_n20190), .Y(new_n23981));
  or_6   g21633(.A(new_n20236), .B(new_n20211), .Y(new_n23982));
  nand_5 g21634(.A(new_n23982), .B(new_n23981), .Y(new_n23983));
  xor_4  g21635(.A(new_n23979), .B(new_n20631), .Y(new_n23984));
  nand_5 g21636(.A(new_n23984), .B(new_n23983), .Y(new_n23985));
  nand_5 g21637(.A(new_n23985), .B(new_n23980), .Y(new_n23986));
  xnor_4 g21638(.A(new_n23986), .B(new_n23978), .Y(po0877));
  xor_4  g21639(.A(new_n19217), .B(new_n15187), .Y(po0878));
  nor_5  g21640(.A(new_n21540), .B(new_n15737), .Y(new_n23989));
  nor_5  g21641(.A(new_n21593), .B(new_n23989), .Y(new_n23990));
  nor_5  g21642(.A(new_n21595), .B(new_n21540), .Y(new_n23991));
  nor_5  g21643(.A(new_n23991), .B(new_n23990), .Y(po0879));
  xor_4  g21644(.A(new_n19195), .B(new_n14062), .Y(po0880));
  xor_4  g21645(.A(new_n14061), .B(new_n12257), .Y(po0881));
  xor_4  g21646(.A(new_n18494), .B(new_n7134), .Y(po0882));
  xor_4  g21647(.A(new_n21224), .B(new_n19860), .Y(new_n23996));
  not_8  g21648(.A(new_n23996), .Y(new_n23997));
  nand_5 g21649(.A(new_n21237), .B(new_n21227), .Y(new_n23998));
  nand_5 g21650(.A(new_n21238), .B(new_n19860), .Y(new_n23999));
  nand_5 g21651(.A(new_n23999), .B(new_n23998), .Y(new_n24000));
  xor_4  g21652(.A(new_n24000), .B(new_n23997), .Y(po0883));
  nand_5 g21653(.A(new_n13823), .B(new_n13822), .Y(new_n24002));
  xor_4  g21654(.A(new_n24002), .B(new_n13829), .Y(po0884));
  nor_5  g21655(.A(new_n17334), .B(new_n12402), .Y(po0885));
  xnor_4 g21656(.A(new_n23396), .B(new_n23395), .Y(po0886));
  nor_5  g21657(.A(new_n22322), .B(new_n21219), .Y(new_n24006));
  nand_5 g21658(.A(new_n22322), .B(new_n21219), .Y(new_n24007));
  nand_5 g21659(.A(new_n24007), .B(new_n21222), .Y(new_n24008));
  nor_5  g21660(.A(new_n24008), .B(new_n24006), .Y(new_n24009));
  not_8  g21661(.A(new_n21221), .Y(new_n24010));
  nand_5 g21662(.A(new_n22323), .B(new_n24010), .Y(new_n24011));
  nor_5  g21663(.A(new_n22322), .B(new_n21220), .Y(new_n24012));
  nand_5 g21664(.A(new_n21223), .B(new_n21220), .Y(new_n24013));
  nor_5  g21665(.A(new_n24013), .B(new_n22321), .Y(new_n24014));
  nor_5  g21666(.A(new_n24014), .B(new_n24012), .Y(new_n24015));
  nand_5 g21667(.A(new_n24015), .B(new_n24011), .Y(new_n24016));
  nor_5  g21668(.A(new_n24016), .B(new_n24009), .Y(po0887));
  nand_5 g21669(.A(new_n16753), .B(new_n12073), .Y(new_n24018));
  nand_5 g21670(.A(new_n23069), .B(new_n23066), .Y(new_n24019));
  nand_5 g21671(.A(new_n24019), .B(new_n24018), .Y(new_n24020));
  nand_5 g21672(.A(new_n24020), .B(new_n8986), .Y(new_n24021));
  xor_4  g21673(.A(new_n24020), .B(pi800), .Y(new_n24022));
  or_6   g21674(.A(new_n24022), .B(new_n16752), .Y(new_n24023));
  nand_5 g21675(.A(new_n24023), .B(new_n24021), .Y(new_n24024));
  nor_5  g21676(.A(new_n24024), .B(new_n23153), .Y(new_n24025));
  not_8  g21677(.A(new_n24025), .Y(new_n24026));
  xor_4  g21678(.A(new_n24024), .B(new_n23153), .Y(new_n24027));
  not_8  g21679(.A(new_n23065), .Y(new_n24028));
  nor_5  g21680(.A(new_n23070), .B(new_n24028), .Y(new_n24029));
  nor_5  g21681(.A(new_n23071), .B(new_n23059), .Y(new_n24030));
  nor_5  g21682(.A(new_n24030), .B(new_n24029), .Y(new_n24031));
  xor_4  g21683(.A(new_n24022), .B(new_n16752), .Y(new_n24032));
  or_6   g21684(.A(new_n24032), .B(new_n24031), .Y(new_n24033));
  not_8  g21685(.A(new_n23171), .Y(new_n24034));
  xor_4  g21686(.A(new_n24032), .B(new_n24031), .Y(new_n24035));
  nand_5 g21687(.A(new_n24035), .B(new_n24034), .Y(new_n24036));
  nand_5 g21688(.A(new_n24036), .B(new_n24033), .Y(new_n24037));
  nand_5 g21689(.A(new_n24037), .B(new_n23299), .Y(new_n24038));
  nor_5  g21690(.A(new_n24037), .B(new_n23299), .Y(new_n24039));
  not_8  g21691(.A(new_n24039), .Y(new_n24040));
  nand_5 g21692(.A(new_n24040), .B(new_n24038), .Y(new_n24041));
  or_6   g21693(.A(new_n24041), .B(new_n24027), .Y(new_n24042));
  nand_5 g21694(.A(new_n24042), .B(new_n23916), .Y(new_n24043));
  not_8  g21695(.A(new_n24043), .Y(new_n24044));
  nor_5  g21696(.A(new_n24027), .B(new_n23916), .Y(new_n24045));
  nand_5 g21697(.A(new_n24045), .B(new_n24038), .Y(new_n24046));
  nand_5 g21698(.A(new_n24046), .B(new_n24040), .Y(new_n24047));
  nor_5  g21699(.A(new_n24047), .B(new_n24044), .Y(new_n24048));
  xor_4  g21700(.A(new_n24048), .B(new_n24026), .Y(po0888));
  nand_5 g21701(.A(new_n23496), .B(new_n23490), .Y(new_n24050));
  not_8  g21702(.A(new_n23484), .Y(new_n24051));
  nand_5 g21703(.A(new_n24051), .B(new_n18759), .Y(new_n24052));
  nor_5  g21704(.A(new_n23483), .B(new_n18759), .Y(new_n24053));
  nor_5  g21705(.A(new_n24053), .B(new_n22245), .Y(new_n24054));
  nand_5 g21706(.A(new_n24054), .B(new_n24052), .Y(new_n24055));
  nand_5 g21707(.A(new_n23486), .B(new_n18760), .Y(new_n24056));
  nor_5  g21708(.A(new_n23482), .B(new_n18760), .Y(new_n24057));
  nor_5  g21709(.A(new_n24057), .B(new_n23487), .Y(new_n24058));
  nand_5 g21710(.A(new_n24058), .B(new_n24056), .Y(new_n24059));
  nand_5 g21711(.A(new_n24059), .B(new_n24055), .Y(new_n24060));
  or_6   g21712(.A(new_n23486), .B(new_n24051), .Y(new_n24061));
  not_8  g21713(.A(new_n23493), .Y(new_n24062));
  nand_5 g21714(.A(new_n24062), .B(new_n23488), .Y(new_n24063));
  nor_5  g21715(.A(new_n24063), .B(new_n24061), .Y(new_n24064));
  nor_5  g21716(.A(new_n24064), .B(new_n5753), .Y(new_n24065));
  nand_5 g21717(.A(new_n24065), .B(new_n24060), .Y(new_n24066));
  nand_5 g21718(.A(new_n24066), .B(new_n24050), .Y(po0889));
  nand_5 g21719(.A(new_n23740), .B(new_n23739), .Y(new_n24068));
  xor_4  g21720(.A(new_n24068), .B(new_n23743), .Y(po0890));
  not_8  g21721(.A(new_n23158), .Y(new_n24070));
  nand_5 g21722(.A(new_n24070), .B(new_n23155), .Y(new_n24071));
  nand_5 g21723(.A(new_n23160), .B(new_n23150), .Y(new_n24072));
  nand_5 g21724(.A(new_n24072), .B(new_n24071), .Y(new_n24073));
  nand_5 g21725(.A(new_n23153), .B(new_n6386), .Y(new_n24074));
  or_6   g21726(.A(new_n23154), .B(new_n12083), .Y(new_n24075));
  nand_5 g21727(.A(new_n24075), .B(new_n24074), .Y(new_n24076));
  xnor_4 g21728(.A(new_n24076), .B(new_n24073), .Y(po0891));
  xnor_4 g21729(.A(new_n17836), .B(new_n17835), .Y(po0892));
  xor_4  g21730(.A(new_n15406), .B(new_n15380), .Y(po0893));
  xnor_4 g21731(.A(new_n16852), .B(new_n8255), .Y(po0894));
  xnor_4 g21732(.A(new_n12709), .B(new_n12708), .Y(po0895));
  xor_4  g21733(.A(new_n21256), .B(new_n11416), .Y(po0896));
  xnor_4 g21734(.A(new_n21340), .B(new_n21336), .Y(po0897));
  xor_4  g21735(.A(new_n19322), .B(new_n19321), .Y(po0898));
  xor_4  g21736(.A(new_n3866), .B(new_n3865), .Y(po0899));
  xor_4  g21737(.A(new_n6909), .B(new_n6899), .Y(po0900));
  nand_5 g21738(.A(new_n8484), .B(new_n8483), .Y(new_n24087));
  xnor_4 g21739(.A(new_n24087), .B(new_n8495), .Y(po0901));
  xnor_4 g21740(.A(new_n17596), .B(new_n17595), .Y(po0902));
  xnor_4 g21741(.A(new_n10381), .B(new_n10380), .Y(po0903));
  nand_5 g21742(.A(new_n20845), .B(new_n18033), .Y(new_n24091));
  not_8  g21743(.A(new_n20846), .Y(new_n24092));
  nand_5 g21744(.A(new_n24092), .B(new_n20844), .Y(new_n24093));
  nand_5 g21745(.A(new_n24093), .B(new_n24091), .Y(po0904));
  xor_4  g21746(.A(new_n17604), .B(new_n17568), .Y(po0905));
  xor_4  g21747(.A(new_n21721), .B(new_n17650), .Y(po0906));
  xor_4  g21748(.A(new_n6612), .B(new_n6610), .Y(po0907));
  xor_4  g21749(.A(new_n19430), .B(new_n19397), .Y(po0908));
  xor_4  g21750(.A(new_n20347), .B(new_n9481), .Y(po0909));
  xnor_4 g21751(.A(new_n13810), .B(new_n13808), .Y(po0910));
  xor_4  g21752(.A(new_n22532), .B(new_n22524), .Y(po0911));
  xnor_4 g21753(.A(new_n24041), .B(new_n24027), .Y(po0912));
  xnor_4 g21754(.A(new_n8435), .B(new_n8434), .Y(po0913));
  xor_4  g21755(.A(new_n21246), .B(new_n14204), .Y(po0914));
  xor_4  g21756(.A(new_n12190), .B(new_n12135), .Y(po0916));
  xnor_4 g21757(.A(new_n17838), .B(new_n17824), .Y(po0917));
  xor_4  g21758(.A(new_n14381), .B(new_n14322), .Y(new_n24107));
  xor_4  g21759(.A(new_n24107), .B(new_n14451), .Y(po0918));
  xor_4  g21760(.A(new_n20232), .B(new_n20222), .Y(po0919));
  nor_5  g21761(.A(new_n15097), .B(new_n22974), .Y(new_n24110));
  xor_4  g21762(.A(new_n15098), .B(new_n11290), .Y(new_n24111));
  not_8  g21763(.A(new_n24111), .Y(new_n24112));
  nand_5 g21764(.A(new_n20908), .B(new_n20891), .Y(new_n24113));
  nand_5 g21765(.A(new_n24113), .B(new_n20890), .Y(new_n24114));
  nor_5  g21766(.A(new_n24114), .B(new_n24112), .Y(new_n24115));
  nor_5  g21767(.A(new_n24115), .B(new_n24110), .Y(po0920));
  xnor_4 g21768(.A(new_n4676), .B(new_n4674), .Y(po0921));
  xor_4  g21769(.A(new_n13086), .B(new_n13083), .Y(po0922));
  xor_4  g21770(.A(new_n22609), .B(new_n3767), .Y(po0923));
  xor_4  g21771(.A(new_n15898), .B(new_n15896), .Y(po0924));
  xor_4  g21772(.A(new_n10930), .B(new_n9351), .Y(po0925));
  nand_5 g21773(.A(new_n6025), .B(new_n6027), .Y(new_n24122));
  xor_4  g21774(.A(new_n24122), .B(new_n5779), .Y(po0926));
  nand_5 g21775(.A(new_n10419), .B(new_n10399), .Y(new_n24124));
  nor_5  g21776(.A(new_n10416), .B(new_n10396), .Y(new_n24125));
  nand_5 g21777(.A(new_n22038), .B(new_n10421), .Y(new_n24126));
  nand_5 g21778(.A(new_n24126), .B(new_n10398), .Y(new_n24127));
  nand_5 g21779(.A(new_n10423), .B(new_n10395), .Y(new_n24128));
  nand_5 g21780(.A(new_n24128), .B(new_n24127), .Y(new_n24129));
  nor_5  g21781(.A(new_n24129), .B(new_n24125), .Y(new_n24130));
  nand_5 g21782(.A(new_n24130), .B(new_n24124), .Y(po0927));
  xnor_4 g21783(.A(new_n19505), .B(new_n19479), .Y(po0928));
  xor_4  g21784(.A(new_n22047), .B(new_n21234), .Y(po0929));
  xnor_4 g21785(.A(new_n22804), .B(new_n22803), .Y(po0930));
  xnor_4 g21786(.A(new_n7673), .B(new_n7639), .Y(po0931));
  xnor_4 g21787(.A(new_n22774), .B(new_n4882), .Y(po0932));
  nor_5  g21788(.A(new_n2529), .B(new_n2489), .Y(new_n24137));
  xor_4  g21789(.A(new_n24137), .B(new_n2523), .Y(po0933));
  xor_4  g21790(.A(new_n6927), .B(new_n6871), .Y(po0934));
  xor_4  g21791(.A(new_n14449), .B(new_n14388), .Y(po0935));
  xor_4  g21792(.A(new_n22726), .B(new_n22725), .Y(po0936));
  xor_4  g21793(.A(new_n10675), .B(new_n10671), .Y(po0937));
  xnor_4 g21794(.A(new_n6192), .B(new_n6191), .Y(po0938));
  xor_4  g21795(.A(new_n7937), .B(new_n7936), .Y(po0939));
  xnor_4 g21796(.A(new_n16977), .B(new_n16969), .Y(po0940));
  xor_4  g21797(.A(new_n3100), .B(new_n3056), .Y(po0941));
  xnor_4 g21798(.A(new_n22317), .B(new_n22316), .Y(po0942));
  xor_4  g21799(.A(new_n5069), .B(new_n5068), .Y(po0943));
  xor_4  g21800(.A(new_n8289), .B(new_n8288), .Y(po0944));
  nand_5 g21801(.A(new_n22222), .B(new_n18403), .Y(new_n24150));
  nor_5  g21802(.A(new_n22221), .B(new_n18408), .Y(new_n24151));
  nor_5  g21803(.A(new_n24151), .B(new_n22230), .Y(new_n24152));
  nand_5 g21804(.A(new_n24152), .B(new_n24150), .Y(po0945));
  nand_5 g21805(.A(new_n16457), .B(new_n16458), .Y(new_n24154));
  xor_4  g21806(.A(new_n24154), .B(new_n16468), .Y(po0946));
  xor_4  g21807(.A(new_n8417), .B(new_n3642), .Y(po0947));
  xnor_4 g21808(.A(new_n19433), .B(new_n19432), .Y(po0948));
  xor_4  g21809(.A(new_n13601), .B(new_n13576), .Y(po0949));
  xnor_4 g21810(.A(new_n15395), .B(new_n13808), .Y(po0950));
  xnor_4 g21811(.A(new_n20840), .B(new_n20839), .Y(po0951));
  xnor_4 g21812(.A(new_n17263), .B(new_n17240), .Y(po0952));
  xnor_4 g21813(.A(new_n4635), .B(new_n4603), .Y(po0953));
  xnor_4 g21814(.A(new_n13478), .B(new_n13476), .Y(po0954));
  xor_4  g21815(.A(new_n9819), .B(new_n9817), .Y(po0955));
  xor_4  g21816(.A(new_n13370), .B(new_n13368), .Y(new_n24165));
  xor_4  g21817(.A(new_n24165), .B(new_n13333), .Y(po0956));
  xor_4  g21818(.A(new_n23255), .B(new_n19357), .Y(po0957));
  xor_4  g21819(.A(new_n22612), .B(new_n22611), .Y(new_n24168));
  xor_4  g21820(.A(new_n24168), .B(new_n16990), .Y(po0958));
  xor_4  g21821(.A(new_n20442), .B(new_n20441), .Y(po0959));
  xor_4  g21822(.A(new_n11616), .B(new_n11075), .Y(po0960));
  xnor_4 g21823(.A(new_n19674), .B(new_n19671), .Y(po0961));
  xor_4  g21824(.A(new_n18889), .B(new_n18888), .Y(po0962));
  nor_5  g21825(.A(new_n15515), .B(new_n15514), .Y(new_n24174));
  xor_4  g21826(.A(new_n24174), .B(new_n15516), .Y(po0963));
  xnor_4 g21827(.A(new_n10625), .B(new_n10624), .Y(po0964));
  xor_4  g21828(.A(new_n11250), .B(new_n11249), .Y(po0965));
  nand_5 g21829(.A(new_n19866), .B(new_n19837), .Y(new_n24178));
  nand_5 g21830(.A(new_n19867), .B(new_n19863), .Y(new_n24179));
  nand_5 g21831(.A(new_n24179), .B(new_n24178), .Y(po0966));
  xor_4  g21832(.A(new_n11837), .B(new_n11799), .Y(po0967));
  xnor_4 g21833(.A(new_n2805), .B(new_n2804), .Y(po0968));
  nand_5 g21834(.A(new_n22428), .B(new_n22426), .Y(new_n24183));
  xnor_4 g21835(.A(new_n24183), .B(new_n3389), .Y(po0969));
  not_8  g21836(.A(new_n22455), .Y(new_n24185));
  nand_5 g21837(.A(new_n24185), .B(new_n22445), .Y(new_n24186));
  nor_5  g21838(.A(new_n22446), .B(new_n22388), .Y(new_n24187));
  nand_5 g21839(.A(new_n24187), .B(new_n23722), .Y(new_n24188));
  nor_5  g21840(.A(new_n22440), .B(new_n22442), .Y(new_n24189));
  nor_5  g21841(.A(new_n24189), .B(new_n22449), .Y(new_n24190));
  nor_5  g21842(.A(new_n24190), .B(new_n22454), .Y(new_n24191));
  nand_5 g21843(.A(new_n24191), .B(new_n24188), .Y(new_n24192));
  nand_5 g21844(.A(new_n24192), .B(new_n24186), .Y(po0970));
  xor_4  g21845(.A(new_n14420), .B(new_n13540), .Y(po0971));
  xor_4  g21846(.A(new_n13241), .B(new_n5059), .Y(po0972));
  xnor_4 g21847(.A(new_n19428), .B(new_n19427), .Y(po0973));
  xnor_4 g21848(.A(new_n22728), .B(new_n22703), .Y(po0974));
  xnor_4 g21849(.A(new_n12313), .B(new_n6488), .Y(po0975));
  xnor_4 g21850(.A(new_n21570), .B(new_n21549), .Y(po0976));
  xor_4  g21851(.A(new_n7134), .B(new_n4597), .Y(po0977));
  xor_4  g21852(.A(new_n8502), .B(new_n13084), .Y(po0978));
  nor_5  g21853(.A(new_n7505), .B(new_n7392), .Y(new_n24202));
  nor_5  g21854(.A(new_n24202), .B(new_n19170), .Y(new_n24203));
  nor_5  g21855(.A(new_n24202), .B(new_n7511), .Y(new_n24204));
  nor_5  g21856(.A(new_n24204), .B(new_n24203), .Y(po0979));
  xnor_4 g21857(.A(new_n23695), .B(new_n23694), .Y(po0980));
  xnor_4 g21858(.A(new_n13687), .B(new_n13677), .Y(po0981));
  xor_4  g21859(.A(new_n22078), .B(new_n16441), .Y(po0982));
  xor_4  g21860(.A(new_n23002), .B(new_n17805), .Y(po0983));
  xnor_4 g21861(.A(new_n5731), .B(new_n5730), .Y(po0984));
  xor_4  g21862(.A(new_n15250), .B(new_n5772), .Y(po0985));
  xnor_4 g21863(.A(new_n16868), .B(new_n16828), .Y(po0986));
  xor_4  g21864(.A(new_n14439), .B(new_n14407), .Y(po0987));
  xnor_4 g21865(.A(new_n8424), .B(new_n8408), .Y(po0988));
  xor_4  g21866(.A(new_n20234), .B(new_n20217), .Y(po0989));
  xnor_4 g21867(.A(new_n14022), .B(new_n13983), .Y(po0990));
  xor_4  g21868(.A(new_n22284), .B(new_n22263), .Y(po0991));
  nor_5  g21869(.A(new_n21686), .B(new_n21667), .Y(new_n24218));
  and_6  g21870(.A(new_n24218), .B(new_n21682), .Y(new_n24219));
  nand_5 g21871(.A(new_n21812), .B(new_n21674), .Y(new_n24220));
  xor_4  g21872(.A(new_n24218), .B(new_n21682), .Y(new_n24221));
  nand_5 g21873(.A(new_n24221), .B(new_n21672), .Y(new_n24222));
  nand_5 g21874(.A(new_n24222), .B(new_n24220), .Y(new_n24223));
  nor_5  g21875(.A(new_n24223), .B(new_n24219), .Y(po0992));
  xor_4  g21876(.A(new_n15610), .B(new_n15607), .Y(po0993));
  xnor_4 g21877(.A(new_n23459), .B(new_n23458), .Y(po0994));
  xnor_4 g21878(.A(new_n19037), .B(new_n19018), .Y(po0995));
  xor_4  g21879(.A(new_n14437), .B(new_n14413), .Y(po0996));
  nand_5 g21880(.A(new_n4939), .B(new_n4870), .Y(new_n24229));
  not_8  g21881(.A(new_n4939), .Y(new_n24230));
  nand_5 g21882(.A(new_n24230), .B(new_n4871), .Y(new_n24231));
  nand_5 g21883(.A(new_n24231), .B(new_n24229), .Y(new_n24232));
  nor_5  g21884(.A(new_n4940), .B(new_n4752), .Y(new_n24233));
  nor_5  g21885(.A(new_n5019), .B(new_n4942), .Y(new_n24234));
  or_6   g21886(.A(new_n24234), .B(new_n24233), .Y(new_n24235));
  not_8  g21887(.A(new_n24235), .Y(new_n24236));
  or_6   g21888(.A(new_n24236), .B(new_n24232), .Y(new_n24237));
  and_6  g21889(.A(new_n24237), .B(new_n24229), .Y(po0997));
  xnor_4 g21890(.A(new_n15821), .B(new_n15820), .Y(po0998));
  nor_5  g21891(.A(new_n23363), .B(new_n23359), .Y(new_n24240));
  not_8  g21892(.A(new_n23361), .Y(new_n24241));
  nand_5 g21893(.A(new_n23348), .B(new_n24241), .Y(new_n24242));
  nand_5 g21894(.A(new_n24242), .B(new_n23360), .Y(new_n24243));
  nor_5  g21895(.A(new_n24243), .B(new_n24240), .Y(po0999));
  xnor_4 g21896(.A(new_n22718), .B(new_n22715), .Y(po1000));
  xor_4  g21897(.A(new_n22789), .B(new_n4877), .Y(po1001));
  xor_4  g21898(.A(new_n7932), .B(new_n7931), .Y(po1002));
  xor_4  g21899(.A(new_n16031), .B(new_n11458), .Y(po1003));
  nor_5  g21900(.A(new_n13044), .B(new_n13035), .Y(new_n24249));
  nand_5 g21901(.A(new_n24249), .B(new_n13042), .Y(new_n24250));
  nand_5 g21902(.A(new_n13043), .B(new_n13035), .Y(new_n24251));
  nand_5 g21903(.A(new_n24251), .B(new_n24250), .Y(po1004));
  nor_5  g21904(.A(new_n13305), .B(new_n13306), .Y(new_n24253));
  nor_5  g21905(.A(new_n13307), .B(new_n7222), .Y(new_n24254));
  nor_5  g21906(.A(new_n24254), .B(new_n24253), .Y(new_n24255));
  nand_5 g21907(.A(pi785), .B(new_n16216), .Y(new_n24256));
  nand_5 g21908(.A(new_n17845), .B(new_n17841), .Y(new_n24257));
  nand_5 g21909(.A(new_n24257), .B(new_n24256), .Y(new_n24258));
  and_6  g21910(.A(new_n24258), .B(new_n13370), .Y(new_n24259));
  or_6   g21911(.A(new_n17846), .B(new_n13336), .Y(new_n24260));
  nand_5 g21912(.A(new_n17847), .B(new_n17840), .Y(new_n24261));
  nand_5 g21913(.A(new_n24261), .B(new_n24260), .Y(new_n24262));
  and_6  g21914(.A(new_n24262), .B(new_n24259), .Y(new_n24263));
  or_6   g21915(.A(new_n24258), .B(new_n13370), .Y(new_n24264));
  nor_5  g21916(.A(new_n24264), .B(new_n24262), .Y(new_n24265));
  nor_5  g21917(.A(new_n24265), .B(new_n24263), .Y(new_n24266));
  nor_5  g21918(.A(new_n24266), .B(new_n24255), .Y(po1005));
  xor_4  g21919(.A(new_n7169), .B(new_n7168), .Y(po1006));
  xor_4  g21920(.A(new_n6135), .B(new_n6442), .Y(new_n24269));
  xor_4  g21921(.A(new_n24269), .B(new_n2754), .Y(po1007));
  xor_4  g21922(.A(new_n21189), .B(new_n21144), .Y(po1008));
  xnor_4 g21923(.A(new_n22643), .B(new_n20872), .Y(po1009));
  xor_4  g21924(.A(new_n3874), .B(new_n12039), .Y(po1010));
  nand_5 g21925(.A(new_n20832), .B(new_n20833), .Y(new_n24274));
  xor_4  g21926(.A(new_n24274), .B(new_n20835), .Y(po1011));
  xnor_4 g21927(.A(new_n3409), .B(new_n3408), .Y(po1012));
  xor_4  g21928(.A(new_n10182), .B(new_n10164), .Y(po1013));
  xor_4  g21929(.A(new_n22082), .B(new_n21614), .Y(po1014));
  nand_5 g21930(.A(new_n7665), .B(new_n7650), .Y(new_n24279));
  xnor_4 g21931(.A(new_n24279), .B(new_n7663), .Y(po1015));
  nor_5  g21932(.A(new_n11893), .B(new_n11888), .Y(new_n24281));
  xor_4  g21933(.A(new_n24281), .B(new_n11871), .Y(po1016));
  xor_4  g21934(.A(new_n17265), .B(new_n17236), .Y(po1017));
  xnor_4 g21935(.A(new_n18875), .B(new_n18872), .Y(po1018));
  xnor_4 g21936(.A(new_n21565), .B(new_n21564), .Y(po1019));
  xnor_4 g21937(.A(new_n22282), .B(new_n22266), .Y(po1020));
  xor_4  g21938(.A(new_n17326), .B(new_n12399), .Y(po1021));
  xor_4  g21939(.A(new_n22619), .B(new_n17009), .Y(po1022));
  xnor_4 g21940(.A(new_n13721), .B(new_n13709), .Y(po1023));
  xor_4  g21941(.A(new_n6614), .B(new_n6613), .Y(po1024));
  nand_5 g21942(.A(new_n17940), .B(new_n17939), .Y(new_n24291));
  xnor_4 g21943(.A(new_n24291), .B(new_n17956), .Y(po1025));
  xor_4  g21944(.A(new_n5444), .B(new_n5441), .Y(po1026));
  xnor_4 g21945(.A(new_n22807), .B(new_n22806), .Y(po1027));
  xor_4  g21946(.A(new_n19750), .B(new_n19748), .Y(po1028));
  xor_4  g21947(.A(new_n18464), .B(new_n6893), .Y(po1029));
  xnor_4 g21948(.A(new_n5014), .B(new_n4952), .Y(po1030));
  xor_4  g21949(.A(new_n4039), .B(new_n4038), .Y(po1031));
  xnor_4 g21950(.A(new_n17083), .B(new_n17072), .Y(po1032));
  xnor_4 g21951(.A(new_n14964), .B(new_n14963), .Y(po1033));
  nand_5 g21952(.A(new_n8227), .B(new_n8226), .Y(new_n24301));
  xor_4  g21953(.A(new_n24301), .B(new_n8272), .Y(po1034));
  xnor_4 g21954(.A(new_n20625), .B(new_n20576), .Y(po1035));
  xnor_4 g21955(.A(new_n11332), .B(new_n11329), .Y(po1036));
  nor_5  g21956(.A(new_n6877), .B(new_n6876), .Y(new_n24305));
  xor_4  g21957(.A(new_n24305), .B(new_n6925), .Y(po1037));
  xor_4  g21958(.A(new_n18903), .B(new_n18847), .Y(po1038));
  xor_4  g21959(.A(new_n19213), .B(new_n19192), .Y(po1039));
  xor_4  g21960(.A(new_n14223), .B(new_n9031), .Y(new_n24309));
  nand_5 g21961(.A(new_n14234), .B(new_n14231), .Y(new_n24310));
  xor_4  g21962(.A(new_n24310), .B(new_n24309), .Y(po1040));
  xnor_4 g21963(.A(new_n15404), .B(new_n15402), .Y(po1041));
  xor_4  g21964(.A(new_n16312), .B(new_n16283), .Y(po1042));
  nor_5  g21965(.A(new_n24044), .B(new_n24026), .Y(new_n24314));
  nor_5  g21966(.A(new_n24047), .B(new_n24025), .Y(new_n24315));
  nor_5  g21967(.A(new_n24315), .B(new_n24314), .Y(po1043));
  xor_4  g21968(.A(new_n21717), .B(new_n17645), .Y(po1044));
  nor_5  g21969(.A(new_n23135), .B(new_n23133), .Y(new_n24318));
  xor_4  g21970(.A(new_n24318), .B(new_n17937), .Y(po1045));
  xor_4  g21971(.A(new_n20342), .B(new_n20341), .Y(po1046));
  xor_4  g21972(.A(new_n20799), .B(new_n6021), .Y(po1047));
  xnor_4 g21973(.A(new_n22657), .B(new_n22656), .Y(po1048));
  nor_5  g21974(.A(new_n6708), .B(new_n6709), .Y(new_n24323));
  xor_4  g21975(.A(new_n24323), .B(new_n3367), .Y(po1049));
  xnor_4 g21976(.A(new_n3689), .B(new_n3688), .Y(po1050));
  nand_5 g21977(.A(new_n20949), .B(new_n20936), .Y(new_n24326));
  xnor_4 g21978(.A(new_n24326), .B(new_n20948), .Y(po1051));
  xor_4  g21979(.A(new_n3098), .B(new_n3060), .Y(po1052));
  nand_5 g21980(.A(new_n23511), .B(new_n23507), .Y(new_n24329));
  xnor_4 g21981(.A(new_n24329), .B(new_n23505), .Y(po1053));
  xor_4  g21982(.A(new_n19049), .B(new_n4945), .Y(po1054));
  xor_4  g21983(.A(new_n21372), .B(new_n21371), .Y(po1055));
  xor_4  g21984(.A(new_n16857), .B(new_n8232), .Y(po1056));
  xor_4  g21985(.A(new_n19990), .B(new_n19988), .Y(po1057));
  or_6   g21986(.A(new_n7691), .B(new_n7688), .Y(new_n24335));
  and_6  g21987(.A(new_n24335), .B(new_n7696), .Y(new_n24336));
  nor_5  g21988(.A(new_n24336), .B(new_n7692), .Y(po1058));
  xnor_4 g21989(.A(new_n11058), .B(new_n11042), .Y(po1059));
  xnor_4 g21990(.A(new_n13135), .B(new_n11244), .Y(po1060));
  xnor_4 g21991(.A(new_n12172), .B(new_n12159), .Y(po1061));
  xnor_4 g21992(.A(new_n3093), .B(new_n3092), .Y(po1062));
  xor_4  g21993(.A(new_n10023), .B(new_n10022), .Y(po1063));
  xor_4  g21994(.A(new_n17606), .B(new_n17564), .Y(po1064));
  xor_4  g21995(.A(new_n4527), .B(new_n4525), .Y(po1065));
  xor_4  g21996(.A(new_n22003), .B(new_n6939), .Y(po1066));
  xor_4  g21997(.A(new_n16848), .B(new_n16847), .Y(po1067));
  xor_4  g21998(.A(new_n8954), .B(new_n8953), .Y(po1068));
  xnor_4 g21999(.A(new_n12625), .B(new_n12624), .Y(po1069));
  xor_4  g22000(.A(new_n23903), .B(new_n23902), .Y(new_n24349));
  xor_4  g22001(.A(new_n24349), .B(new_n4868), .Y(po1070));
  xor_4  g22002(.A(new_n23332), .B(new_n23331), .Y(po1071));
  xor_4  g22003(.A(new_n17332), .B(new_n17330), .Y(po1072));
  xor_4  g22004(.A(new_n15521), .B(new_n10023), .Y(po1073));
  xor_4  g22005(.A(new_n21456), .B(new_n21426), .Y(po1074));
  xor_4  g22006(.A(new_n5744), .B(new_n23479), .Y(po1075));
  xor_4  g22007(.A(new_n15252), .B(new_n15243), .Y(po1076));
  xor_4  g22008(.A(new_n5739), .B(new_n5681), .Y(po1077));
  nor_5  g22009(.A(new_n17718), .B(new_n14389), .Y(new_n24358));
  nor_5  g22010(.A(new_n19084), .B(new_n19083), .Y(new_n24359));
  nor_5  g22011(.A(new_n24359), .B(new_n24358), .Y(new_n24360));
  nor_5  g22012(.A(new_n24360), .B(new_n17714), .Y(new_n24361));
  xor_4  g22013(.A(new_n24360), .B(new_n17714), .Y(new_n24362));
  not_8  g22014(.A(new_n24362), .Y(new_n24363));
  nor_5  g22015(.A(new_n24363), .B(new_n14384), .Y(new_n24364));
  or_6   g22016(.A(new_n24364), .B(new_n24361), .Y(new_n24365));
  or_6   g22017(.A(new_n24365), .B(new_n17733), .Y(new_n24366));
  nand_5 g22018(.A(new_n24365), .B(new_n17733), .Y(new_n24367));
  nand_5 g22019(.A(new_n24367), .B(new_n24366), .Y(new_n24368));
  xor_4  g22020(.A(new_n24368), .B(new_n14322), .Y(po1078));
  xor_4  g22021(.A(new_n8430), .B(new_n8398), .Y(po1079));
  xor_4  g22022(.A(new_n21636), .B(new_n16390), .Y(po1080));
  xor_4  g22023(.A(new_n22623), .B(new_n17007), .Y(po1081));
  xnor_4 g22024(.A(new_n20718), .B(new_n20717), .Y(po1082));
  xnor_4 g22025(.A(new_n7968), .B(new_n7912), .Y(po1083));
  xnor_4 g22026(.A(new_n11475), .B(new_n4662), .Y(po1084));
  xor_4  g22027(.A(new_n17590), .B(new_n17589), .Y(po1085));
  xor_4  g22028(.A(new_n15975), .B(new_n15957), .Y(po1086));
  xor_4  g22029(.A(new_n13120), .B(new_n6081), .Y(po1087));
  xnor_4 g22030(.A(new_n8958), .B(new_n8956), .Y(po1088));
  xnor_4 g22031(.A(new_n10944), .B(new_n10943), .Y(po1089));
  xor_4  g22032(.A(new_n13657), .B(new_n3480), .Y(po1090));
  xor_4  g22033(.A(new_n22422), .B(new_n3336), .Y(po1091));
  not_8  g22034(.A(new_n17707), .Y(new_n24383));
  nand_5 g22035(.A(new_n18170), .B(new_n24383), .Y(new_n24384));
  not_8  g22036(.A(new_n24384), .Y(new_n24385));
  nand_5 g22037(.A(new_n24385), .B(new_n10211), .Y(new_n24386));
  nand_5 g22038(.A(new_n17736), .B(new_n17711), .Y(new_n24387));
  nand_5 g22039(.A(new_n17737), .B(new_n10219), .Y(new_n24388));
  nand_5 g22040(.A(new_n24388), .B(new_n24387), .Y(new_n24389));
  xor_4  g22041(.A(new_n24384), .B(new_n10210), .Y(new_n24390));
  nand_5 g22042(.A(new_n24390), .B(new_n24389), .Y(new_n24391));
  nand_5 g22043(.A(new_n24391), .B(new_n24386), .Y(po1092));
  xor_4  g22044(.A(new_n17285), .B(new_n17283), .Y(po1093));
  xor_4  g22045(.A(new_n11267), .B(new_n8808), .Y(po1094));
  xnor_4 g22046(.A(new_n19586), .B(new_n19585), .Y(po1095));
  xor_4  g22047(.A(new_n17436), .B(new_n17350), .Y(po1096));
  xnor_4 g22048(.A(new_n16744), .B(new_n16709), .Y(po1097));
  xor_4  g22049(.A(new_n22919), .B(new_n22910), .Y(po1098));
  xor_4  g22050(.A(new_n19773), .B(new_n19772), .Y(po1099));
  xor_4  g22051(.A(new_n22021), .B(new_n22009), .Y(new_n24400));
  xor_4  g22052(.A(new_n24400), .B(new_n17352), .Y(po1100));
  nor_5  g22053(.A(new_n24385), .B(new_n14321), .Y(new_n24402));
  xor_4  g22054(.A(new_n24384), .B(new_n14320), .Y(new_n24403));
  not_8  g22055(.A(new_n24403), .Y(new_n24404));
  nand_5 g22056(.A(new_n17711), .B(new_n14456), .Y(new_n24405));
  xor_4  g22057(.A(new_n17711), .B(new_n14456), .Y(new_n24406));
  nand_5 g22058(.A(new_n24367), .B(new_n14322), .Y(new_n24407));
  nand_5 g22059(.A(new_n24407), .B(new_n24366), .Y(new_n24408));
  nand_5 g22060(.A(new_n24408), .B(new_n24406), .Y(new_n24409));
  nand_5 g22061(.A(new_n24409), .B(new_n24405), .Y(new_n24410));
  nor_5  g22062(.A(new_n24410), .B(new_n24404), .Y(new_n24411));
  nor_5  g22063(.A(new_n24411), .B(new_n24402), .Y(po1101));
  xor_4  g22064(.A(new_n15613), .B(new_n15612), .Y(po1102));
  xnor_4 g22065(.A(new_n8279), .B(new_n8278), .Y(po1103));
  xnor_4 g22066(.A(new_n15572), .B(new_n13077), .Y(po1104));
  xnor_4 g22067(.A(new_n4497), .B(new_n4496), .Y(po1105));
  nand_5 g22068(.A(new_n12274), .B(new_n12270), .Y(new_n24417));
  xor_4  g22069(.A(new_n24417), .B(new_n12273), .Y(po1106));
  nand_5 g22070(.A(new_n12690), .B(new_n12689), .Y(new_n24419));
  xnor_4 g22071(.A(new_n24419), .B(new_n12701), .Y(po1107));
  nand_5 g22072(.A(new_n14020), .B(new_n14019), .Y(new_n24421));
  xor_4  g22073(.A(new_n24421), .B(new_n12926), .Y(po1108));
  xor_4  g22074(.A(new_n22965), .B(new_n22964), .Y(po1109));
  nand_5 g22075(.A(new_n22734), .B(new_n22732), .Y(new_n24424));
  xor_4  g22076(.A(new_n24424), .B(new_n22730), .Y(po1110));
  xnor_4 g22077(.A(new_n16310), .B(new_n16286), .Y(po1111));
  nand_5 g22078(.A(new_n20423), .B(new_n20422), .Y(new_n24427));
  xnor_4 g22079(.A(new_n24427), .B(new_n20439), .Y(po1112));
  not_8  g22080(.A(new_n22920), .Y(new_n24429));
  nand_5 g22081(.A(new_n22922), .B(new_n24429), .Y(new_n24430));
  nand_5 g22082(.A(new_n22920), .B(new_n22907), .Y(new_n24431));
  nand_5 g22083(.A(new_n24431), .B(new_n24430), .Y(po1113));
  xor_4  g22084(.A(new_n15304), .B(new_n11626), .Y(po1114));
  xor_4  g22085(.A(new_n12263), .B(new_n17770), .Y(po1115));
  xnor_4 g22086(.A(new_n3412), .B(new_n3411), .Y(po1116));
  xor_4  g22087(.A(new_n23544), .B(new_n23521), .Y(po1117));
  xor_4  g22088(.A(new_n21168), .B(new_n21167), .Y(po1118));
  xnor_4 g22089(.A(new_n16975), .B(new_n16972), .Y(po1119));
  nor_5  g22090(.A(new_n18938), .B(new_n18928), .Y(new_n24439));
  nor_5  g22091(.A(new_n24439), .B(new_n18937), .Y(new_n24440));
  nor_5  g22092(.A(new_n18936), .B(new_n18928), .Y(new_n24441));
  nor_5  g22093(.A(new_n24441), .B(new_n24440), .Y(po1120));
  xor_4  g22094(.A(new_n20437), .B(new_n20426), .Y(po1121));
  xor_4  g22095(.A(new_n21178), .B(new_n2789), .Y(po1122));
  nand_5 g22096(.A(new_n19443), .B(new_n19441), .Y(new_n24445));
  xor_4  g22097(.A(new_n24445), .B(new_n19435), .Y(po1123));
  xnor_4 g22098(.A(new_n6398), .B(new_n6395), .Y(po1124));
  xnor_4 g22099(.A(new_n19953), .B(new_n17237), .Y(po1125));
  nand_5 g22100(.A(new_n21275), .B(new_n22041), .Y(new_n24449));
  nand_5 g22101(.A(new_n22039), .B(new_n21276), .Y(new_n24450));
  nand_5 g22102(.A(new_n24450), .B(new_n24449), .Y(po1126));
  xnor_4 g22103(.A(new_n21365), .B(new_n7810), .Y(po1127));
  xor_4  g22104(.A(new_n18892), .B(new_n18891), .Y(po1128));
  xor_4  g22105(.A(new_n14138), .B(new_n6565), .Y(po1129));
  xor_4  g22106(.A(new_n18430), .B(new_n18427), .Y(po1130));
  not_8  g22107(.A(new_n14924), .Y(new_n24456));
  nand_5 g22108(.A(new_n14929), .B(new_n24456), .Y(po1131));
  xnor_4 g22109(.A(new_n19846), .B(new_n19845), .Y(po1132));
  xor_4  g22110(.A(new_n13607), .B(new_n13606), .Y(po1133));
  xor_4  g22111(.A(new_n11841), .B(new_n11840), .Y(po1134));
  xnor_4 g22112(.A(new_n21810), .B(new_n21807), .Y(po1135));
  xor_4  g22113(.A(new_n12188), .B(new_n12139), .Y(po1136));
  nand_5 g22114(.A(new_n17797), .B(new_n17795), .Y(new_n24463));
  xor_4  g22115(.A(new_n24463), .B(new_n12231), .Y(po1137));
  nand_5 g22116(.A(new_n23145), .B(new_n23141), .Y(new_n24465));
  not_8  g22117(.A(new_n23145), .Y(new_n24466));
  nand_5 g22118(.A(new_n24466), .B(new_n23139), .Y(new_n24467));
  nand_5 g22119(.A(new_n24467), .B(new_n24465), .Y(po1138));
  xor_4  g22120(.A(new_n20971), .B(new_n19813), .Y(po1139));
  nor_5  g22121(.A(new_n8291), .B(new_n8214), .Y(new_n24470));
  nor_5  g22122(.A(new_n24470), .B(new_n22539), .Y(po1140));
  xnor_4 g22123(.A(new_n12184), .B(new_n12183), .Y(po1141));
  not_8  g22124(.A(new_n10633), .Y(new_n24473));
  nor_5  g22125(.A(new_n24473), .B(new_n10560), .Y(new_n24474));
  nor_5  g22126(.A(new_n10633), .B(new_n10559), .Y(new_n24475));
  nor_5  g22127(.A(new_n24475), .B(new_n24474), .Y(po1142));
  xor_4  g22128(.A(new_n11359), .B(new_n5161), .Y(po1143));
  xor_4  g22129(.A(new_n19626), .B(new_n19623), .Y(po1144));
  xnor_4 g22130(.A(new_n22785), .B(new_n22767), .Y(po1145));
  xnor_4 g22131(.A(new_n15787), .B(new_n15785), .Y(po1146));
  xor_4  g22132(.A(new_n13511), .B(new_n5782), .Y(po1147));
  xor_4  g22133(.A(new_n20808), .B(new_n6014), .Y(po1148));
  xor_4  g22134(.A(new_n8244), .B(new_n8243), .Y(po1149));
  xor_4  g22135(.A(new_n7691), .B(new_n7688), .Y(po1150));
  xnor_4 g22136(.A(new_n5017), .B(new_n5016), .Y(po1151));
  nand_5 g22137(.A(new_n20712), .B(new_n20711), .Y(new_n24486));
  xor_4  g22138(.A(new_n24486), .B(new_n20713), .Y(po1153));
  nand_5 g22139(.A(new_n15823), .B(new_n15739), .Y(new_n24488));
  not_8  g22140(.A(new_n15823), .Y(new_n24489));
  nand_5 g22141(.A(new_n24489), .B(new_n15738), .Y(new_n24490));
  nand_5 g22142(.A(new_n24490), .B(new_n24488), .Y(po1154));
  nand_5 g22143(.A(new_n23549), .B(new_n23547), .Y(new_n24492));
  nand_5 g22144(.A(new_n24492), .B(new_n23545), .Y(po1155));
  xor_4  g22145(.A(new_n18258), .B(new_n18256), .Y(po1156));
  xor_4  g22146(.A(new_n20113), .B(new_n20085), .Y(po1157));
  xnor_4 g22147(.A(new_n3353), .B(new_n3352), .Y(po1158));
  xor_4  g22148(.A(new_n16842), .B(new_n16841), .Y(po1159));
  xnor_4 g22149(.A(new_n6523), .B(new_n6522), .Y(po1160));
  nand_5 g22150(.A(new_n21201), .B(new_n21203), .Y(new_n24499));
  xnor_4 g22151(.A(new_n24499), .B(new_n21200), .Y(po1161));
  xor_4  g22152(.A(new_n14133), .B(new_n6536), .Y(po1162));
  xnor_4 g22153(.A(new_n8515), .B(new_n8514), .Y(po1163));
  nand_5 g22154(.A(new_n21187), .B(new_n21186), .Y(new_n24503));
  xor_4  g22155(.A(new_n24503), .B(new_n2741), .Y(po1164));
  nor_5  g22156(.A(new_n15318), .B(new_n11558), .Y(new_n24505));
  nor_5  g22157(.A(new_n15320), .B(new_n15288), .Y(new_n24506));
  nor_5  g22158(.A(new_n24506), .B(new_n24505), .Y(po1165));
  not_8  g22159(.A(new_n4117), .Y(new_n24508));
  xor_4  g22160(.A(new_n6182), .B(new_n24508), .Y(po1166));
  xor_4  g22161(.A(new_n24266), .B(new_n13310), .Y(po1167));
  xnor_4 g22162(.A(new_n16308), .B(new_n16289), .Y(po1168));
  xnor_4 g22163(.A(new_n23250), .B(new_n18610), .Y(po1169));
  xor_4  g22164(.A(new_n22274), .B(new_n22271), .Y(po1170));
  nor_5  g22165(.A(new_n10111), .B(new_n10110), .Y(new_n24514));
  xor_4  g22166(.A(new_n24514), .B(new_n10134), .Y(po1171));
  xnor_4 g22167(.A(new_n15215), .B(new_n15190), .Y(po1172));
  xnor_4 g22168(.A(new_n8707), .B(new_n6672), .Y(po1173));
  or_6   g22169(.A(new_n20048), .B(new_n20046), .Y(new_n24518));
  nand_5 g22170(.A(new_n23823), .B(new_n20026), .Y(new_n24519));
  nor_5  g22171(.A(new_n24519), .B(new_n24518), .Y(new_n24520));
  nand_5 g22172(.A(new_n23824), .B(new_n20025), .Y(new_n24521));
  not_8  g22173(.A(new_n24521), .Y(new_n24522));
  nand_5 g22174(.A(new_n24522), .B(new_n20048), .Y(new_n24523));
  nor_5  g22175(.A(new_n24523), .B(new_n20046), .Y(new_n24524));
  or_6   g22176(.A(new_n24524), .B(new_n24520), .Y(po1174));
  nand_5 g22177(.A(new_n23140), .B(new_n23120), .Y(new_n24526));
  xor_4  g22178(.A(new_n24526), .B(new_n23137), .Y(po1175));
  xor_4  g22179(.A(new_n5422), .B(new_n5421), .Y(po1176));
  xor_4  g22180(.A(new_n20829), .B(new_n20828), .Y(po1177));
  xor_4  g22181(.A(new_n24410), .B(new_n24404), .Y(po1178));
  nor_5  g22182(.A(new_n23788), .B(new_n23783), .Y(new_n24531));
  nor_5  g22183(.A(new_n23785), .B(new_n22652), .Y(new_n24532));
  nor_5  g22184(.A(new_n24532), .B(new_n24531), .Y(po1179));
  not_8  g22185(.A(new_n20877), .Y(new_n24534));
  nand_5 g22186(.A(new_n20880), .B(new_n24534), .Y(new_n24535));
  xor_4  g22187(.A(new_n24535), .B(new_n20868), .Y(po1180));
  xor_4  g22188(.A(new_n24236), .B(new_n24232), .Y(po1181));
  xor_4  g22189(.A(new_n23462), .B(new_n23453), .Y(po1182));
  xnor_4 g22190(.A(new_n6213), .B(new_n6212), .Y(po1183));
  nand_5 g22191(.A(new_n7295), .B(pi068), .Y(new_n24540));
  not_8  g22192(.A(new_n24540), .Y(new_n24541));
  nand_5 g22193(.A(pi582), .B(new_n16941), .Y(new_n24542));
  not_8  g22194(.A(new_n24542), .Y(new_n24543));
  nand_5 g22195(.A(new_n2978), .B(pi349), .Y(new_n24544));
  not_8  g22196(.A(new_n24544), .Y(new_n24545));
  nor_5  g22197(.A(new_n22299), .B(new_n22294), .Y(new_n24546));
  nor_5  g22198(.A(new_n24546), .B(new_n24545), .Y(new_n24547));
  nor_5  g22199(.A(new_n24547), .B(new_n24543), .Y(new_n24548));
  nor_5  g22200(.A(new_n24548), .B(new_n24541), .Y(new_n24549));
  nand_5 g22201(.A(new_n24549), .B(new_n23349), .Y(new_n24550));
  not_8  g22202(.A(new_n22154), .Y(new_n24551));
  nand_5 g22203(.A(new_n24542), .B(new_n24540), .Y(new_n24552));
  xor_4  g22204(.A(new_n24552), .B(new_n24547), .Y(new_n24553));
  or_6   g22205(.A(new_n24553), .B(new_n24551), .Y(new_n24554));
  or_6   g22206(.A(new_n22300), .B(new_n20458), .Y(new_n24555));
  nand_5 g22207(.A(new_n22301), .B(new_n22292), .Y(new_n24556));
  nand_5 g22208(.A(new_n24556), .B(new_n24555), .Y(new_n24557));
  xor_4  g22209(.A(new_n24553), .B(new_n24551), .Y(new_n24558));
  nand_5 g22210(.A(new_n24558), .B(new_n24557), .Y(new_n24559));
  nand_5 g22211(.A(new_n24559), .B(new_n24554), .Y(new_n24560));
  not_8  g22212(.A(new_n24560), .Y(new_n24561));
  nor_5  g22213(.A(new_n24561), .B(new_n24550), .Y(new_n24562));
  not_8  g22214(.A(new_n23349), .Y(new_n24563));
  nand_5 g22215(.A(new_n24561), .B(new_n24563), .Y(new_n24564));
  not_8  g22216(.A(new_n24564), .Y(new_n24565));
  nor_5  g22217(.A(new_n24565), .B(new_n24562), .Y(new_n24566));
  nor_5  g22218(.A(new_n24549), .B(new_n23363), .Y(new_n24567));
  or_6   g22219(.A(new_n24549), .B(new_n23349), .Y(new_n24568));
  and_6  g22220(.A(new_n24568), .B(new_n23363), .Y(new_n24569));
  nor_5  g22221(.A(new_n24569), .B(new_n24567), .Y(new_n24570));
  nand_5 g22222(.A(new_n24568), .B(new_n24550), .Y(new_n24571));
  nand_5 g22223(.A(new_n24571), .B(new_n24570), .Y(new_n24572));
  nor_5  g22224(.A(new_n24572), .B(new_n24566), .Y(po1184));
  xnor_4 g22225(.A(new_n22723), .B(new_n22708), .Y(po1185));
  xor_4  g22226(.A(new_n17312), .B(new_n14419), .Y(po1186));
  xnor_4 g22227(.A(new_n19984), .B(new_n19982), .Y(po1187));
  nor_5  g22228(.A(new_n23887), .B(new_n22138), .Y(new_n24577));
  nor_5  g22229(.A(new_n23893), .B(new_n24577), .Y(po1188));
  xor_4  g22230(.A(new_n22887), .B(new_n22886), .Y(po1189));
  xnor_4 g22231(.A(new_n8626), .B(new_n8625), .Y(po1190));
  nor_5  g22232(.A(new_n23631), .B(new_n23518), .Y(new_n24581));
  or_6   g22233(.A(new_n24581), .B(po0712), .Y(new_n24582));
  not_8  g22234(.A(new_n23519), .Y(new_n24583));
  nor_5  g22235(.A(new_n23623), .B(new_n24583), .Y(new_n24584));
  nand_5 g22236(.A(new_n24584), .B(new_n23629), .Y(new_n24585));
  nand_5 g22237(.A(new_n24585), .B(new_n24582), .Y(po1191));
  xor_4  g22238(.A(new_n9878), .B(new_n7931), .Y(po1192));
  xor_4  g22239(.A(new_n15076), .B(new_n15063), .Y(po1193));
  xor_4  g22240(.A(new_n19316), .B(new_n19289), .Y(po1194));
  xor_4  g22241(.A(new_n15920), .B(new_n10507), .Y(po1195));
  xor_4  g22242(.A(new_n21771), .B(new_n9843), .Y(po1196));
  xor_4  g22243(.A(new_n7435), .B(new_n7427), .Y(po1197));
  xor_4  g22244(.A(new_n4487), .B(new_n4486), .Y(po1198));
  xor_4  g22245(.A(new_n14769), .B(new_n14748), .Y(po1199));
  nand_5 g22246(.A(new_n22736), .B(new_n21832), .Y(new_n24595));
  nand_5 g22247(.A(new_n22739), .B(new_n21831), .Y(new_n24596));
  nand_5 g22248(.A(new_n24596), .B(new_n24595), .Y(po1200));
  xor_4  g22249(.A(new_n9634), .B(new_n9624), .Y(po1201));
  xor_4  g22250(.A(new_n16837), .B(new_n16836), .Y(po1202));
  xor_4  g22251(.A(new_n20381), .B(new_n19558), .Y(po1203));
  xor_4  g22252(.A(new_n14142), .B(new_n14140), .Y(po1204));
  xnor_4 g22253(.A(new_n20621), .B(new_n20585), .Y(po1205));
  xor_4  g22254(.A(new_n20326), .B(new_n9446), .Y(po1206));
  xnor_4 g22255(.A(new_n20434), .B(new_n20433), .Y(po1207));
  nor_5  g22256(.A(new_n16473), .B(new_n16472), .Y(new_n24605));
  xor_4  g22257(.A(new_n24605), .B(new_n4244), .Y(po1208));
  xor_4  g22258(.A(new_n15575), .B(new_n15574), .Y(po1209));
  xor_4  g22259(.A(new_n12060), .B(new_n12025), .Y(po1210));
  xnor_4 g22260(.A(new_n7682), .B(new_n7681), .Y(po1211));
  xnor_4 g22261(.A(new_n3419), .B(new_n3414), .Y(po1212));
  nand_5 g22262(.A(new_n8524), .B(new_n8523), .Y(new_n24611));
  xnor_4 g22263(.A(new_n24611), .B(new_n8530), .Y(po1213));
  nand_5 g22264(.A(new_n11892), .B(new_n11887), .Y(new_n24613));
  xor_4  g22265(.A(new_n24613), .B(new_n11891), .Y(po1214));
  xnor_4 g22266(.A(new_n7477), .B(new_n7476), .Y(po1215));
  xnor_4 g22267(.A(new_n17651), .B(new_n17650), .Y(po1216));
  xnor_4 g22268(.A(new_n20230), .B(new_n20227), .Y(po1217));
  nand_5 g22269(.A(new_n24466), .B(new_n13821), .Y(new_n24618));
  nand_5 g22270(.A(new_n17984), .B(new_n17981), .Y(new_n24619));
  nand_5 g22271(.A(new_n24619), .B(new_n17965), .Y(new_n24620));
  xor_4  g22272(.A(new_n23145), .B(new_n13820), .Y(new_n24621));
  nand_5 g22273(.A(new_n24621), .B(new_n24620), .Y(new_n24622));
  nand_5 g22274(.A(new_n24622), .B(new_n24618), .Y(po1218));
  nor_5  g22275(.A(new_n22345), .B(new_n21834), .Y(new_n24624));
  xor_4  g22276(.A(new_n22345), .B(new_n21840), .Y(new_n24625));
  nand_5 g22277(.A(new_n22350), .B(new_n21834), .Y(new_n24626));
  nand_5 g22278(.A(new_n23754), .B(new_n23751), .Y(new_n24627));
  nand_5 g22279(.A(new_n24627), .B(new_n24626), .Y(new_n24628));
  not_8  g22280(.A(new_n24628), .Y(new_n24629));
  nor_5  g22281(.A(new_n24629), .B(new_n24625), .Y(new_n24630));
  nor_5  g22282(.A(new_n24630), .B(new_n24624), .Y(po1219));
  xnor_4 g22283(.A(new_n22277), .B(new_n22276), .Y(po1220));
  xor_4  g22284(.A(new_n12315), .B(new_n6513), .Y(po1221));
  xor_4  g22285(.A(new_n15317), .B(new_n15316), .Y(po1222));
  xor_4  g22286(.A(new_n22801), .B(new_n4935), .Y(po1223));
  xnor_4 g22287(.A(new_n19039), .B(new_n19014), .Y(po1224));
  xnor_4 g22288(.A(new_n17299), .B(new_n13471), .Y(po1225));
  xnor_4 g22289(.A(new_n19027), .B(new_n19026), .Y(po1226));
  xor_4  g22290(.A(new_n22546), .B(new_n22542), .Y(po1227));
  xnor_4 g22291(.A(new_n24558), .B(new_n24557), .Y(po1228));
  xor_4  g22292(.A(new_n4214), .B(new_n4212), .Y(po1229));
  xor_4  g22293(.A(new_n19966), .B(new_n17229), .Y(po1230));
  xnor_4 g22294(.A(new_n13609), .B(new_n13594), .Y(po1231));
  xor_4  g22295(.A(new_n16481), .B(new_n5443), .Y(po1232));
  xnor_4 g22296(.A(new_n7144), .B(new_n7132), .Y(po1233));
  xnor_4 g22297(.A(new_n11488), .B(new_n11457), .Y(po1234));
  xor_4  g22298(.A(new_n11272), .B(new_n8804), .Y(po1235));
  xor_4  g22299(.A(new_n19031), .B(new_n4970), .Y(po1236));
  xor_4  g22300(.A(new_n13472), .B(new_n13471), .Y(po1237));
  xor_4  g22301(.A(new_n4119), .B(new_n24508), .Y(po1238));
  xnor_4 g22302(.A(new_n21760), .B(new_n21759), .Y(po1239));
  nor_5  g22303(.A(new_n21243), .B(new_n20861), .Y(new_n24652));
  nor_5  g22304(.A(new_n21266), .B(new_n21245), .Y(new_n24653));
  nor_5  g22305(.A(new_n24653), .B(new_n24652), .Y(po1240));
  xor_4  g22306(.A(new_n23329), .B(new_n23328), .Y(po1241));
  nand_5 g22307(.A(new_n18132), .B(new_n18131), .Y(new_n24656));
  xor_4  g22308(.A(new_n24656), .B(new_n18147), .Y(po1242));
  and_6  g22309(.A(new_n21224), .B(new_n19860), .Y(new_n24658));
  nor_5  g22310(.A(new_n24000), .B(new_n23997), .Y(new_n24659));
  nor_5  g22311(.A(new_n24659), .B(new_n24658), .Y(po1244));
  not_8  g22312(.A(new_n24566), .Y(new_n24661));
  nor_5  g22313(.A(new_n24661), .B(new_n23363), .Y(new_n24662));
  nand_5 g22314(.A(new_n24570), .B(new_n24561), .Y(new_n24663));
  nand_5 g22315(.A(new_n24562), .B(new_n23363), .Y(new_n24664));
  nand_5 g22316(.A(new_n24664), .B(new_n24663), .Y(new_n24665));
  nor_5  g22317(.A(new_n24665), .B(new_n24662), .Y(po1245));
  nand_5 g22318(.A(new_n18357), .B(new_n18356), .Y(new_n24667));
  xor_4  g22319(.A(new_n24667), .B(new_n18360), .Y(po1246));
  xnor_4 g22320(.A(new_n23745), .B(new_n23736), .Y(po1247));
  xnor_4 g22321(.A(new_n20168), .B(new_n20167), .Y(po1248));
  xor_4  g22322(.A(new_n24363), .B(new_n14384), .Y(po1249));
  xor_4  g22323(.A(new_n10610), .B(new_n10603), .Y(po1250));
  xnor_4 g22324(.A(new_n20897), .B(new_n15016), .Y(po1251));
  xnor_4 g22325(.A(new_n8961), .B(new_n8960), .Y(po1252));
  xor_4  g22326(.A(new_n17895), .B(new_n17894), .Y(po1253));
  nand_5 g22327(.A(new_n7233), .B(new_n7217), .Y(new_n24676));
  nor_5  g22328(.A(new_n7238), .B(new_n7216), .Y(new_n24677));
  nand_5 g22329(.A(new_n24677), .B(new_n24676), .Y(new_n24678));
  not_8  g22330(.A(new_n7235), .Y(new_n24679));
  nand_5 g22331(.A(new_n24679), .B(new_n7216), .Y(new_n24680));
  nand_5 g22332(.A(new_n24680), .B(new_n24678), .Y(new_n24681));
  not_8  g22333(.A(new_n7241), .Y(new_n24682));
  nand_5 g22334(.A(new_n24682), .B(new_n7216), .Y(new_n24683));
  nor_5  g22335(.A(new_n7236), .B(new_n7215), .Y(new_n24684));
  nand_5 g22336(.A(new_n24684), .B(new_n24683), .Y(new_n24685));
  not_8  g22337(.A(new_n7236), .Y(new_n24686));
  nor_5  g22338(.A(new_n24686), .B(new_n7213), .Y(new_n24687));
  nand_5 g22339(.A(new_n7238), .B(new_n7215), .Y(new_n24688));
  nor_5  g22340(.A(new_n24688), .B(new_n24687), .Y(new_n24689));
  nand_5 g22341(.A(new_n24689), .B(new_n7235), .Y(new_n24690));
  nand_5 g22342(.A(new_n24690), .B(new_n24685), .Y(new_n24691));
  nor_5  g22343(.A(new_n24691), .B(new_n24681), .Y(po1254));
  xor_4  g22344(.A(new_n17892), .B(new_n17891), .Y(po1255));
  xor_4  g22345(.A(new_n10368), .B(new_n10358), .Y(po1256));
  xor_4  g22346(.A(pi708), .B(new_n4088), .Y(new_n24695));
  xor_4  g22347(.A(new_n24695), .B(new_n8928), .Y(po1257));
  xnor_4 g22348(.A(new_n4505), .B(new_n4435), .Y(po1258));
  xor_4  g22349(.A(new_n8438), .B(new_n8437), .Y(po1259));
  xnor_4 g22350(.A(new_n10618), .B(new_n10590), .Y(po1260));
  xor_4  g22351(.A(new_n23246), .B(new_n23242), .Y(po1261));
  not_8  g22352(.A(new_n18302), .Y(new_n24701));
  nor_5  g22353(.A(new_n18376), .B(new_n24701), .Y(po1262));
  xnor_4 g22354(.A(new_n24408), .B(new_n24406), .Y(po1263));
  xor_4  g22355(.A(new_n8504), .B(new_n8502), .Y(po1264));
  xnor_4 g22356(.A(new_n17413), .B(new_n17412), .Y(po1265));
  xor_4  g22357(.A(new_n8945), .B(new_n8919), .Y(po1266));
  xor_4  g22358(.A(new_n12196), .B(new_n12197), .Y(po1267));
  xor_4  g22359(.A(new_n19503), .B(new_n19502), .Y(po1268));
  xor_4  g22360(.A(new_n23273), .B(new_n24028), .Y(po1269));
  xor_4  g22361(.A(new_n2548), .B(new_n2547), .Y(po1270));
  xor_4  g22362(.A(new_n23806), .B(new_n9066), .Y(po1272));
  xor_4  g22363(.A(new_n9826), .B(new_n9825), .Y(po1273));
  xor_4  g22364(.A(new_n20100), .B(new_n16796), .Y(po1274));
  xor_4  g22365(.A(new_n10389), .B(new_n10327), .Y(po1275));
  xnor_4 g22366(.A(new_n14792), .B(new_n14791), .Y(po1276));
  nand_5 g22367(.A(new_n7154), .B(new_n7155), .Y(new_n24716));
  xor_4  g22368(.A(new_n24716), .B(new_n7157), .Y(po1277));
  xnor_4 g22369(.A(new_n12676), .B(new_n12559), .Y(po1278));
  xor_4  g22370(.A(new_n5763), .B(new_n5689), .Y(po1279));
  xor_4  g22371(.A(new_n19630), .B(new_n4522), .Y(new_n24720));
  xor_4  g22372(.A(new_n24720), .B(new_n19629), .Y(po1280));
  xor_4  g22373(.A(new_n13139), .B(new_n4145), .Y(po1282));
  xnor_4 g22374(.A(new_n18566), .B(new_n18565), .Y(po1283));
  xor_4  g22375(.A(new_n17277), .B(new_n17211), .Y(po1284));
  xor_4  g22376(.A(new_n24629), .B(new_n24625), .Y(po1285));
  xor_4  g22377(.A(new_n17954), .B(new_n7913), .Y(po1286));
  xor_4  g22378(.A(new_n14804), .B(new_n10469), .Y(new_n24727));
  xor_4  g22379(.A(new_n24727), .B(new_n18966), .Y(po1288));
  xnor_4 g22380(.A(new_n16466), .B(new_n5421), .Y(po1289));
  nand_5 g22381(.A(new_n17731), .B(new_n17730), .Y(new_n24730));
  xor_4  g22382(.A(new_n24730), .B(new_n17734), .Y(po1290));
  xnor_4 g22383(.A(new_n15397), .B(new_n15390), .Y(po1291));
  xor_4  g22384(.A(new_n17785), .B(new_n12278), .Y(po1292));
  xor_4  g22385(.A(new_n23352), .B(new_n24563), .Y(new_n24734));
  xor_4  g22386(.A(new_n24734), .B(new_n23356), .Y(po1293));
  xnor_4 g22387(.A(new_n5447), .B(new_n5446), .Y(po1294));
  xnor_4 g22388(.A(new_n21562), .B(new_n21559), .Y(po1295));
  xor_4  g22389(.A(new_n9456), .B(new_n4887), .Y(po1296));
  and_6  g22390(.A(new_n21914), .B(new_n7581), .Y(new_n24739));
  or_6   g22391(.A(new_n24739), .B(new_n21936), .Y(new_n24740));
  and_6  g22392(.A(new_n24740), .B(new_n21939), .Y(po1297));
  xor_4  g22393(.A(new_n19719), .B(new_n15419), .Y(po1298));
  xnor_4 g22394(.A(new_n15803), .B(new_n15801), .Y(po1299));
  xor_4  g22395(.A(new_n13465), .B(new_n13464), .Y(po1300));
  xor_4  g22396(.A(new_n17792), .B(new_n17766), .Y(po1301));
  nand_5 g22397(.A(new_n20642), .B(new_n22175), .Y(new_n24746));
  nand_5 g22398(.A(new_n24746), .B(new_n22173), .Y(new_n24747));
  nand_5 g22399(.A(new_n22174), .B(new_n20642), .Y(new_n24748));
  and_6  g22400(.A(new_n24748), .B(new_n24747), .Y(po1302));
  xnor_4 g22401(.A(new_n18881), .B(new_n18867), .Y(po1303));
  or_6   g22402(.A(new_n22322), .B(new_n21226), .Y(new_n24751));
  nand_5 g22403(.A(new_n24014), .B(new_n21221), .Y(new_n24752));
  nand_5 g22404(.A(new_n24752), .B(new_n24751), .Y(po1304));
  xnor_4 g22405(.A(new_n17275), .B(new_n17274), .Y(po1305));
  xnor_4 g22406(.A(new_n21576), .B(new_n21575), .Y(po1306));
  nand_5 g22407(.A(new_n18173), .B(new_n18170), .Y(new_n24756));
  nor_5  g22408(.A(new_n24756), .B(new_n8047), .Y(new_n24757));
  nand_5 g22409(.A(new_n24757), .B(new_n18187), .Y(new_n24758));
  nand_5 g22410(.A(new_n18192), .B(new_n18177), .Y(new_n24759));
  and_6  g22411(.A(new_n24759), .B(new_n24758), .Y(new_n24760));
  and_6  g22412(.A(new_n24760), .B(po0242), .Y(po1307));
  nand_5 g22413(.A(new_n21162), .B(new_n21149), .Y(new_n24762));
  xnor_4 g22414(.A(new_n24762), .B(new_n21161), .Y(po1308));
  xor_4  g22415(.A(new_n7452), .B(new_n7451), .Y(po1309));
  xor_4  g22416(.A(new_n20095), .B(new_n20094), .Y(po1310));
  xor_4  g22417(.A(new_n21454), .B(new_n21429), .Y(po1311));
  xnor_4 g22418(.A(new_n3090), .B(new_n3074), .Y(po1312));
  xnor_4 g22419(.A(new_n12052), .B(new_n12040), .Y(po1313));
  xor_4  g22420(.A(new_n22433), .B(new_n3394), .Y(po1314));
  xnor_4 g22421(.A(new_n23055), .B(new_n23053), .Y(po1315));
  xnor_4 g22422(.A(new_n12054), .B(new_n12035), .Y(po1316));
  xnor_4 g22423(.A(new_n13366), .B(new_n13365), .Y(po1317));
  xnor_4 g22424(.A(new_n19423), .B(new_n19406), .Y(po1318));
  xor_4  g22425(.A(new_n22797), .B(new_n4928), .Y(po1319));
  nor_5  g22426(.A(new_n24076), .B(new_n24073), .Y(po1320));
  nand_5 g22427(.A(new_n21870), .B(new_n21869), .Y(new_n24776));
  xnor_4 g22428(.A(new_n24776), .B(new_n21874), .Y(po1321));
  xor_4  g22429(.A(new_n7445), .B(new_n7422), .Y(po1323));
  xnor_4 g22430(.A(new_n3377), .B(new_n3376), .Y(po1325));
  xor_4  g22431(.A(new_n15246), .B(new_n9626), .Y(po1326));
  xor_4  g22432(.A(new_n13114), .B(new_n6063), .Y(po1327));
  xor_4  g22433(.A(new_n16933), .B(new_n16923), .Y(po1328));
  xnor_4 g22434(.A(new_n13361), .B(new_n13360), .Y(po1329));
  nand_5 g22435(.A(new_n18008), .B(new_n18007), .Y(new_n24784));
  xnor_4 g22436(.A(new_n24784), .B(new_n18019), .Y(po1330));
  xnor_4 g22437(.A(new_n19127), .B(new_n19107), .Y(po1331));
  xor_4  g22438(.A(new_n22952), .B(new_n18633), .Y(po1332));
  xor_4  g22439(.A(new_n17318), .B(new_n14417), .Y(po1333));
  nand_5 g22440(.A(new_n13268), .B(new_n13266), .Y(new_n24789));
  xor_4  g22441(.A(new_n24789), .B(new_n13256), .Y(po1334));
  xnor_4 g22442(.A(new_n23984), .B(new_n23983), .Y(po1335));
  xor_4  g22443(.A(new_n20814), .B(new_n6043), .Y(po1336));
  xor_4  g22444(.A(new_n15909), .B(new_n10510), .Y(po1337));
  xor_4  g22445(.A(new_n12387), .B(new_n11170), .Y(po1338));
  nand_5 g22446(.A(new_n12027), .B(new_n12028), .Y(new_n24795));
  xor_4  g22447(.A(new_n24795), .B(new_n12058), .Y(po1339));
  nand_5 g22448(.A(new_n18548), .B(new_n18547), .Y(new_n24797));
  xor_4  g22449(.A(new_n24797), .B(new_n16098), .Y(po1340));
  xor_4  g22450(.A(new_n15311), .B(new_n11564), .Y(po1341));
  xor_4  g22451(.A(new_n20357), .B(new_n19571), .Y(po1342));
  nand_5 g22452(.A(new_n21817), .B(new_n21815), .Y(new_n24801));
  xnor_4 g22453(.A(new_n24801), .B(new_n21816), .Y(po1343));
  xnor_4 g22454(.A(new_n22493), .B(new_n22492), .Y(po1344));
  xnor_4 g22455(.A(new_n13008), .B(new_n13007), .Y(po1345));
  xor_4  g22456(.A(new_n24258), .B(new_n13370), .Y(new_n24805));
  xor_4  g22457(.A(new_n24805), .B(new_n24262), .Y(po1346));
  xor_4  g22458(.A(new_n9369), .B(new_n9368), .Y(po1347));
  nor_5  g22459(.A(new_n20951), .B(new_n20930), .Y(po1348));
  xor_4  g22460(.A(new_n14772), .B(new_n14771), .Y(po1349));
  xor_4  g22461(.A(new_n24114), .B(new_n24112), .Y(po1350));
  xor_4  g22462(.A(new_n17898), .B(new_n17897), .Y(po1351));
  nand_5 g22463(.A(new_n24689), .B(new_n18665), .Y(new_n24812));
  nand_5 g22464(.A(new_n24812), .B(new_n24683), .Y(po1352));
  xnor_4 g22465(.A(new_n19508), .B(new_n19507), .Y(po1353));
  xnor_4 g22466(.A(new_n4649), .B(new_n4648), .Y(po1354));
  xor_4  g22467(.A(new_n12048), .B(new_n3857), .Y(po1355));
  nand_5 g22468(.A(new_n2519), .B(new_n2518), .Y(new_n24817));
  xnor_4 g22469(.A(new_n24817), .B(new_n2539), .Y(po1356));
  xor_4  g22470(.A(new_n16477), .B(new_n5435), .Y(po1357));
  xor_4  g22471(.A(new_n9638), .B(new_n9623), .Y(po1358));
  xnor_4 g22472(.A(new_n5012), .B(new_n4957), .Y(po1359));
  xor_4  g22473(.A(new_n18496), .B(new_n7133), .Y(po1360));
  nor_5  g22474(.A(new_n14059), .B(new_n14058), .Y(new_n24823));
  xor_4  g22475(.A(new_n24823), .B(new_n14072), .Y(po1361));
  xor_4  g22476(.A(new_n10938), .B(new_n10935), .Y(po1362));
  xor_4  g22477(.A(new_n13908), .B(new_n13879), .Y(po1363));
  xnor_4 g22478(.A(new_n12181), .B(new_n12179), .Y(po1364));
  xor_4  g22479(.A(new_n8452), .B(new_n22873), .Y(new_n24828));
  xor_4  g22480(.A(new_n24828), .B(new_n23368), .Y(po1365));
  xnor_4 g22481(.A(new_n10383), .B(new_n10341), .Y(po1366));
  xor_4  g22482(.A(new_n13800), .B(new_n13799), .Y(po1367));
  xnor_4 g22483(.A(new_n18582), .B(new_n18579), .Y(po1368));
  xnor_4 g22484(.A(new_n4663), .B(new_n4662), .Y(po1369));
  nand_5 g22485(.A(new_n2749), .B(new_n2751), .Y(new_n24834));
  xor_4  g22486(.A(new_n24834), .B(new_n2754), .Y(po1370));
  xnor_4 g22487(.A(new_n2760), .B(new_n2759), .Y(po1371));
  xor_4  g22488(.A(new_n20906), .B(new_n11283), .Y(po1372));
  xnor_4 g22489(.A(new_n14608), .B(new_n14607), .Y(po1373));
  xor_4  g22490(.A(new_n24061), .B(new_n22246), .Y(po1374));
  nand_5 g22491(.A(new_n22510), .B(new_n22499), .Y(new_n24840));
  nand_5 g22492(.A(new_n22531), .B(new_n24840), .Y(new_n24841));
  and_6  g22493(.A(new_n22522), .B(new_n22514), .Y(new_n24842));
  nand_5 g22494(.A(new_n24842), .B(new_n24841), .Y(new_n24843));
  nor_5  g22495(.A(new_n22535), .B(new_n22523), .Y(new_n24844));
  nand_5 g22496(.A(new_n24844), .B(new_n24843), .Y(po1375));
  xnor_4 g22497(.A(new_n22280), .B(new_n22279), .Y(po1376));
  xor_4  g22498(.A(new_n21999), .B(new_n21998), .Y(po1377));
  xor_4  g22499(.A(new_n20842), .B(new_n20787), .Y(po1378));
  nor_5  g22500(.A(new_n17289), .B(new_n17173), .Y(new_n24849));
  xnor_4 g22501(.A(new_n24849), .B(new_n17287), .Y(po1379));
  xor_4  g22502(.A(new_n20820), .B(new_n6052), .Y(po1380));
  xnor_4 g22503(.A(new_n23575), .B(new_n23574), .Y(po1381));
  not_8  g22504(.A(new_n15767), .Y(new_n24853));
  xor_4  g22505(.A(new_n16632), .B(new_n24853), .Y(po1382));
  xor_4  g22506(.A(new_n18067), .B(new_n7925), .Y(po1383));
  xnor_4 g22507(.A(new_n7676), .B(new_n7675), .Y(po1384));
  xor_4  g22508(.A(new_n10016), .B(new_n10015), .Y(po1385));
  nor_5  g22509(.A(new_n5154), .B(new_n5155), .Y(new_n24858));
  xor_4  g22510(.A(new_n24858), .B(new_n5170), .Y(po1386));
  xnor_4 g22511(.A(new_n3095), .B(new_n3065), .Y(po1387));
  xnor_4 g22512(.A(new_n6194), .B(new_n6180), .Y(po1388));
  xnor_4 g22513(.A(new_n9356), .B(new_n9355), .Y(po1389));
  xor_4  g22514(.A(new_n7492), .B(new_n7394), .Y(new_n24863));
  nand_5 g22515(.A(new_n7499), .B(new_n7495), .Y(new_n24864));
  xor_4  g22516(.A(new_n24864), .B(new_n7497), .Y(new_n24865));
  xor_4  g22517(.A(new_n24865), .B(new_n24863), .Y(po1390));
  xor_4  g22518(.A(new_n11831), .B(new_n11810), .Y(po1391));
  xor_4  g22519(.A(new_n21262), .B(new_n14179), .Y(po1392));
  xor_4  g22520(.A(new_n16581), .B(new_n12082), .Y(new_n24869));
  nand_5 g22521(.A(new_n16587), .B(new_n16574), .Y(new_n24870));
  xor_4  g22522(.A(new_n24870), .B(new_n24869), .Y(po1393));
  xor_4  g22523(.A(new_n24849), .B(new_n19997), .Y(po1394));
  xor_4  g22524(.A(new_n13352), .B(new_n13348), .Y(po1395));
  nor_5  g22525(.A(new_n18192), .B(new_n18186), .Y(new_n24874));
  xor_4  g22526(.A(new_n18175), .B(new_n8048), .Y(new_n24875));
  xor_4  g22527(.A(new_n24875), .B(new_n24874), .Y(po1396));
  xor_4  g22528(.A(new_n18884), .B(new_n18883), .Y(po1397));
  xor_4  g22529(.A(new_n24571), .B(new_n24561), .Y(po1398));
  xnor_4 g22530(.A(new_n21264), .B(new_n21248), .Y(po1399));
  xnor_4 g22531(.A(new_n15448), .B(new_n15445), .Y(po1401));
  xor_4  g22532(.A(new_n18668), .B(new_n18663), .Y(po1402));
  xor_4  g22533(.A(new_n18270), .B(new_n15360), .Y(po1403));
  xor_4  g22534(.A(new_n21460), .B(new_n21458), .Y(po1404));
  nor_5  g22535(.A(new_n23954), .B(new_n23950), .Y(new_n24884));
  xor_4  g22536(.A(new_n24884), .B(new_n23939), .Y(po1405));
  xor_4  g22537(.A(new_n21448), .B(new_n21434), .Y(po1406));
  xor_4  g22538(.A(new_n11234), .B(new_n4206), .Y(po1407));
  nor_5  g22539(.A(new_n23592), .B(new_n20993), .Y(po1408));
  xnor_4 g22540(.A(new_n11612), .B(new_n11611), .Y(po1409));
  xnor_4 g22541(.A(new_n9117), .B(new_n9116), .Y(po1410));
  xnor_4 g22542(.A(new_n14899), .B(new_n14877), .Y(po1411));
  xor_4  g22543(.A(new_n24853), .B(new_n15766), .Y(po1412));
  xor_4  g22544(.A(new_n7457), .B(new_n16897), .Y(po1413));
  xnor_4 g22545(.A(new_n14901), .B(new_n14873), .Y(po1414));
  xnor_4 g22546(.A(new_n20330), .B(new_n20328), .Y(po1415));
  xor_4  g22547(.A(new_n12382), .B(new_n8906), .Y(po1416));
  xnor_4 g22548(.A(new_n13673), .B(new_n3477), .Y(po1417));
  xor_4  g22549(.A(new_n20732), .B(new_n20730), .Y(po1418));
  xor_4  g22550(.A(new_n17397), .B(new_n21294), .Y(po1419));
  xor_4  g22551(.A(new_n21568), .B(new_n21567), .Y(po1420));
  xor_4  g22552(.A(new_n5413), .B(new_n5363), .Y(po1421));
  xor_4  g22553(.A(new_n13110), .B(new_n6055), .Y(po1422));
  nand_5 g22554(.A(new_n24521), .B(new_n24519), .Y(new_n24903));
  not_8  g22555(.A(new_n24903), .Y(new_n24904));
  nor_5  g22556(.A(new_n24904), .B(new_n23827), .Y(po1423));
  xnor_4 g22557(.A(new_n9364), .B(new_n9325), .Y(po1424));
  nand_5 g22558(.A(new_n20045), .B(new_n20027), .Y(new_n24907));
  and_6  g22559(.A(new_n23823), .B(new_n24907), .Y(new_n24908));
  nand_5 g22560(.A(new_n24908), .B(new_n24518), .Y(new_n24909));
  nor_5  g22561(.A(new_n24903), .B(new_n24518), .Y(new_n24910));
  nor_5  g22562(.A(new_n24910), .B(new_n24524), .Y(new_n24911));
  nand_5 g22563(.A(new_n24911), .B(new_n24909), .Y(po1425));
  xnor_4 g22564(.A(new_n9849), .B(new_n9799), .Y(po1426));
  nor_5  g22565(.A(new_n24255), .B(new_n13375), .Y(po1427));
  xor_4  g22566(.A(new_n15246), .B(new_n5773), .Y(po1428));
  xor_4  g22567(.A(new_n21349), .B(new_n18085), .Y(po1429));
  xor_4  g22568(.A(new_n8428), .B(new_n8401), .Y(po1430));
  xor_4  g22569(.A(new_n6923), .B(new_n6881), .Y(po1431));
  xor_4  g22570(.A(new_n6256), .B(new_n6227), .Y(po1432));
  xor_4  g22571(.A(new_n15626), .B(new_n12608), .Y(po1433));
  xnor_4 g22572(.A(new_n14447), .B(new_n14446), .Y(po1434));
  xor_4  g22573(.A(new_n8264), .B(new_n8263), .Y(po1435));
  xnor_4 g22574(.A(new_n24621), .B(new_n24620), .Y(po1436));
  xor_4  g22575(.A(new_n21782), .B(new_n9796), .Y(po1437));
  xnor_4 g22576(.A(new_n22135), .B(new_n22134), .Y(po1438));
  nor_5  g22577(.A(new_n14233), .B(new_n14225), .Y(new_n24926));
  xor_4  g22578(.A(new_n24926), .B(new_n9022), .Y(po1439));
  nor_5  g22579(.A(new_n18829), .B(new_n18758), .Y(new_n24928));
  nor_5  g22580(.A(new_n18905), .B(new_n18831), .Y(new_n24929));
  nor_5  g22581(.A(new_n24929), .B(new_n24928), .Y(po1440));
  xnor_4 g22582(.A(new_n23584), .B(new_n23583), .Y(po1441));
  nand_5 g22583(.A(new_n11766), .B(new_n11660), .Y(new_n24932));
  nor_5  g22584(.A(new_n11855), .B(new_n24932), .Y(po1442));
  xnor_4 g22585(.A(new_n11835), .B(new_n11803), .Y(po1443));
  xor_4  g22586(.A(new_n20852), .B(new_n11259), .Y(po1444));
  xor_4  g22587(.A(new_n17600), .B(new_n17578), .Y(po1445));
  xnor_4 g22588(.A(new_n3684), .B(new_n3683), .Y(po1446));
  xor_4  g22589(.A(new_n14421), .B(new_n14420), .Y(po1447));
  nand_5 g22590(.A(new_n23623), .B(new_n23625), .Y(new_n24939));
  xor_4  g22591(.A(new_n24939), .B(new_n23521), .Y(new_n24940));
  xor_4  g22592(.A(new_n24940), .B(new_n23628), .Y(po1448));
  xnor_4 g22593(.A(new_n12996), .B(new_n12994), .Y(po1449));
  xor_4  g22594(.A(new_n16155), .B(new_n16140), .Y(po1450));
  xor_4  g22595(.A(new_n21844), .B(new_n21841), .Y(po1451));
  xor_4  g22596(.A(new_n16179), .B(new_n16176), .Y(new_n24945));
  xor_4  g22597(.A(new_n24945), .B(new_n16193), .Y(po1452));
  nand_5 g22598(.A(new_n21271), .B(new_n10423), .Y(new_n24947));
  nand_5 g22599(.A(new_n24947), .B(new_n10416), .Y(new_n24948));
  and_6  g22600(.A(new_n24948), .B(new_n21274), .Y(new_n24949));
  nand_5 g22601(.A(new_n21277), .B(new_n10420), .Y(new_n24950));
  nand_5 g22602(.A(new_n24126), .B(new_n21276), .Y(new_n24951));
  nand_5 g22603(.A(new_n24951), .B(new_n24950), .Y(new_n24952));
  nor_5  g22604(.A(new_n24952), .B(new_n24949), .Y(po1453));
  or_6   g22605(.A(new_n19176), .B(new_n7392), .Y(new_n24954));
  nand_5 g22606(.A(new_n24954), .B(new_n19171), .Y(po1454));
  xor_4  g22607(.A(new_n20901), .B(new_n11276), .Y(po1455));
  nor_5  g22608(.A(new_n23977), .B(new_n22175), .Y(new_n24957));
  and_6  g22609(.A(new_n23986), .B(new_n23978), .Y(new_n24958));
  nor_5  g22610(.A(new_n24958), .B(new_n24957), .Y(po1456));
  xor_4  g22611(.A(pi718), .B(pi364), .Y(new_n24960));
  xor_4  g22612(.A(new_n24960), .B(new_n5347), .Y(po1457));
  xnor_4 g22613(.A(new_n14966), .B(new_n14951), .Y(po1458));
  xor_4  g22614(.A(new_n7211), .B(new_n7192), .Y(po1459));
  xor_4  g22615(.A(new_n21155), .B(new_n21154), .Y(po1460));
  xnor_4 g22616(.A(new_n10374), .B(new_n10351), .Y(po1461));
  xor_4  g22617(.A(new_n2545), .B(new_n2543), .Y(po1462));
  xor_4  g22618(.A(new_n15400), .B(new_n15386), .Y(po1463));
  xor_4  g22619(.A(new_n17251), .B(new_n5345), .Y(po1464));
  nand_5 g22620(.A(new_n23953), .B(new_n23949), .Y(new_n24969));
  xor_4  g22621(.A(new_n24969), .B(new_n22121), .Y(po1465));
  nand_5 g22622(.A(new_n23914), .B(new_n23915), .Y(new_n24971));
  nor_5  g22623(.A(new_n24971), .B(new_n23917), .Y(new_n24972));
  nand_5 g22624(.A(new_n23311), .B(new_n23298), .Y(new_n24973));
  nand_5 g22625(.A(new_n23918), .B(new_n24973), .Y(new_n24974));
  nor_5  g22626(.A(new_n24974), .B(new_n24972), .Y(po1466));
  xor_4  g22627(.A(new_n11824), .B(new_n4016), .Y(po1467));
  xnor_4 g22628(.A(new_n9722), .B(new_n9721), .Y(po1468));
  xnor_4 g22629(.A(new_n21180), .B(new_n21147), .Y(po1469));
  nand_5 g22630(.A(new_n5753), .B(new_n5749), .Y(new_n24979));
  and_6  g22631(.A(new_n24979), .B(new_n5751), .Y(new_n24980));
  nand_5 g22632(.A(new_n5753), .B(new_n5746), .Y(new_n24981));
  nand_5 g22633(.A(new_n24981), .B(new_n5633), .Y(new_n24982));
  nor_5  g22634(.A(new_n24982), .B(new_n24980), .Y(po1470));
  xor_4  g22635(.A(new_n15213), .B(new_n15195), .Y(po1471));
  xor_4  g22636(.A(new_n15893), .B(new_n5788), .Y(po1472));
  xnor_4 g22637(.A(new_n24390), .B(new_n24389), .Y(po1473));
  xor_4  g22638(.A(new_n9359), .B(new_n9358), .Y(po1474));
  nand_5 g22639(.A(new_n22185), .B(new_n19804), .Y(new_n24988));
  nand_5 g22640(.A(new_n22190), .B(new_n22186), .Y(new_n24989));
  nand_5 g22641(.A(new_n24989), .B(new_n24988), .Y(po1475));
  xor_4  g22642(.A(new_n22212), .B(new_n22208), .Y(po1476));
  xor_4  g22643(.A(new_n7956), .B(new_n11320), .Y(po1477));
  xor_4  g22644(.A(new_n13109), .B(new_n10695), .Y(po1478));
  xnor_4 g22645(.A(new_n22646), .B(new_n22645), .Y(po1479));
  xnor_4 g22646(.A(new_n3406), .B(new_n3404), .Y(po1480));
  xor_4  g22647(.A(new_n10955), .B(new_n10912), .Y(po1481));
  xnor_4 g22648(.A(new_n11339), .B(new_n11338), .Y(po1482));
  xor_4  g22649(.A(new_n24035), .B(new_n24034), .Y(po1483));
  nor_5  g22650(.A(new_n24203), .B(new_n7511), .Y(new_n24999));
  not_8  g22651(.A(new_n7384), .Y(new_n25000));
  nor_5  g22652(.A(new_n7511), .B(new_n25000), .Y(new_n25001));
  nand_5 g22653(.A(new_n19181), .B(new_n7505), .Y(new_n25002));
  nor_5  g22654(.A(new_n25002), .B(new_n25001), .Y(new_n25003));
  nor_5  g22655(.A(new_n25003), .B(new_n24999), .Y(po1484));
  xor_4  g22656(.A(new_n19327), .B(new_n19326), .Y(po1485));
  xnor_4 g22657(.A(new_n17833), .B(new_n17830), .Y(po1486));
  xnor_4 g22658(.A(new_n8270), .B(new_n8269), .Y(po1487));
  xor_4  g22659(.A(new_n23010), .B(new_n22995), .Y(po1488));
  xnor_4 g22660(.A(new_n13041), .B(new_n13012), .Y(po1490));
  xnor_4 g22661(.A(new_n16174), .B(new_n16162), .Y(po1491));
  xnor_4 g22662(.A(new_n14904), .B(new_n14903), .Y(po1492));
  xor_4  g22663(.A(new_n21725), .B(new_n22073), .Y(po1493));
  xor_4  g22664(.A(new_n10631), .B(new_n10629), .Y(po1494));
  xor_4  g22665(.A(new_n19994), .B(new_n19933), .Y(po1495));
  not_8  g22666(.A(new_n4984), .Y(new_n25015));
  xnor_4 g22667(.A(new_n4980), .B(new_n4733), .Y(new_n25016));
  nor_5  g22668(.A(new_n25016), .B(new_n25015), .Y(new_n25017));
  nand_5 g22669(.A(new_n25016), .B(new_n4994), .Y(new_n25018));
  nand_5 g22670(.A(new_n25018), .B(new_n4999), .Y(new_n25019));
  nor_5  g22671(.A(new_n25019), .B(new_n25017), .Y(new_n25020));
  not_8  g22672(.A(new_n4993), .Y(new_n25021));
  nand_5 g22673(.A(new_n4998), .B(new_n25021), .Y(new_n25022));
  nand_5 g22674(.A(new_n25022), .B(new_n5000), .Y(new_n25023));
  nor_5  g22675(.A(new_n25023), .B(new_n25020), .Y(po1496));
  nand_5 g22676(.A(new_n22738), .B(new_n22700), .Y(new_n25025));
  xor_4  g22677(.A(new_n25025), .B(new_n22737), .Y(po1497));
  xnor_4 g22678(.A(new_n17724), .B(new_n17723), .Y(po1498));
  xnor_4 g22679(.A(new_n15807), .B(new_n15748), .Y(po1499));
  xor_4  g22680(.A(new_n4207), .B(new_n4206), .Y(po1500));
  xor_4  g22681(.A(new_n14599), .B(new_n14581), .Y(po1501));
  xor_4  g22682(.A(new_n13996), .B(new_n12950), .Y(po1502));
  or_6   g22683(.A(new_n23013), .B(new_n22521), .Y(new_n25032));
  xor_4  g22684(.A(new_n25032), .B(new_n23022), .Y(po1503));
  xor_4  g22685(.A(new_n16567), .B(new_n16559), .Y(po1504));
  or_6   g22686(.A(new_n17022), .B(new_n17105), .Y(new_n25035));
  nand_5 g22687(.A(new_n22378), .B(new_n22377), .Y(new_n25036));
  nand_5 g22688(.A(new_n25036), .B(new_n25035), .Y(po1505));
  xor_4  g22689(.A(new_n21961), .B(new_n16316), .Y(po1506));
  nand_5 g22690(.A(new_n21684), .B(new_n21673), .Y(new_n25039));
  nor_5  g22691(.A(new_n25039), .B(new_n24221), .Y(new_n25040));
  nor_5  g22692(.A(new_n25040), .B(new_n24223), .Y(po1507));
endmodule


