// Benchmark "top_810222779_843330999_776144567_776418743_1234615" written by ABC on Sun Aug 18 19:24:06 2024

module top_810222779_843330999_776144567_776418743_1234615 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107;
  wire new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1306, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1330,
    new_n1331, new_n1332;
  nand_5     g0000(.A(pi123), .B(pi000), .Y(new_n316));
  nand_5 g0001(.A(pi054), .B(pi054), .Y(new_n317));
  nand_5     g0002(.A(pi150), .B(new_n317), .Y(new_n318));
  nand_5     g0003(.A(new_n318), .B(new_n316), .Y(new_n319));
  nand_5     g0004(.A(new_n319), .B(pi050), .Y(new_n320));
  nand_5 g0005(.A(pi115), .B(pi115), .Y(new_n321));
  nand_5     g0006(.A(pi150), .B(new_n321), .Y(new_n322));
  nand_5     g0007(.A(new_n322), .B(new_n316), .Y(new_n323));
  nand_5     g0008(.A(new_n323), .B(pi056), .Y(new_n324));
  nand_5 g0009(.A(new_n324), .B(new_n324), .Y(new_n325));
  nand_5 g0010(.A(pi056), .B(pi056), .Y(new_n326));
  xor_4      g0011(.A(new_n323), .B(new_n326), .Y(new_n327));
  nand_5 g0012(.A(pi150), .B(pi150), .Y(new_n328));
  or_6       g0013(.A(pi154), .B(new_n328), .Y(new_n329));
  nand_5     g0014(.A(new_n329), .B(new_n316), .Y(new_n330));
  or_6       g0015(.A(new_n330), .B(pi122), .Y(new_n331));
  xor_4      g0016(.A(new_n330), .B(pi122), .Y(new_n332));
  or_6       g0017(.A(pi175), .B(new_n328), .Y(new_n333));
  nand_5     g0018(.A(new_n333), .B(new_n316), .Y(new_n334));
  or_6       g0019(.A(new_n334), .B(pi047), .Y(new_n335));
  xor_4      g0020(.A(new_n334), .B(pi047), .Y(new_n336));
  nand_5 g0021(.A(pi196), .B(pi196), .Y(new_n337));
  nand_5 g0022(.A(pi186), .B(pi186), .Y(new_n338));
  nand_5     g0023(.A(new_n338), .B(new_n328), .Y(new_n339));
  nand_5 g0024(.A(new_n339), .B(new_n339), .Y(new_n340));
  nor_5      g0025(.A(pi182), .B(new_n328), .Y(new_n341));
  nor_5      g0026(.A(new_n341), .B(new_n340), .Y(new_n342));
  nor_5      g0027(.A(new_n342), .B(new_n337), .Y(new_n343));
  and_6      g0028(.A(new_n342), .B(new_n337), .Y(new_n344));
  nand_5 g0029(.A(pi199), .B(pi199), .Y(new_n345));
  nand_5     g0030(.A(pi150), .B(pi009), .Y(new_n346));
  nand_5     g0031(.A(pi177), .B(new_n328), .Y(new_n347));
  nand_5     g0032(.A(new_n347), .B(new_n346), .Y(new_n348));
  nand_5     g0033(.A(new_n348), .B(new_n345), .Y(new_n349));
  xor_4      g0034(.A(new_n348), .B(new_n345), .Y(new_n350));
  nand_5 g0035(.A(pi178), .B(pi178), .Y(new_n351));
  nand_5     g0036(.A(pi150), .B(pi080), .Y(new_n352));
  nand_5     g0037(.A(pi203), .B(new_n328), .Y(new_n353));
  nand_5     g0038(.A(new_n353), .B(new_n352), .Y(new_n354));
  nand_5     g0039(.A(new_n354), .B(new_n351), .Y(new_n355));
  or_6       g0040(.A(new_n354), .B(new_n351), .Y(new_n356));
  nand_5 g0041(.A(pi162), .B(pi162), .Y(new_n357));
  nand_5     g0042(.A(pi151), .B(new_n328), .Y(new_n358));
  nand_5     g0043(.A(pi172), .B(pi150), .Y(new_n359));
  nand_5     g0044(.A(new_n359), .B(new_n358), .Y(new_n360));
  nand_5     g0045(.A(new_n360), .B(new_n357), .Y(new_n361));
  nand_5 g0046(.A(new_n361), .B(new_n361), .Y(new_n362));
  nand_5 g0047(.A(pi160), .B(pi160), .Y(new_n363));
  nand_5     g0048(.A(new_n328), .B(pi034), .Y(new_n364));
  nand_5     g0049(.A(pi164), .B(pi150), .Y(new_n365));
  nand_5     g0050(.A(new_n365), .B(new_n364), .Y(new_n366));
  nand_5     g0051(.A(new_n366), .B(new_n363), .Y(new_n367));
  nand_5 g0052(.A(new_n367), .B(new_n367), .Y(new_n368));
  nand_5 g0053(.A(pi192), .B(pi192), .Y(new_n369));
  nand_5     g0054(.A(new_n328), .B(pi139), .Y(new_n370));
  nand_5     g0055(.A(pi150), .B(pi090), .Y(new_n371));
  nand_5     g0056(.A(new_n371), .B(new_n370), .Y(new_n372));
  or_6       g0057(.A(new_n372), .B(new_n369), .Y(new_n373));
  xor_4      g0058(.A(new_n372), .B(new_n369), .Y(new_n374));
  nand_5 g0059(.A(pi116), .B(pi116), .Y(new_n375));
  nand_5     g0060(.A(pi158), .B(pi150), .Y(new_n376));
  nand_5     g0061(.A(new_n328), .B(pi146), .Y(new_n377));
  nand_5     g0062(.A(new_n377), .B(new_n376), .Y(new_n378));
  or_6       g0063(.A(new_n378), .B(new_n375), .Y(new_n379));
  nand_5     g0064(.A(new_n378), .B(new_n375), .Y(new_n380));
  nand_5 g0065(.A(pi039), .B(pi039), .Y(new_n381));
  nand_5     g0066(.A(new_n328), .B(pi086), .Y(new_n382));
  nand_5     g0067(.A(pi150), .B(pi030), .Y(new_n383));
  nand_5     g0068(.A(new_n383), .B(new_n382), .Y(new_n384));
  nand_5     g0069(.A(new_n384), .B(new_n381), .Y(new_n385));
  nand_5 g0070(.A(new_n385), .B(new_n385), .Y(new_n386));
  nand_5 g0071(.A(pi057), .B(pi057), .Y(new_n387));
  nand_5     g0072(.A(new_n328), .B(pi142), .Y(new_n388));
  nand_5     g0073(.A(pi150), .B(pi032), .Y(new_n389));
  nand_5     g0074(.A(new_n389), .B(new_n388), .Y(new_n390));
  or_6       g0075(.A(new_n390), .B(new_n387), .Y(new_n391));
  nand_5 g0076(.A(pi107), .B(pi107), .Y(new_n392));
  nand_5     g0077(.A(pi189), .B(new_n328), .Y(new_n393));
  nand_5     g0078(.A(pi150), .B(pi106), .Y(new_n394));
  nand_5     g0079(.A(new_n394), .B(new_n393), .Y(new_n395));
  or_6       g0080(.A(new_n395), .B(new_n392), .Y(new_n396));
  xor_4      g0081(.A(new_n395), .B(new_n392), .Y(new_n397));
  nand_5     g0082(.A(pi194), .B(pi150), .Y(new_n398));
  nand_5     g0083(.A(pi156), .B(new_n328), .Y(new_n399));
  nand_5     g0084(.A(new_n399), .B(new_n398), .Y(new_n400));
  nand_5 g0085(.A(new_n400), .B(new_n400), .Y(new_n401));
  nand_5     g0086(.A(new_n401), .B(pi020), .Y(new_n402));
  nand_5 g0087(.A(pi020), .B(pi020), .Y(new_n403));
  nand_5     g0088(.A(new_n400), .B(new_n403), .Y(new_n404));
  nand_5 g0089(.A(pi170), .B(pi170), .Y(new_n405));
  nand_5     g0090(.A(pi150), .B(pi012), .Y(new_n406));
  nand_5     g0091(.A(new_n328), .B(pi131), .Y(new_n407));
  nand_5     g0092(.A(new_n407), .B(new_n406), .Y(new_n408));
  or_6       g0093(.A(new_n408), .B(new_n405), .Y(new_n409));
  xor_4      g0094(.A(new_n408), .B(new_n405), .Y(new_n410));
  nand_5 g0095(.A(pi051), .B(pi051), .Y(new_n411));
  nand_5     g0096(.A(pi150), .B(pi087), .Y(new_n412));
  nand_5     g0097(.A(new_n328), .B(pi014), .Y(new_n413));
  nand_5     g0098(.A(new_n413), .B(new_n412), .Y(new_n414));
  or_6       g0099(.A(new_n414), .B(new_n411), .Y(new_n415));
  nand_5 g0100(.A(pi074), .B(pi074), .Y(new_n416));
  nand_5 g0101(.A(pi180), .B(pi180), .Y(new_n417));
  nand_5     g0102(.A(pi169), .B(pi150), .Y(new_n418));
  nand_5     g0103(.A(new_n328), .B(pi033), .Y(new_n419));
  nand_5     g0104(.A(new_n419), .B(new_n418), .Y(new_n420));
  nand_5     g0105(.A(new_n420), .B(new_n417), .Y(new_n421));
  nand_5 g0106(.A(pi027), .B(pi027), .Y(new_n422));
  nand_5     g0107(.A(new_n328), .B(pi042), .Y(new_n423));
  nand_5     g0108(.A(pi150), .B(pi044), .Y(new_n424));
  nand_5     g0109(.A(new_n424), .B(new_n423), .Y(new_n425));
  nand_5     g0110(.A(new_n425), .B(new_n422), .Y(new_n426));
  nand_5 g0111(.A(pi083), .B(pi083), .Y(new_n427));
  nand_5     g0112(.A(new_n328), .B(pi007), .Y(new_n428));
  nand_5     g0113(.A(pi197), .B(pi150), .Y(new_n429));
  nand_5     g0114(.A(new_n429), .B(new_n428), .Y(new_n430));
  nand_5     g0115(.A(new_n430), .B(new_n427), .Y(new_n431));
  nand_5 g0116(.A(pi132), .B(pi132), .Y(new_n432));
  nand_5     g0117(.A(new_n328), .B(pi143), .Y(new_n433));
  nand_5     g0118(.A(pi150), .B(pi043), .Y(new_n434));
  nand_5     g0119(.A(new_n434), .B(new_n433), .Y(new_n435));
  nand_5     g0120(.A(new_n435), .B(new_n432), .Y(new_n436));
  xor_4      g0121(.A(new_n435), .B(new_n432), .Y(new_n437));
  nand_5 g0122(.A(pi004), .B(pi004), .Y(new_n438));
  nand_5     g0123(.A(new_n328), .B(pi058), .Y(new_n439));
  nand_5     g0124(.A(pi150), .B(pi025), .Y(new_n440));
  nand_5     g0125(.A(new_n440), .B(new_n439), .Y(new_n441));
  nand_5     g0126(.A(new_n441), .B(new_n438), .Y(new_n442));
  or_6       g0127(.A(new_n441), .B(new_n438), .Y(new_n443));
  nand_5     g0128(.A(new_n443), .B(new_n442), .Y(new_n444));
  nand_5 g0129(.A(pi092), .B(pi092), .Y(new_n445));
  nand_5     g0130(.A(pi193), .B(pi150), .Y(new_n446));
  nand_5     g0131(.A(pi152), .B(new_n328), .Y(new_n447));
  nand_5     g0132(.A(new_n447), .B(new_n446), .Y(new_n448));
  nand_5     g0133(.A(new_n448), .B(new_n445), .Y(new_n449));
  nand_5 g0134(.A(new_n449), .B(new_n449), .Y(new_n450));
  nand_5 g0135(.A(pi069), .B(pi069), .Y(new_n451));
  nand_5 g0136(.A(pi147), .B(pi147), .Y(new_n452));
  nand_5     g0137(.A(new_n452), .B(new_n451), .Y(new_n453));
  nand_5     g0138(.A(pi147), .B(pi069), .Y(new_n454));
  nand_5     g0139(.A(new_n454), .B(new_n328), .Y(new_n455));
  nand_5 g0140(.A(new_n455), .B(new_n455), .Y(new_n456));
  nand_5     g0141(.A(new_n456), .B(new_n453), .Y(new_n457));
  nand_5     g0142(.A(new_n457), .B(pi070), .Y(new_n458));
  nand_5     g0143(.A(new_n456), .B(pi069), .Y(new_n459));
  nand_5     g0144(.A(new_n459), .B(new_n458), .Y(new_n460));
  nand_5 g0145(.A(new_n460), .B(new_n460), .Y(new_n461));
  xor_4      g0146(.A(new_n448), .B(pi092), .Y(new_n462));
  nor_5      g0147(.A(new_n462), .B(new_n461), .Y(new_n463));
  nor_5      g0148(.A(new_n463), .B(new_n450), .Y(new_n464));
  or_6       g0149(.A(new_n464), .B(new_n444), .Y(new_n465));
  nand_5     g0150(.A(new_n465), .B(new_n442), .Y(new_n466));
  nand_5     g0151(.A(new_n466), .B(new_n437), .Y(new_n467));
  nand_5     g0152(.A(new_n467), .B(new_n436), .Y(new_n468));
  xor_4      g0153(.A(new_n430), .B(pi083), .Y(new_n469));
  nand_5 g0154(.A(new_n469), .B(new_n469), .Y(new_n470));
  nand_5     g0155(.A(new_n470), .B(new_n468), .Y(new_n471));
  nand_5     g0156(.A(new_n471), .B(new_n431), .Y(new_n472));
  nand_5 g0157(.A(new_n472), .B(new_n472), .Y(new_n473));
  xor_4      g0158(.A(new_n425), .B(pi027), .Y(new_n474));
  or_6       g0159(.A(new_n474), .B(new_n473), .Y(new_n475));
  nand_5     g0160(.A(new_n475), .B(new_n426), .Y(new_n476));
  xor_4      g0161(.A(new_n420), .B(new_n417), .Y(new_n477));
  nand_5     g0162(.A(new_n477), .B(new_n476), .Y(new_n478));
  nand_5     g0163(.A(new_n478), .B(new_n421), .Y(new_n479));
  or_6       g0164(.A(new_n479), .B(new_n416), .Y(new_n480));
  nand_5     g0165(.A(new_n328), .B(pi081), .Y(new_n481));
  nand_5     g0166(.A(pi150), .B(pi035), .Y(new_n482));
  nand_5     g0167(.A(new_n482), .B(new_n481), .Y(new_n483));
  nand_5     g0168(.A(new_n479), .B(new_n416), .Y(new_n484));
  nand_5     g0169(.A(new_n484), .B(new_n480), .Y(new_n485));
  or_6       g0170(.A(new_n485), .B(new_n483), .Y(new_n486));
  nand_5     g0171(.A(new_n486), .B(new_n480), .Y(new_n487));
  xor_4      g0172(.A(new_n414), .B(new_n411), .Y(new_n488));
  nand_5     g0173(.A(new_n488), .B(new_n487), .Y(new_n489));
  nand_5     g0174(.A(new_n489), .B(new_n415), .Y(new_n490));
  nand_5     g0175(.A(new_n490), .B(new_n410), .Y(new_n491));
  nand_5     g0176(.A(new_n491), .B(new_n409), .Y(new_n492));
  nand_5     g0177(.A(new_n492), .B(new_n404), .Y(new_n493));
  nand_5     g0178(.A(new_n493), .B(new_n402), .Y(new_n494));
  nand_5     g0179(.A(new_n494), .B(new_n397), .Y(new_n495));
  nand_5     g0180(.A(new_n495), .B(new_n396), .Y(new_n496));
  nand_5     g0181(.A(new_n496), .B(pi183), .Y(new_n497));
  or_6       g0182(.A(new_n496), .B(pi183), .Y(new_n498));
  nand_5     g0183(.A(new_n498), .B(new_n497), .Y(new_n499));
  nand_5     g0184(.A(pi187), .B(pi150), .Y(new_n500));
  nand_5     g0185(.A(new_n328), .B(pi094), .Y(new_n501));
  nand_5     g0186(.A(new_n501), .B(new_n500), .Y(new_n502));
  or_6       g0187(.A(new_n502), .B(new_n499), .Y(new_n503));
  nand_5     g0188(.A(new_n503), .B(new_n497), .Y(new_n504));
  xor_4      g0189(.A(new_n390), .B(new_n387), .Y(new_n505));
  nand_5     g0190(.A(new_n505), .B(new_n504), .Y(new_n506));
  nand_5     g0191(.A(new_n506), .B(new_n391), .Y(new_n507));
  xor_4      g0192(.A(new_n384), .B(pi039), .Y(new_n508));
  nor_5      g0193(.A(new_n508), .B(new_n507), .Y(new_n509));
  nor_5      g0194(.A(new_n509), .B(new_n386), .Y(new_n510));
  nand_5     g0195(.A(new_n510), .B(new_n380), .Y(new_n511));
  nand_5     g0196(.A(new_n511), .B(new_n379), .Y(new_n512));
  nand_5     g0197(.A(new_n512), .B(new_n374), .Y(new_n513));
  nand_5     g0198(.A(new_n513), .B(new_n373), .Y(new_n514));
  xor_4      g0199(.A(new_n366), .B(pi160), .Y(new_n515));
  nor_5      g0200(.A(new_n515), .B(new_n514), .Y(new_n516));
  nor_5      g0201(.A(new_n516), .B(new_n368), .Y(new_n517));
  xor_4      g0202(.A(new_n360), .B(pi162), .Y(new_n518));
  nor_5      g0203(.A(new_n518), .B(new_n517), .Y(new_n519));
  nor_5      g0204(.A(new_n519), .B(new_n362), .Y(new_n520));
  nand_5 g0205(.A(new_n520), .B(new_n520), .Y(new_n521));
  nand_5     g0206(.A(new_n521), .B(new_n356), .Y(new_n522));
  nand_5     g0207(.A(new_n522), .B(new_n355), .Y(new_n523));
  nand_5     g0208(.A(new_n523), .B(new_n350), .Y(new_n524));
  nand_5     g0209(.A(new_n524), .B(new_n349), .Y(new_n525));
  nor_5      g0210(.A(new_n525), .B(new_n344), .Y(new_n526));
  nor_5      g0211(.A(new_n526), .B(new_n343), .Y(new_n527));
  nand_5     g0212(.A(new_n527), .B(new_n336), .Y(new_n528));
  nand_5     g0213(.A(new_n528), .B(new_n335), .Y(new_n529));
  nand_5     g0214(.A(new_n529), .B(new_n332), .Y(new_n530));
  nand_5     g0215(.A(new_n530), .B(new_n331), .Y(new_n531));
  nor_5      g0216(.A(new_n531), .B(new_n327), .Y(new_n532));
  nor_5      g0217(.A(new_n532), .B(new_n325), .Y(new_n533));
  or_6       g0218(.A(new_n319), .B(pi050), .Y(new_n534));
  nand_5     g0219(.A(new_n534), .B(new_n320), .Y(new_n535));
  or_6       g0220(.A(new_n535), .B(new_n533), .Y(new_n536));
  and_6      g0221(.A(new_n536), .B(new_n320), .Y(new_n537));
  nand_5 g0222(.A(pi153), .B(pi153), .Y(new_n538));
  or_6       g0223(.A(new_n328), .B(pi026), .Y(new_n539));
  nand_5     g0224(.A(new_n539), .B(new_n316), .Y(new_n540));
  xor_4      g0225(.A(new_n540), .B(new_n538), .Y(new_n541));
  xnor_4     g0226(.A(new_n541), .B(new_n537), .Y(po000));
  nand_5 g0227(.A(pi165), .B(pi165), .Y(new_n543));
  nand_5     g0228(.A(pi167), .B(new_n543), .Y(po003));
  xor_4      g0229(.A(new_n508), .B(new_n507), .Y(po005));
  nand_5     g0230(.A(pi075), .B(pi037), .Y(new_n546));
  nand_5     g0231(.A(pi198), .B(pi188), .Y(new_n547));
  nor_5      g0232(.A(new_n547), .B(new_n546), .Y(new_n548));
  nand_5 g0233(.A(new_n548), .B(new_n548), .Y(po006));
  nand_5 g0234(.A(new_n316), .B(new_n316), .Y(new_n550));
  nor_5      g0235(.A(new_n328), .B(pi028), .Y(new_n551));
  nor_5      g0236(.A(new_n551), .B(new_n550), .Y(new_n552));
  nand_5 g0237(.A(pi041), .B(pi041), .Y(new_n553));
  nand_5     g0238(.A(new_n328), .B(new_n553), .Y(new_n554));
  nand_5 g0239(.A(new_n554), .B(new_n554), .Y(new_n555));
  nand_5 g0240(.A(pi181), .B(pi181), .Y(new_n556));
  nor_5      g0241(.A(new_n556), .B(new_n328), .Y(new_n557));
  nor_5      g0242(.A(new_n557), .B(new_n555), .Y(new_n558));
  nor_5      g0243(.A(new_n558), .B(new_n552), .Y(new_n559));
  nand_5     g0244(.A(pi203), .B(pi140), .Y(new_n560));
  nand_5     g0245(.A(pi186), .B(pi161), .Y(new_n561));
  nand_5 g0246(.A(new_n561), .B(new_n561), .Y(new_n562));
  nand_5     g0247(.A(pi177), .B(pi173), .Y(new_n563));
  nand_5     g0248(.A(new_n563), .B(new_n328), .Y(new_n564));
  nor_5      g0249(.A(new_n564), .B(new_n562), .Y(new_n565));
  and_6      g0250(.A(new_n565), .B(new_n560), .Y(new_n566));
  nand_5     g0251(.A(new_n316), .B(pi110), .Y(new_n567));
  or_6       g0252(.A(new_n567), .B(pi047), .Y(new_n568));
  nand_5 g0253(.A(pi119), .B(pi119), .Y(new_n569));
  nor_5      g0254(.A(pi196), .B(new_n569), .Y(new_n570));
  nor_5      g0255(.A(new_n570), .B(new_n328), .Y(new_n571));
  nand_5     g0256(.A(new_n571), .B(new_n568), .Y(new_n572));
  nand_5     g0257(.A(new_n351), .B(pi174), .Y(new_n573));
  nand_5     g0258(.A(new_n345), .B(pi006), .Y(new_n574));
  nand_5     g0259(.A(new_n574), .B(new_n573), .Y(new_n575));
  nor_5      g0260(.A(new_n575), .B(new_n572), .Y(new_n576));
  nor_5      g0261(.A(new_n576), .B(new_n566), .Y(new_n577));
  nand_5 g0262(.A(pi055), .B(pi055), .Y(new_n578));
  nor_5      g0263(.A(pi083), .B(new_n578), .Y(new_n579));
  nor_5      g0264(.A(new_n432), .B(pi089), .Y(new_n580));
  nand_5     g0265(.A(pi103), .B(pi091), .Y(new_n581));
  nand_5     g0266(.A(new_n581), .B(pi092), .Y(new_n582));
  nand_5 g0267(.A(pi091), .B(pi091), .Y(new_n583));
  nand_5 g0268(.A(pi103), .B(pi103), .Y(new_n584));
  nand_5     g0269(.A(new_n584), .B(new_n583), .Y(new_n585));
  nand_5     g0270(.A(new_n585), .B(new_n582), .Y(new_n586));
  nor_5      g0271(.A(new_n438), .B(pi002), .Y(new_n587));
  nor_5      g0272(.A(new_n587), .B(new_n586), .Y(new_n588));
  nand_5     g0273(.A(new_n438), .B(pi002), .Y(new_n589));
  nand_5     g0274(.A(new_n432), .B(pi089), .Y(new_n590));
  nand_5     g0275(.A(new_n590), .B(new_n589), .Y(new_n591));
  nor_5      g0276(.A(new_n591), .B(new_n588), .Y(new_n592));
  nor_5      g0277(.A(new_n592), .B(new_n580), .Y(new_n593));
  nor_5      g0278(.A(new_n593), .B(new_n579), .Y(new_n594));
  or_6       g0279(.A(pi067), .B(new_n422), .Y(new_n595));
  nand_5     g0280(.A(pi083), .B(new_n578), .Y(new_n596));
  nand_5     g0281(.A(new_n596), .B(new_n595), .Y(new_n597));
  nor_5      g0282(.A(new_n597), .B(new_n594), .Y(new_n598));
  nand_5     g0283(.A(new_n417), .B(pi059), .Y(new_n599));
  nand_5     g0284(.A(pi067), .B(new_n422), .Y(new_n600));
  nand_5     g0285(.A(new_n600), .B(new_n599), .Y(new_n601));
  nor_5      g0286(.A(new_n601), .B(new_n598), .Y(new_n602));
  nand_5 g0287(.A(pi059), .B(pi059), .Y(new_n603));
  nand_5     g0288(.A(pi180), .B(new_n603), .Y(new_n604));
  or_6       g0289(.A(new_n416), .B(pi038), .Y(new_n605));
  nand_5     g0290(.A(new_n605), .B(new_n604), .Y(new_n606));
  nor_5      g0291(.A(new_n606), .B(new_n602), .Y(new_n607));
  nand_5     g0292(.A(new_n416), .B(pi038), .Y(new_n608));
  nand_5     g0293(.A(pi206), .B(new_n411), .Y(new_n609));
  nand_5     g0294(.A(new_n609), .B(new_n608), .Y(new_n610));
  nor_5      g0295(.A(new_n610), .B(new_n607), .Y(new_n611));
  nand_5 g0296(.A(pi049), .B(pi049), .Y(new_n612));
  nand_5     g0297(.A(pi170), .B(new_n612), .Y(new_n613));
  or_6       g0298(.A(pi206), .B(new_n411), .Y(new_n614));
  nand_5     g0299(.A(new_n614), .B(new_n613), .Y(new_n615));
  nor_5      g0300(.A(new_n615), .B(new_n611), .Y(new_n616));
  nand_5     g0301(.A(pi135), .B(new_n403), .Y(new_n617));
  nand_5     g0302(.A(new_n405), .B(pi049), .Y(new_n618));
  nand_5     g0303(.A(new_n618), .B(new_n617), .Y(new_n619));
  nor_5      g0304(.A(new_n619), .B(new_n616), .Y(new_n620));
  nor_5      g0305(.A(pi135), .B(new_n403), .Y(new_n621));
  nor_5      g0306(.A(new_n392), .B(pi011), .Y(new_n622));
  or_6       g0307(.A(new_n622), .B(new_n621), .Y(new_n623));
  nor_5      g0308(.A(new_n623), .B(new_n620), .Y(new_n624));
  nand_5 g0309(.A(pi195), .B(pi195), .Y(new_n625));
  or_6       g0310(.A(new_n625), .B(pi183), .Y(new_n626));
  nand_5     g0311(.A(new_n392), .B(pi011), .Y(new_n627));
  nand_5     g0312(.A(new_n627), .B(new_n626), .Y(new_n628));
  nor_5      g0313(.A(new_n628), .B(new_n624), .Y(new_n629));
  nand_5     g0314(.A(new_n625), .B(pi183), .Y(new_n630));
  or_6       g0315(.A(pi097), .B(new_n387), .Y(new_n631));
  nand_5     g0316(.A(new_n631), .B(new_n630), .Y(new_n632));
  nor_5      g0317(.A(new_n632), .B(new_n629), .Y(new_n633));
  nand_5     g0318(.A(new_n381), .B(pi005), .Y(new_n634));
  nand_5     g0319(.A(pi097), .B(new_n387), .Y(new_n635));
  nand_5     g0320(.A(new_n635), .B(new_n634), .Y(new_n636));
  nor_5      g0321(.A(new_n636), .B(new_n633), .Y(new_n637));
  nor_5      g0322(.A(new_n375), .B(pi114), .Y(new_n638));
  nor_5      g0323(.A(new_n381), .B(pi005), .Y(new_n639));
  or_6       g0324(.A(new_n639), .B(new_n638), .Y(new_n640));
  nor_5      g0325(.A(new_n640), .B(new_n637), .Y(new_n641));
  nand_5     g0326(.A(new_n369), .B(pi036), .Y(new_n642));
  nand_5     g0327(.A(new_n375), .B(pi114), .Y(new_n643));
  nand_5     g0328(.A(new_n643), .B(new_n642), .Y(new_n644));
  nor_5      g0329(.A(new_n644), .B(new_n641), .Y(new_n645));
  nor_5      g0330(.A(new_n369), .B(pi036), .Y(new_n646));
  nor_5      g0331(.A(new_n363), .B(pi052), .Y(new_n647));
  or_6       g0332(.A(new_n647), .B(new_n646), .Y(new_n648));
  nor_5      g0333(.A(new_n648), .B(new_n645), .Y(new_n649));
  nand_5     g0334(.A(new_n363), .B(pi052), .Y(new_n650));
  nand_5     g0335(.A(new_n650), .B(pi150), .Y(new_n651));
  nor_5      g0336(.A(new_n651), .B(new_n649), .Y(new_n652));
  or_6       g0337(.A(pi142), .B(pi138), .Y(new_n653));
  nand_5 g0338(.A(pi081), .B(pi081), .Y(new_n654));
  nand_5 g0339(.A(pi117), .B(pi117), .Y(new_n655));
  nor_5      g0340(.A(new_n655), .B(new_n654), .Y(new_n656));
  nor_5      g0341(.A(pi033), .B(pi023), .Y(new_n657));
  nor_5      g0342(.A(new_n583), .B(new_n451), .Y(new_n658));
  nor_5      g0343(.A(new_n658), .B(pi096), .Y(new_n659));
  or_6       g0344(.A(pi152), .B(pi066), .Y(new_n660));
  nand_5     g0345(.A(new_n583), .B(new_n451), .Y(new_n661));
  nand_5     g0346(.A(new_n661), .B(new_n660), .Y(new_n662));
  nor_5      g0347(.A(new_n662), .B(new_n659), .Y(new_n663));
  nand_5     g0348(.A(pi152), .B(pi066), .Y(new_n664));
  nand_5     g0349(.A(pi111), .B(pi058), .Y(new_n665));
  nand_5     g0350(.A(new_n665), .B(new_n664), .Y(new_n666));
  nor_5      g0351(.A(new_n666), .B(new_n663), .Y(new_n667));
  nor_5      g0352(.A(pi111), .B(pi058), .Y(new_n668));
  nor_5      g0353(.A(pi143), .B(pi048), .Y(new_n669));
  or_6       g0354(.A(new_n669), .B(new_n668), .Y(new_n670));
  nor_5      g0355(.A(new_n670), .B(new_n667), .Y(new_n671));
  nand_5     g0356(.A(pi143), .B(pi048), .Y(new_n672));
  nand_5     g0357(.A(pi098), .B(pi007), .Y(new_n673));
  nand_5     g0358(.A(new_n673), .B(new_n672), .Y(new_n674));
  nor_5      g0359(.A(new_n674), .B(new_n671), .Y(new_n675));
  nor_5      g0360(.A(pi098), .B(pi007), .Y(new_n676));
  nor_5      g0361(.A(pi042), .B(pi029), .Y(new_n677));
  or_6       g0362(.A(new_n677), .B(new_n676), .Y(new_n678));
  nor_5      g0363(.A(new_n678), .B(new_n675), .Y(new_n679));
  nand_5     g0364(.A(pi042), .B(pi029), .Y(new_n680));
  nand_5     g0365(.A(pi033), .B(pi023), .Y(new_n681));
  nand_5     g0366(.A(new_n681), .B(new_n680), .Y(new_n682));
  nor_5      g0367(.A(new_n682), .B(new_n679), .Y(new_n683));
  nor_5      g0368(.A(new_n683), .B(new_n657), .Y(new_n684));
  nor_5      g0369(.A(new_n684), .B(new_n656), .Y(new_n685));
  nand_5     g0370(.A(new_n655), .B(new_n654), .Y(new_n686));
  or_6       g0371(.A(pi100), .B(pi014), .Y(new_n687));
  nand_5     g0372(.A(new_n687), .B(new_n686), .Y(new_n688));
  nor_5      g0373(.A(new_n688), .B(new_n685), .Y(new_n689));
  nand_5     g0374(.A(pi149), .B(pi131), .Y(new_n690));
  nand_5     g0375(.A(pi100), .B(pi014), .Y(new_n691));
  nand_5     g0376(.A(new_n691), .B(new_n690), .Y(new_n692));
  nor_5      g0377(.A(new_n692), .B(new_n689), .Y(new_n693));
  nor_5      g0378(.A(pi149), .B(pi131), .Y(new_n694));
  nor_5      g0379(.A(pi201), .B(pi156), .Y(new_n695));
  or_6       g0380(.A(new_n695), .B(new_n694), .Y(new_n696));
  nor_5      g0381(.A(new_n696), .B(new_n693), .Y(new_n697));
  nand_5     g0382(.A(pi201), .B(pi156), .Y(new_n698));
  nand_5     g0383(.A(pi189), .B(pi113), .Y(new_n699));
  nand_5     g0384(.A(new_n699), .B(new_n698), .Y(new_n700));
  nor_5      g0385(.A(new_n700), .B(new_n697), .Y(new_n701));
  nor_5      g0386(.A(pi189), .B(pi113), .Y(new_n702));
  nor_5      g0387(.A(pi166), .B(pi094), .Y(new_n703));
  or_6       g0388(.A(new_n703), .B(new_n702), .Y(new_n704));
  or_6       g0389(.A(new_n704), .B(new_n701), .Y(new_n705));
  nand_5     g0390(.A(pi166), .B(pi094), .Y(new_n706));
  nand_5     g0391(.A(new_n706), .B(new_n705), .Y(new_n707));
  nand_5     g0392(.A(new_n707), .B(new_n653), .Y(new_n708));
  nand_5     g0393(.A(pi179), .B(pi086), .Y(new_n709));
  nand_5     g0394(.A(pi142), .B(pi138), .Y(new_n710));
  and_6      g0395(.A(new_n710), .B(new_n709), .Y(new_n711));
  nand_5     g0396(.A(new_n711), .B(new_n708), .Y(new_n712));
  nor_5      g0397(.A(pi146), .B(pi016), .Y(new_n713));
  nor_5      g0398(.A(pi179), .B(pi086), .Y(new_n714));
  nor_5      g0399(.A(new_n714), .B(new_n713), .Y(new_n715));
  and_6      g0400(.A(new_n715), .B(new_n712), .Y(new_n716));
  nand_5     g0401(.A(pi139), .B(pi068), .Y(new_n717));
  nand_5     g0402(.A(pi146), .B(pi016), .Y(new_n718));
  nand_5     g0403(.A(new_n718), .B(new_n717), .Y(new_n719));
  nor_5      g0404(.A(new_n719), .B(new_n716), .Y(new_n720));
  nor_5      g0405(.A(pi104), .B(pi034), .Y(new_n721));
  nor_5      g0406(.A(pi139), .B(pi068), .Y(new_n722));
  or_6       g0407(.A(new_n722), .B(new_n721), .Y(new_n723));
  nor_5      g0408(.A(new_n723), .B(new_n720), .Y(new_n724));
  nand_5     g0409(.A(pi104), .B(pi034), .Y(new_n725));
  nand_5     g0410(.A(new_n725), .B(new_n328), .Y(new_n726));
  nor_5      g0411(.A(new_n726), .B(new_n724), .Y(new_n727));
  nor_5      g0412(.A(new_n727), .B(new_n652), .Y(po084));
  nand_5 g0413(.A(pi082), .B(pi082), .Y(new_n729));
  nor_5      g0414(.A(new_n328), .B(new_n729), .Y(new_n730));
  nand_5     g0415(.A(new_n730), .B(new_n357), .Y(new_n731));
  nand_5 g0416(.A(pi121), .B(pi121), .Y(new_n732));
  or_6       g0417(.A(new_n358), .B(new_n732), .Y(new_n733));
  nand_5     g0418(.A(new_n733), .B(new_n731), .Y(new_n734));
  nor_5      g0419(.A(new_n734), .B(po084), .Y(new_n735));
  or_6       g0420(.A(new_n351), .B(pi174), .Y(new_n736));
  nand_5     g0421(.A(pi162), .B(new_n729), .Y(new_n737));
  nand_5     g0422(.A(new_n737), .B(new_n736), .Y(new_n738));
  nand_5     g0423(.A(new_n738), .B(pi150), .Y(new_n739));
  nand_5     g0424(.A(new_n328), .B(new_n732), .Y(new_n740));
  or_6       g0425(.A(new_n740), .B(pi151), .Y(new_n741));
  nand_5     g0426(.A(new_n741), .B(new_n739), .Y(new_n742));
  nor_5      g0427(.A(new_n742), .B(new_n735), .Y(new_n743));
  nor_5      g0428(.A(new_n743), .B(new_n577), .Y(new_n744));
  nor_5      g0429(.A(pi088), .B(pi073), .Y(new_n745));
  nor_5      g0430(.A(pi141), .B(pi112), .Y(new_n746));
  nand_5     g0431(.A(new_n746), .B(new_n745), .Y(new_n747));
  nor_5      g0432(.A(pi065), .B(pi003), .Y(new_n748));
  nand_5 g0433(.A(new_n748), .B(new_n748), .Y(new_n749));
  nor_5      g0434(.A(pi019), .B(pi010), .Y(new_n750));
  nand_5     g0435(.A(new_n750), .B(new_n555), .Y(new_n751));
  nor_5      g0436(.A(new_n751), .B(new_n749), .Y(new_n752));
  nand_5 g0437(.A(new_n752), .B(new_n752), .Y(new_n753));
  nor_5      g0438(.A(new_n753), .B(new_n747), .Y(new_n754));
  nand_5 g0439(.A(new_n754), .B(new_n754), .Y(new_n755));
  nand_5 g0440(.A(pi018), .B(pi018), .Y(new_n756));
  nand_5     g0441(.A(new_n326), .B(new_n756), .Y(new_n757));
  nor_5      g0442(.A(new_n757), .B(pi101), .Y(new_n758));
  nand_5 g0443(.A(pi085), .B(pi085), .Y(new_n759));
  nand_5 g0444(.A(pi204), .B(pi204), .Y(new_n760));
  nand_5     g0445(.A(new_n760), .B(new_n759), .Y(new_n761));
  nand_5 g0446(.A(pi050), .B(pi050), .Y(new_n762));
  nand_5     g0447(.A(new_n538), .B(new_n762), .Y(new_n763));
  nor_5      g0448(.A(new_n763), .B(new_n761), .Y(new_n764));
  nand_5     g0449(.A(new_n764), .B(new_n758), .Y(new_n765));
  nand_5 g0450(.A(pi101), .B(pi101), .Y(new_n766));
  nor_5      g0451(.A(pi159), .B(new_n766), .Y(new_n767));
  nor_5      g0452(.A(new_n756), .B(pi013), .Y(new_n768));
  nor_5      g0453(.A(new_n768), .B(new_n767), .Y(new_n769));
  nand_5 g0454(.A(pi095), .B(pi095), .Y(new_n770));
  nand_5     g0455(.A(pi153), .B(new_n770), .Y(new_n771));
  and_6      g0456(.A(new_n771), .B(new_n316), .Y(new_n772));
  nand_5     g0457(.A(new_n772), .B(new_n769), .Y(new_n773));
  nand_5     g0458(.A(new_n773), .B(new_n765), .Y(new_n774));
  nand_5 g0459(.A(pi185), .B(pi185), .Y(new_n775));
  nand_5     g0460(.A(new_n775), .B(pi085), .Y(new_n776));
  nand_5     g0461(.A(new_n776), .B(pi150), .Y(new_n777));
  nand_5 g0462(.A(pi015), .B(pi015), .Y(new_n778));
  nand_5     g0463(.A(pi050), .B(new_n778), .Y(new_n779));
  or_6       g0464(.A(pi105), .B(new_n326), .Y(new_n780));
  nand_5     g0465(.A(new_n780), .B(new_n779), .Y(new_n781));
  nor_5      g0466(.A(new_n781), .B(new_n777), .Y(new_n782));
  nand_5     g0467(.A(new_n782), .B(new_n774), .Y(new_n783));
  nand_5     g0468(.A(pi088), .B(pi019), .Y(new_n784));
  nand_5     g0469(.A(pi112), .B(pi073), .Y(new_n785));
  nor_5      g0470(.A(new_n785), .B(new_n784), .Y(new_n786));
  nand_5     g0471(.A(new_n328), .B(pi141), .Y(new_n787));
  nand_5     g0472(.A(pi065), .B(pi003), .Y(new_n788));
  nor_5      g0473(.A(new_n788), .B(new_n787), .Y(new_n789));
  nand_5     g0474(.A(new_n789), .B(new_n786), .Y(new_n790));
  nand_5     g0475(.A(new_n790), .B(new_n783), .Y(new_n791));
  nand_5 g0476(.A(pi122), .B(pi122), .Y(new_n792));
  nand_5 g0477(.A(pi047), .B(pi047), .Y(new_n793));
  nand_5     g0478(.A(pi150), .B(new_n793), .Y(new_n794));
  nand_5     g0479(.A(new_n794), .B(new_n567), .Y(new_n795));
  nand_5     g0480(.A(new_n795), .B(new_n792), .Y(new_n796));
  nand_5 g0481(.A(pi190), .B(pi190), .Y(new_n797));
  nand_5     g0482(.A(new_n328), .B(pi010), .Y(new_n798));
  nor_5      g0483(.A(new_n798), .B(new_n797), .Y(new_n799));
  nor_5      g0484(.A(pi110), .B(new_n793), .Y(new_n800));
  nand_5     g0485(.A(new_n316), .B(pi084), .Y(new_n801));
  nor_5      g0486(.A(new_n801), .B(new_n800), .Y(new_n802));
  nor_5      g0487(.A(new_n802), .B(new_n799), .Y(new_n803));
  nand_5     g0488(.A(new_n803), .B(new_n796), .Y(new_n804));
  nand_5     g0489(.A(new_n804), .B(new_n791), .Y(new_n805));
  nand_5     g0490(.A(new_n805), .B(new_n755), .Y(new_n806));
  nor_5      g0491(.A(new_n337), .B(pi119), .Y(new_n807));
  nor_5      g0492(.A(new_n345), .B(pi006), .Y(new_n808));
  nor_5      g0493(.A(new_n808), .B(new_n807), .Y(new_n809));
  nor_5      g0494(.A(new_n809), .B(new_n572), .Y(new_n810));
  or_6       g0495(.A(new_n339), .B(pi161), .Y(new_n811));
  nor_5      g0496(.A(pi177), .B(pi173), .Y(new_n812));
  nor_5      g0497(.A(pi203), .B(pi140), .Y(new_n813));
  or_6       g0498(.A(new_n813), .B(new_n812), .Y(new_n814));
  nand_5     g0499(.A(new_n814), .B(new_n565), .Y(new_n815));
  nand_5     g0500(.A(new_n815), .B(new_n811), .Y(new_n816));
  nor_5      g0501(.A(new_n816), .B(new_n810), .Y(new_n817));
  nand_5     g0502(.A(new_n817), .B(new_n806), .Y(new_n818));
  nor_5      g0503(.A(new_n818), .B(new_n744), .Y(new_n819));
  nand_5     g0504(.A(new_n754), .B(pi190), .Y(new_n820));
  nand_5     g0505(.A(new_n792), .B(pi084), .Y(new_n821));
  nand_5     g0506(.A(pi105), .B(new_n326), .Y(new_n822));
  nand_5     g0507(.A(new_n822), .B(new_n821), .Y(new_n823));
  nand_5     g0508(.A(new_n823), .B(new_n791), .Y(new_n824));
  nand_5     g0509(.A(pi159), .B(new_n766), .Y(new_n825));
  nor_5      g0510(.A(pi050), .B(new_n778), .Y(new_n826));
  nand_5     g0511(.A(new_n826), .B(new_n771), .Y(new_n827));
  nor_5      g0512(.A(pi153), .B(new_n770), .Y(new_n828));
  nand_5     g0513(.A(pi185), .B(new_n759), .Y(new_n829));
  nand_5     g0514(.A(new_n829), .B(pi204), .Y(new_n830));
  nor_5      g0515(.A(new_n830), .B(new_n828), .Y(new_n831));
  nand_5     g0516(.A(new_n831), .B(new_n827), .Y(new_n832));
  nand_5     g0517(.A(new_n832), .B(new_n776), .Y(new_n833));
  nand_5     g0518(.A(new_n833), .B(new_n825), .Y(new_n834));
  nand_5     g0519(.A(new_n834), .B(new_n769), .Y(new_n835));
  nand_5 g0520(.A(pi013), .B(pi013), .Y(new_n836));
  nor_5      g0521(.A(pi018), .B(new_n836), .Y(new_n837));
  nor_5      g0522(.A(new_n557), .B(new_n551), .Y(new_n838));
  nor_5      g0523(.A(new_n838), .B(new_n837), .Y(new_n839));
  nand_5     g0524(.A(new_n839), .B(new_n835), .Y(new_n840));
  nand_5     g0525(.A(new_n840), .B(new_n755), .Y(new_n841));
  nand_5     g0526(.A(new_n841), .B(new_n824), .Y(new_n842));
  nand_5     g0527(.A(new_n842), .B(new_n316), .Y(new_n843));
  nand_5     g0528(.A(new_n843), .B(new_n820), .Y(new_n844));
  nor_5      g0529(.A(new_n844), .B(new_n819), .Y(new_n845));
  nor_5      g0530(.A(new_n845), .B(new_n559), .Y(new_n846));
  nand_5 g0531(.A(pi124), .B(pi124), .Y(new_n847));
  nand_5 g0532(.A(pi022), .B(pi022), .Y(new_n848));
  nand_5 g0533(.A(pi071), .B(pi071), .Y(new_n849));
  nand_5 g0534(.A(pi078), .B(pi078), .Y(new_n850));
  nand_5     g0535(.A(new_n850), .B(new_n849), .Y(new_n851));
  nor_5      g0536(.A(new_n851), .B(new_n848), .Y(new_n852));
  nor_5      g0537(.A(new_n852), .B(new_n847), .Y(new_n853));
  nor_5      g0538(.A(new_n853), .B(new_n846), .Y(new_n854));
  nor_5      g0539(.A(new_n850), .B(new_n849), .Y(new_n855));
  nand_5     g0540(.A(new_n847), .B(pi022), .Y(new_n856));
  nor_5      g0541(.A(new_n856), .B(new_n855), .Y(new_n857));
  nor_5      g0542(.A(new_n857), .B(new_n854), .Y(po008));
  xor_4      g0543(.A(new_n527), .B(new_n336), .Y(po009));
  xor_4      g0544(.A(new_n529), .B(new_n332), .Y(po011));
  nand_5 g0545(.A(pi145), .B(pi145), .Y(new_n861));
  nand_5     g0546(.A(pi150), .B(new_n861), .Y(new_n862));
  nand_5     g0547(.A(new_n862), .B(new_n316), .Y(new_n863));
  nand_5     g0548(.A(new_n863), .B(pi085), .Y(new_n864));
  xor_4      g0549(.A(new_n863), .B(pi085), .Y(new_n865));
  nand_5     g0550(.A(new_n540), .B(pi153), .Y(new_n866));
  or_6       g0551(.A(new_n541), .B(new_n537), .Y(new_n867));
  nand_5     g0552(.A(new_n867), .B(new_n866), .Y(new_n868));
  nand_5     g0553(.A(new_n868), .B(pi204), .Y(new_n869));
  nor_5      g0554(.A(new_n328), .B(pi061), .Y(new_n870));
  nor_5      g0555(.A(new_n870), .B(new_n550), .Y(new_n871));
  xor_4      g0556(.A(new_n868), .B(new_n760), .Y(new_n872));
  or_6       g0557(.A(new_n872), .B(new_n871), .Y(new_n873));
  nand_5     g0558(.A(new_n873), .B(new_n869), .Y(new_n874));
  nand_5     g0559(.A(new_n874), .B(new_n865), .Y(new_n875));
  nand_5     g0560(.A(new_n875), .B(new_n864), .Y(new_n876));
  or_6       g0561(.A(new_n328), .B(pi062), .Y(new_n877));
  nand_5     g0562(.A(new_n877), .B(new_n316), .Y(new_n878));
  xor_4      g0563(.A(new_n878), .B(pi101), .Y(new_n879));
  xnor_4     g0564(.A(new_n879), .B(new_n876), .Y(po013));
  xor_4      g0565(.A(pi092), .B(new_n411), .Y(new_n881));
  xor_4      g0566(.A(pi180), .B(pi083), .Y(new_n882));
  xor_4      g0567(.A(new_n882), .B(pi132), .Y(new_n883));
  xor_4      g0568(.A(new_n883), .B(new_n881), .Y(new_n884));
  or_6       g0569(.A(new_n431), .B(new_n426), .Y(new_n885));
  nor_5      g0570(.A(new_n425), .B(new_n422), .Y(new_n886));
  nand_5     g0571(.A(new_n886), .B(new_n431), .Y(new_n887));
  nand_5     g0572(.A(new_n887), .B(new_n885), .Y(new_n888));
  or_6       g0573(.A(new_n888), .B(new_n468), .Y(new_n889));
  nor_5      g0574(.A(new_n430), .B(new_n427), .Y(new_n890));
  or_6       g0575(.A(new_n890), .B(new_n426), .Y(new_n891));
  nand_5     g0576(.A(new_n886), .B(new_n890), .Y(new_n892));
  nand_5     g0577(.A(new_n892), .B(new_n891), .Y(new_n893));
  nand_5     g0578(.A(new_n893), .B(new_n468), .Y(new_n894));
  nand_5     g0579(.A(new_n894), .B(new_n889), .Y(new_n895));
  xor_4      g0580(.A(pi043), .B(pi035), .Y(new_n896));
  xor_4      g0581(.A(pi197), .B(pi193), .Y(new_n897));
  xor_4      g0582(.A(pi169), .B(pi087), .Y(new_n898));
  xnor_4     g0583(.A(new_n898), .B(new_n897), .Y(new_n899));
  xor_4      g0584(.A(new_n899), .B(new_n896), .Y(new_n900));
  nand_5     g0585(.A(new_n900), .B(pi150), .Y(new_n901));
  xor_4      g0586(.A(new_n451), .B(pi033), .Y(new_n902));
  xor_4      g0587(.A(new_n902), .B(pi007), .Y(new_n903));
  xor_4      g0588(.A(pi143), .B(pi081), .Y(new_n904));
  xnor_4     g0589(.A(pi152), .B(pi014), .Y(new_n905));
  xor_4      g0590(.A(new_n905), .B(new_n904), .Y(new_n906));
  xor_4      g0591(.A(new_n906), .B(new_n903), .Y(new_n907));
  nand_5 g0592(.A(pi070), .B(pi070), .Y(new_n908));
  nand_5     g0593(.A(new_n453), .B(new_n908), .Y(new_n909));
  nand_5     g0594(.A(new_n909), .B(new_n454), .Y(new_n910));
  xnor_4     g0595(.A(new_n910), .B(new_n907), .Y(new_n911));
  nand_5     g0596(.A(new_n911), .B(new_n328), .Y(new_n912));
  nand_5     g0597(.A(new_n912), .B(new_n901), .Y(new_n913));
  xor_4      g0598(.A(new_n913), .B(new_n895), .Y(new_n914));
  xor_4      g0599(.A(new_n914), .B(new_n884), .Y(new_n915));
  nand_5     g0600(.A(new_n464), .B(new_n443), .Y(new_n916));
  nand_5 g0601(.A(new_n464), .B(new_n464), .Y(new_n917));
  nand_5     g0602(.A(new_n917), .B(new_n442), .Y(new_n918));
  nand_5     g0603(.A(new_n918), .B(new_n916), .Y(new_n919));
  nand_5     g0604(.A(new_n486), .B(new_n484), .Y(new_n920));
  xnor_4     g0605(.A(new_n920), .B(new_n919), .Y(new_n921));
  xor_4      g0606(.A(new_n921), .B(new_n915), .Y(po015));
  xnor_4     g0607(.A(new_n502), .B(new_n499), .Y(po016));
  nand_5 g0608(.A(pi125), .B(pi125), .Y(po017));
  and_6      g0609(.A(pi109), .B(pi060), .Y(po020));
  nand_5 g0610(.A(new_n533), .B(new_n533), .Y(new_n926));
  xor_4      g0611(.A(new_n535), .B(new_n926), .Y(po024));
  xnor_4     g0612(.A(new_n505), .B(new_n504), .Y(po025));
  or_6       g0613(.A(new_n328), .B(pi077), .Y(new_n929));
  nand_5     g0614(.A(new_n929), .B(new_n316), .Y(new_n930));
  and_6      g0615(.A(new_n930), .B(pi181), .Y(new_n931));
  nand_5     g0616(.A(new_n878), .B(pi101), .Y(new_n932));
  nand_5     g0617(.A(new_n879), .B(new_n876), .Y(new_n933));
  nand_5     g0618(.A(new_n933), .B(new_n932), .Y(new_n934));
  or_6       g0619(.A(new_n934), .B(pi018), .Y(new_n935));
  nor_5      g0620(.A(pi184), .B(new_n328), .Y(new_n936));
  nor_5      g0621(.A(new_n936), .B(new_n550), .Y(new_n937));
  nand_5     g0622(.A(new_n934), .B(pi018), .Y(new_n938));
  and_6      g0623(.A(new_n938), .B(new_n935), .Y(new_n939));
  nand_5     g0624(.A(new_n939), .B(new_n937), .Y(new_n940));
  nand_5     g0625(.A(new_n940), .B(new_n935), .Y(new_n941));
  xor_4      g0626(.A(new_n930), .B(new_n556), .Y(new_n942));
  nor_5      g0627(.A(new_n942), .B(new_n941), .Y(new_n943));
  nor_5      g0628(.A(new_n943), .B(new_n931), .Y(new_n944));
  nand_5     g0629(.A(new_n944), .B(new_n847), .Y(new_n945));
  or_6       g0630(.A(new_n944), .B(new_n847), .Y(new_n946));
  nand_5     g0631(.A(new_n946), .B(new_n945), .Y(new_n947));
  nand_5     g0632(.A(pi064), .B(pi022), .Y(new_n948));
  nor_5      g0633(.A(new_n948), .B(new_n947), .Y(new_n949));
  xor_4      g0634(.A(pi064), .B(pi024), .Y(new_n950));
  nand_5     g0635(.A(new_n950), .B(pi022), .Y(new_n951));
  nor_5      g0636(.A(new_n951), .B(new_n946), .Y(new_n952));
  nand_5 g0637(.A(new_n951), .B(new_n951), .Y(new_n953));
  nor_5      g0638(.A(new_n953), .B(new_n945), .Y(new_n954));
  or_6       g0639(.A(new_n954), .B(new_n952), .Y(new_n955));
  nor_5      g0640(.A(new_n955), .B(new_n949), .Y(po029));
  nand_5     g0641(.A(new_n940), .B(new_n938), .Y(new_n957));
  nand_5 g0642(.A(new_n865), .B(new_n865), .Y(new_n958));
  or_6       g0643(.A(new_n868), .B(pi204), .Y(new_n959));
  nand_5     g0644(.A(new_n959), .B(new_n958), .Y(new_n960));
  xor_4      g0645(.A(new_n960), .B(new_n957), .Y(new_n961));
  xor_4      g0646(.A(new_n961), .B(po029), .Y(new_n962));
  nand_5     g0647(.A(pi024), .B(pi022), .Y(new_n963));
  xor_4      g0648(.A(new_n963), .B(new_n947), .Y(po030));
  xor_4      g0649(.A(pi181), .B(new_n766), .Y(new_n965));
  xor_4      g0650(.A(pi184), .B(pi077), .Y(new_n966));
  xor_4      g0651(.A(new_n966), .B(pi062), .Y(new_n967));
  nand_5     g0652(.A(pi145), .B(pi061), .Y(new_n968));
  or_6       g0653(.A(pi145), .B(pi061), .Y(new_n969));
  nand_5     g0654(.A(new_n969), .B(new_n759), .Y(new_n970));
  nand_5     g0655(.A(new_n970), .B(new_n968), .Y(new_n971));
  nand_5     g0656(.A(new_n971), .B(new_n967), .Y(new_n972));
  nor_5      g0657(.A(new_n971), .B(new_n967), .Y(new_n973));
  nand_5     g0658(.A(new_n316), .B(pi150), .Y(new_n974));
  nor_5      g0659(.A(new_n974), .B(new_n973), .Y(new_n975));
  nand_5     g0660(.A(new_n975), .B(new_n972), .Y(new_n976));
  nand_5     g0661(.A(new_n871), .B(new_n958), .Y(new_n977));
  nand_5     g0662(.A(new_n977), .B(new_n872), .Y(new_n978));
  xor_4      g0663(.A(new_n978), .B(new_n976), .Y(new_n979));
  xor_4      g0664(.A(new_n979), .B(new_n965), .Y(new_n980));
  xor_4      g0665(.A(new_n980), .B(po030), .Y(new_n981));
  xor_4      g0666(.A(new_n981), .B(new_n962), .Y(po026));
  xnor_4     g0667(.A(new_n531), .B(new_n327), .Y(po027));
  xor_4      g0668(.A(new_n515), .B(new_n514), .Y(po038));
  xor_4      g0669(.A(new_n523), .B(new_n350), .Y(po039));
  nand_5 g0670(.A(pi064), .B(pi064), .Y(new_n986));
  nor_5      g0671(.A(new_n963), .B(new_n986), .Y(new_n987));
  nor_5      g0672(.A(new_n987), .B(new_n847), .Y(new_n988));
  nor_5      g0673(.A(new_n988), .B(new_n944), .Y(new_n989));
  nor_5      g0674(.A(pi064), .B(pi024), .Y(new_n990));
  nor_5      g0675(.A(new_n990), .B(new_n856), .Y(new_n991));
  nor_5      g0676(.A(new_n991), .B(new_n989), .Y(po040));
  xor_4      g0677(.A(new_n457), .B(pi070), .Y(po043));
  xor_4      g0678(.A(pi192), .B(pi107), .Y(new_n994));
  xor_4      g0679(.A(new_n994), .B(new_n387), .Y(new_n995));
  xnor_4     g0680(.A(new_n490), .B(new_n410), .Y(po069));
  xor_4      g0681(.A(po069), .B(new_n995), .Y(new_n997));
  xor_4      g0682(.A(new_n997), .B(po005), .Y(new_n998));
  xor_4      g0683(.A(new_n998), .B(po038), .Y(new_n999));
  nand_5 g0684(.A(new_n379), .B(new_n379), .Y(new_n1000));
  nand_5     g0685(.A(new_n510), .B(new_n1000), .Y(new_n1001));
  or_6       g0686(.A(new_n510), .B(new_n380), .Y(new_n1002));
  nand_5     g0687(.A(new_n1002), .B(new_n1001), .Y(new_n1003));
  nand_5     g0688(.A(pi189), .B(pi139), .Y(new_n1004));
  nand_5     g0689(.A(new_n393), .B(new_n370), .Y(new_n1005));
  nand_5     g0690(.A(new_n1005), .B(new_n1004), .Y(new_n1006));
  nand_5     g0691(.A(new_n1006), .B(new_n394), .Y(new_n1007));
  xor_4      g0692(.A(pi142), .B(pi094), .Y(new_n1008));
  or_6       g0693(.A(new_n1008), .B(pi150), .Y(new_n1009));
  xnor_4     g0694(.A(pi187), .B(pi090), .Y(new_n1010));
  nand_5     g0695(.A(new_n1010), .B(pi032), .Y(new_n1011));
  nor_5      g0696(.A(new_n1010), .B(pi032), .Y(new_n1012));
  nor_5      g0697(.A(new_n1012), .B(new_n328), .Y(new_n1013));
  nand_5     g0698(.A(new_n1013), .B(new_n1011), .Y(new_n1014));
  nand_5     g0699(.A(new_n1014), .B(new_n1009), .Y(new_n1015));
  xnor_4     g0700(.A(new_n1015), .B(new_n1007), .Y(new_n1016));
  nand_5     g0701(.A(new_n503), .B(new_n498), .Y(new_n1017));
  or_6       g0702(.A(new_n492), .B(new_n404), .Y(new_n1018));
  nand_5 g0703(.A(new_n402), .B(new_n402), .Y(new_n1019));
  nand_5     g0704(.A(new_n492), .B(new_n1019), .Y(new_n1020));
  nand_5     g0705(.A(new_n1020), .B(new_n1018), .Y(new_n1021));
  xor_4      g0706(.A(new_n1021), .B(new_n1017), .Y(new_n1022));
  xor_4      g0707(.A(new_n1022), .B(new_n1016), .Y(new_n1023));
  xor_4      g0708(.A(new_n1023), .B(new_n1003), .Y(new_n1024));
  xnor_4     g0709(.A(new_n1024), .B(new_n999), .Y(po044));
  nand_5     g0710(.A(pi126), .B(pi046), .Y(new_n1026));
  nand_5     g0711(.A(pi191), .B(pi176), .Y(new_n1027));
  nor_5      g0712(.A(new_n1027), .B(new_n1026), .Y(new_n1028));
  nand_5 g0713(.A(new_n1028), .B(new_n1028), .Y(po047));
  nand_5     g0714(.A(new_n1020), .B(new_n494), .Y(new_n1030));
  nand_5     g0715(.A(new_n1030), .B(new_n1018), .Y(po048));
  xnor_4     g0716(.A(new_n488), .B(new_n487), .Y(po049));
  or_6       g0717(.A(pi165), .B(pi148), .Y(po050));
  xor_4      g0718(.A(new_n464), .B(new_n444), .Y(po054));
  nand_5     g0719(.A(new_n525), .B(new_n344), .Y(new_n1035));
  nand_5 g0720(.A(new_n527), .B(new_n527), .Y(new_n1036));
  nand_5 g0721(.A(new_n525), .B(new_n525), .Y(new_n1037));
  nand_5     g0722(.A(new_n1037), .B(new_n343), .Y(new_n1038));
  nand_5     g0723(.A(new_n1038), .B(new_n1036), .Y(new_n1039));
  nand_5     g0724(.A(new_n1039), .B(new_n1035), .Y(po057));
  xnor_4     g0725(.A(new_n872), .B(new_n871), .Y(po058));
  xor_4      g0726(.A(pi084), .B(new_n778), .Y(new_n1042));
  xor_4      g0727(.A(pi110), .B(pi105), .Y(new_n1043));
  xor_4      g0728(.A(new_n1043), .B(new_n770), .Y(new_n1044));
  nand_5     g0729(.A(new_n1044), .B(new_n1042), .Y(new_n1045));
  nor_5      g0730(.A(new_n1044), .B(new_n1042), .Y(new_n1046));
  nor_5      g0731(.A(new_n1046), .B(new_n550), .Y(new_n1047));
  nand_5     g0732(.A(new_n1047), .B(new_n1045), .Y(new_n1048));
  xor_4      g0733(.A(pi174), .B(new_n569), .Y(new_n1049));
  xor_4      g0734(.A(new_n1049), .B(pi127), .Y(new_n1050));
  xor_4      g0735(.A(pi082), .B(pi006), .Y(new_n1051));
  xor_4      g0736(.A(new_n1051), .B(new_n1050), .Y(new_n1052));
  xor_4      g0737(.A(new_n1052), .B(new_n1048), .Y(new_n1053));
  xor_4      g0738(.A(pi028), .B(new_n836), .Y(new_n1054));
  xor_4      g0739(.A(new_n1054), .B(pi008), .Y(new_n1055));
  xor_4      g0740(.A(new_n775), .B(pi168), .Y(new_n1056));
  xor_4      g0741(.A(pi159), .B(pi031), .Y(new_n1057));
  xor_4      g0742(.A(new_n1057), .B(new_n1056), .Y(new_n1058));
  xor_4      g0743(.A(new_n1058), .B(new_n1055), .Y(new_n1059));
  nor_5      g0744(.A(new_n1059), .B(new_n550), .Y(new_n1060));
  nor_5      g0745(.A(new_n1060), .B(new_n328), .Y(new_n1061));
  nand_5     g0746(.A(new_n1061), .B(new_n1053), .Y(new_n1062));
  xor_4      g0747(.A(pi072), .B(pi052), .Y(new_n1063));
  nand_5     g0748(.A(pi036), .B(pi011), .Y(new_n1064));
  nor_5      g0749(.A(pi036), .B(pi011), .Y(new_n1065));
  nor_5      g0750(.A(new_n1065), .B(new_n328), .Y(new_n1066));
  nand_5     g0751(.A(new_n1066), .B(new_n1064), .Y(new_n1067));
  nand_5     g0752(.A(new_n1067), .B(new_n1006), .Y(new_n1068));
  nand_5     g0753(.A(new_n625), .B(pi097), .Y(new_n1069));
  nor_5      g0754(.A(new_n625), .B(pi097), .Y(new_n1070));
  nor_5      g0755(.A(new_n1070), .B(new_n328), .Y(new_n1071));
  nand_5     g0756(.A(new_n1071), .B(new_n1069), .Y(new_n1072));
  nand_5     g0757(.A(new_n1072), .B(new_n1009), .Y(new_n1073));
  xnor_4     g0758(.A(new_n1073), .B(new_n1068), .Y(new_n1074));
  xor_4      g0759(.A(pi114), .B(pi005), .Y(new_n1075));
  nor_5      g0760(.A(new_n1075), .B(new_n328), .Y(new_n1076));
  xor_4      g0761(.A(pi146), .B(pi086), .Y(new_n1077));
  nor_5      g0762(.A(new_n1077), .B(pi150), .Y(new_n1078));
  nor_5      g0763(.A(new_n1078), .B(new_n1076), .Y(new_n1079));
  xor_4      g0764(.A(new_n1079), .B(new_n1074), .Y(new_n1080));
  xor_4      g0765(.A(pi135), .B(new_n612), .Y(new_n1081));
  nand_5     g0766(.A(new_n1081), .B(pi150), .Y(new_n1082));
  xnor_4     g0767(.A(pi156), .B(pi131), .Y(new_n1083));
  nand_5     g0768(.A(new_n1083), .B(new_n328), .Y(new_n1084));
  nand_5     g0769(.A(new_n1084), .B(new_n1082), .Y(new_n1085));
  xor_4      g0770(.A(new_n1085), .B(new_n1080), .Y(new_n1086));
  xor_4      g0771(.A(new_n1086), .B(new_n1063), .Y(new_n1087));
  nor_5      g0772(.A(new_n1087), .B(new_n1062), .Y(new_n1088));
  xnor_4     g0773(.A(pi136), .B(pi034), .Y(new_n1089));
  nor_5      g0774(.A(new_n1086), .B(new_n1089), .Y(new_n1090));
  xor_4      g0775(.A(pi203), .B(new_n338), .Y(new_n1091));
  xor_4      g0776(.A(new_n1091), .B(pi134), .Y(new_n1092));
  xor_4      g0777(.A(pi177), .B(pi151), .Y(new_n1093));
  xor_4      g0778(.A(new_n1093), .B(new_n550), .Y(new_n1094));
  nor_5      g0779(.A(new_n1094), .B(new_n1092), .Y(new_n1095));
  nand_5     g0780(.A(new_n1094), .B(new_n1092), .Y(new_n1096));
  nand_5     g0781(.A(new_n1096), .B(new_n328), .Y(new_n1097));
  nor_5      g0782(.A(new_n1097), .B(new_n1095), .Y(new_n1098));
  nand_5     g0783(.A(new_n1086), .B(new_n1089), .Y(new_n1099));
  nand_5     g0784(.A(new_n1099), .B(new_n1098), .Y(new_n1100));
  nor_5      g0785(.A(new_n1100), .B(new_n1090), .Y(new_n1101));
  nor_5      g0786(.A(new_n1101), .B(new_n1088), .Y(new_n1102));
  nand_5     g0787(.A(new_n903), .B(new_n328), .Y(new_n1103));
  xor_4      g0788(.A(pi171), .B(new_n603), .Y(new_n1104));
  nand_5     g0789(.A(new_n1104), .B(pi150), .Y(new_n1105));
  nand_5     g0790(.A(new_n1105), .B(new_n1103), .Y(new_n1106));
  xor_4      g0791(.A(pi206), .B(new_n584), .Y(new_n1107));
  nand_5     g0792(.A(new_n1107), .B(pi150), .Y(new_n1108));
  nand_5     g0793(.A(new_n905), .B(new_n328), .Y(new_n1109));
  nand_5     g0794(.A(new_n1109), .B(new_n1108), .Y(new_n1110));
  nor_5      g0795(.A(pi067), .B(pi038), .Y(new_n1111));
  nand_5     g0796(.A(pi067), .B(pi038), .Y(new_n1112));
  nand_5     g0797(.A(new_n1112), .B(pi150), .Y(new_n1113));
  nor_5      g0798(.A(new_n1113), .B(new_n1111), .Y(new_n1114));
  nor_5      g0799(.A(new_n423), .B(pi081), .Y(new_n1115));
  nor_5      g0800(.A(new_n481), .B(pi042), .Y(new_n1116));
  or_6       g0801(.A(new_n1116), .B(new_n1115), .Y(new_n1117));
  nor_5      g0802(.A(new_n1117), .B(new_n1114), .Y(new_n1118));
  xnor_4     g0803(.A(pi129), .B(pi089), .Y(new_n1119));
  nor_5      g0804(.A(new_n1119), .B(new_n328), .Y(new_n1120));
  nor_5      g0805(.A(pi143), .B(pi040), .Y(new_n1121));
  nand_5     g0806(.A(pi143), .B(pi040), .Y(new_n1122));
  nand_5     g0807(.A(new_n1122), .B(new_n328), .Y(new_n1123));
  nor_5      g0808(.A(new_n1123), .B(new_n1121), .Y(new_n1124));
  or_6       g0809(.A(new_n1124), .B(new_n1120), .Y(new_n1125));
  nand_5     g0810(.A(pi055), .B(pi002), .Y(new_n1126));
  nor_5      g0811(.A(pi055), .B(pi002), .Y(new_n1127));
  nor_5      g0812(.A(new_n1127), .B(new_n328), .Y(new_n1128));
  nand_5     g0813(.A(new_n1128), .B(new_n1126), .Y(new_n1129));
  nand_5     g0814(.A(new_n1129), .B(new_n439), .Y(new_n1130));
  xor_4      g0815(.A(new_n1130), .B(new_n1125), .Y(new_n1131));
  xor_4      g0816(.A(new_n1131), .B(new_n1118), .Y(new_n1132));
  xor_4      g0817(.A(new_n1132), .B(new_n1110), .Y(new_n1133));
  xor_4      g0818(.A(new_n1133), .B(new_n1106), .Y(new_n1134));
  nor_5      g0819(.A(new_n1134), .B(new_n1102), .Y(new_n1135));
  xor_4      g0820(.A(pi183), .B(pi170), .Y(new_n1136));
  nand_5     g0821(.A(new_n1136), .B(pi150), .Y(new_n1137));
  nand_5     g0822(.A(pi166), .B(pi149), .Y(new_n1138));
  nor_5      g0823(.A(pi166), .B(pi149), .Y(new_n1139));
  nor_5      g0824(.A(new_n1139), .B(pi150), .Y(new_n1140));
  nand_5     g0825(.A(new_n1140), .B(new_n1138), .Y(new_n1141));
  nand_5     g0826(.A(new_n1141), .B(new_n1137), .Y(new_n1142));
  xor_4      g0827(.A(pi160), .B(new_n403), .Y(new_n1143));
  nor_5      g0828(.A(new_n1143), .B(new_n328), .Y(new_n1144));
  nor_5      g0829(.A(pi201), .B(pi104), .Y(new_n1145));
  nand_5     g0830(.A(pi201), .B(pi104), .Y(new_n1146));
  nand_5     g0831(.A(new_n1146), .B(new_n328), .Y(new_n1147));
  nor_5      g0832(.A(new_n1147), .B(new_n1145), .Y(new_n1148));
  or_6       g0833(.A(new_n1148), .B(new_n1144), .Y(new_n1149));
  xor_4      g0834(.A(pi116), .B(new_n381), .Y(new_n1150));
  nor_5      g0835(.A(new_n1150), .B(new_n328), .Y(new_n1151));
  nor_5      g0836(.A(pi179), .B(pi016), .Y(new_n1152));
  nand_5     g0837(.A(pi179), .B(pi016), .Y(new_n1153));
  nand_5     g0838(.A(new_n1153), .B(new_n328), .Y(new_n1154));
  nor_5      g0839(.A(new_n1154), .B(new_n1152), .Y(new_n1155));
  nor_5      g0840(.A(new_n1155), .B(new_n1151), .Y(new_n1156));
  xor_4      g0841(.A(new_n1156), .B(new_n1149), .Y(new_n1157));
  xor_4      g0842(.A(new_n1157), .B(new_n1142), .Y(new_n1158));
  xor_4      g0843(.A(pi113), .B(pi068), .Y(new_n1159));
  xor_4      g0844(.A(pi205), .B(pi138), .Y(new_n1160));
  xor_4      g0845(.A(new_n1160), .B(new_n1159), .Y(new_n1161));
  xor_4      g0846(.A(new_n1161), .B(new_n1158), .Y(new_n1162));
  xor_4      g0847(.A(pi112), .B(new_n553), .Y(new_n1163));
  xor_4      g0848(.A(pi108), .B(new_n756), .Y(new_n1164));
  nor_5      g0849(.A(new_n1164), .B(new_n328), .Y(new_n1165));
  nor_5      g0850(.A(pi163), .B(pi073), .Y(new_n1166));
  nand_5     g0851(.A(pi163), .B(pi073), .Y(new_n1167));
  nand_5     g0852(.A(new_n1167), .B(new_n328), .Y(new_n1168));
  nor_5      g0853(.A(new_n1168), .B(new_n1166), .Y(new_n1169));
  nor_5      g0854(.A(new_n1169), .B(new_n1165), .Y(new_n1170));
  nand_5     g0855(.A(new_n950), .B(pi150), .Y(new_n1171));
  nand_5     g0856(.A(new_n851), .B(new_n328), .Y(new_n1172));
  or_6       g0857(.A(new_n1172), .B(new_n855), .Y(new_n1173));
  nand_5     g0858(.A(new_n1173), .B(new_n1171), .Y(new_n1174));
  xor_4      g0859(.A(pi204), .B(new_n759), .Y(new_n1175));
  nand_5     g0860(.A(new_n1175), .B(pi150), .Y(new_n1176));
  xor_4      g0861(.A(pi088), .B(pi019), .Y(new_n1177));
  or_6       g0862(.A(new_n1177), .B(pi150), .Y(new_n1178));
  nand_5     g0863(.A(new_n1178), .B(new_n1176), .Y(new_n1179));
  xnor_4     g0864(.A(new_n1179), .B(new_n1174), .Y(new_n1180));
  xor_4      g0865(.A(new_n1180), .B(new_n1170), .Y(new_n1181));
  nor_5      g0866(.A(new_n1181), .B(new_n1163), .Y(new_n1182));
  nand_5     g0867(.A(new_n1181), .B(new_n1163), .Y(new_n1183));
  xnor_4     g0868(.A(pi098), .B(pi096), .Y(new_n1184));
  xor_4      g0869(.A(new_n1184), .B(pi066), .Y(new_n1185));
  xor_4      g0870(.A(pi023), .B(pi021), .Y(new_n1186));
  xor_4      g0871(.A(new_n1186), .B(new_n1185), .Y(new_n1187));
  xor_4      g0872(.A(pi048), .B(pi029), .Y(new_n1188));
  xor_4      g0873(.A(pi111), .B(pi100), .Y(new_n1189));
  xor_4      g0874(.A(new_n1189), .B(pi117), .Y(new_n1190));
  xor_4      g0875(.A(new_n1190), .B(new_n1188), .Y(new_n1191));
  xor_4      g0876(.A(new_n1191), .B(new_n1187), .Y(new_n1192));
  nor_5      g0877(.A(new_n1192), .B(pi150), .Y(new_n1193));
  nand_5     g0878(.A(new_n1193), .B(new_n1183), .Y(new_n1194));
  or_6       g0879(.A(new_n1194), .B(new_n1182), .Y(new_n1195));
  nor_5      g0880(.A(new_n1195), .B(new_n1162), .Y(new_n1196));
  xor_4      g0881(.A(pi074), .B(new_n438), .Y(new_n1197));
  xor_4      g0882(.A(pi147), .B(pi137), .Y(new_n1198));
  xor_4      g0883(.A(new_n1198), .B(pi027), .Y(new_n1199));
  xor_4      g0884(.A(new_n1199), .B(new_n884), .Y(new_n1200));
  xor_4      g0885(.A(new_n1200), .B(new_n1197), .Y(new_n1201));
  nand_5     g0886(.A(new_n1201), .B(pi150), .Y(new_n1202));
  xor_4      g0887(.A(new_n1181), .B(new_n965), .Y(new_n1203));
  xor_4      g0888(.A(new_n995), .B(pi118), .Y(new_n1204));
  xor_4      g0889(.A(new_n1204), .B(new_n1158), .Y(new_n1205));
  nand_5     g0890(.A(new_n1205), .B(new_n1203), .Y(new_n1206));
  nor_5      g0891(.A(new_n1206), .B(new_n1202), .Y(new_n1207));
  or_6       g0892(.A(new_n1207), .B(new_n1196), .Y(new_n1208));
  xor_4      g0893(.A(pi178), .B(new_n357), .Y(new_n1209));
  nand_5     g0894(.A(new_n1209), .B(pi150), .Y(new_n1210));
  nand_5     g0895(.A(pi140), .B(new_n732), .Y(new_n1211));
  nor_5      g0896(.A(pi140), .B(new_n732), .Y(new_n1212));
  nor_5      g0897(.A(new_n1212), .B(pi150), .Y(new_n1213));
  nand_5     g0898(.A(new_n1213), .B(new_n1211), .Y(new_n1214));
  nand_5     g0899(.A(new_n1214), .B(new_n1210), .Y(new_n1215));
  nand_5     g0900(.A(pi141), .B(pi010), .Y(new_n1216));
  nand_5     g0901(.A(new_n798), .B(new_n787), .Y(new_n1217));
  nand_5     g0902(.A(new_n1217), .B(new_n1216), .Y(new_n1218));
  nand_5     g0903(.A(pi122), .B(pi056), .Y(new_n1219));
  nor_5      g0904(.A(pi122), .B(pi056), .Y(new_n1220));
  nor_5      g0905(.A(new_n1220), .B(new_n328), .Y(new_n1221));
  nand_5     g0906(.A(new_n1221), .B(new_n1219), .Y(new_n1222));
  nand_5     g0907(.A(new_n1222), .B(new_n1218), .Y(new_n1223));
  xor_4      g0908(.A(pi196), .B(pi001), .Y(new_n1224));
  nand_5     g0909(.A(new_n1224), .B(pi150), .Y(new_n1225));
  nand_5     g0910(.A(pi202), .B(pi161), .Y(new_n1226));
  nor_5      g0911(.A(pi202), .B(pi161), .Y(new_n1227));
  nor_5      g0912(.A(new_n1227), .B(pi150), .Y(new_n1228));
  nand_5     g0913(.A(new_n1228), .B(new_n1226), .Y(new_n1229));
  nand_5     g0914(.A(new_n1229), .B(new_n1225), .Y(new_n1230));
  xnor_4     g0915(.A(new_n1230), .B(new_n1223), .Y(new_n1231));
  xor_4      g0916(.A(new_n1231), .B(new_n1215), .Y(new_n1232));
  xor_4      g0917(.A(pi199), .B(new_n793), .Y(new_n1233));
  nand_5     g0918(.A(new_n1233), .B(pi150), .Y(new_n1234));
  xor_4      g0919(.A(new_n797), .B(pi173), .Y(new_n1235));
  nand_5     g0920(.A(new_n1235), .B(new_n328), .Y(new_n1236));
  nand_5     g0921(.A(new_n1236), .B(new_n1234), .Y(new_n1237));
  xor_4      g0922(.A(pi153), .B(new_n762), .Y(new_n1238));
  nand_5     g0923(.A(new_n1238), .B(pi150), .Y(new_n1239));
  nand_5     g0924(.A(new_n788), .B(new_n749), .Y(new_n1240));
  nand_5     g0925(.A(new_n1240), .B(new_n328), .Y(new_n1241));
  nand_5     g0926(.A(new_n1241), .B(new_n1239), .Y(new_n1242));
  xor_4      g0927(.A(new_n1242), .B(new_n1237), .Y(new_n1243));
  xor_4      g0928(.A(new_n1243), .B(new_n1232), .Y(new_n1244));
  nand_5     g0929(.A(new_n1244), .B(new_n1208), .Y(po086));
  xor_4      g0930(.A(pi058), .B(pi042), .Y(new_n1246));
  xor_4      g0931(.A(new_n1246), .B(pi040), .Y(new_n1247));
  xor_4      g0932(.A(new_n1247), .B(new_n907), .Y(new_n1248));
  nand_5     g0933(.A(new_n1248), .B(new_n1098), .Y(new_n1249));
  xor_4      g0934(.A(pi200), .B(new_n861), .Y(new_n1250));
  xor_4      g0935(.A(pi102), .B(pi061), .Y(new_n1251));
  xor_4      g0936(.A(new_n1251), .B(new_n1250), .Y(new_n1252));
  nand_5     g0937(.A(new_n1252), .B(new_n967), .Y(new_n1253));
  nor_5      g0938(.A(new_n1252), .B(new_n967), .Y(new_n1254));
  nor_5      g0939(.A(new_n1254), .B(new_n550), .Y(new_n1255));
  nand_5     g0940(.A(new_n1255), .B(new_n1253), .Y(new_n1256));
  nand_5     g0941(.A(new_n1256), .B(pi150), .Y(new_n1257));
  xor_4      g0942(.A(pi155), .B(pi120), .Y(new_n1258));
  xor_4      g0943(.A(pi044), .B(pi025), .Y(new_n1259));
  xnor_4     g0944(.A(new_n1259), .B(new_n1258), .Y(new_n1260));
  xnor_4     g0945(.A(new_n1260), .B(new_n900), .Y(new_n1261));
  nor_5      g0946(.A(new_n1261), .B(new_n1257), .Y(new_n1262));
  xor_4      g0947(.A(pi182), .B(pi009), .Y(new_n1263));
  xor_4      g0948(.A(new_n1263), .B(pi017), .Y(new_n1264));
  xor_4      g0949(.A(pi175), .B(pi026), .Y(new_n1265));
  xor_4      g0950(.A(new_n1265), .B(new_n317), .Y(new_n1266));
  xor_4      g0951(.A(pi154), .B(new_n321), .Y(new_n1267));
  nor_5      g0952(.A(new_n1267), .B(new_n1266), .Y(new_n1268));
  nand_5     g0953(.A(new_n1267), .B(new_n1266), .Y(new_n1269));
  nand_5     g0954(.A(new_n1269), .B(new_n316), .Y(new_n1270));
  nor_5      g0955(.A(new_n1270), .B(new_n1268), .Y(new_n1271));
  xor_4      g0956(.A(pi172), .B(pi080), .Y(new_n1272));
  xor_4      g0957(.A(new_n1272), .B(new_n1271), .Y(new_n1273));
  xor_4      g0958(.A(new_n1273), .B(new_n1264), .Y(new_n1274));
  nand_5     g0959(.A(new_n1274), .B(new_n1262), .Y(new_n1275));
  nand_5     g0960(.A(new_n1275), .B(new_n1249), .Y(new_n1276));
  xor_4      g0961(.A(pi194), .B(pi164), .Y(new_n1277));
  xor_4      g0962(.A(pi158), .B(pi045), .Y(new_n1278));
  xor_4      g0963(.A(pi030), .B(pi012), .Y(new_n1279));
  xnor_4     g0964(.A(new_n1279), .B(new_n1278), .Y(new_n1280));
  xor_4      g0965(.A(new_n1280), .B(new_n1277), .Y(new_n1281));
  or_6       g0966(.A(new_n1281), .B(new_n328), .Y(new_n1282));
  xor_4      g0967(.A(new_n1083), .B(new_n1089), .Y(new_n1283));
  xor_4      g0968(.A(new_n1283), .B(new_n1077), .Y(new_n1284));
  nand_5     g0969(.A(new_n1284), .B(new_n328), .Y(new_n1285));
  nand_5     g0970(.A(new_n1285), .B(new_n1282), .Y(new_n1286));
  xor_4      g0971(.A(new_n1286), .B(new_n1016), .Y(new_n1287));
  nand_5     g0972(.A(new_n1287), .B(new_n1276), .Y(po080));
  nor_5      g0973(.A(po047), .B(po006), .Y(new_n1289));
  nand_5     g0974(.A(pi076), .B(pi063), .Y(new_n1290));
  nand_5     g0975(.A(pi133), .B(pi099), .Y(new_n1291));
  nor_5      g0976(.A(new_n1291), .B(new_n1290), .Y(new_n1292));
  nand_5 g0977(.A(new_n1292), .B(new_n1292), .Y(po107));
  nand_5     g0978(.A(pi128), .B(pi079), .Y(new_n1294));
  nand_5     g0979(.A(pi157), .B(pi130), .Y(new_n1295));
  nor_5      g0980(.A(new_n1295), .B(new_n1294), .Y(new_n1296));
  nand_5 g0981(.A(new_n1296), .B(new_n1296), .Y(po100));
  nor_5      g0982(.A(po100), .B(po107), .Y(new_n1298));
  nand_5     g0983(.A(new_n1298), .B(new_n1289), .Y(new_n1299));
  or_6       g0984(.A(new_n1299), .B(po080), .Y(new_n1300));
  nor_5      g0985(.A(new_n1300), .B(po086), .Y(new_n1301));
  nand_5     g0986(.A(new_n1301), .B(new_n1135), .Y(po059));
  xnor_4     g0987(.A(new_n494), .B(new_n397), .Y(po060));
  xnor_4     g0988(.A(new_n942), .B(new_n941), .Y(po061));
  xor_4      g0989(.A(new_n474), .B(new_n473), .Y(po062));
  nand_5     g0990(.A(pi093), .B(pi053), .Y(new_n1306));
  or_6       g0991(.A(new_n1306), .B(pi165), .Y(po065));
  nor_5      g0992(.A(new_n521), .B(new_n356), .Y(new_n1308));
  nand_5 g0993(.A(new_n1308), .B(new_n1308), .Y(new_n1309));
  nor_5      g0994(.A(new_n520), .B(new_n355), .Y(new_n1310));
  nand_5 g0995(.A(new_n1310), .B(new_n1310), .Y(new_n1311));
  nand_5     g0996(.A(new_n1311), .B(new_n523), .Y(new_n1312));
  and_6      g0997(.A(new_n1312), .B(new_n1309), .Y(po066));
  xor_4      g0998(.A(new_n466), .B(new_n437), .Y(po067));
  nand_5     g0999(.A(new_n1001), .B(new_n512), .Y(new_n1315));
  nand_5     g1000(.A(new_n1315), .B(new_n1002), .Y(po068));
  nand_5     g1001(.A(new_n1311), .B(new_n1309), .Y(new_n1317));
  nand_5 g1002(.A(new_n974), .B(new_n974), .Y(new_n1318));
  nand_5     g1003(.A(new_n1265), .B(new_n1318), .Y(new_n1319));
  xor_4      g1004(.A(new_n1319), .B(new_n1317), .Y(new_n1320));
  xor_4      g1005(.A(new_n348), .B(pi153), .Y(new_n1321));
  xor_4      g1006(.A(new_n1321), .B(po011), .Y(new_n1322));
  xor_4      g1007(.A(new_n1322), .B(new_n1320), .Y(new_n1323));
  xor_4      g1008(.A(new_n1233), .B(po027), .Y(new_n1324));
  xor_4      g1009(.A(new_n1324), .B(new_n1323), .Y(new_n1325));
  nand_5     g1010(.A(new_n534), .B(new_n533), .Y(new_n1326));
  nand_5     g1011(.A(new_n926), .B(new_n320), .Y(new_n1327));
  nand_5     g1012(.A(new_n1327), .B(new_n1326), .Y(new_n1328));
  xor_4      g1013(.A(new_n518), .B(new_n517), .Y(po095));
  nand_5     g1014(.A(new_n1038), .B(new_n1035), .Y(new_n1330));
  xor_4      g1015(.A(new_n1330), .B(po095), .Y(new_n1331));
  xor_4      g1016(.A(new_n1331), .B(new_n1328), .Y(new_n1332));
  xor_4      g1017(.A(new_n1332), .B(new_n1325), .Y(po070));
  xnor_4     g1018(.A(new_n485), .B(new_n483), .Y(po073));
  xor_4      g1019(.A(new_n874), .B(new_n958), .Y(po083));
  nand_5 g1020(.A(new_n1135), .B(new_n1135), .Y(po090));
  xor_4      g1021(.A(new_n939), .B(new_n937), .Y(po091));
  xor_4      g1022(.A(new_n462), .B(new_n461), .Y(po092));
  xor_4      g1023(.A(new_n477), .B(new_n476), .Y(po094));
  xor_4      g1024(.A(new_n470), .B(new_n468), .Y(po102));
  xnor_4     g1025(.A(new_n512), .B(new_n374), .Y(po104));
  buf_8      g1026(.A(pi050), .Y(po001));
  buf_8      g1027(.A(pi118), .Y(po002));
  buf_8      g1028(.A(pi020), .Y(po004));
  buf_8      g1029(.A(pi196), .Y(po007));
  buf_8      g1030(.A(pi107), .Y(po010));
  buf_8      g1031(.A(pi060), .Y(po012));
  buf_8      g1032(.A(pi108), .Y(po014));
  buf_8      g1033(.A(pi057), .Y(po018));
  buf_8      g1034(.A(pi047), .Y(po019));
  buf_8      g1035(.A(pi085), .Y(po021));
  buf_8      g1036(.A(pi180), .Y(po022));
  buf_8      g1037(.A(po003), .Y(po023));
  buf_8      g1038(.A(pi056), .Y(po028));
  buf_8      g1039(.A(po008), .Y(po031));
  buf_8      g1040(.A(pi001), .Y(po032));
  buf_8      g1041(.A(pi204), .Y(po033));
  buf_8      g1042(.A(pi039), .Y(po034));
  buf_8      g1043(.A(pi024), .Y(po035));
  buf_8      g1044(.A(pi101), .Y(po036));
  buf_8      g1045(.A(pi144), .Y(po037));
  buf_8      g1046(.A(po040), .Y(po041));
  buf_8      g1047(.A(pi160), .Y(po042));
  buf_8      g1048(.A(pi060), .Y(po045));
  buf_8      g1049(.A(pi162), .Y(po046));
  buf_8      g1050(.A(po017), .Y(po051));
  buf_8      g1051(.A(pi122), .Y(po052));
  buf_8      g1052(.A(pi027), .Y(po053));
  buf_8      g1053(.A(pi051), .Y(po055));
  buf_8      g1054(.A(pi147), .Y(po056));
  buf_8      g1055(.A(pi183), .Y(po063));
  buf_8      g1056(.A(pi192), .Y(po064));
  buf_8      g1057(.A(pi064), .Y(po071));
  buf_8      g1058(.A(po040), .Y(po072));
  buf_8      g1059(.A(pi132), .Y(po074));
  buf_8      g1060(.A(po008), .Y(po075));
  buf_8      g1061(.A(pi181), .Y(po076));
  buf_8      g1062(.A(pi083), .Y(po077));
  buf_8      g1063(.A(po065), .Y(po078));
  buf_8      g1064(.A(pi170), .Y(po079));
  buf_8      g1065(.A(pi199), .Y(po081));
  buf_8      g1066(.A(po017), .Y(po082));
  buf_8      g1067(.A(pi153), .Y(po085));
  buf_8      g1068(.A(pi137), .Y(po087));
  buf_8      g1069(.A(po030), .Y(po088));
  buf_8      g1070(.A(pi060), .Y(po089));
  buf_8      g1071(.A(pi092), .Y(po093));
  buf_8      g1072(.A(pi116), .Y(po096));
  buf_8      g1073(.A(pi060), .Y(po097));
  buf_8      g1074(.A(pi074), .Y(po098));
  buf_8      g1075(.A(po029), .Y(po099));
  buf_8      g1076(.A(po040), .Y(po101));
  buf_8      g1077(.A(pi178), .Y(po103));
  buf_8      g1078(.A(pi018), .Y(po105));
  buf_8      g1079(.A(pi004), .Y(po106));
endmodule


