// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Wed Aug 14 23:00:42 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119;
  wire new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n385, new_n386, new_n387, new_n388, new_n389, new_n390, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1875, new_n1876, new_n1877, new_n1878, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1890, new_n1891, new_n1892,
    new_n1893, new_n1894, new_n1895, new_n1896, new_n1897, new_n1898,
    new_n1899, new_n1900, new_n1901, new_n1902, new_n1903, new_n1904,
    new_n1905, new_n1906, new_n1907, new_n1908, new_n1909, new_n1910,
    new_n1911, new_n1912, new_n1913, new_n1914, new_n1915, new_n1916,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019,
    new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025,
    new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031,
    new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055,
    new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061,
    new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067,
    new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896,
    new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914,
    new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944,
    new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956,
    new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962,
    new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046,
    new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052,
    new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058,
    new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064,
    new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070,
    new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076,
    new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088,
    new_n3089, new_n3090, new_n3091, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3101, new_n3102, new_n3103, new_n3104, new_n3105, new_n3106,
    new_n3107, new_n3108, new_n3109, new_n3110, new_n3111, new_n3112,
    new_n3113, new_n3114, new_n3115, new_n3116, new_n3117, new_n3118,
    new_n3119, new_n3120, new_n3121, new_n3122, new_n3123, new_n3124,
    new_n3125, new_n3126, new_n3127, new_n3128, new_n3129, new_n3130,
    new_n3131, new_n3132, new_n3133, new_n3134, new_n3135, new_n3136,
    new_n3137, new_n3138, new_n3139, new_n3140, new_n3141, new_n3142,
    new_n3143, new_n3144, new_n3145, new_n3146, new_n3147, new_n3148,
    new_n3149, new_n3150, new_n3151, new_n3152, new_n3153, new_n3154,
    new_n3155, new_n3156, new_n3158, new_n3159, new_n3160, new_n3161,
    new_n3162, new_n3163, new_n3164, new_n3165, new_n3166, new_n3167,
    new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173,
    new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179,
    new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185,
    new_n3186, new_n3187, new_n3188, new_n3189, new_n3190, new_n3191,
    new_n3192, new_n3193, new_n3194, new_n3195, new_n3196, new_n3197,
    new_n3198, new_n3199, new_n3200, new_n3201, new_n3202, new_n3203,
    new_n3204, new_n3205, new_n3206, new_n3207, new_n3208, new_n3209,
    new_n3210, new_n3211, new_n3212, new_n3213, new_n3214, new_n3215,
    new_n3216, new_n3217, new_n3218, new_n3219, new_n3220, new_n3221,
    new_n3222, new_n3223, new_n3224, new_n3225, new_n3226, new_n3227,
    new_n3228, new_n3229, new_n3230, new_n3231, new_n3232, new_n3233,
    new_n3234, new_n3235, new_n3236, new_n3237, new_n3238, new_n3239,
    new_n3240, new_n3241, new_n3242, new_n3243, new_n3244, new_n3245,
    new_n3246, new_n3247, new_n3248, new_n3249, new_n3250, new_n3251,
    new_n3252, new_n3253, new_n3254, new_n3255, new_n3256, new_n3257,
    new_n3258, new_n3259, new_n3260, new_n3261, new_n3262, new_n3263,
    new_n3264, new_n3265, new_n3266, new_n3267, new_n3268, new_n3269,
    new_n3270, new_n3271, new_n3272, new_n3273, new_n3274, new_n3275,
    new_n3276, new_n3277, new_n3278, new_n3279, new_n3280, new_n3281,
    new_n3282, new_n3283, new_n3284, new_n3285, new_n3286, new_n3287,
    new_n3288, new_n3289, new_n3290, new_n3291, new_n3292, new_n3293,
    new_n3294, new_n3295, new_n3296, new_n3297, new_n3298, new_n3299,
    new_n3300, new_n3301, new_n3302, new_n3303, new_n3304, new_n3305,
    new_n3306, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516,
    new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552,
    new_n3553, new_n3555, new_n3556, new_n3557, new_n3558, new_n3559,
    new_n3560, new_n3564, new_n3565, new_n3566, new_n3567, new_n3568,
    new_n3569, new_n3570, new_n3571, new_n3572, new_n3573, new_n3574,
    new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577,
    new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583,
    new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589,
    new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595,
    new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601,
    new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607,
    new_n4608, new_n4609, new_n4610, new_n4611, new_n4612, new_n4613,
    new_n4614, new_n4615, new_n4616, new_n4617, new_n4618, new_n4619,
    new_n4620, new_n4621, new_n4622, new_n4623, new_n4624, new_n4625,
    new_n4626, new_n4627, new_n4628, new_n4629, new_n4630, new_n4631,
    new_n4632, new_n4633, new_n4634, new_n4635, new_n4636, new_n4637,
    new_n4638, new_n4639, new_n4640, new_n4641, new_n4642, new_n4643,
    new_n4644, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4886, new_n4887, new_n4888, new_n4889, new_n4890, new_n4891,
    new_n4892, new_n4893, new_n4894, new_n4895, new_n4896, new_n4897,
    new_n4898, new_n4899, new_n4900, new_n4901, new_n4902, new_n4903,
    new_n4904, new_n4905, new_n4906, new_n4907, new_n4908, new_n4909,
    new_n4910, new_n4911, new_n4912, new_n4913, new_n4914, new_n4915,
    new_n4916, new_n4917, new_n4918, new_n4919, new_n4920, new_n4921,
    new_n4922, new_n4923, new_n4924, new_n4925, new_n4926, new_n4927,
    new_n4928, new_n4929, new_n4930, new_n4931, new_n4932, new_n4933,
    new_n4934, new_n4935, new_n4936, new_n4937, new_n4938, new_n4939,
    new_n4940, new_n4941, new_n4942, new_n4943, new_n4944, new_n4945,
    new_n4946, new_n4947, new_n4948, new_n4949, new_n4950, new_n4951,
    new_n4952, new_n4953, new_n4954, new_n4955, new_n4956, new_n4957,
    new_n4958, new_n4959, new_n4960, new_n4961, new_n4962, new_n4963,
    new_n4964, new_n4965, new_n4966, new_n4967, new_n4968, new_n4969,
    new_n4970, new_n4971, new_n4972, new_n4973, new_n4974, new_n4975,
    new_n4976, new_n4977, new_n4978, new_n4979, new_n4980, new_n4981,
    new_n4982, new_n4983, new_n4984, new_n4985, new_n4986, new_n4987,
    new_n4988, new_n4989, new_n4990, new_n4991, new_n4992, new_n4993,
    new_n4994, new_n4995, new_n4996, new_n4997, new_n4998, new_n4999,
    new_n5000, new_n5001, new_n5002, new_n5003, new_n5004, new_n5005,
    new_n5006, new_n5007, new_n5008, new_n5009, new_n5010, new_n5011,
    new_n5012, new_n5013, new_n5014, new_n5015, new_n5016, new_n5017,
    new_n5018, new_n5019, new_n5020, new_n5021, new_n5022, new_n5023,
    new_n5024, new_n5025, new_n5026, new_n5027, new_n5028, new_n5029,
    new_n5030, new_n5031, new_n5033, new_n5034, new_n5035, new_n5036,
    new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5043, new_n5044, new_n5045, new_n5046, new_n5047, new_n5048,
    new_n5049, new_n5050, new_n5051, new_n5052, new_n5053, new_n5054,
    new_n5055, new_n5056, new_n5057, new_n5058, new_n5059, new_n5060,
    new_n5061, new_n5062, new_n5063, new_n5064, new_n5065, new_n5066,
    new_n5067, new_n5068, new_n5069, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6478, new_n6479, new_n6480, new_n6481,
    new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487,
    new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493,
    new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523,
    new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559,
    new_n6560, new_n6561, new_n6562, new_n6563, new_n6564, new_n6565,
    new_n6566, new_n6567, new_n6568, new_n6569, new_n6570, new_n6571,
    new_n6572, new_n6573, new_n6574, new_n6575, new_n6576, new_n6577,
    new_n6578, new_n6579, new_n6580, new_n6581, new_n6582, new_n6583,
    new_n6584, new_n6585, new_n6586, new_n6587, new_n6588, new_n6589,
    new_n6590, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595,
    new_n6596, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601,
    new_n6602, new_n6603, new_n6604, new_n6605, new_n6606, new_n6607,
    new_n6608, new_n6609, new_n6610, new_n6611, new_n6612, new_n6613,
    new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619,
    new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6628,
    new_n6629, new_n6630, new_n6631, new_n6632, new_n6633, new_n6634,
    new_n6635, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654,
    new_n6655, new_n6656, new_n6657, new_n6658, new_n6659, new_n6660,
    new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672,
    new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684,
    new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690,
    new_n6691, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229, new_n7230, new_n7231, new_n7232, new_n7233,
    new_n7234, new_n7235, new_n7236, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253, new_n7254, new_n7255, new_n7256, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7265, new_n7266, new_n7267, new_n7268, new_n7269,
    new_n7270, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275,
    new_n7276, new_n7277, new_n7278, new_n7279, new_n7280, new_n7281,
    new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287,
    new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293,
    new_n7294, new_n7295, new_n7296, new_n7297, new_n7298, new_n7299,
    new_n7300, new_n7301, new_n7302, new_n7303, new_n7304, new_n7305,
    new_n7306, new_n7307, new_n7308, new_n7309, new_n7310, new_n7311,
    new_n7312, new_n7313, new_n7314, new_n7315, new_n7316, new_n7317,
    new_n7318, new_n7319, new_n7320, new_n7321, new_n7322, new_n7323,
    new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329,
    new_n7330, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335,
    new_n7336, new_n7337, new_n7338, new_n7339, new_n7340, new_n7341,
    new_n7342, new_n7343, new_n7344, new_n7345, new_n7346, new_n7347,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717, new_n8718, new_n8719, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744, new_n8745, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9533, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763, new_n9764, new_n9765, new_n9766, new_n9767,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9831, new_n9832, new_n9833, new_n9834, new_n9835,
    new_n9836, new_n9837, new_n9838, new_n9839, new_n9840, new_n9841,
    new_n9842, new_n9843, new_n9844, new_n9845, new_n9846, new_n9847,
    new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865,
    new_n9866, new_n9867, new_n9868, new_n9869, new_n9870, new_n9871,
    new_n9872, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877,
    new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883,
    new_n9884, new_n9885, new_n9886, new_n9887, new_n9888, new_n9889,
    new_n9890, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895,
    new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901,
    new_n9902, new_n9903, new_n9904, new_n9905, new_n9906, new_n9907,
    new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915, new_n9916, new_n9917, new_n9918, new_n9919,
    new_n9920, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937,
    new_n9938, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997,
    new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003,
    new_n10004, new_n10005, new_n10014, new_n10015, new_n10016, new_n10017,
    new_n10018, new_n10019, new_n10020, new_n10021, new_n10022, new_n10023,
    new_n10024, new_n10025, new_n10026, new_n10027, new_n10028, new_n10029,
    new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035,
    new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041,
    new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047,
    new_n10048, new_n10049, new_n10050, new_n10051, new_n10052, new_n10053,
    new_n10054, new_n10055, new_n10056, new_n10057, new_n10058, new_n10059,
    new_n10060, new_n10061, new_n10062, new_n10063, new_n10064, new_n10065,
    new_n10066, new_n10067, new_n10068, new_n10069, new_n10070, new_n10071,
    new_n10072, new_n10073, new_n10074, new_n10075, new_n10076, new_n10077,
    new_n10078, new_n10079, new_n10080, new_n10081, new_n10082, new_n10083,
    new_n10084, new_n10085, new_n10086, new_n10087, new_n10088, new_n10089,
    new_n10090, new_n10091, new_n10092, new_n10093, new_n10094, new_n10095,
    new_n10096, new_n10097, new_n10098, new_n10099, new_n10100, new_n10101,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111, new_n10112, new_n10113,
    new_n10114, new_n10115, new_n10116, new_n10117, new_n10118, new_n10119,
    new_n10120, new_n10121, new_n10122, new_n10123, new_n10124, new_n10125,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10133, new_n10134, new_n10135, new_n10136, new_n10137,
    new_n10138, new_n10139, new_n10140, new_n10141, new_n10142, new_n10143,
    new_n10144, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158, new_n10159, new_n10160, new_n10161,
    new_n10162, new_n10163, new_n10164, new_n10165, new_n10166, new_n10167,
    new_n10168, new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174, new_n10175, new_n10176, new_n10177, new_n10178, new_n10179,
    new_n10180, new_n10181, new_n10182, new_n10183, new_n10184, new_n10185,
    new_n10186, new_n10187, new_n10188, new_n10189, new_n10190, new_n10191,
    new_n10192, new_n10193, new_n10194, new_n10195, new_n10196, new_n10197,
    new_n10198, new_n10199, new_n10200, new_n10201, new_n10202, new_n10203,
    new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209,
    new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215,
    new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236, new_n10237, new_n10238, new_n10239,
    new_n10240, new_n10241, new_n10242, new_n10243, new_n10244, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250, new_n10251,
    new_n10252, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10263,
    new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274, new_n10275,
    new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283, new_n10284, new_n10285, new_n10286, new_n10287,
    new_n10288, new_n10289, new_n10290, new_n10291, new_n10292, new_n10293,
    new_n10294, new_n10295, new_n10296, new_n10297, new_n10298, new_n10299,
    new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305,
    new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311,
    new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317,
    new_n10318, new_n10319, new_n10320, new_n10321, new_n10322, new_n10335,
    new_n10336, new_n10337, new_n10338, new_n10339, new_n10340, new_n10341,
    new_n10342, new_n10343, new_n10344, new_n10345, new_n10346, new_n10347,
    new_n10348, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377,
    new_n10378, new_n10379, new_n10380, new_n10381, new_n10382, new_n10383,
    new_n10384, new_n10385, new_n10386, new_n10387, new_n10388, new_n10389,
    new_n10390, new_n10391, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439, new_n10440, new_n10441, new_n10442, new_n10443,
    new_n10444, new_n10445, new_n10446, new_n10447, new_n10448, new_n10449,
    new_n10450, new_n10451, new_n10452, new_n10453, new_n10454, new_n10455,
    new_n10456, new_n10457, new_n10458, new_n10459, new_n10460, new_n10461,
    new_n10462, new_n10463, new_n10464, new_n10465, new_n10466, new_n10467,
    new_n10468, new_n10469, new_n10470, new_n10471, new_n10472, new_n10473,
    new_n10474, new_n10475, new_n10476, new_n10477, new_n10478, new_n10479,
    new_n10480, new_n10481, new_n10482, new_n10483, new_n10484, new_n10485,
    new_n10486, new_n10487, new_n10488, new_n10489, new_n10490, new_n10491,
    new_n10492, new_n10493, new_n10494, new_n10495, new_n10496, new_n10497,
    new_n10498, new_n10499, new_n10500, new_n10501, new_n10502, new_n10503,
    new_n10504, new_n10505, new_n10506, new_n10507, new_n10510, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545, new_n10546, new_n10547,
    new_n10548, new_n10549, new_n10550, new_n10551, new_n10552, new_n10553,
    new_n10554, new_n10555, new_n10556, new_n10557, new_n10558, new_n10559,
    new_n10560, new_n10561, new_n10562, new_n10563, new_n10564, new_n10565,
    new_n10566, new_n10567, new_n10568, new_n10569, new_n10570, new_n10571,
    new_n10572, new_n10573, new_n10574, new_n10575, new_n10576, new_n10577,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588, new_n10589,
    new_n10590, new_n10591, new_n10592, new_n10593, new_n10594, new_n10595,
    new_n10596, new_n10597, new_n10598, new_n10599, new_n10600, new_n10601,
    new_n10602, new_n10603, new_n10604, new_n10605, new_n10606, new_n10607,
    new_n10608, new_n10609, new_n10610, new_n10611, new_n10612, new_n10613,
    new_n10614, new_n10615, new_n10616, new_n10617, new_n10618, new_n10619,
    new_n10620, new_n10621, new_n10622, new_n10623, new_n10624, new_n10625,
    new_n10626, new_n10627, new_n10628, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647, new_n10648, new_n10649,
    new_n10650, new_n10651, new_n10652, new_n10653, new_n10654, new_n10655,
    new_n10656, new_n10657, new_n10658, new_n10659, new_n10660, new_n10661,
    new_n10662, new_n10663, new_n10664, new_n10665, new_n10666, new_n10667,
    new_n10668, new_n10669, new_n10670, new_n10671, new_n10672, new_n10673,
    new_n10674, new_n10675, new_n10676, new_n10677, new_n10678, new_n10679,
    new_n10680, new_n10681, new_n10682, new_n10683, new_n10695, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923, new_n10924,
    new_n10925, new_n10926, new_n10927, new_n10928, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954,
    new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961, new_n10962, new_n10963, new_n10964, new_n10965, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990,
    new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996,
    new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002,
    new_n11003, new_n11004, new_n11005, new_n11006, new_n11007, new_n11008,
    new_n11009, new_n11010, new_n11011, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023, new_n11024, new_n11025, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054;
  nand_5 g00000(.A(pi168), .B(pi147), .Y(new_n377));
  and_6  g00001(.A(pi236), .B(pi027), .Y(new_n378));
  not_8  g00002(.A(new_n378), .Y(new_n379));
  nand_5 g00003(.A(pi213), .B(pi164), .Y(new_n380));
  xor_4  g00004(.A(new_n380), .B(new_n379), .Y(new_n381));
  xor_4  g00005(.A(new_n381), .B(new_n377), .Y(new_n382));
  nand_5 g00006(.A(pi131), .B(pi119), .Y(new_n383));
  xor_4  g00007(.A(new_n383), .B(new_n382), .Y(po000));
  nand_5 g00008(.A(pi103), .B(pi072), .Y(new_n385));
  nand_5 g00009(.A(pi103), .B(pi044), .Y(new_n386));
  nand_5 g00010(.A(pi250), .B(pi103), .Y(new_n387));
  nand_5 g00011(.A(pi117), .B(pi045), .Y(new_n388));
  nand_5 g00012(.A(new_n388), .B(new_n387), .Y(new_n389));
  nand_5 g00013(.A(pi119), .B(pi016), .Y(new_n390));
  xor_4  g00014(.A(new_n388), .B(new_n387), .Y(new_n391));
  nand_5 g00015(.A(new_n391), .B(new_n390), .Y(new_n392));
  nand_5 g00016(.A(new_n392), .B(new_n389), .Y(new_n393));
  nor_5  g00017(.A(new_n393), .B(new_n386), .Y(new_n394));
  nand_5 g00018(.A(pi250), .B(pi117), .Y(new_n395));
  nand_5 g00019(.A(pi119), .B(pi080), .Y(new_n396));
  nand_5 g00020(.A(pi045), .B(pi016), .Y(new_n397));
  xor_4  g00021(.A(new_n397), .B(new_n396), .Y(new_n398));
  xor_4  g00022(.A(new_n398), .B(new_n395), .Y(new_n399));
  xor_4  g00023(.A(new_n393), .B(new_n386), .Y(new_n400));
  not_8  g00024(.A(new_n400), .Y(new_n401));
  nor_5  g00025(.A(new_n401), .B(new_n399), .Y(new_n402));
  nor_5  g00026(.A(new_n402), .B(new_n394), .Y(new_n403));
  nand_5 g00027(.A(pi103), .B(pi054), .Y(new_n404));
  nand_5 g00028(.A(pi250), .B(pi016), .Y(new_n405));
  nand_5 g00029(.A(pi080), .B(pi045), .Y(new_n406));
  nand_5 g00030(.A(pi247), .B(pi119), .Y(new_n407));
  xor_4  g00031(.A(new_n407), .B(new_n406), .Y(new_n408));
  xor_4  g00032(.A(new_n408), .B(new_n405), .Y(new_n409));
  nand_5 g00033(.A(new_n397), .B(new_n396), .Y(new_n410));
  nand_5 g00034(.A(new_n398), .B(new_n395), .Y(new_n411));
  nand_5 g00035(.A(new_n411), .B(new_n410), .Y(new_n412));
  nand_5 g00036(.A(pi117), .B(pi044), .Y(new_n413));
  xor_4  g00037(.A(new_n413), .B(new_n412), .Y(new_n414));
  xor_4  g00038(.A(new_n414), .B(new_n409), .Y(new_n415));
  xnor_4 g00039(.A(new_n415), .B(new_n404), .Y(new_n416));
  xor_4  g00040(.A(new_n416), .B(new_n403), .Y(new_n417));
  xor_4  g00041(.A(new_n391), .B(new_n390), .Y(new_n418));
  nand_5 g00042(.A(pi119), .B(pi103), .Y(new_n419));
  nor_5  g00043(.A(new_n419), .B(new_n388), .Y(new_n420));
  not_8  g00044(.A(new_n420), .Y(new_n421));
  or_6   g00045(.A(new_n421), .B(new_n418), .Y(new_n422));
  xor_4  g00046(.A(new_n400), .B(new_n399), .Y(new_n423));
  nor_5  g00047(.A(new_n423), .B(new_n422), .Y(new_n424));
  nand_5 g00048(.A(new_n424), .B(new_n417), .Y(new_n425));
  nand_5 g00049(.A(new_n425), .B(new_n385), .Y(new_n426));
  xor_4  g00050(.A(new_n425), .B(new_n385), .Y(new_n427));
  nor_5  g00051(.A(new_n415), .B(new_n404), .Y(new_n428));
  nor_5  g00052(.A(new_n416), .B(new_n403), .Y(new_n429));
  or_6   g00053(.A(new_n429), .B(new_n428), .Y(new_n430));
  nand_5 g00054(.A(new_n413), .B(new_n412), .Y(new_n431));
  nand_5 g00055(.A(new_n414), .B(new_n409), .Y(new_n432));
  nand_5 g00056(.A(new_n432), .B(new_n431), .Y(new_n433));
  nand_5 g00057(.A(pi117), .B(pi054), .Y(new_n434));
  nand_5 g00058(.A(pi044), .B(pi016), .Y(new_n435));
  and_6  g00059(.A(new_n435), .B(new_n434), .Y(new_n436));
  nand_5 g00060(.A(pi054), .B(pi016), .Y(new_n437));
  nor_5  g00061(.A(new_n437), .B(new_n413), .Y(new_n438));
  or_6   g00062(.A(new_n438), .B(new_n436), .Y(new_n439));
  nand_5 g00063(.A(pi247), .B(pi045), .Y(new_n440));
  nand_5 g00064(.A(pi234), .B(pi119), .Y(new_n441));
  nand_5 g00065(.A(new_n441), .B(new_n440), .Y(new_n442));
  nand_5 g00066(.A(pi234), .B(pi045), .Y(new_n443));
  nor_5  g00067(.A(new_n443), .B(new_n407), .Y(new_n444));
  not_8  g00068(.A(new_n444), .Y(new_n445));
  nand_5 g00069(.A(new_n445), .B(new_n442), .Y(new_n446));
  nand_5 g00070(.A(pi250), .B(pi080), .Y(new_n447));
  nand_5 g00071(.A(new_n407), .B(new_n406), .Y(new_n448));
  nand_5 g00072(.A(new_n408), .B(new_n405), .Y(new_n449));
  nand_5 g00073(.A(new_n449), .B(new_n448), .Y(new_n450));
  xor_4  g00074(.A(new_n450), .B(new_n447), .Y(new_n451));
  xor_4  g00075(.A(new_n451), .B(new_n446), .Y(new_n452));
  xor_4  g00076(.A(new_n452), .B(new_n439), .Y(new_n453));
  xor_4  g00077(.A(new_n453), .B(new_n433), .Y(new_n454));
  xor_4  g00078(.A(new_n454), .B(new_n430), .Y(new_n455));
  nand_5 g00079(.A(new_n455), .B(new_n427), .Y(new_n456));
  nand_5 g00080(.A(new_n456), .B(new_n426), .Y(new_n457));
  not_8  g00081(.A(new_n454), .Y(new_n458));
  nand_5 g00082(.A(new_n458), .B(new_n430), .Y(new_n459));
  not_8  g00083(.A(new_n453), .Y(new_n460));
  nor_5  g00084(.A(new_n460), .B(new_n433), .Y(new_n461));
  and_6  g00085(.A(new_n461), .B(new_n438), .Y(new_n462));
  nor_5  g00086(.A(new_n452), .B(new_n439), .Y(new_n463));
  nor_5  g00087(.A(new_n463), .B(new_n438), .Y(new_n464));
  not_8  g00088(.A(new_n464), .Y(new_n465));
  nor_5  g00089(.A(new_n465), .B(new_n461), .Y(new_n466));
  or_6   g00090(.A(new_n466), .B(new_n462), .Y(new_n467));
  nand_5 g00091(.A(pi080), .B(pi044), .Y(new_n468));
  xor_4  g00092(.A(new_n468), .B(new_n444), .Y(new_n469));
  nand_5 g00093(.A(pi250), .B(pi247), .Y(new_n470));
  nand_5 g00094(.A(pi214), .B(pi119), .Y(new_n471));
  xor_4  g00095(.A(new_n471), .B(new_n470), .Y(new_n472));
  xor_4  g00096(.A(new_n472), .B(new_n443), .Y(new_n473));
  xor_4  g00097(.A(new_n473), .B(new_n469), .Y(new_n474));
  nand_5 g00098(.A(new_n450), .B(new_n447), .Y(new_n475));
  nand_5 g00099(.A(new_n451), .B(new_n446), .Y(new_n476));
  nand_5 g00100(.A(new_n476), .B(new_n475), .Y(new_n477));
  nand_5 g00101(.A(pi248), .B(pi103), .Y(new_n478));
  nand_5 g00102(.A(pi117), .B(pi072), .Y(new_n479));
  xor_4  g00103(.A(new_n479), .B(new_n437), .Y(new_n480));
  xor_4  g00104(.A(new_n480), .B(new_n478), .Y(new_n481));
  xnor_4 g00105(.A(new_n481), .B(new_n477), .Y(new_n482));
  xor_4  g00106(.A(new_n482), .B(new_n474), .Y(new_n483));
  xor_4  g00107(.A(new_n483), .B(new_n467), .Y(new_n484));
  xor_4  g00108(.A(new_n484), .B(new_n459), .Y(new_n485));
  xnor_4 g00109(.A(new_n485), .B(new_n457), .Y(new_n486));
  nand_5 g00110(.A(pi175), .B(pi075), .Y(new_n487));
  nand_5 g00111(.A(pi151), .B(pi134), .Y(new_n488));
  not_8  g00112(.A(new_n488), .Y(new_n489));
  nand_5 g00113(.A(pi240), .B(pi147), .Y(new_n490));
  nand_5 g00114(.A(pi175), .B(pi019), .Y(new_n491));
  nor_5  g00115(.A(new_n491), .B(new_n490), .Y(new_n492));
  or_6   g00116(.A(new_n492), .B(new_n489), .Y(new_n493));
  nand_5 g00117(.A(new_n491), .B(new_n490), .Y(new_n494));
  nand_5 g00118(.A(new_n494), .B(new_n493), .Y(new_n495));
  nand_5 g00119(.A(pi175), .B(pi097), .Y(new_n496));
  nor_5  g00120(.A(new_n496), .B(new_n495), .Y(new_n497));
  nand_5 g00121(.A(pi149), .B(pi147), .Y(new_n498));
  nand_5 g00122(.A(pi134), .B(pi019), .Y(new_n499));
  nand_5 g00123(.A(pi240), .B(pi151), .Y(new_n500));
  xor_4  g00124(.A(new_n500), .B(new_n499), .Y(new_n501));
  xor_4  g00125(.A(new_n501), .B(new_n498), .Y(new_n502));
  not_8  g00126(.A(new_n502), .Y(new_n503));
  xor_4  g00127(.A(new_n496), .B(new_n495), .Y(new_n504));
  and_6  g00128(.A(new_n504), .B(new_n503), .Y(new_n505));
  nor_5  g00129(.A(new_n505), .B(new_n497), .Y(new_n506));
  xor_4  g00130(.A(new_n506), .B(new_n487), .Y(new_n507));
  nand_5 g00131(.A(pi240), .B(pi019), .Y(new_n508));
  nand_5 g00132(.A(pi167), .B(pi147), .Y(new_n509));
  nand_5 g00133(.A(pi151), .B(pi149), .Y(new_n510));
  xor_4  g00134(.A(new_n510), .B(new_n509), .Y(new_n511));
  xor_4  g00135(.A(new_n511), .B(new_n508), .Y(new_n512));
  nand_5 g00136(.A(pi134), .B(pi097), .Y(new_n513));
  nand_5 g00137(.A(new_n500), .B(new_n499), .Y(new_n514));
  nand_5 g00138(.A(new_n501), .B(new_n498), .Y(new_n515));
  nand_5 g00139(.A(new_n515), .B(new_n514), .Y(new_n516));
  xor_4  g00140(.A(new_n516), .B(new_n513), .Y(new_n517));
  xnor_4 g00141(.A(new_n517), .B(new_n512), .Y(new_n518));
  xor_4  g00142(.A(new_n518), .B(new_n507), .Y(new_n519));
  nand_5 g00143(.A(pi175), .B(pi147), .Y(new_n520));
  and_6  g00144(.A(new_n520), .B(new_n489), .Y(new_n521));
  nor_5  g00145(.A(new_n521), .B(new_n494), .Y(new_n522));
  nor_5  g00146(.A(new_n522), .B(new_n492), .Y(new_n523));
  nor_5  g00147(.A(new_n523), .B(new_n488), .Y(new_n524));
  not_8  g00148(.A(new_n524), .Y(new_n525));
  xor_4  g00149(.A(new_n504), .B(new_n502), .Y(new_n526));
  nor_5  g00150(.A(new_n526), .B(new_n525), .Y(new_n527));
  nand_5 g00151(.A(new_n527), .B(new_n519), .Y(new_n528));
  not_8  g00152(.A(new_n528), .Y(new_n529));
  nand_5 g00153(.A(pi175), .B(pi093), .Y(new_n530));
  nand_5 g00154(.A(new_n516), .B(new_n513), .Y(new_n531));
  nand_5 g00155(.A(new_n517), .B(new_n512), .Y(new_n532));
  nand_5 g00156(.A(new_n532), .B(new_n531), .Y(new_n533));
  nand_5 g00157(.A(pi240), .B(pi097), .Y(new_n534));
  nand_5 g00158(.A(pi134), .B(pi075), .Y(new_n535));
  and_6  g00159(.A(new_n535), .B(new_n534), .Y(new_n536));
  nand_5 g00160(.A(pi240), .B(pi075), .Y(new_n537));
  nor_5  g00161(.A(new_n537), .B(new_n513), .Y(new_n538));
  or_6   g00162(.A(new_n538), .B(new_n536), .Y(new_n539));
  nand_5 g00163(.A(new_n510), .B(new_n509), .Y(new_n540));
  nand_5 g00164(.A(new_n511), .B(new_n508), .Y(new_n541));
  nand_5 g00165(.A(new_n541), .B(new_n540), .Y(new_n542));
  nand_5 g00166(.A(pi149), .B(pi019), .Y(new_n543));
  nand_5 g00167(.A(pi181), .B(pi151), .Y(new_n544));
  nor_5  g00168(.A(new_n544), .B(new_n509), .Y(new_n545));
  not_8  g00169(.A(new_n545), .Y(new_n546));
  nand_5 g00170(.A(pi167), .B(pi151), .Y(new_n547));
  nand_5 g00171(.A(pi181), .B(pi147), .Y(new_n548));
  nand_5 g00172(.A(new_n548), .B(new_n547), .Y(new_n549));
  nand_5 g00173(.A(new_n549), .B(new_n546), .Y(new_n550));
  xor_4  g00174(.A(new_n550), .B(new_n543), .Y(new_n551));
  xor_4  g00175(.A(new_n551), .B(new_n542), .Y(new_n552));
  xnor_4 g00176(.A(new_n552), .B(new_n539), .Y(new_n553));
  xor_4  g00177(.A(new_n553), .B(new_n533), .Y(new_n554));
  or_6   g00178(.A(new_n506), .B(new_n487), .Y(new_n555));
  nand_5 g00179(.A(new_n518), .B(new_n507), .Y(new_n556));
  nand_5 g00180(.A(new_n556), .B(new_n555), .Y(new_n557));
  xnor_4 g00181(.A(new_n557), .B(new_n554), .Y(new_n558));
  xor_4  g00182(.A(new_n558), .B(new_n530), .Y(new_n559));
  xor_4  g00183(.A(new_n559), .B(new_n529), .Y(new_n560));
  not_8  g00184(.A(pi026), .Y(new_n561));
  not_8  g00185(.A(pi171), .Y(new_n562));
  nor_5  g00186(.A(new_n562), .B(new_n561), .Y(new_n563));
  not_8  g00187(.A(new_n563), .Y(new_n564));
  nand_5 g00188(.A(pi049), .B(pi027), .Y(new_n565));
  nand_5 g00189(.A(pi107), .B(pi008), .Y(new_n566));
  nor_5  g00190(.A(new_n566), .B(new_n565), .Y(new_n567));
  nand_5 g00191(.A(pi107), .B(pi027), .Y(new_n568));
  and_6  g00192(.A(new_n568), .B(new_n563), .Y(new_n569));
  nand_5 g00193(.A(new_n566), .B(new_n565), .Y(new_n570));
  nor_5  g00194(.A(new_n570), .B(new_n569), .Y(new_n571));
  nor_5  g00195(.A(new_n571), .B(new_n567), .Y(new_n572));
  nor_5  g00196(.A(new_n572), .B(new_n564), .Y(new_n573));
  nand_5 g00197(.A(pi245), .B(pi027), .Y(new_n574));
  nand_5 g00198(.A(pi049), .B(pi026), .Y(new_n575));
  nand_5 g00199(.A(pi171), .B(pi008), .Y(new_n576));
  xor_4  g00200(.A(new_n576), .B(new_n575), .Y(new_n577));
  xor_4  g00201(.A(new_n577), .B(new_n574), .Y(new_n578));
  or_6   g00202(.A(new_n567), .B(new_n563), .Y(new_n579));
  nand_5 g00203(.A(new_n579), .B(new_n570), .Y(new_n580));
  nand_5 g00204(.A(pi107), .B(pi056), .Y(new_n581));
  xnor_4 g00205(.A(new_n581), .B(new_n580), .Y(new_n582));
  xor_4  g00206(.A(new_n582), .B(new_n578), .Y(new_n583));
  and_6  g00207(.A(new_n583), .B(new_n573), .Y(new_n584));
  nand_5 g00208(.A(pi136), .B(pi107), .Y(new_n585));
  nor_5  g00209(.A(new_n581), .B(new_n580), .Y(new_n586));
  nor_5  g00210(.A(new_n582), .B(new_n578), .Y(new_n587));
  nor_5  g00211(.A(new_n587), .B(new_n586), .Y(new_n588));
  xor_4  g00212(.A(new_n588), .B(new_n585), .Y(new_n589));
  nand_5 g00213(.A(pi201), .B(pi027), .Y(new_n590));
  nand_5 g00214(.A(pi049), .B(pi008), .Y(new_n591));
  nand_5 g00215(.A(pi245), .B(pi026), .Y(new_n592));
  xor_4  g00216(.A(new_n592), .B(new_n591), .Y(new_n593));
  xor_4  g00217(.A(new_n593), .B(new_n590), .Y(new_n594));
  nand_5 g00218(.A(new_n576), .B(new_n575), .Y(new_n595));
  nand_5 g00219(.A(new_n577), .B(new_n574), .Y(new_n596));
  nand_5 g00220(.A(new_n596), .B(new_n595), .Y(new_n597));
  nand_5 g00221(.A(pi171), .B(pi056), .Y(new_n598));
  xor_4  g00222(.A(new_n598), .B(new_n597), .Y(new_n599));
  xnor_4 g00223(.A(new_n599), .B(new_n594), .Y(new_n600));
  xor_4  g00224(.A(new_n600), .B(new_n589), .Y(new_n601));
  xor_4  g00225(.A(new_n601), .B(new_n584), .Y(new_n602));
  nand_5 g00226(.A(new_n570), .B(new_n569), .Y(new_n603));
  nand_5 g00227(.A(new_n603), .B(new_n572), .Y(new_n604));
  nand_5 g00228(.A(pi206), .B(pi148), .Y(new_n605));
  nand_5 g00229(.A(pi164), .B(pi163), .Y(new_n606));
  or_6   g00230(.A(new_n606), .B(new_n605), .Y(new_n607));
  nand_5 g00231(.A(pi206), .B(pi163), .Y(new_n608));
  nand_5 g00232(.A(pi164), .B(pi148), .Y(new_n609));
  nand_5 g00233(.A(new_n609), .B(new_n608), .Y(new_n610));
  and_6  g00234(.A(new_n610), .B(new_n607), .Y(new_n611));
  nand_5 g00235(.A(pi107), .B(pi026), .Y(new_n612));
  nand_5 g00236(.A(pi171), .B(pi027), .Y(new_n613));
  xor_4  g00237(.A(new_n613), .B(new_n612), .Y(new_n614));
  nor_5  g00238(.A(new_n614), .B(new_n611), .Y(new_n615));
  nor_5  g00239(.A(new_n606), .B(new_n568), .Y(new_n616));
  nand_5 g00240(.A(new_n610), .B(new_n607), .Y(new_n617));
  xor_4  g00241(.A(new_n614), .B(new_n617), .Y(new_n618));
  nor_5  g00242(.A(new_n618), .B(new_n616), .Y(new_n619));
  nor_5  g00243(.A(new_n619), .B(new_n615), .Y(new_n620));
  not_8  g00244(.A(new_n620), .Y(new_n621));
  nand_5 g00245(.A(new_n621), .B(new_n604), .Y(new_n622));
  nand_5 g00246(.A(pi228), .B(pi164), .Y(new_n623));
  nand_5 g00247(.A(pi163), .B(pi032), .Y(new_n624));
  xor_4  g00248(.A(new_n624), .B(new_n605), .Y(new_n625));
  xor_4  g00249(.A(new_n625), .B(new_n623), .Y(new_n626));
  xor_4  g00250(.A(new_n626), .B(new_n607), .Y(new_n627));
  xor_4  g00251(.A(new_n620), .B(new_n604), .Y(new_n628));
  or_6   g00252(.A(new_n628), .B(new_n627), .Y(new_n629));
  nand_5 g00253(.A(new_n629), .B(new_n622), .Y(new_n630));
  xnor_4 g00254(.A(new_n583), .B(new_n573), .Y(new_n631));
  and_6  g00255(.A(new_n631), .B(new_n630), .Y(new_n632));
  nor_5  g00256(.A(new_n626), .B(new_n607), .Y(new_n633));
  nand_5 g00257(.A(pi228), .B(pi206), .Y(new_n634));
  nand_5 g00258(.A(pi148), .B(pi032), .Y(new_n635));
  nand_5 g00259(.A(pi164), .B(pi039), .Y(new_n636));
  xor_4  g00260(.A(new_n636), .B(new_n635), .Y(new_n637));
  xor_4  g00261(.A(new_n637), .B(new_n634), .Y(new_n638));
  nand_5 g00262(.A(pi163), .B(pi145), .Y(new_n639));
  nand_5 g00263(.A(new_n624), .B(new_n605), .Y(new_n640));
  nand_5 g00264(.A(new_n625), .B(new_n623), .Y(new_n641));
  nand_5 g00265(.A(new_n641), .B(new_n640), .Y(new_n642));
  xor_4  g00266(.A(new_n642), .B(new_n639), .Y(new_n643));
  xnor_4 g00267(.A(new_n643), .B(new_n638), .Y(new_n644));
  xor_4  g00268(.A(new_n644), .B(new_n633), .Y(new_n645));
  xnor_4 g00269(.A(new_n631), .B(new_n630), .Y(new_n646));
  nor_5  g00270(.A(new_n646), .B(new_n645), .Y(new_n647));
  nor_5  g00271(.A(new_n647), .B(new_n632), .Y(new_n648));
  nor_5  g00272(.A(new_n648), .B(new_n602), .Y(new_n649));
  and_6  g00273(.A(new_n644), .B(new_n633), .Y(new_n650));
  nand_5 g00274(.A(pi246), .B(pi163), .Y(new_n651));
  nand_5 g00275(.A(new_n642), .B(new_n639), .Y(new_n652));
  nand_5 g00276(.A(new_n643), .B(new_n638), .Y(new_n653));
  nand_5 g00277(.A(new_n653), .B(new_n652), .Y(new_n654));
  xor_4  g00278(.A(new_n654), .B(new_n651), .Y(new_n655));
  nand_5 g00279(.A(pi164), .B(pi116), .Y(new_n656));
  nand_5 g00280(.A(pi228), .B(pi032), .Y(new_n657));
  nand_5 g00281(.A(pi206), .B(pi039), .Y(new_n658));
  xor_4  g00282(.A(new_n658), .B(new_n657), .Y(new_n659));
  xor_4  g00283(.A(new_n659), .B(new_n656), .Y(new_n660));
  nand_5 g00284(.A(new_n636), .B(new_n635), .Y(new_n661));
  nand_5 g00285(.A(new_n637), .B(new_n634), .Y(new_n662));
  nand_5 g00286(.A(new_n662), .B(new_n661), .Y(new_n663));
  nand_5 g00287(.A(pi148), .B(pi145), .Y(new_n664));
  xnor_4 g00288(.A(new_n664), .B(new_n663), .Y(new_n665));
  xor_4  g00289(.A(new_n665), .B(new_n660), .Y(new_n666));
  xor_4  g00290(.A(new_n666), .B(new_n655), .Y(new_n667));
  xor_4  g00291(.A(new_n667), .B(new_n650), .Y(new_n668));
  xnor_4 g00292(.A(new_n648), .B(new_n602), .Y(new_n669));
  nor_5  g00293(.A(new_n669), .B(new_n668), .Y(new_n670));
  nor_5  g00294(.A(new_n670), .B(new_n649), .Y(new_n671));
  or_6   g00295(.A(new_n588), .B(new_n585), .Y(new_n672));
  nand_5 g00296(.A(new_n600), .B(new_n589), .Y(new_n673));
  nand_5 g00297(.A(new_n673), .B(new_n672), .Y(new_n674));
  nand_5 g00298(.A(new_n592), .B(new_n591), .Y(new_n675));
  nand_5 g00299(.A(new_n593), .B(new_n590), .Y(new_n676));
  nand_5 g00300(.A(new_n676), .B(new_n675), .Y(new_n677));
  nand_5 g00301(.A(pi245), .B(pi008), .Y(new_n678));
  nand_5 g00302(.A(pi156), .B(pi027), .Y(new_n679));
  nand_5 g00303(.A(pi201), .B(pi026), .Y(new_n680));
  nand_5 g00304(.A(new_n680), .B(new_n679), .Y(new_n681));
  nand_5 g00305(.A(pi156), .B(pi026), .Y(new_n682));
  nor_5  g00306(.A(new_n682), .B(new_n590), .Y(new_n683));
  not_8  g00307(.A(new_n683), .Y(new_n684));
  nand_5 g00308(.A(new_n684), .B(new_n681), .Y(new_n685));
  xor_4  g00309(.A(new_n685), .B(new_n678), .Y(new_n686));
  xor_4  g00310(.A(new_n686), .B(new_n677), .Y(new_n687));
  nand_5 g00311(.A(new_n598), .B(new_n597), .Y(new_n688));
  nand_5 g00312(.A(new_n599), .B(new_n594), .Y(new_n689));
  nand_5 g00313(.A(new_n689), .B(new_n688), .Y(new_n690));
  nand_5 g00314(.A(pi056), .B(pi049), .Y(new_n691));
  nand_5 g00315(.A(pi171), .B(pi136), .Y(new_n692));
  nand_5 g00316(.A(new_n692), .B(new_n691), .Y(new_n693));
  nand_5 g00317(.A(pi136), .B(pi049), .Y(new_n694));
  nor_5  g00318(.A(new_n694), .B(new_n598), .Y(new_n695));
  not_8  g00319(.A(new_n695), .Y(new_n696));
  nand_5 g00320(.A(new_n696), .B(new_n693), .Y(new_n697));
  xor_4  g00321(.A(new_n697), .B(new_n690), .Y(new_n698));
  xnor_4 g00322(.A(new_n698), .B(new_n687), .Y(new_n699));
  xor_4  g00323(.A(new_n699), .B(new_n674), .Y(new_n700));
  nand_5 g00324(.A(new_n601), .B(new_n584), .Y(new_n701));
  nand_5 g00325(.A(pi107), .B(pi096), .Y(new_n702));
  xnor_4 g00326(.A(new_n702), .B(new_n701), .Y(new_n703));
  xor_4  g00327(.A(new_n703), .B(new_n700), .Y(new_n704));
  or_6   g00328(.A(new_n654), .B(new_n651), .Y(new_n705));
  nand_5 g00329(.A(new_n666), .B(new_n655), .Y(new_n706));
  and_6  g00330(.A(new_n706), .B(new_n705), .Y(new_n707));
  nand_5 g00331(.A(pi039), .B(pi032), .Y(new_n708));
  nand_5 g00332(.A(pi206), .B(pi116), .Y(new_n709));
  nand_5 g00333(.A(pi164), .B(pi070), .Y(new_n710));
  nand_5 g00334(.A(new_n710), .B(new_n709), .Y(new_n711));
  nand_5 g00335(.A(pi206), .B(pi070), .Y(new_n712));
  nor_5  g00336(.A(new_n712), .B(new_n656), .Y(new_n713));
  not_8  g00337(.A(new_n713), .Y(new_n714));
  nand_5 g00338(.A(new_n714), .B(new_n711), .Y(new_n715));
  xor_4  g00339(.A(new_n715), .B(new_n708), .Y(new_n716));
  nand_5 g00340(.A(new_n658), .B(new_n657), .Y(new_n717));
  nand_5 g00341(.A(new_n659), .B(new_n656), .Y(new_n718));
  nand_5 g00342(.A(new_n718), .B(new_n717), .Y(new_n719));
  xor_4  g00343(.A(new_n719), .B(new_n716), .Y(new_n720));
  nand_5 g00344(.A(pi228), .B(pi145), .Y(new_n721));
  nand_5 g00345(.A(pi246), .B(pi148), .Y(new_n722));
  and_6  g00346(.A(new_n722), .B(new_n721), .Y(new_n723));
  nand_5 g00347(.A(pi246), .B(pi228), .Y(new_n724));
  nor_5  g00348(.A(new_n724), .B(new_n664), .Y(new_n725));
  or_6   g00349(.A(new_n725), .B(new_n723), .Y(new_n726));
  xnor_4 g00350(.A(new_n726), .B(new_n720), .Y(new_n727));
  nand_5 g00351(.A(new_n664), .B(new_n663), .Y(new_n728));
  not_8  g00352(.A(new_n660), .Y(new_n729));
  or_6   g00353(.A(new_n665), .B(new_n729), .Y(new_n730));
  nand_5 g00354(.A(new_n730), .B(new_n728), .Y(new_n731));
  xnor_4 g00355(.A(new_n731), .B(new_n727), .Y(new_n732));
  xnor_4 g00356(.A(new_n732), .B(new_n707), .Y(new_n733));
  nand_5 g00357(.A(new_n667), .B(new_n650), .Y(new_n734));
  nand_5 g00358(.A(pi163), .B(pi114), .Y(new_n735));
  xor_4  g00359(.A(new_n735), .B(new_n734), .Y(new_n736));
  xor_4  g00360(.A(new_n736), .B(new_n733), .Y(new_n737));
  xor_4  g00361(.A(new_n737), .B(new_n704), .Y(new_n738));
  xor_4  g00362(.A(new_n738), .B(new_n671), .Y(new_n739));
  nand_5 g00363(.A(new_n739), .B(new_n560), .Y(new_n740));
  xor_4  g00364(.A(new_n527), .B(new_n519), .Y(new_n741));
  not_8  g00365(.A(new_n741), .Y(new_n742));
  nand_5 g00366(.A(new_n521), .B(new_n494), .Y(new_n743));
  nand_5 g00367(.A(new_n743), .B(new_n523), .Y(new_n744));
  not_8  g00368(.A(new_n744), .Y(new_n745));
  not_8  g00369(.A(new_n627), .Y(new_n746));
  xor_4  g00370(.A(new_n628), .B(new_n746), .Y(new_n747));
  and_6  g00371(.A(new_n747), .B(new_n745), .Y(new_n748));
  nand_5 g00372(.A(pi175), .B(pi151), .Y(new_n749));
  nand_5 g00373(.A(pi147), .B(pi134), .Y(new_n750));
  xor_4  g00374(.A(new_n750), .B(new_n749), .Y(new_n751));
  xnor_4 g00375(.A(new_n606), .B(new_n568), .Y(new_n752));
  nor_5  g00376(.A(new_n752), .B(new_n520), .Y(new_n753));
  and_6  g00377(.A(new_n753), .B(new_n751), .Y(new_n754));
  xor_4  g00378(.A(new_n618), .B(new_n616), .Y(new_n755));
  xnor_4 g00379(.A(new_n753), .B(new_n751), .Y(new_n756));
  nor_5  g00380(.A(new_n756), .B(new_n755), .Y(new_n757));
  nor_5  g00381(.A(new_n757), .B(new_n754), .Y(new_n758));
  xor_4  g00382(.A(new_n747), .B(new_n744), .Y(new_n759));
  nor_5  g00383(.A(new_n759), .B(new_n758), .Y(new_n760));
  nor_5  g00384(.A(new_n760), .B(new_n748), .Y(new_n761));
  xor_4  g00385(.A(new_n526), .B(new_n524), .Y(new_n762));
  nor_5  g00386(.A(new_n762), .B(new_n761), .Y(new_n763));
  xor_4  g00387(.A(new_n762), .B(new_n761), .Y(new_n764));
  xnor_4 g00388(.A(new_n646), .B(new_n645), .Y(new_n765));
  and_6  g00389(.A(new_n765), .B(new_n764), .Y(new_n766));
  nor_5  g00390(.A(new_n766), .B(new_n763), .Y(new_n767));
  nor_5  g00391(.A(new_n767), .B(new_n742), .Y(new_n768));
  xor_4  g00392(.A(new_n669), .B(new_n668), .Y(new_n769));
  xor_4  g00393(.A(new_n767), .B(new_n741), .Y(new_n770));
  nor_5  g00394(.A(new_n770), .B(new_n769), .Y(new_n771));
  nor_5  g00395(.A(new_n771), .B(new_n768), .Y(new_n772));
  xnor_4 g00396(.A(new_n739), .B(new_n560), .Y(new_n773));
  or_6   g00397(.A(new_n773), .B(new_n772), .Y(new_n774));
  nand_5 g00398(.A(new_n774), .B(new_n740), .Y(new_n775));
  nand_5 g00399(.A(new_n702), .B(new_n701), .Y(new_n776));
  or_6   g00400(.A(new_n703), .B(new_n700), .Y(new_n777));
  nand_5 g00401(.A(new_n777), .B(new_n776), .Y(new_n778));
  and_6  g00402(.A(new_n699), .B(new_n674), .Y(new_n779));
  nand_5 g00403(.A(new_n685), .B(new_n678), .Y(new_n780));
  nand_5 g00404(.A(new_n686), .B(new_n677), .Y(new_n781));
  nand_5 g00405(.A(new_n781), .B(new_n780), .Y(new_n782));
  nand_5 g00406(.A(pi171), .B(pi096), .Y(new_n783));
  nand_5 g00407(.A(pi235), .B(pi107), .Y(new_n784));
  xor_4  g00408(.A(new_n784), .B(new_n783), .Y(new_n785));
  xor_4  g00409(.A(new_n785), .B(new_n694), .Y(new_n786));
  xor_4  g00410(.A(new_n786), .B(new_n782), .Y(new_n787));
  nand_5 g00411(.A(pi245), .B(pi056), .Y(new_n788));
  xor_4  g00412(.A(new_n788), .B(new_n684), .Y(new_n789));
  nand_5 g00413(.A(pi201), .B(pi008), .Y(new_n790));
  nand_5 g00414(.A(pi063), .B(pi027), .Y(new_n791));
  xor_4  g00415(.A(new_n791), .B(new_n790), .Y(new_n792));
  xor_4  g00416(.A(new_n792), .B(new_n682), .Y(new_n793));
  xor_4  g00417(.A(new_n793), .B(new_n789), .Y(new_n794));
  xnor_4 g00418(.A(new_n794), .B(new_n787), .Y(new_n795));
  nand_5 g00419(.A(new_n697), .B(new_n690), .Y(new_n796));
  nand_5 g00420(.A(new_n698), .B(new_n687), .Y(new_n797));
  nand_5 g00421(.A(new_n797), .B(new_n796), .Y(new_n798));
  xor_4  g00422(.A(new_n798), .B(new_n696), .Y(new_n799));
  xor_4  g00423(.A(new_n799), .B(new_n795), .Y(new_n800));
  xnor_4 g00424(.A(new_n800), .B(new_n779), .Y(new_n801));
  xor_4  g00425(.A(new_n801), .B(new_n778), .Y(new_n802));
  nand_5 g00426(.A(new_n735), .B(new_n734), .Y(new_n803));
  nand_5 g00427(.A(new_n736), .B(new_n733), .Y(new_n804));
  nand_5 g00428(.A(new_n804), .B(new_n803), .Y(new_n805));
  or_6   g00429(.A(new_n732), .B(new_n707), .Y(new_n806));
  not_8  g00430(.A(new_n806), .Y(new_n807));
  nand_5 g00431(.A(pi148), .B(pi114), .Y(new_n808));
  nand_5 g00432(.A(pi163), .B(pi091), .Y(new_n809));
  xor_4  g00433(.A(new_n809), .B(new_n808), .Y(new_n810));
  xor_4  g00434(.A(new_n810), .B(new_n724), .Y(new_n811));
  nand_5 g00435(.A(new_n715), .B(new_n708), .Y(new_n812));
  nand_5 g00436(.A(new_n719), .B(new_n716), .Y(new_n813));
  nand_5 g00437(.A(new_n813), .B(new_n812), .Y(new_n814));
  xor_4  g00438(.A(new_n814), .B(new_n811), .Y(new_n815));
  nand_5 g00439(.A(pi164), .B(pi115), .Y(new_n816));
  nand_5 g00440(.A(pi116), .B(pi032), .Y(new_n817));
  xor_4  g00441(.A(new_n817), .B(new_n816), .Y(new_n818));
  xor_4  g00442(.A(new_n818), .B(new_n712), .Y(new_n819));
  nand_5 g00443(.A(pi145), .B(pi039), .Y(new_n820));
  xor_4  g00444(.A(new_n820), .B(new_n713), .Y(new_n821));
  xnor_4 g00445(.A(new_n821), .B(new_n819), .Y(new_n822));
  xnor_4 g00446(.A(new_n822), .B(new_n815), .Y(new_n823));
  nor_5  g00447(.A(new_n726), .B(new_n720), .Y(new_n824));
  nor_5  g00448(.A(new_n731), .B(new_n727), .Y(new_n825));
  xor_4  g00449(.A(new_n825), .B(new_n725), .Y(new_n826));
  nor_5  g00450(.A(new_n826), .B(new_n824), .Y(new_n827));
  not_8  g00451(.A(new_n827), .Y(new_n828));
  xor_4  g00452(.A(new_n828), .B(new_n823), .Y(new_n829));
  or_6   g00453(.A(new_n829), .B(new_n807), .Y(new_n830));
  nand_5 g00454(.A(new_n829), .B(new_n807), .Y(new_n831));
  nand_5 g00455(.A(new_n831), .B(new_n830), .Y(new_n832));
  xor_4  g00456(.A(new_n832), .B(new_n805), .Y(new_n833));
  xor_4  g00457(.A(new_n833), .B(new_n802), .Y(new_n834));
  nand_5 g00458(.A(new_n737), .B(new_n704), .Y(new_n835));
  nor_5  g00459(.A(new_n737), .B(new_n704), .Y(new_n836));
  or_6   g00460(.A(new_n836), .B(new_n671), .Y(new_n837));
  and_6  g00461(.A(new_n837), .B(new_n835), .Y(new_n838));
  xor_4  g00462(.A(new_n838), .B(new_n834), .Y(new_n839));
  nand_5 g00463(.A(new_n557), .B(new_n554), .Y(new_n840));
  nor_5  g00464(.A(new_n552), .B(new_n539), .Y(new_n841));
  nor_5  g00465(.A(new_n553), .B(new_n533), .Y(new_n842));
  xor_4  g00466(.A(new_n842), .B(new_n538), .Y(new_n843));
  nor_5  g00467(.A(new_n843), .B(new_n841), .Y(new_n844));
  nand_5 g00468(.A(new_n550), .B(new_n543), .Y(new_n845));
  nand_5 g00469(.A(new_n551), .B(new_n542), .Y(new_n846));
  nand_5 g00470(.A(new_n846), .B(new_n845), .Y(new_n847));
  nand_5 g00471(.A(pi134), .B(pi093), .Y(new_n848));
  nand_5 g00472(.A(pi175), .B(pi166), .Y(new_n849));
  xor_4  g00473(.A(new_n849), .B(new_n848), .Y(new_n850));
  xor_4  g00474(.A(new_n850), .B(new_n537), .Y(new_n851));
  xor_4  g00475(.A(new_n851), .B(new_n847), .Y(new_n852));
  nand_5 g00476(.A(pi149), .B(pi097), .Y(new_n853));
  xor_4  g00477(.A(new_n853), .B(new_n546), .Y(new_n854));
  nand_5 g00478(.A(pi167), .B(pi019), .Y(new_n855));
  nand_5 g00479(.A(pi200), .B(pi147), .Y(new_n856));
  xor_4  g00480(.A(new_n856), .B(new_n855), .Y(new_n857));
  xnor_4 g00481(.A(new_n857), .B(new_n544), .Y(new_n858));
  xnor_4 g00482(.A(new_n858), .B(new_n854), .Y(new_n859));
  xor_4  g00483(.A(new_n859), .B(new_n852), .Y(new_n860));
  xor_4  g00484(.A(new_n860), .B(new_n844), .Y(new_n861));
  xor_4  g00485(.A(new_n861), .B(new_n840), .Y(new_n862));
  nor_5  g00486(.A(new_n558), .B(new_n530), .Y(new_n863));
  and_6  g00487(.A(new_n559), .B(new_n529), .Y(new_n864));
  nor_5  g00488(.A(new_n864), .B(new_n863), .Y(new_n865));
  xor_4  g00489(.A(new_n865), .B(new_n862), .Y(new_n866));
  xnor_4 g00490(.A(new_n866), .B(new_n839), .Y(new_n867));
  xor_4  g00491(.A(new_n867), .B(new_n775), .Y(new_n868));
  xor_4  g00492(.A(new_n868), .B(new_n486), .Y(new_n869));
  xor_4  g00493(.A(new_n765), .B(new_n764), .Y(new_n870));
  xor_4  g00494(.A(new_n423), .B(new_n422), .Y(new_n871));
  or_6   g00495(.A(new_n871), .B(new_n870), .Y(new_n872));
  xor_4  g00496(.A(new_n871), .B(new_n870), .Y(new_n873));
  xor_4  g00497(.A(new_n421), .B(new_n418), .Y(new_n874));
  not_8  g00498(.A(new_n874), .Y(new_n875));
  xnor_4 g00499(.A(new_n752), .B(new_n520), .Y(new_n876));
  or_6   g00500(.A(new_n876), .B(new_n419), .Y(new_n877));
  nand_5 g00501(.A(pi103), .B(pi045), .Y(new_n878));
  nand_5 g00502(.A(pi119), .B(pi117), .Y(new_n879));
  nand_5 g00503(.A(new_n879), .B(new_n878), .Y(new_n880));
  nand_5 g00504(.A(new_n880), .B(new_n421), .Y(new_n881));
  nand_5 g00505(.A(new_n881), .B(new_n877), .Y(new_n882));
  xnor_4 g00506(.A(new_n756), .B(new_n755), .Y(new_n883));
  xor_4  g00507(.A(new_n881), .B(new_n877), .Y(new_n884));
  nand_5 g00508(.A(new_n884), .B(new_n883), .Y(new_n885));
  nand_5 g00509(.A(new_n885), .B(new_n882), .Y(new_n886));
  nand_5 g00510(.A(new_n886), .B(new_n875), .Y(new_n887));
  xor_4  g00511(.A(new_n886), .B(new_n875), .Y(new_n888));
  xnor_4 g00512(.A(new_n759), .B(new_n758), .Y(new_n889));
  nand_5 g00513(.A(new_n889), .B(new_n888), .Y(new_n890));
  nand_5 g00514(.A(new_n890), .B(new_n887), .Y(new_n891));
  nand_5 g00515(.A(new_n891), .B(new_n873), .Y(new_n892));
  nand_5 g00516(.A(new_n892), .B(new_n872), .Y(new_n893));
  xor_4  g00517(.A(new_n424), .B(new_n417), .Y(new_n894));
  not_8  g00518(.A(new_n894), .Y(new_n895));
  or_6   g00519(.A(new_n895), .B(new_n893), .Y(new_n896));
  xor_4  g00520(.A(new_n770), .B(new_n769), .Y(new_n897));
  xor_4  g00521(.A(new_n895), .B(new_n893), .Y(new_n898));
  nand_5 g00522(.A(new_n898), .B(new_n897), .Y(new_n899));
  and_6  g00523(.A(new_n899), .B(new_n896), .Y(new_n900));
  xor_4  g00524(.A(new_n455), .B(new_n427), .Y(new_n901));
  nand_5 g00525(.A(new_n901), .B(new_n900), .Y(new_n902));
  xor_4  g00526(.A(new_n901), .B(new_n900), .Y(new_n903));
  xnor_4 g00527(.A(new_n773), .B(new_n772), .Y(new_n904));
  nand_5 g00528(.A(new_n904), .B(new_n903), .Y(new_n905));
  nand_5 g00529(.A(new_n905), .B(new_n902), .Y(new_n906));
  xnor_4 g00530(.A(new_n906), .B(new_n869), .Y(po001));
  nand_5 g00531(.A(pi134), .B(pi033), .Y(new_n908));
  not_8  g00532(.A(new_n908), .Y(new_n909));
  nand_5 g00533(.A(pi175), .B(pi162), .Y(new_n910));
  and_6  g00534(.A(new_n910), .B(new_n909), .Y(new_n911));
  nand_5 g00535(.A(pi179), .B(pi175), .Y(new_n912));
  nand_5 g00536(.A(pi240), .B(pi162), .Y(new_n913));
  nand_5 g00537(.A(new_n913), .B(new_n912), .Y(new_n914));
  nor_5  g00538(.A(new_n914), .B(new_n911), .Y(new_n915));
  nor_5  g00539(.A(new_n913), .B(new_n912), .Y(new_n916));
  nor_5  g00540(.A(new_n916), .B(new_n915), .Y(new_n917));
  nor_5  g00541(.A(new_n917), .B(new_n908), .Y(new_n918));
  nand_5 g00542(.A(pi179), .B(pi134), .Y(new_n919));
  nand_5 g00543(.A(pi162), .B(pi149), .Y(new_n920));
  nand_5 g00544(.A(pi240), .B(pi033), .Y(new_n921));
  xor_4  g00545(.A(new_n921), .B(new_n920), .Y(new_n922));
  xor_4  g00546(.A(new_n922), .B(new_n919), .Y(new_n923));
  not_8  g00547(.A(new_n914), .Y(new_n924));
  nor_5  g00548(.A(new_n916), .B(new_n909), .Y(new_n925));
  nor_5  g00549(.A(new_n925), .B(new_n924), .Y(new_n926));
  nand_5 g00550(.A(pi175), .B(pi048), .Y(new_n927));
  xor_4  g00551(.A(new_n927), .B(new_n926), .Y(new_n928));
  xor_4  g00552(.A(new_n928), .B(new_n923), .Y(new_n929));
  xor_4  g00553(.A(new_n929), .B(new_n918), .Y(new_n930));
  nand_5 g00554(.A(pi107), .B(pi051), .Y(new_n931));
  nand_5 g00555(.A(pi171), .B(pi042), .Y(new_n932));
  nor_5  g00556(.A(new_n932), .B(new_n931), .Y(new_n933));
  nand_5 g00557(.A(pi171), .B(pi051), .Y(new_n934));
  nand_5 g00558(.A(pi107), .B(pi042), .Y(new_n935));
  and_6  g00559(.A(new_n935), .B(new_n934), .Y(new_n936));
  or_6   g00560(.A(new_n936), .B(new_n933), .Y(new_n937));
  nand_5 g00561(.A(pi188), .B(pi163), .Y(new_n938));
  nand_5 g00562(.A(pi178), .B(pi148), .Y(new_n939));
  nor_5  g00563(.A(new_n939), .B(new_n938), .Y(new_n940));
  nand_5 g00564(.A(pi188), .B(pi148), .Y(new_n941));
  nand_5 g00565(.A(pi178), .B(pi163), .Y(new_n942));
  and_6  g00566(.A(new_n942), .B(new_n941), .Y(new_n943));
  or_6   g00567(.A(new_n943), .B(new_n940), .Y(new_n944));
  nand_5 g00568(.A(new_n944), .B(new_n937), .Y(new_n945));
  or_6   g00569(.A(new_n938), .B(new_n931), .Y(new_n946));
  xor_4  g00570(.A(new_n944), .B(new_n937), .Y(new_n947));
  nand_5 g00571(.A(new_n947), .B(new_n946), .Y(new_n948));
  nand_5 g00572(.A(new_n948), .B(new_n945), .Y(new_n949));
  nand_5 g00573(.A(pi051), .B(pi049), .Y(new_n950));
  nand_5 g00574(.A(pi108), .B(pi107), .Y(new_n951));
  xor_4  g00575(.A(new_n951), .B(new_n932), .Y(new_n952));
  xor_4  g00576(.A(new_n952), .B(new_n950), .Y(new_n953));
  xor_4  g00577(.A(new_n953), .B(new_n933), .Y(new_n954));
  nand_5 g00578(.A(pi228), .B(pi188), .Y(new_n955));
  nand_5 g00579(.A(pi163), .B(pi061), .Y(new_n956));
  xor_4  g00580(.A(new_n956), .B(new_n939), .Y(new_n957));
  xnor_4 g00581(.A(new_n957), .B(new_n955), .Y(new_n958));
  xor_4  g00582(.A(new_n958), .B(new_n940), .Y(new_n959));
  xor_4  g00583(.A(new_n959), .B(new_n954), .Y(new_n960));
  xnor_4 g00584(.A(new_n960), .B(new_n949), .Y(new_n961));
  nand_5 g00585(.A(new_n914), .B(new_n911), .Y(new_n962));
  nand_5 g00586(.A(new_n962), .B(new_n917), .Y(new_n963));
  or_6   g00587(.A(new_n963), .B(new_n961), .Y(new_n964));
  xnor_4 g00588(.A(new_n938), .B(new_n931), .Y(new_n965));
  nor_5  g00589(.A(new_n965), .B(new_n910), .Y(new_n966));
  nand_5 g00590(.A(pi162), .B(pi134), .Y(new_n967));
  nand_5 g00591(.A(pi175), .B(pi033), .Y(new_n968));
  xor_4  g00592(.A(new_n968), .B(new_n967), .Y(new_n969));
  nand_5 g00593(.A(new_n969), .B(new_n966), .Y(new_n970));
  xnor_4 g00594(.A(new_n947), .B(new_n946), .Y(new_n971));
  xor_4  g00595(.A(new_n969), .B(new_n966), .Y(new_n972));
  nand_5 g00596(.A(new_n972), .B(new_n971), .Y(new_n973));
  nand_5 g00597(.A(new_n973), .B(new_n970), .Y(new_n974));
  nand_5 g00598(.A(new_n963), .B(new_n961), .Y(new_n975));
  nand_5 g00599(.A(new_n975), .B(new_n974), .Y(new_n976));
  nand_5 g00600(.A(new_n976), .B(new_n964), .Y(new_n977));
  xor_4  g00601(.A(new_n977), .B(new_n930), .Y(new_n978));
  not_8  g00602(.A(new_n959), .Y(new_n979));
  nor_5  g00603(.A(new_n979), .B(new_n954), .Y(new_n980));
  nor_5  g00604(.A(new_n960), .B(new_n949), .Y(new_n981));
  or_6   g00605(.A(new_n981), .B(new_n980), .Y(new_n982));
  not_8  g00606(.A(new_n953), .Y(new_n983));
  nand_5 g00607(.A(new_n983), .B(new_n933), .Y(new_n984));
  nand_5 g00608(.A(pi171), .B(pi108), .Y(new_n985));
  nand_5 g00609(.A(pi245), .B(pi051), .Y(new_n986));
  nand_5 g00610(.A(pi049), .B(pi042), .Y(new_n987));
  xor_4  g00611(.A(new_n987), .B(new_n986), .Y(new_n988));
  xor_4  g00612(.A(new_n988), .B(new_n985), .Y(new_n989));
  nand_5 g00613(.A(pi107), .B(pi007), .Y(new_n990));
  nand_5 g00614(.A(new_n951), .B(new_n932), .Y(new_n991));
  nand_5 g00615(.A(new_n952), .B(new_n950), .Y(new_n992));
  nand_5 g00616(.A(new_n992), .B(new_n991), .Y(new_n993));
  xnor_4 g00617(.A(new_n993), .B(new_n990), .Y(new_n994));
  xnor_4 g00618(.A(new_n994), .B(new_n989), .Y(new_n995));
  xor_4  g00619(.A(new_n995), .B(new_n984), .Y(new_n996));
  nand_5 g00620(.A(new_n958), .B(new_n940), .Y(new_n997));
  nand_5 g00621(.A(pi148), .B(pi061), .Y(new_n998));
  nand_5 g00622(.A(pi188), .B(pi039), .Y(new_n999));
  nand_5 g00623(.A(pi228), .B(pi178), .Y(new_n1000));
  xor_4  g00624(.A(new_n1000), .B(new_n999), .Y(new_n1001));
  xor_4  g00625(.A(new_n1001), .B(new_n998), .Y(new_n1002));
  nand_5 g00626(.A(pi163), .B(pi012), .Y(new_n1003));
  nand_5 g00627(.A(new_n956), .B(new_n939), .Y(new_n1004));
  nand_5 g00628(.A(new_n957), .B(new_n955), .Y(new_n1005));
  nand_5 g00629(.A(new_n1005), .B(new_n1004), .Y(new_n1006));
  xor_4  g00630(.A(new_n1006), .B(new_n1003), .Y(new_n1007));
  xor_4  g00631(.A(new_n1007), .B(new_n1002), .Y(new_n1008));
  xor_4  g00632(.A(new_n1008), .B(new_n997), .Y(new_n1009));
  xor_4  g00633(.A(new_n1009), .B(new_n996), .Y(new_n1010));
  xnor_4 g00634(.A(new_n1010), .B(new_n982), .Y(new_n1011));
  xor_4  g00635(.A(new_n1011), .B(new_n978), .Y(new_n1012));
  nand_5 g00636(.A(pi143), .B(pi016), .Y(new_n1013));
  nand_5 g00637(.A(pi117), .B(pi057), .Y(new_n1014));
  nand_5 g00638(.A(pi194), .B(pi103), .Y(new_n1015));
  xor_4  g00639(.A(new_n1015), .B(new_n1014), .Y(new_n1016));
  xor_4  g00640(.A(new_n1016), .B(new_n1013), .Y(new_n1017));
  nand_5 g00641(.A(pi143), .B(pi103), .Y(new_n1018));
  or_6   g00642(.A(new_n1018), .B(new_n1014), .Y(new_n1019));
  or_6   g00643(.A(new_n1019), .B(new_n1017), .Y(new_n1020));
  not_8  g00644(.A(new_n1020), .Y(new_n1021));
  nand_5 g00645(.A(pi143), .B(pi080), .Y(new_n1022));
  nand_5 g00646(.A(pi194), .B(pi117), .Y(new_n1023));
  nand_5 g00647(.A(pi057), .B(pi016), .Y(new_n1024));
  xor_4  g00648(.A(new_n1024), .B(new_n1023), .Y(new_n1025));
  xor_4  g00649(.A(new_n1025), .B(new_n1022), .Y(new_n1026));
  nand_5 g00650(.A(pi103), .B(pi085), .Y(new_n1027));
  nand_5 g00651(.A(new_n1015), .B(new_n1014), .Y(new_n1028));
  nand_5 g00652(.A(new_n1016), .B(new_n1013), .Y(new_n1029));
  nand_5 g00653(.A(new_n1029), .B(new_n1028), .Y(new_n1030));
  xor_4  g00654(.A(new_n1030), .B(new_n1027), .Y(new_n1031));
  xor_4  g00655(.A(new_n1031), .B(new_n1026), .Y(new_n1032));
  xor_4  g00656(.A(new_n1032), .B(new_n1021), .Y(new_n1033));
  xnor_4 g00657(.A(new_n965), .B(new_n910), .Y(new_n1034));
  or_6   g00658(.A(new_n1034), .B(new_n1018), .Y(new_n1035));
  nand_5 g00659(.A(pi103), .B(pi057), .Y(new_n1036));
  nand_5 g00660(.A(pi143), .B(pi117), .Y(new_n1037));
  nand_5 g00661(.A(new_n1037), .B(new_n1036), .Y(new_n1038));
  nand_5 g00662(.A(new_n1038), .B(new_n1019), .Y(new_n1039));
  nand_5 g00663(.A(new_n1039), .B(new_n1035), .Y(new_n1040));
  xnor_4 g00664(.A(new_n972), .B(new_n971), .Y(new_n1041));
  xor_4  g00665(.A(new_n1039), .B(new_n1035), .Y(new_n1042));
  nand_5 g00666(.A(new_n1042), .B(new_n1041), .Y(new_n1043));
  nand_5 g00667(.A(new_n1043), .B(new_n1040), .Y(new_n1044));
  xnor_4 g00668(.A(new_n1019), .B(new_n1017), .Y(new_n1045));
  nor_5  g00669(.A(new_n1045), .B(new_n1044), .Y(new_n1046));
  nand_5 g00670(.A(new_n975), .B(new_n964), .Y(new_n1047));
  xor_4  g00671(.A(new_n1047), .B(new_n974), .Y(new_n1048));
  xnor_4 g00672(.A(new_n1045), .B(new_n1044), .Y(new_n1049));
  nor_5  g00673(.A(new_n1049), .B(new_n1048), .Y(new_n1050));
  nor_5  g00674(.A(new_n1050), .B(new_n1046), .Y(new_n1051));
  xnor_4 g00675(.A(new_n1051), .B(new_n1033), .Y(new_n1052));
  xor_4  g00676(.A(new_n1052), .B(new_n1012), .Y(po002));
  nand_5 g00677(.A(pi160), .B(pi119), .Y(new_n1054));
  nand_5 g00678(.A(pi147), .B(pi138), .Y(new_n1055));
  nand_5 g00679(.A(pi087), .B(pi027), .Y(new_n1056));
  nand_5 g00680(.A(pi164), .B(pi142), .Y(new_n1057));
  xor_4  g00681(.A(new_n1057), .B(new_n1056), .Y(new_n1058));
  xor_4  g00682(.A(new_n1058), .B(new_n1055), .Y(new_n1059));
  xor_4  g00683(.A(new_n1059), .B(new_n1054), .Y(po003));
  nand_5 g00684(.A(pi217), .B(pi131), .Y(new_n1061));
  nand_5 g00685(.A(pi249), .B(pi168), .Y(new_n1062));
  not_8  g00686(.A(pi236), .Y(new_n1063));
  not_8  g00687(.A(pi242), .Y(new_n1064));
  nor_5  g00688(.A(new_n1064), .B(new_n1063), .Y(new_n1065));
  not_8  g00689(.A(pi210), .Y(new_n1066));
  not_8  g00690(.A(pi213), .Y(new_n1067));
  nor_5  g00691(.A(new_n1067), .B(new_n1066), .Y(new_n1068));
  xnor_4 g00692(.A(new_n1068), .B(new_n1065), .Y(new_n1069));
  xnor_4 g00693(.A(new_n1069), .B(new_n1062), .Y(new_n1070));
  or_6   g00694(.A(new_n1070), .B(new_n1061), .Y(new_n1071));
  not_8  g00695(.A(new_n1071), .Y(new_n1072));
  nand_5 g00696(.A(pi131), .B(pi100), .Y(new_n1073));
  nand_5 g00697(.A(pi217), .B(pi052), .Y(new_n1074));
  xor_4  g00698(.A(new_n1074), .B(new_n1073), .Y(new_n1075));
  nor_5  g00699(.A(new_n1075), .B(new_n1072), .Y(new_n1076));
  nand_5 g00700(.A(new_n1068), .B(new_n1065), .Y(new_n1077));
  nand_5 g00701(.A(pi242), .B(pi241), .Y(new_n1078));
  nand_5 g00702(.A(pi236), .B(pi140), .Y(new_n1079));
  xor_4  g00703(.A(new_n1079), .B(new_n1078), .Y(new_n1080));
  nand_5 g00704(.A(pi212), .B(pi210), .Y(new_n1081));
  nand_5 g00705(.A(pi213), .B(pi111), .Y(new_n1082));
  xor_4  g00706(.A(new_n1082), .B(new_n1081), .Y(new_n1083));
  xor_4  g00707(.A(new_n1083), .B(new_n1080), .Y(new_n1084));
  xor_4  g00708(.A(new_n1084), .B(new_n1077), .Y(new_n1085));
  or_6   g00709(.A(new_n1069), .B(new_n1062), .Y(new_n1086));
  nand_5 g00710(.A(pi222), .B(pi208), .Y(new_n1087));
  or_6   g00711(.A(new_n1087), .B(new_n1062), .Y(new_n1088));
  nand_5 g00712(.A(pi249), .B(pi208), .Y(new_n1089));
  nand_5 g00713(.A(pi222), .B(pi168), .Y(new_n1090));
  nand_5 g00714(.A(new_n1090), .B(new_n1089), .Y(new_n1091));
  nand_5 g00715(.A(new_n1091), .B(new_n1088), .Y(new_n1092));
  xnor_4 g00716(.A(new_n1092), .B(new_n1086), .Y(new_n1093));
  xor_4  g00717(.A(new_n1093), .B(new_n1085), .Y(new_n1094));
  xor_4  g00718(.A(new_n1075), .B(new_n1071), .Y(new_n1095));
  nor_5  g00719(.A(new_n1095), .B(new_n1094), .Y(new_n1096));
  nor_5  g00720(.A(new_n1096), .B(new_n1076), .Y(new_n1097));
  not_8  g00721(.A(new_n1097), .Y(new_n1098));
  nand_5 g00722(.A(pi217), .B(pi077), .Y(new_n1099));
  nand_5 g00723(.A(pi227), .B(pi131), .Y(new_n1100));
  nor_5  g00724(.A(new_n1100), .B(new_n1099), .Y(new_n1101));
  nand_5 g00725(.A(new_n1100), .B(new_n1099), .Y(new_n1102));
  nand_5 g00726(.A(pi100), .B(pi052), .Y(new_n1103));
  not_8  g00727(.A(new_n1103), .Y(new_n1104));
  and_6  g00728(.A(new_n1104), .B(new_n1061), .Y(new_n1105));
  nor_5  g00729(.A(new_n1105), .B(new_n1102), .Y(new_n1106));
  nor_5  g00730(.A(new_n1106), .B(new_n1101), .Y(new_n1107));
  nand_5 g00731(.A(new_n1105), .B(new_n1102), .Y(new_n1108));
  nand_5 g00732(.A(new_n1108), .B(new_n1107), .Y(new_n1109));
  nand_5 g00733(.A(new_n1109), .B(new_n1098), .Y(new_n1110));
  xor_4  g00734(.A(new_n1109), .B(new_n1097), .Y(new_n1111));
  or_6   g00735(.A(new_n1083), .B(new_n1080), .Y(new_n1112));
  nand_5 g00736(.A(new_n1084), .B(new_n1077), .Y(new_n1113));
  nand_5 g00737(.A(new_n1113), .B(new_n1112), .Y(new_n1114));
  nand_5 g00738(.A(pi241), .B(pi140), .Y(new_n1115));
  nor_5  g00739(.A(new_n1115), .B(new_n1065), .Y(new_n1116));
  nand_5 g00740(.A(pi242), .B(pi161), .Y(new_n1117));
  nand_5 g00741(.A(pi252), .B(pi236), .Y(new_n1118));
  nand_5 g00742(.A(new_n1118), .B(new_n1117), .Y(new_n1119));
  nand_5 g00743(.A(new_n1119), .B(new_n1116), .Y(new_n1120));
  nor_5  g00744(.A(new_n1118), .B(new_n1117), .Y(new_n1121));
  nor_5  g00745(.A(new_n1119), .B(new_n1116), .Y(new_n1122));
  nor_5  g00746(.A(new_n1122), .B(new_n1121), .Y(new_n1123));
  nand_5 g00747(.A(new_n1123), .B(new_n1120), .Y(new_n1124));
  nand_5 g00748(.A(pi210), .B(pi104), .Y(new_n1125));
  nand_5 g00749(.A(pi213), .B(pi024), .Y(new_n1126));
  nand_5 g00750(.A(new_n1126), .B(new_n1125), .Y(new_n1127));
  nand_5 g00751(.A(pi212), .B(pi111), .Y(new_n1128));
  nor_5  g00752(.A(new_n1128), .B(new_n1068), .Y(new_n1129));
  nand_5 g00753(.A(new_n1129), .B(new_n1127), .Y(new_n1130));
  nor_5  g00754(.A(new_n1126), .B(new_n1125), .Y(new_n1131));
  nor_5  g00755(.A(new_n1129), .B(new_n1127), .Y(new_n1132));
  nor_5  g00756(.A(new_n1132), .B(new_n1131), .Y(new_n1133));
  nand_5 g00757(.A(new_n1133), .B(new_n1130), .Y(new_n1134));
  xor_4  g00758(.A(new_n1134), .B(new_n1124), .Y(new_n1135));
  xor_4  g00759(.A(new_n1135), .B(new_n1114), .Y(new_n1136));
  nand_5 g00760(.A(pi249), .B(pi139), .Y(new_n1137));
  nand_5 g00761(.A(pi168), .B(pi125), .Y(new_n1138));
  xor_4  g00762(.A(new_n1138), .B(new_n1087), .Y(new_n1139));
  xor_4  g00763(.A(new_n1139), .B(new_n1137), .Y(new_n1140));
  xnor_4 g00764(.A(new_n1140), .B(new_n1088), .Y(new_n1141));
  xnor_4 g00765(.A(new_n1141), .B(new_n1136), .Y(new_n1142));
  nor_5  g00766(.A(new_n1092), .B(new_n1086), .Y(new_n1143));
  nor_5  g00767(.A(new_n1093), .B(new_n1085), .Y(new_n1144));
  nor_5  g00768(.A(new_n1144), .B(new_n1143), .Y(new_n1145));
  xor_4  g00769(.A(new_n1145), .B(new_n1142), .Y(new_n1146));
  or_6   g00770(.A(new_n1146), .B(new_n1111), .Y(new_n1147));
  nand_5 g00771(.A(new_n1147), .B(new_n1110), .Y(new_n1148));
  nand_5 g00772(.A(pi100), .B(pi077), .Y(new_n1149));
  nand_5 g00773(.A(pi217), .B(pi133), .Y(new_n1150));
  nand_5 g00774(.A(pi227), .B(pi052), .Y(new_n1151));
  xor_4  g00775(.A(new_n1151), .B(new_n1150), .Y(new_n1152));
  xor_4  g00776(.A(new_n1152), .B(new_n1149), .Y(new_n1153));
  not_8  g00777(.A(new_n1102), .Y(new_n1154));
  nor_5  g00778(.A(new_n1104), .B(new_n1101), .Y(new_n1155));
  nor_5  g00779(.A(new_n1155), .B(new_n1154), .Y(new_n1156));
  not_8  g00780(.A(new_n1156), .Y(new_n1157));
  nand_5 g00781(.A(pi131), .B(pi081), .Y(new_n1158));
  xor_4  g00782(.A(new_n1158), .B(new_n1157), .Y(new_n1159));
  xor_4  g00783(.A(new_n1159), .B(new_n1153), .Y(new_n1160));
  nor_5  g00784(.A(new_n1107), .B(new_n1103), .Y(new_n1161));
  xor_4  g00785(.A(new_n1161), .B(new_n1160), .Y(new_n1162));
  xnor_4 g00786(.A(new_n1162), .B(new_n1148), .Y(new_n1163));
  nor_5  g00787(.A(new_n1141), .B(new_n1136), .Y(new_n1164));
  nor_5  g00788(.A(new_n1145), .B(new_n1142), .Y(new_n1165));
  nor_5  g00789(.A(new_n1165), .B(new_n1164), .Y(new_n1166));
  nor_5  g00790(.A(new_n1140), .B(new_n1088), .Y(new_n1167));
  not_8  g00791(.A(new_n1167), .Y(new_n1168));
  nand_5 g00792(.A(pi208), .B(pi125), .Y(new_n1169));
  nand_5 g00793(.A(pi249), .B(pi035), .Y(new_n1170));
  nand_5 g00794(.A(pi222), .B(pi139), .Y(new_n1171));
  xor_4  g00795(.A(new_n1171), .B(new_n1170), .Y(new_n1172));
  xor_4  g00796(.A(new_n1172), .B(new_n1169), .Y(new_n1173));
  nand_5 g00797(.A(pi176), .B(pi168), .Y(new_n1174));
  nand_5 g00798(.A(new_n1138), .B(new_n1087), .Y(new_n1175));
  nand_5 g00799(.A(new_n1139), .B(new_n1137), .Y(new_n1176));
  nand_5 g00800(.A(new_n1176), .B(new_n1175), .Y(new_n1177));
  xor_4  g00801(.A(new_n1177), .B(new_n1174), .Y(new_n1178));
  xor_4  g00802(.A(new_n1178), .B(new_n1173), .Y(new_n1179));
  xor_4  g00803(.A(new_n1179), .B(new_n1168), .Y(new_n1180));
  nand_5 g00804(.A(new_n1134), .B(new_n1124), .Y(new_n1181));
  nand_5 g00805(.A(new_n1135), .B(new_n1114), .Y(new_n1182));
  nand_5 g00806(.A(new_n1182), .B(new_n1181), .Y(new_n1183));
  nor_5  g00807(.A(new_n1133), .B(new_n1128), .Y(new_n1184));
  nand_5 g00808(.A(pi111), .B(pi104), .Y(new_n1185));
  nand_5 g00809(.A(pi210), .B(pi013), .Y(new_n1186));
  nand_5 g00810(.A(pi212), .B(pi024), .Y(new_n1187));
  xor_4  g00811(.A(new_n1187), .B(new_n1186), .Y(new_n1188));
  xor_4  g00812(.A(new_n1188), .B(new_n1185), .Y(new_n1189));
  not_8  g00813(.A(new_n1128), .Y(new_n1190));
  or_6   g00814(.A(new_n1131), .B(new_n1190), .Y(new_n1191));
  nand_5 g00815(.A(new_n1191), .B(new_n1127), .Y(new_n1192));
  nand_5 g00816(.A(pi224), .B(pi213), .Y(new_n1193));
  xor_4  g00817(.A(new_n1193), .B(new_n1192), .Y(new_n1194));
  xnor_4 g00818(.A(new_n1194), .B(new_n1189), .Y(new_n1195));
  xor_4  g00819(.A(new_n1195), .B(new_n1184), .Y(new_n1196));
  nor_5  g00820(.A(new_n1123), .B(new_n1115), .Y(new_n1197));
  nand_5 g00821(.A(pi161), .B(pi140), .Y(new_n1198));
  nand_5 g00822(.A(pi242), .B(pi141), .Y(new_n1199));
  nand_5 g00823(.A(pi252), .B(pi241), .Y(new_n1200));
  xnor_4 g00824(.A(new_n1200), .B(new_n1199), .Y(new_n1201));
  xor_4  g00825(.A(new_n1201), .B(new_n1198), .Y(new_n1202));
  not_8  g00826(.A(new_n1115), .Y(new_n1203));
  or_6   g00827(.A(new_n1121), .B(new_n1203), .Y(new_n1204));
  nand_5 g00828(.A(new_n1204), .B(new_n1119), .Y(new_n1205));
  nand_5 g00829(.A(pi236), .B(pi121), .Y(new_n1206));
  xor_4  g00830(.A(new_n1206), .B(new_n1205), .Y(new_n1207));
  xor_4  g00831(.A(new_n1207), .B(new_n1202), .Y(new_n1208));
  xor_4  g00832(.A(new_n1208), .B(new_n1197), .Y(new_n1209));
  nand_5 g00833(.A(new_n1209), .B(new_n1196), .Y(new_n1210));
  or_6   g00834(.A(new_n1209), .B(new_n1196), .Y(new_n1211));
  nand_5 g00835(.A(new_n1211), .B(new_n1210), .Y(new_n1212));
  xnor_4 g00836(.A(new_n1212), .B(new_n1183), .Y(new_n1213));
  xor_4  g00837(.A(new_n1213), .B(new_n1180), .Y(new_n1214));
  xor_4  g00838(.A(new_n1214), .B(new_n1166), .Y(new_n1215));
  xnor_4 g00839(.A(new_n1215), .B(new_n1163), .Y(po004));
  nand_5 g00840(.A(pi093), .B(pi041), .Y(new_n1217));
  nand_5 g00841(.A(pi045), .B(pi020), .Y(new_n1218));
  nand_5 g00842(.A(pi119), .B(pi060), .Y(new_n1219));
  nand_5 g00843(.A(pi250), .B(pi160), .Y(new_n1220));
  nand_5 g00844(.A(new_n1220), .B(new_n1219), .Y(new_n1221));
  not_8  g00845(.A(new_n1218), .Y(new_n1222));
  and_6  g00846(.A(new_n1222), .B(new_n1054), .Y(new_n1223));
  nor_5  g00847(.A(new_n1223), .B(new_n1221), .Y(new_n1224));
  nor_5  g00848(.A(new_n1220), .B(new_n1219), .Y(new_n1225));
  nor_5  g00849(.A(new_n1225), .B(new_n1224), .Y(new_n1226));
  nor_5  g00850(.A(new_n1226), .B(new_n1218), .Y(new_n1227));
  or_6   g00851(.A(new_n1225), .B(new_n1222), .Y(new_n1228));
  nand_5 g00852(.A(new_n1228), .B(new_n1221), .Y(new_n1229));
  nand_5 g00853(.A(pi160), .B(pi044), .Y(new_n1230));
  xor_4  g00854(.A(new_n1230), .B(new_n1229), .Y(new_n1231));
  nand_5 g00855(.A(pi250), .B(pi020), .Y(new_n1232));
  nand_5 g00856(.A(pi060), .B(pi045), .Y(new_n1233));
  nand_5 g00857(.A(pi223), .B(pi119), .Y(new_n1234));
  xor_4  g00858(.A(new_n1234), .B(new_n1233), .Y(new_n1235));
  xor_4  g00859(.A(new_n1235), .B(new_n1232), .Y(new_n1236));
  xor_4  g00860(.A(new_n1236), .B(new_n1231), .Y(new_n1237));
  not_8  g00861(.A(new_n1237), .Y(new_n1238));
  xor_4  g00862(.A(new_n1238), .B(new_n1227), .Y(new_n1239));
  nor_5  g00863(.A(new_n1059), .B(new_n1054), .Y(new_n1240));
  nand_5 g00864(.A(pi160), .B(pi045), .Y(new_n1241));
  nand_5 g00865(.A(pi119), .B(pi020), .Y(new_n1242));
  xor_4  g00866(.A(new_n1242), .B(new_n1241), .Y(new_n1243));
  nor_5  g00867(.A(new_n1243), .B(new_n1240), .Y(new_n1244));
  not_8  g00868(.A(new_n1055), .Y(new_n1245));
  nand_5 g00869(.A(new_n1058), .B(new_n1245), .Y(new_n1246));
  nand_5 g00870(.A(pi151), .B(pi138), .Y(new_n1247));
  nand_5 g00871(.A(pi182), .B(pi147), .Y(new_n1248));
  and_6  g00872(.A(new_n1248), .B(new_n1247), .Y(new_n1249));
  nand_5 g00873(.A(pi182), .B(pi151), .Y(new_n1250));
  nor_5  g00874(.A(new_n1250), .B(new_n1055), .Y(new_n1251));
  or_6   g00875(.A(new_n1251), .B(new_n1249), .Y(new_n1252));
  xnor_4 g00876(.A(new_n1252), .B(new_n1246), .Y(new_n1253));
  nor_5  g00877(.A(new_n1057), .B(new_n1056), .Y(new_n1254));
  nand_5 g00878(.A(pi087), .B(pi026), .Y(new_n1255));
  nand_5 g00879(.A(pi219), .B(pi027), .Y(new_n1256));
  and_6  g00880(.A(new_n1256), .B(new_n1255), .Y(new_n1257));
  nand_5 g00881(.A(pi219), .B(pi026), .Y(new_n1258));
  nor_5  g00882(.A(new_n1258), .B(new_n1056), .Y(new_n1259));
  or_6   g00883(.A(new_n1259), .B(new_n1257), .Y(new_n1260));
  nand_5 g00884(.A(pi164), .B(pi071), .Y(new_n1261));
  nand_5 g00885(.A(pi206), .B(pi142), .Y(new_n1262));
  xnor_4 g00886(.A(new_n1262), .B(new_n1261), .Y(new_n1263));
  xnor_4 g00887(.A(new_n1263), .B(new_n1260), .Y(new_n1264));
  xor_4  g00888(.A(new_n1264), .B(new_n1254), .Y(new_n1265));
  xor_4  g00889(.A(new_n1265), .B(new_n1253), .Y(new_n1266));
  xnor_4 g00890(.A(new_n1243), .B(new_n1240), .Y(new_n1267));
  nor_5  g00891(.A(new_n1267), .B(new_n1266), .Y(new_n1268));
  or_6   g00892(.A(new_n1268), .B(new_n1244), .Y(new_n1269));
  nand_5 g00893(.A(pi102), .B(pi027), .Y(new_n1270));
  nand_5 g00894(.A(pi087), .B(pi008), .Y(new_n1271));
  xor_4  g00895(.A(new_n1271), .B(new_n1258), .Y(new_n1272));
  xor_4  g00896(.A(new_n1272), .B(new_n1270), .Y(new_n1273));
  xor_4  g00897(.A(new_n1273), .B(new_n1259), .Y(new_n1274));
  nand_5 g00898(.A(pi169), .B(pi164), .Y(new_n1275));
  nand_5 g00899(.A(pi142), .B(pi032), .Y(new_n1276));
  nand_5 g00900(.A(new_n1276), .B(new_n1275), .Y(new_n1277));
  not_8  g00901(.A(new_n1057), .Y(new_n1278));
  nand_5 g00902(.A(pi206), .B(pi071), .Y(new_n1279));
  nor_5  g00903(.A(new_n1279), .B(new_n1278), .Y(new_n1280));
  nand_5 g00904(.A(new_n1280), .B(new_n1277), .Y(new_n1281));
  or_6   g00905(.A(new_n1276), .B(new_n1275), .Y(new_n1282));
  and_6  g00906(.A(new_n1282), .B(new_n1277), .Y(new_n1283));
  or_6   g00907(.A(new_n1283), .B(new_n1280), .Y(new_n1284));
  nand_5 g00908(.A(new_n1284), .B(new_n1281), .Y(new_n1285));
  nand_5 g00909(.A(new_n1263), .B(new_n1260), .Y(new_n1286));
  or_6   g00910(.A(new_n1264), .B(new_n1254), .Y(new_n1287));
  nand_5 g00911(.A(new_n1287), .B(new_n1286), .Y(new_n1288));
  xor_4  g00912(.A(new_n1288), .B(new_n1285), .Y(new_n1289));
  xor_4  g00913(.A(new_n1289), .B(new_n1274), .Y(new_n1290));
  nand_5 g00914(.A(pi147), .B(pi041), .Y(new_n1291));
  nand_5 g00915(.A(pi138), .B(pi019), .Y(new_n1292));
  xor_4  g00916(.A(new_n1292), .B(new_n1250), .Y(new_n1293));
  xnor_4 g00917(.A(new_n1293), .B(new_n1291), .Y(new_n1294));
  xor_4  g00918(.A(new_n1294), .B(new_n1251), .Y(new_n1295));
  nor_5  g00919(.A(new_n1252), .B(new_n1246), .Y(new_n1296));
  nor_5  g00920(.A(new_n1265), .B(new_n1253), .Y(new_n1297));
  nor_5  g00921(.A(new_n1297), .B(new_n1296), .Y(new_n1298));
  xor_4  g00922(.A(new_n1298), .B(new_n1295), .Y(new_n1299));
  xnor_4 g00923(.A(new_n1299), .B(new_n1290), .Y(new_n1300));
  nor_5  g00924(.A(new_n1300), .B(new_n1269), .Y(new_n1301));
  xnor_4 g00925(.A(new_n1300), .B(new_n1269), .Y(new_n1302));
  nand_5 g00926(.A(new_n1223), .B(new_n1221), .Y(new_n1303));
  nand_5 g00927(.A(new_n1303), .B(new_n1226), .Y(new_n1304));
  nor_5  g00928(.A(new_n1304), .B(new_n1302), .Y(new_n1305));
  or_6   g00929(.A(new_n1305), .B(new_n1301), .Y(new_n1306));
  nor_5  g00930(.A(new_n1306), .B(new_n1239), .Y(new_n1307));
  not_8  g00931(.A(new_n1295), .Y(new_n1308));
  nor_5  g00932(.A(new_n1298), .B(new_n1308), .Y(new_n1309));
  nor_5  g00933(.A(new_n1299), .B(new_n1290), .Y(new_n1310));
  nor_5  g00934(.A(new_n1310), .B(new_n1309), .Y(new_n1311));
  nand_5 g00935(.A(new_n1294), .B(new_n1251), .Y(new_n1312));
  nand_5 g00936(.A(pi182), .B(pi019), .Y(new_n1313));
  nand_5 g00937(.A(pi216), .B(pi147), .Y(new_n1314));
  nand_5 g00938(.A(pi151), .B(pi041), .Y(new_n1315));
  xor_4  g00939(.A(new_n1315), .B(new_n1314), .Y(new_n1316));
  xor_4  g00940(.A(new_n1316), .B(new_n1313), .Y(new_n1317));
  not_8  g00941(.A(new_n1317), .Y(new_n1318));
  nand_5 g00942(.A(pi138), .B(pi097), .Y(new_n1319));
  nand_5 g00943(.A(new_n1292), .B(new_n1250), .Y(new_n1320));
  nand_5 g00944(.A(new_n1293), .B(new_n1291), .Y(new_n1321));
  nand_5 g00945(.A(new_n1321), .B(new_n1320), .Y(new_n1322));
  xor_4  g00946(.A(new_n1322), .B(new_n1319), .Y(new_n1323));
  xor_4  g00947(.A(new_n1323), .B(new_n1318), .Y(new_n1324));
  xor_4  g00948(.A(new_n1324), .B(new_n1312), .Y(new_n1325));
  xor_4  g00949(.A(new_n1325), .B(new_n1311), .Y(new_n1326));
  nand_5 g00950(.A(pi071), .B(pi032), .Y(new_n1327));
  nand_5 g00951(.A(pi164), .B(pi123), .Y(new_n1328));
  nand_5 g00952(.A(pi206), .B(pi169), .Y(new_n1329));
  xor_4  g00953(.A(new_n1329), .B(new_n1328), .Y(new_n1330));
  xor_4  g00954(.A(new_n1330), .B(new_n1327), .Y(new_n1331));
  nand_5 g00955(.A(new_n1282), .B(new_n1279), .Y(new_n1332));
  nand_5 g00956(.A(new_n1332), .B(new_n1277), .Y(new_n1333));
  nand_5 g00957(.A(pi145), .B(pi142), .Y(new_n1334));
  xor_4  g00958(.A(new_n1334), .B(new_n1333), .Y(new_n1335));
  xnor_4 g00959(.A(new_n1335), .B(new_n1331), .Y(new_n1336));
  nor_5  g00960(.A(new_n1284), .B(new_n1279), .Y(new_n1337));
  xor_4  g00961(.A(new_n1337), .B(new_n1336), .Y(new_n1338));
  not_8  g00962(.A(new_n1259), .Y(new_n1339));
  nor_5  g00963(.A(new_n1273), .B(new_n1339), .Y(new_n1340));
  nand_5 g00964(.A(pi219), .B(pi008), .Y(new_n1341));
  nand_5 g00965(.A(pi027), .B(pi001), .Y(new_n1342));
  nand_5 g00966(.A(pi102), .B(pi026), .Y(new_n1343));
  xor_4  g00967(.A(new_n1343), .B(new_n1342), .Y(new_n1344));
  xor_4  g00968(.A(new_n1344), .B(new_n1341), .Y(new_n1345));
  nand_5 g00969(.A(pi087), .B(pi056), .Y(new_n1346));
  nand_5 g00970(.A(new_n1271), .B(new_n1258), .Y(new_n1347));
  nand_5 g00971(.A(new_n1272), .B(new_n1270), .Y(new_n1348));
  nand_5 g00972(.A(new_n1348), .B(new_n1347), .Y(new_n1349));
  xor_4  g00973(.A(new_n1349), .B(new_n1346), .Y(new_n1350));
  xor_4  g00974(.A(new_n1350), .B(new_n1345), .Y(new_n1351));
  xor_4  g00975(.A(new_n1351), .B(new_n1340), .Y(new_n1352));
  nand_5 g00976(.A(new_n1288), .B(new_n1285), .Y(new_n1353));
  nand_5 g00977(.A(new_n1289), .B(new_n1274), .Y(new_n1354));
  nand_5 g00978(.A(new_n1354), .B(new_n1353), .Y(new_n1355));
  xnor_4 g00979(.A(new_n1355), .B(new_n1352), .Y(new_n1356));
  xnor_4 g00980(.A(new_n1356), .B(new_n1338), .Y(new_n1357));
  xor_4  g00981(.A(new_n1357), .B(new_n1326), .Y(new_n1358));
  xnor_4 g00982(.A(new_n1306), .B(new_n1239), .Y(new_n1359));
  nor_5  g00983(.A(new_n1359), .B(new_n1358), .Y(new_n1360));
  nor_5  g00984(.A(new_n1360), .B(new_n1307), .Y(new_n1361));
  nand_5 g00985(.A(new_n1238), .B(new_n1227), .Y(new_n1362));
  nand_5 g00986(.A(pi250), .B(pi060), .Y(new_n1363));
  nand_5 g00987(.A(pi119), .B(pi101), .Y(new_n1364));
  xor_4  g00988(.A(new_n1364), .B(new_n1363), .Y(new_n1365));
  nand_5 g00989(.A(pi223), .B(pi045), .Y(new_n1366));
  xor_4  g00990(.A(new_n1366), .B(new_n1365), .Y(new_n1367));
  nand_5 g00991(.A(pi044), .B(pi020), .Y(new_n1368));
  nand_5 g00992(.A(new_n1234), .B(new_n1233), .Y(new_n1369));
  nand_5 g00993(.A(new_n1235), .B(new_n1232), .Y(new_n1370));
  nand_5 g00994(.A(new_n1370), .B(new_n1369), .Y(new_n1371));
  xor_4  g00995(.A(new_n1371), .B(new_n1368), .Y(new_n1372));
  xor_4  g00996(.A(new_n1372), .B(new_n1367), .Y(new_n1373));
  nand_5 g00997(.A(pi160), .B(pi054), .Y(new_n1374));
  xor_4  g00998(.A(new_n1374), .B(new_n1373), .Y(new_n1375));
  nor_5  g00999(.A(new_n1230), .B(new_n1229), .Y(new_n1376));
  not_8  g01000(.A(new_n1236), .Y(new_n1377));
  nand_5 g01001(.A(new_n1377), .B(new_n1231), .Y(new_n1378));
  not_8  g01002(.A(new_n1378), .Y(new_n1379));
  nor_5  g01003(.A(new_n1379), .B(new_n1376), .Y(new_n1380));
  xor_4  g01004(.A(new_n1380), .B(new_n1375), .Y(new_n1381));
  xor_4  g01005(.A(new_n1381), .B(new_n1362), .Y(new_n1382));
  nand_5 g01006(.A(new_n1382), .B(new_n1361), .Y(new_n1383));
  or_6   g01007(.A(new_n1325), .B(new_n1311), .Y(new_n1384));
  nand_5 g01008(.A(new_n1357), .B(new_n1326), .Y(new_n1385));
  nand_5 g01009(.A(new_n1385), .B(new_n1384), .Y(new_n1386));
  not_8  g01010(.A(new_n1324), .Y(new_n1387));
  nor_5  g01011(.A(new_n1387), .B(new_n1312), .Y(new_n1388));
  not_8  g01012(.A(new_n1388), .Y(new_n1389));
  nand_5 g01013(.A(pi216), .B(pi151), .Y(new_n1390));
  nand_5 g01014(.A(pi041), .B(pi019), .Y(new_n1391));
  nand_5 g01015(.A(pi147), .B(pi076), .Y(new_n1392));
  xor_4  g01016(.A(new_n1392), .B(new_n1391), .Y(new_n1393));
  xor_4  g01017(.A(new_n1393), .B(new_n1390), .Y(new_n1394));
  nand_5 g01018(.A(new_n1315), .B(new_n1314), .Y(new_n1395));
  nand_5 g01019(.A(new_n1316), .B(new_n1313), .Y(new_n1396));
  nand_5 g01020(.A(new_n1396), .B(new_n1395), .Y(new_n1397));
  nand_5 g01021(.A(pi182), .B(pi097), .Y(new_n1398));
  xor_4  g01022(.A(new_n1398), .B(new_n1397), .Y(new_n1399));
  xor_4  g01023(.A(new_n1399), .B(new_n1394), .Y(new_n1400));
  nand_5 g01024(.A(pi138), .B(pi075), .Y(new_n1401));
  nor_5  g01025(.A(new_n1322), .B(new_n1319), .Y(new_n1402));
  nand_5 g01026(.A(new_n1323), .B(new_n1318), .Y(new_n1403));
  not_8  g01027(.A(new_n1403), .Y(new_n1404));
  or_6   g01028(.A(new_n1404), .B(new_n1402), .Y(new_n1405));
  xor_4  g01029(.A(new_n1405), .B(new_n1401), .Y(new_n1406));
  xnor_4 g01030(.A(new_n1406), .B(new_n1400), .Y(new_n1407));
  xor_4  g01031(.A(new_n1407), .B(new_n1389), .Y(new_n1408));
  not_8  g01032(.A(new_n1340), .Y(new_n1409));
  nor_5  g01033(.A(new_n1351), .B(new_n1409), .Y(new_n1410));
  nor_5  g01034(.A(new_n1349), .B(new_n1346), .Y(new_n1411));
  not_8  g01035(.A(new_n1350), .Y(new_n1412));
  nor_5  g01036(.A(new_n1412), .B(new_n1345), .Y(new_n1413));
  nor_5  g01037(.A(new_n1413), .B(new_n1411), .Y(new_n1414));
  nand_5 g01038(.A(pi136), .B(pi087), .Y(new_n1415));
  nand_5 g01039(.A(pi102), .B(pi008), .Y(new_n1416));
  nand_5 g01040(.A(pi122), .B(pi027), .Y(new_n1417));
  nand_5 g01041(.A(pi026), .B(pi001), .Y(new_n1418));
  xor_4  g01042(.A(new_n1418), .B(new_n1417), .Y(new_n1419));
  xor_4  g01043(.A(new_n1419), .B(new_n1416), .Y(new_n1420));
  nand_5 g01044(.A(pi219), .B(pi056), .Y(new_n1421));
  nand_5 g01045(.A(new_n1343), .B(new_n1342), .Y(new_n1422));
  nand_5 g01046(.A(new_n1344), .B(new_n1341), .Y(new_n1423));
  nand_5 g01047(.A(new_n1423), .B(new_n1422), .Y(new_n1424));
  xor_4  g01048(.A(new_n1424), .B(new_n1421), .Y(new_n1425));
  xor_4  g01049(.A(new_n1425), .B(new_n1420), .Y(new_n1426));
  xnor_4 g01050(.A(new_n1426), .B(new_n1415), .Y(new_n1427));
  xor_4  g01051(.A(new_n1427), .B(new_n1414), .Y(new_n1428));
  xnor_4 g01052(.A(new_n1428), .B(new_n1410), .Y(new_n1429));
  nand_5 g01053(.A(new_n1337), .B(new_n1336), .Y(new_n1430));
  not_8  g01054(.A(new_n1430), .Y(new_n1431));
  nand_5 g01055(.A(pi246), .B(pi142), .Y(new_n1432));
  nand_5 g01056(.A(new_n1334), .B(new_n1333), .Y(new_n1433));
  nand_5 g01057(.A(new_n1335), .B(new_n1331), .Y(new_n1434));
  nand_5 g01058(.A(new_n1434), .B(new_n1433), .Y(new_n1435));
  xor_4  g01059(.A(new_n1435), .B(new_n1432), .Y(new_n1436));
  nand_5 g01060(.A(pi169), .B(pi032), .Y(new_n1437));
  nand_5 g01061(.A(pi206), .B(pi123), .Y(new_n1438));
  nand_5 g01062(.A(pi164), .B(pi099), .Y(new_n1439));
  xor_4  g01063(.A(new_n1439), .B(new_n1438), .Y(new_n1440));
  xor_4  g01064(.A(new_n1440), .B(new_n1437), .Y(new_n1441));
  nand_5 g01065(.A(pi145), .B(pi071), .Y(new_n1442));
  nand_5 g01066(.A(new_n1329), .B(new_n1328), .Y(new_n1443));
  nand_5 g01067(.A(new_n1330), .B(new_n1327), .Y(new_n1444));
  nand_5 g01068(.A(new_n1444), .B(new_n1443), .Y(new_n1445));
  xor_4  g01069(.A(new_n1445), .B(new_n1442), .Y(new_n1446));
  xnor_4 g01070(.A(new_n1446), .B(new_n1441), .Y(new_n1447));
  xor_4  g01071(.A(new_n1447), .B(new_n1436), .Y(new_n1448));
  xor_4  g01072(.A(new_n1448), .B(new_n1431), .Y(new_n1449));
  and_6  g01073(.A(new_n1355), .B(new_n1352), .Y(new_n1450));
  nor_5  g01074(.A(new_n1356), .B(new_n1338), .Y(new_n1451));
  nor_5  g01075(.A(new_n1451), .B(new_n1450), .Y(new_n1452));
  xnor_4 g01076(.A(new_n1452), .B(new_n1449), .Y(new_n1453));
  xor_4  g01077(.A(new_n1453), .B(new_n1429), .Y(new_n1454));
  xnor_4 g01078(.A(new_n1454), .B(new_n1408), .Y(new_n1455));
  xnor_4 g01079(.A(new_n1455), .B(new_n1386), .Y(new_n1456));
  xor_4  g01080(.A(new_n1382), .B(new_n1361), .Y(new_n1457));
  nand_5 g01081(.A(new_n1457), .B(new_n1456), .Y(new_n1458));
  nand_5 g01082(.A(new_n1458), .B(new_n1383), .Y(new_n1459));
  nor_5  g01083(.A(new_n1374), .B(new_n1373), .Y(new_n1460));
  not_8  g01084(.A(new_n1375), .Y(new_n1461));
  nor_5  g01085(.A(new_n1380), .B(new_n1461), .Y(new_n1462));
  nor_5  g01086(.A(new_n1462), .B(new_n1460), .Y(new_n1463));
  nand_5 g01087(.A(pi250), .B(pi223), .Y(new_n1464));
  nand_5 g01088(.A(new_n1364), .B(new_n1363), .Y(new_n1465));
  nand_5 g01089(.A(new_n1366), .B(new_n1365), .Y(new_n1466));
  nand_5 g01090(.A(new_n1466), .B(new_n1465), .Y(new_n1467));
  nand_5 g01091(.A(pi225), .B(pi119), .Y(new_n1468));
  nand_5 g01092(.A(pi101), .B(pi045), .Y(new_n1469));
  nand_5 g01093(.A(new_n1469), .B(new_n1468), .Y(new_n1470));
  nand_5 g01094(.A(pi225), .B(pi045), .Y(new_n1471));
  nor_5  g01095(.A(new_n1471), .B(new_n1364), .Y(new_n1472));
  not_8  g01096(.A(new_n1472), .Y(new_n1473));
  nand_5 g01097(.A(new_n1473), .B(new_n1470), .Y(new_n1474));
  xor_4  g01098(.A(new_n1474), .B(new_n1467), .Y(new_n1475));
  xor_4  g01099(.A(new_n1475), .B(new_n1464), .Y(new_n1476));
  nand_5 g01100(.A(new_n1371), .B(new_n1368), .Y(new_n1477));
  nand_5 g01101(.A(new_n1372), .B(new_n1367), .Y(new_n1478));
  nand_5 g01102(.A(new_n1478), .B(new_n1477), .Y(new_n1479));
  nand_5 g01103(.A(pi060), .B(pi044), .Y(new_n1480));
  nand_5 g01104(.A(pi054), .B(pi020), .Y(new_n1481));
  nand_5 g01105(.A(new_n1481), .B(new_n1480), .Y(new_n1482));
  nand_5 g01106(.A(pi060), .B(pi054), .Y(new_n1483));
  nor_5  g01107(.A(new_n1483), .B(new_n1368), .Y(new_n1484));
  not_8  g01108(.A(new_n1484), .Y(new_n1485));
  nand_5 g01109(.A(new_n1485), .B(new_n1482), .Y(new_n1486));
  xor_4  g01110(.A(new_n1486), .B(new_n1479), .Y(new_n1487));
  xor_4  g01111(.A(new_n1487), .B(new_n1476), .Y(new_n1488));
  xor_4  g01112(.A(new_n1488), .B(new_n1463), .Y(new_n1489));
  nor_5  g01113(.A(new_n1381), .B(new_n1362), .Y(new_n1490));
  nand_5 g01114(.A(pi160), .B(pi072), .Y(new_n1491));
  xor_4  g01115(.A(new_n1491), .B(new_n1490), .Y(new_n1492));
  xor_4  g01116(.A(new_n1492), .B(new_n1489), .Y(new_n1493));
  not_8  g01117(.A(new_n1493), .Y(new_n1494));
  nor_5  g01118(.A(new_n1494), .B(new_n1459), .Y(new_n1495));
  xor_4  g01119(.A(new_n1493), .B(new_n1459), .Y(new_n1496));
  nor_5  g01120(.A(new_n1454), .B(new_n1408), .Y(new_n1497));
  nor_5  g01121(.A(new_n1455), .B(new_n1386), .Y(new_n1498));
  or_6   g01122(.A(new_n1498), .B(new_n1497), .Y(new_n1499));
  nor_5  g01123(.A(new_n1435), .B(new_n1432), .Y(new_n1500));
  nand_5 g01124(.A(new_n1447), .B(new_n1436), .Y(new_n1501));
  not_8  g01125(.A(new_n1501), .Y(new_n1502));
  or_6   g01126(.A(new_n1502), .B(new_n1500), .Y(new_n1503));
  nand_5 g01127(.A(new_n1445), .B(new_n1442), .Y(new_n1504));
  nand_5 g01128(.A(new_n1446), .B(new_n1441), .Y(new_n1505));
  nand_5 g01129(.A(new_n1505), .B(new_n1504), .Y(new_n1506));
  nand_5 g01130(.A(pi246), .B(pi071), .Y(new_n1507));
  nand_5 g01131(.A(pi169), .B(pi145), .Y(new_n1508));
  nand_5 g01132(.A(new_n1508), .B(new_n1507), .Y(new_n1509));
  nand_5 g01133(.A(pi246), .B(pi169), .Y(new_n1510));
  nor_5  g01134(.A(new_n1510), .B(new_n1442), .Y(new_n1511));
  not_8  g01135(.A(new_n1511), .Y(new_n1512));
  nand_5 g01136(.A(new_n1512), .B(new_n1509), .Y(new_n1513));
  nand_5 g01137(.A(pi164), .B(pi023), .Y(new_n1514));
  nand_5 g01138(.A(pi206), .B(pi099), .Y(new_n1515));
  nand_5 g01139(.A(new_n1515), .B(new_n1514), .Y(new_n1516));
  nand_5 g01140(.A(pi206), .B(pi023), .Y(new_n1517));
  nor_5  g01141(.A(new_n1517), .B(new_n1439), .Y(new_n1518));
  not_8  g01142(.A(new_n1518), .Y(new_n1519));
  nand_5 g01143(.A(new_n1519), .B(new_n1516), .Y(new_n1520));
  nand_5 g01144(.A(pi123), .B(pi032), .Y(new_n1521));
  nand_5 g01145(.A(new_n1439), .B(new_n1438), .Y(new_n1522));
  nand_5 g01146(.A(new_n1440), .B(new_n1437), .Y(new_n1523));
  nand_5 g01147(.A(new_n1523), .B(new_n1522), .Y(new_n1524));
  xor_4  g01148(.A(new_n1524), .B(new_n1521), .Y(new_n1525));
  xor_4  g01149(.A(new_n1525), .B(new_n1520), .Y(new_n1526));
  xor_4  g01150(.A(new_n1526), .B(new_n1513), .Y(new_n1527));
  xor_4  g01151(.A(new_n1527), .B(new_n1506), .Y(new_n1528));
  xor_4  g01152(.A(new_n1528), .B(new_n1503), .Y(new_n1529));
  nand_5 g01153(.A(new_n1448), .B(new_n1431), .Y(new_n1530));
  nand_5 g01154(.A(pi142), .B(pi114), .Y(new_n1531));
  xor_4  g01155(.A(new_n1531), .B(new_n1530), .Y(new_n1532));
  xor_4  g01156(.A(new_n1532), .B(new_n1529), .Y(new_n1533));
  nor_5  g01157(.A(new_n1452), .B(new_n1449), .Y(new_n1534));
  not_8  g01158(.A(new_n1429), .Y(new_n1535));
  nor_5  g01159(.A(new_n1453), .B(new_n1535), .Y(new_n1536));
  nor_5  g01160(.A(new_n1536), .B(new_n1534), .Y(new_n1537));
  and_6  g01161(.A(new_n1428), .B(new_n1410), .Y(new_n1538));
  nand_5 g01162(.A(pi096), .B(pi087), .Y(new_n1539));
  xor_4  g01163(.A(new_n1539), .B(new_n1538), .Y(new_n1540));
  nor_5  g01164(.A(new_n1426), .B(new_n1415), .Y(new_n1541));
  or_6   g01165(.A(new_n1427), .B(new_n1414), .Y(new_n1542));
  not_8  g01166(.A(new_n1542), .Y(new_n1543));
  or_6   g01167(.A(new_n1543), .B(new_n1541), .Y(new_n1544));
  nand_5 g01168(.A(pi219), .B(pi136), .Y(new_n1545));
  nand_5 g01169(.A(pi102), .B(pi056), .Y(new_n1546));
  and_6  g01170(.A(new_n1546), .B(new_n1545), .Y(new_n1547));
  nand_5 g01171(.A(pi136), .B(pi102), .Y(new_n1548));
  nor_5  g01172(.A(new_n1548), .B(new_n1421), .Y(new_n1549));
  or_6   g01173(.A(new_n1549), .B(new_n1547), .Y(new_n1550));
  nand_5 g01174(.A(new_n1418), .B(new_n1417), .Y(new_n1551));
  nand_5 g01175(.A(new_n1419), .B(new_n1416), .Y(new_n1552));
  nand_5 g01176(.A(new_n1552), .B(new_n1551), .Y(new_n1553));
  nand_5 g01177(.A(pi008), .B(pi001), .Y(new_n1554));
  nand_5 g01178(.A(pi122), .B(pi026), .Y(new_n1555));
  nand_5 g01179(.A(pi135), .B(pi027), .Y(new_n1556));
  nand_5 g01180(.A(new_n1556), .B(new_n1555), .Y(new_n1557));
  nand_5 g01181(.A(pi135), .B(pi026), .Y(new_n1558));
  nor_5  g01182(.A(new_n1558), .B(new_n1417), .Y(new_n1559));
  not_8  g01183(.A(new_n1559), .Y(new_n1560));
  nand_5 g01184(.A(new_n1560), .B(new_n1557), .Y(new_n1561));
  xor_4  g01185(.A(new_n1561), .B(new_n1554), .Y(new_n1562));
  xor_4  g01186(.A(new_n1562), .B(new_n1553), .Y(new_n1563));
  xor_4  g01187(.A(new_n1563), .B(new_n1550), .Y(new_n1564));
  nand_5 g01188(.A(new_n1424), .B(new_n1421), .Y(new_n1565));
  nand_5 g01189(.A(new_n1425), .B(new_n1420), .Y(new_n1566));
  nand_5 g01190(.A(new_n1566), .B(new_n1565), .Y(new_n1567));
  xor_4  g01191(.A(new_n1567), .B(new_n1564), .Y(new_n1568));
  xor_4  g01192(.A(new_n1568), .B(new_n1544), .Y(new_n1569));
  xor_4  g01193(.A(new_n1569), .B(new_n1540), .Y(new_n1570));
  xor_4  g01194(.A(new_n1570), .B(new_n1537), .Y(new_n1571));
  xor_4  g01195(.A(new_n1571), .B(new_n1533), .Y(new_n1572));
  or_6   g01196(.A(new_n1407), .B(new_n1389), .Y(new_n1573));
  nand_5 g01197(.A(pi138), .B(pi093), .Y(new_n1574));
  xor_4  g01198(.A(new_n1574), .B(new_n1573), .Y(new_n1575));
  nand_5 g01199(.A(new_n1398), .B(new_n1397), .Y(new_n1576));
  nand_5 g01200(.A(new_n1399), .B(new_n1394), .Y(new_n1577));
  nand_5 g01201(.A(new_n1577), .B(new_n1576), .Y(new_n1578));
  nand_5 g01202(.A(pi097), .B(pi041), .Y(new_n1579));
  nand_5 g01203(.A(pi182), .B(pi075), .Y(new_n1580));
  and_6  g01204(.A(new_n1580), .B(new_n1579), .Y(new_n1581));
  nand_5 g01205(.A(pi075), .B(pi041), .Y(new_n1582));
  nor_5  g01206(.A(new_n1582), .B(new_n1398), .Y(new_n1583));
  or_6   g01207(.A(new_n1583), .B(new_n1581), .Y(new_n1584));
  nand_5 g01208(.A(pi216), .B(pi019), .Y(new_n1585));
  nand_5 g01209(.A(new_n1392), .B(new_n1391), .Y(new_n1586));
  nand_5 g01210(.A(new_n1393), .B(new_n1390), .Y(new_n1587));
  nand_5 g01211(.A(new_n1587), .B(new_n1586), .Y(new_n1588));
  nand_5 g01212(.A(pi147), .B(pi079), .Y(new_n1589));
  nand_5 g01213(.A(pi151), .B(pi076), .Y(new_n1590));
  nand_5 g01214(.A(new_n1590), .B(new_n1589), .Y(new_n1591));
  nand_5 g01215(.A(pi151), .B(pi079), .Y(new_n1592));
  nor_5  g01216(.A(new_n1592), .B(new_n1392), .Y(new_n1593));
  not_8  g01217(.A(new_n1593), .Y(new_n1594));
  nand_5 g01218(.A(new_n1594), .B(new_n1591), .Y(new_n1595));
  xor_4  g01219(.A(new_n1595), .B(new_n1588), .Y(new_n1596));
  xor_4  g01220(.A(new_n1596), .B(new_n1585), .Y(new_n1597));
  xor_4  g01221(.A(new_n1597), .B(new_n1584), .Y(new_n1598));
  not_8  g01222(.A(new_n1598), .Y(new_n1599));
  xor_4  g01223(.A(new_n1599), .B(new_n1578), .Y(new_n1600));
  not_8  g01224(.A(new_n1405), .Y(new_n1601));
  nor_5  g01225(.A(new_n1601), .B(new_n1401), .Y(new_n1602));
  nor_5  g01226(.A(new_n1406), .B(new_n1400), .Y(new_n1603));
  nor_5  g01227(.A(new_n1603), .B(new_n1602), .Y(new_n1604));
  xor_4  g01228(.A(new_n1604), .B(new_n1600), .Y(new_n1605));
  xor_4  g01229(.A(new_n1605), .B(new_n1575), .Y(new_n1606));
  xnor_4 g01230(.A(new_n1606), .B(new_n1572), .Y(new_n1607));
  xor_4  g01231(.A(new_n1607), .B(new_n1499), .Y(new_n1608));
  nor_5  g01232(.A(new_n1608), .B(new_n1496), .Y(new_n1609));
  or_6   g01233(.A(new_n1609), .B(new_n1495), .Y(new_n1610));
  not_8  g01234(.A(new_n1490), .Y(new_n1611));
  nand_5 g01235(.A(new_n1491), .B(new_n1611), .Y(new_n1612));
  not_8  g01236(.A(new_n1612), .Y(new_n1613));
  nor_5  g01237(.A(new_n1492), .B(new_n1489), .Y(new_n1614));
  nor_5  g01238(.A(new_n1614), .B(new_n1613), .Y(new_n1615));
  nor_5  g01239(.A(new_n1488), .B(new_n1463), .Y(new_n1616));
  nand_5 g01240(.A(pi177), .B(pi119), .Y(new_n1617));
  xor_4  g01241(.A(new_n1617), .B(new_n1471), .Y(new_n1618));
  nand_5 g01242(.A(pi250), .B(pi101), .Y(new_n1619));
  xor_4  g01243(.A(new_n1619), .B(new_n1618), .Y(new_n1620));
  nand_5 g01244(.A(pi223), .B(pi044), .Y(new_n1621));
  xor_4  g01245(.A(new_n1621), .B(new_n1472), .Y(new_n1622));
  xnor_4 g01246(.A(new_n1622), .B(new_n1620), .Y(new_n1623));
  nand_5 g01247(.A(new_n1474), .B(new_n1467), .Y(new_n1624));
  nand_5 g01248(.A(new_n1475), .B(new_n1464), .Y(new_n1625));
  nand_5 g01249(.A(new_n1625), .B(new_n1624), .Y(new_n1626));
  nand_5 g01250(.A(pi248), .B(pi160), .Y(new_n1627));
  nand_5 g01251(.A(pi072), .B(pi020), .Y(new_n1628));
  xor_4  g01252(.A(new_n1628), .B(new_n1627), .Y(new_n1629));
  xor_4  g01253(.A(new_n1629), .B(new_n1483), .Y(new_n1630));
  xnor_4 g01254(.A(new_n1630), .B(new_n1626), .Y(new_n1631));
  xor_4  g01255(.A(new_n1631), .B(new_n1623), .Y(new_n1632));
  not_8  g01256(.A(new_n1632), .Y(new_n1633));
  nand_5 g01257(.A(new_n1486), .B(new_n1479), .Y(new_n1634));
  nand_5 g01258(.A(new_n1487), .B(new_n1476), .Y(new_n1635));
  nand_5 g01259(.A(new_n1635), .B(new_n1634), .Y(new_n1636));
  xor_4  g01260(.A(new_n1636), .B(new_n1484), .Y(new_n1637));
  xor_4  g01261(.A(new_n1637), .B(new_n1633), .Y(new_n1638));
  xor_4  g01262(.A(new_n1638), .B(new_n1616), .Y(new_n1639));
  xnor_4 g01263(.A(new_n1639), .B(new_n1615), .Y(new_n1640));
  nor_5  g01264(.A(new_n1640), .B(new_n1610), .Y(new_n1641));
  nor_5  g01265(.A(new_n1606), .B(new_n1572), .Y(new_n1642));
  nor_5  g01266(.A(new_n1607), .B(new_n1499), .Y(new_n1643));
  or_6   g01267(.A(new_n1643), .B(new_n1642), .Y(new_n1644));
  nand_5 g01268(.A(new_n1574), .B(new_n1573), .Y(new_n1645));
  nand_5 g01269(.A(new_n1605), .B(new_n1575), .Y(new_n1646));
  nand_5 g01270(.A(new_n1646), .B(new_n1645), .Y(new_n1647));
  not_8  g01271(.A(new_n1600), .Y(new_n1648));
  nor_5  g01272(.A(new_n1604), .B(new_n1648), .Y(new_n1649));
  nand_5 g01273(.A(pi216), .B(pi097), .Y(new_n1650));
  xor_4  g01274(.A(new_n1650), .B(new_n1593), .Y(new_n1651));
  nand_5 g01275(.A(pi251), .B(pi147), .Y(new_n1652));
  nand_5 g01276(.A(pi076), .B(pi019), .Y(new_n1653));
  xor_4  g01277(.A(new_n1653), .B(new_n1652), .Y(new_n1654));
  xor_4  g01278(.A(new_n1654), .B(new_n1592), .Y(new_n1655));
  xor_4  g01279(.A(new_n1655), .B(new_n1651), .Y(new_n1656));
  not_8  g01280(.A(new_n1656), .Y(new_n1657));
  nand_5 g01281(.A(new_n1595), .B(new_n1588), .Y(new_n1658));
  nand_5 g01282(.A(new_n1596), .B(new_n1585), .Y(new_n1659));
  nand_5 g01283(.A(new_n1659), .B(new_n1658), .Y(new_n1660));
  nand_5 g01284(.A(pi166), .B(pi138), .Y(new_n1661));
  nand_5 g01285(.A(pi182), .B(pi093), .Y(new_n1662));
  xor_4  g01286(.A(new_n1662), .B(new_n1661), .Y(new_n1663));
  xor_4  g01287(.A(new_n1663), .B(new_n1582), .Y(new_n1664));
  xor_4  g01288(.A(new_n1664), .B(new_n1660), .Y(new_n1665));
  xor_4  g01289(.A(new_n1665), .B(new_n1657), .Y(new_n1666));
  nor_5  g01290(.A(new_n1599), .B(new_n1578), .Y(new_n1667));
  and_6  g01291(.A(new_n1667), .B(new_n1583), .Y(new_n1668));
  nor_5  g01292(.A(new_n1597), .B(new_n1584), .Y(new_n1669));
  nor_5  g01293(.A(new_n1669), .B(new_n1583), .Y(new_n1670));
  not_8  g01294(.A(new_n1670), .Y(new_n1671));
  nor_5  g01295(.A(new_n1671), .B(new_n1667), .Y(new_n1672));
  or_6   g01296(.A(new_n1672), .B(new_n1668), .Y(new_n1673));
  xor_4  g01297(.A(new_n1673), .B(new_n1666), .Y(new_n1674));
  xor_4  g01298(.A(new_n1674), .B(new_n1649), .Y(new_n1675));
  xor_4  g01299(.A(new_n1675), .B(new_n1647), .Y(new_n1676));
  not_8  g01300(.A(new_n1676), .Y(new_n1677));
  xor_4  g01301(.A(new_n1677), .B(new_n1644), .Y(new_n1678));
  or_6   g01302(.A(new_n1570), .B(new_n1537), .Y(new_n1679));
  nand_5 g01303(.A(new_n1571), .B(new_n1533), .Y(new_n1680));
  nand_5 g01304(.A(new_n1680), .B(new_n1679), .Y(new_n1681));
  not_8  g01305(.A(new_n1538), .Y(new_n1682));
  nand_5 g01306(.A(new_n1539), .B(new_n1682), .Y(new_n1683));
  not_8  g01307(.A(new_n1540), .Y(new_n1684));
  nand_5 g01308(.A(new_n1569), .B(new_n1684), .Y(new_n1685));
  nand_5 g01309(.A(new_n1685), .B(new_n1683), .Y(new_n1686));
  not_8  g01310(.A(new_n1544), .Y(new_n1687));
  nor_5  g01311(.A(new_n1568), .B(new_n1687), .Y(new_n1688));
  nand_5 g01312(.A(pi056), .B(pi001), .Y(new_n1689));
  xor_4  g01313(.A(new_n1689), .B(new_n1560), .Y(new_n1690));
  nand_5 g01314(.A(pi122), .B(pi008), .Y(new_n1691));
  nand_5 g01315(.A(pi059), .B(pi027), .Y(new_n1692));
  xor_4  g01316(.A(new_n1692), .B(new_n1691), .Y(new_n1693));
  xor_4  g01317(.A(new_n1693), .B(new_n1558), .Y(new_n1694));
  xor_4  g01318(.A(new_n1694), .B(new_n1690), .Y(new_n1695));
  nand_5 g01319(.A(new_n1561), .B(new_n1554), .Y(new_n1696));
  nand_5 g01320(.A(new_n1562), .B(new_n1553), .Y(new_n1697));
  nand_5 g01321(.A(new_n1697), .B(new_n1696), .Y(new_n1698));
  nand_5 g01322(.A(pi235), .B(pi087), .Y(new_n1699));
  nand_5 g01323(.A(pi219), .B(pi096), .Y(new_n1700));
  xor_4  g01324(.A(new_n1700), .B(new_n1548), .Y(new_n1701));
  xor_4  g01325(.A(new_n1701), .B(new_n1699), .Y(new_n1702));
  xor_4  g01326(.A(new_n1702), .B(new_n1698), .Y(new_n1703));
  xor_4  g01327(.A(new_n1703), .B(new_n1695), .Y(new_n1704));
  nor_5  g01328(.A(new_n1563), .B(new_n1550), .Y(new_n1705));
  not_8  g01329(.A(new_n1564), .Y(new_n1706));
  nor_5  g01330(.A(new_n1567), .B(new_n1706), .Y(new_n1707));
  xor_4  g01331(.A(new_n1707), .B(new_n1549), .Y(new_n1708));
  nor_5  g01332(.A(new_n1708), .B(new_n1705), .Y(new_n1709));
  xor_4  g01333(.A(new_n1709), .B(new_n1704), .Y(new_n1710));
  xor_4  g01334(.A(new_n1710), .B(new_n1688), .Y(new_n1711));
  xor_4  g01335(.A(new_n1711), .B(new_n1686), .Y(new_n1712));
  xnor_4 g01336(.A(new_n1712), .B(new_n1681), .Y(new_n1713));
  not_8  g01337(.A(new_n1503), .Y(new_n1714));
  or_6   g01338(.A(new_n1528), .B(new_n1714), .Y(new_n1715));
  nand_5 g01339(.A(pi114), .B(pi071), .Y(new_n1716));
  nand_5 g01340(.A(pi142), .B(pi091), .Y(new_n1717));
  xor_4  g01341(.A(new_n1717), .B(new_n1716), .Y(new_n1718));
  xor_4  g01342(.A(new_n1718), .B(new_n1510), .Y(new_n1719));
  nand_5 g01343(.A(new_n1524), .B(new_n1521), .Y(new_n1720));
  nand_5 g01344(.A(new_n1525), .B(new_n1520), .Y(new_n1721));
  nand_5 g01345(.A(new_n1721), .B(new_n1720), .Y(new_n1722));
  xor_4  g01346(.A(new_n1722), .B(new_n1719), .Y(new_n1723));
  nand_5 g01347(.A(pi145), .B(pi123), .Y(new_n1724));
  xor_4  g01348(.A(new_n1724), .B(new_n1519), .Y(new_n1725));
  nand_5 g01349(.A(pi099), .B(pi032), .Y(new_n1726));
  nand_5 g01350(.A(pi164), .B(pi155), .Y(new_n1727));
  xor_4  g01351(.A(new_n1727), .B(new_n1517), .Y(new_n1728));
  xnor_4 g01352(.A(new_n1728), .B(new_n1726), .Y(new_n1729));
  xnor_4 g01353(.A(new_n1729), .B(new_n1725), .Y(new_n1730));
  xnor_4 g01354(.A(new_n1730), .B(new_n1723), .Y(new_n1731));
  nand_5 g01355(.A(new_n1526), .B(new_n1513), .Y(new_n1732));
  nand_5 g01356(.A(new_n1527), .B(new_n1506), .Y(new_n1733));
  nand_5 g01357(.A(new_n1733), .B(new_n1732), .Y(new_n1734));
  xor_4  g01358(.A(new_n1734), .B(new_n1512), .Y(new_n1735));
  xor_4  g01359(.A(new_n1735), .B(new_n1731), .Y(new_n1736));
  xor_4  g01360(.A(new_n1736), .B(new_n1715), .Y(new_n1737));
  nand_5 g01361(.A(new_n1531), .B(new_n1530), .Y(new_n1738));
  nand_5 g01362(.A(new_n1532), .B(new_n1529), .Y(new_n1739));
  nand_5 g01363(.A(new_n1739), .B(new_n1738), .Y(new_n1740));
  xor_4  g01364(.A(new_n1740), .B(new_n1737), .Y(new_n1741));
  xor_4  g01365(.A(new_n1741), .B(new_n1713), .Y(new_n1742));
  xor_4  g01366(.A(new_n1742), .B(new_n1678), .Y(new_n1743));
  xnor_4 g01367(.A(new_n1640), .B(new_n1610), .Y(new_n1744));
  nor_5  g01368(.A(new_n1744), .B(new_n1743), .Y(new_n1745));
  nor_5  g01369(.A(new_n1745), .B(new_n1641), .Y(new_n1746));
  nand_5 g01370(.A(new_n1692), .B(new_n1691), .Y(new_n1747));
  nand_5 g01371(.A(new_n1693), .B(new_n1558), .Y(new_n1748));
  nand_5 g01372(.A(new_n1748), .B(new_n1747), .Y(new_n1749));
  nand_5 g01373(.A(pi079), .B(pi019), .Y(new_n1750));
  nand_5 g01374(.A(pi182), .B(pi166), .Y(new_n1751));
  xor_4  g01375(.A(new_n1751), .B(new_n1750), .Y(new_n1752));
  xor_4  g01376(.A(new_n1752), .B(new_n1749), .Y(new_n1753));
  xor_4  g01377(.A(new_n1753), .B(new_n1746), .Y(new_n1754));
  nand_5 g01378(.A(pi251), .B(pi151), .Y(new_n1755));
  nand_5 g01379(.A(pi032), .B(pi023), .Y(new_n1756));
  xor_4  g01380(.A(new_n1756), .B(new_n1755), .Y(new_n1757));
  nand_5 g01381(.A(pi164), .B(pi086), .Y(new_n1758));
  nand_5 g01382(.A(new_n1664), .B(new_n1660), .Y(new_n1759));
  nand_5 g01383(.A(new_n1665), .B(new_n1657), .Y(new_n1760));
  nand_5 g01384(.A(new_n1760), .B(new_n1759), .Y(new_n1761));
  xor_4  g01385(.A(new_n1761), .B(new_n1758), .Y(new_n1762));
  not_8  g01386(.A(new_n1666), .Y(new_n1763));
  nor_5  g01387(.A(new_n1673), .B(new_n1763), .Y(new_n1764));
  nor_5  g01388(.A(new_n1764), .B(new_n1672), .Y(new_n1765));
  xor_4  g01389(.A(new_n1765), .B(new_n1762), .Y(new_n1766));
  xor_4  g01390(.A(new_n1766), .B(new_n1757), .Y(new_n1767));
  nand_5 g01391(.A(pi138), .B(pi011), .Y(new_n1768));
  nand_5 g01392(.A(new_n1628), .B(new_n1627), .Y(new_n1769));
  nand_5 g01393(.A(new_n1629), .B(new_n1483), .Y(new_n1770));
  nand_5 g01394(.A(new_n1770), .B(new_n1769), .Y(new_n1771));
  xor_4  g01395(.A(new_n1771), .B(new_n1768), .Y(new_n1772));
  nand_5 g01396(.A(pi097), .B(pi076), .Y(new_n1773));
  nand_5 g01397(.A(pi248), .B(pi020), .Y(new_n1774));
  nand_5 g01398(.A(pi216), .B(pi075), .Y(new_n1775));
  xor_4  g01399(.A(new_n1775), .B(new_n1774), .Y(new_n1776));
  xor_4  g01400(.A(new_n1776), .B(new_n1773), .Y(new_n1777));
  xor_4  g01401(.A(new_n1777), .B(new_n1772), .Y(new_n1778));
  xor_4  g01402(.A(new_n1778), .B(new_n1767), .Y(new_n1779));
  xor_4  g01403(.A(new_n1779), .B(new_n1754), .Y(new_n1780));
  xor_4  g01404(.A(new_n1780), .B(new_n1217), .Y(new_n1781));
  or_6   g01405(.A(new_n1724), .B(new_n1519), .Y(new_n1782));
  nand_5 g01406(.A(new_n1729), .B(new_n1725), .Y(new_n1783));
  nand_5 g01407(.A(new_n1783), .B(new_n1782), .Y(new_n1784));
  nand_5 g01408(.A(new_n1702), .B(new_n1698), .Y(new_n1785));
  nand_5 g01409(.A(new_n1703), .B(new_n1695), .Y(new_n1786));
  nand_5 g01410(.A(new_n1786), .B(new_n1785), .Y(new_n1787));
  xor_4  g01411(.A(new_n1787), .B(new_n1784), .Y(new_n1788));
  nand_5 g01412(.A(new_n1617), .B(new_n1471), .Y(new_n1789));
  nand_5 g01413(.A(new_n1619), .B(new_n1618), .Y(new_n1790));
  nand_5 g01414(.A(new_n1790), .B(new_n1789), .Y(new_n1791));
  nand_5 g01415(.A(new_n1722), .B(new_n1719), .Y(new_n1792));
  nand_5 g01416(.A(new_n1730), .B(new_n1723), .Y(new_n1793));
  nand_5 g01417(.A(new_n1793), .B(new_n1792), .Y(new_n1794));
  xor_4  g01418(.A(new_n1794), .B(new_n1791), .Y(new_n1795));
  xor_4  g01419(.A(new_n1795), .B(new_n1788), .Y(new_n1796));
  nand_5 g01420(.A(new_n1700), .B(new_n1548), .Y(new_n1797));
  nand_5 g01421(.A(new_n1701), .B(new_n1699), .Y(new_n1798));
  nand_5 g01422(.A(new_n1798), .B(new_n1797), .Y(new_n1799));
  nand_5 g01423(.A(pi091), .B(pi071), .Y(new_n1800));
  nand_5 g01424(.A(pi094), .B(pi027), .Y(new_n1801));
  xor_4  g01425(.A(new_n1801), .B(new_n1800), .Y(new_n1802));
  xor_4  g01426(.A(new_n1802), .B(new_n1799), .Y(new_n1803));
  and_6  g01427(.A(new_n1707), .B(new_n1549), .Y(new_n1804));
  nor_5  g01428(.A(new_n1709), .B(new_n1704), .Y(new_n1805));
  nor_5  g01429(.A(new_n1805), .B(new_n1804), .Y(new_n1806));
  xor_4  g01430(.A(new_n1806), .B(new_n1803), .Y(new_n1807));
  nor_5  g01431(.A(new_n1621), .B(new_n1473), .Y(new_n1808));
  nor_5  g01432(.A(new_n1622), .B(new_n1620), .Y(new_n1809));
  nor_5  g01433(.A(new_n1809), .B(new_n1808), .Y(new_n1810));
  nand_5 g01434(.A(pi136), .B(pi001), .Y(new_n1811));
  xor_4  g01435(.A(new_n1811), .B(new_n1810), .Y(new_n1812));
  nand_5 g01436(.A(pi169), .B(pi114), .Y(new_n1813));
  nand_5 g01437(.A(new_n1717), .B(new_n1716), .Y(new_n1814));
  nand_5 g01438(.A(new_n1718), .B(new_n1510), .Y(new_n1815));
  nand_5 g01439(.A(new_n1815), .B(new_n1814), .Y(new_n1816));
  xor_4  g01440(.A(new_n1816), .B(new_n1813), .Y(new_n1817));
  xor_4  g01441(.A(new_n1817), .B(new_n1812), .Y(new_n1818));
  xor_4  g01442(.A(new_n1818), .B(new_n1807), .Y(new_n1819));
  xor_4  g01443(.A(new_n1819), .B(new_n1796), .Y(new_n1820));
  nand_5 g01444(.A(new_n1727), .B(new_n1517), .Y(new_n1821));
  nand_5 g01445(.A(new_n1728), .B(new_n1726), .Y(new_n1822));
  nand_5 g01446(.A(new_n1822), .B(new_n1821), .Y(new_n1823));
  nand_5 g01447(.A(pi110), .B(pi087), .Y(new_n1824));
  and_6  g01448(.A(new_n1674), .B(new_n1649), .Y(new_n1825));
  not_8  g01449(.A(new_n1675), .Y(new_n1826));
  nor_5  g01450(.A(new_n1826), .B(new_n1647), .Y(new_n1827));
  nor_5  g01451(.A(new_n1827), .B(new_n1825), .Y(new_n1828));
  xor_4  g01452(.A(new_n1828), .B(new_n1824), .Y(new_n1829));
  xor_4  g01453(.A(new_n1829), .B(new_n1823), .Y(new_n1830));
  xor_4  g01454(.A(new_n1830), .B(new_n1820), .Y(new_n1831));
  nand_5 g01455(.A(new_n1653), .B(new_n1652), .Y(new_n1832));
  nand_5 g01456(.A(new_n1654), .B(new_n1592), .Y(new_n1833));
  nand_5 g01457(.A(new_n1833), .B(new_n1832), .Y(new_n1834));
  nand_5 g01458(.A(pi160), .B(pi009), .Y(new_n1835));
  nand_5 g01459(.A(pi246), .B(pi123), .Y(new_n1836));
  xor_4  g01460(.A(new_n1836), .B(new_n1835), .Y(new_n1837));
  nand_5 g01461(.A(pi145), .B(pi099), .Y(new_n1838));
  xor_4  g01462(.A(new_n1838), .B(new_n1837), .Y(new_n1839));
  xor_4  g01463(.A(new_n1839), .B(new_n1834), .Y(new_n1840));
  xor_4  g01464(.A(new_n1840), .B(new_n1831), .Y(new_n1841));
  nand_5 g01465(.A(pi192), .B(pi147), .Y(new_n1842));
  nand_5 g01466(.A(pi250), .B(pi225), .Y(new_n1843));
  xor_4  g01467(.A(new_n1843), .B(new_n1842), .Y(new_n1844));
  nand_5 g01468(.A(new_n1638), .B(new_n1616), .Y(new_n1845));
  nand_5 g01469(.A(new_n1639), .B(new_n1615), .Y(new_n1846));
  nand_5 g01470(.A(new_n1846), .B(new_n1845), .Y(new_n1847));
  xor_4  g01471(.A(new_n1847), .B(new_n1844), .Y(new_n1848));
  nand_5 g01472(.A(pi135), .B(pi008), .Y(new_n1849));
  nand_5 g01473(.A(pi059), .B(pi026), .Y(new_n1850));
  nand_5 g01474(.A(pi223), .B(pi054), .Y(new_n1851));
  or_6   g01475(.A(new_n1689), .B(new_n1560), .Y(new_n1852));
  not_8  g01476(.A(new_n1694), .Y(new_n1853));
  nand_5 g01477(.A(new_n1853), .B(new_n1690), .Y(new_n1854));
  nand_5 g01478(.A(new_n1854), .B(new_n1852), .Y(new_n1855));
  xor_4  g01479(.A(new_n1855), .B(new_n1851), .Y(new_n1856));
  xor_4  g01480(.A(new_n1856), .B(new_n1850), .Y(new_n1857));
  xor_4  g01481(.A(new_n1857), .B(new_n1849), .Y(new_n1858));
  xor_4  g01482(.A(new_n1858), .B(new_n1848), .Y(new_n1859));
  nand_5 g01483(.A(pi122), .B(pi056), .Y(new_n1860));
  nor_5  g01484(.A(new_n1636), .B(new_n1485), .Y(new_n1861));
  nor_5  g01485(.A(new_n1637), .B(new_n1633), .Y(new_n1862));
  or_6   g01486(.A(new_n1862), .B(new_n1861), .Y(new_n1863));
  nand_5 g01487(.A(pi102), .B(pi096), .Y(new_n1864));
  nand_5 g01488(.A(pi235), .B(pi219), .Y(new_n1865));
  xor_4  g01489(.A(new_n1865), .B(new_n1864), .Y(new_n1866));
  xor_4  g01490(.A(new_n1866), .B(new_n1863), .Y(new_n1867));
  xor_4  g01491(.A(new_n1867), .B(new_n1860), .Y(new_n1868));
  xor_4  g01492(.A(new_n1868), .B(new_n1859), .Y(new_n1869));
  xor_4  g01493(.A(new_n1869), .B(new_n1841), .Y(new_n1870));
  nand_5 g01494(.A(pi177), .B(pi045), .Y(new_n1871));
  nand_5 g01495(.A(pi142), .B(pi031), .Y(new_n1872));
  xor_4  g01496(.A(new_n1872), .B(new_n1871), .Y(new_n1873));
  nand_5 g01497(.A(pi101), .B(pi044), .Y(new_n1874));
  nand_5 g01498(.A(pi206), .B(pi155), .Y(new_n1875));
  nand_5 g01499(.A(pi072), .B(pi060), .Y(new_n1876));
  xor_4  g01500(.A(new_n1876), .B(new_n1875), .Y(new_n1877));
  xor_4  g01501(.A(new_n1877), .B(new_n1874), .Y(new_n1878));
  nand_5 g01502(.A(new_n1662), .B(new_n1661), .Y(new_n1879));
  nand_5 g01503(.A(new_n1663), .B(new_n1582), .Y(new_n1880));
  nand_5 g01504(.A(new_n1880), .B(new_n1879), .Y(new_n1881));
  nor_5  g01505(.A(new_n1650), .B(new_n1594), .Y(new_n1882));
  nor_5  g01506(.A(new_n1655), .B(new_n1651), .Y(new_n1883));
  nor_5  g01507(.A(new_n1883), .B(new_n1882), .Y(new_n1884));
  xor_4  g01508(.A(new_n1884), .B(new_n1881), .Y(new_n1885));
  nand_5 g01509(.A(pi137), .B(pi119), .Y(new_n1886));
  nor_5  g01510(.A(new_n1710), .B(new_n1688), .Y(new_n1887));
  and_6  g01511(.A(new_n1711), .B(new_n1686), .Y(new_n1888));
  nor_5  g01512(.A(new_n1888), .B(new_n1887), .Y(new_n1889));
  xor_4  g01513(.A(new_n1889), .B(new_n1886), .Y(new_n1890));
  xor_4  g01514(.A(new_n1890), .B(new_n1885), .Y(new_n1891));
  xor_4  g01515(.A(new_n1891), .B(new_n1878), .Y(new_n1892));
  xor_4  g01516(.A(new_n1892), .B(new_n1873), .Y(new_n1893));
  xor_4  g01517(.A(new_n1893), .B(new_n1870), .Y(new_n1894));
  not_8  g01518(.A(new_n1736), .Y(new_n1895));
  nor_5  g01519(.A(new_n1895), .B(new_n1715), .Y(new_n1896));
  nor_5  g01520(.A(new_n1740), .B(new_n1737), .Y(new_n1897));
  nor_5  g01521(.A(new_n1897), .B(new_n1896), .Y(new_n1898));
  or_6   g01522(.A(new_n1677), .B(new_n1644), .Y(new_n1899));
  nand_5 g01523(.A(new_n1742), .B(new_n1678), .Y(new_n1900));
  nand_5 g01524(.A(new_n1900), .B(new_n1899), .Y(new_n1901));
  xor_4  g01525(.A(new_n1901), .B(new_n1898), .Y(new_n1902));
  nor_5  g01526(.A(new_n1712), .B(new_n1681), .Y(new_n1903));
  not_8  g01527(.A(new_n1741), .Y(new_n1904));
  nor_5  g01528(.A(new_n1904), .B(new_n1713), .Y(new_n1905));
  nor_5  g01529(.A(new_n1905), .B(new_n1903), .Y(new_n1906));
  xor_4  g01530(.A(new_n1906), .B(new_n1902), .Y(new_n1907));
  or_6   g01531(.A(new_n1734), .B(new_n1512), .Y(new_n1908));
  nand_5 g01532(.A(new_n1735), .B(new_n1731), .Y(new_n1909));
  nand_5 g01533(.A(new_n1909), .B(new_n1908), .Y(new_n1910));
  nor_5  g01534(.A(new_n1630), .B(new_n1626), .Y(new_n1911));
  nor_5  g01535(.A(new_n1631), .B(new_n1623), .Y(new_n1912));
  nor_5  g01536(.A(new_n1912), .B(new_n1911), .Y(new_n1913));
  xor_4  g01537(.A(new_n1913), .B(new_n1910), .Y(new_n1914));
  xor_4  g01538(.A(new_n1914), .B(new_n1907), .Y(new_n1915));
  xor_4  g01539(.A(new_n1915), .B(new_n1894), .Y(new_n1916));
  xor_4  g01540(.A(new_n1916), .B(new_n1781), .Y(po005));
  nand_5 g01541(.A(pi175), .B(pi165), .Y(new_n1918));
  nand_5 g01542(.A(pi134), .B(pi062), .Y(new_n1919));
  nand_5 g01543(.A(pi175), .B(pi120), .Y(new_n1920));
  nand_5 g01544(.A(pi240), .B(pi065), .Y(new_n1921));
  or_6   g01545(.A(new_n1921), .B(new_n1920), .Y(new_n1922));
  nand_5 g01546(.A(new_n1922), .B(new_n1919), .Y(new_n1923));
  nand_5 g01547(.A(new_n1921), .B(new_n1920), .Y(new_n1924));
  nand_5 g01548(.A(new_n1924), .B(new_n1923), .Y(new_n1925));
  nand_5 g01549(.A(pi175), .B(pi172), .Y(new_n1926));
  nor_5  g01550(.A(new_n1926), .B(new_n1925), .Y(new_n1927));
  nand_5 g01551(.A(pi134), .B(pi120), .Y(new_n1928));
  nand_5 g01552(.A(pi149), .B(pi065), .Y(new_n1929));
  not_8  g01553(.A(pi062), .Y(new_n1930));
  not_8  g01554(.A(pi240), .Y(new_n1931));
  nor_5  g01555(.A(new_n1931), .B(new_n1930), .Y(new_n1932));
  xor_4  g01556(.A(new_n1932), .B(new_n1929), .Y(new_n1933));
  xor_4  g01557(.A(new_n1933), .B(new_n1928), .Y(new_n1934));
  xor_4  g01558(.A(new_n1926), .B(new_n1925), .Y(new_n1935));
  nand_5 g01559(.A(new_n1935), .B(new_n1934), .Y(new_n1936));
  not_8  g01560(.A(new_n1936), .Y(new_n1937));
  nor_5  g01561(.A(new_n1937), .B(new_n1927), .Y(new_n1938));
  nand_5 g01562(.A(pi198), .B(pi175), .Y(new_n1939));
  nand_5 g01563(.A(pi167), .B(pi065), .Y(new_n1940));
  nand_5 g01564(.A(pi240), .B(pi120), .Y(new_n1941));
  nand_5 g01565(.A(pi149), .B(pi062), .Y(new_n1942));
  xor_4  g01566(.A(new_n1942), .B(new_n1941), .Y(new_n1943));
  xor_4  g01567(.A(new_n1943), .B(new_n1940), .Y(new_n1944));
  nand_5 g01568(.A(pi172), .B(pi134), .Y(new_n1945));
  not_8  g01569(.A(new_n1929), .Y(new_n1946));
  nor_5  g01570(.A(new_n1932), .B(new_n1946), .Y(new_n1947));
  not_8  g01571(.A(new_n1928), .Y(new_n1948));
  nor_5  g01572(.A(new_n1933), .B(new_n1948), .Y(new_n1949));
  or_6   g01573(.A(new_n1949), .B(new_n1947), .Y(new_n1950));
  xor_4  g01574(.A(new_n1950), .B(new_n1945), .Y(new_n1951));
  xor_4  g01575(.A(new_n1951), .B(new_n1944), .Y(new_n1952));
  xnor_4 g01576(.A(new_n1952), .B(new_n1939), .Y(new_n1953));
  xor_4  g01577(.A(new_n1953), .B(new_n1938), .Y(new_n1954));
  nand_5 g01578(.A(pi175), .B(pi065), .Y(new_n1955));
  not_8  g01579(.A(new_n1955), .Y(new_n1956));
  nor_5  g01580(.A(new_n1956), .B(new_n1919), .Y(new_n1957));
  or_6   g01581(.A(new_n1957), .B(new_n1924), .Y(new_n1958));
  and_6  g01582(.A(new_n1958), .B(new_n1922), .Y(new_n1959));
  nor_5  g01583(.A(new_n1959), .B(new_n1919), .Y(new_n1960));
  not_8  g01584(.A(new_n1960), .Y(new_n1961));
  xnor_4 g01585(.A(new_n1935), .B(new_n1934), .Y(new_n1962));
  nor_5  g01586(.A(new_n1962), .B(new_n1961), .Y(new_n1963));
  nand_5 g01587(.A(new_n1963), .B(new_n1954), .Y(new_n1964));
  xnor_4 g01588(.A(new_n1964), .B(new_n1918), .Y(new_n1965));
  nor_5  g01589(.A(new_n1952), .B(new_n1939), .Y(new_n1966));
  nor_5  g01590(.A(new_n1953), .B(new_n1938), .Y(new_n1967));
  nor_5  g01591(.A(new_n1967), .B(new_n1966), .Y(new_n1968));
  nand_5 g01592(.A(new_n1950), .B(new_n1945), .Y(new_n1969));
  nand_5 g01593(.A(new_n1951), .B(new_n1944), .Y(new_n1970));
  nand_5 g01594(.A(new_n1970), .B(new_n1969), .Y(new_n1971));
  nand_5 g01595(.A(pi240), .B(pi172), .Y(new_n1972));
  nand_5 g01596(.A(pi198), .B(pi134), .Y(new_n1973));
  nand_5 g01597(.A(new_n1973), .B(new_n1972), .Y(new_n1974));
  nand_5 g01598(.A(pi240), .B(pi198), .Y(new_n1975));
  nor_5  g01599(.A(new_n1975), .B(new_n1945), .Y(new_n1976));
  not_8  g01600(.A(new_n1976), .Y(new_n1977));
  nand_5 g01601(.A(new_n1977), .B(new_n1974), .Y(new_n1978));
  nand_5 g01602(.A(new_n1942), .B(new_n1941), .Y(new_n1979));
  nand_5 g01603(.A(new_n1943), .B(new_n1940), .Y(new_n1980));
  nand_5 g01604(.A(new_n1980), .B(new_n1979), .Y(new_n1981));
  nand_5 g01605(.A(pi149), .B(pi120), .Y(new_n1982));
  nand_5 g01606(.A(pi167), .B(pi062), .Y(new_n1983));
  nand_5 g01607(.A(pi181), .B(pi065), .Y(new_n1984));
  nand_5 g01608(.A(new_n1984), .B(new_n1983), .Y(new_n1985));
  nand_5 g01609(.A(pi181), .B(pi062), .Y(new_n1986));
  nor_5  g01610(.A(new_n1986), .B(new_n1940), .Y(new_n1987));
  not_8  g01611(.A(new_n1987), .Y(new_n1988));
  nand_5 g01612(.A(new_n1988), .B(new_n1985), .Y(new_n1989));
  xor_4  g01613(.A(new_n1989), .B(new_n1982), .Y(new_n1990));
  xor_4  g01614(.A(new_n1990), .B(new_n1981), .Y(new_n1991));
  xor_4  g01615(.A(new_n1991), .B(new_n1978), .Y(new_n1992));
  xor_4  g01616(.A(new_n1992), .B(new_n1971), .Y(new_n1993));
  xor_4  g01617(.A(new_n1993), .B(new_n1968), .Y(new_n1994));
  xnor_4 g01618(.A(new_n1994), .B(new_n1965), .Y(new_n1995));
  xnor_4 g01619(.A(new_n1963), .B(new_n1954), .Y(new_n1996));
  nand_5 g01620(.A(pi148), .B(pi004), .Y(new_n1997));
  nand_5 g01621(.A(pi163), .B(pi073), .Y(new_n1998));
  nand_5 g01622(.A(pi228), .B(pi170), .Y(new_n1999));
  nor_5  g01623(.A(new_n1999), .B(new_n1998), .Y(new_n2000));
  and_6  g01624(.A(pi170), .B(pi163), .Y(new_n2001));
  nor_5  g01625(.A(new_n2001), .B(new_n1997), .Y(new_n2002));
  nand_5 g01626(.A(new_n1999), .B(new_n1998), .Y(new_n2003));
  nor_5  g01627(.A(new_n2003), .B(new_n2002), .Y(new_n2004));
  nor_5  g01628(.A(new_n2004), .B(new_n2000), .Y(new_n2005));
  nor_5  g01629(.A(new_n2005), .B(new_n1997), .Y(new_n2006));
  nand_5 g01630(.A(pi170), .B(pi039), .Y(new_n2007));
  nand_5 g01631(.A(pi228), .B(pi004), .Y(new_n2008));
  nand_5 g01632(.A(pi148), .B(pi073), .Y(new_n2009));
  xor_4  g01633(.A(new_n2009), .B(new_n2008), .Y(new_n2010));
  xnor_4 g01634(.A(new_n2010), .B(new_n2007), .Y(new_n2011));
  not_8  g01635(.A(new_n1997), .Y(new_n2012));
  or_6   g01636(.A(new_n2000), .B(new_n2012), .Y(new_n2013));
  nand_5 g01637(.A(new_n2013), .B(new_n2003), .Y(new_n2014));
  nand_5 g01638(.A(pi163), .B(pi003), .Y(new_n2015));
  xnor_4 g01639(.A(new_n2015), .B(new_n2014), .Y(new_n2016));
  xnor_4 g01640(.A(new_n2016), .B(new_n2011), .Y(new_n2017));
  nand_5 g01641(.A(new_n2017), .B(new_n2006), .Y(new_n2018));
  nand_5 g01642(.A(pi163), .B(pi130), .Y(new_n2019));
  nand_5 g01643(.A(new_n2015), .B(new_n2014), .Y(new_n2020));
  or_6   g01644(.A(new_n2016), .B(new_n2011), .Y(new_n2021));
  nand_5 g01645(.A(new_n2021), .B(new_n2020), .Y(new_n2022));
  xnor_4 g01646(.A(new_n2022), .B(new_n2019), .Y(new_n2023));
  nand_5 g01647(.A(pi039), .B(pi004), .Y(new_n2024));
  nand_5 g01648(.A(pi228), .B(pi073), .Y(new_n2025));
  nand_5 g01649(.A(pi170), .B(pi116), .Y(new_n2026));
  xor_4  g01650(.A(new_n2026), .B(new_n2025), .Y(new_n2027));
  xor_4  g01651(.A(new_n2027), .B(new_n2024), .Y(new_n2028));
  nand_5 g01652(.A(pi148), .B(pi003), .Y(new_n2029));
  nand_5 g01653(.A(new_n2009), .B(new_n2008), .Y(new_n2030));
  nand_5 g01654(.A(new_n2010), .B(new_n2007), .Y(new_n2031));
  nand_5 g01655(.A(new_n2031), .B(new_n2030), .Y(new_n2032));
  xor_4  g01656(.A(new_n2032), .B(new_n2029), .Y(new_n2033));
  xor_4  g01657(.A(new_n2033), .B(new_n2028), .Y(new_n2034));
  xnor_4 g01658(.A(new_n2034), .B(new_n2023), .Y(new_n2035));
  xor_4  g01659(.A(new_n2035), .B(new_n2018), .Y(new_n2036));
  nand_5 g01660(.A(pi171), .B(pi158), .Y(new_n2037));
  nand_5 g01661(.A(pi254), .B(pi049), .Y(new_n2038));
  nand_5 g01662(.A(pi107), .B(pi089), .Y(new_n2039));
  nor_5  g01663(.A(new_n2039), .B(new_n2038), .Y(new_n2040));
  and_6  g01664(.A(pi254), .B(pi107), .Y(new_n2041));
  nor_5  g01665(.A(new_n2041), .B(new_n2037), .Y(new_n2042));
  nand_5 g01666(.A(new_n2039), .B(new_n2038), .Y(new_n2043));
  nor_5  g01667(.A(new_n2043), .B(new_n2042), .Y(new_n2044));
  nor_5  g01668(.A(new_n2044), .B(new_n2040), .Y(new_n2045));
  nor_5  g01669(.A(new_n2045), .B(new_n2037), .Y(new_n2046));
  nand_5 g01670(.A(pi158), .B(pi049), .Y(new_n2047));
  nand_5 g01671(.A(pi171), .B(pi089), .Y(new_n2048));
  nand_5 g01672(.A(pi254), .B(pi245), .Y(new_n2049));
  xor_4  g01673(.A(new_n2049), .B(new_n2048), .Y(new_n2050));
  xor_4  g01674(.A(new_n2050), .B(new_n2047), .Y(new_n2051));
  not_8  g01675(.A(new_n2037), .Y(new_n2052));
  or_6   g01676(.A(new_n2040), .B(new_n2052), .Y(new_n2053));
  nand_5 g01677(.A(new_n2053), .B(new_n2043), .Y(new_n2054));
  nand_5 g01678(.A(pi154), .B(pi107), .Y(new_n2055));
  xnor_4 g01679(.A(new_n2055), .B(new_n2054), .Y(new_n2056));
  xor_4  g01680(.A(new_n2056), .B(new_n2051), .Y(new_n2057));
  xor_4  g01681(.A(new_n2057), .B(new_n2046), .Y(new_n2058));
  nand_5 g01682(.A(new_n2043), .B(new_n2042), .Y(new_n2059));
  nand_5 g01683(.A(new_n2059), .B(new_n2045), .Y(new_n2060));
  nand_5 g01684(.A(new_n2003), .B(new_n2002), .Y(new_n2061));
  nand_5 g01685(.A(new_n2061), .B(new_n2005), .Y(new_n2062));
  nand_5 g01686(.A(new_n2062), .B(new_n2060), .Y(new_n2063));
  or_6   g01687(.A(new_n2062), .B(new_n2060), .Y(new_n2064));
  and_6  g01688(.A(new_n2041), .B(new_n2001), .Y(new_n2065));
  nand_5 g01689(.A(pi254), .B(pi171), .Y(new_n2066));
  nand_5 g01690(.A(pi158), .B(pi107), .Y(new_n2067));
  xor_4  g01691(.A(new_n2067), .B(new_n2066), .Y(new_n2068));
  nand_5 g01692(.A(new_n2068), .B(new_n2065), .Y(new_n2069));
  xor_4  g01693(.A(new_n2068), .B(new_n2065), .Y(new_n2070));
  nand_5 g01694(.A(pi163), .B(pi004), .Y(new_n2071));
  nand_5 g01695(.A(pi170), .B(pi148), .Y(new_n2072));
  xor_4  g01696(.A(new_n2072), .B(new_n2071), .Y(new_n2073));
  nand_5 g01697(.A(new_n2073), .B(new_n2070), .Y(new_n2074));
  and_6  g01698(.A(new_n2074), .B(new_n2069), .Y(new_n2075));
  nand_5 g01699(.A(new_n2075), .B(new_n2064), .Y(new_n2076));
  and_6  g01700(.A(new_n2076), .B(new_n2063), .Y(new_n2077));
  nor_5  g01701(.A(new_n2077), .B(new_n2058), .Y(new_n2078));
  xor_4  g01702(.A(new_n2017), .B(new_n2006), .Y(new_n2079));
  nand_5 g01703(.A(new_n2076), .B(new_n2063), .Y(new_n2080));
  xor_4  g01704(.A(new_n2080), .B(new_n2058), .Y(new_n2081));
  nor_5  g01705(.A(new_n2081), .B(new_n2079), .Y(new_n2082));
  nor_5  g01706(.A(new_n2082), .B(new_n2078), .Y(new_n2083));
  nand_5 g01707(.A(new_n2057), .B(new_n2046), .Y(new_n2084));
  nand_5 g01708(.A(pi171), .B(pi154), .Y(new_n2085));
  nand_5 g01709(.A(new_n2049), .B(new_n2048), .Y(new_n2086));
  nand_5 g01710(.A(new_n2050), .B(new_n2047), .Y(new_n2087));
  nand_5 g01711(.A(new_n2087), .B(new_n2086), .Y(new_n2088));
  xor_4  g01712(.A(new_n2088), .B(new_n2085), .Y(new_n2089));
  nand_5 g01713(.A(pi089), .B(pi049), .Y(new_n2090));
  nand_5 g01714(.A(pi254), .B(pi201), .Y(new_n2091));
  nand_5 g01715(.A(pi245), .B(pi158), .Y(new_n2092));
  xor_4  g01716(.A(new_n2092), .B(new_n2091), .Y(new_n2093));
  xor_4  g01717(.A(new_n2093), .B(new_n2090), .Y(new_n2094));
  xnor_4 g01718(.A(new_n2094), .B(new_n2089), .Y(new_n2095));
  nand_5 g01719(.A(pi107), .B(pi095), .Y(new_n2096));
  nor_5  g01720(.A(new_n2055), .B(new_n2054), .Y(new_n2097));
  nor_5  g01721(.A(new_n2056), .B(new_n2051), .Y(new_n2098));
  nor_5  g01722(.A(new_n2098), .B(new_n2097), .Y(new_n2099));
  xor_4  g01723(.A(new_n2099), .B(new_n2096), .Y(new_n2100));
  xor_4  g01724(.A(new_n2100), .B(new_n2095), .Y(new_n2101));
  xor_4  g01725(.A(new_n2101), .B(new_n2084), .Y(new_n2102));
  xor_4  g01726(.A(new_n2102), .B(new_n2083), .Y(new_n2103));
  xor_4  g01727(.A(new_n2103), .B(new_n2036), .Y(new_n2104));
  or_6   g01728(.A(new_n2104), .B(new_n1996), .Y(new_n2105));
  xor_4  g01729(.A(new_n2104), .B(new_n1996), .Y(new_n2106));
  xor_4  g01730(.A(new_n2081), .B(new_n2079), .Y(new_n2107));
  xor_4  g01731(.A(new_n1962), .B(new_n1960), .Y(new_n2108));
  nand_5 g01732(.A(new_n2108), .B(new_n2107), .Y(new_n2109));
  xor_4  g01733(.A(new_n2108), .B(new_n2107), .Y(new_n2110));
  nand_5 g01734(.A(new_n1957), .B(new_n1924), .Y(new_n2111));
  nand_5 g01735(.A(new_n2111), .B(new_n1959), .Y(new_n2112));
  nand_5 g01736(.A(new_n2064), .B(new_n2063), .Y(new_n2113));
  xnor_4 g01737(.A(new_n2113), .B(new_n2075), .Y(new_n2114));
  nor_5  g01738(.A(new_n2114), .B(new_n2112), .Y(new_n2115));
  nand_5 g01739(.A(pi175), .B(pi062), .Y(new_n2116));
  nand_5 g01740(.A(pi134), .B(pi065), .Y(new_n2117));
  xor_4  g01741(.A(new_n2117), .B(new_n2116), .Y(new_n2118));
  xnor_4 g01742(.A(new_n2041), .B(new_n2001), .Y(new_n2119));
  nor_5  g01743(.A(new_n2119), .B(new_n1955), .Y(new_n2120));
  nor_5  g01744(.A(new_n2120), .B(new_n2118), .Y(new_n2121));
  xnor_4 g01745(.A(new_n2120), .B(new_n2118), .Y(new_n2122));
  xor_4  g01746(.A(new_n2073), .B(new_n2070), .Y(new_n2123));
  nor_5  g01747(.A(new_n2123), .B(new_n2122), .Y(new_n2124));
  nor_5  g01748(.A(new_n2124), .B(new_n2121), .Y(new_n2125));
  xor_4  g01749(.A(new_n2114), .B(new_n2112), .Y(new_n2126));
  and_6  g01750(.A(new_n2126), .B(new_n2125), .Y(new_n2127));
  nor_5  g01751(.A(new_n2127), .B(new_n2115), .Y(new_n2128));
  nand_5 g01752(.A(new_n2128), .B(new_n2110), .Y(new_n2129));
  and_6  g01753(.A(new_n2129), .B(new_n2109), .Y(new_n2130));
  nand_5 g01754(.A(new_n2130), .B(new_n2106), .Y(new_n2131));
  nand_5 g01755(.A(new_n2131), .B(new_n2105), .Y(new_n2132));
  or_6   g01756(.A(new_n2132), .B(new_n1995), .Y(new_n2133));
  xor_4  g01757(.A(new_n2132), .B(new_n1995), .Y(new_n2134));
  nor_5  g01758(.A(new_n2035), .B(new_n2018), .Y(new_n2135));
  nor_5  g01759(.A(new_n2022), .B(new_n2019), .Y(new_n2136));
  nor_5  g01760(.A(new_n2034), .B(new_n2023), .Y(new_n2137));
  or_6   g01761(.A(new_n2137), .B(new_n2136), .Y(new_n2138));
  nand_5 g01762(.A(new_n2032), .B(new_n2029), .Y(new_n2139));
  nand_5 g01763(.A(new_n2033), .B(new_n2028), .Y(new_n2140));
  nand_5 g01764(.A(new_n2140), .B(new_n2139), .Y(new_n2141));
  nand_5 g01765(.A(pi148), .B(pi130), .Y(new_n2142));
  nand_5 g01766(.A(pi228), .B(pi003), .Y(new_n2143));
  and_6  g01767(.A(new_n2143), .B(new_n2142), .Y(new_n2144));
  nand_5 g01768(.A(pi228), .B(pi130), .Y(new_n2145));
  nor_5  g01769(.A(new_n2145), .B(new_n2029), .Y(new_n2146));
  or_6   g01770(.A(new_n2146), .B(new_n2144), .Y(new_n2147));
  nand_5 g01771(.A(pi170), .B(pi070), .Y(new_n2148));
  nand_5 g01772(.A(pi116), .B(pi004), .Y(new_n2149));
  nand_5 g01773(.A(new_n2149), .B(new_n2148), .Y(new_n2150));
  nand_5 g01774(.A(pi070), .B(pi004), .Y(new_n2151));
  nor_5  g01775(.A(new_n2151), .B(new_n2026), .Y(new_n2152));
  not_8  g01776(.A(new_n2152), .Y(new_n2153));
  nand_5 g01777(.A(new_n2153), .B(new_n2150), .Y(new_n2154));
  nand_5 g01778(.A(pi073), .B(pi039), .Y(new_n2155));
  nand_5 g01779(.A(new_n2026), .B(new_n2025), .Y(new_n2156));
  nand_5 g01780(.A(new_n2027), .B(new_n2024), .Y(new_n2157));
  nand_5 g01781(.A(new_n2157), .B(new_n2156), .Y(new_n2158));
  xor_4  g01782(.A(new_n2158), .B(new_n2155), .Y(new_n2159));
  xor_4  g01783(.A(new_n2159), .B(new_n2154), .Y(new_n2160));
  xnor_4 g01784(.A(new_n2160), .B(new_n2147), .Y(new_n2161));
  xor_4  g01785(.A(new_n2161), .B(new_n2141), .Y(new_n2162));
  xnor_4 g01786(.A(new_n2162), .B(new_n2138), .Y(new_n2163));
  nand_5 g01787(.A(pi163), .B(pi124), .Y(new_n2164));
  xor_4  g01788(.A(new_n2164), .B(new_n2163), .Y(new_n2165));
  xor_4  g01789(.A(new_n2165), .B(new_n2135), .Y(new_n2166));
  not_8  g01790(.A(new_n2084), .Y(new_n2167));
  nand_5 g01791(.A(new_n2101), .B(new_n2167), .Y(new_n2168));
  nand_5 g01792(.A(pi107), .B(pi006), .Y(new_n2169));
  xor_4  g01793(.A(new_n2169), .B(new_n2168), .Y(new_n2170));
  nor_5  g01794(.A(new_n2099), .B(new_n2096), .Y(new_n2171));
  and_6  g01795(.A(new_n2100), .B(new_n2095), .Y(new_n2172));
  nor_5  g01796(.A(new_n2172), .B(new_n2171), .Y(new_n2173));
  nand_5 g01797(.A(new_n2088), .B(new_n2085), .Y(new_n2174));
  nand_5 g01798(.A(new_n2094), .B(new_n2089), .Y(new_n2175));
  nand_5 g01799(.A(new_n2175), .B(new_n2174), .Y(new_n2176));
  nand_5 g01800(.A(pi154), .B(pi049), .Y(new_n2177));
  nand_5 g01801(.A(pi171), .B(pi095), .Y(new_n2178));
  nand_5 g01802(.A(new_n2178), .B(new_n2177), .Y(new_n2179));
  nand_5 g01803(.A(pi095), .B(pi049), .Y(new_n2180));
  nor_5  g01804(.A(new_n2180), .B(new_n2085), .Y(new_n2181));
  not_8  g01805(.A(new_n2181), .Y(new_n2182));
  nand_5 g01806(.A(new_n2182), .B(new_n2179), .Y(new_n2183));
  nand_5 g01807(.A(new_n2092), .B(new_n2091), .Y(new_n2184));
  nand_5 g01808(.A(new_n2093), .B(new_n2090), .Y(new_n2185));
  nand_5 g01809(.A(new_n2185), .B(new_n2184), .Y(new_n2186));
  nand_5 g01810(.A(pi245), .B(pi089), .Y(new_n2187));
  nand_5 g01811(.A(pi201), .B(pi158), .Y(new_n2188));
  nand_5 g01812(.A(pi254), .B(pi156), .Y(new_n2189));
  nand_5 g01813(.A(new_n2189), .B(new_n2188), .Y(new_n2190));
  nand_5 g01814(.A(pi158), .B(pi156), .Y(new_n2191));
  nor_5  g01815(.A(new_n2191), .B(new_n2091), .Y(new_n2192));
  not_8  g01816(.A(new_n2192), .Y(new_n2193));
  nand_5 g01817(.A(new_n2193), .B(new_n2190), .Y(new_n2194));
  xor_4  g01818(.A(new_n2194), .B(new_n2187), .Y(new_n2195));
  xor_4  g01819(.A(new_n2195), .B(new_n2186), .Y(new_n2196));
  xor_4  g01820(.A(new_n2196), .B(new_n2183), .Y(new_n2197));
  xor_4  g01821(.A(new_n2197), .B(new_n2176), .Y(new_n2198));
  xnor_4 g01822(.A(new_n2198), .B(new_n2173), .Y(new_n2199));
  xnor_4 g01823(.A(new_n2199), .B(new_n2170), .Y(new_n2200));
  xnor_4 g01824(.A(new_n2200), .B(new_n2166), .Y(new_n2201));
  not_8  g01825(.A(new_n2083), .Y(new_n2202));
  nand_5 g01826(.A(new_n2102), .B(new_n2202), .Y(new_n2203));
  or_6   g01827(.A(new_n2103), .B(new_n2036), .Y(new_n2204));
  nand_5 g01828(.A(new_n2204), .B(new_n2203), .Y(new_n2205));
  xnor_4 g01829(.A(new_n2205), .B(new_n2201), .Y(new_n2206));
  nand_5 g01830(.A(new_n2206), .B(new_n2134), .Y(new_n2207));
  nand_5 g01831(.A(new_n2207), .B(new_n2133), .Y(new_n2208));
  nand_5 g01832(.A(new_n2200), .B(new_n2166), .Y(new_n2209));
  or_6   g01833(.A(new_n2205), .B(new_n2201), .Y(new_n2210));
  nand_5 g01834(.A(new_n2210), .B(new_n2209), .Y(new_n2211));
  nand_5 g01835(.A(new_n2169), .B(new_n2168), .Y(new_n2212));
  nand_5 g01836(.A(new_n2199), .B(new_n2170), .Y(new_n2213));
  nand_5 g01837(.A(new_n2213), .B(new_n2212), .Y(new_n2214));
  nor_5  g01838(.A(new_n2198), .B(new_n2173), .Y(new_n2215));
  nand_5 g01839(.A(pi171), .B(pi006), .Y(new_n2216));
  nand_5 g01840(.A(pi209), .B(pi107), .Y(new_n2217));
  xor_4  g01841(.A(new_n2217), .B(new_n2216), .Y(new_n2218));
  xor_4  g01842(.A(new_n2218), .B(new_n2180), .Y(new_n2219));
  nand_5 g01843(.A(new_n2194), .B(new_n2187), .Y(new_n2220));
  nand_5 g01844(.A(new_n2195), .B(new_n2186), .Y(new_n2221));
  nand_5 g01845(.A(new_n2221), .B(new_n2220), .Y(new_n2222));
  xor_4  g01846(.A(new_n2222), .B(new_n2219), .Y(new_n2223));
  nand_5 g01847(.A(pi245), .B(pi154), .Y(new_n2224));
  xor_4  g01848(.A(new_n2224), .B(new_n2192), .Y(new_n2225));
  nand_5 g01849(.A(pi201), .B(pi089), .Y(new_n2226));
  nand_5 g01850(.A(pi254), .B(pi063), .Y(new_n2227));
  xor_4  g01851(.A(new_n2227), .B(new_n2226), .Y(new_n2228));
  xor_4  g01852(.A(new_n2228), .B(new_n2191), .Y(new_n2229));
  xnor_4 g01853(.A(new_n2229), .B(new_n2225), .Y(new_n2230));
  xor_4  g01854(.A(new_n2230), .B(new_n2223), .Y(new_n2231));
  nand_5 g01855(.A(new_n2196), .B(new_n2183), .Y(new_n2232));
  nand_5 g01856(.A(new_n2197), .B(new_n2176), .Y(new_n2233));
  nand_5 g01857(.A(new_n2233), .B(new_n2232), .Y(new_n2234));
  xor_4  g01858(.A(new_n2234), .B(new_n2181), .Y(new_n2235));
  xnor_4 g01859(.A(new_n2235), .B(new_n2231), .Y(new_n2236));
  xor_4  g01860(.A(new_n2236), .B(new_n2215), .Y(new_n2237));
  xor_4  g01861(.A(new_n2237), .B(new_n2214), .Y(new_n2238));
  nand_5 g01862(.A(new_n2162), .B(new_n2138), .Y(new_n2239));
  nor_5  g01863(.A(new_n2161), .B(new_n2141), .Y(new_n2240));
  nand_5 g01864(.A(new_n2240), .B(new_n2146), .Y(new_n2241));
  or_6   g01865(.A(new_n2161), .B(new_n2141), .Y(new_n2242));
  nor_5  g01866(.A(new_n2160), .B(new_n2147), .Y(new_n2243));
  nor_5  g01867(.A(new_n2243), .B(new_n2146), .Y(new_n2244));
  nand_5 g01868(.A(new_n2244), .B(new_n2242), .Y(new_n2245));
  nand_5 g01869(.A(new_n2245), .B(new_n2241), .Y(new_n2246));
  nand_5 g01870(.A(new_n2158), .B(new_n2155), .Y(new_n2247));
  nand_5 g01871(.A(new_n2159), .B(new_n2154), .Y(new_n2248));
  nand_5 g01872(.A(new_n2248), .B(new_n2247), .Y(new_n2249));
  nand_5 g01873(.A(pi148), .B(pi124), .Y(new_n2250));
  nand_5 g01874(.A(pi215), .B(pi163), .Y(new_n2251));
  xor_4  g01875(.A(new_n2251), .B(new_n2145), .Y(new_n2252));
  xor_4  g01876(.A(new_n2252), .B(new_n2250), .Y(new_n2253));
  xor_4  g01877(.A(new_n2253), .B(new_n2249), .Y(new_n2254));
  nand_5 g01878(.A(pi039), .B(pi003), .Y(new_n2255));
  xor_4  g01879(.A(new_n2255), .B(new_n2152), .Y(new_n2256));
  nand_5 g01880(.A(pi116), .B(pi073), .Y(new_n2257));
  nand_5 g01881(.A(pi170), .B(pi115), .Y(new_n2258));
  xor_4  g01882(.A(new_n2258), .B(new_n2257), .Y(new_n2259));
  xor_4  g01883(.A(new_n2259), .B(new_n2151), .Y(new_n2260));
  xnor_4 g01884(.A(new_n2260), .B(new_n2256), .Y(new_n2261));
  xor_4  g01885(.A(new_n2261), .B(new_n2254), .Y(new_n2262));
  not_8  g01886(.A(new_n2262), .Y(new_n2263));
  xor_4  g01887(.A(new_n2263), .B(new_n2246), .Y(new_n2264));
  xor_4  g01888(.A(new_n2264), .B(new_n2239), .Y(new_n2265));
  nor_5  g01889(.A(new_n2164), .B(new_n2163), .Y(new_n2266));
  and_6  g01890(.A(new_n2165), .B(new_n2135), .Y(new_n2267));
  nor_5  g01891(.A(new_n2267), .B(new_n2266), .Y(new_n2268));
  xor_4  g01892(.A(new_n2268), .B(new_n2265), .Y(new_n2269));
  xor_4  g01893(.A(new_n2269), .B(new_n2238), .Y(new_n2270));
  xor_4  g01894(.A(new_n2270), .B(new_n2211), .Y(new_n2271));
  nand_5 g01895(.A(new_n2271), .B(new_n2208), .Y(new_n2272));
  nand_5 g01896(.A(new_n1964), .B(new_n1918), .Y(new_n2273));
  or_6   g01897(.A(new_n1994), .B(new_n1965), .Y(new_n2274));
  nand_5 g01898(.A(new_n2274), .B(new_n2273), .Y(new_n2275));
  or_6   g01899(.A(new_n1993), .B(new_n1968), .Y(new_n2276));
  nand_5 g01900(.A(pi172), .B(pi149), .Y(new_n2277));
  xor_4  g01901(.A(new_n2277), .B(new_n1987), .Y(new_n2278));
  nand_5 g01902(.A(pi200), .B(pi065), .Y(new_n2279));
  nand_5 g01903(.A(pi167), .B(pi120), .Y(new_n2280));
  xor_4  g01904(.A(new_n2280), .B(new_n2279), .Y(new_n2281));
  xor_4  g01905(.A(new_n2281), .B(new_n1986), .Y(new_n2282));
  xor_4  g01906(.A(new_n2282), .B(new_n2278), .Y(new_n2283));
  nand_5 g01907(.A(new_n1989), .B(new_n1982), .Y(new_n2284));
  nand_5 g01908(.A(new_n1990), .B(new_n1981), .Y(new_n2285));
  nand_5 g01909(.A(new_n2285), .B(new_n2284), .Y(new_n2286));
  nand_5 g01910(.A(pi165), .B(pi134), .Y(new_n2287));
  nand_5 g01911(.A(pi197), .B(pi175), .Y(new_n2288));
  xor_4  g01912(.A(new_n2288), .B(new_n2287), .Y(new_n2289));
  xor_4  g01913(.A(new_n2289), .B(new_n1975), .Y(new_n2290));
  xor_4  g01914(.A(new_n2290), .B(new_n2286), .Y(new_n2291));
  not_8  g01915(.A(new_n2291), .Y(new_n2292));
  xor_4  g01916(.A(new_n2292), .B(new_n2283), .Y(new_n2293));
  nand_5 g01917(.A(new_n1991), .B(new_n1978), .Y(new_n2294));
  nand_5 g01918(.A(new_n1992), .B(new_n1971), .Y(new_n2295));
  nand_5 g01919(.A(new_n2295), .B(new_n2294), .Y(new_n2296));
  xor_4  g01920(.A(new_n2296), .B(new_n1977), .Y(new_n2297));
  xor_4  g01921(.A(new_n2297), .B(new_n2293), .Y(new_n2298));
  xor_4  g01922(.A(new_n2298), .B(new_n2276), .Y(new_n2299));
  xor_4  g01923(.A(new_n2299), .B(new_n2275), .Y(new_n2300));
  xor_4  g01924(.A(new_n2271), .B(new_n2208), .Y(new_n2301));
  nand_5 g01925(.A(new_n2301), .B(new_n2300), .Y(new_n2302));
  nand_5 g01926(.A(new_n2302), .B(new_n2272), .Y(new_n2303));
  not_8  g01927(.A(new_n2269), .Y(new_n2304));
  nand_5 g01928(.A(new_n2304), .B(new_n2238), .Y(new_n2305));
  not_8  g01929(.A(new_n2270), .Y(new_n2306));
  nand_5 g01930(.A(new_n2306), .B(new_n2211), .Y(new_n2307));
  nand_5 g01931(.A(new_n2307), .B(new_n2305), .Y(new_n2308));
  xor_4  g01932(.A(new_n2308), .B(new_n2303), .Y(new_n2309));
  nor_5  g01933(.A(new_n2234), .B(new_n2182), .Y(new_n2310));
  nor_5  g01934(.A(new_n2235), .B(new_n2231), .Y(new_n2311));
  nor_5  g01935(.A(new_n2311), .B(new_n2310), .Y(new_n2312));
  nand_5 g01936(.A(pi220), .B(pi103), .Y(new_n2313));
  xor_4  g01937(.A(new_n2313), .B(new_n2312), .Y(new_n2314));
  nand_5 g01938(.A(pi053), .B(pi016), .Y(new_n2315));
  not_8  g01939(.A(new_n2315), .Y(new_n2316));
  nand_5 g01940(.A(pi117), .B(pi067), .Y(new_n2317));
  not_8  g01941(.A(new_n2317), .Y(new_n2318));
  nand_5 g01942(.A(new_n2318), .B(new_n2316), .Y(new_n2319));
  not_8  g01943(.A(new_n2319), .Y(new_n2320));
  nand_5 g01944(.A(pi067), .B(pi016), .Y(new_n2321));
  nand_5 g01945(.A(pi117), .B(pi053), .Y(new_n2322));
  nand_5 g01946(.A(new_n2322), .B(new_n2321), .Y(new_n2323));
  nand_5 g01947(.A(new_n2323), .B(new_n2319), .Y(new_n2324));
  nand_5 g01948(.A(pi234), .B(pi190), .Y(new_n2325));
  nand_5 g01949(.A(pi247), .B(pi092), .Y(new_n2326));
  nand_5 g01950(.A(new_n2326), .B(new_n2325), .Y(new_n2327));
  nand_5 g01951(.A(pi247), .B(pi190), .Y(new_n2328));
  nand_5 g01952(.A(pi234), .B(pi092), .Y(new_n2329));
  nor_5  g01953(.A(new_n2329), .B(new_n2328), .Y(new_n2330));
  not_8  g01954(.A(new_n2330), .Y(new_n2331));
  nand_5 g01955(.A(new_n2331), .B(new_n2327), .Y(new_n2332));
  nand_5 g01956(.A(pi229), .B(pi080), .Y(new_n2333));
  nand_5 g01957(.A(pi229), .B(pi016), .Y(new_n2334));
  nand_5 g01958(.A(pi092), .B(pi080), .Y(new_n2335));
  nand_5 g01959(.A(new_n2335), .B(new_n2334), .Y(new_n2336));
  xor_4  g01960(.A(new_n2335), .B(new_n2334), .Y(new_n2337));
  nand_5 g01961(.A(new_n2337), .B(new_n2328), .Y(new_n2338));
  nand_5 g01962(.A(new_n2338), .B(new_n2336), .Y(new_n2339));
  xor_4  g01963(.A(new_n2339), .B(new_n2333), .Y(new_n2340));
  xor_4  g01964(.A(new_n2340), .B(new_n2332), .Y(new_n2341));
  xor_4  g01965(.A(new_n2341), .B(new_n2324), .Y(new_n2342));
  not_8  g01966(.A(new_n2342), .Y(new_n2343));
  nand_5 g01967(.A(pi092), .B(pi016), .Y(new_n2344));
  nand_5 g01968(.A(pi190), .B(pi080), .Y(new_n2345));
  nand_5 g01969(.A(new_n2345), .B(new_n2344), .Y(new_n2346));
  nand_5 g01970(.A(pi229), .B(pi117), .Y(new_n2347));
  xor_4  g01971(.A(new_n2345), .B(new_n2344), .Y(new_n2348));
  nand_5 g01972(.A(new_n2348), .B(new_n2347), .Y(new_n2349));
  nand_5 g01973(.A(new_n2349), .B(new_n2346), .Y(new_n2350));
  nand_5 g01974(.A(new_n2350), .B(new_n2317), .Y(new_n2351));
  xor_4  g01975(.A(new_n2337), .B(new_n2328), .Y(new_n2352));
  xor_4  g01976(.A(new_n2350), .B(new_n2318), .Y(new_n2353));
  not_8  g01977(.A(new_n2353), .Y(new_n2354));
  nand_5 g01978(.A(new_n2354), .B(new_n2352), .Y(new_n2355));
  nand_5 g01979(.A(new_n2355), .B(new_n2351), .Y(new_n2356));
  nor_5  g01980(.A(new_n2356), .B(new_n2343), .Y(new_n2357));
  and_6  g01981(.A(new_n2357), .B(new_n2320), .Y(new_n2358));
  nor_5  g01982(.A(new_n2341), .B(new_n2324), .Y(new_n2359));
  xor_4  g01983(.A(new_n2357), .B(new_n2320), .Y(new_n2360));
  nor_5  g01984(.A(new_n2360), .B(new_n2359), .Y(new_n2361));
  nand_5 g01985(.A(pi080), .B(pi067), .Y(new_n2362));
  xor_4  g01986(.A(new_n2362), .B(new_n2330), .Y(new_n2363));
  nand_5 g01987(.A(pi214), .B(pi190), .Y(new_n2364));
  nand_5 g01988(.A(pi247), .B(pi229), .Y(new_n2365));
  xor_4  g01989(.A(new_n2365), .B(new_n2364), .Y(new_n2366));
  xor_4  g01990(.A(new_n2366), .B(new_n2329), .Y(new_n2367));
  xor_4  g01991(.A(new_n2367), .B(new_n2363), .Y(new_n2368));
  nand_5 g01992(.A(new_n2339), .B(new_n2333), .Y(new_n2369));
  nand_5 g01993(.A(new_n2340), .B(new_n2332), .Y(new_n2370));
  nand_5 g01994(.A(new_n2370), .B(new_n2369), .Y(new_n2371));
  nand_5 g01995(.A(pi103), .B(pi030), .Y(new_n2372));
  nand_5 g01996(.A(pi185), .B(pi117), .Y(new_n2373));
  xor_4  g01997(.A(new_n2373), .B(new_n2372), .Y(new_n2374));
  xor_4  g01998(.A(new_n2374), .B(new_n2316), .Y(new_n2375));
  xor_4  g01999(.A(new_n2375), .B(new_n2371), .Y(new_n2376));
  xor_4  g02000(.A(new_n2376), .B(new_n2368), .Y(new_n2377));
  nor_5  g02001(.A(new_n2377), .B(new_n2361), .Y(new_n2378));
  nor_5  g02002(.A(new_n2378), .B(new_n2358), .Y(new_n2379));
  nand_5 g02003(.A(new_n2280), .B(new_n2279), .Y(new_n2380));
  nand_5 g02004(.A(new_n2281), .B(new_n1986), .Y(new_n2381));
  nand_5 g02005(.A(new_n2381), .B(new_n2380), .Y(new_n2382));
  xor_4  g02006(.A(new_n2382), .B(new_n2379), .Y(new_n2383));
  nand_5 g02007(.A(pi197), .B(pi134), .Y(new_n2384));
  nand_5 g02008(.A(new_n2365), .B(new_n2364), .Y(new_n2385));
  nand_5 g02009(.A(new_n2366), .B(new_n2329), .Y(new_n2386));
  nand_5 g02010(.A(new_n2386), .B(new_n2385), .Y(new_n2387));
  xor_4  g02011(.A(new_n2387), .B(new_n2384), .Y(new_n2388));
  not_8  g02012(.A(new_n2375), .Y(new_n2389));
  nand_5 g02013(.A(new_n2389), .B(new_n2371), .Y(new_n2390));
  or_6   g02014(.A(new_n2376), .B(new_n2368), .Y(new_n2391));
  nand_5 g02015(.A(new_n2391), .B(new_n2390), .Y(new_n2392));
  nand_5 g02016(.A(pi175), .B(pi078), .Y(new_n2393));
  xor_4  g02017(.A(new_n2393), .B(new_n2392), .Y(new_n2394));
  nand_5 g02018(.A(new_n2290), .B(new_n2286), .Y(new_n2395));
  or_6   g02019(.A(new_n2292), .B(new_n2283), .Y(new_n2396));
  nand_5 g02020(.A(new_n2396), .B(new_n2395), .Y(new_n2397));
  nand_5 g02021(.A(pi163), .B(pi022), .Y(new_n2398));
  xor_4  g02022(.A(new_n2398), .B(new_n2397), .Y(new_n2399));
  xor_4  g02023(.A(new_n2399), .B(new_n2394), .Y(new_n2400));
  xor_4  g02024(.A(new_n2400), .B(new_n2388), .Y(new_n2401));
  xor_4  g02025(.A(new_n2401), .B(new_n2383), .Y(new_n2402));
  xor_4  g02026(.A(new_n2402), .B(new_n2314), .Y(new_n2403));
  nand_5 g02027(.A(pi049), .B(pi006), .Y(new_n2404));
  nor_5  g02028(.A(new_n2264), .B(new_n2239), .Y(new_n2405));
  not_8  g02029(.A(new_n2265), .Y(new_n2406));
  nor_5  g02030(.A(new_n2268), .B(new_n2406), .Y(new_n2407));
  nor_5  g02031(.A(new_n2407), .B(new_n2405), .Y(new_n2408));
  nand_5 g02032(.A(new_n2253), .B(new_n2249), .Y(new_n2409));
  nand_5 g02033(.A(new_n2261), .B(new_n2254), .Y(new_n2410));
  nand_5 g02034(.A(new_n2410), .B(new_n2409), .Y(new_n2411));
  xor_4  g02035(.A(new_n2411), .B(new_n2408), .Y(new_n2412));
  nand_5 g02036(.A(new_n2222), .B(new_n2219), .Y(new_n2413));
  nand_5 g02037(.A(new_n2230), .B(new_n2223), .Y(new_n2414));
  nand_5 g02038(.A(new_n2414), .B(new_n2413), .Y(new_n2415));
  xor_4  g02039(.A(new_n2415), .B(new_n2412), .Y(new_n2416));
  nand_5 g02040(.A(new_n2258), .B(new_n2257), .Y(new_n2417));
  nand_5 g02041(.A(new_n2259), .B(new_n2151), .Y(new_n2418));
  nand_5 g02042(.A(new_n2418), .B(new_n2417), .Y(new_n2419));
  nand_5 g02043(.A(pi245), .B(pi095), .Y(new_n2420));
  nor_5  g02044(.A(new_n2224), .B(new_n2193), .Y(new_n2421));
  nor_5  g02045(.A(new_n2229), .B(new_n2225), .Y(new_n2422));
  nor_5  g02046(.A(new_n2422), .B(new_n2421), .Y(new_n2423));
  xor_4  g02047(.A(new_n2423), .B(new_n2420), .Y(new_n2424));
  xor_4  g02048(.A(new_n2424), .B(new_n2419), .Y(new_n2425));
  xor_4  g02049(.A(new_n2425), .B(new_n2416), .Y(new_n2426));
  xor_4  g02050(.A(new_n2426), .B(new_n2404), .Y(new_n2427));
  xor_4  g02051(.A(new_n2427), .B(new_n2403), .Y(new_n2428));
  xor_4  g02052(.A(new_n2428), .B(new_n2309), .Y(new_n2429));
  or_6   g02053(.A(new_n2263), .B(new_n2246), .Y(new_n2430));
  nand_5 g02054(.A(new_n2430), .B(new_n2245), .Y(new_n2431));
  nand_5 g02055(.A(pi198), .B(pi149), .Y(new_n2432));
  not_8  g02056(.A(new_n2215), .Y(new_n2433));
  nand_5 g02057(.A(new_n2236), .B(new_n2433), .Y(new_n2434));
  not_8  g02058(.A(new_n2237), .Y(new_n2435));
  nand_5 g02059(.A(new_n2435), .B(new_n2214), .Y(new_n2436));
  nand_5 g02060(.A(new_n2436), .B(new_n2434), .Y(new_n2437));
  nand_5 g02061(.A(new_n2217), .B(new_n2216), .Y(new_n2438));
  nand_5 g02062(.A(new_n2218), .B(new_n2180), .Y(new_n2439));
  nand_5 g02063(.A(new_n2439), .B(new_n2438), .Y(new_n2440));
  xor_4  g02064(.A(new_n2440), .B(new_n2437), .Y(new_n2441));
  nand_5 g02065(.A(new_n2288), .B(new_n2287), .Y(new_n2442));
  nand_5 g02066(.A(new_n2289), .B(new_n1975), .Y(new_n2443));
  nand_5 g02067(.A(new_n2443), .B(new_n2442), .Y(new_n2444));
  nor_5  g02068(.A(new_n2277), .B(new_n1988), .Y(new_n2445));
  nor_5  g02069(.A(new_n2282), .B(new_n2278), .Y(new_n2446));
  nor_5  g02070(.A(new_n2446), .B(new_n2445), .Y(new_n2447));
  xor_4  g02071(.A(new_n2447), .B(new_n2444), .Y(new_n2448));
  xor_4  g02072(.A(new_n2448), .B(new_n2441), .Y(new_n2449));
  xor_4  g02073(.A(new_n2449), .B(new_n2432), .Y(new_n2450));
  nor_5  g02074(.A(new_n2255), .B(new_n2153), .Y(new_n2451));
  nor_5  g02075(.A(new_n2260), .B(new_n2256), .Y(new_n2452));
  nor_5  g02076(.A(new_n2452), .B(new_n2451), .Y(new_n2453));
  nand_5 g02077(.A(pi228), .B(pi124), .Y(new_n2454));
  xor_4  g02078(.A(new_n2454), .B(new_n2453), .Y(new_n2455));
  xor_4  g02079(.A(new_n2455), .B(new_n2450), .Y(new_n2456));
  nand_5 g02080(.A(pi202), .B(pi190), .Y(new_n2457));
  nand_5 g02081(.A(new_n2227), .B(new_n2226), .Y(new_n2458));
  nand_5 g02082(.A(new_n2228), .B(new_n2191), .Y(new_n2459));
  nand_5 g02083(.A(new_n2459), .B(new_n2458), .Y(new_n2460));
  xor_4  g02084(.A(new_n2460), .B(new_n2457), .Y(new_n2461));
  nand_5 g02085(.A(pi156), .B(pi089), .Y(new_n2462));
  nand_5 g02086(.A(new_n2251), .B(new_n2145), .Y(new_n2463));
  nand_5 g02087(.A(new_n2252), .B(new_n2250), .Y(new_n2464));
  nand_5 g02088(.A(new_n2464), .B(new_n2463), .Y(new_n2465));
  xor_4  g02089(.A(new_n2465), .B(new_n2462), .Y(new_n2466));
  xor_4  g02090(.A(new_n2377), .B(new_n2361), .Y(new_n2467));
  nand_5 g02091(.A(pi103), .B(pi053), .Y(new_n2468));
  xor_4  g02092(.A(new_n2353), .B(new_n2352), .Y(new_n2469));
  not_8  g02093(.A(new_n2469), .Y(new_n2470));
  nor_5  g02094(.A(new_n2470), .B(new_n2468), .Y(new_n2471));
  nand_5 g02095(.A(pi103), .B(pi067), .Y(new_n2472));
  nand_5 g02096(.A(pi229), .B(pi103), .Y(new_n2473));
  nand_5 g02097(.A(pi117), .B(pi092), .Y(new_n2474));
  nand_5 g02098(.A(new_n2474), .B(new_n2473), .Y(new_n2475));
  nand_5 g02099(.A(pi190), .B(pi016), .Y(new_n2476));
  xor_4  g02100(.A(new_n2474), .B(new_n2473), .Y(new_n2477));
  nand_5 g02101(.A(new_n2477), .B(new_n2476), .Y(new_n2478));
  nand_5 g02102(.A(new_n2478), .B(new_n2475), .Y(new_n2479));
  nor_5  g02103(.A(new_n2479), .B(new_n2472), .Y(new_n2480));
  xor_4  g02104(.A(new_n2348), .B(new_n2347), .Y(new_n2481));
  xor_4  g02105(.A(new_n2479), .B(new_n2472), .Y(new_n2482));
  not_8  g02106(.A(new_n2482), .Y(new_n2483));
  nor_5  g02107(.A(new_n2483), .B(new_n2481), .Y(new_n2484));
  nor_5  g02108(.A(new_n2484), .B(new_n2480), .Y(new_n2485));
  xor_4  g02109(.A(new_n2469), .B(new_n2468), .Y(new_n2486));
  or_6   g02110(.A(new_n2486), .B(new_n2485), .Y(new_n2487));
  not_8  g02111(.A(new_n2487), .Y(new_n2488));
  nor_5  g02112(.A(new_n2488), .B(new_n2471), .Y(new_n2489));
  xor_4  g02113(.A(new_n2356), .B(new_n2342), .Y(new_n2490));
  nor_5  g02114(.A(new_n2490), .B(new_n2489), .Y(new_n2491));
  or_6   g02115(.A(new_n2491), .B(new_n2467), .Y(new_n2492));
  xor_4  g02116(.A(new_n2491), .B(new_n2467), .Y(new_n2493));
  nand_5 g02117(.A(pi185), .B(pi103), .Y(new_n2494));
  xor_4  g02118(.A(new_n2486), .B(new_n2485), .Y(new_n2495));
  xor_4  g02119(.A(new_n2477), .B(new_n2476), .Y(new_n2496));
  nand_5 g02120(.A(pi190), .B(pi103), .Y(new_n2497));
  nor_5  g02121(.A(new_n2497), .B(new_n2474), .Y(new_n2498));
  not_8  g02122(.A(new_n2498), .Y(new_n2499));
  nor_5  g02123(.A(new_n2499), .B(new_n2496), .Y(new_n2500));
  not_8  g02124(.A(new_n2500), .Y(new_n2501));
  xor_4  g02125(.A(new_n2482), .B(new_n2481), .Y(new_n2502));
  nor_5  g02126(.A(new_n2502), .B(new_n2501), .Y(new_n2503));
  nand_5 g02127(.A(new_n2503), .B(new_n2495), .Y(new_n2504));
  nand_5 g02128(.A(new_n2504), .B(new_n2494), .Y(new_n2505));
  xor_4  g02129(.A(new_n2504), .B(new_n2494), .Y(new_n2506));
  xnor_4 g02130(.A(new_n2490), .B(new_n2489), .Y(new_n2507));
  nand_5 g02131(.A(new_n2507), .B(new_n2506), .Y(new_n2508));
  nand_5 g02132(.A(new_n2508), .B(new_n2505), .Y(new_n2509));
  nand_5 g02133(.A(new_n2509), .B(new_n2493), .Y(new_n2510));
  nand_5 g02134(.A(new_n2510), .B(new_n2492), .Y(new_n2511));
  nand_5 g02135(.A(pi234), .B(pi229), .Y(new_n2512));
  xor_4  g02136(.A(new_n2512), .B(new_n2511), .Y(new_n2513));
  nand_5 g02137(.A(pi158), .B(pi063), .Y(new_n2514));
  nand_5 g02138(.A(pi254), .B(pi083), .Y(new_n2515));
  xor_4  g02139(.A(new_n2515), .B(new_n2514), .Y(new_n2516));
  nand_5 g02140(.A(pi130), .B(pi039), .Y(new_n2517));
  xor_4  g02141(.A(new_n2517), .B(new_n2516), .Y(new_n2518));
  xor_4  g02142(.A(new_n2518), .B(new_n2513), .Y(new_n2519));
  xor_4  g02143(.A(new_n2519), .B(new_n2466), .Y(new_n2520));
  xor_4  g02144(.A(new_n2520), .B(new_n2461), .Y(new_n2521));
  xor_4  g02145(.A(new_n2521), .B(new_n2456), .Y(new_n2522));
  nand_5 g02146(.A(pi209), .B(pi171), .Y(new_n2523));
  nand_5 g02147(.A(pi153), .B(pi107), .Y(new_n2524));
  nand_5 g02148(.A(pi215), .B(pi148), .Y(new_n2525));
  nand_5 g02149(.A(pi201), .B(pi154), .Y(new_n2526));
  xor_4  g02150(.A(new_n2526), .B(new_n2525), .Y(new_n2527));
  nand_5 g02151(.A(pi116), .B(pi003), .Y(new_n2528));
  xor_4  g02152(.A(new_n2528), .B(new_n2527), .Y(new_n2529));
  xor_4  g02153(.A(new_n2529), .B(new_n2524), .Y(new_n2530));
  xor_4  g02154(.A(new_n2530), .B(new_n2523), .Y(new_n2531));
  xor_4  g02155(.A(new_n2531), .B(new_n2522), .Y(new_n2532));
  xor_4  g02156(.A(new_n2532), .B(new_n2431), .Y(new_n2533));
  xor_4  g02157(.A(new_n2533), .B(new_n2429), .Y(new_n2534));
  nand_5 g02158(.A(pi117), .B(pi030), .Y(new_n2535));
  nand_5 g02159(.A(pi240), .B(pi165), .Y(new_n2536));
  xor_4  g02160(.A(new_n2536), .B(new_n2535), .Y(new_n2537));
  nand_5 g02161(.A(pi185), .B(pi016), .Y(new_n2538));
  xor_4  g02162(.A(new_n2538), .B(new_n2537), .Y(new_n2539));
  xor_4  g02163(.A(new_n2539), .B(new_n2534), .Y(new_n2540));
  nand_5 g02164(.A(pi172), .B(pi167), .Y(new_n2541));
  nand_5 g02165(.A(new_n2298), .B(new_n2276), .Y(new_n2542));
  nand_5 g02166(.A(new_n2299), .B(new_n2275), .Y(new_n2543));
  nand_5 g02167(.A(new_n2543), .B(new_n2542), .Y(new_n2544));
  xor_4  g02168(.A(new_n2544), .B(new_n2541), .Y(new_n2545));
  xnor_4 g02169(.A(new_n2509), .B(new_n2493), .Y(new_n2546));
  xnor_4 g02170(.A(new_n2301), .B(new_n2300), .Y(new_n2547));
  nand_5 g02171(.A(new_n2547), .B(new_n2546), .Y(new_n2548));
  xor_4  g02172(.A(new_n2547), .B(new_n2546), .Y(new_n2549));
  xor_4  g02173(.A(new_n2507), .B(new_n2506), .Y(new_n2550));
  not_8  g02174(.A(new_n2550), .Y(new_n2551));
  xnor_4 g02175(.A(new_n2206), .B(new_n2134), .Y(new_n2552));
  nand_5 g02176(.A(new_n2552), .B(new_n2551), .Y(new_n2553));
  xor_4  g02177(.A(new_n2552), .B(new_n2551), .Y(new_n2554));
  xnor_4 g02178(.A(new_n2128), .B(new_n2110), .Y(new_n2555));
  xor_4  g02179(.A(new_n2502), .B(new_n2500), .Y(new_n2556));
  not_8  g02180(.A(new_n2556), .Y(new_n2557));
  nor_5  g02181(.A(new_n2557), .B(new_n2555), .Y(new_n2558));
  xor_4  g02182(.A(new_n2119), .B(new_n1956), .Y(new_n2559));
  or_6   g02183(.A(new_n2559), .B(new_n2497), .Y(new_n2560));
  nand_5 g02184(.A(pi103), .B(pi092), .Y(new_n2561));
  nand_5 g02185(.A(pi190), .B(pi117), .Y(new_n2562));
  nand_5 g02186(.A(new_n2562), .B(new_n2561), .Y(new_n2563));
  nand_5 g02187(.A(new_n2563), .B(new_n2499), .Y(new_n2564));
  nor_5  g02188(.A(new_n2564), .B(new_n2560), .Y(new_n2565));
  xor_4  g02189(.A(new_n2564), .B(new_n2560), .Y(new_n2566));
  xor_4  g02190(.A(new_n2123), .B(new_n2122), .Y(new_n2567));
  not_8  g02191(.A(new_n2567), .Y(new_n2568));
  nand_5 g02192(.A(new_n2568), .B(new_n2566), .Y(new_n2569));
  not_8  g02193(.A(new_n2569), .Y(new_n2570));
  nor_5  g02194(.A(new_n2570), .B(new_n2565), .Y(new_n2571));
  xor_4  g02195(.A(new_n2498), .B(new_n2496), .Y(new_n2572));
  nor_5  g02196(.A(new_n2572), .B(new_n2571), .Y(new_n2573));
  not_8  g02197(.A(new_n2573), .Y(new_n2574));
  xor_4  g02198(.A(new_n2572), .B(new_n2571), .Y(new_n2575));
  xor_4  g02199(.A(new_n2126), .B(new_n2125), .Y(new_n2576));
  nand_5 g02200(.A(new_n2576), .B(new_n2575), .Y(new_n2577));
  nand_5 g02201(.A(new_n2577), .B(new_n2574), .Y(new_n2578));
  xor_4  g02202(.A(new_n2556), .B(new_n2555), .Y(new_n2579));
  nor_5  g02203(.A(new_n2579), .B(new_n2578), .Y(new_n2580));
  nor_5  g02204(.A(new_n2580), .B(new_n2558), .Y(new_n2581));
  xnor_4 g02205(.A(new_n2130), .B(new_n2106), .Y(new_n2582));
  xnor_4 g02206(.A(new_n2503), .B(new_n2495), .Y(new_n2583));
  nor_5  g02207(.A(new_n2583), .B(new_n2582), .Y(new_n2584));
  nor_5  g02208(.A(new_n2584), .B(new_n2581), .Y(new_n2585));
  and_6  g02209(.A(new_n2583), .B(new_n2582), .Y(new_n2586));
  nor_5  g02210(.A(new_n2586), .B(new_n2585), .Y(new_n2587));
  nand_5 g02211(.A(new_n2587), .B(new_n2554), .Y(new_n2588));
  nand_5 g02212(.A(new_n2588), .B(new_n2553), .Y(new_n2589));
  nand_5 g02213(.A(new_n2589), .B(new_n2549), .Y(new_n2590));
  nand_5 g02214(.A(new_n2590), .B(new_n2548), .Y(new_n2591));
  nand_5 g02215(.A(pi181), .B(pi120), .Y(new_n2592));
  xor_4  g02216(.A(new_n2592), .B(new_n2591), .Y(new_n2593));
  nand_5 g02217(.A(pi214), .B(pi092), .Y(new_n2594));
  nor_5  g02218(.A(new_n2296), .B(new_n1977), .Y(new_n2595));
  not_8  g02219(.A(new_n2297), .Y(new_n2596));
  nor_5  g02220(.A(new_n2596), .B(new_n2293), .Y(new_n2597));
  nor_5  g02221(.A(new_n2597), .B(new_n2595), .Y(new_n2598));
  xor_4  g02222(.A(new_n2598), .B(new_n2594), .Y(new_n2599));
  nand_5 g02223(.A(pi247), .B(pi067), .Y(new_n2600));
  xor_4  g02224(.A(new_n2600), .B(new_n2599), .Y(new_n2601));
  xor_4  g02225(.A(new_n2601), .B(new_n2593), .Y(new_n2602));
  xor_4  g02226(.A(new_n2602), .B(new_n2545), .Y(new_n2603));
  nand_5 g02227(.A(pi115), .B(pi004), .Y(new_n2604));
  nand_5 g02228(.A(new_n2373), .B(new_n2372), .Y(new_n2605));
  nand_5 g02229(.A(new_n2374), .B(new_n2315), .Y(new_n2606));
  nand_5 g02230(.A(new_n2606), .B(new_n2605), .Y(new_n2607));
  nand_5 g02231(.A(pi200), .B(pi062), .Y(new_n2608));
  xnor_4 g02232(.A(new_n2608), .B(new_n2607), .Y(new_n2609));
  xor_4  g02233(.A(new_n2609), .B(new_n2604), .Y(new_n2610));
  nand_5 g02234(.A(pi203), .B(pi065), .Y(new_n2611));
  nand_5 g02235(.A(pi170), .B(pi000), .Y(new_n2612));
  nand_5 g02236(.A(pi073), .B(pi070), .Y(new_n2613));
  xor_4  g02237(.A(new_n2613), .B(new_n2612), .Y(new_n2614));
  xor_4  g02238(.A(new_n2614), .B(new_n2611), .Y(new_n2615));
  xor_4  g02239(.A(new_n2615), .B(new_n2610), .Y(new_n2616));
  nor_5  g02240(.A(new_n2362), .B(new_n2331), .Y(new_n2617));
  nor_5  g02241(.A(new_n2367), .B(new_n2363), .Y(new_n2618));
  nor_5  g02242(.A(new_n2618), .B(new_n2617), .Y(new_n2619));
  nand_5 g02243(.A(pi080), .B(pi053), .Y(new_n2620));
  xor_4  g02244(.A(new_n2620), .B(new_n2619), .Y(new_n2621));
  xor_4  g02245(.A(new_n2621), .B(new_n2616), .Y(new_n2622));
  xor_4  g02246(.A(new_n2622), .B(new_n2603), .Y(new_n2623));
  xor_4  g02247(.A(new_n2623), .B(new_n2540), .Y(po006));
  nand_5 g02248(.A(pi065), .B(pi041), .Y(new_n2625));
  nand_5 g02249(.A(pi182), .B(pi062), .Y(new_n2626));
  nand_5 g02250(.A(pi138), .B(pi120), .Y(new_n2627));
  xor_4  g02251(.A(new_n2627), .B(new_n2626), .Y(new_n2628));
  xor_4  g02252(.A(new_n2628), .B(new_n2625), .Y(new_n2629));
  nand_5 g02253(.A(pi138), .B(pi065), .Y(new_n2630));
  or_6   g02254(.A(new_n2630), .B(new_n2626), .Y(new_n2631));
  or_6   g02255(.A(new_n2631), .B(new_n2629), .Y(new_n2632));
  nand_5 g02256(.A(pi182), .B(pi120), .Y(new_n2633));
  nand_5 g02257(.A(pi062), .B(pi041), .Y(new_n2634));
  nand_5 g02258(.A(pi216), .B(pi065), .Y(new_n2635));
  xor_4  g02259(.A(new_n2635), .B(new_n2634), .Y(new_n2636));
  xor_4  g02260(.A(new_n2636), .B(new_n2633), .Y(new_n2637));
  nand_5 g02261(.A(pi172), .B(pi138), .Y(new_n2638));
  nand_5 g02262(.A(new_n2627), .B(new_n2626), .Y(new_n2639));
  nand_5 g02263(.A(new_n2628), .B(new_n2625), .Y(new_n2640));
  nand_5 g02264(.A(new_n2640), .B(new_n2639), .Y(new_n2641));
  xor_4  g02265(.A(new_n2641), .B(new_n2638), .Y(new_n2642));
  xor_4  g02266(.A(new_n2642), .B(new_n2637), .Y(new_n2643));
  xor_4  g02267(.A(new_n2643), .B(new_n2632), .Y(new_n2644));
  nand_5 g02268(.A(pi071), .B(pi004), .Y(new_n2645));
  nand_5 g02269(.A(pi170), .B(pi142), .Y(new_n2646));
  not_8  g02270(.A(new_n2646), .Y(new_n2647));
  nor_5  g02271(.A(new_n2647), .B(new_n2645), .Y(new_n2648));
  nand_5 g02272(.A(pi170), .B(pi169), .Y(new_n2649));
  nand_5 g02273(.A(pi142), .B(pi073), .Y(new_n2650));
  or_6   g02274(.A(new_n2650), .B(new_n2649), .Y(new_n2651));
  nand_5 g02275(.A(new_n2650), .B(new_n2649), .Y(new_n2652));
  and_6  g02276(.A(new_n2652), .B(new_n2651), .Y(new_n2653));
  or_6   g02277(.A(new_n2653), .B(new_n2648), .Y(new_n2654));
  nand_5 g02278(.A(new_n2652), .B(new_n2648), .Y(new_n2655));
  nand_5 g02279(.A(new_n2655), .B(new_n2654), .Y(new_n2656));
  nand_5 g02280(.A(pi219), .B(pi158), .Y(new_n2657));
  nand_5 g02281(.A(pi254), .B(pi087), .Y(new_n2658));
  not_8  g02282(.A(new_n2658), .Y(new_n2659));
  nor_5  g02283(.A(new_n2659), .B(new_n2657), .Y(new_n2660));
  nand_5 g02284(.A(pi254), .B(pi102), .Y(new_n2661));
  nand_5 g02285(.A(pi089), .B(pi087), .Y(new_n2662));
  or_6   g02286(.A(new_n2662), .B(new_n2661), .Y(new_n2663));
  nand_5 g02287(.A(new_n2662), .B(new_n2661), .Y(new_n2664));
  and_6  g02288(.A(new_n2664), .B(new_n2663), .Y(new_n2665));
  or_6   g02289(.A(new_n2665), .B(new_n2660), .Y(new_n2666));
  nand_5 g02290(.A(new_n2660), .B(new_n2664), .Y(new_n2667));
  nand_5 g02291(.A(new_n2667), .B(new_n2666), .Y(new_n2668));
  nand_5 g02292(.A(new_n2668), .B(new_n2656), .Y(new_n2669));
  xnor_4 g02293(.A(new_n2668), .B(new_n2656), .Y(new_n2670));
  nor_5  g02294(.A(new_n2658), .B(new_n2646), .Y(new_n2671));
  nand_5 g02295(.A(pi158), .B(pi087), .Y(new_n2672));
  nand_5 g02296(.A(pi254), .B(pi219), .Y(new_n2673));
  xor_4  g02297(.A(new_n2673), .B(new_n2672), .Y(new_n2674));
  nand_5 g02298(.A(new_n2674), .B(new_n2671), .Y(new_n2675));
  nand_5 g02299(.A(pi142), .B(pi004), .Y(new_n2676));
  nand_5 g02300(.A(pi170), .B(pi071), .Y(new_n2677));
  xor_4  g02301(.A(new_n2677), .B(new_n2676), .Y(new_n2678));
  xor_4  g02302(.A(new_n2674), .B(new_n2671), .Y(new_n2679));
  nand_5 g02303(.A(new_n2679), .B(new_n2678), .Y(new_n2680));
  nand_5 g02304(.A(new_n2680), .B(new_n2675), .Y(new_n2681));
  or_6   g02305(.A(new_n2681), .B(new_n2670), .Y(new_n2682));
  nand_5 g02306(.A(new_n2682), .B(new_n2669), .Y(new_n2683));
  or_6   g02307(.A(new_n2666), .B(new_n2657), .Y(new_n2684));
  nand_5 g02308(.A(pi254), .B(pi001), .Y(new_n2685));
  nand_5 g02309(.A(pi158), .B(pi102), .Y(new_n2686));
  nand_5 g02310(.A(pi219), .B(pi089), .Y(new_n2687));
  xor_4  g02311(.A(new_n2687), .B(new_n2686), .Y(new_n2688));
  xor_4  g02312(.A(new_n2688), .B(new_n2685), .Y(new_n2689));
  nand_5 g02313(.A(new_n2657), .B(new_n2663), .Y(new_n2690));
  nand_5 g02314(.A(new_n2690), .B(new_n2664), .Y(new_n2691));
  nand_5 g02315(.A(pi154), .B(pi087), .Y(new_n2692));
  xor_4  g02316(.A(new_n2692), .B(new_n2691), .Y(new_n2693));
  xor_4  g02317(.A(new_n2693), .B(new_n2689), .Y(new_n2694));
  xnor_4 g02318(.A(new_n2694), .B(new_n2684), .Y(new_n2695));
  xor_4  g02319(.A(new_n2695), .B(new_n2683), .Y(new_n2696));
  nor_5  g02320(.A(new_n2654), .B(new_n2645), .Y(new_n2697));
  nand_5 g02321(.A(pi170), .B(pi123), .Y(new_n2698));
  nand_5 g02322(.A(pi169), .B(pi004), .Y(new_n2699));
  nand_5 g02323(.A(pi073), .B(pi071), .Y(new_n2700));
  xor_4  g02324(.A(new_n2700), .B(new_n2699), .Y(new_n2701));
  xor_4  g02325(.A(new_n2701), .B(new_n2698), .Y(new_n2702));
  nand_5 g02326(.A(new_n2645), .B(new_n2651), .Y(new_n2703));
  nand_5 g02327(.A(new_n2703), .B(new_n2652), .Y(new_n2704));
  nand_5 g02328(.A(pi142), .B(pi003), .Y(new_n2705));
  xor_4  g02329(.A(new_n2705), .B(new_n2704), .Y(new_n2706));
  xor_4  g02330(.A(new_n2706), .B(new_n2702), .Y(new_n2707));
  xor_4  g02331(.A(new_n2707), .B(new_n2697), .Y(new_n2708));
  xnor_4 g02332(.A(new_n2708), .B(new_n2696), .Y(new_n2709));
  or_6   g02333(.A(new_n2709), .B(new_n2644), .Y(new_n2710));
  xor_4  g02334(.A(new_n2709), .B(new_n2644), .Y(new_n2711));
  xor_4  g02335(.A(new_n2659), .B(new_n2646), .Y(new_n2712));
  or_6   g02336(.A(new_n2712), .B(new_n2630), .Y(new_n2713));
  nand_5 g02337(.A(pi138), .B(pi062), .Y(new_n2714));
  nand_5 g02338(.A(pi182), .B(pi065), .Y(new_n2715));
  nand_5 g02339(.A(new_n2715), .B(new_n2714), .Y(new_n2716));
  nand_5 g02340(.A(new_n2716), .B(new_n2631), .Y(new_n2717));
  nand_5 g02341(.A(new_n2717), .B(new_n2713), .Y(new_n2718));
  xnor_4 g02342(.A(new_n2717), .B(new_n2713), .Y(new_n2719));
  xor_4  g02343(.A(new_n2679), .B(new_n2678), .Y(new_n2720));
  or_6   g02344(.A(new_n2720), .B(new_n2719), .Y(new_n2721));
  nand_5 g02345(.A(new_n2721), .B(new_n2718), .Y(new_n2722));
  xnor_4 g02346(.A(new_n2631), .B(new_n2629), .Y(new_n2723));
  nor_5  g02347(.A(new_n2723), .B(new_n2722), .Y(new_n2724));
  xor_4  g02348(.A(new_n2681), .B(new_n2670), .Y(new_n2725));
  xnor_4 g02349(.A(new_n2723), .B(new_n2722), .Y(new_n2726));
  nor_5  g02350(.A(new_n2726), .B(new_n2725), .Y(new_n2727));
  nor_5  g02351(.A(new_n2727), .B(new_n2724), .Y(new_n2728));
  nand_5 g02352(.A(new_n2728), .B(new_n2711), .Y(new_n2729));
  nand_5 g02353(.A(new_n2729), .B(new_n2710), .Y(new_n2730));
  nor_5  g02354(.A(new_n2643), .B(new_n2632), .Y(new_n2731));
  nand_5 g02355(.A(pi198), .B(pi138), .Y(new_n2732));
  nand_5 g02356(.A(pi216), .B(pi062), .Y(new_n2733));
  nand_5 g02357(.A(pi076), .B(pi065), .Y(new_n2734));
  nand_5 g02358(.A(pi120), .B(pi041), .Y(new_n2735));
  xor_4  g02359(.A(new_n2735), .B(new_n2734), .Y(new_n2736));
  xor_4  g02360(.A(new_n2736), .B(new_n2733), .Y(new_n2737));
  nand_5 g02361(.A(pi182), .B(pi172), .Y(new_n2738));
  nand_5 g02362(.A(new_n2635), .B(new_n2634), .Y(new_n2739));
  nand_5 g02363(.A(new_n2636), .B(new_n2633), .Y(new_n2740));
  nand_5 g02364(.A(new_n2740), .B(new_n2739), .Y(new_n2741));
  xor_4  g02365(.A(new_n2741), .B(new_n2738), .Y(new_n2742));
  xor_4  g02366(.A(new_n2742), .B(new_n2737), .Y(new_n2743));
  xor_4  g02367(.A(new_n2743), .B(new_n2732), .Y(new_n2744));
  nor_5  g02368(.A(new_n2641), .B(new_n2638), .Y(new_n2745));
  not_8  g02369(.A(new_n2642), .Y(new_n2746));
  nor_5  g02370(.A(new_n2746), .B(new_n2637), .Y(new_n2747));
  nor_5  g02371(.A(new_n2747), .B(new_n2745), .Y(new_n2748));
  xor_4  g02372(.A(new_n2748), .B(new_n2744), .Y(new_n2749));
  xor_4  g02373(.A(new_n2749), .B(new_n2731), .Y(new_n2750));
  nand_5 g02374(.A(new_n2750), .B(new_n2730), .Y(new_n2751));
  nand_5 g02375(.A(new_n2695), .B(new_n2683), .Y(new_n2752));
  nand_5 g02376(.A(new_n2708), .B(new_n2696), .Y(new_n2753));
  nand_5 g02377(.A(new_n2753), .B(new_n2752), .Y(new_n2754));
  nor_5  g02378(.A(new_n2694), .B(new_n2684), .Y(new_n2755));
  nor_5  g02379(.A(new_n2692), .B(new_n2691), .Y(new_n2756));
  not_8  g02380(.A(new_n2693), .Y(new_n2757));
  nor_5  g02381(.A(new_n2757), .B(new_n2689), .Y(new_n2758));
  or_6   g02382(.A(new_n2758), .B(new_n2756), .Y(new_n2759));
  nand_5 g02383(.A(pi095), .B(pi087), .Y(new_n2760));
  nand_5 g02384(.A(pi102), .B(pi089), .Y(new_n2761));
  nand_5 g02385(.A(pi254), .B(pi122), .Y(new_n2762));
  nand_5 g02386(.A(pi158), .B(pi001), .Y(new_n2763));
  xor_4  g02387(.A(new_n2763), .B(new_n2762), .Y(new_n2764));
  xor_4  g02388(.A(new_n2764), .B(new_n2761), .Y(new_n2765));
  nand_5 g02389(.A(pi219), .B(pi154), .Y(new_n2766));
  nand_5 g02390(.A(new_n2687), .B(new_n2686), .Y(new_n2767));
  nand_5 g02391(.A(new_n2688), .B(new_n2685), .Y(new_n2768));
  nand_5 g02392(.A(new_n2768), .B(new_n2767), .Y(new_n2769));
  xor_4  g02393(.A(new_n2769), .B(new_n2766), .Y(new_n2770));
  xor_4  g02394(.A(new_n2770), .B(new_n2765), .Y(new_n2771));
  xor_4  g02395(.A(new_n2771), .B(new_n2760), .Y(new_n2772));
  xor_4  g02396(.A(new_n2772), .B(new_n2759), .Y(new_n2773));
  xor_4  g02397(.A(new_n2773), .B(new_n2755), .Y(new_n2774));
  not_8  g02398(.A(new_n2697), .Y(new_n2775));
  nor_5  g02399(.A(new_n2707), .B(new_n2775), .Y(new_n2776));
  or_6   g02400(.A(new_n2705), .B(new_n2704), .Y(new_n2777));
  not_8  g02401(.A(new_n2702), .Y(new_n2778));
  nand_5 g02402(.A(new_n2706), .B(new_n2778), .Y(new_n2779));
  nand_5 g02403(.A(new_n2779), .B(new_n2777), .Y(new_n2780));
  nand_5 g02404(.A(pi142), .B(pi130), .Y(new_n2781));
  nand_5 g02405(.A(pi170), .B(pi099), .Y(new_n2782));
  nand_5 g02406(.A(pi169), .B(pi073), .Y(new_n2783));
  nand_5 g02407(.A(pi123), .B(pi004), .Y(new_n2784));
  xor_4  g02408(.A(new_n2784), .B(new_n2783), .Y(new_n2785));
  xor_4  g02409(.A(new_n2785), .B(new_n2782), .Y(new_n2786));
  nand_5 g02410(.A(pi071), .B(pi003), .Y(new_n2787));
  nand_5 g02411(.A(new_n2700), .B(new_n2699), .Y(new_n2788));
  nand_5 g02412(.A(new_n2701), .B(new_n2698), .Y(new_n2789));
  nand_5 g02413(.A(new_n2789), .B(new_n2788), .Y(new_n2790));
  xor_4  g02414(.A(new_n2790), .B(new_n2787), .Y(new_n2791));
  xor_4  g02415(.A(new_n2791), .B(new_n2786), .Y(new_n2792));
  xor_4  g02416(.A(new_n2792), .B(new_n2781), .Y(new_n2793));
  xor_4  g02417(.A(new_n2793), .B(new_n2780), .Y(new_n2794));
  xor_4  g02418(.A(new_n2794), .B(new_n2776), .Y(new_n2795));
  xnor_4 g02419(.A(new_n2795), .B(new_n2774), .Y(new_n2796));
  xnor_4 g02420(.A(new_n2796), .B(new_n2754), .Y(new_n2797));
  not_8  g02421(.A(new_n2797), .Y(new_n2798));
  xnor_4 g02422(.A(new_n2750), .B(new_n2730), .Y(new_n2799));
  or_6   g02423(.A(new_n2799), .B(new_n2798), .Y(new_n2800));
  nand_5 g02424(.A(new_n2800), .B(new_n2751), .Y(new_n2801));
  nand_5 g02425(.A(new_n2795), .B(new_n2774), .Y(new_n2802));
  or_6   g02426(.A(new_n2796), .B(new_n2754), .Y(new_n2803));
  nand_5 g02427(.A(new_n2803), .B(new_n2802), .Y(new_n2804));
  nor_5  g02428(.A(new_n2792), .B(new_n2781), .Y(new_n2805));
  and_6  g02429(.A(new_n2793), .B(new_n2780), .Y(new_n2806));
  nor_5  g02430(.A(new_n2806), .B(new_n2805), .Y(new_n2807));
  nand_5 g02431(.A(new_n2790), .B(new_n2787), .Y(new_n2808));
  nand_5 g02432(.A(new_n2791), .B(new_n2786), .Y(new_n2809));
  nand_5 g02433(.A(new_n2809), .B(new_n2808), .Y(new_n2810));
  nand_5 g02434(.A(pi169), .B(pi130), .Y(new_n2811));
  nor_5  g02435(.A(new_n2811), .B(new_n2787), .Y(new_n2812));
  nand_5 g02436(.A(pi130), .B(pi071), .Y(new_n2813));
  nand_5 g02437(.A(pi169), .B(pi003), .Y(new_n2814));
  nand_5 g02438(.A(new_n2814), .B(new_n2813), .Y(new_n2815));
  not_8  g02439(.A(new_n2815), .Y(new_n2816));
  nor_5  g02440(.A(new_n2816), .B(new_n2812), .Y(new_n2817));
  not_8  g02441(.A(new_n2817), .Y(new_n2818));
  nand_5 g02442(.A(pi099), .B(pi004), .Y(new_n2819));
  nand_5 g02443(.A(pi170), .B(pi023), .Y(new_n2820));
  nand_5 g02444(.A(new_n2820), .B(new_n2819), .Y(new_n2821));
  nand_5 g02445(.A(pi023), .B(pi004), .Y(new_n2822));
  nor_5  g02446(.A(new_n2822), .B(new_n2782), .Y(new_n2823));
  not_8  g02447(.A(new_n2823), .Y(new_n2824));
  nand_5 g02448(.A(new_n2824), .B(new_n2821), .Y(new_n2825));
  nand_5 g02449(.A(pi123), .B(pi073), .Y(new_n2826));
  nand_5 g02450(.A(new_n2784), .B(new_n2783), .Y(new_n2827));
  nand_5 g02451(.A(new_n2785), .B(new_n2782), .Y(new_n2828));
  nand_5 g02452(.A(new_n2828), .B(new_n2827), .Y(new_n2829));
  xor_4  g02453(.A(new_n2829), .B(new_n2826), .Y(new_n2830));
  xor_4  g02454(.A(new_n2830), .B(new_n2825), .Y(new_n2831));
  xor_4  g02455(.A(new_n2831), .B(new_n2818), .Y(new_n2832));
  xor_4  g02456(.A(new_n2832), .B(new_n2810), .Y(new_n2833));
  xor_4  g02457(.A(new_n2833), .B(new_n2807), .Y(new_n2834));
  and_6  g02458(.A(new_n2794), .B(new_n2776), .Y(new_n2835));
  nand_5 g02459(.A(pi142), .B(pi124), .Y(new_n2836));
  xor_4  g02460(.A(new_n2836), .B(new_n2835), .Y(new_n2837));
  xor_4  g02461(.A(new_n2837), .B(new_n2834), .Y(new_n2838));
  nand_5 g02462(.A(new_n2773), .B(new_n2755), .Y(new_n2839));
  nand_5 g02463(.A(pi087), .B(pi006), .Y(new_n2840));
  xor_4  g02464(.A(new_n2840), .B(new_n2839), .Y(new_n2841));
  nor_5  g02465(.A(new_n2771), .B(new_n2760), .Y(new_n2842));
  and_6  g02466(.A(new_n2772), .B(new_n2759), .Y(new_n2843));
  or_6   g02467(.A(new_n2843), .B(new_n2842), .Y(new_n2844));
  nand_5 g02468(.A(pi219), .B(pi095), .Y(new_n2845));
  nand_5 g02469(.A(pi154), .B(pi102), .Y(new_n2846));
  and_6  g02470(.A(new_n2846), .B(new_n2845), .Y(new_n2847));
  nand_5 g02471(.A(pi102), .B(pi095), .Y(new_n2848));
  nor_5  g02472(.A(new_n2848), .B(new_n2766), .Y(new_n2849));
  or_6   g02473(.A(new_n2849), .B(new_n2847), .Y(new_n2850));
  nand_5 g02474(.A(pi158), .B(pi122), .Y(new_n2851));
  nand_5 g02475(.A(pi254), .B(pi135), .Y(new_n2852));
  nand_5 g02476(.A(new_n2852), .B(new_n2851), .Y(new_n2853));
  nand_5 g02477(.A(pi158), .B(pi135), .Y(new_n2854));
  nor_5  g02478(.A(new_n2854), .B(new_n2762), .Y(new_n2855));
  not_8  g02479(.A(new_n2855), .Y(new_n2856));
  nand_5 g02480(.A(new_n2856), .B(new_n2853), .Y(new_n2857));
  nand_5 g02481(.A(pi089), .B(pi001), .Y(new_n2858));
  nand_5 g02482(.A(new_n2763), .B(new_n2762), .Y(new_n2859));
  nand_5 g02483(.A(new_n2764), .B(new_n2761), .Y(new_n2860));
  nand_5 g02484(.A(new_n2860), .B(new_n2859), .Y(new_n2861));
  xor_4  g02485(.A(new_n2861), .B(new_n2858), .Y(new_n2862));
  xor_4  g02486(.A(new_n2862), .B(new_n2857), .Y(new_n2863));
  xnor_4 g02487(.A(new_n2863), .B(new_n2850), .Y(new_n2864));
  nand_5 g02488(.A(new_n2769), .B(new_n2766), .Y(new_n2865));
  nand_5 g02489(.A(new_n2770), .B(new_n2765), .Y(new_n2866));
  nand_5 g02490(.A(new_n2866), .B(new_n2865), .Y(new_n2867));
  xor_4  g02491(.A(new_n2867), .B(new_n2864), .Y(new_n2868));
  xnor_4 g02492(.A(new_n2868), .B(new_n2844), .Y(new_n2869));
  xor_4  g02493(.A(new_n2869), .B(new_n2841), .Y(new_n2870));
  xnor_4 g02494(.A(new_n2870), .B(new_n2838), .Y(new_n2871));
  xor_4  g02495(.A(new_n2871), .B(new_n2804), .Y(new_n2872));
  nor_5  g02496(.A(new_n2743), .B(new_n2732), .Y(new_n2873));
  not_8  g02497(.A(new_n2744), .Y(new_n2874));
  nor_5  g02498(.A(new_n2748), .B(new_n2874), .Y(new_n2875));
  nor_5  g02499(.A(new_n2875), .B(new_n2873), .Y(new_n2876));
  nand_5 g02500(.A(pi172), .B(pi041), .Y(new_n2877));
  nand_5 g02501(.A(pi198), .B(pi182), .Y(new_n2878));
  and_6  g02502(.A(new_n2878), .B(new_n2877), .Y(new_n2879));
  nand_5 g02503(.A(pi198), .B(pi041), .Y(new_n2880));
  nor_5  g02504(.A(new_n2880), .B(new_n2738), .Y(new_n2881));
  or_6   g02505(.A(new_n2881), .B(new_n2879), .Y(new_n2882));
  nand_5 g02506(.A(new_n2735), .B(new_n2734), .Y(new_n2883));
  nand_5 g02507(.A(new_n2736), .B(new_n2733), .Y(new_n2884));
  nand_5 g02508(.A(new_n2884), .B(new_n2883), .Y(new_n2885));
  nand_5 g02509(.A(pi216), .B(pi120), .Y(new_n2886));
  nand_5 g02510(.A(pi076), .B(pi062), .Y(new_n2887));
  nand_5 g02511(.A(pi079), .B(pi065), .Y(new_n2888));
  nand_5 g02512(.A(new_n2888), .B(new_n2887), .Y(new_n2889));
  nand_5 g02513(.A(pi079), .B(pi062), .Y(new_n2890));
  nor_5  g02514(.A(new_n2890), .B(new_n2734), .Y(new_n2891));
  not_8  g02515(.A(new_n2891), .Y(new_n2892));
  nand_5 g02516(.A(new_n2892), .B(new_n2889), .Y(new_n2893));
  xor_4  g02517(.A(new_n2893), .B(new_n2886), .Y(new_n2894));
  xor_4  g02518(.A(new_n2894), .B(new_n2885), .Y(new_n2895));
  xor_4  g02519(.A(new_n2895), .B(new_n2882), .Y(new_n2896));
  nand_5 g02520(.A(new_n2741), .B(new_n2738), .Y(new_n2897));
  nand_5 g02521(.A(new_n2742), .B(new_n2737), .Y(new_n2898));
  nand_5 g02522(.A(new_n2898), .B(new_n2897), .Y(new_n2899));
  xor_4  g02523(.A(new_n2899), .B(new_n2896), .Y(new_n2900));
  xor_4  g02524(.A(new_n2900), .B(new_n2876), .Y(new_n2901));
  not_8  g02525(.A(new_n2731), .Y(new_n2902));
  nor_5  g02526(.A(new_n2749), .B(new_n2902), .Y(new_n2903));
  nand_5 g02527(.A(pi165), .B(pi138), .Y(new_n2904));
  xor_4  g02528(.A(new_n2904), .B(new_n2903), .Y(new_n2905));
  xor_4  g02529(.A(new_n2905), .B(new_n2901), .Y(new_n2906));
  xnor_4 g02530(.A(new_n2906), .B(new_n2872), .Y(new_n2907));
  xor_4  g02531(.A(new_n2907), .B(new_n2801), .Y(new_n2908));
  nand_5 g02532(.A(pi092), .B(pi020), .Y(new_n2909));
  nand_5 g02533(.A(pi190), .B(pi060), .Y(new_n2910));
  nand_5 g02534(.A(pi229), .B(pi160), .Y(new_n2911));
  or_6   g02535(.A(new_n2911), .B(new_n2910), .Y(new_n2912));
  nand_5 g02536(.A(new_n2912), .B(new_n2909), .Y(new_n2913));
  nand_5 g02537(.A(new_n2911), .B(new_n2910), .Y(new_n2914));
  nand_5 g02538(.A(new_n2914), .B(new_n2913), .Y(new_n2915));
  nand_5 g02539(.A(pi160), .B(pi067), .Y(new_n2916));
  xor_4  g02540(.A(new_n2916), .B(new_n2915), .Y(new_n2917));
  nand_5 g02541(.A(pi223), .B(pi190), .Y(new_n2918));
  nand_5 g02542(.A(pi229), .B(pi020), .Y(new_n2919));
  nand_5 g02543(.A(pi092), .B(pi060), .Y(new_n2920));
  xor_4  g02544(.A(new_n2920), .B(new_n2919), .Y(new_n2921));
  xor_4  g02545(.A(new_n2921), .B(new_n2918), .Y(new_n2922));
  not_8  g02546(.A(new_n2922), .Y(new_n2923));
  xor_4  g02547(.A(new_n2923), .B(new_n2917), .Y(new_n2924));
  nand_5 g02548(.A(pi190), .B(pi160), .Y(new_n2925));
  not_8  g02549(.A(new_n2925), .Y(new_n2926));
  nor_5  g02550(.A(new_n2926), .B(new_n2909), .Y(new_n2927));
  and_6  g02551(.A(new_n2914), .B(new_n2912), .Y(new_n2928));
  or_6   g02552(.A(new_n2928), .B(new_n2927), .Y(new_n2929));
  nor_5  g02553(.A(new_n2929), .B(new_n2909), .Y(new_n2930));
  nand_5 g02554(.A(new_n2930), .B(new_n2924), .Y(new_n2931));
  not_8  g02555(.A(new_n2931), .Y(new_n2932));
  nor_5  g02556(.A(new_n2916), .B(new_n2915), .Y(new_n2933));
  nand_5 g02557(.A(new_n2923), .B(new_n2917), .Y(new_n2934));
  not_8  g02558(.A(new_n2934), .Y(new_n2935));
  nor_5  g02559(.A(new_n2935), .B(new_n2933), .Y(new_n2936));
  not_8  g02560(.A(new_n2936), .Y(new_n2937));
  nand_5 g02561(.A(pi160), .B(pi053), .Y(new_n2938));
  nand_5 g02562(.A(pi190), .B(pi101), .Y(new_n2939));
  nand_5 g02563(.A(pi229), .B(pi060), .Y(new_n2940));
  nand_5 g02564(.A(pi223), .B(pi092), .Y(new_n2941));
  xor_4  g02565(.A(new_n2941), .B(new_n2940), .Y(new_n2942));
  xor_4  g02566(.A(new_n2942), .B(new_n2939), .Y(new_n2943));
  nand_5 g02567(.A(pi067), .B(pi020), .Y(new_n2944));
  nand_5 g02568(.A(new_n2920), .B(new_n2919), .Y(new_n2945));
  nand_5 g02569(.A(new_n2921), .B(new_n2918), .Y(new_n2946));
  nand_5 g02570(.A(new_n2946), .B(new_n2945), .Y(new_n2947));
  xor_4  g02571(.A(new_n2947), .B(new_n2944), .Y(new_n2948));
  xor_4  g02572(.A(new_n2948), .B(new_n2943), .Y(new_n2949));
  xor_4  g02573(.A(new_n2949), .B(new_n2938), .Y(new_n2950));
  xor_4  g02574(.A(new_n2950), .B(new_n2937), .Y(new_n2951));
  nand_5 g02575(.A(new_n2951), .B(new_n2932), .Y(new_n2952));
  nand_5 g02576(.A(pi185), .B(pi160), .Y(new_n2953));
  xor_4  g02577(.A(new_n2953), .B(new_n2952), .Y(new_n2954));
  nand_5 g02578(.A(new_n2947), .B(new_n2944), .Y(new_n2955));
  nand_5 g02579(.A(new_n2948), .B(new_n2943), .Y(new_n2956));
  nand_5 g02580(.A(new_n2956), .B(new_n2955), .Y(new_n2957));
  nand_5 g02581(.A(pi229), .B(pi223), .Y(new_n2958));
  nand_5 g02582(.A(new_n2941), .B(new_n2940), .Y(new_n2959));
  nand_5 g02583(.A(new_n2942), .B(new_n2939), .Y(new_n2960));
  nand_5 g02584(.A(new_n2960), .B(new_n2959), .Y(new_n2961));
  nand_5 g02585(.A(pi225), .B(pi092), .Y(new_n2962));
  nor_5  g02586(.A(new_n2962), .B(new_n2939), .Y(new_n2963));
  not_8  g02587(.A(new_n2963), .Y(new_n2964));
  nand_5 g02588(.A(pi225), .B(pi190), .Y(new_n2965));
  nand_5 g02589(.A(pi101), .B(pi092), .Y(new_n2966));
  nand_5 g02590(.A(new_n2966), .B(new_n2965), .Y(new_n2967));
  nand_5 g02591(.A(new_n2967), .B(new_n2964), .Y(new_n2968));
  xnor_4 g02592(.A(new_n2968), .B(new_n2961), .Y(new_n2969));
  xor_4  g02593(.A(new_n2969), .B(new_n2958), .Y(new_n2970));
  not_8  g02594(.A(new_n2970), .Y(new_n2971));
  xor_4  g02595(.A(new_n2971), .B(new_n2957), .Y(new_n2972));
  nand_5 g02596(.A(pi060), .B(pi053), .Y(new_n2973));
  nor_5  g02597(.A(new_n2973), .B(new_n2944), .Y(new_n2974));
  not_8  g02598(.A(new_n2974), .Y(new_n2975));
  nand_5 g02599(.A(pi067), .B(pi060), .Y(new_n2976));
  nand_5 g02600(.A(pi053), .B(pi020), .Y(new_n2977));
  nand_5 g02601(.A(new_n2977), .B(new_n2976), .Y(new_n2978));
  nand_5 g02602(.A(new_n2978), .B(new_n2975), .Y(new_n2979));
  xor_4  g02603(.A(new_n2979), .B(new_n2972), .Y(new_n2980));
  nor_5  g02604(.A(new_n2949), .B(new_n2938), .Y(new_n2981));
  and_6  g02605(.A(new_n2950), .B(new_n2937), .Y(new_n2982));
  nor_5  g02606(.A(new_n2982), .B(new_n2981), .Y(new_n2983));
  xor_4  g02607(.A(new_n2983), .B(new_n2980), .Y(new_n2984));
  xor_4  g02608(.A(new_n2984), .B(new_n2954), .Y(new_n2985));
  nand_5 g02609(.A(new_n2985), .B(new_n2908), .Y(new_n2986));
  xor_4  g02610(.A(new_n2930), .B(new_n2924), .Y(new_n2987));
  not_8  g02611(.A(new_n2987), .Y(new_n2988));
  xnor_4 g02612(.A(new_n2712), .B(new_n2630), .Y(new_n2989));
  nor_5  g02613(.A(new_n2989), .B(new_n2925), .Y(new_n2990));
  nand_5 g02614(.A(pi160), .B(pi092), .Y(new_n2991));
  nand_5 g02615(.A(pi190), .B(pi020), .Y(new_n2992));
  xor_4  g02616(.A(new_n2992), .B(new_n2991), .Y(new_n2993));
  nand_5 g02617(.A(new_n2993), .B(new_n2990), .Y(new_n2994));
  xor_4  g02618(.A(new_n2720), .B(new_n2719), .Y(new_n2995));
  xnor_4 g02619(.A(new_n2993), .B(new_n2990), .Y(new_n2996));
  or_6   g02620(.A(new_n2996), .B(new_n2995), .Y(new_n2997));
  and_6  g02621(.A(new_n2997), .B(new_n2994), .Y(new_n2998));
  nand_5 g02622(.A(new_n2927), .B(new_n2914), .Y(new_n2999));
  nand_5 g02623(.A(new_n2999), .B(new_n2929), .Y(new_n3000));
  and_6  g02624(.A(new_n3000), .B(new_n2998), .Y(new_n3001));
  xnor_4 g02625(.A(new_n3000), .B(new_n2998), .Y(new_n3002));
  xor_4  g02626(.A(new_n2726), .B(new_n2725), .Y(new_n3003));
  nor_5  g02627(.A(new_n3003), .B(new_n3002), .Y(new_n3004));
  or_6   g02628(.A(new_n3004), .B(new_n3001), .Y(new_n3005));
  nor_5  g02629(.A(new_n3005), .B(new_n2988), .Y(new_n3006));
  xor_4  g02630(.A(new_n2728), .B(new_n2711), .Y(new_n3007));
  xor_4  g02631(.A(new_n3005), .B(new_n2987), .Y(new_n3008));
  nor_5  g02632(.A(new_n3008), .B(new_n3007), .Y(new_n3009));
  nor_5  g02633(.A(new_n3009), .B(new_n3006), .Y(new_n3010));
  xor_4  g02634(.A(new_n2951), .B(new_n2931), .Y(new_n3011));
  or_6   g02635(.A(new_n3011), .B(new_n3010), .Y(new_n3012));
  xor_4  g02636(.A(new_n3011), .B(new_n3010), .Y(new_n3013));
  xor_4  g02637(.A(new_n2799), .B(new_n2797), .Y(new_n3014));
  nand_5 g02638(.A(new_n3014), .B(new_n3013), .Y(new_n3015));
  nand_5 g02639(.A(new_n3015), .B(new_n3012), .Y(new_n3016));
  xor_4  g02640(.A(new_n2985), .B(new_n2908), .Y(new_n3017));
  nand_5 g02641(.A(new_n3017), .B(new_n3016), .Y(new_n3018));
  nand_5 g02642(.A(new_n3018), .B(new_n2986), .Y(new_n3019));
  nor_5  g02643(.A(new_n2906), .B(new_n2872), .Y(new_n3020));
  nor_5  g02644(.A(new_n2907), .B(new_n2801), .Y(new_n3021));
  nor_5  g02645(.A(new_n3021), .B(new_n3020), .Y(new_n3022));
  not_8  g02646(.A(new_n2836), .Y(new_n3023));
  nor_5  g02647(.A(new_n3023), .B(new_n2835), .Y(new_n3024));
  not_8  g02648(.A(new_n3024), .Y(new_n3025));
  or_6   g02649(.A(new_n2837), .B(new_n2834), .Y(new_n3026));
  nand_5 g02650(.A(new_n3026), .B(new_n3025), .Y(new_n3027));
  nor_5  g02651(.A(new_n2833), .B(new_n2807), .Y(new_n3028));
  not_8  g02652(.A(new_n3028), .Y(new_n3029));
  nand_5 g02653(.A(new_n2829), .B(new_n2826), .Y(new_n3030));
  nand_5 g02654(.A(new_n2830), .B(new_n2825), .Y(new_n3031));
  nand_5 g02655(.A(new_n3031), .B(new_n3030), .Y(new_n3032));
  nand_5 g02656(.A(pi215), .B(pi142), .Y(new_n3033));
  nand_5 g02657(.A(pi124), .B(pi071), .Y(new_n3034));
  xor_4  g02658(.A(new_n3034), .B(new_n3033), .Y(new_n3035));
  xor_4  g02659(.A(new_n3035), .B(new_n2811), .Y(new_n3036));
  xor_4  g02660(.A(new_n3036), .B(new_n3032), .Y(new_n3037));
  nand_5 g02661(.A(pi123), .B(pi003), .Y(new_n3038));
  xor_4  g02662(.A(new_n3038), .B(new_n2823), .Y(new_n3039));
  nand_5 g02663(.A(pi099), .B(pi073), .Y(new_n3040));
  nand_5 g02664(.A(pi170), .B(pi155), .Y(new_n3041));
  xor_4  g02665(.A(new_n3041), .B(new_n3040), .Y(new_n3042));
  xor_4  g02666(.A(new_n3042), .B(new_n2822), .Y(new_n3043));
  xor_4  g02667(.A(new_n3043), .B(new_n3039), .Y(new_n3044));
  xor_4  g02668(.A(new_n3044), .B(new_n3037), .Y(new_n3045));
  nand_5 g02669(.A(new_n2831), .B(new_n2818), .Y(new_n3046));
  nand_5 g02670(.A(new_n2832), .B(new_n2810), .Y(new_n3047));
  nand_5 g02671(.A(new_n3047), .B(new_n3046), .Y(new_n3048));
  xor_4  g02672(.A(new_n3048), .B(new_n2812), .Y(new_n3049));
  xor_4  g02673(.A(new_n3049), .B(new_n3045), .Y(new_n3050));
  xor_4  g02674(.A(new_n3050), .B(new_n3029), .Y(new_n3051));
  xor_4  g02675(.A(new_n3051), .B(new_n3027), .Y(new_n3052));
  nand_5 g02676(.A(new_n2840), .B(new_n2839), .Y(new_n3053));
  nand_5 g02677(.A(new_n2869), .B(new_n2841), .Y(new_n3054));
  nand_5 g02678(.A(new_n3054), .B(new_n3053), .Y(new_n3055));
  nand_5 g02679(.A(new_n2868), .B(new_n2844), .Y(new_n3056));
  nand_5 g02680(.A(pi154), .B(pi001), .Y(new_n3057));
  xor_4  g02681(.A(new_n3057), .B(new_n2855), .Y(new_n3058));
  nand_5 g02682(.A(pi122), .B(pi089), .Y(new_n3059));
  nand_5 g02683(.A(pi254), .B(pi059), .Y(new_n3060));
  xor_4  g02684(.A(new_n3060), .B(new_n3059), .Y(new_n3061));
  xor_4  g02685(.A(new_n3061), .B(new_n2854), .Y(new_n3062));
  xor_4  g02686(.A(new_n3062), .B(new_n3058), .Y(new_n3063));
  nand_5 g02687(.A(new_n2861), .B(new_n2858), .Y(new_n3064));
  nand_5 g02688(.A(new_n2862), .B(new_n2857), .Y(new_n3065));
  nand_5 g02689(.A(new_n3065), .B(new_n3064), .Y(new_n3066));
  nand_5 g02690(.A(pi209), .B(pi087), .Y(new_n3067));
  nand_5 g02691(.A(pi219), .B(pi006), .Y(new_n3068));
  xor_4  g02692(.A(new_n3068), .B(new_n2848), .Y(new_n3069));
  xor_4  g02693(.A(new_n3069), .B(new_n3067), .Y(new_n3070));
  xor_4  g02694(.A(new_n3070), .B(new_n3066), .Y(new_n3071));
  xor_4  g02695(.A(new_n3071), .B(new_n3063), .Y(new_n3072));
  nor_5  g02696(.A(new_n2867), .B(new_n2864), .Y(new_n3073));
  nand_5 g02697(.A(new_n3073), .B(new_n2849), .Y(new_n3074));
  or_6   g02698(.A(new_n2867), .B(new_n2864), .Y(new_n3075));
  nor_5  g02699(.A(new_n2863), .B(new_n2850), .Y(new_n3076));
  nor_5  g02700(.A(new_n3076), .B(new_n2849), .Y(new_n3077));
  nand_5 g02701(.A(new_n3077), .B(new_n3075), .Y(new_n3078));
  nand_5 g02702(.A(new_n3078), .B(new_n3074), .Y(new_n3079));
  xor_4  g02703(.A(new_n3079), .B(new_n3072), .Y(new_n3080));
  xor_4  g02704(.A(new_n3080), .B(new_n3056), .Y(new_n3081));
  xor_4  g02705(.A(new_n3081), .B(new_n3055), .Y(new_n3082));
  xor_4  g02706(.A(new_n3082), .B(new_n3052), .Y(new_n3083));
  nor_5  g02707(.A(new_n2870), .B(new_n2838), .Y(new_n3084));
  not_8  g02708(.A(new_n2804), .Y(new_n3085));
  nor_5  g02709(.A(new_n2871), .B(new_n3085), .Y(new_n3086));
  or_6   g02710(.A(new_n3086), .B(new_n3084), .Y(new_n3087));
  xnor_4 g02711(.A(new_n3087), .B(new_n3083), .Y(new_n3088));
  or_6   g02712(.A(new_n2900), .B(new_n2876), .Y(new_n3089));
  not_8  g02713(.A(new_n2896), .Y(new_n3090));
  nor_5  g02714(.A(new_n2899), .B(new_n3090), .Y(new_n3091));
  not_8  g02715(.A(new_n3091), .Y(new_n3092));
  nor_5  g02716(.A(new_n2895), .B(new_n2882), .Y(new_n3093));
  nor_5  g02717(.A(new_n3093), .B(new_n2881), .Y(new_n3094));
  nand_5 g02718(.A(new_n3094), .B(new_n3092), .Y(new_n3095));
  nand_5 g02719(.A(new_n3091), .B(new_n2881), .Y(new_n3096));
  nand_5 g02720(.A(new_n3096), .B(new_n3095), .Y(new_n3097));
  nand_5 g02721(.A(pi120), .B(pi076), .Y(new_n3098));
  nand_5 g02722(.A(pi251), .B(pi065), .Y(new_n3099));
  xor_4  g02723(.A(new_n3099), .B(new_n3098), .Y(new_n3100));
  xor_4  g02724(.A(new_n3100), .B(new_n2890), .Y(new_n3101));
  nand_5 g02725(.A(pi216), .B(pi172), .Y(new_n3102));
  xor_4  g02726(.A(new_n3102), .B(new_n2891), .Y(new_n3103));
  xor_4  g02727(.A(new_n3103), .B(new_n3101), .Y(new_n3104));
  nand_5 g02728(.A(new_n2893), .B(new_n2886), .Y(new_n3105));
  nand_5 g02729(.A(new_n2894), .B(new_n2885), .Y(new_n3106));
  nand_5 g02730(.A(new_n3106), .B(new_n3105), .Y(new_n3107));
  nand_5 g02731(.A(pi197), .B(pi138), .Y(new_n3108));
  nand_5 g02732(.A(pi182), .B(pi165), .Y(new_n3109));
  xor_4  g02733(.A(new_n3109), .B(new_n3108), .Y(new_n3110));
  xor_4  g02734(.A(new_n3110), .B(new_n2880), .Y(new_n3111));
  xnor_4 g02735(.A(new_n3111), .B(new_n3107), .Y(new_n3112));
  xor_4  g02736(.A(new_n3112), .B(new_n3104), .Y(new_n3113));
  not_8  g02737(.A(new_n3113), .Y(new_n3114));
  xor_4  g02738(.A(new_n3114), .B(new_n3097), .Y(new_n3115));
  xor_4  g02739(.A(new_n3115), .B(new_n3089), .Y(new_n3116));
  not_8  g02740(.A(new_n2903), .Y(new_n3117));
  nand_5 g02741(.A(new_n2904), .B(new_n3117), .Y(new_n3118));
  or_6   g02742(.A(new_n2905), .B(new_n2901), .Y(new_n3119));
  nand_5 g02743(.A(new_n3119), .B(new_n3118), .Y(new_n3120));
  xor_4  g02744(.A(new_n3120), .B(new_n3116), .Y(new_n3121));
  xnor_4 g02745(.A(new_n3121), .B(new_n3088), .Y(new_n3122));
  xor_4  g02746(.A(new_n3122), .B(new_n3022), .Y(new_n3123));
  nand_5 g02747(.A(new_n2953), .B(new_n2952), .Y(new_n3124));
  not_8  g02748(.A(new_n2984), .Y(new_n3125));
  nand_5 g02749(.A(new_n3125), .B(new_n2954), .Y(new_n3126));
  nand_5 g02750(.A(new_n3126), .B(new_n3124), .Y(new_n3127));
  nor_5  g02751(.A(new_n2983), .B(new_n2980), .Y(new_n3128));
  nand_5 g02752(.A(new_n2971), .B(new_n2957), .Y(new_n3129));
  nand_5 g02753(.A(new_n2979), .B(new_n2972), .Y(new_n3130));
  nand_5 g02754(.A(new_n3130), .B(new_n3129), .Y(new_n3131));
  nand_5 g02755(.A(new_n3131), .B(new_n2975), .Y(new_n3132));
  nor_5  g02756(.A(new_n2971), .B(new_n2957), .Y(new_n3133));
  nand_5 g02757(.A(new_n2974), .B(new_n3133), .Y(new_n3134));
  nand_5 g02758(.A(new_n3134), .B(new_n3132), .Y(new_n3135));
  nand_5 g02759(.A(pi223), .B(pi067), .Y(new_n3136));
  xor_4  g02760(.A(new_n3136), .B(new_n2963), .Y(new_n3137));
  nand_5 g02761(.A(pi190), .B(pi177), .Y(new_n3138));
  nand_5 g02762(.A(pi229), .B(pi101), .Y(new_n3139));
  xor_4  g02763(.A(new_n3139), .B(new_n3138), .Y(new_n3140));
  xor_4  g02764(.A(new_n3140), .B(new_n2962), .Y(new_n3141));
  xor_4  g02765(.A(new_n3141), .B(new_n3137), .Y(new_n3142));
  nand_5 g02766(.A(pi160), .B(pi030), .Y(new_n3143));
  nand_5 g02767(.A(pi185), .B(pi020), .Y(new_n3144));
  xor_4  g02768(.A(new_n3144), .B(new_n3143), .Y(new_n3145));
  xnor_4 g02769(.A(new_n3145), .B(new_n2973), .Y(new_n3146));
  nor_5  g02770(.A(new_n2968), .B(new_n2961), .Y(new_n3147));
  nor_5  g02771(.A(new_n2969), .B(new_n2958), .Y(new_n3148));
  nor_5  g02772(.A(new_n3148), .B(new_n3147), .Y(new_n3149));
  xor_4  g02773(.A(new_n3149), .B(new_n3146), .Y(new_n3150));
  xor_4  g02774(.A(new_n3150), .B(new_n3142), .Y(new_n3151));
  not_8  g02775(.A(new_n3151), .Y(new_n3152));
  xor_4  g02776(.A(new_n3152), .B(new_n3135), .Y(new_n3153));
  xor_4  g02777(.A(new_n3153), .B(new_n3128), .Y(new_n3154));
  xor_4  g02778(.A(new_n3154), .B(new_n3127), .Y(new_n3155));
  xnor_4 g02779(.A(new_n3155), .B(new_n3123), .Y(new_n3156));
  xnor_4 g02780(.A(new_n3156), .B(new_n3019), .Y(po007));
  nand_5 g02781(.A(pi208), .B(pi186), .Y(new_n3158));
  nand_5 g02782(.A(pi168), .B(pi132), .Y(new_n3159));
  or_6   g02783(.A(new_n3159), .B(new_n3158), .Y(new_n3160));
  nand_5 g02784(.A(pi186), .B(pi168), .Y(new_n3161));
  nand_5 g02785(.A(pi208), .B(pi132), .Y(new_n3162));
  nand_5 g02786(.A(new_n3162), .B(new_n3161), .Y(new_n3163));
  nand_5 g02787(.A(new_n3163), .B(new_n3160), .Y(new_n3164));
  nand_5 g02788(.A(pi236), .B(pi109), .Y(new_n3165));
  not_8  g02789(.A(new_n3165), .Y(new_n3166));
  nand_5 g02790(.A(pi226), .B(pi213), .Y(new_n3167));
  xor_4  g02791(.A(new_n3167), .B(new_n3166), .Y(new_n3168));
  or_6   g02792(.A(new_n3168), .B(new_n3159), .Y(new_n3169));
  nor_5  g02793(.A(new_n3169), .B(new_n3164), .Y(new_n3170));
  nor_5  g02794(.A(new_n3167), .B(new_n3165), .Y(new_n3171));
  not_8  g02795(.A(new_n3171), .Y(new_n3172));
  nand_5 g02796(.A(pi212), .B(pi207), .Y(new_n3173));
  or_6   g02797(.A(new_n3173), .B(new_n3167), .Y(new_n3174));
  nand_5 g02798(.A(pi213), .B(pi207), .Y(new_n3175));
  nand_5 g02799(.A(pi226), .B(pi212), .Y(new_n3176));
  nand_5 g02800(.A(new_n3176), .B(new_n3175), .Y(new_n3177));
  nand_5 g02801(.A(new_n3177), .B(new_n3174), .Y(new_n3178));
  nand_5 g02802(.A(pi241), .B(pi014), .Y(new_n3179));
  or_6   g02803(.A(new_n3179), .B(new_n3165), .Y(new_n3180));
  nand_5 g02804(.A(pi241), .B(pi109), .Y(new_n3181));
  nand_5 g02805(.A(pi236), .B(pi014), .Y(new_n3182));
  nand_5 g02806(.A(new_n3182), .B(new_n3181), .Y(new_n3183));
  nand_5 g02807(.A(new_n3183), .B(new_n3180), .Y(new_n3184));
  xor_4  g02808(.A(new_n3184), .B(new_n3178), .Y(new_n3185));
  xor_4  g02809(.A(new_n3185), .B(new_n3172), .Y(new_n3186));
  xnor_4 g02810(.A(new_n3169), .B(new_n3164), .Y(new_n3187));
  nor_5  g02811(.A(new_n3187), .B(new_n3186), .Y(new_n3188));
  nor_5  g02812(.A(new_n3188), .B(new_n3170), .Y(new_n3189));
  nand_5 g02813(.A(pi139), .B(pi132), .Y(new_n3190));
  nand_5 g02814(.A(pi168), .B(pi058), .Y(new_n3191));
  xor_4  g02815(.A(new_n3191), .B(new_n3158), .Y(new_n3192));
  xor_4  g02816(.A(new_n3192), .B(new_n3190), .Y(new_n3193));
  xnor_4 g02817(.A(new_n3193), .B(new_n3160), .Y(new_n3194));
  nor_5  g02818(.A(new_n3194), .B(new_n3189), .Y(new_n3195));
  xor_4  g02819(.A(new_n3194), .B(new_n3189), .Y(new_n3196));
  nand_5 g02820(.A(pi226), .B(pi104), .Y(new_n3197));
  nand_5 g02821(.A(pi213), .B(pi066), .Y(new_n3198));
  xor_4  g02822(.A(new_n3198), .B(new_n3173), .Y(new_n3199));
  xor_4  g02823(.A(new_n3199), .B(new_n3197), .Y(new_n3200));
  xnor_4 g02824(.A(new_n3200), .B(new_n3174), .Y(new_n3201));
  nand_5 g02825(.A(new_n3184), .B(new_n3178), .Y(new_n3202));
  nand_5 g02826(.A(new_n3185), .B(new_n3172), .Y(new_n3203));
  nand_5 g02827(.A(new_n3203), .B(new_n3202), .Y(new_n3204));
  xor_4  g02828(.A(new_n3204), .B(new_n3201), .Y(new_n3205));
  nand_5 g02829(.A(pi236), .B(pi173), .Y(new_n3206));
  nand_5 g02830(.A(pi161), .B(pi109), .Y(new_n3207));
  xor_4  g02831(.A(new_n3207), .B(new_n3206), .Y(new_n3208));
  nor_5  g02832(.A(new_n3208), .B(new_n3179), .Y(new_n3209));
  nand_5 g02833(.A(new_n3209), .B(new_n3166), .Y(new_n3210));
  not_8  g02834(.A(new_n3210), .Y(new_n3211));
  nand_5 g02835(.A(new_n3208), .B(new_n3179), .Y(new_n3212));
  nand_5 g02836(.A(new_n3212), .B(new_n3180), .Y(new_n3213));
  nor_5  g02837(.A(new_n3213), .B(new_n3209), .Y(new_n3214));
  nor_5  g02838(.A(new_n3214), .B(new_n3211), .Y(new_n3215));
  xor_4  g02839(.A(new_n3215), .B(new_n3205), .Y(new_n3216));
  and_6  g02840(.A(new_n3216), .B(new_n3196), .Y(new_n3217));
  nor_5  g02841(.A(new_n3217), .B(new_n3195), .Y(new_n3218));
  nor_5  g02842(.A(new_n3193), .B(new_n3160), .Y(new_n3219));
  nand_5 g02843(.A(pi132), .B(pi035), .Y(new_n3220));
  nand_5 g02844(.A(pi208), .B(pi058), .Y(new_n3221));
  nand_5 g02845(.A(pi186), .B(pi139), .Y(new_n3222));
  xor_4  g02846(.A(new_n3222), .B(new_n3221), .Y(new_n3223));
  xor_4  g02847(.A(new_n3223), .B(new_n3220), .Y(new_n3224));
  not_8  g02848(.A(new_n3224), .Y(new_n3225));
  nand_5 g02849(.A(pi211), .B(pi168), .Y(new_n3226));
  nand_5 g02850(.A(new_n3191), .B(new_n3158), .Y(new_n3227));
  nand_5 g02851(.A(new_n3192), .B(new_n3190), .Y(new_n3228));
  nand_5 g02852(.A(new_n3228), .B(new_n3227), .Y(new_n3229));
  xor_4  g02853(.A(new_n3229), .B(new_n3226), .Y(new_n3230));
  xor_4  g02854(.A(new_n3230), .B(new_n3225), .Y(new_n3231));
  xnor_4 g02855(.A(new_n3231), .B(new_n3219), .Y(new_n3232));
  xnor_4 g02856(.A(new_n3232), .B(new_n3218), .Y(new_n3233));
  nand_5 g02857(.A(new_n3204), .B(new_n3201), .Y(new_n3234));
  not_8  g02858(.A(new_n3215), .Y(new_n3235));
  nand_5 g02859(.A(new_n3235), .B(new_n3205), .Y(new_n3236));
  nand_5 g02860(.A(new_n3236), .B(new_n3234), .Y(new_n3237));
  nor_5  g02861(.A(new_n3200), .B(new_n3174), .Y(new_n3238));
  nand_5 g02862(.A(pi212), .B(pi066), .Y(new_n3239));
  nand_5 g02863(.A(pi207), .B(pi104), .Y(new_n3240));
  nand_5 g02864(.A(pi226), .B(pi013), .Y(new_n3241));
  xor_4  g02865(.A(new_n3241), .B(new_n3240), .Y(new_n3242));
  xor_4  g02866(.A(new_n3242), .B(new_n3239), .Y(new_n3243));
  nand_5 g02867(.A(pi213), .B(pi055), .Y(new_n3244));
  nand_5 g02868(.A(new_n3198), .B(new_n3173), .Y(new_n3245));
  nand_5 g02869(.A(new_n3199), .B(new_n3197), .Y(new_n3246));
  nand_5 g02870(.A(new_n3246), .B(new_n3245), .Y(new_n3247));
  xor_4  g02871(.A(new_n3247), .B(new_n3244), .Y(new_n3248));
  xor_4  g02872(.A(new_n3248), .B(new_n3243), .Y(new_n3249));
  xor_4  g02873(.A(new_n3249), .B(new_n3238), .Y(new_n3250));
  nand_5 g02874(.A(pi161), .B(pi014), .Y(new_n3251));
  nand_5 g02875(.A(pi141), .B(pi109), .Y(new_n3252));
  nand_5 g02876(.A(pi241), .B(pi173), .Y(new_n3253));
  xor_4  g02877(.A(new_n3253), .B(new_n3252), .Y(new_n3254));
  xor_4  g02878(.A(new_n3254), .B(new_n3251), .Y(new_n3255));
  nand_5 g02879(.A(pi236), .B(pi230), .Y(new_n3256));
  nand_5 g02880(.A(new_n3207), .B(new_n3206), .Y(new_n3257));
  nand_5 g02881(.A(new_n3212), .B(new_n3257), .Y(new_n3258));
  xor_4  g02882(.A(new_n3258), .B(new_n3256), .Y(new_n3259));
  xor_4  g02883(.A(new_n3259), .B(new_n3255), .Y(new_n3260));
  xor_4  g02884(.A(new_n3260), .B(new_n3211), .Y(new_n3261));
  nand_5 g02885(.A(new_n3261), .B(new_n3250), .Y(new_n3262));
  or_6   g02886(.A(new_n3261), .B(new_n3250), .Y(new_n3263));
  nand_5 g02887(.A(new_n3263), .B(new_n3262), .Y(new_n3264));
  xor_4  g02888(.A(new_n3264), .B(new_n3237), .Y(new_n3265));
  xnor_4 g02889(.A(new_n3265), .B(new_n3233), .Y(new_n3266));
  nand_5 g02890(.A(pi077), .B(pi029), .Y(new_n3267));
  nand_5 g02891(.A(pi069), .B(pi052), .Y(new_n3268));
  nand_5 g02892(.A(pi244), .B(pi131), .Y(new_n3269));
  xor_4  g02893(.A(new_n3269), .B(new_n3268), .Y(new_n3270));
  xor_4  g02894(.A(new_n3270), .B(new_n3267), .Y(new_n3271));
  nand_5 g02895(.A(pi131), .B(pi029), .Y(new_n3272));
  nor_5  g02896(.A(new_n3272), .B(new_n3268), .Y(new_n3273));
  not_8  g02897(.A(new_n3273), .Y(new_n3274));
  xor_4  g02898(.A(new_n3274), .B(new_n3271), .Y(new_n3275));
  not_8  g02899(.A(new_n3275), .Y(new_n3276));
  xnor_4 g02900(.A(new_n3168), .B(new_n3159), .Y(new_n3277));
  or_6   g02901(.A(new_n3277), .B(new_n3272), .Y(new_n3278));
  nand_5 g02902(.A(pi131), .B(pi069), .Y(new_n3279));
  nand_5 g02903(.A(pi052), .B(pi029), .Y(new_n3280));
  nand_5 g02904(.A(new_n3280), .B(new_n3279), .Y(new_n3281));
  nand_5 g02905(.A(new_n3281), .B(new_n3274), .Y(new_n3282));
  nand_5 g02906(.A(new_n3282), .B(new_n3278), .Y(new_n3283));
  xnor_4 g02907(.A(new_n3187), .B(new_n3186), .Y(new_n3284));
  xor_4  g02908(.A(new_n3282), .B(new_n3278), .Y(new_n3285));
  nand_5 g02909(.A(new_n3285), .B(new_n3284), .Y(new_n3286));
  nand_5 g02910(.A(new_n3286), .B(new_n3283), .Y(new_n3287));
  nand_5 g02911(.A(new_n3287), .B(new_n3276), .Y(new_n3288));
  xor_4  g02912(.A(new_n3216), .B(new_n3196), .Y(new_n3289));
  xor_4  g02913(.A(new_n3287), .B(new_n3275), .Y(new_n3290));
  or_6   g02914(.A(new_n3290), .B(new_n3289), .Y(new_n3291));
  nand_5 g02915(.A(new_n3291), .B(new_n3288), .Y(new_n3292));
  or_6   g02916(.A(new_n3274), .B(new_n3271), .Y(new_n3293));
  nand_5 g02917(.A(pi133), .B(pi029), .Y(new_n3294));
  nand_5 g02918(.A(pi244), .B(pi052), .Y(new_n3295));
  nand_5 g02919(.A(pi077), .B(pi069), .Y(new_n3296));
  xor_4  g02920(.A(new_n3296), .B(new_n3295), .Y(new_n3297));
  xor_4  g02921(.A(new_n3297), .B(new_n3294), .Y(new_n3298));
  nand_5 g02922(.A(pi150), .B(pi131), .Y(new_n3299));
  nand_5 g02923(.A(new_n3269), .B(new_n3268), .Y(new_n3300));
  nand_5 g02924(.A(new_n3270), .B(new_n3267), .Y(new_n3301));
  nand_5 g02925(.A(new_n3301), .B(new_n3300), .Y(new_n3302));
  xor_4  g02926(.A(new_n3302), .B(new_n3299), .Y(new_n3303));
  xor_4  g02927(.A(new_n3303), .B(new_n3298), .Y(new_n3304));
  xnor_4 g02928(.A(new_n3304), .B(new_n3293), .Y(new_n3305));
  xor_4  g02929(.A(new_n3305), .B(new_n3292), .Y(new_n3306));
  xor_4  g02930(.A(new_n3306), .B(new_n3266), .Y(po008));
  nand_5 g02931(.A(pi208), .B(pi062), .Y(new_n3308));
  nand_5 g02932(.A(pi168), .B(pi120), .Y(new_n3309));
  xor_4  g02933(.A(new_n3309), .B(new_n3308), .Y(new_n3310));
  nand_5 g02934(.A(pi139), .B(pi065), .Y(new_n3311));
  xor_4  g02935(.A(new_n3311), .B(new_n3310), .Y(new_n3312));
  nand_5 g02936(.A(pi168), .B(pi065), .Y(new_n3313));
  nor_5  g02937(.A(new_n3313), .B(new_n3308), .Y(new_n3314));
  not_8  g02938(.A(new_n3314), .Y(new_n3315));
  nor_5  g02939(.A(new_n3315), .B(new_n3312), .Y(new_n3316));
  not_8  g02940(.A(new_n3316), .Y(new_n3317));
  nand_5 g02941(.A(pi208), .B(pi120), .Y(new_n3318));
  nand_5 g02942(.A(pi065), .B(pi035), .Y(new_n3319));
  nand_5 g02943(.A(pi139), .B(pi062), .Y(new_n3320));
  xor_4  g02944(.A(new_n3320), .B(new_n3319), .Y(new_n3321));
  xor_4  g02945(.A(new_n3321), .B(new_n3318), .Y(new_n3322));
  nand_5 g02946(.A(pi172), .B(pi168), .Y(new_n3323));
  nand_5 g02947(.A(new_n3309), .B(new_n3308), .Y(new_n3324));
  nand_5 g02948(.A(new_n3311), .B(new_n3310), .Y(new_n3325));
  nand_5 g02949(.A(new_n3325), .B(new_n3324), .Y(new_n3326));
  xor_4  g02950(.A(new_n3326), .B(new_n3323), .Y(new_n3327));
  xor_4  g02951(.A(new_n3327), .B(new_n3322), .Y(new_n3328));
  xor_4  g02952(.A(new_n3328), .B(new_n3317), .Y(new_n3329));
  nand_5 g02953(.A(pi254), .B(pi161), .Y(new_n3330));
  nand_5 g02954(.A(pi241), .B(pi158), .Y(new_n3331));
  nand_5 g02955(.A(pi236), .B(pi089), .Y(new_n3332));
  xor_4  g02956(.A(new_n3332), .B(new_n3331), .Y(new_n3333));
  xnor_4 g02957(.A(new_n3333), .B(new_n3330), .Y(new_n3334));
  nand_5 g02958(.A(pi254), .B(pi236), .Y(new_n3335));
  or_6   g02959(.A(new_n3335), .B(new_n3331), .Y(new_n3336));
  not_8  g02960(.A(new_n3336), .Y(new_n3337));
  xor_4  g02961(.A(new_n3337), .B(new_n3334), .Y(new_n3338));
  not_8  g02962(.A(new_n3338), .Y(new_n3339));
  nand_5 g02963(.A(pi170), .B(pi104), .Y(new_n3340));
  nand_5 g02964(.A(pi213), .B(pi073), .Y(new_n3341));
  nor_5  g02965(.A(new_n3341), .B(new_n3340), .Y(new_n3342));
  nand_5 g02966(.A(pi212), .B(pi004), .Y(new_n3343));
  not_8  g02967(.A(new_n3343), .Y(new_n3344));
  nand_5 g02968(.A(pi213), .B(pi170), .Y(new_n3345));
  and_6  g02969(.A(new_n3345), .B(new_n3344), .Y(new_n3346));
  nand_5 g02970(.A(new_n3341), .B(new_n3340), .Y(new_n3347));
  nor_5  g02971(.A(new_n3347), .B(new_n3346), .Y(new_n3348));
  nor_5  g02972(.A(new_n3348), .B(new_n3342), .Y(new_n3349));
  nand_5 g02973(.A(new_n3347), .B(new_n3346), .Y(new_n3350));
  nand_5 g02974(.A(new_n3350), .B(new_n3349), .Y(new_n3351));
  nor_5  g02975(.A(new_n3351), .B(new_n3339), .Y(new_n3352));
  xor_4  g02976(.A(new_n3351), .B(new_n3338), .Y(new_n3353));
  nand_5 g02977(.A(pi236), .B(pi158), .Y(new_n3354));
  nand_5 g02978(.A(pi254), .B(pi241), .Y(new_n3355));
  nand_5 g02979(.A(new_n3355), .B(new_n3354), .Y(new_n3356));
  nand_5 g02980(.A(new_n3356), .B(new_n3336), .Y(new_n3357));
  nand_5 g02981(.A(pi213), .B(pi004), .Y(new_n3358));
  and_6  g02982(.A(pi212), .B(pi170), .Y(new_n3359));
  xor_4  g02983(.A(new_n3359), .B(new_n3358), .Y(new_n3360));
  nand_5 g02984(.A(new_n3360), .B(new_n3357), .Y(new_n3361));
  nor_5  g02985(.A(new_n3345), .B(new_n3335), .Y(new_n3362));
  xor_4  g02986(.A(new_n3360), .B(new_n3357), .Y(new_n3363));
  not_8  g02987(.A(new_n3363), .Y(new_n3364));
  or_6   g02988(.A(new_n3364), .B(new_n3362), .Y(new_n3365));
  nand_5 g02989(.A(new_n3365), .B(new_n3361), .Y(new_n3366));
  nor_5  g02990(.A(new_n3366), .B(new_n3353), .Y(new_n3367));
  nor_5  g02991(.A(new_n3367), .B(new_n3352), .Y(new_n3368));
  nand_5 g02992(.A(new_n3337), .B(new_n3334), .Y(new_n3369));
  nand_5 g02993(.A(pi161), .B(pi158), .Y(new_n3370));
  nand_5 g02994(.A(pi241), .B(pi089), .Y(new_n3371));
  nand_5 g02995(.A(pi254), .B(pi141), .Y(new_n3372));
  xor_4  g02996(.A(new_n3372), .B(new_n3371), .Y(new_n3373));
  xor_4  g02997(.A(new_n3373), .B(new_n3370), .Y(new_n3374));
  nand_5 g02998(.A(pi236), .B(pi154), .Y(new_n3375));
  nand_5 g02999(.A(new_n3332), .B(new_n3331), .Y(new_n3376));
  nand_5 g03000(.A(new_n3333), .B(new_n3330), .Y(new_n3377));
  nand_5 g03001(.A(new_n3377), .B(new_n3376), .Y(new_n3378));
  xnor_4 g03002(.A(new_n3378), .B(new_n3375), .Y(new_n3379));
  xnor_4 g03003(.A(new_n3379), .B(new_n3374), .Y(new_n3380));
  xnor_4 g03004(.A(new_n3380), .B(new_n3369), .Y(new_n3381));
  nor_5  g03005(.A(new_n3349), .B(new_n3343), .Y(new_n3382));
  nand_5 g03006(.A(pi170), .B(pi013), .Y(new_n3383));
  nand_5 g03007(.A(pi212), .B(pi073), .Y(new_n3384));
  nand_5 g03008(.A(pi104), .B(pi004), .Y(new_n3385));
  xor_4  g03009(.A(new_n3385), .B(new_n3384), .Y(new_n3386));
  xor_4  g03010(.A(new_n3386), .B(new_n3383), .Y(new_n3387));
  nand_5 g03011(.A(pi213), .B(pi003), .Y(new_n3388));
  or_6   g03012(.A(new_n3344), .B(new_n3342), .Y(new_n3389));
  nand_5 g03013(.A(new_n3389), .B(new_n3347), .Y(new_n3390));
  xnor_4 g03014(.A(new_n3390), .B(new_n3388), .Y(new_n3391));
  xnor_4 g03015(.A(new_n3391), .B(new_n3387), .Y(new_n3392));
  xor_4  g03016(.A(new_n3392), .B(new_n3382), .Y(new_n3393));
  xnor_4 g03017(.A(new_n3393), .B(new_n3381), .Y(new_n3394));
  xor_4  g03018(.A(new_n3394), .B(new_n3368), .Y(new_n3395));
  nor_5  g03019(.A(new_n3395), .B(new_n3329), .Y(new_n3396));
  xor_4  g03020(.A(new_n3314), .B(new_n3312), .Y(new_n3397));
  xnor_4 g03021(.A(new_n3366), .B(new_n3353), .Y(new_n3398));
  nand_5 g03022(.A(new_n3398), .B(new_n3397), .Y(new_n3399));
  xor_4  g03023(.A(new_n3398), .B(new_n3397), .Y(new_n3400));
  not_8  g03024(.A(new_n3313), .Y(new_n3401));
  xor_4  g03025(.A(new_n3345), .B(new_n3335), .Y(new_n3402));
  nand_5 g03026(.A(new_n3402), .B(new_n3401), .Y(new_n3403));
  nand_5 g03027(.A(pi168), .B(pi062), .Y(new_n3404));
  nand_5 g03028(.A(pi208), .B(pi065), .Y(new_n3405));
  nand_5 g03029(.A(new_n3405), .B(new_n3404), .Y(new_n3406));
  nand_5 g03030(.A(new_n3406), .B(new_n3315), .Y(new_n3407));
  nor_5  g03031(.A(new_n3407), .B(new_n3403), .Y(new_n3408));
  xnor_4 g03032(.A(new_n3407), .B(new_n3403), .Y(new_n3409));
  xor_4  g03033(.A(new_n3364), .B(new_n3362), .Y(new_n3410));
  nor_5  g03034(.A(new_n3410), .B(new_n3409), .Y(new_n3411));
  nor_5  g03035(.A(new_n3411), .B(new_n3408), .Y(new_n3412));
  nand_5 g03036(.A(new_n3412), .B(new_n3400), .Y(new_n3413));
  nand_5 g03037(.A(new_n3413), .B(new_n3399), .Y(new_n3414));
  not_8  g03038(.A(new_n3414), .Y(new_n3415));
  xnor_4 g03039(.A(new_n3395), .B(new_n3329), .Y(new_n3416));
  nor_5  g03040(.A(new_n3416), .B(new_n3415), .Y(new_n3417));
  or_6   g03041(.A(new_n3417), .B(new_n3396), .Y(new_n3418));
  nor_5  g03042(.A(new_n3328), .B(new_n3317), .Y(new_n3419));
  nand_5 g03043(.A(pi198), .B(pi168), .Y(new_n3420));
  nor_5  g03044(.A(new_n3326), .B(new_n3323), .Y(new_n3421));
  not_8  g03045(.A(new_n3327), .Y(new_n3422));
  nor_5  g03046(.A(new_n3422), .B(new_n3322), .Y(new_n3423));
  nor_5  g03047(.A(new_n3423), .B(new_n3421), .Y(new_n3424));
  xor_4  g03048(.A(new_n3424), .B(new_n3420), .Y(new_n3425));
  nand_5 g03049(.A(pi139), .B(pi120), .Y(new_n3426));
  nand_5 g03050(.A(pi062), .B(pi035), .Y(new_n3427));
  nand_5 g03051(.A(pi065), .B(pi015), .Y(new_n3428));
  xor_4  g03052(.A(new_n3428), .B(new_n3427), .Y(new_n3429));
  xor_4  g03053(.A(new_n3429), .B(new_n3426), .Y(new_n3430));
  nand_5 g03054(.A(pi208), .B(pi172), .Y(new_n3431));
  nand_5 g03055(.A(new_n3320), .B(new_n3319), .Y(new_n3432));
  nand_5 g03056(.A(new_n3321), .B(new_n3318), .Y(new_n3433));
  nand_5 g03057(.A(new_n3433), .B(new_n3432), .Y(new_n3434));
  xor_4  g03058(.A(new_n3434), .B(new_n3431), .Y(new_n3435));
  xnor_4 g03059(.A(new_n3435), .B(new_n3430), .Y(new_n3436));
  xor_4  g03060(.A(new_n3436), .B(new_n3425), .Y(new_n3437));
  xor_4  g03061(.A(new_n3437), .B(new_n3419), .Y(new_n3438));
  not_8  g03062(.A(new_n3438), .Y(new_n3439));
  xor_4  g03063(.A(new_n3439), .B(new_n3418), .Y(new_n3440));
  nor_5  g03064(.A(new_n3393), .B(new_n3381), .Y(new_n3441));
  nor_5  g03065(.A(new_n3394), .B(new_n3368), .Y(new_n3442));
  nor_5  g03066(.A(new_n3442), .B(new_n3441), .Y(new_n3443));
  nor_5  g03067(.A(new_n3380), .B(new_n3369), .Y(new_n3444));
  nand_5 g03068(.A(pi236), .B(pi095), .Y(new_n3445));
  nor_5  g03069(.A(new_n3378), .B(new_n3375), .Y(new_n3446));
  nor_5  g03070(.A(new_n3379), .B(new_n3374), .Y(new_n3447));
  nor_5  g03071(.A(new_n3447), .B(new_n3446), .Y(new_n3448));
  xor_4  g03072(.A(new_n3448), .B(new_n3445), .Y(new_n3449));
  nand_5 g03073(.A(pi158), .B(pi141), .Y(new_n3450));
  nand_5 g03074(.A(pi254), .B(pi090), .Y(new_n3451));
  nand_5 g03075(.A(pi161), .B(pi089), .Y(new_n3452));
  xor_4  g03076(.A(new_n3452), .B(new_n3451), .Y(new_n3453));
  xor_4  g03077(.A(new_n3453), .B(new_n3450), .Y(new_n3454));
  nand_5 g03078(.A(pi241), .B(pi154), .Y(new_n3455));
  and_6  g03079(.A(new_n3372), .B(new_n3371), .Y(new_n3456));
  and_6  g03080(.A(new_n3373), .B(new_n3370), .Y(new_n3457));
  or_6   g03081(.A(new_n3457), .B(new_n3456), .Y(new_n3458));
  xor_4  g03082(.A(new_n3458), .B(new_n3455), .Y(new_n3459));
  xnor_4 g03083(.A(new_n3459), .B(new_n3454), .Y(new_n3460));
  xor_4  g03084(.A(new_n3460), .B(new_n3449), .Y(new_n3461));
  xnor_4 g03085(.A(new_n3461), .B(new_n3444), .Y(new_n3462));
  xor_4  g03086(.A(new_n3462), .B(new_n3443), .Y(new_n3463));
  not_8  g03087(.A(new_n3382), .Y(new_n3464));
  nor_5  g03088(.A(new_n3392), .B(new_n3464), .Y(new_n3465));
  nand_5 g03089(.A(pi213), .B(pi130), .Y(new_n3466));
  nor_5  g03090(.A(new_n3390), .B(new_n3388), .Y(new_n3467));
  nor_5  g03091(.A(new_n3391), .B(new_n3387), .Y(new_n3468));
  nor_5  g03092(.A(new_n3468), .B(new_n3467), .Y(new_n3469));
  xor_4  g03093(.A(new_n3469), .B(new_n3466), .Y(new_n3470));
  nand_5 g03094(.A(pi104), .B(pi073), .Y(new_n3471));
  nand_5 g03095(.A(pi013), .B(pi004), .Y(new_n3472));
  nand_5 g03096(.A(pi170), .B(pi112), .Y(new_n3473));
  xor_4  g03097(.A(new_n3473), .B(new_n3472), .Y(new_n3474));
  xor_4  g03098(.A(new_n3474), .B(new_n3471), .Y(new_n3475));
  nand_5 g03099(.A(new_n3385), .B(new_n3384), .Y(new_n3476));
  nand_5 g03100(.A(new_n3386), .B(new_n3383), .Y(new_n3477));
  nand_5 g03101(.A(new_n3477), .B(new_n3476), .Y(new_n3478));
  nand_5 g03102(.A(pi212), .B(pi003), .Y(new_n3479));
  xor_4  g03103(.A(new_n3479), .B(new_n3478), .Y(new_n3480));
  xor_4  g03104(.A(new_n3480), .B(new_n3475), .Y(new_n3481));
  xnor_4 g03105(.A(new_n3481), .B(new_n3470), .Y(new_n3482));
  xnor_4 g03106(.A(new_n3482), .B(new_n3465), .Y(new_n3483));
  xnor_4 g03107(.A(new_n3483), .B(new_n3463), .Y(new_n3484));
  xor_4  g03108(.A(new_n3484), .B(new_n3440), .Y(new_n3485));
  nand_5 g03109(.A(pi131), .B(pi053), .Y(new_n3486));
  nand_5 g03110(.A(pi131), .B(pi067), .Y(new_n3487));
  nand_5 g03111(.A(pi229), .B(pi131), .Y(new_n3488));
  nand_5 g03112(.A(pi092), .B(pi052), .Y(new_n3489));
  nand_5 g03113(.A(new_n3489), .B(new_n3488), .Y(new_n3490));
  nand_5 g03114(.A(pi190), .B(pi077), .Y(new_n3491));
  xor_4  g03115(.A(new_n3489), .B(new_n3488), .Y(new_n3492));
  nand_5 g03116(.A(new_n3492), .B(new_n3491), .Y(new_n3493));
  nand_5 g03117(.A(new_n3493), .B(new_n3490), .Y(new_n3494));
  nor_5  g03118(.A(new_n3494), .B(new_n3487), .Y(new_n3495));
  nand_5 g03119(.A(pi229), .B(pi052), .Y(new_n3496));
  nand_5 g03120(.A(pi190), .B(pi133), .Y(new_n3497));
  nand_5 g03121(.A(pi092), .B(pi077), .Y(new_n3498));
  xor_4  g03122(.A(new_n3498), .B(new_n3497), .Y(new_n3499));
  xor_4  g03123(.A(new_n3499), .B(new_n3496), .Y(new_n3500));
  xor_4  g03124(.A(new_n3494), .B(new_n3487), .Y(new_n3501));
  not_8  g03125(.A(new_n3501), .Y(new_n3502));
  nor_5  g03126(.A(new_n3502), .B(new_n3500), .Y(new_n3503));
  nor_5  g03127(.A(new_n3503), .B(new_n3495), .Y(new_n3504));
  xor_4  g03128(.A(new_n3504), .B(new_n3486), .Y(new_n3505));
  nand_5 g03129(.A(pi229), .B(pi077), .Y(new_n3506));
  nand_5 g03130(.A(pi133), .B(pi092), .Y(new_n3507));
  nand_5 g03131(.A(pi190), .B(pi189), .Y(new_n3508));
  xor_4  g03132(.A(new_n3508), .B(new_n3507), .Y(new_n3509));
  xor_4  g03133(.A(new_n3509), .B(new_n3506), .Y(new_n3510));
  nand_5 g03134(.A(pi067), .B(pi052), .Y(new_n3511));
  nand_5 g03135(.A(new_n3498), .B(new_n3497), .Y(new_n3512));
  nand_5 g03136(.A(new_n3499), .B(new_n3496), .Y(new_n3513));
  nand_5 g03137(.A(new_n3513), .B(new_n3512), .Y(new_n3514));
  xor_4  g03138(.A(new_n3514), .B(new_n3511), .Y(new_n3515));
  xor_4  g03139(.A(new_n3515), .B(new_n3510), .Y(new_n3516));
  not_8  g03140(.A(new_n3516), .Y(new_n3517));
  xor_4  g03141(.A(new_n3517), .B(new_n3505), .Y(new_n3518));
  xor_4  g03142(.A(new_n3492), .B(new_n3491), .Y(new_n3519));
  not_8  g03143(.A(new_n3519), .Y(new_n3520));
  nand_5 g03144(.A(pi190), .B(pi131), .Y(new_n3521));
  nor_5  g03145(.A(new_n3521), .B(new_n3489), .Y(new_n3522));
  nand_5 g03146(.A(new_n3522), .B(new_n3520), .Y(new_n3523));
  xor_4  g03147(.A(new_n3501), .B(new_n3500), .Y(new_n3524));
  nor_5  g03148(.A(new_n3524), .B(new_n3523), .Y(new_n3525));
  xor_4  g03149(.A(new_n3525), .B(new_n3518), .Y(new_n3526));
  xor_4  g03150(.A(new_n3524), .B(new_n3523), .Y(new_n3527));
  xor_4  g03151(.A(new_n3416), .B(new_n3414), .Y(new_n3528));
  nor_5  g03152(.A(new_n3528), .B(new_n3527), .Y(new_n3529));
  xor_4  g03153(.A(new_n3402), .B(new_n3313), .Y(new_n3530));
  nor_5  g03154(.A(new_n3530), .B(new_n3521), .Y(new_n3531));
  not_8  g03155(.A(new_n3531), .Y(new_n3532));
  nand_5 g03156(.A(pi131), .B(pi092), .Y(new_n3533));
  nand_5 g03157(.A(pi190), .B(pi052), .Y(new_n3534));
  and_6  g03158(.A(new_n3534), .B(new_n3533), .Y(new_n3535));
  or_6   g03159(.A(new_n3535), .B(new_n3522), .Y(new_n3536));
  nand_5 g03160(.A(new_n3536), .B(new_n3532), .Y(new_n3537));
  xor_4  g03161(.A(new_n3536), .B(new_n3532), .Y(new_n3538));
  not_8  g03162(.A(new_n3538), .Y(new_n3539));
  xor_4  g03163(.A(new_n3410), .B(new_n3409), .Y(new_n3540));
  or_6   g03164(.A(new_n3540), .B(new_n3539), .Y(new_n3541));
  nand_5 g03165(.A(new_n3541), .B(new_n3537), .Y(new_n3542));
  xor_4  g03166(.A(new_n3522), .B(new_n3519), .Y(new_n3543));
  nor_5  g03167(.A(new_n3543), .B(new_n3542), .Y(new_n3544));
  not_8  g03168(.A(new_n3544), .Y(new_n3545));
  xor_4  g03169(.A(new_n3543), .B(new_n3542), .Y(new_n3546));
  xnor_4 g03170(.A(new_n3412), .B(new_n3400), .Y(new_n3547));
  nand_5 g03171(.A(new_n3547), .B(new_n3546), .Y(new_n3548));
  nand_5 g03172(.A(new_n3548), .B(new_n3545), .Y(new_n3549));
  xnor_4 g03173(.A(new_n3528), .B(new_n3527), .Y(new_n3550));
  nor_5  g03174(.A(new_n3550), .B(new_n3549), .Y(new_n3551));
  nor_5  g03175(.A(new_n3551), .B(new_n3529), .Y(new_n3552));
  xnor_4 g03176(.A(new_n3552), .B(new_n3526), .Y(new_n3553));
  xnor_4 g03177(.A(new_n3553), .B(new_n3485), .Y(po009));
  nand_5 g03178(.A(pi168), .B(pi162), .Y(new_n3555));
  nand_5 g03179(.A(pi236), .B(pi051), .Y(new_n3556));
  nand_5 g03180(.A(pi213), .B(pi188), .Y(new_n3557));
  xnor_4 g03181(.A(new_n3557), .B(new_n3556), .Y(new_n3558));
  xnor_4 g03182(.A(new_n3558), .B(new_n3555), .Y(new_n3559));
  nand_5 g03183(.A(pi143), .B(pi131), .Y(new_n3560));
  xor_4  g03184(.A(new_n3560), .B(new_n3559), .Y(po010));
  xnor_4 g03185(.A(new_n1608), .B(new_n1496), .Y(po011));
  xnor_4 g03186(.A(new_n3550), .B(new_n3549), .Y(po012));
  nand_5 g03187(.A(pi173), .B(pi135), .Y(new_n3564));
  nand_5 g03188(.A(pi059), .B(pi014), .Y(new_n3565));
  xor_4  g03189(.A(new_n3565), .B(new_n3564), .Y(new_n3566));
  nand_5 g03190(.A(pi211), .B(pi076), .Y(new_n3567));
  nand_5 g03191(.A(pi079), .B(pi058), .Y(new_n3568));
  xor_4  g03192(.A(new_n3568), .B(new_n3567), .Y(new_n3569));
  nand_5 g03193(.A(pi226), .B(pi086), .Y(new_n3570));
  nand_5 g03194(.A(pi207), .B(pi155), .Y(new_n3571));
  xnor_4 g03195(.A(new_n3571), .B(new_n3570), .Y(new_n3572));
  xor_4  g03196(.A(new_n3572), .B(new_n3569), .Y(new_n3573));
  xor_4  g03197(.A(new_n3573), .B(new_n3566), .Y(new_n3574));
  nand_5 g03198(.A(pi221), .B(pi060), .Y(new_n3575));
  nand_5 g03199(.A(pi196), .B(pi020), .Y(new_n3576));
  nand_5 g03200(.A(pi184), .B(pi160), .Y(new_n3577));
  xor_4  g03201(.A(new_n3577), .B(new_n3576), .Y(new_n3578));
  xor_4  g03202(.A(new_n3578), .B(new_n3575), .Y(new_n3579));
  nand_5 g03203(.A(pi225), .B(pi029), .Y(new_n3580));
  nand_5 g03204(.A(pi101), .B(pi069), .Y(new_n3581));
  nand_5 g03205(.A(new_n3581), .B(new_n3580), .Y(new_n3582));
  nand_5 g03206(.A(pi101), .B(pi029), .Y(new_n3583));
  nand_5 g03207(.A(pi225), .B(pi069), .Y(new_n3584));
  nor_5  g03208(.A(new_n3584), .B(new_n3583), .Y(new_n3585));
  not_8  g03209(.A(new_n3585), .Y(new_n3586));
  nand_5 g03210(.A(new_n3586), .B(new_n3582), .Y(new_n3587));
  nand_5 g03211(.A(pi244), .B(pi223), .Y(new_n3588));
  nand_5 g03212(.A(new_n3588), .B(new_n3587), .Y(new_n3589));
  nand_5 g03213(.A(pi223), .B(pi069), .Y(new_n3590));
  nand_5 g03214(.A(new_n3590), .B(new_n3583), .Y(new_n3591));
  nand_5 g03215(.A(pi244), .B(pi060), .Y(new_n3592));
  xor_4  g03216(.A(new_n3590), .B(new_n3583), .Y(new_n3593));
  nand_5 g03217(.A(new_n3593), .B(new_n3592), .Y(new_n3594));
  nand_5 g03218(.A(new_n3594), .B(new_n3591), .Y(new_n3595));
  xor_4  g03219(.A(new_n3588), .B(new_n3587), .Y(new_n3596));
  nand_5 g03220(.A(new_n3596), .B(new_n3595), .Y(new_n3597));
  nand_5 g03221(.A(new_n3597), .B(new_n3589), .Y(new_n3598));
  nand_5 g03222(.A(new_n3598), .B(new_n3579), .Y(new_n3599));
  xor_4  g03223(.A(new_n3598), .B(new_n3579), .Y(new_n3600));
  nand_5 g03224(.A(pi177), .B(pi029), .Y(new_n3601));
  nand_5 g03225(.A(pi244), .B(pi101), .Y(new_n3602));
  xor_4  g03226(.A(new_n3602), .B(new_n3601), .Y(new_n3603));
  xor_4  g03227(.A(new_n3603), .B(new_n3584), .Y(new_n3604));
  nand_5 g03228(.A(pi223), .B(pi150), .Y(new_n3605));
  xor_4  g03229(.A(new_n3605), .B(new_n3585), .Y(new_n3606));
  xor_4  g03230(.A(new_n3606), .B(new_n3604), .Y(new_n3607));
  not_8  g03231(.A(new_n3607), .Y(new_n3608));
  nand_5 g03232(.A(new_n3608), .B(new_n3600), .Y(new_n3609));
  nand_5 g03233(.A(new_n3609), .B(new_n3599), .Y(new_n3610));
  nand_5 g03234(.A(pi218), .B(pi138), .Y(new_n3611));
  nand_5 g03235(.A(pi195), .B(pi182), .Y(new_n3612));
  nand_5 g03236(.A(new_n3612), .B(new_n3611), .Y(new_n3613));
  nand_5 g03237(.A(pi199), .B(pi041), .Y(new_n3614));
  xor_4  g03238(.A(new_n3612), .B(new_n3611), .Y(new_n3615));
  nand_5 g03239(.A(new_n3615), .B(new_n3614), .Y(new_n3616));
  nand_5 g03240(.A(new_n3616), .B(new_n3613), .Y(new_n3617));
  xor_4  g03241(.A(new_n3617), .B(new_n3610), .Y(new_n3618));
  nand_5 g03242(.A(pi135), .B(pi014), .Y(new_n3619));
  nand_5 g03243(.A(pi122), .B(pi109), .Y(new_n3620));
  nor_5  g03244(.A(new_n3620), .B(new_n3619), .Y(new_n3621));
  not_8  g03245(.A(new_n3621), .Y(new_n3622));
  nand_5 g03246(.A(pi230), .B(pi001), .Y(new_n3623));
  or_6   g03247(.A(new_n3623), .B(new_n3622), .Y(new_n3624));
  xor_4  g03248(.A(new_n3623), .B(new_n3622), .Y(new_n3625));
  nand_5 g03249(.A(pi173), .B(pi122), .Y(new_n3626));
  nand_5 g03250(.A(pi109), .B(pi059), .Y(new_n3627));
  xor_4  g03251(.A(new_n3627), .B(new_n3626), .Y(new_n3628));
  xor_4  g03252(.A(new_n3628), .B(new_n3619), .Y(new_n3629));
  not_8  g03253(.A(new_n3629), .Y(new_n3630));
  nand_5 g03254(.A(new_n3630), .B(new_n3625), .Y(new_n3631));
  nand_5 g03255(.A(new_n3631), .B(new_n3624), .Y(new_n3632));
  nand_5 g03256(.A(pi137), .B(pi029), .Y(new_n3633));
  nand_5 g03257(.A(pi169), .B(pi025), .Y(new_n3634));
  nand_5 g03258(.A(pi071), .B(pi025), .Y(new_n3635));
  nand_5 g03259(.A(pi239), .B(pi142), .Y(new_n3636));
  nand_5 g03260(.A(new_n3636), .B(new_n3635), .Y(new_n3637));
  nand_5 g03261(.A(pi169), .B(pi002), .Y(new_n3638));
  xor_4  g03262(.A(new_n3636), .B(new_n3635), .Y(new_n3639));
  nand_5 g03263(.A(new_n3639), .B(new_n3638), .Y(new_n3640));
  nand_5 g03264(.A(new_n3640), .B(new_n3637), .Y(new_n3641));
  xor_4  g03265(.A(new_n3641), .B(new_n3634), .Y(new_n3642));
  xor_4  g03266(.A(new_n3642), .B(new_n3633), .Y(new_n3643));
  xor_4  g03267(.A(new_n3643), .B(new_n3632), .Y(new_n3644));
  xor_4  g03268(.A(new_n3644), .B(new_n3618), .Y(new_n3645));
  nand_5 g03269(.A(pi066), .B(pi023), .Y(new_n3646));
  nand_5 g03270(.A(pi216), .B(pi199), .Y(new_n3647));
  xor_4  g03271(.A(new_n3647), .B(new_n3646), .Y(new_n3648));
  nand_5 g03272(.A(pi186), .B(pi079), .Y(new_n3649));
  nand_5 g03273(.A(pi076), .B(pi058), .Y(new_n3650));
  nand_5 g03274(.A(new_n3650), .B(new_n3649), .Y(new_n3651));
  nand_5 g03275(.A(pi251), .B(pi132), .Y(new_n3652));
  xor_4  g03276(.A(new_n3650), .B(new_n3649), .Y(new_n3653));
  nand_5 g03277(.A(new_n3653), .B(new_n3652), .Y(new_n3654));
  nand_5 g03278(.A(new_n3654), .B(new_n3651), .Y(new_n3655));
  nand_5 g03279(.A(pi218), .B(pi182), .Y(new_n3656));
  nand_5 g03280(.A(pi243), .B(pi142), .Y(new_n3657));
  xor_4  g03281(.A(new_n3657), .B(new_n3656), .Y(new_n3658));
  xor_4  g03282(.A(new_n3658), .B(new_n3655), .Y(new_n3659));
  nand_5 g03283(.A(pi199), .B(pi138), .Y(new_n3660));
  nand_5 g03284(.A(pi211), .B(pi138), .Y(new_n3661));
  nand_5 g03285(.A(pi186), .B(pi182), .Y(new_n3662));
  nand_5 g03286(.A(pi138), .B(pi058), .Y(new_n3663));
  nand_5 g03287(.A(new_n3663), .B(new_n3662), .Y(new_n3664));
  xor_4  g03288(.A(new_n3663), .B(new_n3662), .Y(new_n3665));
  nand_5 g03289(.A(pi132), .B(pi041), .Y(new_n3666));
  nand_5 g03290(.A(new_n3666), .B(new_n3665), .Y(new_n3667));
  nand_5 g03291(.A(new_n3667), .B(new_n3664), .Y(new_n3668));
  nor_5  g03292(.A(new_n3668), .B(new_n3661), .Y(new_n3669));
  xor_4  g03293(.A(new_n3668), .B(new_n3661), .Y(new_n3670));
  nand_5 g03294(.A(pi182), .B(pi058), .Y(new_n3671));
  nand_5 g03295(.A(pi186), .B(pi041), .Y(new_n3672));
  nand_5 g03296(.A(pi216), .B(pi132), .Y(new_n3673));
  xor_4  g03297(.A(new_n3673), .B(new_n3672), .Y(new_n3674));
  xor_4  g03298(.A(new_n3674), .B(new_n3671), .Y(new_n3675));
  not_8  g03299(.A(new_n3675), .Y(new_n3676));
  and_6  g03300(.A(new_n3676), .B(new_n3670), .Y(new_n3677));
  nor_5  g03301(.A(new_n3677), .B(new_n3669), .Y(new_n3678));
  nor_5  g03302(.A(new_n3678), .B(new_n3660), .Y(new_n3679));
  xnor_4 g03303(.A(new_n3678), .B(new_n3660), .Y(new_n3680));
  nand_5 g03304(.A(pi132), .B(pi076), .Y(new_n3681));
  nand_5 g03305(.A(pi058), .B(pi041), .Y(new_n3682));
  nand_5 g03306(.A(pi216), .B(pi186), .Y(new_n3683));
  xor_4  g03307(.A(new_n3683), .B(new_n3682), .Y(new_n3684));
  xor_4  g03308(.A(new_n3684), .B(new_n3681), .Y(new_n3685));
  nand_5 g03309(.A(pi211), .B(pi182), .Y(new_n3686));
  nand_5 g03310(.A(new_n3673), .B(new_n3672), .Y(new_n3687));
  nand_5 g03311(.A(new_n3674), .B(new_n3671), .Y(new_n3688));
  nand_5 g03312(.A(new_n3688), .B(new_n3687), .Y(new_n3689));
  xor_4  g03313(.A(new_n3689), .B(new_n3686), .Y(new_n3690));
  xor_4  g03314(.A(new_n3690), .B(new_n3685), .Y(new_n3691));
  nor_5  g03315(.A(new_n3691), .B(new_n3680), .Y(new_n3692));
  nor_5  g03316(.A(new_n3692), .B(new_n3679), .Y(new_n3693));
  nand_5 g03317(.A(new_n3689), .B(new_n3686), .Y(new_n3694));
  nand_5 g03318(.A(new_n3690), .B(new_n3685), .Y(new_n3695));
  nand_5 g03319(.A(new_n3695), .B(new_n3694), .Y(new_n3696));
  nand_5 g03320(.A(pi211), .B(pi041), .Y(new_n3697));
  nand_5 g03321(.A(pi199), .B(pi182), .Y(new_n3698));
  and_6  g03322(.A(new_n3698), .B(new_n3697), .Y(new_n3699));
  nor_5  g03323(.A(new_n3686), .B(new_n3614), .Y(new_n3700));
  or_6   g03324(.A(new_n3700), .B(new_n3699), .Y(new_n3701));
  nand_5 g03325(.A(new_n3683), .B(new_n3682), .Y(new_n3702));
  nand_5 g03326(.A(new_n3684), .B(new_n3681), .Y(new_n3703));
  nand_5 g03327(.A(new_n3703), .B(new_n3702), .Y(new_n3704));
  nand_5 g03328(.A(pi132), .B(pi079), .Y(new_n3705));
  nand_5 g03329(.A(pi186), .B(pi076), .Y(new_n3706));
  nand_5 g03330(.A(new_n3706), .B(new_n3705), .Y(new_n3707));
  nor_5  g03331(.A(new_n3681), .B(new_n3649), .Y(new_n3708));
  not_8  g03332(.A(new_n3708), .Y(new_n3709));
  nand_5 g03333(.A(new_n3709), .B(new_n3707), .Y(new_n3710));
  nand_5 g03334(.A(pi216), .B(pi058), .Y(new_n3711));
  xor_4  g03335(.A(new_n3711), .B(new_n3710), .Y(new_n3712));
  xor_4  g03336(.A(new_n3712), .B(new_n3704), .Y(new_n3713));
  xor_4  g03337(.A(new_n3713), .B(new_n3701), .Y(new_n3714));
  xor_4  g03338(.A(new_n3714), .B(new_n3696), .Y(new_n3715));
  or_6   g03339(.A(new_n3715), .B(new_n3693), .Y(new_n3716));
  nand_5 g03340(.A(new_n3711), .B(new_n3710), .Y(new_n3717));
  nand_5 g03341(.A(new_n3712), .B(new_n3704), .Y(new_n3718));
  nand_5 g03342(.A(new_n3718), .B(new_n3717), .Y(new_n3719));
  xor_4  g03343(.A(new_n3615), .B(new_n3614), .Y(new_n3720));
  xor_4  g03344(.A(new_n3720), .B(new_n3719), .Y(new_n3721));
  not_8  g03345(.A(new_n3721), .Y(new_n3722));
  nand_5 g03346(.A(pi216), .B(pi211), .Y(new_n3723));
  xor_4  g03347(.A(new_n3723), .B(new_n3708), .Y(new_n3724));
  xor_4  g03348(.A(new_n3653), .B(new_n3652), .Y(new_n3725));
  xnor_4 g03349(.A(new_n3725), .B(new_n3724), .Y(new_n3726));
  xor_4  g03350(.A(new_n3726), .B(new_n3722), .Y(new_n3727));
  not_8  g03351(.A(new_n3714), .Y(new_n3728));
  nor_5  g03352(.A(new_n3728), .B(new_n3696), .Y(new_n3729));
  nand_5 g03353(.A(new_n3729), .B(new_n3700), .Y(new_n3730));
  nor_5  g03354(.A(new_n3713), .B(new_n3701), .Y(new_n3731));
  nor_5  g03355(.A(new_n3731), .B(new_n3700), .Y(new_n3732));
  not_8  g03356(.A(new_n3732), .Y(new_n3733));
  nor_5  g03357(.A(new_n3733), .B(new_n3729), .Y(new_n3734));
  not_8  g03358(.A(new_n3734), .Y(new_n3735));
  nand_5 g03359(.A(new_n3735), .B(new_n3730), .Y(new_n3736));
  xor_4  g03360(.A(new_n3736), .B(new_n3727), .Y(new_n3737));
  nor_5  g03361(.A(new_n3737), .B(new_n3716), .Y(new_n3738));
  xor_4  g03362(.A(new_n3737), .B(new_n3716), .Y(new_n3739));
  not_8  g03363(.A(new_n3739), .Y(new_n3740));
  nand_5 g03364(.A(pi195), .B(pi138), .Y(new_n3741));
  xor_4  g03365(.A(new_n3715), .B(new_n3693), .Y(new_n3742));
  not_8  g03366(.A(new_n3742), .Y(new_n3743));
  nor_5  g03367(.A(new_n3743), .B(new_n3741), .Y(new_n3744));
  xor_4  g03368(.A(new_n3691), .B(new_n3680), .Y(new_n3745));
  xor_4  g03369(.A(new_n3675), .B(new_n3670), .Y(new_n3746));
  xor_4  g03370(.A(new_n3666), .B(new_n3665), .Y(new_n3747));
  nand_5 g03371(.A(pi138), .B(pi132), .Y(new_n3748));
  or_6   g03372(.A(new_n3748), .B(new_n3662), .Y(new_n3749));
  nor_5  g03373(.A(new_n3749), .B(new_n3747), .Y(new_n3750));
  not_8  g03374(.A(new_n3750), .Y(new_n3751));
  nor_5  g03375(.A(new_n3751), .B(new_n3746), .Y(new_n3752));
  nand_5 g03376(.A(new_n3752), .B(new_n3745), .Y(new_n3753));
  xor_4  g03377(.A(new_n3742), .B(new_n3741), .Y(new_n3754));
  nor_5  g03378(.A(new_n3754), .B(new_n3753), .Y(new_n3755));
  nor_5  g03379(.A(new_n3755), .B(new_n3744), .Y(new_n3756));
  nor_5  g03380(.A(new_n3756), .B(new_n3740), .Y(new_n3757));
  nor_5  g03381(.A(new_n3757), .B(new_n3738), .Y(new_n3758));
  nand_5 g03382(.A(new_n3602), .B(new_n3601), .Y(new_n3759));
  nand_5 g03383(.A(new_n3603), .B(new_n3584), .Y(new_n3760));
  nand_5 g03384(.A(new_n3760), .B(new_n3759), .Y(new_n3761));
  nand_5 g03385(.A(pi196), .B(pi060), .Y(new_n3762));
  xor_4  g03386(.A(new_n3762), .B(new_n3761), .Y(new_n3763));
  xor_4  g03387(.A(new_n3763), .B(new_n3758), .Y(new_n3764));
  nand_5 g03388(.A(pi192), .B(pi132), .Y(new_n3765));
  xor_4  g03389(.A(new_n3765), .B(new_n3764), .Y(new_n3766));
  xor_4  g03390(.A(new_n3766), .B(new_n3659), .Y(new_n3767));
  xor_4  g03391(.A(new_n3767), .B(new_n3648), .Y(new_n3768));
  xor_4  g03392(.A(new_n3768), .B(new_n3645), .Y(new_n3769));
  nand_5 g03393(.A(pi219), .B(pi074), .Y(new_n3770));
  nand_5 g03394(.A(pi239), .B(pi071), .Y(new_n3771));
  xor_4  g03395(.A(new_n3771), .B(new_n3770), .Y(new_n3772));
  nand_5 g03396(.A(pi087), .B(pi074), .Y(new_n3773));
  nand_5 g03397(.A(pi253), .B(pi219), .Y(new_n3774));
  nand_5 g03398(.A(new_n3774), .B(new_n3773), .Y(new_n3775));
  nand_5 g03399(.A(pi102), .B(pi050), .Y(new_n3776));
  xor_4  g03400(.A(new_n3774), .B(new_n3773), .Y(new_n3777));
  nand_5 g03401(.A(new_n3777), .B(new_n3776), .Y(new_n3778));
  nand_5 g03402(.A(new_n3778), .B(new_n3775), .Y(new_n3779));
  nand_5 g03403(.A(pi205), .B(pi087), .Y(new_n3780));
  xor_4  g03404(.A(new_n3780), .B(new_n3779), .Y(new_n3781));
  nand_5 g03405(.A(pi207), .B(pi023), .Y(new_n3782));
  nand_5 g03406(.A(pi226), .B(pi155), .Y(new_n3783));
  nand_5 g03407(.A(new_n3783), .B(new_n3782), .Y(new_n3784));
  xor_4  g03408(.A(new_n3783), .B(new_n3782), .Y(new_n3785));
  nand_5 g03409(.A(pi099), .B(pi066), .Y(new_n3786));
  nand_5 g03410(.A(new_n3786), .B(new_n3785), .Y(new_n3787));
  nand_5 g03411(.A(new_n3787), .B(new_n3784), .Y(new_n3788));
  xor_4  g03412(.A(new_n3788), .B(new_n3781), .Y(new_n3789));
  xor_4  g03413(.A(new_n3789), .B(new_n3772), .Y(new_n3790));
  nand_5 g03414(.A(pi226), .B(pi023), .Y(new_n3791));
  nand_5 g03415(.A(pi207), .B(pi099), .Y(new_n3792));
  nand_5 g03416(.A(new_n3792), .B(new_n3791), .Y(new_n3793));
  nand_5 g03417(.A(pi226), .B(pi099), .Y(new_n3794));
  nor_5  g03418(.A(new_n3794), .B(new_n3782), .Y(new_n3795));
  not_8  g03419(.A(new_n3795), .Y(new_n3796));
  nand_5 g03420(.A(new_n3796), .B(new_n3793), .Y(new_n3797));
  nand_5 g03421(.A(pi123), .B(pi066), .Y(new_n3798));
  nand_5 g03422(.A(new_n3798), .B(new_n3797), .Y(new_n3799));
  nand_5 g03423(.A(pi169), .B(pi066), .Y(new_n3800));
  nand_5 g03424(.A(new_n3800), .B(new_n3794), .Y(new_n3801));
  xor_4  g03425(.A(new_n3800), .B(new_n3794), .Y(new_n3802));
  nand_5 g03426(.A(pi207), .B(pi123), .Y(new_n3803));
  nand_5 g03427(.A(new_n3803), .B(new_n3802), .Y(new_n3804));
  nand_5 g03428(.A(new_n3804), .B(new_n3801), .Y(new_n3805));
  xor_4  g03429(.A(new_n3798), .B(new_n3797), .Y(new_n3806));
  nand_5 g03430(.A(new_n3806), .B(new_n3805), .Y(new_n3807));
  nand_5 g03431(.A(new_n3807), .B(new_n3799), .Y(new_n3808));
  xor_4  g03432(.A(new_n3639), .B(new_n3638), .Y(new_n3809));
  nand_5 g03433(.A(new_n3809), .B(new_n3808), .Y(new_n3810));
  xor_4  g03434(.A(new_n3786), .B(new_n3785), .Y(new_n3811));
  nand_5 g03435(.A(pi123), .B(pi055), .Y(new_n3812));
  xor_4  g03436(.A(new_n3812), .B(new_n3795), .Y(new_n3813));
  xor_4  g03437(.A(new_n3813), .B(new_n3811), .Y(new_n3814));
  not_8  g03438(.A(new_n3814), .Y(new_n3815));
  xor_4  g03439(.A(new_n3809), .B(new_n3808), .Y(new_n3816));
  nand_5 g03440(.A(new_n3816), .B(new_n3815), .Y(new_n3817));
  nand_5 g03441(.A(new_n3817), .B(new_n3810), .Y(new_n3818));
  nand_5 g03442(.A(pi230), .B(pi122), .Y(new_n3819));
  xor_4  g03443(.A(new_n3819), .B(new_n3818), .Y(new_n3820));
  xor_4  g03444(.A(new_n3820), .B(new_n3790), .Y(new_n3821));
  nand_5 g03445(.A(pi138), .B(pi037), .Y(new_n3822));
  nand_5 g03446(.A(pi251), .B(pi186), .Y(new_n3823));
  nand_5 g03447(.A(pi109), .B(pi094), .Y(new_n3824));
  xor_4  g03448(.A(new_n3824), .B(new_n3823), .Y(new_n3825));
  xor_4  g03449(.A(new_n3825), .B(new_n3822), .Y(new_n3826));
  nand_5 g03450(.A(pi150), .B(pi101), .Y(new_n3827));
  nand_5 g03451(.A(pi177), .B(pi069), .Y(new_n3828));
  xor_4  g03452(.A(new_n3828), .B(new_n3827), .Y(new_n3829));
  nand_5 g03453(.A(pi142), .B(pi002), .Y(new_n3830));
  nand_5 g03454(.A(pi142), .B(pi055), .Y(new_n3831));
  nand_5 g03455(.A(pi142), .B(pi066), .Y(new_n3832));
  nand_5 g03456(.A(pi207), .B(pi071), .Y(new_n3833));
  nand_5 g03457(.A(new_n3833), .B(new_n3832), .Y(new_n3834));
  nand_5 g03458(.A(pi226), .B(pi169), .Y(new_n3835));
  xor_4  g03459(.A(new_n3833), .B(new_n3832), .Y(new_n3836));
  nand_5 g03460(.A(new_n3836), .B(new_n3835), .Y(new_n3837));
  nand_5 g03461(.A(new_n3837), .B(new_n3834), .Y(new_n3838));
  nor_5  g03462(.A(new_n3838), .B(new_n3831), .Y(new_n3839));
  xor_4  g03463(.A(new_n3838), .B(new_n3831), .Y(new_n3840));
  nand_5 g03464(.A(pi207), .B(pi169), .Y(new_n3841));
  nand_5 g03465(.A(pi071), .B(pi066), .Y(new_n3842));
  nand_5 g03466(.A(pi226), .B(pi123), .Y(new_n3843));
  xor_4  g03467(.A(new_n3843), .B(new_n3842), .Y(new_n3844));
  xor_4  g03468(.A(new_n3844), .B(new_n3841), .Y(new_n3845));
  not_8  g03469(.A(new_n3845), .Y(new_n3846));
  and_6  g03470(.A(new_n3846), .B(new_n3840), .Y(new_n3847));
  nor_5  g03471(.A(new_n3847), .B(new_n3839), .Y(new_n3848));
  nor_5  g03472(.A(new_n3848), .B(new_n3830), .Y(new_n3849));
  xor_4  g03473(.A(new_n3803), .B(new_n3802), .Y(new_n3850));
  nand_5 g03474(.A(pi071), .B(pi055), .Y(new_n3851));
  nand_5 g03475(.A(new_n3843), .B(new_n3842), .Y(new_n3852));
  nand_5 g03476(.A(new_n3844), .B(new_n3841), .Y(new_n3853));
  nand_5 g03477(.A(new_n3853), .B(new_n3852), .Y(new_n3854));
  xor_4  g03478(.A(new_n3854), .B(new_n3851), .Y(new_n3855));
  xor_4  g03479(.A(new_n3855), .B(new_n3850), .Y(new_n3856));
  xnor_4 g03480(.A(new_n3848), .B(new_n3830), .Y(new_n3857));
  nor_5  g03481(.A(new_n3857), .B(new_n3856), .Y(new_n3858));
  nor_5  g03482(.A(new_n3858), .B(new_n3849), .Y(new_n3859));
  xor_4  g03483(.A(new_n3806), .B(new_n3805), .Y(new_n3860));
  nand_5 g03484(.A(new_n3854), .B(new_n3851), .Y(new_n3861));
  not_8  g03485(.A(new_n3861), .Y(new_n3862));
  and_6  g03486(.A(new_n3855), .B(new_n3850), .Y(new_n3863));
  nor_5  g03487(.A(new_n3863), .B(new_n3862), .Y(new_n3864));
  nand_5 g03488(.A(pi071), .B(pi002), .Y(new_n3865));
  nand_5 g03489(.A(pi169), .B(pi055), .Y(new_n3866));
  nand_5 g03490(.A(new_n3866), .B(new_n3865), .Y(new_n3867));
  nor_5  g03491(.A(new_n3851), .B(new_n3638), .Y(new_n3868));
  not_8  g03492(.A(new_n3868), .Y(new_n3869));
  nand_5 g03493(.A(new_n3869), .B(new_n3867), .Y(new_n3870));
  xor_4  g03494(.A(new_n3870), .B(new_n3864), .Y(new_n3871));
  xor_4  g03495(.A(new_n3871), .B(new_n3860), .Y(new_n3872));
  not_8  g03496(.A(new_n3872), .Y(new_n3873));
  nor_5  g03497(.A(new_n3873), .B(new_n3859), .Y(new_n3874));
  not_8  g03498(.A(new_n3874), .Y(new_n3875));
  xor_4  g03499(.A(new_n3816), .B(new_n3814), .Y(new_n3876));
  not_8  g03500(.A(new_n3864), .Y(new_n3877));
  nand_5 g03501(.A(new_n3870), .B(new_n3877), .Y(new_n3878));
  not_8  g03502(.A(new_n3871), .Y(new_n3879));
  nand_5 g03503(.A(new_n3879), .B(new_n3860), .Y(new_n3880));
  nand_5 g03504(.A(new_n3880), .B(new_n3878), .Y(new_n3881));
  xor_4  g03505(.A(new_n3881), .B(new_n3868), .Y(new_n3882));
  xor_4  g03506(.A(new_n3882), .B(new_n3876), .Y(new_n3883));
  nor_5  g03507(.A(new_n3883), .B(new_n3875), .Y(new_n3884));
  nand_5 g03508(.A(pi142), .B(pi025), .Y(new_n3885));
  xor_4  g03509(.A(new_n3872), .B(new_n3859), .Y(new_n3886));
  nor_5  g03510(.A(new_n3886), .B(new_n3885), .Y(new_n3887));
  xor_4  g03511(.A(new_n3845), .B(new_n3840), .Y(new_n3888));
  xnor_4 g03512(.A(new_n3836), .B(new_n3835), .Y(new_n3889));
  nand_5 g03513(.A(pi207), .B(pi142), .Y(new_n3890));
  nand_5 g03514(.A(pi226), .B(pi071), .Y(new_n3891));
  nor_5  g03515(.A(new_n3891), .B(new_n3890), .Y(new_n3892));
  nand_5 g03516(.A(new_n3892), .B(new_n3889), .Y(new_n3893));
  nor_5  g03517(.A(new_n3893), .B(new_n3888), .Y(new_n3894));
  xor_4  g03518(.A(new_n3857), .B(new_n3856), .Y(new_n3895));
  nand_5 g03519(.A(new_n3895), .B(new_n3894), .Y(new_n3896));
  not_8  g03520(.A(new_n3896), .Y(new_n3897));
  xor_4  g03521(.A(new_n3886), .B(new_n3885), .Y(new_n3898));
  and_6  g03522(.A(new_n3898), .B(new_n3897), .Y(new_n3899));
  nor_5  g03523(.A(new_n3899), .B(new_n3887), .Y(new_n3900));
  xor_4  g03524(.A(new_n3883), .B(new_n3874), .Y(new_n3901));
  nor_5  g03525(.A(new_n3901), .B(new_n3900), .Y(new_n3902));
  nor_5  g03526(.A(new_n3902), .B(new_n3884), .Y(new_n3903));
  nand_5 g03527(.A(pi253), .B(pi102), .Y(new_n3904));
  nor_5  g03528(.A(new_n3605), .B(new_n3586), .Y(new_n3905));
  nor_5  g03529(.A(new_n3606), .B(new_n3604), .Y(new_n3906));
  nor_5  g03530(.A(new_n3906), .B(new_n3905), .Y(new_n3907));
  xor_4  g03531(.A(new_n3907), .B(new_n3904), .Y(new_n3908));
  xor_4  g03532(.A(new_n3908), .B(new_n3903), .Y(new_n3909));
  nor_5  g03533(.A(new_n3720), .B(new_n3719), .Y(new_n3910));
  nor_5  g03534(.A(new_n3726), .B(new_n3722), .Y(new_n3911));
  nor_5  g03535(.A(new_n3911), .B(new_n3910), .Y(new_n3912));
  nand_5 g03536(.A(pi184), .B(pi020), .Y(new_n3913));
  xor_4  g03537(.A(new_n3913), .B(new_n3912), .Y(new_n3914));
  xor_4  g03538(.A(new_n3914), .B(new_n3909), .Y(new_n3915));
  xor_4  g03539(.A(new_n3915), .B(new_n3829), .Y(new_n3916));
  xnor_4 g03540(.A(new_n3901), .B(new_n3900), .Y(new_n3917));
  nand_5 g03541(.A(pi253), .B(pi087), .Y(new_n3918));
  nand_5 g03542(.A(pi219), .B(pi014), .Y(new_n3919));
  nand_5 g03543(.A(pi173), .B(pi087), .Y(new_n3920));
  nand_5 g03544(.A(pi109), .B(pi102), .Y(new_n3921));
  nor_5  g03545(.A(new_n3921), .B(new_n3920), .Y(new_n3922));
  nand_5 g03546(.A(new_n3921), .B(new_n3920), .Y(new_n3923));
  and_6  g03547(.A(pi109), .B(pi087), .Y(new_n3924));
  nor_5  g03548(.A(new_n3924), .B(new_n3919), .Y(new_n3925));
  nor_5  g03549(.A(new_n3925), .B(new_n3923), .Y(new_n3926));
  nor_5  g03550(.A(new_n3926), .B(new_n3922), .Y(new_n3927));
  nor_5  g03551(.A(new_n3927), .B(new_n3919), .Y(new_n3928));
  nand_5 g03552(.A(pi109), .B(pi001), .Y(new_n3929));
  nand_5 g03553(.A(pi219), .B(pi173), .Y(new_n3930));
  nand_5 g03554(.A(pi102), .B(pi014), .Y(new_n3931));
  xor_4  g03555(.A(new_n3931), .B(new_n3930), .Y(new_n3932));
  xor_4  g03556(.A(new_n3932), .B(new_n3929), .Y(new_n3933));
  not_8  g03557(.A(new_n3933), .Y(new_n3934));
  not_8  g03558(.A(new_n3919), .Y(new_n3935));
  or_6   g03559(.A(new_n3922), .B(new_n3935), .Y(new_n3936));
  nand_5 g03560(.A(new_n3936), .B(new_n3923), .Y(new_n3937));
  nand_5 g03561(.A(pi230), .B(pi087), .Y(new_n3938));
  xor_4  g03562(.A(new_n3938), .B(new_n3937), .Y(new_n3939));
  xor_4  g03563(.A(new_n3939), .B(new_n3934), .Y(new_n3940));
  nand_5 g03564(.A(new_n3940), .B(new_n3928), .Y(new_n3941));
  nand_5 g03565(.A(pi087), .B(pi050), .Y(new_n3942));
  nor_5  g03566(.A(new_n3938), .B(new_n3937), .Y(new_n3943));
  and_6  g03567(.A(new_n3939), .B(new_n3934), .Y(new_n3944));
  nor_5  g03568(.A(new_n3944), .B(new_n3943), .Y(new_n3945));
  xor_4  g03569(.A(new_n3945), .B(new_n3942), .Y(new_n3946));
  nand_5 g03570(.A(pi173), .B(pi102), .Y(new_n3947));
  nand_5 g03571(.A(pi014), .B(pi001), .Y(new_n3948));
  xor_4  g03572(.A(new_n3948), .B(new_n3620), .Y(new_n3949));
  xor_4  g03573(.A(new_n3949), .B(new_n3947), .Y(new_n3950));
  nand_5 g03574(.A(pi230), .B(pi219), .Y(new_n3951));
  nand_5 g03575(.A(new_n3931), .B(new_n3930), .Y(new_n3952));
  nand_5 g03576(.A(new_n3932), .B(new_n3929), .Y(new_n3953));
  nand_5 g03577(.A(new_n3953), .B(new_n3952), .Y(new_n3954));
  xor_4  g03578(.A(new_n3954), .B(new_n3951), .Y(new_n3955));
  xnor_4 g03579(.A(new_n3955), .B(new_n3950), .Y(new_n3956));
  xnor_4 g03580(.A(new_n3956), .B(new_n3946), .Y(new_n3957));
  or_6   g03581(.A(new_n3957), .B(new_n3941), .Y(new_n3958));
  nand_5 g03582(.A(new_n3958), .B(new_n3918), .Y(new_n3959));
  xor_4  g03583(.A(new_n3958), .B(new_n3918), .Y(new_n3960));
  not_8  g03584(.A(new_n3960), .Y(new_n3961));
  nand_5 g03585(.A(new_n3954), .B(new_n3951), .Y(new_n3962));
  nand_5 g03586(.A(new_n3955), .B(new_n3950), .Y(new_n3963));
  nand_5 g03587(.A(new_n3963), .B(new_n3962), .Y(new_n3964));
  nand_5 g03588(.A(pi230), .B(pi102), .Y(new_n3965));
  nand_5 g03589(.A(pi219), .B(pi050), .Y(new_n3966));
  nand_5 g03590(.A(new_n3966), .B(new_n3965), .Y(new_n3967));
  nor_5  g03591(.A(new_n3951), .B(new_n3776), .Y(new_n3968));
  not_8  g03592(.A(new_n3968), .Y(new_n3969));
  nand_5 g03593(.A(new_n3969), .B(new_n3967), .Y(new_n3970));
  nand_5 g03594(.A(pi122), .B(pi014), .Y(new_n3971));
  nand_5 g03595(.A(pi135), .B(pi109), .Y(new_n3972));
  nand_5 g03596(.A(new_n3972), .B(new_n3971), .Y(new_n3973));
  nand_5 g03597(.A(new_n3973), .B(new_n3622), .Y(new_n3974));
  nand_5 g03598(.A(pi173), .B(pi001), .Y(new_n3975));
  nand_5 g03599(.A(new_n3948), .B(new_n3620), .Y(new_n3976));
  nand_5 g03600(.A(new_n3949), .B(new_n3947), .Y(new_n3977));
  nand_5 g03601(.A(new_n3977), .B(new_n3976), .Y(new_n3978));
  xor_4  g03602(.A(new_n3978), .B(new_n3975), .Y(new_n3979));
  xor_4  g03603(.A(new_n3979), .B(new_n3974), .Y(new_n3980));
  xnor_4 g03604(.A(new_n3980), .B(new_n3970), .Y(new_n3981));
  xor_4  g03605(.A(new_n3981), .B(new_n3964), .Y(new_n3982));
  not_8  g03606(.A(new_n3982), .Y(new_n3983));
  nor_5  g03607(.A(new_n3945), .B(new_n3942), .Y(new_n3984));
  and_6  g03608(.A(new_n3956), .B(new_n3946), .Y(new_n3985));
  nor_5  g03609(.A(new_n3985), .B(new_n3984), .Y(new_n3986));
  xor_4  g03610(.A(new_n3986), .B(new_n3983), .Y(new_n3987));
  or_6   g03611(.A(new_n3987), .B(new_n3961), .Y(new_n3988));
  nand_5 g03612(.A(new_n3988), .B(new_n3959), .Y(new_n3989));
  nor_5  g03613(.A(new_n3986), .B(new_n3983), .Y(new_n3990));
  nor_5  g03614(.A(new_n3980), .B(new_n3970), .Y(new_n3991));
  nor_5  g03615(.A(new_n3981), .B(new_n3964), .Y(new_n3992));
  xor_4  g03616(.A(new_n3992), .B(new_n3969), .Y(new_n3993));
  not_8  g03617(.A(new_n3993), .Y(new_n3994));
  nor_5  g03618(.A(new_n3994), .B(new_n3991), .Y(new_n3995));
  nand_5 g03619(.A(new_n3978), .B(new_n3975), .Y(new_n3996));
  nand_5 g03620(.A(new_n3979), .B(new_n3974), .Y(new_n3997));
  nand_5 g03621(.A(new_n3997), .B(new_n3996), .Y(new_n3998));
  xor_4  g03622(.A(new_n3777), .B(new_n3776), .Y(new_n3999));
  xor_4  g03623(.A(new_n3999), .B(new_n3998), .Y(new_n4000));
  xor_4  g03624(.A(new_n3629), .B(new_n3625), .Y(new_n4001));
  xor_4  g03625(.A(new_n4001), .B(new_n4000), .Y(new_n4002));
  xor_4  g03626(.A(new_n4002), .B(new_n3995), .Y(new_n4003));
  xor_4  g03627(.A(new_n4003), .B(new_n3990), .Y(new_n4004));
  xor_4  g03628(.A(new_n4004), .B(new_n3989), .Y(new_n4005));
  or_6   g03629(.A(new_n4005), .B(new_n3917), .Y(new_n4006));
  xor_4  g03630(.A(new_n3898), .B(new_n3897), .Y(new_n4007));
  xor_4  g03631(.A(new_n3987), .B(new_n3960), .Y(new_n4008));
  nand_5 g03632(.A(new_n4008), .B(new_n4007), .Y(new_n4009));
  xor_4  g03633(.A(new_n3893), .B(new_n3888), .Y(new_n4010));
  nand_5 g03634(.A(pi109), .B(pi087), .Y(new_n4011));
  nand_5 g03635(.A(pi226), .B(pi142), .Y(new_n4012));
  nor_5  g03636(.A(new_n4012), .B(new_n4011), .Y(new_n4013));
  xor_4  g03637(.A(new_n3891), .B(new_n3890), .Y(new_n4014));
  nor_5  g03638(.A(new_n4014), .B(new_n4013), .Y(new_n4015));
  nand_5 g03639(.A(pi219), .B(pi109), .Y(new_n4016));
  nand_5 g03640(.A(pi087), .B(pi014), .Y(new_n4017));
  xor_4  g03641(.A(new_n4017), .B(new_n4016), .Y(new_n4018));
  xnor_4 g03642(.A(new_n4014), .B(new_n4013), .Y(new_n4019));
  nor_5  g03643(.A(new_n4019), .B(new_n4018), .Y(new_n4020));
  nor_5  g03644(.A(new_n4020), .B(new_n4015), .Y(new_n4021));
  nand_5 g03645(.A(new_n3925), .B(new_n3923), .Y(new_n4022));
  nand_5 g03646(.A(new_n4022), .B(new_n3927), .Y(new_n4023));
  not_8  g03647(.A(new_n4023), .Y(new_n4024));
  nor_5  g03648(.A(new_n4024), .B(new_n4021), .Y(new_n4025));
  xor_4  g03649(.A(new_n3892), .B(new_n3889), .Y(new_n4026));
  xor_4  g03650(.A(new_n4023), .B(new_n4021), .Y(new_n4027));
  nor_5  g03651(.A(new_n4027), .B(new_n4026), .Y(new_n4028));
  nor_5  g03652(.A(new_n4028), .B(new_n4025), .Y(new_n4029));
  nor_5  g03653(.A(new_n4029), .B(new_n4010), .Y(new_n4030));
  xor_4  g03654(.A(new_n3940), .B(new_n3928), .Y(new_n4031));
  xnor_4 g03655(.A(new_n4029), .B(new_n4010), .Y(new_n4032));
  nor_5  g03656(.A(new_n4032), .B(new_n4031), .Y(new_n4033));
  nor_5  g03657(.A(new_n4033), .B(new_n4030), .Y(new_n4034));
  xor_4  g03658(.A(new_n3957), .B(new_n3941), .Y(new_n4035));
  or_6   g03659(.A(new_n4035), .B(new_n4034), .Y(new_n4036));
  xnor_4 g03660(.A(new_n3895), .B(new_n3894), .Y(new_n4037));
  xor_4  g03661(.A(new_n4035), .B(new_n4034), .Y(new_n4038));
  nand_5 g03662(.A(new_n4038), .B(new_n4037), .Y(new_n4039));
  nand_5 g03663(.A(new_n4039), .B(new_n4036), .Y(new_n4040));
  xnor_4 g03664(.A(new_n4008), .B(new_n4007), .Y(new_n4041));
  or_6   g03665(.A(new_n4041), .B(new_n4040), .Y(new_n4042));
  nand_5 g03666(.A(new_n4042), .B(new_n4009), .Y(new_n4043));
  xor_4  g03667(.A(new_n4005), .B(new_n3917), .Y(new_n4044));
  nand_5 g03668(.A(new_n4044), .B(new_n4043), .Y(new_n4045));
  nand_5 g03669(.A(new_n4045), .B(new_n4006), .Y(new_n4046));
  nor_5  g03670(.A(new_n3723), .B(new_n3709), .Y(new_n4047));
  nor_5  g03671(.A(new_n3725), .B(new_n3724), .Y(new_n4048));
  nor_5  g03672(.A(new_n4048), .B(new_n4047), .Y(new_n4049));
  nand_5 g03673(.A(new_n3881), .B(new_n3869), .Y(new_n4050));
  or_6   g03674(.A(new_n3882), .B(new_n3876), .Y(new_n4051));
  nand_5 g03675(.A(new_n4051), .B(new_n4050), .Y(new_n4052));
  xor_4  g03676(.A(new_n4052), .B(new_n4049), .Y(new_n4053));
  nand_5 g03677(.A(pi244), .B(pi225), .Y(new_n4054));
  xor_4  g03678(.A(new_n4054), .B(new_n4053), .Y(new_n4055));
  xor_4  g03679(.A(new_n4055), .B(new_n4046), .Y(new_n4056));
  xor_4  g03680(.A(new_n4056), .B(new_n3916), .Y(new_n4057));
  xor_4  g03681(.A(new_n4057), .B(new_n3826), .Y(new_n4058));
  xor_4  g03682(.A(new_n4058), .B(new_n3821), .Y(new_n4059));
  xor_4  g03683(.A(new_n4059), .B(new_n3769), .Y(new_n4060));
  xor_4  g03684(.A(new_n3752), .B(new_n3745), .Y(new_n4061));
  xor_4  g03685(.A(new_n4032), .B(new_n4031), .Y(new_n4062));
  xor_4  g03686(.A(new_n3750), .B(new_n3746), .Y(new_n4063));
  and_6  g03687(.A(new_n4063), .B(new_n4062), .Y(new_n4064));
  xor_4  g03688(.A(new_n4012), .B(new_n3924), .Y(new_n4065));
  or_6   g03689(.A(new_n4065), .B(new_n3748), .Y(new_n4066));
  nand_5 g03690(.A(pi186), .B(pi138), .Y(new_n4067));
  nand_5 g03691(.A(pi182), .B(pi132), .Y(new_n4068));
  nand_5 g03692(.A(new_n4068), .B(new_n4067), .Y(new_n4069));
  nand_5 g03693(.A(new_n4069), .B(new_n3749), .Y(new_n4070));
  nor_5  g03694(.A(new_n4070), .B(new_n4066), .Y(new_n4071));
  xor_4  g03695(.A(new_n4019), .B(new_n4018), .Y(new_n4072));
  xnor_4 g03696(.A(new_n4070), .B(new_n4066), .Y(new_n4073));
  nor_5  g03697(.A(new_n4073), .B(new_n4072), .Y(new_n4074));
  nor_5  g03698(.A(new_n4074), .B(new_n4071), .Y(new_n4075));
  xnor_4 g03699(.A(new_n3749), .B(new_n3747), .Y(new_n4076));
  or_6   g03700(.A(new_n4076), .B(new_n4075), .Y(new_n4077));
  xnor_4 g03701(.A(new_n4076), .B(new_n4075), .Y(new_n4078));
  xor_4  g03702(.A(new_n4027), .B(new_n4026), .Y(new_n4079));
  or_6   g03703(.A(new_n4079), .B(new_n4078), .Y(new_n4080));
  nand_5 g03704(.A(new_n4080), .B(new_n4077), .Y(new_n4081));
  not_8  g03705(.A(new_n4081), .Y(new_n4082));
  xor_4  g03706(.A(new_n4063), .B(new_n4062), .Y(new_n4083));
  and_6  g03707(.A(new_n4083), .B(new_n4082), .Y(new_n4084));
  nor_5  g03708(.A(new_n4084), .B(new_n4064), .Y(new_n4085));
  nand_5 g03709(.A(new_n4085), .B(new_n4061), .Y(new_n4086));
  xor_4  g03710(.A(new_n4085), .B(new_n4061), .Y(new_n4087));
  xnor_4 g03711(.A(new_n4038), .B(new_n4037), .Y(new_n4088));
  nand_5 g03712(.A(new_n4088), .B(new_n4087), .Y(new_n4089));
  and_6  g03713(.A(new_n4089), .B(new_n4086), .Y(new_n4090));
  xnor_4 g03714(.A(new_n3754), .B(new_n3753), .Y(new_n4091));
  nor_5  g03715(.A(new_n4091), .B(new_n4090), .Y(new_n4092));
  xnor_4 g03716(.A(new_n4041), .B(new_n4040), .Y(new_n4093));
  xnor_4 g03717(.A(new_n4091), .B(new_n4090), .Y(new_n4094));
  nor_5  g03718(.A(new_n4094), .B(new_n4093), .Y(new_n4095));
  nor_5  g03719(.A(new_n4095), .B(new_n4092), .Y(new_n4096));
  xor_4  g03720(.A(new_n3756), .B(new_n3739), .Y(new_n4097));
  nand_5 g03721(.A(new_n4097), .B(new_n4096), .Y(new_n4098));
  xnor_4 g03722(.A(new_n4044), .B(new_n4043), .Y(new_n4099));
  xor_4  g03723(.A(new_n4097), .B(new_n4096), .Y(new_n4100));
  nand_5 g03724(.A(new_n4100), .B(new_n4099), .Y(new_n4101));
  nand_5 g03725(.A(new_n4101), .B(new_n4098), .Y(new_n4102));
  nand_5 g03726(.A(new_n3992), .B(new_n3968), .Y(new_n4103));
  or_6   g03727(.A(new_n4002), .B(new_n3995), .Y(new_n4104));
  nand_5 g03728(.A(new_n4104), .B(new_n4103), .Y(new_n4105));
  xor_4  g03729(.A(new_n4105), .B(new_n4102), .Y(new_n4106));
  nand_5 g03730(.A(pi099), .B(pi055), .Y(new_n4107));
  nand_5 g03731(.A(pi050), .B(pi001), .Y(new_n4108));
  xor_4  g03732(.A(new_n4108), .B(new_n4107), .Y(new_n4109));
  nand_5 g03733(.A(new_n3577), .B(new_n3576), .Y(new_n4110));
  nand_5 g03734(.A(new_n3578), .B(new_n3575), .Y(new_n4111));
  nand_5 g03735(.A(new_n4111), .B(new_n4110), .Y(new_n4112));
  xor_4  g03736(.A(new_n4112), .B(new_n4109), .Y(new_n4113));
  nand_5 g03737(.A(pi160), .B(pi010), .Y(new_n4114));
  nand_5 g03738(.A(pi223), .B(pi221), .Y(new_n4115));
  or_6   g03739(.A(new_n3736), .B(new_n3727), .Y(new_n4116));
  nand_5 g03740(.A(new_n4116), .B(new_n3735), .Y(new_n4117));
  xor_4  g03741(.A(new_n4117), .B(new_n4115), .Y(new_n4118));
  nand_5 g03742(.A(new_n4003), .B(new_n3990), .Y(new_n4119));
  not_8  g03743(.A(new_n4004), .Y(new_n4120));
  or_6   g03744(.A(new_n4120), .B(new_n3989), .Y(new_n4121));
  nand_5 g03745(.A(new_n4121), .B(new_n4119), .Y(new_n4122));
  nand_5 g03746(.A(pi123), .B(pi002), .Y(new_n4123));
  xor_4  g03747(.A(new_n4123), .B(new_n4122), .Y(new_n4124));
  nor_5  g03748(.A(new_n3999), .B(new_n3998), .Y(new_n4125));
  not_8  g03749(.A(new_n4000), .Y(new_n4126));
  nor_5  g03750(.A(new_n4001), .B(new_n4126), .Y(new_n4127));
  or_6   g03751(.A(new_n4127), .B(new_n4125), .Y(new_n4128));
  nor_5  g03752(.A(new_n3812), .B(new_n3796), .Y(new_n4129));
  nor_5  g03753(.A(new_n3813), .B(new_n3811), .Y(new_n4130));
  nor_5  g03754(.A(new_n4130), .B(new_n4129), .Y(new_n4131));
  xor_4  g03755(.A(new_n4131), .B(new_n4128), .Y(new_n4132));
  xor_4  g03756(.A(new_n4132), .B(new_n4124), .Y(new_n4133));
  xor_4  g03757(.A(new_n4133), .B(new_n4118), .Y(new_n4134));
  xor_4  g03758(.A(new_n4134), .B(new_n4114), .Y(new_n4135));
  xor_4  g03759(.A(new_n4135), .B(new_n4113), .Y(new_n4136));
  xor_4  g03760(.A(new_n4136), .B(new_n4106), .Y(new_n4137));
  nand_5 g03761(.A(pi150), .B(pi020), .Y(new_n4138));
  nand_5 g03762(.A(pi223), .B(pi029), .Y(new_n4139));
  nand_5 g03763(.A(pi244), .B(pi020), .Y(new_n4140));
  nand_5 g03764(.A(new_n4140), .B(new_n4139), .Y(new_n4141));
  nand_5 g03765(.A(pi069), .B(pi060), .Y(new_n4142));
  xor_4  g03766(.A(new_n4140), .B(new_n4139), .Y(new_n4143));
  nand_5 g03767(.A(new_n4143), .B(new_n4142), .Y(new_n4144));
  nand_5 g03768(.A(new_n4144), .B(new_n4141), .Y(new_n4145));
  nand_5 g03769(.A(new_n4145), .B(new_n4138), .Y(new_n4146));
  xor_4  g03770(.A(new_n3593), .B(new_n3592), .Y(new_n4147));
  xor_4  g03771(.A(new_n4145), .B(new_n4138), .Y(new_n4148));
  nand_5 g03772(.A(new_n4148), .B(new_n4147), .Y(new_n4149));
  nand_5 g03773(.A(new_n4149), .B(new_n4146), .Y(new_n4150));
  nor_5  g03774(.A(new_n4138), .B(new_n3575), .Y(new_n4151));
  nand_5 g03775(.A(pi150), .B(pi060), .Y(new_n4152));
  nand_5 g03776(.A(pi221), .B(pi020), .Y(new_n4153));
  and_6  g03777(.A(new_n4153), .B(new_n4152), .Y(new_n4154));
  or_6   g03778(.A(new_n4154), .B(new_n4151), .Y(new_n4155));
  xor_4  g03779(.A(new_n3596), .B(new_n3595), .Y(new_n4156));
  xor_4  g03780(.A(new_n4156), .B(new_n4155), .Y(new_n4157));
  xor_4  g03781(.A(new_n4157), .B(new_n4150), .Y(new_n4158));
  nand_5 g03782(.A(pi221), .B(pi160), .Y(new_n4159));
  xor_4  g03783(.A(new_n4148), .B(new_n4147), .Y(new_n4160));
  nand_5 g03784(.A(new_n4160), .B(new_n4159), .Y(new_n4161));
  or_6   g03785(.A(new_n4160), .B(new_n4159), .Y(new_n4162));
  nand_5 g03786(.A(pi160), .B(pi150), .Y(new_n4163));
  nand_5 g03787(.A(pi244), .B(pi160), .Y(new_n4164));
  nand_5 g03788(.A(pi069), .B(pi020), .Y(new_n4165));
  nand_5 g03789(.A(new_n4165), .B(new_n4164), .Y(new_n4166));
  nand_5 g03790(.A(pi060), .B(pi029), .Y(new_n4167));
  xor_4  g03791(.A(new_n4165), .B(new_n4164), .Y(new_n4168));
  nand_5 g03792(.A(new_n4168), .B(new_n4167), .Y(new_n4169));
  nand_5 g03793(.A(new_n4169), .B(new_n4166), .Y(new_n4170));
  nand_5 g03794(.A(new_n4170), .B(new_n4163), .Y(new_n4171));
  xor_4  g03795(.A(new_n4143), .B(new_n4142), .Y(new_n4172));
  xor_4  g03796(.A(new_n4170), .B(new_n4163), .Y(new_n4173));
  nand_5 g03797(.A(new_n4173), .B(new_n4172), .Y(new_n4174));
  nand_5 g03798(.A(new_n4174), .B(new_n4171), .Y(new_n4175));
  nand_5 g03799(.A(new_n4175), .B(new_n4162), .Y(new_n4176));
  nand_5 g03800(.A(new_n4176), .B(new_n4161), .Y(new_n4177));
  nor_5  g03801(.A(new_n4177), .B(new_n4158), .Y(new_n4178));
  not_8  g03802(.A(new_n4178), .Y(new_n4179));
  not_8  g03803(.A(new_n4157), .Y(new_n4180));
  nor_5  g03804(.A(new_n4180), .B(new_n4150), .Y(new_n4181));
  nor_5  g03805(.A(new_n4156), .B(new_n4155), .Y(new_n4182));
  nor_5  g03806(.A(new_n4182), .B(new_n4151), .Y(new_n4183));
  not_8  g03807(.A(new_n4183), .Y(new_n4184));
  nor_5  g03808(.A(new_n4184), .B(new_n4181), .Y(new_n4185));
  and_6  g03809(.A(new_n4181), .B(new_n4151), .Y(new_n4186));
  or_6   g03810(.A(new_n4186), .B(new_n4185), .Y(new_n4187));
  xor_4  g03811(.A(new_n3607), .B(new_n3600), .Y(new_n4188));
  xor_4  g03812(.A(new_n4188), .B(new_n4187), .Y(new_n4189));
  nor_5  g03813(.A(new_n4189), .B(new_n4179), .Y(new_n4190));
  nand_5 g03814(.A(pi196), .B(pi160), .Y(new_n4191));
  xor_4  g03815(.A(new_n4168), .B(new_n4167), .Y(new_n4192));
  nand_5 g03816(.A(pi160), .B(pi029), .Y(new_n4193));
  or_6   g03817(.A(new_n4193), .B(new_n4165), .Y(new_n4194));
  or_6   g03818(.A(new_n4194), .B(new_n4192), .Y(new_n4195));
  not_8  g03819(.A(new_n4195), .Y(new_n4196));
  xor_4  g03820(.A(new_n4173), .B(new_n4172), .Y(new_n4197));
  not_8  g03821(.A(new_n4197), .Y(new_n4198));
  nand_5 g03822(.A(new_n4198), .B(new_n4196), .Y(new_n4199));
  not_8  g03823(.A(new_n4199), .Y(new_n4200));
  nand_5 g03824(.A(new_n4162), .B(new_n4161), .Y(new_n4201));
  xor_4  g03825(.A(new_n4201), .B(new_n4175), .Y(new_n4202));
  nand_5 g03826(.A(new_n4202), .B(new_n4200), .Y(new_n4203));
  nand_5 g03827(.A(new_n4203), .B(new_n4191), .Y(new_n4204));
  xor_4  g03828(.A(new_n4177), .B(new_n4158), .Y(new_n4205));
  not_8  g03829(.A(new_n4205), .Y(new_n4206));
  xor_4  g03830(.A(new_n4203), .B(new_n4191), .Y(new_n4207));
  nand_5 g03831(.A(new_n4207), .B(new_n4206), .Y(new_n4208));
  nand_5 g03832(.A(new_n4208), .B(new_n4204), .Y(new_n4209));
  xor_4  g03833(.A(new_n4189), .B(new_n4178), .Y(new_n4210));
  nor_5  g03834(.A(new_n4210), .B(new_n4209), .Y(new_n4211));
  or_6   g03835(.A(new_n4211), .B(new_n4190), .Y(new_n4212));
  xor_4  g03836(.A(new_n4210), .B(new_n4209), .Y(new_n4213));
  xor_4  g03837(.A(new_n4194), .B(new_n4192), .Y(new_n4214));
  xor_4  g03838(.A(new_n4079), .B(new_n4078), .Y(new_n4215));
  or_6   g03839(.A(new_n4215), .B(new_n4214), .Y(new_n4216));
  xnor_4 g03840(.A(new_n4065), .B(new_n3748), .Y(new_n4217));
  or_6   g03841(.A(new_n4217), .B(new_n4193), .Y(new_n4218));
  nand_5 g03842(.A(pi029), .B(pi020), .Y(new_n4219));
  nand_5 g03843(.A(pi160), .B(pi069), .Y(new_n4220));
  nand_5 g03844(.A(new_n4220), .B(new_n4219), .Y(new_n4221));
  nand_5 g03845(.A(new_n4221), .B(new_n4194), .Y(new_n4222));
  nand_5 g03846(.A(new_n4222), .B(new_n4218), .Y(new_n4223));
  xnor_4 g03847(.A(new_n4073), .B(new_n4072), .Y(new_n4224));
  xor_4  g03848(.A(new_n4222), .B(new_n4218), .Y(new_n4225));
  nand_5 g03849(.A(new_n4225), .B(new_n4224), .Y(new_n4226));
  nand_5 g03850(.A(new_n4226), .B(new_n4223), .Y(new_n4227));
  xor_4  g03851(.A(new_n4215), .B(new_n4214), .Y(new_n4228));
  nand_5 g03852(.A(new_n4228), .B(new_n4227), .Y(new_n4229));
  nand_5 g03853(.A(new_n4229), .B(new_n4216), .Y(new_n4230));
  xor_4  g03854(.A(new_n4197), .B(new_n4196), .Y(new_n4231));
  or_6   g03855(.A(new_n4231), .B(new_n4230), .Y(new_n4232));
  xor_4  g03856(.A(new_n4231), .B(new_n4230), .Y(new_n4233));
  xor_4  g03857(.A(new_n4083), .B(new_n4081), .Y(new_n4234));
  nand_5 g03858(.A(new_n4234), .B(new_n4233), .Y(new_n4235));
  nand_5 g03859(.A(new_n4235), .B(new_n4232), .Y(new_n4236));
  xor_4  g03860(.A(new_n4202), .B(new_n4199), .Y(new_n4237));
  not_8  g03861(.A(new_n4237), .Y(new_n4238));
  nor_5  g03862(.A(new_n4238), .B(new_n4236), .Y(new_n4239));
  xor_4  g03863(.A(new_n4088), .B(new_n4087), .Y(new_n4240));
  xor_4  g03864(.A(new_n4237), .B(new_n4236), .Y(new_n4241));
  nor_5  g03865(.A(new_n4241), .B(new_n4240), .Y(new_n4242));
  nor_5  g03866(.A(new_n4242), .B(new_n4239), .Y(new_n4243));
  xor_4  g03867(.A(new_n4207), .B(new_n4205), .Y(new_n4244));
  nand_5 g03868(.A(new_n4244), .B(new_n4243), .Y(new_n4245));
  xor_4  g03869(.A(new_n4244), .B(new_n4243), .Y(new_n4246));
  xor_4  g03870(.A(new_n4094), .B(new_n4093), .Y(new_n4247));
  nand_5 g03871(.A(new_n4247), .B(new_n4246), .Y(new_n4248));
  nand_5 g03872(.A(new_n4248), .B(new_n4245), .Y(new_n4249));
  nand_5 g03873(.A(new_n4249), .B(new_n4213), .Y(new_n4250));
  xor_4  g03874(.A(new_n4249), .B(new_n4213), .Y(new_n4251));
  xnor_4 g03875(.A(new_n4100), .B(new_n4099), .Y(new_n4252));
  nand_5 g03876(.A(new_n4252), .B(new_n4251), .Y(new_n4253));
  nand_5 g03877(.A(new_n4253), .B(new_n4250), .Y(new_n4254));
  xor_4  g03878(.A(new_n4254), .B(new_n4212), .Y(new_n4255));
  nor_5  g03879(.A(new_n4188), .B(new_n4187), .Y(new_n4256));
  nor_5  g03880(.A(new_n4256), .B(new_n4185), .Y(new_n4257));
  nand_5 g03881(.A(new_n3627), .B(new_n3626), .Y(new_n4258));
  nand_5 g03882(.A(new_n3628), .B(new_n3619), .Y(new_n4259));
  nand_5 g03883(.A(new_n4259), .B(new_n4258), .Y(new_n4260));
  nand_5 g03884(.A(pi195), .B(pi041), .Y(new_n4261));
  xor_4  g03885(.A(new_n4261), .B(new_n4260), .Y(new_n4262));
  xor_4  g03886(.A(new_n4262), .B(new_n4257), .Y(new_n4263));
  xor_4  g03887(.A(new_n4263), .B(new_n4255), .Y(new_n4264));
  xor_4  g03888(.A(new_n4264), .B(new_n4137), .Y(new_n4265));
  xor_4  g03889(.A(new_n4265), .B(new_n4060), .Y(new_n4266));
  xor_4  g03890(.A(new_n4266), .B(new_n3574), .Y(po013));
  or_6   g03891(.A(new_n977), .B(new_n930), .Y(new_n4268));
  nand_5 g03892(.A(new_n1011), .B(new_n978), .Y(new_n4269));
  nand_5 g03893(.A(new_n4269), .B(new_n4268), .Y(new_n4270));
  nand_5 g03894(.A(new_n929), .B(new_n918), .Y(new_n4271));
  nand_5 g03895(.A(pi237), .B(pi175), .Y(new_n4272));
  not_8  g03896(.A(new_n926), .Y(new_n4273));
  nor_5  g03897(.A(new_n927), .B(new_n4273), .Y(new_n4274));
  nor_5  g03898(.A(new_n928), .B(new_n923), .Y(new_n4275));
  nor_5  g03899(.A(new_n4275), .B(new_n4274), .Y(new_n4276));
  xor_4  g03900(.A(new_n4276), .B(new_n4272), .Y(new_n4277));
  nand_5 g03901(.A(pi167), .B(pi162), .Y(new_n4278));
  nand_5 g03902(.A(pi240), .B(pi179), .Y(new_n4279));
  nand_5 g03903(.A(pi149), .B(pi033), .Y(new_n4280));
  xor_4  g03904(.A(new_n4280), .B(new_n4279), .Y(new_n4281));
  xor_4  g03905(.A(new_n4281), .B(new_n4278), .Y(new_n4282));
  nand_5 g03906(.A(new_n921), .B(new_n920), .Y(new_n4283));
  nand_5 g03907(.A(new_n922), .B(new_n919), .Y(new_n4284));
  nand_5 g03908(.A(new_n4284), .B(new_n4283), .Y(new_n4285));
  nand_5 g03909(.A(pi134), .B(pi048), .Y(new_n4286));
  xor_4  g03910(.A(new_n4286), .B(new_n4285), .Y(new_n4287));
  xnor_4 g03911(.A(new_n4287), .B(new_n4282), .Y(new_n4288));
  xor_4  g03912(.A(new_n4288), .B(new_n4277), .Y(new_n4289));
  xor_4  g03913(.A(new_n4289), .B(new_n4271), .Y(new_n4290));
  or_6   g03914(.A(new_n4290), .B(new_n4270), .Y(new_n4291));
  nor_5  g03915(.A(new_n1008), .B(new_n997), .Y(new_n4292));
  nand_5 g03916(.A(pi163), .B(pi144), .Y(new_n4293));
  nand_5 g03917(.A(pi228), .B(pi061), .Y(new_n4294));
  nand_5 g03918(.A(pi178), .B(pi039), .Y(new_n4295));
  nand_5 g03919(.A(pi188), .B(pi116), .Y(new_n4296));
  xor_4  g03920(.A(new_n4296), .B(new_n4295), .Y(new_n4297));
  xor_4  g03921(.A(new_n4297), .B(new_n4294), .Y(new_n4298));
  nand_5 g03922(.A(new_n1000), .B(new_n999), .Y(new_n4299));
  nand_5 g03923(.A(new_n1001), .B(new_n998), .Y(new_n4300));
  nand_5 g03924(.A(new_n4300), .B(new_n4299), .Y(new_n4301));
  nand_5 g03925(.A(pi148), .B(pi012), .Y(new_n4302));
  xor_4  g03926(.A(new_n4302), .B(new_n4301), .Y(new_n4303));
  xor_4  g03927(.A(new_n4303), .B(new_n4298), .Y(new_n4304));
  xnor_4 g03928(.A(new_n4304), .B(new_n4293), .Y(new_n4305));
  nand_5 g03929(.A(new_n1006), .B(new_n1003), .Y(new_n4306));
  nand_5 g03930(.A(new_n1007), .B(new_n1002), .Y(new_n4307));
  nand_5 g03931(.A(new_n4307), .B(new_n4306), .Y(new_n4308));
  xor_4  g03932(.A(new_n4308), .B(new_n4305), .Y(new_n4309));
  xor_4  g03933(.A(new_n4309), .B(new_n4292), .Y(new_n4310));
  nand_5 g03934(.A(new_n1009), .B(new_n996), .Y(new_n4311));
  nand_5 g03935(.A(new_n1010), .B(new_n982), .Y(new_n4312));
  nand_5 g03936(.A(new_n4312), .B(new_n4311), .Y(new_n4313));
  nor_5  g03937(.A(new_n995), .B(new_n984), .Y(new_n4314));
  nand_5 g03938(.A(pi118), .B(pi107), .Y(new_n4315));
  nor_5  g03939(.A(new_n993), .B(new_n990), .Y(new_n4316));
  nor_5  g03940(.A(new_n994), .B(new_n989), .Y(new_n4317));
  nor_5  g03941(.A(new_n4317), .B(new_n4316), .Y(new_n4318));
  xor_4  g03942(.A(new_n4318), .B(new_n4315), .Y(new_n4319));
  nand_5 g03943(.A(pi108), .B(pi049), .Y(new_n4320));
  nand_5 g03944(.A(pi245), .B(pi042), .Y(new_n4321));
  nand_5 g03945(.A(pi201), .B(pi051), .Y(new_n4322));
  xor_4  g03946(.A(new_n4322), .B(new_n4321), .Y(new_n4323));
  xor_4  g03947(.A(new_n4323), .B(new_n4320), .Y(new_n4324));
  nand_5 g03948(.A(pi171), .B(pi007), .Y(new_n4325));
  nand_5 g03949(.A(new_n987), .B(new_n986), .Y(new_n4326));
  nand_5 g03950(.A(new_n988), .B(new_n985), .Y(new_n4327));
  nand_5 g03951(.A(new_n4327), .B(new_n4326), .Y(new_n4328));
  xor_4  g03952(.A(new_n4328), .B(new_n4325), .Y(new_n4329));
  xnor_4 g03953(.A(new_n4329), .B(new_n4324), .Y(new_n4330));
  xor_4  g03954(.A(new_n4330), .B(new_n4319), .Y(new_n4331));
  xnor_4 g03955(.A(new_n4331), .B(new_n4314), .Y(new_n4332));
  xor_4  g03956(.A(new_n4332), .B(new_n4313), .Y(new_n4333));
  xnor_4 g03957(.A(new_n4333), .B(new_n4310), .Y(new_n4334));
  xor_4  g03958(.A(new_n4290), .B(new_n4270), .Y(new_n4335));
  nand_5 g03959(.A(new_n4335), .B(new_n4334), .Y(new_n4336));
  nand_5 g03960(.A(new_n4336), .B(new_n4291), .Y(new_n4337));
  not_8  g03961(.A(new_n4271), .Y(new_n4338));
  nand_5 g03962(.A(new_n4289), .B(new_n4338), .Y(new_n4339));
  nand_5 g03963(.A(pi238), .B(pi175), .Y(new_n4340));
  xor_4  g03964(.A(new_n4340), .B(new_n4339), .Y(new_n4341));
  nand_5 g03965(.A(new_n4286), .B(new_n4285), .Y(new_n4342));
  nand_5 g03966(.A(new_n4287), .B(new_n4282), .Y(new_n4343));
  nand_5 g03967(.A(new_n4343), .B(new_n4342), .Y(new_n4344));
  nand_5 g03968(.A(pi167), .B(pi033), .Y(new_n4345));
  nand_5 g03969(.A(pi181), .B(pi162), .Y(new_n4346));
  nand_5 g03970(.A(new_n4346), .B(new_n4345), .Y(new_n4347));
  nand_5 g03971(.A(pi181), .B(pi033), .Y(new_n4348));
  nor_5  g03972(.A(new_n4348), .B(new_n4278), .Y(new_n4349));
  not_8  g03973(.A(new_n4349), .Y(new_n4350));
  nand_5 g03974(.A(new_n4350), .B(new_n4347), .Y(new_n4351));
  nand_5 g03975(.A(pi179), .B(pi149), .Y(new_n4352));
  nand_5 g03976(.A(new_n4280), .B(new_n4279), .Y(new_n4353));
  nand_5 g03977(.A(new_n4281), .B(new_n4278), .Y(new_n4354));
  nand_5 g03978(.A(new_n4354), .B(new_n4353), .Y(new_n4355));
  xnor_4 g03979(.A(new_n4355), .B(new_n4352), .Y(new_n4356));
  xor_4  g03980(.A(new_n4356), .B(new_n4351), .Y(new_n4357));
  nand_5 g03981(.A(pi240), .B(pi048), .Y(new_n4358));
  nand_5 g03982(.A(pi237), .B(pi134), .Y(new_n4359));
  and_6  g03983(.A(new_n4359), .B(new_n4358), .Y(new_n4360));
  nand_5 g03984(.A(pi240), .B(pi237), .Y(new_n4361));
  nor_5  g03985(.A(new_n4361), .B(new_n4286), .Y(new_n4362));
  or_6   g03986(.A(new_n4362), .B(new_n4360), .Y(new_n4363));
  xor_4  g03987(.A(new_n4363), .B(new_n4357), .Y(new_n4364));
  xor_4  g03988(.A(new_n4364), .B(new_n4344), .Y(new_n4365));
  nor_5  g03989(.A(new_n4276), .B(new_n4272), .Y(new_n4366));
  nand_5 g03990(.A(new_n4288), .B(new_n4277), .Y(new_n4367));
  not_8  g03991(.A(new_n4367), .Y(new_n4368));
  nor_5  g03992(.A(new_n4368), .B(new_n4366), .Y(new_n4369));
  xor_4  g03993(.A(new_n4369), .B(new_n4365), .Y(new_n4370));
  xnor_4 g03994(.A(new_n4370), .B(new_n4341), .Y(new_n4371));
  nand_5 g03995(.A(new_n4371), .B(new_n4337), .Y(new_n4372));
  xor_4  g03996(.A(new_n4371), .B(new_n4337), .Y(new_n4373));
  not_8  g03997(.A(new_n4332), .Y(new_n4374));
  nor_5  g03998(.A(new_n4374), .B(new_n4313), .Y(new_n4375));
  nor_5  g03999(.A(new_n4333), .B(new_n4310), .Y(new_n4376));
  nor_5  g04000(.A(new_n4376), .B(new_n4375), .Y(new_n4377));
  nand_5 g04001(.A(new_n4309), .B(new_n4292), .Y(new_n4378));
  nand_5 g04002(.A(pi163), .B(pi098), .Y(new_n4379));
  nor_5  g04003(.A(new_n4304), .B(new_n4293), .Y(new_n4380));
  nor_5  g04004(.A(new_n4308), .B(new_n4305), .Y(new_n4381));
  nor_5  g04005(.A(new_n4381), .B(new_n4380), .Y(new_n4382));
  nand_5 g04006(.A(new_n4302), .B(new_n4301), .Y(new_n4383));
  nand_5 g04007(.A(new_n4303), .B(new_n4298), .Y(new_n4384));
  nand_5 g04008(.A(new_n4384), .B(new_n4383), .Y(new_n4385));
  nand_5 g04009(.A(pi228), .B(pi012), .Y(new_n4386));
  nand_5 g04010(.A(pi148), .B(pi144), .Y(new_n4387));
  and_6  g04011(.A(new_n4387), .B(new_n4386), .Y(new_n4388));
  nand_5 g04012(.A(pi228), .B(pi144), .Y(new_n4389));
  nor_5  g04013(.A(new_n4389), .B(new_n4302), .Y(new_n4390));
  or_6   g04014(.A(new_n4390), .B(new_n4388), .Y(new_n4391));
  nand_5 g04015(.A(new_n4296), .B(new_n4295), .Y(new_n4392));
  nand_5 g04016(.A(new_n4297), .B(new_n4294), .Y(new_n4393));
  nand_5 g04017(.A(new_n4393), .B(new_n4392), .Y(new_n4394));
  nand_5 g04018(.A(pi061), .B(pi039), .Y(new_n4395));
  nand_5 g04019(.A(pi178), .B(pi116), .Y(new_n4396));
  nand_5 g04020(.A(pi188), .B(pi070), .Y(new_n4397));
  nand_5 g04021(.A(new_n4397), .B(new_n4396), .Y(new_n4398));
  nand_5 g04022(.A(pi178), .B(pi070), .Y(new_n4399));
  nor_5  g04023(.A(new_n4399), .B(new_n4296), .Y(new_n4400));
  not_8  g04024(.A(new_n4400), .Y(new_n4401));
  nand_5 g04025(.A(new_n4401), .B(new_n4398), .Y(new_n4402));
  xor_4  g04026(.A(new_n4402), .B(new_n4395), .Y(new_n4403));
  xor_4  g04027(.A(new_n4403), .B(new_n4394), .Y(new_n4404));
  xor_4  g04028(.A(new_n4404), .B(new_n4391), .Y(new_n4405));
  not_8  g04029(.A(new_n4405), .Y(new_n4406));
  xor_4  g04030(.A(new_n4406), .B(new_n4385), .Y(new_n4407));
  xor_4  g04031(.A(new_n4407), .B(new_n4382), .Y(new_n4408));
  xor_4  g04032(.A(new_n4408), .B(new_n4379), .Y(new_n4409));
  xor_4  g04033(.A(new_n4409), .B(new_n4378), .Y(new_n4410));
  nand_5 g04034(.A(new_n4331), .B(new_n4314), .Y(new_n4411));
  nand_5 g04035(.A(pi113), .B(pi107), .Y(new_n4412));
  xor_4  g04036(.A(new_n4412), .B(new_n4411), .Y(new_n4413));
  nand_5 g04037(.A(pi245), .B(pi108), .Y(new_n4414));
  nand_5 g04038(.A(pi201), .B(pi042), .Y(new_n4415));
  nand_5 g04039(.A(pi156), .B(pi051), .Y(new_n4416));
  nand_5 g04040(.A(new_n4416), .B(new_n4415), .Y(new_n4417));
  nand_5 g04041(.A(pi156), .B(pi042), .Y(new_n4418));
  nor_5  g04042(.A(new_n4418), .B(new_n4322), .Y(new_n4419));
  not_8  g04043(.A(new_n4419), .Y(new_n4420));
  nand_5 g04044(.A(new_n4420), .B(new_n4417), .Y(new_n4421));
  xor_4  g04045(.A(new_n4421), .B(new_n4414), .Y(new_n4422));
  nand_5 g04046(.A(new_n4322), .B(new_n4321), .Y(new_n4423));
  nand_5 g04047(.A(new_n4323), .B(new_n4320), .Y(new_n4424));
  nand_5 g04048(.A(new_n4424), .B(new_n4423), .Y(new_n4425));
  xor_4  g04049(.A(new_n4425), .B(new_n4422), .Y(new_n4426));
  nand_5 g04050(.A(pi049), .B(pi007), .Y(new_n4427));
  nand_5 g04051(.A(pi171), .B(pi118), .Y(new_n4428));
  and_6  g04052(.A(new_n4428), .B(new_n4427), .Y(new_n4429));
  nand_5 g04053(.A(pi118), .B(pi049), .Y(new_n4430));
  nor_5  g04054(.A(new_n4430), .B(new_n4325), .Y(new_n4431));
  or_6   g04055(.A(new_n4431), .B(new_n4429), .Y(new_n4432));
  xor_4  g04056(.A(new_n4432), .B(new_n4426), .Y(new_n4433));
  not_8  g04057(.A(new_n4433), .Y(new_n4434));
  nand_5 g04058(.A(new_n4328), .B(new_n4325), .Y(new_n4435));
  nand_5 g04059(.A(new_n4329), .B(new_n4324), .Y(new_n4436));
  nand_5 g04060(.A(new_n4436), .B(new_n4435), .Y(new_n4437));
  xor_4  g04061(.A(new_n4437), .B(new_n4434), .Y(new_n4438));
  nor_5  g04062(.A(new_n4318), .B(new_n4315), .Y(new_n4439));
  nand_5 g04063(.A(new_n4330), .B(new_n4319), .Y(new_n4440));
  not_8  g04064(.A(new_n4440), .Y(new_n4441));
  nor_5  g04065(.A(new_n4441), .B(new_n4439), .Y(new_n4442));
  xor_4  g04066(.A(new_n4442), .B(new_n4438), .Y(new_n4443));
  xor_4  g04067(.A(new_n4443), .B(new_n4413), .Y(new_n4444));
  xor_4  g04068(.A(new_n4444), .B(new_n4410), .Y(new_n4445));
  xor_4  g04069(.A(new_n4445), .B(new_n4377), .Y(new_n4446));
  nand_5 g04070(.A(new_n4446), .B(new_n4373), .Y(new_n4447));
  nand_5 g04071(.A(new_n4447), .B(new_n4372), .Y(new_n4448));
  or_6   g04072(.A(new_n4444), .B(new_n4410), .Y(new_n4449));
  nand_5 g04073(.A(new_n4445), .B(new_n4377), .Y(new_n4450));
  nand_5 g04074(.A(new_n4450), .B(new_n4449), .Y(new_n4451));
  nand_5 g04075(.A(new_n4412), .B(new_n4411), .Y(new_n4452));
  nand_5 g04076(.A(new_n4443), .B(new_n4413), .Y(new_n4453));
  nand_5 g04077(.A(new_n4453), .B(new_n4452), .Y(new_n4454));
  not_8  g04078(.A(new_n4438), .Y(new_n4455));
  nor_5  g04079(.A(new_n4442), .B(new_n4455), .Y(new_n4456));
  nor_5  g04080(.A(new_n4432), .B(new_n4426), .Y(new_n4457));
  nor_5  g04081(.A(new_n4437), .B(new_n4434), .Y(new_n4458));
  xor_4  g04082(.A(new_n4458), .B(new_n4431), .Y(new_n4459));
  nor_5  g04083(.A(new_n4459), .B(new_n4457), .Y(new_n4460));
  nand_5 g04084(.A(pi063), .B(pi051), .Y(new_n4461));
  nand_5 g04085(.A(pi201), .B(pi108), .Y(new_n4462));
  xor_4  g04086(.A(new_n4462), .B(new_n4461), .Y(new_n4463));
  xor_4  g04087(.A(new_n4463), .B(new_n4418), .Y(new_n4464));
  nand_5 g04088(.A(pi245), .B(pi007), .Y(new_n4465));
  xor_4  g04089(.A(new_n4465), .B(new_n4419), .Y(new_n4466));
  xor_4  g04090(.A(new_n4466), .B(new_n4464), .Y(new_n4467));
  nand_5 g04091(.A(new_n4421), .B(new_n4414), .Y(new_n4468));
  nand_5 g04092(.A(new_n4425), .B(new_n4422), .Y(new_n4469));
  nand_5 g04093(.A(new_n4469), .B(new_n4468), .Y(new_n4470));
  nand_5 g04094(.A(pi107), .B(pi038), .Y(new_n4471));
  nand_5 g04095(.A(pi171), .B(pi113), .Y(new_n4472));
  xor_4  g04096(.A(new_n4472), .B(new_n4471), .Y(new_n4473));
  xor_4  g04097(.A(new_n4473), .B(new_n4430), .Y(new_n4474));
  xor_4  g04098(.A(new_n4474), .B(new_n4470), .Y(new_n4475));
  xnor_4 g04099(.A(new_n4475), .B(new_n4467), .Y(new_n4476));
  xor_4  g04100(.A(new_n4476), .B(new_n4460), .Y(new_n4477));
  xor_4  g04101(.A(new_n4477), .B(new_n4456), .Y(new_n4478));
  xnor_4 g04102(.A(new_n4478), .B(new_n4454), .Y(new_n4479));
  nand_5 g04103(.A(new_n4408), .B(new_n4379), .Y(new_n4480));
  nand_5 g04104(.A(new_n4409), .B(new_n4378), .Y(new_n4481));
  nand_5 g04105(.A(new_n4481), .B(new_n4480), .Y(new_n4482));
  not_8  g04106(.A(new_n4407), .Y(new_n4483));
  nor_5  g04107(.A(new_n4483), .B(new_n4382), .Y(new_n4484));
  nand_5 g04108(.A(pi188), .B(pi115), .Y(new_n4485));
  nand_5 g04109(.A(pi116), .B(pi061), .Y(new_n4486));
  xor_4  g04110(.A(new_n4486), .B(new_n4485), .Y(new_n4487));
  xor_4  g04111(.A(new_n4487), .B(new_n4399), .Y(new_n4488));
  nand_5 g04112(.A(pi039), .B(pi012), .Y(new_n4489));
  xor_4  g04113(.A(new_n4489), .B(new_n4400), .Y(new_n4490));
  xor_4  g04114(.A(new_n4490), .B(new_n4488), .Y(new_n4491));
  nand_5 g04115(.A(new_n4402), .B(new_n4395), .Y(new_n4492));
  nand_5 g04116(.A(new_n4403), .B(new_n4394), .Y(new_n4493));
  nand_5 g04117(.A(new_n4493), .B(new_n4492), .Y(new_n4494));
  nand_5 g04118(.A(pi148), .B(pi098), .Y(new_n4495));
  nand_5 g04119(.A(pi163), .B(pi043), .Y(new_n4496));
  xor_4  g04120(.A(new_n4496), .B(new_n4495), .Y(new_n4497));
  xnor_4 g04121(.A(new_n4497), .B(new_n4389), .Y(new_n4498));
  xor_4  g04122(.A(new_n4498), .B(new_n4494), .Y(new_n4499));
  xor_4  g04123(.A(new_n4499), .B(new_n4491), .Y(new_n4500));
  nor_5  g04124(.A(new_n4404), .B(new_n4391), .Y(new_n4501));
  nor_5  g04125(.A(new_n4406), .B(new_n4385), .Y(new_n4502));
  xor_4  g04126(.A(new_n4502), .B(new_n4390), .Y(new_n4503));
  nor_5  g04127(.A(new_n4503), .B(new_n4501), .Y(new_n4504));
  xor_4  g04128(.A(new_n4504), .B(new_n4500), .Y(new_n4505));
  xor_4  g04129(.A(new_n4505), .B(new_n4484), .Y(new_n4506));
  xor_4  g04130(.A(new_n4506), .B(new_n4482), .Y(new_n4507));
  xor_4  g04131(.A(new_n4507), .B(new_n4479), .Y(new_n4508));
  xnor_4 g04132(.A(new_n4508), .B(new_n4451), .Y(new_n4509));
  nand_5 g04133(.A(new_n4340), .B(new_n4339), .Y(new_n4510));
  nand_5 g04134(.A(new_n4370), .B(new_n4341), .Y(new_n4511));
  nand_5 g04135(.A(new_n4511), .B(new_n4510), .Y(new_n4512));
  not_8  g04136(.A(new_n4365), .Y(new_n4513));
  nor_5  g04137(.A(new_n4369), .B(new_n4513), .Y(new_n4514));
  nor_5  g04138(.A(new_n4355), .B(new_n4352), .Y(new_n4515));
  nor_5  g04139(.A(new_n4356), .B(new_n4351), .Y(new_n4516));
  nor_5  g04140(.A(new_n4516), .B(new_n4515), .Y(new_n4517));
  nand_5 g04141(.A(pi238), .B(pi134), .Y(new_n4518));
  nand_5 g04142(.A(pi193), .B(pi175), .Y(new_n4519));
  xor_4  g04143(.A(new_n4519), .B(new_n4518), .Y(new_n4520));
  xor_4  g04144(.A(new_n4520), .B(new_n4361), .Y(new_n4521));
  xor_4  g04145(.A(new_n4521), .B(new_n4517), .Y(new_n4522));
  nand_5 g04146(.A(pi149), .B(pi048), .Y(new_n4523));
  xor_4  g04147(.A(new_n4523), .B(new_n4349), .Y(new_n4524));
  nand_5 g04148(.A(pi200), .B(pi162), .Y(new_n4525));
  nand_5 g04149(.A(pi179), .B(pi167), .Y(new_n4526));
  xor_4  g04150(.A(new_n4526), .B(new_n4525), .Y(new_n4527));
  xor_4  g04151(.A(new_n4527), .B(new_n4348), .Y(new_n4528));
  xor_4  g04152(.A(new_n4528), .B(new_n4524), .Y(new_n4529));
  not_8  g04153(.A(new_n4529), .Y(new_n4530));
  xor_4  g04154(.A(new_n4530), .B(new_n4522), .Y(new_n4531));
  not_8  g04155(.A(new_n4357), .Y(new_n4532));
  nor_5  g04156(.A(new_n4363), .B(new_n4532), .Y(new_n4533));
  nor_5  g04157(.A(new_n4364), .B(new_n4344), .Y(new_n4534));
  xor_4  g04158(.A(new_n4534), .B(new_n4362), .Y(new_n4535));
  nor_5  g04159(.A(new_n4535), .B(new_n4533), .Y(new_n4536));
  xor_4  g04160(.A(new_n4536), .B(new_n4531), .Y(new_n4537));
  xnor_4 g04161(.A(new_n4537), .B(new_n4514), .Y(new_n4538));
  xor_4  g04162(.A(new_n4538), .B(new_n4512), .Y(new_n4539));
  xor_4  g04163(.A(new_n4539), .B(new_n4509), .Y(new_n4540));
  xor_4  g04164(.A(new_n4540), .B(new_n4448), .Y(new_n4541));
  nor_5  g04165(.A(new_n1051), .B(new_n1033), .Y(new_n4542));
  nor_5  g04166(.A(new_n1052), .B(new_n1012), .Y(new_n4543));
  nor_5  g04167(.A(new_n4543), .B(new_n4542), .Y(new_n4544));
  not_8  g04168(.A(new_n1032), .Y(new_n4545));
  nand_5 g04169(.A(new_n4545), .B(new_n1021), .Y(new_n4546));
  nand_5 g04170(.A(pi180), .B(pi103), .Y(new_n4547));
  nand_5 g04171(.A(new_n1030), .B(new_n1027), .Y(new_n4548));
  nand_5 g04172(.A(new_n1031), .B(new_n1026), .Y(new_n4549));
  nand_5 g04173(.A(new_n4549), .B(new_n4548), .Y(new_n4550));
  xor_4  g04174(.A(new_n4550), .B(new_n4547), .Y(new_n4551));
  nand_5 g04175(.A(pi194), .B(pi016), .Y(new_n4552));
  nand_5 g04176(.A(pi080), .B(pi057), .Y(new_n4553));
  nand_5 g04177(.A(pi247), .B(pi143), .Y(new_n4554));
  xor_4  g04178(.A(new_n4554), .B(new_n4553), .Y(new_n4555));
  xor_4  g04179(.A(new_n4555), .B(new_n4552), .Y(new_n4556));
  nand_5 g04180(.A(pi117), .B(pi085), .Y(new_n4557));
  nand_5 g04181(.A(new_n1024), .B(new_n1023), .Y(new_n4558));
  nand_5 g04182(.A(new_n1025), .B(new_n1022), .Y(new_n4559));
  nand_5 g04183(.A(new_n4559), .B(new_n4558), .Y(new_n4560));
  xor_4  g04184(.A(new_n4560), .B(new_n4557), .Y(new_n4561));
  xor_4  g04185(.A(new_n4561), .B(new_n4556), .Y(new_n4562));
  not_8  g04186(.A(new_n4562), .Y(new_n4563));
  xor_4  g04187(.A(new_n4563), .B(new_n4551), .Y(new_n4564));
  xor_4  g04188(.A(new_n4564), .B(new_n4546), .Y(new_n4565));
  and_6  g04189(.A(new_n4565), .B(new_n4544), .Y(new_n4566));
  xor_4  g04190(.A(new_n4335), .B(new_n4334), .Y(new_n4567));
  xnor_4 g04191(.A(new_n4565), .B(new_n4544), .Y(new_n4568));
  nor_5  g04192(.A(new_n4568), .B(new_n4567), .Y(new_n4569));
  or_6   g04193(.A(new_n4569), .B(new_n4566), .Y(new_n4570));
  not_8  g04194(.A(new_n4546), .Y(new_n4571));
  nand_5 g04195(.A(new_n4564), .B(new_n4571), .Y(new_n4572));
  nand_5 g04196(.A(pi103), .B(pi036), .Y(new_n4573));
  xor_4  g04197(.A(new_n4573), .B(new_n4572), .Y(new_n4574));
  nor_5  g04198(.A(new_n4550), .B(new_n4547), .Y(new_n4575));
  nand_5 g04199(.A(new_n4563), .B(new_n4551), .Y(new_n4576));
  not_8  g04200(.A(new_n4576), .Y(new_n4577));
  nor_5  g04201(.A(new_n4577), .B(new_n4575), .Y(new_n4578));
  nand_5 g04202(.A(pi085), .B(pi016), .Y(new_n4579));
  nand_5 g04203(.A(pi180), .B(pi117), .Y(new_n4580));
  nand_5 g04204(.A(new_n4580), .B(new_n4579), .Y(new_n4581));
  nand_5 g04205(.A(pi180), .B(pi016), .Y(new_n4582));
  nor_5  g04206(.A(new_n4582), .B(new_n4557), .Y(new_n4583));
  not_8  g04207(.A(new_n4583), .Y(new_n4584));
  nand_5 g04208(.A(new_n4584), .B(new_n4581), .Y(new_n4585));
  nand_5 g04209(.A(pi194), .B(pi080), .Y(new_n4586));
  nand_5 g04210(.A(new_n4554), .B(new_n4553), .Y(new_n4587));
  nand_5 g04211(.A(new_n4555), .B(new_n4552), .Y(new_n4588));
  nand_5 g04212(.A(new_n4588), .B(new_n4587), .Y(new_n4589));
  xor_4  g04213(.A(new_n4589), .B(new_n4586), .Y(new_n4590));
  nand_5 g04214(.A(pi247), .B(pi057), .Y(new_n4591));
  nand_5 g04215(.A(pi234), .B(pi143), .Y(new_n4592));
  nand_5 g04216(.A(new_n4592), .B(new_n4591), .Y(new_n4593));
  nand_5 g04217(.A(pi234), .B(pi057), .Y(new_n4594));
  nor_5  g04218(.A(new_n4594), .B(new_n4554), .Y(new_n4595));
  not_8  g04219(.A(new_n4595), .Y(new_n4596));
  nand_5 g04220(.A(new_n4596), .B(new_n4593), .Y(new_n4597));
  xor_4  g04221(.A(new_n4597), .B(new_n4590), .Y(new_n4598));
  xor_4  g04222(.A(new_n4598), .B(new_n4585), .Y(new_n4599));
  nand_5 g04223(.A(new_n4560), .B(new_n4557), .Y(new_n4600));
  nand_5 g04224(.A(new_n4561), .B(new_n4556), .Y(new_n4601));
  nand_5 g04225(.A(new_n4601), .B(new_n4600), .Y(new_n4602));
  xor_4  g04226(.A(new_n4602), .B(new_n4599), .Y(new_n4603));
  xnor_4 g04227(.A(new_n4603), .B(new_n4578), .Y(new_n4604));
  xor_4  g04228(.A(new_n4604), .B(new_n4574), .Y(new_n4605));
  and_6  g04229(.A(new_n4605), .B(new_n4570), .Y(new_n4606));
  xor_4  g04230(.A(new_n4446), .B(new_n4373), .Y(new_n4607));
  xnor_4 g04231(.A(new_n4605), .B(new_n4570), .Y(new_n4608));
  nor_5  g04232(.A(new_n4608), .B(new_n4607), .Y(new_n4609));
  nor_5  g04233(.A(new_n4609), .B(new_n4606), .Y(new_n4610));
  nor_5  g04234(.A(new_n4603), .B(new_n4578), .Y(new_n4611));
  not_8  g04235(.A(new_n4611), .Y(new_n4612));
  nor_5  g04236(.A(new_n4598), .B(new_n4585), .Y(new_n4613));
  not_8  g04237(.A(new_n4599), .Y(new_n4614));
  nor_5  g04238(.A(new_n4602), .B(new_n4614), .Y(new_n4615));
  xor_4  g04239(.A(new_n4615), .B(new_n4584), .Y(new_n4616));
  not_8  g04240(.A(new_n4616), .Y(new_n4617));
  nor_5  g04241(.A(new_n4617), .B(new_n4613), .Y(new_n4618));
  nand_5 g04242(.A(pi117), .B(pi036), .Y(new_n4619));
  nand_5 g04243(.A(pi103), .B(pi068), .Y(new_n4620));
  xor_4  g04244(.A(new_n4620), .B(new_n4619), .Y(new_n4621));
  xor_4  g04245(.A(new_n4621), .B(new_n4582), .Y(new_n4622));
  nor_5  g04246(.A(new_n4589), .B(new_n4586), .Y(new_n4623));
  not_8  g04247(.A(new_n4590), .Y(new_n4624));
  nor_5  g04248(.A(new_n4597), .B(new_n4624), .Y(new_n4625));
  nor_5  g04249(.A(new_n4625), .B(new_n4623), .Y(new_n4626));
  xor_4  g04250(.A(new_n4626), .B(new_n4622), .Y(new_n4627));
  nand_5 g04251(.A(pi085), .B(pi080), .Y(new_n4628));
  xor_4  g04252(.A(new_n4628), .B(new_n4596), .Y(new_n4629));
  nand_5 g04253(.A(pi214), .B(pi143), .Y(new_n4630));
  nand_5 g04254(.A(pi247), .B(pi194), .Y(new_n4631));
  xor_4  g04255(.A(new_n4631), .B(new_n4630), .Y(new_n4632));
  xor_4  g04256(.A(new_n4632), .B(new_n4594), .Y(new_n4633));
  xor_4  g04257(.A(new_n4633), .B(new_n4629), .Y(new_n4634));
  xnor_4 g04258(.A(new_n4634), .B(new_n4627), .Y(new_n4635));
  xor_4  g04259(.A(new_n4635), .B(new_n4618), .Y(new_n4636));
  or_6   g04260(.A(new_n4636), .B(new_n4612), .Y(new_n4637));
  nand_5 g04261(.A(new_n4636), .B(new_n4612), .Y(new_n4638));
  nand_5 g04262(.A(new_n4638), .B(new_n4637), .Y(new_n4639));
  nand_5 g04263(.A(new_n4573), .B(new_n4572), .Y(new_n4640));
  nand_5 g04264(.A(new_n4604), .B(new_n4574), .Y(new_n4641));
  nand_5 g04265(.A(new_n4641), .B(new_n4640), .Y(new_n4642));
  xor_4  g04266(.A(new_n4642), .B(new_n4639), .Y(new_n4643));
  xnor_4 g04267(.A(new_n4643), .B(new_n4610), .Y(new_n4644));
  xnor_4 g04268(.A(new_n4644), .B(new_n4541), .Y(po014));
  nand_5 g04269(.A(pi143), .B(pi077), .Y(new_n4646));
  nand_5 g04270(.A(pi057), .B(pi052), .Y(new_n4647));
  nand_5 g04271(.A(pi194), .B(pi131), .Y(new_n4648));
  xor_4  g04272(.A(new_n4648), .B(new_n4647), .Y(new_n4649));
  xor_4  g04273(.A(new_n4649), .B(new_n4646), .Y(new_n4650));
  not_8  g04274(.A(new_n4650), .Y(new_n4651));
  nand_5 g04275(.A(pi131), .B(pi057), .Y(new_n4652));
  nand_5 g04276(.A(pi143), .B(pi052), .Y(new_n4653));
  nor_5  g04277(.A(new_n4653), .B(new_n4652), .Y(new_n4654));
  nand_5 g04278(.A(new_n4654), .B(new_n4651), .Y(new_n4655));
  nand_5 g04279(.A(pi077), .B(pi057), .Y(new_n4656));
  nand_5 g04280(.A(pi194), .B(pi052), .Y(new_n4657));
  nand_5 g04281(.A(pi143), .B(pi133), .Y(new_n4658));
  xor_4  g04282(.A(new_n4658), .B(new_n4657), .Y(new_n4659));
  xor_4  g04283(.A(new_n4659), .B(new_n4656), .Y(new_n4660));
  nand_5 g04284(.A(pi131), .B(pi085), .Y(new_n4661));
  nand_5 g04285(.A(new_n4648), .B(new_n4647), .Y(new_n4662));
  nand_5 g04286(.A(new_n4649), .B(new_n4646), .Y(new_n4663));
  nand_5 g04287(.A(new_n4663), .B(new_n4662), .Y(new_n4664));
  xor_4  g04288(.A(new_n4664), .B(new_n4661), .Y(new_n4665));
  xor_4  g04289(.A(new_n4665), .B(new_n4660), .Y(new_n4666));
  xor_4  g04290(.A(new_n4666), .B(new_n4655), .Y(new_n4667));
  nand_5 g04291(.A(pi162), .B(pi139), .Y(new_n4668));
  nand_5 g04292(.A(pi208), .B(pi033), .Y(new_n4669));
  nand_5 g04293(.A(pi179), .B(pi168), .Y(new_n4670));
  xor_4  g04294(.A(new_n4670), .B(new_n4669), .Y(new_n4671));
  xor_4  g04295(.A(new_n4671), .B(new_n4668), .Y(new_n4672));
  or_6   g04296(.A(new_n4669), .B(new_n3555), .Y(new_n4673));
  or_6   g04297(.A(new_n4673), .B(new_n4672), .Y(new_n4674));
  nand_5 g04298(.A(pi208), .B(pi179), .Y(new_n4675));
  nand_5 g04299(.A(pi162), .B(pi035), .Y(new_n4676));
  nand_5 g04300(.A(pi139), .B(pi033), .Y(new_n4677));
  xor_4  g04301(.A(new_n4677), .B(new_n4676), .Y(new_n4678));
  xor_4  g04302(.A(new_n4678), .B(new_n4675), .Y(new_n4679));
  nand_5 g04303(.A(pi168), .B(pi048), .Y(new_n4680));
  nand_5 g04304(.A(new_n4670), .B(new_n4669), .Y(new_n4681));
  nand_5 g04305(.A(new_n4671), .B(new_n4668), .Y(new_n4682));
  nand_5 g04306(.A(new_n4682), .B(new_n4681), .Y(new_n4683));
  xor_4  g04307(.A(new_n4683), .B(new_n4680), .Y(new_n4684));
  xor_4  g04308(.A(new_n4684), .B(new_n4679), .Y(new_n4685));
  xor_4  g04309(.A(new_n4685), .B(new_n4674), .Y(new_n4686));
  not_8  g04310(.A(new_n4686), .Y(new_n4687));
  nand_5 g04311(.A(pi188), .B(pi104), .Y(new_n4688));
  nand_5 g04312(.A(pi212), .B(pi178), .Y(new_n4689));
  nand_5 g04313(.A(pi213), .B(pi061), .Y(new_n4690));
  xor_4  g04314(.A(new_n4690), .B(new_n4689), .Y(new_n4691));
  xnor_4 g04315(.A(new_n4691), .B(new_n4688), .Y(new_n4692));
  or_6   g04316(.A(new_n4689), .B(new_n3557), .Y(new_n4693));
  not_8  g04317(.A(new_n4693), .Y(new_n4694));
  xor_4  g04318(.A(new_n4694), .B(new_n4692), .Y(new_n4695));
  not_8  g04319(.A(new_n4695), .Y(new_n4696));
  or_6   g04320(.A(new_n3557), .B(new_n3556), .Y(new_n4697));
  nand_5 g04321(.A(pi241), .B(pi042), .Y(new_n4698));
  or_6   g04322(.A(new_n4698), .B(new_n3556), .Y(new_n4699));
  nand_5 g04323(.A(pi236), .B(pi042), .Y(new_n4700));
  nand_5 g04324(.A(pi241), .B(pi051), .Y(new_n4701));
  nand_5 g04325(.A(new_n4701), .B(new_n4700), .Y(new_n4702));
  nand_5 g04326(.A(new_n4702), .B(new_n4699), .Y(new_n4703));
  nand_5 g04327(.A(new_n4703), .B(new_n4697), .Y(new_n4704));
  or_6   g04328(.A(new_n4703), .B(new_n4697), .Y(new_n4705));
  nand_5 g04329(.A(pi213), .B(pi178), .Y(new_n4706));
  nand_5 g04330(.A(pi212), .B(pi188), .Y(new_n4707));
  nand_5 g04331(.A(new_n4707), .B(new_n4706), .Y(new_n4708));
  nand_5 g04332(.A(new_n4708), .B(new_n4693), .Y(new_n4709));
  nand_5 g04333(.A(new_n4709), .B(new_n4705), .Y(new_n4710));
  nand_5 g04334(.A(new_n4710), .B(new_n4704), .Y(new_n4711));
  nand_5 g04335(.A(new_n4711), .B(new_n4696), .Y(new_n4712));
  nand_5 g04336(.A(pi161), .B(pi051), .Y(new_n4713));
  nand_5 g04337(.A(pi236), .B(pi108), .Y(new_n4714));
  xor_4  g04338(.A(new_n4714), .B(new_n4698), .Y(new_n4715));
  xor_4  g04339(.A(new_n4715), .B(new_n4713), .Y(new_n4716));
  xor_4  g04340(.A(new_n4716), .B(new_n4699), .Y(new_n4717));
  xor_4  g04341(.A(new_n4711), .B(new_n4695), .Y(new_n4718));
  or_6   g04342(.A(new_n4718), .B(new_n4717), .Y(new_n4719));
  nand_5 g04343(.A(new_n4719), .B(new_n4712), .Y(new_n4720));
  nor_5  g04344(.A(new_n4716), .B(new_n4699), .Y(new_n4721));
  nand_5 g04345(.A(pi141), .B(pi051), .Y(new_n4722));
  nand_5 g04346(.A(pi241), .B(pi108), .Y(new_n4723));
  nand_5 g04347(.A(pi161), .B(pi042), .Y(new_n4724));
  xor_4  g04348(.A(new_n4724), .B(new_n4723), .Y(new_n4725));
  xor_4  g04349(.A(new_n4725), .B(new_n4722), .Y(new_n4726));
  nand_5 g04350(.A(pi236), .B(pi007), .Y(new_n4727));
  nand_5 g04351(.A(new_n4714), .B(new_n4698), .Y(new_n4728));
  nand_5 g04352(.A(new_n4715), .B(new_n4713), .Y(new_n4729));
  nand_5 g04353(.A(new_n4729), .B(new_n4728), .Y(new_n4730));
  xnor_4 g04354(.A(new_n4730), .B(new_n4727), .Y(new_n4731));
  xnor_4 g04355(.A(new_n4731), .B(new_n4726), .Y(new_n4732));
  xor_4  g04356(.A(new_n4732), .B(new_n4721), .Y(new_n4733));
  nand_5 g04357(.A(new_n4694), .B(new_n4692), .Y(new_n4734));
  nand_5 g04358(.A(pi188), .B(pi013), .Y(new_n4735));
  nand_5 g04359(.A(pi212), .B(pi061), .Y(new_n4736));
  nand_5 g04360(.A(pi178), .B(pi104), .Y(new_n4737));
  xor_4  g04361(.A(new_n4737), .B(new_n4736), .Y(new_n4738));
  xor_4  g04362(.A(new_n4738), .B(new_n4735), .Y(new_n4739));
  nand_5 g04363(.A(pi213), .B(pi012), .Y(new_n4740));
  nand_5 g04364(.A(new_n4690), .B(new_n4689), .Y(new_n4741));
  nand_5 g04365(.A(new_n4691), .B(new_n4688), .Y(new_n4742));
  nand_5 g04366(.A(new_n4742), .B(new_n4741), .Y(new_n4743));
  xor_4  g04367(.A(new_n4743), .B(new_n4740), .Y(new_n4744));
  xnor_4 g04368(.A(new_n4744), .B(new_n4739), .Y(new_n4745));
  xor_4  g04369(.A(new_n4745), .B(new_n4734), .Y(new_n4746));
  xor_4  g04370(.A(new_n4746), .B(new_n4733), .Y(new_n4747));
  xor_4  g04371(.A(new_n4747), .B(new_n4720), .Y(new_n4748));
  xor_4  g04372(.A(new_n4748), .B(new_n4687), .Y(new_n4749));
  xor_4  g04373(.A(new_n4673), .B(new_n4672), .Y(new_n4750));
  not_8  g04374(.A(new_n4750), .Y(new_n4751));
  or_6   g04375(.A(new_n3558), .B(new_n3555), .Y(new_n4752));
  nand_5 g04376(.A(pi168), .B(pi033), .Y(new_n4753));
  nand_5 g04377(.A(pi208), .B(pi162), .Y(new_n4754));
  nand_5 g04378(.A(new_n4754), .B(new_n4753), .Y(new_n4755));
  nand_5 g04379(.A(new_n4755), .B(new_n4673), .Y(new_n4756));
  nand_5 g04380(.A(new_n4756), .B(new_n4752), .Y(new_n4757));
  xor_4  g04381(.A(new_n4756), .B(new_n4752), .Y(new_n4758));
  not_8  g04382(.A(new_n4758), .Y(new_n4759));
  nand_5 g04383(.A(new_n4705), .B(new_n4704), .Y(new_n4760));
  xor_4  g04384(.A(new_n4760), .B(new_n4709), .Y(new_n4761));
  or_6   g04385(.A(new_n4761), .B(new_n4759), .Y(new_n4762));
  nand_5 g04386(.A(new_n4762), .B(new_n4757), .Y(new_n4763));
  nor_5  g04387(.A(new_n4763), .B(new_n4751), .Y(new_n4764));
  xor_4  g04388(.A(new_n4718), .B(new_n4717), .Y(new_n4765));
  xor_4  g04389(.A(new_n4763), .B(new_n4750), .Y(new_n4766));
  nor_5  g04390(.A(new_n4766), .B(new_n4765), .Y(new_n4767));
  nor_5  g04391(.A(new_n4767), .B(new_n4764), .Y(new_n4768));
  xnor_4 g04392(.A(new_n4768), .B(new_n4749), .Y(new_n4769));
  nor_5  g04393(.A(new_n4769), .B(new_n4667), .Y(new_n4770));
  xnor_4 g04394(.A(new_n4766), .B(new_n4765), .Y(new_n4771));
  xor_4  g04395(.A(new_n4654), .B(new_n4650), .Y(new_n4772));
  nor_5  g04396(.A(new_n4772), .B(new_n4771), .Y(new_n4773));
  not_8  g04397(.A(new_n4773), .Y(new_n4774));
  nor_5  g04398(.A(new_n3560), .B(new_n3559), .Y(new_n4775));
  xor_4  g04399(.A(new_n4653), .B(new_n4652), .Y(new_n4776));
  nor_5  g04400(.A(new_n4776), .B(new_n4775), .Y(new_n4777));
  xor_4  g04401(.A(new_n4761), .B(new_n4758), .Y(new_n4778));
  not_8  g04402(.A(new_n4778), .Y(new_n4779));
  xor_4  g04403(.A(new_n4776), .B(new_n4775), .Y(new_n4780));
  nand_5 g04404(.A(new_n4780), .B(new_n4779), .Y(new_n4781));
  not_8  g04405(.A(new_n4781), .Y(new_n4782));
  nor_5  g04406(.A(new_n4782), .B(new_n4777), .Y(new_n4783));
  xor_4  g04407(.A(new_n4772), .B(new_n4771), .Y(new_n4784));
  nand_5 g04408(.A(new_n4784), .B(new_n4783), .Y(new_n4785));
  nand_5 g04409(.A(new_n4785), .B(new_n4774), .Y(new_n4786));
  xnor_4 g04410(.A(new_n4769), .B(new_n4667), .Y(new_n4787));
  nor_5  g04411(.A(new_n4787), .B(new_n4786), .Y(new_n4788));
  nor_5  g04412(.A(new_n4788), .B(new_n4770), .Y(new_n4789));
  nor_5  g04413(.A(new_n4666), .B(new_n4655), .Y(new_n4790));
  nor_5  g04414(.A(new_n4664), .B(new_n4661), .Y(new_n4791));
  not_8  g04415(.A(new_n4665), .Y(new_n4792));
  nor_5  g04416(.A(new_n4792), .B(new_n4660), .Y(new_n4793));
  nor_5  g04417(.A(new_n4793), .B(new_n4791), .Y(new_n4794));
  nand_5 g04418(.A(pi180), .B(pi131), .Y(new_n4795));
  nand_5 g04419(.A(pi133), .B(pi057), .Y(new_n4796));
  nand_5 g04420(.A(pi189), .B(pi143), .Y(new_n4797));
  nand_5 g04421(.A(pi194), .B(pi077), .Y(new_n4798));
  xor_4  g04422(.A(new_n4798), .B(new_n4797), .Y(new_n4799));
  xor_4  g04423(.A(new_n4799), .B(new_n4796), .Y(new_n4800));
  nand_5 g04424(.A(pi085), .B(pi052), .Y(new_n4801));
  nand_5 g04425(.A(new_n4658), .B(new_n4657), .Y(new_n4802));
  nand_5 g04426(.A(new_n4659), .B(new_n4656), .Y(new_n4803));
  nand_5 g04427(.A(new_n4803), .B(new_n4802), .Y(new_n4804));
  xor_4  g04428(.A(new_n4804), .B(new_n4801), .Y(new_n4805));
  xor_4  g04429(.A(new_n4805), .B(new_n4800), .Y(new_n4806));
  xnor_4 g04430(.A(new_n4806), .B(new_n4795), .Y(new_n4807));
  xor_4  g04431(.A(new_n4807), .B(new_n4794), .Y(new_n4808));
  xor_4  g04432(.A(new_n4808), .B(new_n4790), .Y(new_n4809));
  not_8  g04433(.A(new_n4745), .Y(new_n4810));
  nor_5  g04434(.A(new_n4810), .B(new_n4734), .Y(new_n4811));
  not_8  g04435(.A(new_n4811), .Y(new_n4812));
  nand_5 g04436(.A(pi188), .B(pi112), .Y(new_n4813));
  nand_5 g04437(.A(pi104), .B(pi061), .Y(new_n4814));
  nand_5 g04438(.A(pi178), .B(pi013), .Y(new_n4815));
  xor_4  g04439(.A(new_n4815), .B(new_n4814), .Y(new_n4816));
  xor_4  g04440(.A(new_n4816), .B(new_n4813), .Y(new_n4817));
  nand_5 g04441(.A(pi212), .B(pi012), .Y(new_n4818));
  nand_5 g04442(.A(new_n4737), .B(new_n4736), .Y(new_n4819));
  nand_5 g04443(.A(new_n4738), .B(new_n4735), .Y(new_n4820));
  nand_5 g04444(.A(new_n4820), .B(new_n4819), .Y(new_n4821));
  xor_4  g04445(.A(new_n4821), .B(new_n4818), .Y(new_n4822));
  xor_4  g04446(.A(new_n4822), .B(new_n4817), .Y(new_n4823));
  nand_5 g04447(.A(pi213), .B(pi144), .Y(new_n4824));
  nand_5 g04448(.A(new_n4743), .B(new_n4740), .Y(new_n4825));
  nand_5 g04449(.A(new_n4744), .B(new_n4739), .Y(new_n4826));
  nand_5 g04450(.A(new_n4826), .B(new_n4825), .Y(new_n4827));
  xor_4  g04451(.A(new_n4827), .B(new_n4824), .Y(new_n4828));
  xor_4  g04452(.A(new_n4828), .B(new_n4823), .Y(new_n4829));
  xor_4  g04453(.A(new_n4829), .B(new_n4812), .Y(new_n4830));
  not_8  g04454(.A(new_n4721), .Y(new_n4831));
  nor_5  g04455(.A(new_n4732), .B(new_n4831), .Y(new_n4832));
  nand_5 g04456(.A(pi236), .B(pi118), .Y(new_n4833));
  nor_5  g04457(.A(new_n4730), .B(new_n4727), .Y(new_n4834));
  nor_5  g04458(.A(new_n4731), .B(new_n4726), .Y(new_n4835));
  nor_5  g04459(.A(new_n4835), .B(new_n4834), .Y(new_n4836));
  xor_4  g04460(.A(new_n4836), .B(new_n4833), .Y(new_n4837));
  nand_5 g04461(.A(pi161), .B(pi108), .Y(new_n4838));
  nand_5 g04462(.A(pi141), .B(pi042), .Y(new_n4839));
  nand_5 g04463(.A(pi090), .B(pi051), .Y(new_n4840));
  xor_4  g04464(.A(new_n4840), .B(new_n4839), .Y(new_n4841));
  xor_4  g04465(.A(new_n4841), .B(new_n4838), .Y(new_n4842));
  nand_5 g04466(.A(pi241), .B(pi007), .Y(new_n4843));
  nand_5 g04467(.A(new_n4724), .B(new_n4723), .Y(new_n4844));
  nand_5 g04468(.A(new_n4725), .B(new_n4722), .Y(new_n4845));
  nand_5 g04469(.A(new_n4845), .B(new_n4844), .Y(new_n4846));
  xor_4  g04470(.A(new_n4846), .B(new_n4843), .Y(new_n4847));
  xor_4  g04471(.A(new_n4847), .B(new_n4842), .Y(new_n4848));
  not_8  g04472(.A(new_n4848), .Y(new_n4849));
  xor_4  g04473(.A(new_n4849), .B(new_n4837), .Y(new_n4850));
  xor_4  g04474(.A(new_n4850), .B(new_n4832), .Y(new_n4851));
  xnor_4 g04475(.A(new_n4851), .B(new_n4830), .Y(new_n4852));
  nor_5  g04476(.A(new_n4746), .B(new_n4733), .Y(new_n4853));
  not_8  g04477(.A(new_n4747), .Y(new_n4854));
  nor_5  g04478(.A(new_n4854), .B(new_n4720), .Y(new_n4855));
  nor_5  g04479(.A(new_n4855), .B(new_n4853), .Y(new_n4856));
  xnor_4 g04480(.A(new_n4856), .B(new_n4852), .Y(new_n4857));
  nor_5  g04481(.A(new_n4685), .B(new_n4674), .Y(new_n4858));
  nand_5 g04482(.A(pi237), .B(pi168), .Y(new_n4859));
  nor_5  g04483(.A(new_n4683), .B(new_n4680), .Y(new_n4860));
  not_8  g04484(.A(new_n4684), .Y(new_n4861));
  nor_5  g04485(.A(new_n4861), .B(new_n4679), .Y(new_n4862));
  nor_5  g04486(.A(new_n4862), .B(new_n4860), .Y(new_n4863));
  xor_4  g04487(.A(new_n4863), .B(new_n4859), .Y(new_n4864));
  nand_5 g04488(.A(pi179), .B(pi139), .Y(new_n4865));
  nand_5 g04489(.A(pi035), .B(pi033), .Y(new_n4866));
  nand_5 g04490(.A(pi162), .B(pi015), .Y(new_n4867));
  xor_4  g04491(.A(new_n4867), .B(new_n4866), .Y(new_n4868));
  xor_4  g04492(.A(new_n4868), .B(new_n4865), .Y(new_n4869));
  nand_5 g04493(.A(pi208), .B(pi048), .Y(new_n4870));
  nand_5 g04494(.A(new_n4677), .B(new_n4676), .Y(new_n4871));
  nand_5 g04495(.A(new_n4678), .B(new_n4675), .Y(new_n4872));
  nand_5 g04496(.A(new_n4872), .B(new_n4871), .Y(new_n4873));
  xor_4  g04497(.A(new_n4873), .B(new_n4870), .Y(new_n4874));
  xor_4  g04498(.A(new_n4874), .B(new_n4869), .Y(new_n4875));
  not_8  g04499(.A(new_n4875), .Y(new_n4876));
  xor_4  g04500(.A(new_n4876), .B(new_n4864), .Y(new_n4877));
  xor_4  g04501(.A(new_n4877), .B(new_n4858), .Y(new_n4878));
  nand_5 g04502(.A(new_n4748), .B(new_n4687), .Y(new_n4879));
  nand_5 g04503(.A(new_n4768), .B(new_n4749), .Y(new_n4880));
  and_6  g04504(.A(new_n4880), .B(new_n4879), .Y(new_n4881));
  xor_4  g04505(.A(new_n4881), .B(new_n4878), .Y(new_n4882));
  xnor_4 g04506(.A(new_n4882), .B(new_n4857), .Y(new_n4883));
  xor_4  g04507(.A(new_n4883), .B(new_n4809), .Y(new_n4884));
  xor_4  g04508(.A(new_n4884), .B(new_n4789), .Y(po015));
  nand_5 g04509(.A(pi162), .B(pi041), .Y(new_n4886));
  nand_5 g04510(.A(pi182), .B(pi033), .Y(new_n4887));
  nand_5 g04511(.A(pi179), .B(pi138), .Y(new_n4888));
  xor_4  g04512(.A(new_n4888), .B(new_n4887), .Y(new_n4889));
  xor_4  g04513(.A(new_n4889), .B(new_n4886), .Y(new_n4890));
  nand_5 g04514(.A(pi138), .B(pi033), .Y(new_n4891));
  nand_5 g04515(.A(pi182), .B(pi162), .Y(new_n4892));
  nor_5  g04516(.A(new_n4892), .B(new_n4891), .Y(new_n4893));
  not_8  g04517(.A(new_n4893), .Y(new_n4894));
  nor_5  g04518(.A(new_n4894), .B(new_n4890), .Y(new_n4895));
  nand_5 g04519(.A(pi182), .B(pi179), .Y(new_n4896));
  nand_5 g04520(.A(pi041), .B(pi033), .Y(new_n4897));
  nand_5 g04521(.A(pi216), .B(pi162), .Y(new_n4898));
  xor_4  g04522(.A(new_n4898), .B(new_n4897), .Y(new_n4899));
  xor_4  g04523(.A(new_n4899), .B(new_n4896), .Y(new_n4900));
  nand_5 g04524(.A(pi138), .B(pi048), .Y(new_n4901));
  nand_5 g04525(.A(new_n4888), .B(new_n4887), .Y(new_n4902));
  nand_5 g04526(.A(new_n4889), .B(new_n4886), .Y(new_n4903));
  nand_5 g04527(.A(new_n4903), .B(new_n4902), .Y(new_n4904));
  xor_4  g04528(.A(new_n4904), .B(new_n4901), .Y(new_n4905));
  xnor_4 g04529(.A(new_n4905), .B(new_n4900), .Y(new_n4906));
  xor_4  g04530(.A(new_n4906), .B(new_n4895), .Y(new_n4907));
  nand_5 g04531(.A(pi108), .B(pi087), .Y(new_n4908));
  nand_5 g04532(.A(pi102), .B(pi051), .Y(new_n4909));
  nor_5  g04533(.A(new_n4909), .B(new_n4908), .Y(new_n4910));
  nand_5 g04534(.A(new_n4909), .B(new_n4908), .Y(new_n4911));
  nand_5 g04535(.A(pi219), .B(pi042), .Y(new_n4912));
  not_8  g04536(.A(new_n4912), .Y(new_n4913));
  nand_5 g04537(.A(pi087), .B(pi051), .Y(new_n4914));
  and_6  g04538(.A(new_n4914), .B(new_n4913), .Y(new_n4915));
  nor_5  g04539(.A(new_n4915), .B(new_n4911), .Y(new_n4916));
  nor_5  g04540(.A(new_n4916), .B(new_n4910), .Y(new_n4917));
  nand_5 g04541(.A(new_n4915), .B(new_n4911), .Y(new_n4918));
  nand_5 g04542(.A(new_n4918), .B(new_n4917), .Y(new_n4919));
  nand_5 g04543(.A(pi087), .B(pi042), .Y(new_n4920));
  nand_5 g04544(.A(pi219), .B(pi051), .Y(new_n4921));
  xor_4  g04545(.A(new_n4921), .B(new_n4920), .Y(new_n4922));
  nand_5 g04546(.A(pi178), .B(pi142), .Y(new_n4923));
  nand_5 g04547(.A(pi188), .B(pi071), .Y(new_n4924));
  xor_4  g04548(.A(new_n4924), .B(new_n4923), .Y(new_n4925));
  nor_5  g04549(.A(new_n4925), .B(new_n4922), .Y(new_n4926));
  nand_5 g04550(.A(pi188), .B(pi142), .Y(new_n4927));
  nor_5  g04551(.A(new_n4927), .B(new_n4914), .Y(new_n4928));
  xnor_4 g04552(.A(new_n4925), .B(new_n4922), .Y(new_n4929));
  nor_5  g04553(.A(new_n4929), .B(new_n4928), .Y(new_n4930));
  or_6   g04554(.A(new_n4930), .B(new_n4926), .Y(new_n4931));
  not_8  g04555(.A(new_n4927), .Y(new_n4932));
  nand_5 g04556(.A(pi178), .B(pi071), .Y(new_n4933));
  nor_5  g04557(.A(new_n4933), .B(new_n4932), .Y(new_n4934));
  nand_5 g04558(.A(pi188), .B(pi169), .Y(new_n4935));
  nand_5 g04559(.A(pi142), .B(pi061), .Y(new_n4936));
  or_6   g04560(.A(new_n4936), .B(new_n4935), .Y(new_n4937));
  nand_5 g04561(.A(new_n4936), .B(new_n4935), .Y(new_n4938));
  and_6  g04562(.A(new_n4938), .B(new_n4937), .Y(new_n4939));
  or_6   g04563(.A(new_n4939), .B(new_n4934), .Y(new_n4940));
  nand_5 g04564(.A(new_n4938), .B(new_n4934), .Y(new_n4941));
  nand_5 g04565(.A(new_n4941), .B(new_n4940), .Y(new_n4942));
  xnor_4 g04566(.A(new_n4942), .B(new_n4931), .Y(new_n4943));
  xnor_4 g04567(.A(new_n4943), .B(new_n4919), .Y(new_n4944));
  xor_4  g04568(.A(new_n4893), .B(new_n4890), .Y(new_n4945));
  or_6   g04569(.A(new_n4945), .B(new_n4944), .Y(new_n4946));
  xor_4  g04570(.A(new_n4945), .B(new_n4944), .Y(new_n4947));
  and_6  g04571(.A(pi162), .B(pi138), .Y(new_n4948));
  xor_4  g04572(.A(new_n4927), .B(new_n4914), .Y(new_n4949));
  and_6  g04573(.A(new_n4949), .B(new_n4948), .Y(new_n4950));
  xor_4  g04574(.A(new_n4892), .B(new_n4891), .Y(new_n4951));
  nor_5  g04575(.A(new_n4951), .B(new_n4950), .Y(new_n4952));
  xnor_4 g04576(.A(new_n4951), .B(new_n4950), .Y(new_n4953));
  xnor_4 g04577(.A(new_n4929), .B(new_n4928), .Y(new_n4954));
  nor_5  g04578(.A(new_n4954), .B(new_n4953), .Y(new_n4955));
  nor_5  g04579(.A(new_n4955), .B(new_n4952), .Y(new_n4956));
  nand_5 g04580(.A(new_n4956), .B(new_n4947), .Y(new_n4957));
  nand_5 g04581(.A(new_n4957), .B(new_n4946), .Y(new_n4958));
  xor_4  g04582(.A(new_n4958), .B(new_n4907), .Y(new_n4959));
  nor_5  g04583(.A(new_n4917), .B(new_n4912), .Y(new_n4960));
  nand_5 g04584(.A(pi051), .B(pi001), .Y(new_n4961));
  nand_5 g04585(.A(pi219), .B(pi108), .Y(new_n4962));
  nand_5 g04586(.A(pi102), .B(pi042), .Y(new_n4963));
  xor_4  g04587(.A(new_n4963), .B(new_n4962), .Y(new_n4964));
  xor_4  g04588(.A(new_n4964), .B(new_n4961), .Y(new_n4965));
  nand_5 g04589(.A(pi087), .B(pi007), .Y(new_n4966));
  or_6   g04590(.A(new_n4913), .B(new_n4910), .Y(new_n4967));
  nand_5 g04591(.A(new_n4967), .B(new_n4911), .Y(new_n4968));
  xor_4  g04592(.A(new_n4968), .B(new_n4966), .Y(new_n4969));
  xor_4  g04593(.A(new_n4969), .B(new_n4965), .Y(new_n4970));
  xor_4  g04594(.A(new_n4970), .B(new_n4960), .Y(new_n4971));
  nor_5  g04595(.A(new_n4940), .B(new_n4933), .Y(new_n4972));
  nand_5 g04596(.A(new_n4933), .B(new_n4937), .Y(new_n4973));
  nand_5 g04597(.A(new_n4973), .B(new_n4938), .Y(new_n4974));
  nand_5 g04598(.A(pi142), .B(pi012), .Y(new_n4975));
  xor_4  g04599(.A(new_n4975), .B(new_n4974), .Y(new_n4976));
  nand_5 g04600(.A(pi188), .B(pi123), .Y(new_n4977));
  nand_5 g04601(.A(pi071), .B(pi061), .Y(new_n4978));
  nand_5 g04602(.A(pi178), .B(pi169), .Y(new_n4979));
  xor_4  g04603(.A(new_n4979), .B(new_n4978), .Y(new_n4980));
  xor_4  g04604(.A(new_n4980), .B(new_n4977), .Y(new_n4981));
  xor_4  g04605(.A(new_n4981), .B(new_n4976), .Y(new_n4982));
  xor_4  g04606(.A(new_n4982), .B(new_n4972), .Y(new_n4983));
  xor_4  g04607(.A(new_n4983), .B(new_n4971), .Y(new_n4984));
  nor_5  g04608(.A(new_n4942), .B(new_n4931), .Y(new_n4985));
  nor_5  g04609(.A(new_n4943), .B(new_n4919), .Y(new_n4986));
  or_6   g04610(.A(new_n4986), .B(new_n4985), .Y(new_n4987));
  xnor_4 g04611(.A(new_n4987), .B(new_n4984), .Y(new_n4988));
  xnor_4 g04612(.A(new_n4988), .B(new_n4959), .Y(new_n4989));
  nand_5 g04613(.A(pi143), .B(pi060), .Y(new_n4990));
  nand_5 g04614(.A(pi057), .B(pi020), .Y(new_n4991));
  nand_5 g04615(.A(pi194), .B(pi160), .Y(new_n4992));
  xor_4  g04616(.A(new_n4992), .B(new_n4991), .Y(new_n4993));
  xor_4  g04617(.A(new_n4993), .B(new_n4990), .Y(new_n4994));
  nand_5 g04618(.A(pi160), .B(pi143), .Y(new_n4995));
  nor_5  g04619(.A(new_n4995), .B(new_n4991), .Y(new_n4996));
  not_8  g04620(.A(new_n4996), .Y(new_n4997));
  xor_4  g04621(.A(new_n4997), .B(new_n4994), .Y(new_n4998));
  not_8  g04622(.A(new_n4998), .Y(new_n4999));
  xnor_4 g04623(.A(new_n4949), .B(new_n4948), .Y(new_n5000));
  nor_5  g04624(.A(new_n5000), .B(new_n4995), .Y(new_n5001));
  not_8  g04625(.A(new_n5001), .Y(new_n5002));
  nand_5 g04626(.A(pi160), .B(pi057), .Y(new_n5003));
  nand_5 g04627(.A(pi143), .B(pi020), .Y(new_n5004));
  nand_5 g04628(.A(new_n5004), .B(new_n5003), .Y(new_n5005));
  nand_5 g04629(.A(new_n5005), .B(new_n4997), .Y(new_n5006));
  nor_5  g04630(.A(new_n5006), .B(new_n5002), .Y(new_n5007));
  xor_4  g04631(.A(new_n4954), .B(new_n4953), .Y(new_n5008));
  xor_4  g04632(.A(new_n5006), .B(new_n5001), .Y(new_n5009));
  nor_5  g04633(.A(new_n5009), .B(new_n5008), .Y(new_n5010));
  nor_5  g04634(.A(new_n5010), .B(new_n5007), .Y(new_n5011));
  nand_5 g04635(.A(new_n5011), .B(new_n4999), .Y(new_n5012));
  xor_4  g04636(.A(new_n5011), .B(new_n4999), .Y(new_n5013));
  xnor_4 g04637(.A(new_n4956), .B(new_n4947), .Y(new_n5014));
  nand_5 g04638(.A(new_n5014), .B(new_n5013), .Y(new_n5015));
  nand_5 g04639(.A(new_n5015), .B(new_n5012), .Y(new_n5016));
  or_6   g04640(.A(new_n4997), .B(new_n4994), .Y(new_n5017));
  not_8  g04641(.A(new_n5017), .Y(new_n5018));
  nand_5 g04642(.A(pi194), .B(pi020), .Y(new_n5019));
  nand_5 g04643(.A(pi223), .B(pi143), .Y(new_n5020));
  nand_5 g04644(.A(pi060), .B(pi057), .Y(new_n5021));
  xor_4  g04645(.A(new_n5021), .B(new_n5020), .Y(new_n5022));
  xor_4  g04646(.A(new_n5022), .B(new_n5019), .Y(new_n5023));
  nand_5 g04647(.A(pi160), .B(pi085), .Y(new_n5024));
  nand_5 g04648(.A(new_n4992), .B(new_n4991), .Y(new_n5025));
  nand_5 g04649(.A(new_n4993), .B(new_n4990), .Y(new_n5026));
  nand_5 g04650(.A(new_n5026), .B(new_n5025), .Y(new_n5027));
  xor_4  g04651(.A(new_n5027), .B(new_n5024), .Y(new_n5028));
  xor_4  g04652(.A(new_n5028), .B(new_n5023), .Y(new_n5029));
  xor_4  g04653(.A(new_n5029), .B(new_n5018), .Y(new_n5030));
  xor_4  g04654(.A(new_n5030), .B(new_n5016), .Y(new_n5031));
  xor_4  g04655(.A(new_n5031), .B(new_n4989), .Y(po016));
  nand_5 g04656(.A(pi103), .B(pi029), .Y(new_n5033));
  nand_5 g04657(.A(pi175), .B(pi132), .Y(new_n5034));
  nand_5 g04658(.A(pi226), .B(pi163), .Y(new_n5035));
  nand_5 g04659(.A(pi109), .B(pi107), .Y(new_n5036));
  xor_4  g04660(.A(new_n5036), .B(new_n5035), .Y(new_n5037));
  xor_4  g04661(.A(new_n5037), .B(new_n5034), .Y(new_n5038));
  nor_5  g04662(.A(new_n5038), .B(new_n5033), .Y(new_n5039));
  nand_5 g04663(.A(pi117), .B(pi029), .Y(new_n5040));
  nand_5 g04664(.A(pi103), .B(pi069), .Y(new_n5041));
  xor_4  g04665(.A(new_n5041), .B(new_n5040), .Y(new_n5042));
  xor_4  g04666(.A(new_n5042), .B(new_n5039), .Y(new_n5043));
  not_8  g04667(.A(new_n5037), .Y(new_n5044));
  or_6   g04668(.A(new_n5044), .B(new_n5034), .Y(new_n5045));
  nand_5 g04669(.A(pi186), .B(pi134), .Y(new_n5046));
  nor_5  g04670(.A(new_n5046), .B(new_n5034), .Y(new_n5047));
  nand_5 g04671(.A(pi186), .B(pi175), .Y(new_n5048));
  nand_5 g04672(.A(pi134), .B(pi132), .Y(new_n5049));
  and_6  g04673(.A(new_n5049), .B(new_n5048), .Y(new_n5050));
  or_6   g04674(.A(new_n5050), .B(new_n5047), .Y(new_n5051));
  xor_4  g04675(.A(new_n5051), .B(new_n5045), .Y(new_n5052));
  nand_5 g04676(.A(pi171), .B(pi014), .Y(new_n5053));
  or_6   g04677(.A(new_n5053), .B(new_n5036), .Y(new_n5054));
  nand_5 g04678(.A(pi107), .B(pi014), .Y(new_n5055));
  nand_5 g04679(.A(pi171), .B(pi109), .Y(new_n5056));
  nand_5 g04680(.A(new_n5056), .B(new_n5055), .Y(new_n5057));
  nand_5 g04681(.A(new_n5057), .B(new_n5054), .Y(new_n5058));
  or_6   g04682(.A(new_n5036), .B(new_n5035), .Y(new_n5059));
  nand_5 g04683(.A(pi207), .B(pi148), .Y(new_n5060));
  or_6   g04684(.A(new_n5060), .B(new_n5035), .Y(new_n5061));
  nand_5 g04685(.A(pi226), .B(pi148), .Y(new_n5062));
  nand_5 g04686(.A(pi207), .B(pi163), .Y(new_n5063));
  nand_5 g04687(.A(new_n5063), .B(new_n5062), .Y(new_n5064));
  nand_5 g04688(.A(new_n5064), .B(new_n5061), .Y(new_n5065));
  xnor_4 g04689(.A(new_n5065), .B(new_n5059), .Y(new_n5066));
  xnor_4 g04690(.A(new_n5066), .B(new_n5058), .Y(new_n5067));
  xor_4  g04691(.A(new_n5067), .B(new_n5052), .Y(new_n5068));
  not_8  g04692(.A(new_n5068), .Y(new_n5069));
  xor_4  g04693(.A(new_n5069), .B(new_n5043), .Y(po017));
  xor_4  g04694(.A(new_n3014), .B(new_n3013), .Y(po018));
  nor_5  g04695(.A(new_n3260), .B(new_n3210), .Y(new_n5072));
  nor_5  g04696(.A(new_n3258), .B(new_n3256), .Y(new_n5073));
  not_8  g04697(.A(new_n3259), .Y(new_n5074));
  nor_5  g04698(.A(new_n5074), .B(new_n3255), .Y(new_n5075));
  nor_5  g04699(.A(new_n5075), .B(new_n5073), .Y(new_n5076));
  nand_5 g04700(.A(pi236), .B(pi050), .Y(new_n5077));
  nand_5 g04701(.A(pi173), .B(pi161), .Y(new_n5078));
  nand_5 g04702(.A(pi109), .B(pi090), .Y(new_n5079));
  nand_5 g04703(.A(pi141), .B(pi014), .Y(new_n5080));
  xor_4  g04704(.A(new_n5080), .B(new_n5079), .Y(new_n5081));
  xor_4  g04705(.A(new_n5081), .B(new_n5078), .Y(new_n5082));
  nand_5 g04706(.A(new_n3253), .B(new_n3252), .Y(new_n5083));
  nand_5 g04707(.A(new_n3254), .B(new_n3251), .Y(new_n5084));
  nand_5 g04708(.A(new_n5084), .B(new_n5083), .Y(new_n5085));
  nand_5 g04709(.A(pi241), .B(pi230), .Y(new_n5086));
  xor_4  g04710(.A(new_n5086), .B(new_n5085), .Y(new_n5087));
  xor_4  g04711(.A(new_n5087), .B(new_n5082), .Y(new_n5088));
  xnor_4 g04712(.A(new_n5088), .B(new_n5077), .Y(new_n5089));
  xor_4  g04713(.A(new_n5089), .B(new_n5076), .Y(new_n5090));
  nand_5 g04714(.A(new_n5090), .B(new_n5072), .Y(new_n5091));
  nand_5 g04715(.A(pi253), .B(pi236), .Y(new_n5092));
  nand_5 g04716(.A(new_n5092), .B(new_n5091), .Y(new_n5093));
  nor_5  g04717(.A(new_n5088), .B(new_n5077), .Y(new_n5094));
  or_6   g04718(.A(new_n5089), .B(new_n5076), .Y(new_n5095));
  not_8  g04719(.A(new_n5095), .Y(new_n5096));
  nor_5  g04720(.A(new_n5096), .B(new_n5094), .Y(new_n5097));
  nand_5 g04721(.A(pi230), .B(pi161), .Y(new_n5098));
  nand_5 g04722(.A(pi241), .B(pi050), .Y(new_n5099));
  and_6  g04723(.A(new_n5099), .B(new_n5098), .Y(new_n5100));
  nand_5 g04724(.A(pi161), .B(pi050), .Y(new_n5101));
  nor_5  g04725(.A(new_n5101), .B(new_n5086), .Y(new_n5102));
  or_6   g04726(.A(new_n5102), .B(new_n5100), .Y(new_n5103));
  nand_5 g04727(.A(new_n5080), .B(new_n5079), .Y(new_n5104));
  nand_5 g04728(.A(new_n5081), .B(new_n5078), .Y(new_n5105));
  nand_5 g04729(.A(new_n5105), .B(new_n5104), .Y(new_n5106));
  nand_5 g04730(.A(pi173), .B(pi141), .Y(new_n5107));
  nand_5 g04731(.A(pi047), .B(pi014), .Y(new_n5108));
  nor_5  g04732(.A(new_n5108), .B(new_n5079), .Y(new_n5109));
  not_8  g04733(.A(new_n5109), .Y(new_n5110));
  nand_5 g04734(.A(pi090), .B(pi014), .Y(new_n5111));
  nand_5 g04735(.A(pi109), .B(pi047), .Y(new_n5112));
  nand_5 g04736(.A(new_n5112), .B(new_n5111), .Y(new_n5113));
  nand_5 g04737(.A(new_n5113), .B(new_n5110), .Y(new_n5114));
  xor_4  g04738(.A(new_n5114), .B(new_n5107), .Y(new_n5115));
  xor_4  g04739(.A(new_n5115), .B(new_n5106), .Y(new_n5116));
  xor_4  g04740(.A(new_n5116), .B(new_n5103), .Y(new_n5117));
  nand_5 g04741(.A(new_n5086), .B(new_n5085), .Y(new_n5118));
  nand_5 g04742(.A(new_n5087), .B(new_n5082), .Y(new_n5119));
  nand_5 g04743(.A(new_n5119), .B(new_n5118), .Y(new_n5120));
  xor_4  g04744(.A(new_n5120), .B(new_n5117), .Y(new_n5121));
  xnor_4 g04745(.A(new_n5121), .B(new_n5097), .Y(new_n5122));
  not_8  g04746(.A(new_n5122), .Y(new_n5123));
  xnor_4 g04747(.A(new_n5092), .B(new_n5091), .Y(new_n5124));
  or_6   g04748(.A(new_n5124), .B(new_n5123), .Y(new_n5125));
  nand_5 g04749(.A(new_n5125), .B(new_n5093), .Y(new_n5126));
  or_6   g04750(.A(new_n5121), .B(new_n5097), .Y(new_n5127));
  nand_5 g04751(.A(pi230), .B(pi141), .Y(new_n5128));
  xor_4  g04752(.A(new_n5128), .B(new_n5109), .Y(new_n5129));
  nand_5 g04753(.A(pi173), .B(pi090), .Y(new_n5130));
  nand_5 g04754(.A(pi109), .B(pi018), .Y(new_n5131));
  xor_4  g04755(.A(new_n5131), .B(new_n5130), .Y(new_n5132));
  xor_4  g04756(.A(new_n5132), .B(new_n5108), .Y(new_n5133));
  xor_4  g04757(.A(new_n5133), .B(new_n5129), .Y(new_n5134));
  nand_5 g04758(.A(new_n5114), .B(new_n5107), .Y(new_n5135));
  nand_5 g04759(.A(new_n5115), .B(new_n5106), .Y(new_n5136));
  nand_5 g04760(.A(new_n5136), .B(new_n5135), .Y(new_n5137));
  nand_5 g04761(.A(pi253), .B(pi241), .Y(new_n5138));
  nand_5 g04762(.A(pi236), .B(pi074), .Y(new_n5139));
  xor_4  g04763(.A(new_n5139), .B(new_n5138), .Y(new_n5140));
  xor_4  g04764(.A(new_n5140), .B(new_n5101), .Y(new_n5141));
  xor_4  g04765(.A(new_n5141), .B(new_n5137), .Y(new_n5142));
  not_8  g04766(.A(new_n5142), .Y(new_n5143));
  xor_4  g04767(.A(new_n5143), .B(new_n5134), .Y(new_n5144));
  nor_5  g04768(.A(new_n5116), .B(new_n5103), .Y(new_n5145));
  not_8  g04769(.A(new_n5117), .Y(new_n5146));
  nor_5  g04770(.A(new_n5120), .B(new_n5146), .Y(new_n5147));
  xor_4  g04771(.A(new_n5147), .B(new_n5102), .Y(new_n5148));
  nor_5  g04772(.A(new_n5148), .B(new_n5145), .Y(new_n5149));
  xor_4  g04773(.A(new_n5149), .B(new_n5144), .Y(new_n5150));
  xor_4  g04774(.A(new_n5150), .B(new_n5127), .Y(new_n5151));
  xor_4  g04775(.A(new_n5151), .B(new_n5126), .Y(new_n5152));
  nand_5 g04776(.A(pi213), .B(pi025), .Y(new_n5153));
  nand_5 g04777(.A(pi213), .B(pi002), .Y(new_n5154));
  nand_5 g04778(.A(new_n3247), .B(new_n3244), .Y(new_n5155));
  nand_5 g04779(.A(new_n3248), .B(new_n3243), .Y(new_n5156));
  nand_5 g04780(.A(new_n5156), .B(new_n5155), .Y(new_n5157));
  nor_5  g04781(.A(new_n5157), .B(new_n5154), .Y(new_n5158));
  nand_5 g04782(.A(pi226), .B(pi112), .Y(new_n5159));
  nand_5 g04783(.A(pi207), .B(pi013), .Y(new_n5160));
  nand_5 g04784(.A(pi104), .B(pi066), .Y(new_n5161));
  xor_4  g04785(.A(new_n5161), .B(new_n5160), .Y(new_n5162));
  xor_4  g04786(.A(new_n5162), .B(new_n5159), .Y(new_n5163));
  nand_5 g04787(.A(new_n3241), .B(new_n3240), .Y(new_n5164));
  nand_5 g04788(.A(new_n3242), .B(new_n3239), .Y(new_n5165));
  nand_5 g04789(.A(new_n5165), .B(new_n5164), .Y(new_n5166));
  nand_5 g04790(.A(pi212), .B(pi055), .Y(new_n5167));
  xor_4  g04791(.A(new_n5167), .B(new_n5166), .Y(new_n5168));
  xor_4  g04792(.A(new_n5168), .B(new_n5163), .Y(new_n5169));
  xnor_4 g04793(.A(new_n5157), .B(new_n5154), .Y(new_n5170));
  nor_5  g04794(.A(new_n5170), .B(new_n5169), .Y(new_n5171));
  or_6   g04795(.A(new_n5171), .B(new_n5158), .Y(new_n5172));
  nand_5 g04796(.A(new_n5167), .B(new_n5166), .Y(new_n5173));
  nand_5 g04797(.A(new_n5168), .B(new_n5163), .Y(new_n5174));
  nand_5 g04798(.A(new_n5174), .B(new_n5173), .Y(new_n5175));
  nand_5 g04799(.A(pi104), .B(pi055), .Y(new_n5176));
  nand_5 g04800(.A(pi212), .B(pi002), .Y(new_n5177));
  and_6  g04801(.A(new_n5177), .B(new_n5176), .Y(new_n5178));
  nand_5 g04802(.A(pi104), .B(pi002), .Y(new_n5179));
  nor_5  g04803(.A(new_n5179), .B(new_n5167), .Y(new_n5180));
  or_6   g04804(.A(new_n5180), .B(new_n5178), .Y(new_n5181));
  nand_5 g04805(.A(pi066), .B(pi013), .Y(new_n5182));
  nand_5 g04806(.A(new_n5161), .B(new_n5160), .Y(new_n5183));
  nand_5 g04807(.A(new_n5162), .B(new_n5159), .Y(new_n5184));
  nand_5 g04808(.A(new_n5184), .B(new_n5183), .Y(new_n5185));
  nand_5 g04809(.A(pi207), .B(pi105), .Y(new_n5186));
  nor_5  g04810(.A(new_n5186), .B(new_n5159), .Y(new_n5187));
  not_8  g04811(.A(new_n5187), .Y(new_n5188));
  nand_5 g04812(.A(pi226), .B(pi105), .Y(new_n5189));
  nand_5 g04813(.A(pi207), .B(pi112), .Y(new_n5190));
  nand_5 g04814(.A(new_n5190), .B(new_n5189), .Y(new_n5191));
  nand_5 g04815(.A(new_n5191), .B(new_n5188), .Y(new_n5192));
  xor_4  g04816(.A(new_n5192), .B(new_n5185), .Y(new_n5193));
  xor_4  g04817(.A(new_n5193), .B(new_n5182), .Y(new_n5194));
  xor_4  g04818(.A(new_n5194), .B(new_n5181), .Y(new_n5195));
  not_8  g04819(.A(new_n5195), .Y(new_n5196));
  xor_4  g04820(.A(new_n5196), .B(new_n5175), .Y(new_n5197));
  xnor_4 g04821(.A(new_n5197), .B(new_n5172), .Y(new_n5198));
  or_6   g04822(.A(new_n5198), .B(new_n5153), .Y(new_n5199));
  xor_4  g04823(.A(new_n5198), .B(new_n5153), .Y(new_n5200));
  not_8  g04824(.A(new_n3249), .Y(new_n5201));
  nand_5 g04825(.A(new_n5201), .B(new_n3238), .Y(new_n5202));
  xnor_4 g04826(.A(new_n5170), .B(new_n5169), .Y(new_n5203));
  nor_5  g04827(.A(new_n5203), .B(new_n5202), .Y(new_n5204));
  nand_5 g04828(.A(new_n5204), .B(new_n5200), .Y(new_n5205));
  nand_5 g04829(.A(new_n5205), .B(new_n5199), .Y(new_n5206));
  nand_5 g04830(.A(new_n5197), .B(new_n5172), .Y(new_n5207));
  nor_5  g04831(.A(new_n5196), .B(new_n5175), .Y(new_n5208));
  nand_5 g04832(.A(new_n5208), .B(new_n5180), .Y(new_n5209));
  or_6   g04833(.A(new_n5196), .B(new_n5175), .Y(new_n5210));
  nor_5  g04834(.A(new_n5194), .B(new_n5181), .Y(new_n5211));
  nor_5  g04835(.A(new_n5211), .B(new_n5180), .Y(new_n5212));
  nand_5 g04836(.A(new_n5212), .B(new_n5210), .Y(new_n5213));
  nand_5 g04837(.A(new_n5213), .B(new_n5209), .Y(new_n5214));
  nand_5 g04838(.A(pi055), .B(pi013), .Y(new_n5215));
  xor_4  g04839(.A(new_n5215), .B(new_n5188), .Y(new_n5216));
  nand_5 g04840(.A(pi226), .B(pi183), .Y(new_n5217));
  nand_5 g04841(.A(pi112), .B(pi066), .Y(new_n5218));
  xor_4  g04842(.A(new_n5218), .B(new_n5217), .Y(new_n5219));
  xor_4  g04843(.A(new_n5219), .B(new_n5186), .Y(new_n5220));
  not_8  g04844(.A(new_n5220), .Y(new_n5221));
  xor_4  g04845(.A(new_n5221), .B(new_n5216), .Y(new_n5222));
  nand_5 g04846(.A(new_n5192), .B(new_n5185), .Y(new_n5223));
  nand_5 g04847(.A(new_n5193), .B(new_n5182), .Y(new_n5224));
  nand_5 g04848(.A(new_n5224), .B(new_n5223), .Y(new_n5225));
  nand_5 g04849(.A(pi212), .B(pi025), .Y(new_n5226));
  nand_5 g04850(.A(pi239), .B(pi213), .Y(new_n5227));
  xor_4  g04851(.A(new_n5227), .B(new_n5226), .Y(new_n5228));
  xnor_4 g04852(.A(new_n5228), .B(new_n5179), .Y(new_n5229));
  xor_4  g04853(.A(new_n5229), .B(new_n5225), .Y(new_n5230));
  xor_4  g04854(.A(new_n5230), .B(new_n5222), .Y(new_n5231));
  not_8  g04855(.A(new_n5231), .Y(new_n5232));
  xor_4  g04856(.A(new_n5232), .B(new_n5214), .Y(new_n5233));
  xor_4  g04857(.A(new_n5233), .B(new_n5207), .Y(new_n5234));
  xor_4  g04858(.A(new_n5234), .B(new_n5206), .Y(new_n5235));
  xnor_4 g04859(.A(new_n5235), .B(new_n5152), .Y(new_n5236));
  xor_4  g04860(.A(new_n5204), .B(new_n5200), .Y(new_n5237));
  xor_4  g04861(.A(new_n5124), .B(new_n5122), .Y(new_n5238));
  nand_5 g04862(.A(new_n5238), .B(new_n5237), .Y(new_n5239));
  xnor_4 g04863(.A(new_n5090), .B(new_n5072), .Y(new_n5240));
  xnor_4 g04864(.A(new_n5203), .B(new_n5202), .Y(new_n5241));
  nor_5  g04865(.A(new_n5241), .B(new_n5240), .Y(new_n5242));
  xnor_4 g04866(.A(new_n5241), .B(new_n5240), .Y(new_n5243));
  nand_5 g04867(.A(new_n3263), .B(new_n3237), .Y(new_n5244));
  nand_5 g04868(.A(new_n5244), .B(new_n3262), .Y(new_n5245));
  nor_5  g04869(.A(new_n5245), .B(new_n5243), .Y(new_n5246));
  nor_5  g04870(.A(new_n5246), .B(new_n5242), .Y(new_n5247));
  xnor_4 g04871(.A(new_n5238), .B(new_n5237), .Y(new_n5248));
  or_6   g04872(.A(new_n5248), .B(new_n5247), .Y(new_n5249));
  nand_5 g04873(.A(new_n5249), .B(new_n5239), .Y(new_n5250));
  xor_4  g04874(.A(new_n5250), .B(new_n5236), .Y(new_n5251));
  nand_5 g04875(.A(pi199), .B(pi168), .Y(new_n5252));
  nand_5 g04876(.A(pi139), .B(pi058), .Y(new_n5253));
  nand_5 g04877(.A(pi186), .B(pi035), .Y(new_n5254));
  nand_5 g04878(.A(pi132), .B(pi015), .Y(new_n5255));
  xor_4  g04879(.A(new_n5255), .B(new_n5254), .Y(new_n5256));
  xor_4  g04880(.A(new_n5256), .B(new_n5253), .Y(new_n5257));
  nand_5 g04881(.A(pi211), .B(pi208), .Y(new_n5258));
  nand_5 g04882(.A(new_n3222), .B(new_n3221), .Y(new_n5259));
  nand_5 g04883(.A(new_n3223), .B(new_n3220), .Y(new_n5260));
  nand_5 g04884(.A(new_n5260), .B(new_n5259), .Y(new_n5261));
  xor_4  g04885(.A(new_n5261), .B(new_n5258), .Y(new_n5262));
  xor_4  g04886(.A(new_n5262), .B(new_n5257), .Y(new_n5263));
  nor_5  g04887(.A(new_n5263), .B(new_n5252), .Y(new_n5264));
  nor_5  g04888(.A(new_n3229), .B(new_n3226), .Y(new_n5265));
  and_6  g04889(.A(new_n3230), .B(new_n3225), .Y(new_n5266));
  nor_5  g04890(.A(new_n5266), .B(new_n5265), .Y(new_n5267));
  xnor_4 g04891(.A(new_n5263), .B(new_n5252), .Y(new_n5268));
  nor_5  g04892(.A(new_n5268), .B(new_n5267), .Y(new_n5269));
  nor_5  g04893(.A(new_n5269), .B(new_n5264), .Y(new_n5270));
  nand_5 g04894(.A(pi211), .B(pi139), .Y(new_n5271));
  nand_5 g04895(.A(pi208), .B(pi199), .Y(new_n5272));
  and_6  g04896(.A(new_n5272), .B(new_n5271), .Y(new_n5273));
  nand_5 g04897(.A(pi199), .B(pi139), .Y(new_n5274));
  nor_5  g04898(.A(new_n5274), .B(new_n5258), .Y(new_n5275));
  or_6   g04899(.A(new_n5275), .B(new_n5273), .Y(new_n5276));
  nand_5 g04900(.A(new_n5255), .B(new_n5254), .Y(new_n5277));
  nand_5 g04901(.A(new_n5256), .B(new_n5253), .Y(new_n5278));
  nand_5 g04902(.A(new_n5278), .B(new_n5277), .Y(new_n5279));
  nand_5 g04903(.A(pi058), .B(pi035), .Y(new_n5280));
  nand_5 g04904(.A(pi186), .B(pi015), .Y(new_n5281));
  nand_5 g04905(.A(pi204), .B(pi132), .Y(new_n5282));
  nand_5 g04906(.A(new_n5282), .B(new_n5281), .Y(new_n5283));
  nand_5 g04907(.A(pi204), .B(pi186), .Y(new_n5284));
  nor_5  g04908(.A(new_n5284), .B(new_n5255), .Y(new_n5285));
  not_8  g04909(.A(new_n5285), .Y(new_n5286));
  nand_5 g04910(.A(new_n5286), .B(new_n5283), .Y(new_n5287));
  xor_4  g04911(.A(new_n5287), .B(new_n5280), .Y(new_n5288));
  xor_4  g04912(.A(new_n5288), .B(new_n5279), .Y(new_n5289));
  xor_4  g04913(.A(new_n5289), .B(new_n5276), .Y(new_n5290));
  nand_5 g04914(.A(new_n5261), .B(new_n5258), .Y(new_n5291));
  nand_5 g04915(.A(new_n5262), .B(new_n5257), .Y(new_n5292));
  nand_5 g04916(.A(new_n5292), .B(new_n5291), .Y(new_n5293));
  xor_4  g04917(.A(new_n5293), .B(new_n5290), .Y(new_n5294));
  nor_5  g04918(.A(new_n5294), .B(new_n5270), .Y(new_n5295));
  not_8  g04919(.A(new_n5295), .Y(new_n5296));
  nand_5 g04920(.A(new_n3231), .B(new_n3219), .Y(new_n5297));
  not_8  g04921(.A(new_n5297), .Y(new_n5298));
  xor_4  g04922(.A(new_n5268), .B(new_n5267), .Y(new_n5299));
  nand_5 g04923(.A(new_n5299), .B(new_n5298), .Y(new_n5300));
  nand_5 g04924(.A(pi195), .B(pi168), .Y(new_n5301));
  nand_5 g04925(.A(new_n5301), .B(new_n5300), .Y(new_n5302));
  not_8  g04926(.A(new_n5302), .Y(new_n5303));
  xor_4  g04927(.A(new_n5294), .B(new_n5270), .Y(new_n5304));
  xnor_4 g04928(.A(new_n5301), .B(new_n5300), .Y(new_n5305));
  nor_5  g04929(.A(new_n5305), .B(new_n5304), .Y(new_n5306));
  nor_5  g04930(.A(new_n5306), .B(new_n5303), .Y(new_n5307));
  nor_5  g04931(.A(new_n5289), .B(new_n5276), .Y(new_n5308));
  not_8  g04932(.A(new_n5290), .Y(new_n5309));
  nor_5  g04933(.A(new_n5293), .B(new_n5309), .Y(new_n5310));
  xor_4  g04934(.A(new_n5310), .B(new_n5275), .Y(new_n5311));
  nor_5  g04935(.A(new_n5311), .B(new_n5308), .Y(new_n5312));
  nand_5 g04936(.A(new_n5287), .B(new_n5280), .Y(new_n5313));
  nand_5 g04937(.A(new_n5288), .B(new_n5279), .Y(new_n5314));
  nand_5 g04938(.A(new_n5314), .B(new_n5313), .Y(new_n5315));
  nand_5 g04939(.A(pi208), .B(pi195), .Y(new_n5316));
  nand_5 g04940(.A(pi218), .B(pi168), .Y(new_n5317));
  xor_4  g04941(.A(new_n5317), .B(new_n5316), .Y(new_n5318));
  xnor_4 g04942(.A(new_n5318), .B(new_n5274), .Y(new_n5319));
  xor_4  g04943(.A(new_n5319), .B(new_n5315), .Y(new_n5320));
  nand_5 g04944(.A(pi211), .B(pi035), .Y(new_n5321));
  xor_4  g04945(.A(new_n5321), .B(new_n5285), .Y(new_n5322));
  nand_5 g04946(.A(pi146), .B(pi132), .Y(new_n5323));
  nand_5 g04947(.A(pi058), .B(pi015), .Y(new_n5324));
  xor_4  g04948(.A(new_n5324), .B(new_n5323), .Y(new_n5325));
  xor_4  g04949(.A(new_n5325), .B(new_n5284), .Y(new_n5326));
  xor_4  g04950(.A(new_n5326), .B(new_n5322), .Y(new_n5327));
  xnor_4 g04951(.A(new_n5327), .B(new_n5320), .Y(new_n5328));
  xor_4  g04952(.A(new_n5328), .B(new_n5312), .Y(new_n5329));
  not_8  g04953(.A(new_n5329), .Y(new_n5330));
  xor_4  g04954(.A(new_n5330), .B(new_n5307), .Y(new_n5331));
  xor_4  g04955(.A(new_n5331), .B(new_n5296), .Y(new_n5332));
  xor_4  g04956(.A(new_n5332), .B(new_n5251), .Y(new_n5333));
  xor_4  g04957(.A(new_n5305), .B(new_n5304), .Y(new_n5334));
  xnor_4 g04958(.A(new_n5248), .B(new_n5247), .Y(new_n5335));
  or_6   g04959(.A(new_n5335), .B(new_n5334), .Y(new_n5336));
  xor_4  g04960(.A(new_n5245), .B(new_n5243), .Y(new_n5337));
  xor_4  g04961(.A(new_n5299), .B(new_n5298), .Y(new_n5338));
  nand_5 g04962(.A(new_n5338), .B(new_n5337), .Y(new_n5339));
  nand_5 g04963(.A(new_n3232), .B(new_n3218), .Y(new_n5340));
  or_6   g04964(.A(new_n3265), .B(new_n3233), .Y(new_n5341));
  nand_5 g04965(.A(new_n5341), .B(new_n5340), .Y(new_n5342));
  xnor_4 g04966(.A(new_n5338), .B(new_n5337), .Y(new_n5343));
  or_6   g04967(.A(new_n5343), .B(new_n5342), .Y(new_n5344));
  nand_5 g04968(.A(new_n5344), .B(new_n5339), .Y(new_n5345));
  xor_4  g04969(.A(new_n5335), .B(new_n5334), .Y(new_n5346));
  nand_5 g04970(.A(new_n5346), .B(new_n5345), .Y(new_n5347));
  and_6  g04971(.A(new_n5347), .B(new_n5336), .Y(new_n5348));
  xnor_4 g04972(.A(new_n5348), .B(new_n5333), .Y(new_n5349));
  nand_5 g04973(.A(pi150), .B(pi077), .Y(new_n5350));
  nand_5 g04974(.A(pi221), .B(pi052), .Y(new_n5351));
  nand_5 g04975(.A(new_n5351), .B(new_n5350), .Y(new_n5352));
  nand_5 g04976(.A(pi221), .B(pi077), .Y(new_n5353));
  nand_5 g04977(.A(pi150), .B(pi052), .Y(new_n5354));
  nor_5  g04978(.A(new_n5354), .B(new_n5353), .Y(new_n5355));
  not_8  g04979(.A(new_n5355), .Y(new_n5356));
  nand_5 g04980(.A(new_n5356), .B(new_n5352), .Y(new_n5357));
  nand_5 g04981(.A(pi244), .B(pi077), .Y(new_n5358));
  nand_5 g04982(.A(pi133), .B(pi069), .Y(new_n5359));
  nand_5 g04983(.A(new_n5359), .B(new_n5358), .Y(new_n5360));
  nand_5 g04984(.A(pi189), .B(pi029), .Y(new_n5361));
  xor_4  g04985(.A(new_n5359), .B(new_n5358), .Y(new_n5362));
  nand_5 g04986(.A(new_n5362), .B(new_n5361), .Y(new_n5363));
  nand_5 g04987(.A(new_n5363), .B(new_n5360), .Y(new_n5364));
  nand_5 g04988(.A(pi244), .B(pi133), .Y(new_n5365));
  nand_5 g04989(.A(pi069), .B(pi064), .Y(new_n5366));
  nor_5  g04990(.A(new_n5366), .B(new_n5361), .Y(new_n5367));
  not_8  g04991(.A(new_n5367), .Y(new_n5368));
  nand_5 g04992(.A(pi189), .B(pi069), .Y(new_n5369));
  nand_5 g04993(.A(pi064), .B(pi029), .Y(new_n5370));
  nand_5 g04994(.A(new_n5370), .B(new_n5369), .Y(new_n5371));
  nand_5 g04995(.A(new_n5371), .B(new_n5368), .Y(new_n5372));
  xor_4  g04996(.A(new_n5372), .B(new_n5365), .Y(new_n5373));
  xor_4  g04997(.A(new_n5373), .B(new_n5364), .Y(new_n5374));
  nor_5  g04998(.A(new_n5374), .B(new_n5357), .Y(new_n5375));
  nand_5 g04999(.A(new_n3296), .B(new_n3295), .Y(new_n5376));
  nand_5 g05000(.A(new_n3297), .B(new_n3294), .Y(new_n5377));
  nand_5 g05001(.A(new_n5377), .B(new_n5376), .Y(new_n5378));
  nand_5 g05002(.A(new_n5378), .B(new_n5354), .Y(new_n5379));
  xor_4  g05003(.A(new_n5362), .B(new_n5361), .Y(new_n5380));
  xor_4  g05004(.A(new_n5378), .B(new_n5354), .Y(new_n5381));
  nand_5 g05005(.A(new_n5381), .B(new_n5380), .Y(new_n5382));
  nand_5 g05006(.A(new_n5382), .B(new_n5379), .Y(new_n5383));
  xnor_4 g05007(.A(new_n5374), .B(new_n5357), .Y(new_n5384));
  nor_5  g05008(.A(new_n5384), .B(new_n5383), .Y(new_n5385));
  xor_4  g05009(.A(new_n5385), .B(new_n5356), .Y(new_n5386));
  not_8  g05010(.A(new_n5386), .Y(new_n5387));
  nor_5  g05011(.A(new_n5387), .B(new_n5375), .Y(new_n5388));
  nand_5 g05012(.A(pi196), .B(pi052), .Y(new_n5389));
  nand_5 g05013(.A(pi184), .B(pi131), .Y(new_n5390));
  xor_4  g05014(.A(new_n5390), .B(new_n5389), .Y(new_n5391));
  xor_4  g05015(.A(new_n5391), .B(new_n5353), .Y(new_n5392));
  nand_5 g05016(.A(new_n5372), .B(new_n5365), .Y(new_n5393));
  nand_5 g05017(.A(new_n5373), .B(new_n5364), .Y(new_n5394));
  nand_5 g05018(.A(new_n5394), .B(new_n5393), .Y(new_n5395));
  xor_4  g05019(.A(new_n5395), .B(new_n5392), .Y(new_n5396));
  nand_5 g05020(.A(pi150), .B(pi133), .Y(new_n5397));
  xor_4  g05021(.A(new_n5397), .B(new_n5368), .Y(new_n5398));
  nand_5 g05022(.A(pi084), .B(pi029), .Y(new_n5399));
  nand_5 g05023(.A(pi244), .B(pi189), .Y(new_n5400));
  xor_4  g05024(.A(new_n5400), .B(new_n5399), .Y(new_n5401));
  xor_4  g05025(.A(new_n5401), .B(new_n5366), .Y(new_n5402));
  xor_4  g05026(.A(new_n5402), .B(new_n5398), .Y(new_n5403));
  xor_4  g05027(.A(new_n5403), .B(new_n5396), .Y(new_n5404));
  xor_4  g05028(.A(new_n5404), .B(new_n5388), .Y(new_n5405));
  xnor_4 g05029(.A(new_n5384), .B(new_n5383), .Y(new_n5406));
  nand_5 g05030(.A(pi221), .B(pi131), .Y(new_n5407));
  nand_5 g05031(.A(new_n3302), .B(new_n3299), .Y(new_n5408));
  nand_5 g05032(.A(new_n3303), .B(new_n3298), .Y(new_n5409));
  nand_5 g05033(.A(new_n5409), .B(new_n5408), .Y(new_n5410));
  nor_5  g05034(.A(new_n5410), .B(new_n5407), .Y(new_n5411));
  xor_4  g05035(.A(new_n5381), .B(new_n5380), .Y(new_n5412));
  xor_4  g05036(.A(new_n5410), .B(new_n5407), .Y(new_n5413));
  not_8  g05037(.A(new_n5413), .Y(new_n5414));
  nor_5  g05038(.A(new_n5414), .B(new_n5412), .Y(new_n5415));
  nor_5  g05039(.A(new_n5415), .B(new_n5411), .Y(new_n5416));
  nor_5  g05040(.A(new_n5416), .B(new_n5406), .Y(new_n5417));
  xor_4  g05041(.A(new_n5417), .B(new_n5405), .Y(new_n5418));
  nand_5 g05042(.A(pi196), .B(pi131), .Y(new_n5419));
  not_8  g05043(.A(new_n5419), .Y(new_n5420));
  or_6   g05044(.A(new_n3304), .B(new_n3293), .Y(new_n5421));
  xor_4  g05045(.A(new_n5413), .B(new_n5412), .Y(new_n5422));
  nor_5  g05046(.A(new_n5422), .B(new_n5421), .Y(new_n5423));
  nor_5  g05047(.A(new_n5423), .B(new_n5420), .Y(new_n5424));
  xor_4  g05048(.A(new_n5416), .B(new_n5406), .Y(new_n5425));
  xor_4  g05049(.A(new_n5423), .B(new_n5419), .Y(new_n5426));
  nor_5  g05050(.A(new_n5426), .B(new_n5425), .Y(new_n5427));
  nor_5  g05051(.A(new_n5427), .B(new_n5424), .Y(new_n5428));
  xor_4  g05052(.A(new_n5428), .B(new_n5418), .Y(new_n5429));
  xnor_4 g05053(.A(new_n5429), .B(new_n5349), .Y(new_n5430));
  or_6   g05054(.A(new_n3305), .B(new_n3292), .Y(new_n5431));
  nand_5 g05055(.A(new_n3306), .B(new_n3266), .Y(new_n5432));
  nand_5 g05056(.A(new_n5432), .B(new_n5431), .Y(new_n5433));
  xor_4  g05057(.A(new_n5422), .B(new_n5421), .Y(new_n5434));
  nor_5  g05058(.A(new_n5434), .B(new_n5433), .Y(new_n5435));
  xor_4  g05059(.A(new_n5343), .B(new_n5342), .Y(new_n5436));
  xnor_4 g05060(.A(new_n5434), .B(new_n5433), .Y(new_n5437));
  nor_5  g05061(.A(new_n5437), .B(new_n5436), .Y(new_n5438));
  nor_5  g05062(.A(new_n5438), .B(new_n5435), .Y(new_n5439));
  xor_4  g05063(.A(new_n5346), .B(new_n5345), .Y(new_n5440));
  nand_5 g05064(.A(new_n5440), .B(new_n5439), .Y(new_n5441));
  xor_4  g05065(.A(new_n5426), .B(new_n5425), .Y(new_n5442));
  xor_4  g05066(.A(new_n5440), .B(new_n5439), .Y(new_n5443));
  not_8  g05067(.A(new_n5443), .Y(new_n5444));
  or_6   g05068(.A(new_n5444), .B(new_n5442), .Y(new_n5445));
  nand_5 g05069(.A(new_n5445), .B(new_n5441), .Y(new_n5446));
  xnor_4 g05070(.A(new_n5446), .B(new_n5430), .Y(po019));
  xnor_4 g05071(.A(new_n3290), .B(new_n3289), .Y(po020));
  nand_5 g05072(.A(pi113), .B(pi087), .Y(new_n5449));
  nand_5 g05073(.A(pi219), .B(pi007), .Y(new_n5450));
  nand_5 g05074(.A(new_n4963), .B(new_n4962), .Y(new_n5451));
  nand_5 g05075(.A(new_n4964), .B(new_n4961), .Y(new_n5452));
  nand_5 g05076(.A(new_n5452), .B(new_n5451), .Y(new_n5453));
  nand_5 g05077(.A(new_n5453), .B(new_n5450), .Y(new_n5454));
  nand_5 g05078(.A(pi122), .B(pi051), .Y(new_n5455));
  nand_5 g05079(.A(pi108), .B(pi102), .Y(new_n5456));
  nand_5 g05080(.A(pi042), .B(pi001), .Y(new_n5457));
  xor_4  g05081(.A(new_n5457), .B(new_n5456), .Y(new_n5458));
  xor_4  g05082(.A(new_n5458), .B(new_n5455), .Y(new_n5459));
  xor_4  g05083(.A(new_n5453), .B(new_n5450), .Y(new_n5460));
  nand_5 g05084(.A(new_n5460), .B(new_n5459), .Y(new_n5461));
  nand_5 g05085(.A(new_n5461), .B(new_n5454), .Y(new_n5462));
  nand_5 g05086(.A(pi118), .B(pi102), .Y(new_n5463));
  nor_5  g05087(.A(new_n5463), .B(new_n5450), .Y(new_n5464));
  not_8  g05088(.A(new_n5464), .Y(new_n5465));
  nand_5 g05089(.A(pi219), .B(pi118), .Y(new_n5466));
  nand_5 g05090(.A(pi102), .B(pi007), .Y(new_n5467));
  nand_5 g05091(.A(new_n5467), .B(new_n5466), .Y(new_n5468));
  nand_5 g05092(.A(new_n5468), .B(new_n5465), .Y(new_n5469));
  nand_5 g05093(.A(new_n5457), .B(new_n5456), .Y(new_n5470));
  nand_5 g05094(.A(new_n5458), .B(new_n5455), .Y(new_n5471));
  nand_5 g05095(.A(new_n5471), .B(new_n5470), .Y(new_n5472));
  nand_5 g05096(.A(pi108), .B(pi001), .Y(new_n5473));
  nand_5 g05097(.A(pi122), .B(pi042), .Y(new_n5474));
  nand_5 g05098(.A(pi135), .B(pi051), .Y(new_n5475));
  nand_5 g05099(.A(new_n5475), .B(new_n5474), .Y(new_n5476));
  nand_5 g05100(.A(pi135), .B(pi042), .Y(new_n5477));
  nor_5  g05101(.A(new_n5477), .B(new_n5455), .Y(new_n5478));
  not_8  g05102(.A(new_n5478), .Y(new_n5479));
  and_6  g05103(.A(new_n5479), .B(new_n5476), .Y(new_n5480));
  xor_4  g05104(.A(new_n5480), .B(new_n5473), .Y(new_n5481));
  xor_4  g05105(.A(new_n5481), .B(new_n5472), .Y(new_n5482));
  xor_4  g05106(.A(new_n5482), .B(new_n5469), .Y(new_n5483));
  xor_4  g05107(.A(new_n5483), .B(new_n5462), .Y(new_n5484));
  nand_5 g05108(.A(pi118), .B(pi087), .Y(new_n5485));
  nor_5  g05109(.A(new_n4968), .B(new_n4966), .Y(new_n5486));
  not_8  g05110(.A(new_n4965), .Y(new_n5487));
  and_6  g05111(.A(new_n4969), .B(new_n5487), .Y(new_n5488));
  nor_5  g05112(.A(new_n5488), .B(new_n5486), .Y(new_n5489));
  nand_5 g05113(.A(new_n5489), .B(new_n5485), .Y(new_n5490));
  or_6   g05114(.A(new_n5489), .B(new_n5485), .Y(new_n5491));
  xor_4  g05115(.A(new_n5460), .B(new_n5459), .Y(new_n5492));
  nand_5 g05116(.A(new_n5492), .B(new_n5491), .Y(new_n5493));
  nand_5 g05117(.A(new_n5493), .B(new_n5490), .Y(new_n5494));
  xor_4  g05118(.A(new_n5494), .B(new_n5484), .Y(new_n5495));
  xor_4  g05119(.A(new_n5495), .B(new_n5449), .Y(new_n5496));
  not_8  g05120(.A(new_n4970), .Y(new_n5497));
  nand_5 g05121(.A(new_n5497), .B(new_n4960), .Y(new_n5498));
  nand_5 g05122(.A(new_n5491), .B(new_n5490), .Y(new_n5499));
  xnor_4 g05123(.A(new_n5499), .B(new_n5492), .Y(new_n5500));
  nor_5  g05124(.A(new_n5500), .B(new_n5498), .Y(new_n5501));
  xor_4  g05125(.A(new_n5501), .B(new_n5496), .Y(new_n5502));
  nand_5 g05126(.A(pi142), .B(pi098), .Y(new_n5503));
  not_8  g05127(.A(new_n4972), .Y(new_n5504));
  nor_5  g05128(.A(new_n4982), .B(new_n5504), .Y(new_n5505));
  not_8  g05129(.A(new_n5505), .Y(new_n5506));
  nand_5 g05130(.A(pi178), .B(pi123), .Y(new_n5507));
  nand_5 g05131(.A(pi188), .B(pi099), .Y(new_n5508));
  nand_5 g05132(.A(pi169), .B(pi061), .Y(new_n5509));
  xor_4  g05133(.A(new_n5509), .B(new_n5508), .Y(new_n5510));
  xor_4  g05134(.A(new_n5510), .B(new_n5507), .Y(new_n5511));
  nand_5 g05135(.A(pi071), .B(pi012), .Y(new_n5512));
  nand_5 g05136(.A(new_n4979), .B(new_n4978), .Y(new_n5513));
  nand_5 g05137(.A(new_n4980), .B(new_n4977), .Y(new_n5514));
  nand_5 g05138(.A(new_n5514), .B(new_n5513), .Y(new_n5515));
  xor_4  g05139(.A(new_n5515), .B(new_n5512), .Y(new_n5516));
  xor_4  g05140(.A(new_n5516), .B(new_n5511), .Y(new_n5517));
  nand_5 g05141(.A(pi144), .B(pi142), .Y(new_n5518));
  or_6   g05142(.A(new_n4975), .B(new_n4974), .Y(new_n5519));
  not_8  g05143(.A(new_n4981), .Y(new_n5520));
  nand_5 g05144(.A(new_n5520), .B(new_n4976), .Y(new_n5521));
  and_6  g05145(.A(new_n5521), .B(new_n5519), .Y(new_n5522));
  xnor_4 g05146(.A(new_n5522), .B(new_n5518), .Y(new_n5523));
  xnor_4 g05147(.A(new_n5523), .B(new_n5517), .Y(new_n5524));
  or_6   g05148(.A(new_n5524), .B(new_n5506), .Y(new_n5525));
  xor_4  g05149(.A(new_n5525), .B(new_n5503), .Y(new_n5526));
  nand_5 g05150(.A(new_n5515), .B(new_n5512), .Y(new_n5527));
  nand_5 g05151(.A(new_n5516), .B(new_n5511), .Y(new_n5528));
  nand_5 g05152(.A(new_n5528), .B(new_n5527), .Y(new_n5529));
  nand_5 g05153(.A(pi169), .B(pi012), .Y(new_n5530));
  nand_5 g05154(.A(pi144), .B(pi071), .Y(new_n5531));
  and_6  g05155(.A(new_n5531), .B(new_n5530), .Y(new_n5532));
  nand_5 g05156(.A(pi169), .B(pi144), .Y(new_n5533));
  nor_5  g05157(.A(new_n5512), .B(new_n5533), .Y(new_n5534));
  or_6   g05158(.A(new_n5534), .B(new_n5532), .Y(new_n5535));
  nand_5 g05159(.A(new_n5509), .B(new_n5508), .Y(new_n5536));
  nand_5 g05160(.A(new_n5510), .B(new_n5507), .Y(new_n5537));
  nand_5 g05161(.A(new_n5537), .B(new_n5536), .Y(new_n5538));
  nand_5 g05162(.A(pi123), .B(pi061), .Y(new_n5539));
  nand_5 g05163(.A(pi178), .B(pi099), .Y(new_n5540));
  nand_5 g05164(.A(pi188), .B(pi023), .Y(new_n5541));
  nand_5 g05165(.A(new_n5541), .B(new_n5540), .Y(new_n5542));
  nand_5 g05166(.A(pi178), .B(pi023), .Y(new_n5543));
  nor_5  g05167(.A(new_n5543), .B(new_n5508), .Y(new_n5544));
  not_8  g05168(.A(new_n5544), .Y(new_n5545));
  nand_5 g05169(.A(new_n5545), .B(new_n5542), .Y(new_n5546));
  xor_4  g05170(.A(new_n5546), .B(new_n5539), .Y(new_n5547));
  xor_4  g05171(.A(new_n5547), .B(new_n5538), .Y(new_n5548));
  xor_4  g05172(.A(new_n5548), .B(new_n5535), .Y(new_n5549));
  xor_4  g05173(.A(new_n5549), .B(new_n5529), .Y(new_n5550));
  nor_5  g05174(.A(new_n5522), .B(new_n5518), .Y(new_n5551));
  nor_5  g05175(.A(new_n5523), .B(new_n5517), .Y(new_n5552));
  nor_5  g05176(.A(new_n5552), .B(new_n5551), .Y(new_n5553));
  xor_4  g05177(.A(new_n5553), .B(new_n5550), .Y(new_n5554));
  xor_4  g05178(.A(new_n5554), .B(new_n5526), .Y(new_n5555));
  nand_5 g05179(.A(new_n5555), .B(new_n5502), .Y(new_n5556));
  xor_4  g05180(.A(new_n5555), .B(new_n5502), .Y(new_n5557));
  xor_4  g05181(.A(new_n5500), .B(new_n5498), .Y(new_n5558));
  xor_4  g05182(.A(new_n5524), .B(new_n5506), .Y(new_n5559));
  nor_5  g05183(.A(new_n5559), .B(new_n5558), .Y(new_n5560));
  xnor_4 g05184(.A(new_n5559), .B(new_n5558), .Y(new_n5561));
  or_6   g05185(.A(new_n4983), .B(new_n4971), .Y(new_n5562));
  nand_5 g05186(.A(new_n4987), .B(new_n4984), .Y(new_n5563));
  nand_5 g05187(.A(new_n5563), .B(new_n5562), .Y(new_n5564));
  nor_5  g05188(.A(new_n5564), .B(new_n5561), .Y(new_n5565));
  nor_5  g05189(.A(new_n5565), .B(new_n5560), .Y(new_n5566));
  nand_5 g05190(.A(new_n5566), .B(new_n5557), .Y(new_n5567));
  nand_5 g05191(.A(new_n5567), .B(new_n5556), .Y(new_n5568));
  nor_5  g05192(.A(new_n5495), .B(new_n5449), .Y(new_n5569));
  nand_5 g05193(.A(new_n5501), .B(new_n5496), .Y(new_n5570));
  not_8  g05194(.A(new_n5570), .Y(new_n5571));
  or_6   g05195(.A(new_n5571), .B(new_n5569), .Y(new_n5572));
  not_8  g05196(.A(new_n5484), .Y(new_n5573));
  nor_5  g05197(.A(new_n5494), .B(new_n5573), .Y(new_n5574));
  not_8  g05198(.A(new_n5480), .Y(new_n5575));
  nand_5 g05199(.A(new_n5575), .B(new_n5473), .Y(new_n5576));
  not_8  g05200(.A(new_n5481), .Y(new_n5577));
  nand_5 g05201(.A(new_n5577), .B(new_n5472), .Y(new_n5578));
  nand_5 g05202(.A(new_n5578), .B(new_n5576), .Y(new_n5579));
  nand_5 g05203(.A(pi087), .B(pi038), .Y(new_n5580));
  nand_5 g05204(.A(pi219), .B(pi113), .Y(new_n5581));
  xor_4  g05205(.A(new_n5581), .B(new_n5580), .Y(new_n5582));
  xor_4  g05206(.A(new_n5582), .B(new_n5463), .Y(new_n5583));
  xor_4  g05207(.A(new_n5583), .B(new_n5579), .Y(new_n5584));
  nand_5 g05208(.A(pi059), .B(pi051), .Y(new_n5585));
  nand_5 g05209(.A(pi122), .B(pi108), .Y(new_n5586));
  xor_4  g05210(.A(new_n5586), .B(new_n5585), .Y(new_n5587));
  xor_4  g05211(.A(new_n5587), .B(new_n5477), .Y(new_n5588));
  nand_5 g05212(.A(pi007), .B(pi001), .Y(new_n5589));
  xor_4  g05213(.A(new_n5589), .B(new_n5478), .Y(new_n5590));
  xor_4  g05214(.A(new_n5590), .B(new_n5588), .Y(new_n5591));
  xor_4  g05215(.A(new_n5591), .B(new_n5584), .Y(new_n5592));
  not_8  g05216(.A(new_n5482), .Y(new_n5593));
  nor_5  g05217(.A(new_n5593), .B(new_n5469), .Y(new_n5594));
  nor_5  g05218(.A(new_n5483), .B(new_n5462), .Y(new_n5595));
  xor_4  g05219(.A(new_n5595), .B(new_n5465), .Y(new_n5596));
  not_8  g05220(.A(new_n5596), .Y(new_n5597));
  nor_5  g05221(.A(new_n5597), .B(new_n5594), .Y(new_n5598));
  xor_4  g05222(.A(new_n5598), .B(new_n5592), .Y(new_n5599));
  xor_4  g05223(.A(new_n5599), .B(new_n5574), .Y(new_n5600));
  xor_4  g05224(.A(new_n5600), .B(new_n5572), .Y(new_n5601));
  nand_5 g05225(.A(new_n5525), .B(new_n5503), .Y(new_n5602));
  not_8  g05226(.A(new_n5554), .Y(new_n5603));
  nand_5 g05227(.A(new_n5603), .B(new_n5526), .Y(new_n5604));
  nand_5 g05228(.A(new_n5604), .B(new_n5602), .Y(new_n5605));
  nor_5  g05229(.A(new_n5553), .B(new_n5550), .Y(new_n5606));
  nand_5 g05230(.A(pi099), .B(pi061), .Y(new_n5607));
  nand_5 g05231(.A(pi188), .B(pi155), .Y(new_n5608));
  xor_4  g05232(.A(new_n5608), .B(new_n5607), .Y(new_n5609));
  xor_4  g05233(.A(new_n5609), .B(new_n5543), .Y(new_n5610));
  nand_5 g05234(.A(pi123), .B(pi012), .Y(new_n5611));
  xor_4  g05235(.A(new_n5611), .B(new_n5544), .Y(new_n5612));
  xor_4  g05236(.A(new_n5612), .B(new_n5610), .Y(new_n5613));
  nand_5 g05237(.A(new_n5546), .B(new_n5539), .Y(new_n5614));
  nand_5 g05238(.A(new_n5547), .B(new_n5538), .Y(new_n5615));
  nand_5 g05239(.A(new_n5615), .B(new_n5614), .Y(new_n5616));
  nand_5 g05240(.A(pi098), .B(pi071), .Y(new_n5617));
  nand_5 g05241(.A(pi142), .B(pi043), .Y(new_n5618));
  xor_4  g05242(.A(new_n5618), .B(new_n5617), .Y(new_n5619));
  xor_4  g05243(.A(new_n5619), .B(new_n5533), .Y(new_n5620));
  xor_4  g05244(.A(new_n5620), .B(new_n5616), .Y(new_n5621));
  not_8  g05245(.A(new_n5621), .Y(new_n5622));
  xor_4  g05246(.A(new_n5622), .B(new_n5613), .Y(new_n5623));
  nor_5  g05247(.A(new_n5548), .B(new_n5535), .Y(new_n5624));
  not_8  g05248(.A(new_n5549), .Y(new_n5625));
  nor_5  g05249(.A(new_n5625), .B(new_n5529), .Y(new_n5626));
  xor_4  g05250(.A(new_n5626), .B(new_n5534), .Y(new_n5627));
  nor_5  g05251(.A(new_n5627), .B(new_n5624), .Y(new_n5628));
  xor_4  g05252(.A(new_n5628), .B(new_n5623), .Y(new_n5629));
  xnor_4 g05253(.A(new_n5629), .B(new_n5606), .Y(new_n5630));
  xor_4  g05254(.A(new_n5630), .B(new_n5605), .Y(new_n5631));
  xor_4  g05255(.A(new_n5631), .B(new_n5601), .Y(new_n5632));
  xnor_4 g05256(.A(new_n5632), .B(new_n5568), .Y(new_n5633));
  nand_5 g05257(.A(pi238), .B(pi138), .Y(new_n5634));
  nand_5 g05258(.A(new_n4906), .B(new_n4895), .Y(new_n5635));
  not_8  g05259(.A(new_n5635), .Y(new_n5636));
  nand_5 g05260(.A(new_n4904), .B(new_n4901), .Y(new_n5637));
  nand_5 g05261(.A(new_n4905), .B(new_n4900), .Y(new_n5638));
  nand_5 g05262(.A(new_n5638), .B(new_n5637), .Y(new_n5639));
  nand_5 g05263(.A(pi237), .B(pi138), .Y(new_n5640));
  nand_5 g05264(.A(pi162), .B(pi076), .Y(new_n5641));
  nand_5 g05265(.A(pi216), .B(pi033), .Y(new_n5642));
  nand_5 g05266(.A(pi179), .B(pi041), .Y(new_n5643));
  xor_4  g05267(.A(new_n5643), .B(new_n5642), .Y(new_n5644));
  xor_4  g05268(.A(new_n5644), .B(new_n5641), .Y(new_n5645));
  nand_5 g05269(.A(pi182), .B(pi048), .Y(new_n5646));
  nand_5 g05270(.A(new_n4898), .B(new_n4897), .Y(new_n5647));
  nand_5 g05271(.A(new_n4899), .B(new_n4896), .Y(new_n5648));
  nand_5 g05272(.A(new_n5648), .B(new_n5647), .Y(new_n5649));
  xor_4  g05273(.A(new_n5649), .B(new_n5646), .Y(new_n5650));
  xor_4  g05274(.A(new_n5650), .B(new_n5645), .Y(new_n5651));
  xnor_4 g05275(.A(new_n5651), .B(new_n5640), .Y(new_n5652));
  xor_4  g05276(.A(new_n5652), .B(new_n5639), .Y(new_n5653));
  nand_5 g05277(.A(new_n5653), .B(new_n5636), .Y(new_n5654));
  nand_5 g05278(.A(new_n5654), .B(new_n5634), .Y(new_n5655));
  xor_4  g05279(.A(new_n5654), .B(new_n5634), .Y(new_n5656));
  nor_5  g05280(.A(new_n5651), .B(new_n5640), .Y(new_n5657));
  nor_5  g05281(.A(new_n5652), .B(new_n5639), .Y(new_n5658));
  nor_5  g05282(.A(new_n5658), .B(new_n5657), .Y(new_n5659));
  nand_5 g05283(.A(new_n5649), .B(new_n5646), .Y(new_n5660));
  nand_5 g05284(.A(new_n5650), .B(new_n5645), .Y(new_n5661));
  nand_5 g05285(.A(new_n5661), .B(new_n5660), .Y(new_n5662));
  nand_5 g05286(.A(pi237), .B(pi041), .Y(new_n5663));
  nor_5  g05287(.A(new_n5646), .B(new_n5663), .Y(new_n5664));
  not_8  g05288(.A(new_n5664), .Y(new_n5665));
  nand_5 g05289(.A(pi048), .B(pi041), .Y(new_n5666));
  nand_5 g05290(.A(pi237), .B(pi182), .Y(new_n5667));
  nand_5 g05291(.A(new_n5667), .B(new_n5666), .Y(new_n5668));
  nand_5 g05292(.A(new_n5668), .B(new_n5665), .Y(new_n5669));
  nand_5 g05293(.A(new_n5643), .B(new_n5642), .Y(new_n5670));
  nand_5 g05294(.A(new_n5644), .B(new_n5641), .Y(new_n5671));
  nand_5 g05295(.A(new_n5671), .B(new_n5670), .Y(new_n5672));
  nand_5 g05296(.A(pi216), .B(pi179), .Y(new_n5673));
  nand_5 g05297(.A(pi076), .B(pi033), .Y(new_n5674));
  nand_5 g05298(.A(pi162), .B(pi079), .Y(new_n5675));
  nand_5 g05299(.A(new_n5675), .B(new_n5674), .Y(new_n5676));
  nand_5 g05300(.A(pi079), .B(pi033), .Y(new_n5677));
  nor_5  g05301(.A(new_n5677), .B(new_n5641), .Y(new_n5678));
  not_8  g05302(.A(new_n5678), .Y(new_n5679));
  nand_5 g05303(.A(new_n5679), .B(new_n5676), .Y(new_n5680));
  xor_4  g05304(.A(new_n5680), .B(new_n5673), .Y(new_n5681));
  xor_4  g05305(.A(new_n5681), .B(new_n5672), .Y(new_n5682));
  xor_4  g05306(.A(new_n5682), .B(new_n5669), .Y(new_n5683));
  xor_4  g05307(.A(new_n5683), .B(new_n5662), .Y(new_n5684));
  xor_4  g05308(.A(new_n5684), .B(new_n5659), .Y(new_n5685));
  not_8  g05309(.A(new_n5685), .Y(new_n5686));
  nand_5 g05310(.A(new_n5686), .B(new_n5656), .Y(new_n5687));
  nand_5 g05311(.A(new_n5687), .B(new_n5655), .Y(new_n5688));
  nor_5  g05312(.A(new_n5684), .B(new_n5659), .Y(new_n5689));
  nand_5 g05313(.A(pi216), .B(pi048), .Y(new_n5690));
  xor_4  g05314(.A(new_n5690), .B(new_n5679), .Y(new_n5691));
  nand_5 g05315(.A(pi251), .B(pi162), .Y(new_n5692));
  nand_5 g05316(.A(pi179), .B(pi076), .Y(new_n5693));
  xor_4  g05317(.A(new_n5693), .B(new_n5692), .Y(new_n5694));
  xor_4  g05318(.A(new_n5694), .B(new_n5677), .Y(new_n5695));
  xor_4  g05319(.A(new_n5695), .B(new_n5691), .Y(new_n5696));
  nand_5 g05320(.A(new_n5680), .B(new_n5673), .Y(new_n5697));
  nand_5 g05321(.A(new_n5681), .B(new_n5672), .Y(new_n5698));
  nand_5 g05322(.A(new_n5698), .B(new_n5697), .Y(new_n5699));
  nand_5 g05323(.A(pi238), .B(pi182), .Y(new_n5700));
  nand_5 g05324(.A(pi193), .B(pi138), .Y(new_n5701));
  xor_4  g05325(.A(new_n5701), .B(new_n5700), .Y(new_n5702));
  xor_4  g05326(.A(new_n5702), .B(new_n5663), .Y(new_n5703));
  xor_4  g05327(.A(new_n5703), .B(new_n5699), .Y(new_n5704));
  xor_4  g05328(.A(new_n5704), .B(new_n5696), .Y(new_n5705));
  nand_5 g05329(.A(new_n5682), .B(new_n5669), .Y(new_n5706));
  nand_5 g05330(.A(new_n5683), .B(new_n5662), .Y(new_n5707));
  nand_5 g05331(.A(new_n5707), .B(new_n5706), .Y(new_n5708));
  xor_4  g05332(.A(new_n5708), .B(new_n5664), .Y(new_n5709));
  xor_4  g05333(.A(new_n5709), .B(new_n5705), .Y(new_n5710));
  xnor_4 g05334(.A(new_n5710), .B(new_n5689), .Y(new_n5711));
  xor_4  g05335(.A(new_n5711), .B(new_n5688), .Y(new_n5712));
  and_6  g05336(.A(new_n5712), .B(new_n5633), .Y(new_n5713));
  or_6   g05337(.A(new_n4958), .B(new_n4907), .Y(new_n5714));
  nand_5 g05338(.A(new_n4988), .B(new_n4959), .Y(new_n5715));
  nand_5 g05339(.A(new_n5715), .B(new_n5714), .Y(new_n5716));
  xor_4  g05340(.A(new_n5653), .B(new_n5635), .Y(new_n5717));
  or_6   g05341(.A(new_n5717), .B(new_n5716), .Y(new_n5718));
  xor_4  g05342(.A(new_n5564), .B(new_n5561), .Y(new_n5719));
  xnor_4 g05343(.A(new_n5717), .B(new_n5716), .Y(new_n5720));
  or_6   g05344(.A(new_n5720), .B(new_n5719), .Y(new_n5721));
  nand_5 g05345(.A(new_n5721), .B(new_n5718), .Y(new_n5722));
  xor_4  g05346(.A(new_n5566), .B(new_n5557), .Y(new_n5723));
  or_6   g05347(.A(new_n5723), .B(new_n5722), .Y(new_n5724));
  xor_4  g05348(.A(new_n5686), .B(new_n5656), .Y(new_n5725));
  xor_4  g05349(.A(new_n5723), .B(new_n5722), .Y(new_n5726));
  nand_5 g05350(.A(new_n5726), .B(new_n5725), .Y(new_n5727));
  nand_5 g05351(.A(new_n5727), .B(new_n5724), .Y(new_n5728));
  xnor_4 g05352(.A(new_n5712), .B(new_n5633), .Y(new_n5729));
  nor_5  g05353(.A(new_n5729), .B(new_n5728), .Y(new_n5730));
  nor_5  g05354(.A(new_n5730), .B(new_n5713), .Y(new_n5731));
  nand_5 g05355(.A(pi188), .B(pi086), .Y(new_n5732));
  xor_4  g05356(.A(new_n5732), .B(new_n5731), .Y(new_n5733));
  nand_5 g05357(.A(pi238), .B(pi041), .Y(new_n5734));
  nand_5 g05358(.A(pi143), .B(pi137), .Y(new_n5735));
  xor_4  g05359(.A(new_n5735), .B(new_n5734), .Y(new_n5736));
  nor_5  g05360(.A(new_n5611), .B(new_n5545), .Y(new_n5737));
  nor_5  g05361(.A(new_n5612), .B(new_n5610), .Y(new_n5738));
  or_6   g05362(.A(new_n5738), .B(new_n5737), .Y(new_n5739));
  nand_5 g05363(.A(pi118), .B(pi001), .Y(new_n5740));
  xor_4  g05364(.A(new_n5740), .B(new_n5739), .Y(new_n5741));
  nand_5 g05365(.A(pi099), .B(pi012), .Y(new_n5742));
  nand_5 g05366(.A(new_n5620), .B(new_n5616), .Y(new_n5743));
  or_6   g05367(.A(new_n5622), .B(new_n5613), .Y(new_n5744));
  nand_5 g05368(.A(new_n5744), .B(new_n5743), .Y(new_n5745));
  xor_4  g05369(.A(new_n5745), .B(new_n5742), .Y(new_n5746));
  nand_5 g05370(.A(pi169), .B(pi098), .Y(new_n5747));
  nand_5 g05371(.A(pi059), .B(pi042), .Y(new_n5748));
  xor_4  g05372(.A(new_n5748), .B(new_n5747), .Y(new_n5749));
  nand_5 g05373(.A(pi122), .B(pi007), .Y(new_n5750));
  nand_5 g05374(.A(new_n5618), .B(new_n5617), .Y(new_n5751));
  nand_5 g05375(.A(new_n5619), .B(new_n5533), .Y(new_n5752));
  nand_5 g05376(.A(new_n5752), .B(new_n5751), .Y(new_n5753));
  xnor_4 g05377(.A(new_n5753), .B(new_n5750), .Y(new_n5754));
  xor_4  g05378(.A(new_n5754), .B(new_n5749), .Y(new_n5755));
  xor_4  g05379(.A(new_n5755), .B(new_n5746), .Y(new_n5756));
  xor_4  g05380(.A(new_n5756), .B(new_n5741), .Y(new_n5757));
  xor_4  g05381(.A(new_n5757), .B(new_n5736), .Y(new_n5758));
  xor_4  g05382(.A(new_n5758), .B(new_n5733), .Y(new_n5759));
  nand_5 g05383(.A(new_n5710), .B(new_n5689), .Y(new_n5760));
  or_6   g05384(.A(new_n5711), .B(new_n5688), .Y(new_n5761));
  nand_5 g05385(.A(new_n5761), .B(new_n5760), .Y(new_n5762));
  nand_5 g05386(.A(pi193), .B(pi182), .Y(new_n5763));
  nand_5 g05387(.A(pi076), .B(pi048), .Y(new_n5764));
  xor_4  g05388(.A(new_n5764), .B(new_n5763), .Y(new_n5765));
  xor_4  g05389(.A(new_n5765), .B(new_n5762), .Y(new_n5766));
  nor_5  g05390(.A(new_n5708), .B(new_n5665), .Y(new_n5767));
  nor_5  g05391(.A(new_n5709), .B(new_n5705), .Y(new_n5768));
  nor_5  g05392(.A(new_n5768), .B(new_n5767), .Y(new_n5769));
  nand_5 g05393(.A(pi142), .B(pi126), .Y(new_n5770));
  xor_4  g05394(.A(new_n5770), .B(new_n5769), .Y(new_n5771));
  xor_4  g05395(.A(new_n5771), .B(new_n5766), .Y(new_n5772));
  not_8  g05396(.A(new_n5574), .Y(new_n5773));
  nor_5  g05397(.A(new_n5599), .B(new_n5773), .Y(new_n5774));
  not_8  g05398(.A(new_n5572), .Y(new_n5775));
  nor_5  g05399(.A(new_n5600), .B(new_n5775), .Y(new_n5776));
  or_6   g05400(.A(new_n5776), .B(new_n5774), .Y(new_n5777));
  not_8  g05401(.A(new_n5029), .Y(new_n5778));
  nand_5 g05402(.A(new_n5778), .B(new_n5018), .Y(new_n5779));
  not_8  g05403(.A(new_n5779), .Y(new_n5780));
  nand_5 g05404(.A(pi180), .B(pi160), .Y(new_n5781));
  nand_5 g05405(.A(pi194), .B(pi060), .Y(new_n5782));
  nand_5 g05406(.A(pi223), .B(pi057), .Y(new_n5783));
  nand_5 g05407(.A(pi143), .B(pi101), .Y(new_n5784));
  xor_4  g05408(.A(new_n5784), .B(new_n5783), .Y(new_n5785));
  xor_4  g05409(.A(new_n5785), .B(new_n5782), .Y(new_n5786));
  nand_5 g05410(.A(new_n5021), .B(new_n5020), .Y(new_n5787));
  nand_5 g05411(.A(new_n5022), .B(new_n5019), .Y(new_n5788));
  nand_5 g05412(.A(new_n5788), .B(new_n5787), .Y(new_n5789));
  nand_5 g05413(.A(pi085), .B(pi020), .Y(new_n5790));
  xor_4  g05414(.A(new_n5790), .B(new_n5789), .Y(new_n5791));
  xor_4  g05415(.A(new_n5791), .B(new_n5786), .Y(new_n5792));
  nand_5 g05416(.A(new_n5792), .B(new_n5781), .Y(new_n5793));
  or_6   g05417(.A(new_n5792), .B(new_n5781), .Y(new_n5794));
  nand_5 g05418(.A(new_n5794), .B(new_n5793), .Y(new_n5795));
  nand_5 g05419(.A(new_n5027), .B(new_n5024), .Y(new_n5796));
  nand_5 g05420(.A(new_n5028), .B(new_n5023), .Y(new_n5797));
  nand_5 g05421(.A(new_n5797), .B(new_n5796), .Y(new_n5798));
  xor_4  g05422(.A(new_n5798), .B(new_n5795), .Y(new_n5799));
  nand_5 g05423(.A(new_n5799), .B(new_n5780), .Y(new_n5800));
  nand_5 g05424(.A(pi160), .B(pi036), .Y(new_n5801));
  nand_5 g05425(.A(new_n5801), .B(new_n5800), .Y(new_n5802));
  not_8  g05426(.A(new_n5802), .Y(new_n5803));
  xor_4  g05427(.A(new_n5801), .B(new_n5800), .Y(new_n5804));
  not_8  g05428(.A(new_n5804), .Y(new_n5805));
  nand_5 g05429(.A(new_n5790), .B(new_n5789), .Y(new_n5806));
  nand_5 g05430(.A(new_n5791), .B(new_n5786), .Y(new_n5807));
  nand_5 g05431(.A(new_n5807), .B(new_n5806), .Y(new_n5808));
  nand_5 g05432(.A(pi180), .B(pi020), .Y(new_n5809));
  nand_5 g05433(.A(pi085), .B(pi060), .Y(new_n5810));
  nand_5 g05434(.A(new_n5810), .B(new_n5809), .Y(new_n5811));
  nand_5 g05435(.A(pi180), .B(pi060), .Y(new_n5812));
  nor_5  g05436(.A(new_n5812), .B(new_n5790), .Y(new_n5813));
  not_8  g05437(.A(new_n5813), .Y(new_n5814));
  nand_5 g05438(.A(new_n5814), .B(new_n5811), .Y(new_n5815));
  nand_5 g05439(.A(new_n5784), .B(new_n5783), .Y(new_n5816));
  nand_5 g05440(.A(new_n5785), .B(new_n5782), .Y(new_n5817));
  nand_5 g05441(.A(new_n5817), .B(new_n5816), .Y(new_n5818));
  nand_5 g05442(.A(pi223), .B(pi194), .Y(new_n5819));
  nand_5 g05443(.A(pi101), .B(pi057), .Y(new_n5820));
  nand_5 g05444(.A(pi225), .B(pi143), .Y(new_n5821));
  nand_5 g05445(.A(new_n5821), .B(new_n5820), .Y(new_n5822));
  nand_5 g05446(.A(pi225), .B(pi057), .Y(new_n5823));
  nor_5  g05447(.A(new_n5823), .B(new_n5784), .Y(new_n5824));
  not_8  g05448(.A(new_n5824), .Y(new_n5825));
  nand_5 g05449(.A(new_n5825), .B(new_n5822), .Y(new_n5826));
  xor_4  g05450(.A(new_n5826), .B(new_n5819), .Y(new_n5827));
  xor_4  g05451(.A(new_n5827), .B(new_n5818), .Y(new_n5828));
  xnor_4 g05452(.A(new_n5828), .B(new_n5815), .Y(new_n5829));
  xnor_4 g05453(.A(new_n5829), .B(new_n5808), .Y(new_n5830));
  nand_5 g05454(.A(new_n5798), .B(new_n5794), .Y(new_n5831));
  nand_5 g05455(.A(new_n5831), .B(new_n5793), .Y(new_n5832));
  xor_4  g05456(.A(new_n5832), .B(new_n5830), .Y(new_n5833));
  nor_5  g05457(.A(new_n5833), .B(new_n5805), .Y(new_n5834));
  nor_5  g05458(.A(new_n5834), .B(new_n5803), .Y(new_n5835));
  nand_5 g05459(.A(pi177), .B(pi143), .Y(new_n5836));
  nand_5 g05460(.A(pi194), .B(pi101), .Y(new_n5837));
  xor_4  g05461(.A(new_n5837), .B(new_n5836), .Y(new_n5838));
  xor_4  g05462(.A(new_n5838), .B(new_n5823), .Y(new_n5839));
  nand_5 g05463(.A(pi223), .B(pi085), .Y(new_n5840));
  xor_4  g05464(.A(new_n5840), .B(new_n5824), .Y(new_n5841));
  xor_4  g05465(.A(new_n5841), .B(new_n5839), .Y(new_n5842));
  nand_5 g05466(.A(new_n5826), .B(new_n5819), .Y(new_n5843));
  nand_5 g05467(.A(new_n5827), .B(new_n5818), .Y(new_n5844));
  nand_5 g05468(.A(new_n5844), .B(new_n5843), .Y(new_n5845));
  nand_5 g05469(.A(pi160), .B(pi068), .Y(new_n5846));
  nand_5 g05470(.A(pi036), .B(pi020), .Y(new_n5847));
  xor_4  g05471(.A(new_n5847), .B(new_n5846), .Y(new_n5848));
  xor_4  g05472(.A(new_n5848), .B(new_n5812), .Y(new_n5849));
  xor_4  g05473(.A(new_n5849), .B(new_n5845), .Y(new_n5850));
  xor_4  g05474(.A(new_n5850), .B(new_n5842), .Y(new_n5851));
  nor_5  g05475(.A(new_n5828), .B(new_n5815), .Y(new_n5852));
  nor_5  g05476(.A(new_n5829), .B(new_n5808), .Y(new_n5853));
  xor_4  g05477(.A(new_n5853), .B(new_n5814), .Y(new_n5854));
  not_8  g05478(.A(new_n5854), .Y(new_n5855));
  nor_5  g05479(.A(new_n5855), .B(new_n5852), .Y(new_n5856));
  xor_4  g05480(.A(new_n5856), .B(new_n5851), .Y(new_n5857));
  not_8  g05481(.A(new_n5857), .Y(new_n5858));
  nor_5  g05482(.A(new_n5858), .B(new_n5835), .Y(new_n5859));
  nor_5  g05483(.A(new_n5832), .B(new_n5830), .Y(new_n5860));
  xor_4  g05484(.A(new_n5858), .B(new_n5835), .Y(new_n5861));
  not_8  g05485(.A(new_n5861), .Y(new_n5862));
  nor_5  g05486(.A(new_n5862), .B(new_n5860), .Y(new_n5863));
  nor_5  g05487(.A(new_n5863), .B(new_n5859), .Y(new_n5864));
  xor_4  g05488(.A(new_n5864), .B(new_n5777), .Y(new_n5865));
  nand_5 g05489(.A(pi087), .B(pi028), .Y(new_n5866));
  xor_4  g05490(.A(new_n5866), .B(new_n5865), .Y(new_n5867));
  nand_5 g05491(.A(pi071), .B(pi043), .Y(new_n5868));
  nand_5 g05492(.A(pi144), .B(pi123), .Y(new_n5869));
  nand_5 g05493(.A(new_n5595), .B(new_n5464), .Y(new_n5870));
  not_8  g05494(.A(new_n5598), .Y(new_n5871));
  nand_5 g05495(.A(new_n5871), .B(new_n5592), .Y(new_n5872));
  nand_5 g05496(.A(new_n5872), .B(new_n5870), .Y(new_n5873));
  nand_5 g05497(.A(pi135), .B(pi108), .Y(new_n5874));
  xor_4  g05498(.A(new_n5874), .B(new_n5873), .Y(new_n5875));
  xor_4  g05499(.A(new_n5875), .B(new_n5869), .Y(new_n5876));
  xor_4  g05500(.A(new_n5876), .B(new_n5868), .Y(new_n5877));
  xor_4  g05501(.A(new_n5877), .B(new_n5867), .Y(new_n5878));
  xor_4  g05502(.A(new_n5878), .B(new_n5772), .Y(new_n5879));
  xor_4  g05503(.A(new_n5879), .B(new_n5759), .Y(new_n5880));
  nand_5 g05504(.A(pi159), .B(pi138), .Y(new_n5881));
  nand_5 g05505(.A(new_n5703), .B(new_n5699), .Y(new_n5882));
  nand_5 g05506(.A(new_n5704), .B(new_n5696), .Y(new_n5883));
  nand_5 g05507(.A(new_n5883), .B(new_n5882), .Y(new_n5884));
  nor_5  g05508(.A(new_n5629), .B(new_n5606), .Y(new_n5885));
  not_8  g05509(.A(new_n5605), .Y(new_n5886));
  nor_5  g05510(.A(new_n5630), .B(new_n5886), .Y(new_n5887));
  nor_5  g05511(.A(new_n5887), .B(new_n5885), .Y(new_n5888));
  xor_4  g05512(.A(new_n5888), .B(new_n5884), .Y(new_n5889));
  nand_5 g05513(.A(pi192), .B(pi162), .Y(new_n5890));
  or_6   g05514(.A(new_n5690), .B(new_n5679), .Y(new_n5891));
  not_8  g05515(.A(new_n5695), .Y(new_n5892));
  nand_5 g05516(.A(new_n5892), .B(new_n5691), .Y(new_n5893));
  nand_5 g05517(.A(new_n5893), .B(new_n5891), .Y(new_n5894));
  and_6  g05518(.A(new_n5626), .B(new_n5534), .Y(new_n5895));
  nor_5  g05519(.A(new_n5628), .B(new_n5623), .Y(new_n5896));
  nor_5  g05520(.A(new_n5896), .B(new_n5895), .Y(new_n5897));
  xor_4  g05521(.A(new_n5897), .B(new_n5894), .Y(new_n5898));
  xor_4  g05522(.A(new_n5898), .B(new_n5890), .Y(new_n5899));
  xor_4  g05523(.A(new_n5899), .B(new_n5889), .Y(new_n5900));
  xor_4  g05524(.A(new_n5900), .B(new_n5881), .Y(new_n5901));
  xor_4  g05525(.A(new_n5901), .B(new_n5880), .Y(new_n5902));
  nand_5 g05526(.A(pi179), .B(pi079), .Y(new_n5903));
  nand_5 g05527(.A(new_n5693), .B(new_n5692), .Y(new_n5904));
  nand_5 g05528(.A(new_n5694), .B(new_n5677), .Y(new_n5905));
  nand_5 g05529(.A(new_n5905), .B(new_n5904), .Y(new_n5906));
  nand_5 g05530(.A(pi251), .B(pi033), .Y(new_n5907));
  xor_4  g05531(.A(new_n5907), .B(new_n5906), .Y(new_n5908));
  xor_4  g05532(.A(new_n5908), .B(new_n5903), .Y(new_n5909));
  nand_5 g05533(.A(pi061), .B(pi023), .Y(new_n5910));
  nand_5 g05534(.A(pi178), .B(pi155), .Y(new_n5911));
  xor_4  g05535(.A(new_n5911), .B(new_n5910), .Y(new_n5912));
  not_8  g05536(.A(new_n5601), .Y(new_n5913));
  nor_5  g05537(.A(new_n5631), .B(new_n5913), .Y(new_n5914));
  nor_5  g05538(.A(new_n5632), .B(new_n5568), .Y(new_n5915));
  nor_5  g05539(.A(new_n5915), .B(new_n5914), .Y(new_n5916));
  xor_4  g05540(.A(new_n5916), .B(new_n5912), .Y(new_n5917));
  or_6   g05541(.A(new_n5849), .B(new_n5845), .Y(new_n5918));
  nand_5 g05542(.A(new_n5850), .B(new_n5842), .Y(new_n5919));
  nand_5 g05543(.A(new_n5919), .B(new_n5918), .Y(new_n5920));
  nor_5  g05544(.A(new_n5840), .B(new_n5825), .Y(new_n5921));
  nor_5  g05545(.A(new_n5841), .B(new_n5839), .Y(new_n5922));
  nor_5  g05546(.A(new_n5922), .B(new_n5921), .Y(new_n5923));
  nand_5 g05547(.A(pi060), .B(pi036), .Y(new_n5924));
  xor_4  g05548(.A(new_n5924), .B(new_n5923), .Y(new_n5925));
  xor_4  g05549(.A(new_n5925), .B(new_n5920), .Y(new_n5926));
  nand_5 g05550(.A(pi068), .B(pi020), .Y(new_n5927));
  nand_5 g05551(.A(pi101), .B(pi085), .Y(new_n5928));
  xor_4  g05552(.A(new_n5928), .B(new_n5927), .Y(new_n5929));
  nand_5 g05553(.A(pi223), .B(pi180), .Y(new_n5930));
  nand_5 g05554(.A(new_n5837), .B(new_n5836), .Y(new_n5931));
  nand_5 g05555(.A(new_n5838), .B(new_n5823), .Y(new_n5932));
  nand_5 g05556(.A(new_n5932), .B(new_n5931), .Y(new_n5933));
  nand_5 g05557(.A(new_n5847), .B(new_n5846), .Y(new_n5934));
  nand_5 g05558(.A(new_n5848), .B(new_n5812), .Y(new_n5935));
  nand_5 g05559(.A(new_n5935), .B(new_n5934), .Y(new_n5936));
  xor_4  g05560(.A(new_n5936), .B(new_n5933), .Y(new_n5937));
  xor_4  g05561(.A(new_n5937), .B(new_n5930), .Y(new_n5938));
  xor_4  g05562(.A(new_n5938), .B(new_n5929), .Y(new_n5939));
  xor_4  g05563(.A(new_n5939), .B(new_n5926), .Y(new_n5940));
  xor_4  g05564(.A(new_n5940), .B(new_n5917), .Y(new_n5941));
  xor_4  g05565(.A(new_n5941), .B(new_n5909), .Y(new_n5942));
  xor_4  g05566(.A(new_n5833), .B(new_n5805), .Y(new_n5943));
  xor_4  g05567(.A(new_n5726), .B(new_n5725), .Y(new_n5944));
  and_6  g05568(.A(new_n5944), .B(new_n5943), .Y(new_n5945));
  or_6   g05569(.A(new_n5030), .B(new_n5016), .Y(new_n5946));
  nand_5 g05570(.A(new_n5031), .B(new_n4989), .Y(new_n5947));
  nand_5 g05571(.A(new_n5947), .B(new_n5946), .Y(new_n5948));
  xor_4  g05572(.A(new_n5799), .B(new_n5779), .Y(new_n5949));
  not_8  g05573(.A(new_n5949), .Y(new_n5950));
  nor_5  g05574(.A(new_n5950), .B(new_n5948), .Y(new_n5951));
  xor_4  g05575(.A(new_n5949), .B(new_n5948), .Y(new_n5952));
  xor_4  g05576(.A(new_n5720), .B(new_n5719), .Y(new_n5953));
  nor_5  g05577(.A(new_n5953), .B(new_n5952), .Y(new_n5954));
  nor_5  g05578(.A(new_n5954), .B(new_n5951), .Y(new_n5955));
  xnor_4 g05579(.A(new_n5944), .B(new_n5943), .Y(new_n5956));
  nor_5  g05580(.A(new_n5956), .B(new_n5955), .Y(new_n5957));
  nor_5  g05581(.A(new_n5957), .B(new_n5945), .Y(new_n5958));
  xor_4  g05582(.A(new_n5861), .B(new_n5860), .Y(new_n5959));
  or_6   g05583(.A(new_n5959), .B(new_n5958), .Y(new_n5960));
  xnor_4 g05584(.A(new_n5729), .B(new_n5728), .Y(new_n5961));
  xor_4  g05585(.A(new_n5959), .B(new_n5958), .Y(new_n5962));
  nand_5 g05586(.A(new_n5962), .B(new_n5961), .Y(new_n5963));
  nand_5 g05587(.A(new_n5963), .B(new_n5960), .Y(new_n5964));
  nand_5 g05588(.A(pi094), .B(pi051), .Y(new_n5965));
  nand_5 g05589(.A(pi237), .B(pi216), .Y(new_n5966));
  nand_5 g05590(.A(new_n5701), .B(new_n5700), .Y(new_n5967));
  nand_5 g05591(.A(new_n5702), .B(new_n5663), .Y(new_n5968));
  nand_5 g05592(.A(new_n5968), .B(new_n5967), .Y(new_n5969));
  xor_4  g05593(.A(new_n5969), .B(new_n5966), .Y(new_n5970));
  xor_4  g05594(.A(new_n5970), .B(new_n5965), .Y(new_n5971));
  xor_4  g05595(.A(new_n5971), .B(new_n5964), .Y(new_n5972));
  nand_5 g05596(.A(pi160), .B(pi046), .Y(new_n5973));
  nand_5 g05597(.A(new_n5586), .B(new_n5585), .Y(new_n5974));
  nand_5 g05598(.A(new_n5587), .B(new_n5477), .Y(new_n5975));
  nand_5 g05599(.A(new_n5975), .B(new_n5974), .Y(new_n5976));
  xor_4  g05600(.A(new_n5976), .B(new_n5973), .Y(new_n5977));
  or_6   g05601(.A(new_n5583), .B(new_n5579), .Y(new_n5978));
  nand_5 g05602(.A(new_n5591), .B(new_n5584), .Y(new_n5979));
  nand_5 g05603(.A(new_n5979), .B(new_n5978), .Y(new_n5980));
  nor_5  g05604(.A(new_n5589), .B(new_n5479), .Y(new_n5981));
  nor_5  g05605(.A(new_n5590), .B(new_n5588), .Y(new_n5982));
  nor_5  g05606(.A(new_n5982), .B(new_n5981), .Y(new_n5983));
  xor_4  g05607(.A(new_n5983), .B(new_n5980), .Y(new_n5984));
  xor_4  g05608(.A(new_n5984), .B(new_n5977), .Y(new_n5985));
  nand_5 g05609(.A(new_n5853), .B(new_n5813), .Y(new_n5986));
  not_8  g05610(.A(new_n5856), .Y(new_n5987));
  nand_5 g05611(.A(new_n5987), .B(new_n5851), .Y(new_n5988));
  nand_5 g05612(.A(new_n5988), .B(new_n5986), .Y(new_n5989));
  nand_5 g05613(.A(new_n5608), .B(new_n5607), .Y(new_n5990));
  nand_5 g05614(.A(new_n5609), .B(new_n5543), .Y(new_n5991));
  nand_5 g05615(.A(new_n5991), .B(new_n5990), .Y(new_n5992));
  nand_5 g05616(.A(new_n5581), .B(new_n5580), .Y(new_n5993));
  nand_5 g05617(.A(new_n5582), .B(new_n5463), .Y(new_n5994));
  nand_5 g05618(.A(new_n5994), .B(new_n5993), .Y(new_n5995));
  xnor_4 g05619(.A(new_n5995), .B(new_n5992), .Y(new_n5996));
  nand_5 g05620(.A(pi113), .B(pi102), .Y(new_n5997));
  nand_5 g05621(.A(pi219), .B(pi038), .Y(new_n5998));
  xor_4  g05622(.A(new_n5998), .B(new_n5997), .Y(new_n5999));
  xor_4  g05623(.A(new_n5999), .B(new_n5996), .Y(new_n6000));
  xor_4  g05624(.A(new_n6000), .B(new_n5989), .Y(new_n6001));
  xor_4  g05625(.A(new_n6001), .B(new_n5985), .Y(new_n6002));
  nand_5 g05626(.A(pi225), .B(pi194), .Y(new_n6003));
  nand_5 g05627(.A(pi177), .B(pi057), .Y(new_n6004));
  xor_4  g05628(.A(new_n6004), .B(new_n6003), .Y(new_n6005));
  xor_4  g05629(.A(new_n6005), .B(new_n6002), .Y(new_n6006));
  xor_4  g05630(.A(new_n6006), .B(new_n5972), .Y(new_n6007));
  xor_4  g05631(.A(new_n6007), .B(new_n5942), .Y(new_n6008));
  xor_4  g05632(.A(new_n6008), .B(new_n5902), .Y(po021));
  xor_4  g05633(.A(new_n4784), .B(new_n4783), .Y(po022));
  xor_4  g05634(.A(new_n2589), .B(new_n2549), .Y(po023));
  xnor_4 g05635(.A(new_n1359), .B(new_n1358), .Y(po024));
  xnor_4 g05636(.A(new_n4225), .B(new_n4224), .Y(po025));
  xor_4  g05637(.A(new_n5444), .B(new_n5442), .Y(po026));
  nand_5 g05638(.A(pi130), .B(pi104), .Y(new_n6015));
  nand_5 g05639(.A(pi212), .B(pi124), .Y(new_n6016));
  nand_5 g05640(.A(new_n6016), .B(new_n6015), .Y(new_n6017));
  nand_5 g05641(.A(pi215), .B(pi213), .Y(new_n6018));
  xor_4  g05642(.A(new_n6016), .B(new_n6015), .Y(new_n6019));
  nand_5 g05643(.A(new_n6019), .B(new_n6018), .Y(new_n6020));
  nand_5 g05644(.A(new_n6020), .B(new_n6017), .Y(new_n6021));
  nand_5 g05645(.A(pi208), .B(pi197), .Y(new_n6022));
  nand_5 g05646(.A(new_n3461), .B(new_n3444), .Y(new_n6023));
  not_8  g05647(.A(new_n6023), .Y(new_n6024));
  nor_5  g05648(.A(new_n3448), .B(new_n3445), .Y(new_n6025));
  and_6  g05649(.A(new_n3460), .B(new_n3449), .Y(new_n6026));
  nor_5  g05650(.A(new_n6026), .B(new_n6025), .Y(new_n6027));
  nand_5 g05651(.A(pi254), .B(pi047), .Y(new_n6028));
  nand_5 g05652(.A(pi158), .B(pi090), .Y(new_n6029));
  nand_5 g05653(.A(new_n6029), .B(new_n6028), .Y(new_n6030));
  nand_5 g05654(.A(pi158), .B(pi047), .Y(new_n6031));
  nor_5  g05655(.A(new_n6031), .B(new_n3451), .Y(new_n6032));
  not_8  g05656(.A(new_n6032), .Y(new_n6033));
  nand_5 g05657(.A(new_n6033), .B(new_n6030), .Y(new_n6034));
  nand_5 g05658(.A(pi141), .B(pi089), .Y(new_n6035));
  nand_5 g05659(.A(new_n3452), .B(new_n3451), .Y(new_n6036));
  nand_5 g05660(.A(new_n3453), .B(new_n3450), .Y(new_n6037));
  nand_5 g05661(.A(new_n6037), .B(new_n6036), .Y(new_n6038));
  xor_4  g05662(.A(new_n6038), .B(new_n6035), .Y(new_n6039));
  xor_4  g05663(.A(new_n6039), .B(new_n6034), .Y(new_n6040));
  and_6  g05664(.A(new_n3458), .B(new_n3455), .Y(new_n6041));
  and_6  g05665(.A(new_n3459), .B(new_n3454), .Y(new_n6042));
  nor_5  g05666(.A(new_n6042), .B(new_n6041), .Y(new_n6043));
  nand_5 g05667(.A(pi161), .B(pi154), .Y(new_n6044));
  nand_5 g05668(.A(pi241), .B(pi095), .Y(new_n6045));
  nand_5 g05669(.A(new_n6045), .B(new_n6044), .Y(new_n6046));
  nand_5 g05670(.A(pi161), .B(pi095), .Y(new_n6047));
  or_6   g05671(.A(new_n6047), .B(new_n3455), .Y(new_n6048));
  nand_5 g05672(.A(new_n6048), .B(new_n6046), .Y(new_n6049));
  xor_4  g05673(.A(new_n6049), .B(new_n6043), .Y(new_n6050));
  xor_4  g05674(.A(new_n6050), .B(new_n6040), .Y(new_n6051));
  xor_4  g05675(.A(new_n6051), .B(new_n6027), .Y(new_n6052));
  nand_5 g05676(.A(pi236), .B(pi006), .Y(new_n6053));
  xor_4  g05677(.A(new_n6053), .B(new_n6052), .Y(new_n6054));
  xor_4  g05678(.A(new_n6054), .B(new_n6024), .Y(new_n6055));
  and_6  g05679(.A(new_n3482), .B(new_n3465), .Y(new_n6056));
  nand_5 g05680(.A(pi213), .B(pi124), .Y(new_n6057));
  nand_5 g05681(.A(new_n3479), .B(new_n3478), .Y(new_n6058));
  nand_5 g05682(.A(new_n3480), .B(new_n3475), .Y(new_n6059));
  nand_5 g05683(.A(new_n6059), .B(new_n6058), .Y(new_n6060));
  nand_5 g05684(.A(pi212), .B(pi130), .Y(new_n6061));
  nand_5 g05685(.A(pi104), .B(pi003), .Y(new_n6062));
  and_6  g05686(.A(new_n6062), .B(new_n6061), .Y(new_n6063));
  nor_5  g05687(.A(new_n6015), .B(new_n3479), .Y(new_n6064));
  or_6   g05688(.A(new_n6064), .B(new_n6063), .Y(new_n6065));
  nand_5 g05689(.A(new_n3473), .B(new_n3472), .Y(new_n6066));
  nand_5 g05690(.A(new_n3474), .B(new_n3471), .Y(new_n6067));
  nand_5 g05691(.A(new_n6067), .B(new_n6066), .Y(new_n6068));
  nand_5 g05692(.A(pi073), .B(pi013), .Y(new_n6069));
  nand_5 g05693(.A(pi112), .B(pi004), .Y(new_n6070));
  nand_5 g05694(.A(pi170), .B(pi105), .Y(new_n6071));
  nand_5 g05695(.A(new_n6071), .B(new_n6070), .Y(new_n6072));
  nand_5 g05696(.A(pi105), .B(pi004), .Y(new_n6073));
  nor_5  g05697(.A(new_n6073), .B(new_n3473), .Y(new_n6074));
  not_8  g05698(.A(new_n6074), .Y(new_n6075));
  and_6  g05699(.A(new_n6075), .B(new_n6072), .Y(new_n6076));
  xor_4  g05700(.A(new_n6076), .B(new_n6069), .Y(new_n6077));
  xor_4  g05701(.A(new_n6077), .B(new_n6068), .Y(new_n6078));
  xor_4  g05702(.A(new_n6078), .B(new_n6065), .Y(new_n6079));
  xor_4  g05703(.A(new_n6079), .B(new_n6060), .Y(new_n6080));
  nand_5 g05704(.A(new_n3469), .B(new_n3466), .Y(new_n6081));
  nand_5 g05705(.A(new_n3481), .B(new_n3470), .Y(new_n6082));
  nand_5 g05706(.A(new_n6082), .B(new_n6081), .Y(new_n6083));
  xor_4  g05707(.A(new_n6083), .B(new_n6080), .Y(new_n6084));
  xor_4  g05708(.A(new_n6084), .B(new_n6057), .Y(new_n6085));
  xor_4  g05709(.A(new_n6085), .B(new_n6056), .Y(new_n6086));
  and_6  g05710(.A(new_n6086), .B(new_n6055), .Y(new_n6087));
  nand_5 g05711(.A(new_n3462), .B(new_n3443), .Y(new_n6088));
  nand_5 g05712(.A(new_n3483), .B(new_n3463), .Y(new_n6089));
  nand_5 g05713(.A(new_n6089), .B(new_n6088), .Y(new_n6090));
  xnor_4 g05714(.A(new_n6086), .B(new_n6055), .Y(new_n6091));
  nor_5  g05715(.A(new_n6091), .B(new_n6090), .Y(new_n6092));
  nor_5  g05716(.A(new_n6092), .B(new_n6087), .Y(new_n6093));
  not_8  g05717(.A(new_n6080), .Y(new_n6094));
  nor_5  g05718(.A(new_n6083), .B(new_n6094), .Y(new_n6095));
  nand_5 g05719(.A(pi183), .B(pi170), .Y(new_n6096));
  nand_5 g05720(.A(pi112), .B(pi073), .Y(new_n6097));
  xor_4  g05721(.A(new_n6097), .B(new_n6096), .Y(new_n6098));
  xor_4  g05722(.A(new_n6098), .B(new_n6073), .Y(new_n6099));
  nand_5 g05723(.A(pi013), .B(pi003), .Y(new_n6100));
  xor_4  g05724(.A(new_n6100), .B(new_n6074), .Y(new_n6101));
  xor_4  g05725(.A(new_n6101), .B(new_n6099), .Y(new_n6102));
  not_8  g05726(.A(new_n6102), .Y(new_n6103));
  not_8  g05727(.A(new_n6076), .Y(new_n6104));
  nand_5 g05728(.A(new_n6104), .B(new_n6069), .Y(new_n6105));
  not_8  g05729(.A(new_n6077), .Y(new_n6106));
  nand_5 g05730(.A(new_n6106), .B(new_n6068), .Y(new_n6107));
  nand_5 g05731(.A(new_n6107), .B(new_n6105), .Y(new_n6108));
  xor_4  g05732(.A(new_n6019), .B(new_n6018), .Y(new_n6109));
  xor_4  g05733(.A(new_n6109), .B(new_n6108), .Y(new_n6110));
  xor_4  g05734(.A(new_n6110), .B(new_n6103), .Y(new_n6111));
  nor_5  g05735(.A(new_n6079), .B(new_n6060), .Y(new_n6112));
  nand_5 g05736(.A(new_n6112), .B(new_n6064), .Y(new_n6113));
  not_8  g05737(.A(new_n6112), .Y(new_n6114));
  not_8  g05738(.A(new_n6078), .Y(new_n6115));
  nor_5  g05739(.A(new_n6115), .B(new_n6065), .Y(new_n6116));
  nor_5  g05740(.A(new_n6116), .B(new_n6064), .Y(new_n6117));
  nand_5 g05741(.A(new_n6117), .B(new_n6114), .Y(new_n6118));
  nand_5 g05742(.A(new_n6118), .B(new_n6113), .Y(new_n6119));
  xor_4  g05743(.A(new_n6119), .B(new_n6111), .Y(new_n6120));
  xor_4  g05744(.A(new_n6120), .B(new_n6095), .Y(new_n6121));
  nor_5  g05745(.A(new_n6084), .B(new_n6057), .Y(new_n6122));
  and_6  g05746(.A(new_n6085), .B(new_n6056), .Y(new_n6123));
  nor_5  g05747(.A(new_n6123), .B(new_n6122), .Y(new_n6124));
  xor_4  g05748(.A(new_n6124), .B(new_n6121), .Y(new_n6125));
  nor_5  g05749(.A(new_n6125), .B(new_n6093), .Y(new_n6126));
  xnor_4 g05750(.A(new_n6125), .B(new_n6093), .Y(new_n6127));
  not_8  g05751(.A(new_n6051), .Y(new_n6128));
  nor_5  g05752(.A(new_n6128), .B(new_n6027), .Y(new_n6129));
  not_8  g05753(.A(new_n6043), .Y(new_n6130));
  nand_5 g05754(.A(new_n6049), .B(new_n6130), .Y(new_n6131));
  not_8  g05755(.A(new_n6050), .Y(new_n6132));
  nand_5 g05756(.A(new_n6132), .B(new_n6040), .Y(new_n6133));
  nand_5 g05757(.A(new_n6133), .B(new_n6131), .Y(new_n6134));
  xor_4  g05758(.A(new_n6134), .B(new_n6048), .Y(new_n6135));
  nand_5 g05759(.A(pi090), .B(pi089), .Y(new_n6136));
  nand_5 g05760(.A(pi254), .B(pi018), .Y(new_n6137));
  xor_4  g05761(.A(new_n6137), .B(new_n6136), .Y(new_n6138));
  xor_4  g05762(.A(new_n6138), .B(new_n6031), .Y(new_n6139));
  nand_5 g05763(.A(pi154), .B(pi141), .Y(new_n6140));
  xor_4  g05764(.A(new_n6140), .B(new_n6032), .Y(new_n6141));
  xor_4  g05765(.A(new_n6141), .B(new_n6139), .Y(new_n6142));
  nand_5 g05766(.A(new_n6038), .B(new_n6035), .Y(new_n6143));
  nand_5 g05767(.A(new_n6039), .B(new_n6034), .Y(new_n6144));
  nand_5 g05768(.A(new_n6144), .B(new_n6143), .Y(new_n6145));
  nand_5 g05769(.A(pi241), .B(pi006), .Y(new_n6146));
  nand_5 g05770(.A(pi236), .B(pi209), .Y(new_n6147));
  xor_4  g05771(.A(new_n6147), .B(new_n6146), .Y(new_n6148));
  xnor_4 g05772(.A(new_n6148), .B(new_n6047), .Y(new_n6149));
  xor_4  g05773(.A(new_n6149), .B(new_n6145), .Y(new_n6150));
  xor_4  g05774(.A(new_n6150), .B(new_n6142), .Y(new_n6151));
  not_8  g05775(.A(new_n6151), .Y(new_n6152));
  xor_4  g05776(.A(new_n6152), .B(new_n6135), .Y(new_n6153));
  xor_4  g05777(.A(new_n6153), .B(new_n6129), .Y(new_n6154));
  nor_5  g05778(.A(new_n6053), .B(new_n6052), .Y(new_n6155));
  and_6  g05779(.A(new_n6054), .B(new_n6024), .Y(new_n6156));
  nor_5  g05780(.A(new_n6156), .B(new_n6155), .Y(new_n6157));
  xor_4  g05781(.A(new_n6157), .B(new_n6154), .Y(new_n6158));
  nor_5  g05782(.A(new_n6158), .B(new_n6127), .Y(new_n6159));
  or_6   g05783(.A(new_n6159), .B(new_n6126), .Y(new_n6160));
  xor_4  g05784(.A(new_n6160), .B(new_n6022), .Y(new_n6161));
  xor_4  g05785(.A(new_n6161), .B(new_n6021), .Y(new_n6162));
  nand_5 g05786(.A(pi077), .B(pi053), .Y(new_n6163));
  nor_5  g05787(.A(new_n6163), .B(new_n3511), .Y(new_n6164));
  nand_5 g05788(.A(new_n3514), .B(new_n3511), .Y(new_n6165));
  nand_5 g05789(.A(new_n3515), .B(new_n3510), .Y(new_n6166));
  nand_5 g05790(.A(new_n6166), .B(new_n6165), .Y(new_n6167));
  nand_5 g05791(.A(pi077), .B(pi067), .Y(new_n6168));
  nand_5 g05792(.A(pi053), .B(pi052), .Y(new_n6169));
  and_6  g05793(.A(new_n6169), .B(new_n6168), .Y(new_n6170));
  or_6   g05794(.A(new_n6170), .B(new_n6164), .Y(new_n6171));
  nand_5 g05795(.A(pi189), .B(pi092), .Y(new_n6172));
  nand_5 g05796(.A(pi190), .B(pi064), .Y(new_n6173));
  nand_5 g05797(.A(new_n6173), .B(new_n6172), .Y(new_n6174));
  nand_5 g05798(.A(pi092), .B(pi064), .Y(new_n6175));
  nor_5  g05799(.A(new_n6175), .B(new_n3508), .Y(new_n6176));
  not_8  g05800(.A(new_n6176), .Y(new_n6177));
  nand_5 g05801(.A(new_n6177), .B(new_n6174), .Y(new_n6178));
  nand_5 g05802(.A(pi229), .B(pi133), .Y(new_n6179));
  nand_5 g05803(.A(new_n3508), .B(new_n3507), .Y(new_n6180));
  nand_5 g05804(.A(new_n3509), .B(new_n3506), .Y(new_n6181));
  nand_5 g05805(.A(new_n6181), .B(new_n6180), .Y(new_n6182));
  xor_4  g05806(.A(new_n6182), .B(new_n6179), .Y(new_n6183));
  xor_4  g05807(.A(new_n6183), .B(new_n6178), .Y(new_n6184));
  xor_4  g05808(.A(new_n6184), .B(new_n6171), .Y(new_n6185));
  not_8  g05809(.A(new_n6185), .Y(new_n6186));
  nor_5  g05810(.A(new_n6186), .B(new_n6167), .Y(new_n6187));
  and_6  g05811(.A(new_n6187), .B(new_n6164), .Y(new_n6188));
  nand_5 g05812(.A(pi185), .B(pi052), .Y(new_n6189));
  nand_5 g05813(.A(pi131), .B(pi030), .Y(new_n6190));
  xor_4  g05814(.A(new_n6190), .B(new_n6163), .Y(new_n6191));
  xor_4  g05815(.A(new_n6191), .B(new_n6189), .Y(new_n6192));
  nand_5 g05816(.A(new_n6182), .B(new_n6179), .Y(new_n6193));
  nand_5 g05817(.A(new_n6183), .B(new_n6178), .Y(new_n6194));
  nand_5 g05818(.A(new_n6194), .B(new_n6193), .Y(new_n6195));
  xor_4  g05819(.A(new_n6195), .B(new_n6192), .Y(new_n6196));
  nand_5 g05820(.A(pi133), .B(pi067), .Y(new_n6197));
  xor_4  g05821(.A(new_n6197), .B(new_n6177), .Y(new_n6198));
  nand_5 g05822(.A(pi229), .B(pi189), .Y(new_n6199));
  nand_5 g05823(.A(pi190), .B(pi084), .Y(new_n6200));
  xor_4  g05824(.A(new_n6200), .B(new_n6199), .Y(new_n6201));
  xor_4  g05825(.A(new_n6201), .B(new_n6175), .Y(new_n6202));
  xor_4  g05826(.A(new_n6202), .B(new_n6198), .Y(new_n6203));
  xor_4  g05827(.A(new_n6203), .B(new_n6196), .Y(new_n6204));
  nor_5  g05828(.A(new_n6184), .B(new_n6171), .Y(new_n6205));
  xor_4  g05829(.A(new_n6187), .B(new_n6164), .Y(new_n6206));
  nor_5  g05830(.A(new_n6206), .B(new_n6205), .Y(new_n6207));
  nor_5  g05831(.A(new_n6207), .B(new_n6204), .Y(new_n6208));
  nor_5  g05832(.A(new_n6208), .B(new_n6188), .Y(new_n6209));
  nand_5 g05833(.A(pi130), .B(pi013), .Y(new_n6210));
  xor_4  g05834(.A(new_n6210), .B(new_n6209), .Y(new_n6211));
  nand_5 g05835(.A(pi165), .B(pi139), .Y(new_n6212));
  nand_5 g05836(.A(pi152), .B(pi065), .Y(new_n6213));
  nand_5 g05837(.A(new_n6200), .B(new_n6199), .Y(new_n6214));
  nand_5 g05838(.A(new_n6201), .B(new_n6175), .Y(new_n6215));
  nand_5 g05839(.A(new_n6215), .B(new_n6214), .Y(new_n6216));
  xnor_4 g05840(.A(new_n6216), .B(new_n6213), .Y(new_n6217));
  nand_5 g05841(.A(pi198), .B(pi035), .Y(new_n6218));
  xor_4  g05842(.A(new_n6218), .B(new_n6217), .Y(new_n6219));
  xor_4  g05843(.A(new_n6219), .B(new_n6212), .Y(new_n6220));
  xor_4  g05844(.A(new_n6220), .B(new_n6211), .Y(new_n6221));
  xor_4  g05845(.A(new_n6221), .B(new_n6162), .Y(new_n6222));
  xnor_4 g05846(.A(new_n6091), .B(new_n6090), .Y(new_n6223));
  nand_5 g05847(.A(new_n3437), .B(new_n3419), .Y(new_n6224));
  not_8  g05848(.A(new_n6224), .Y(new_n6225));
  nand_5 g05849(.A(pi168), .B(pi165), .Y(new_n6226));
  nor_5  g05850(.A(new_n3424), .B(new_n3420), .Y(new_n6227));
  and_6  g05851(.A(new_n3436), .B(new_n3425), .Y(new_n6228));
  nor_5  g05852(.A(new_n6228), .B(new_n6227), .Y(new_n6229));
  nand_5 g05853(.A(new_n3434), .B(new_n3431), .Y(new_n6230));
  nand_5 g05854(.A(new_n3435), .B(new_n3430), .Y(new_n6231));
  nand_5 g05855(.A(new_n6231), .B(new_n6230), .Y(new_n6232));
  nand_5 g05856(.A(pi172), .B(pi139), .Y(new_n6233));
  nand_5 g05857(.A(pi208), .B(pi198), .Y(new_n6234));
  nand_5 g05858(.A(new_n6234), .B(new_n6233), .Y(new_n6235));
  nand_5 g05859(.A(pi198), .B(pi139), .Y(new_n6236));
  nor_5  g05860(.A(new_n6236), .B(new_n3431), .Y(new_n6237));
  not_8  g05861(.A(new_n6237), .Y(new_n6238));
  nand_5 g05862(.A(new_n6238), .B(new_n6235), .Y(new_n6239));
  nand_5 g05863(.A(pi062), .B(pi015), .Y(new_n6240));
  nand_5 g05864(.A(pi204), .B(pi065), .Y(new_n6241));
  nand_5 g05865(.A(new_n6241), .B(new_n6240), .Y(new_n6242));
  nand_5 g05866(.A(pi204), .B(pi062), .Y(new_n6243));
  nor_5  g05867(.A(new_n6243), .B(new_n3428), .Y(new_n6244));
  not_8  g05868(.A(new_n6244), .Y(new_n6245));
  nand_5 g05869(.A(new_n6245), .B(new_n6242), .Y(new_n6246));
  nand_5 g05870(.A(pi120), .B(pi035), .Y(new_n6247));
  nand_5 g05871(.A(new_n3428), .B(new_n3427), .Y(new_n6248));
  nand_5 g05872(.A(new_n3429), .B(new_n3426), .Y(new_n6249));
  nand_5 g05873(.A(new_n6249), .B(new_n6248), .Y(new_n6250));
  xor_4  g05874(.A(new_n6250), .B(new_n6247), .Y(new_n6251));
  xor_4  g05875(.A(new_n6251), .B(new_n6246), .Y(new_n6252));
  xor_4  g05876(.A(new_n6252), .B(new_n6239), .Y(new_n6253));
  xnor_4 g05877(.A(new_n6253), .B(new_n6232), .Y(new_n6254));
  xor_4  g05878(.A(new_n6254), .B(new_n6229), .Y(new_n6255));
  xor_4  g05879(.A(new_n6255), .B(new_n6226), .Y(new_n6256));
  xor_4  g05880(.A(new_n6256), .B(new_n6225), .Y(new_n6257));
  not_8  g05881(.A(new_n6257), .Y(new_n6258));
  nor_5  g05882(.A(new_n6258), .B(new_n6223), .Y(new_n6259));
  nor_5  g05883(.A(new_n3439), .B(new_n3418), .Y(new_n6260));
  and_6  g05884(.A(new_n3484), .B(new_n3440), .Y(new_n6261));
  nor_5  g05885(.A(new_n6261), .B(new_n6260), .Y(new_n6262));
  xor_4  g05886(.A(new_n6257), .B(new_n6223), .Y(new_n6263));
  nor_5  g05887(.A(new_n6263), .B(new_n6262), .Y(new_n6264));
  or_6   g05888(.A(new_n6264), .B(new_n6259), .Y(new_n6265));
  not_8  g05889(.A(new_n6229), .Y(new_n6266));
  nand_5 g05890(.A(new_n6254), .B(new_n6266), .Y(new_n6267));
  nand_5 g05891(.A(pi172), .B(pi035), .Y(new_n6268));
  xor_4  g05892(.A(new_n6268), .B(new_n6244), .Y(new_n6269));
  nand_5 g05893(.A(pi120), .B(pi015), .Y(new_n6270));
  nand_5 g05894(.A(pi146), .B(pi065), .Y(new_n6271));
  xor_4  g05895(.A(new_n6271), .B(new_n6270), .Y(new_n6272));
  xor_4  g05896(.A(new_n6272), .B(new_n6243), .Y(new_n6273));
  xor_4  g05897(.A(new_n6273), .B(new_n6269), .Y(new_n6274));
  nand_5 g05898(.A(new_n6250), .B(new_n6247), .Y(new_n6275));
  nand_5 g05899(.A(new_n6251), .B(new_n6246), .Y(new_n6276));
  nand_5 g05900(.A(new_n6276), .B(new_n6275), .Y(new_n6277));
  nand_5 g05901(.A(pi197), .B(pi168), .Y(new_n6278));
  nand_5 g05902(.A(pi208), .B(pi165), .Y(new_n6279));
  xor_4  g05903(.A(new_n6279), .B(new_n6278), .Y(new_n6280));
  xnor_4 g05904(.A(new_n6280), .B(new_n6236), .Y(new_n6281));
  xor_4  g05905(.A(new_n6281), .B(new_n6277), .Y(new_n6282));
  xor_4  g05906(.A(new_n6282), .B(new_n6274), .Y(new_n6283));
  not_8  g05907(.A(new_n6283), .Y(new_n6284));
  nand_5 g05908(.A(new_n6252), .B(new_n6239), .Y(new_n6285));
  nand_5 g05909(.A(new_n6253), .B(new_n6232), .Y(new_n6286));
  nand_5 g05910(.A(new_n6286), .B(new_n6285), .Y(new_n6287));
  xor_4  g05911(.A(new_n6287), .B(new_n6238), .Y(new_n6288));
  xor_4  g05912(.A(new_n6288), .B(new_n6284), .Y(new_n6289));
  xor_4  g05913(.A(new_n6289), .B(new_n6267), .Y(new_n6290));
  nor_5  g05914(.A(new_n6255), .B(new_n6226), .Y(new_n6291));
  and_6  g05915(.A(new_n6256), .B(new_n6225), .Y(new_n6292));
  nor_5  g05916(.A(new_n6292), .B(new_n6291), .Y(new_n6293));
  xor_4  g05917(.A(new_n6293), .B(new_n6290), .Y(new_n6294));
  xor_4  g05918(.A(new_n6158), .B(new_n6127), .Y(new_n6295));
  xnor_4 g05919(.A(new_n6295), .B(new_n6294), .Y(new_n6296));
  xnor_4 g05920(.A(new_n6296), .B(new_n6265), .Y(new_n6297));
  nand_5 g05921(.A(new_n3525), .B(new_n3518), .Y(new_n6298));
  nand_5 g05922(.A(pi185), .B(pi131), .Y(new_n6299));
  nand_5 g05923(.A(new_n6299), .B(new_n6298), .Y(new_n6300));
  xor_4  g05924(.A(new_n6299), .B(new_n6298), .Y(new_n6301));
  xor_4  g05925(.A(new_n6186), .B(new_n6167), .Y(new_n6302));
  nor_5  g05926(.A(new_n3504), .B(new_n3486), .Y(new_n6303));
  nand_5 g05927(.A(new_n3517), .B(new_n3505), .Y(new_n6304));
  not_8  g05928(.A(new_n6304), .Y(new_n6305));
  nor_5  g05929(.A(new_n6305), .B(new_n6303), .Y(new_n6306));
  xor_4  g05930(.A(new_n6306), .B(new_n6302), .Y(new_n6307));
  nand_5 g05931(.A(new_n6307), .B(new_n6301), .Y(new_n6308));
  nand_5 g05932(.A(new_n6308), .B(new_n6300), .Y(new_n6309));
  not_8  g05933(.A(new_n6302), .Y(new_n6310));
  nor_5  g05934(.A(new_n6306), .B(new_n6310), .Y(new_n6311));
  xor_4  g05935(.A(new_n6207), .B(new_n6204), .Y(new_n6312));
  nand_5 g05936(.A(new_n6312), .B(new_n6311), .Y(new_n6313));
  or_6   g05937(.A(new_n6312), .B(new_n6311), .Y(new_n6314));
  nand_5 g05938(.A(new_n6314), .B(new_n6313), .Y(new_n6315));
  xor_4  g05939(.A(new_n6315), .B(new_n6309), .Y(new_n6316));
  nand_5 g05940(.A(new_n6316), .B(new_n6297), .Y(new_n6317));
  xor_4  g05941(.A(new_n6316), .B(new_n6297), .Y(new_n6318));
  xor_4  g05942(.A(new_n6263), .B(new_n6262), .Y(new_n6319));
  xnor_4 g05943(.A(new_n6307), .B(new_n6301), .Y(new_n6320));
  nand_5 g05944(.A(new_n6320), .B(new_n6319), .Y(new_n6321));
  xor_4  g05945(.A(new_n6320), .B(new_n6319), .Y(new_n6322));
  nor_5  g05946(.A(new_n3552), .B(new_n3526), .Y(new_n6323));
  nor_5  g05947(.A(new_n3553), .B(new_n3485), .Y(new_n6324));
  nor_5  g05948(.A(new_n6324), .B(new_n6323), .Y(new_n6325));
  nand_5 g05949(.A(new_n6325), .B(new_n6322), .Y(new_n6326));
  nand_5 g05950(.A(new_n6326), .B(new_n6321), .Y(new_n6327));
  nand_5 g05951(.A(new_n6327), .B(new_n6318), .Y(new_n6328));
  nand_5 g05952(.A(new_n6328), .B(new_n6317), .Y(new_n6329));
  nand_5 g05953(.A(new_n6271), .B(new_n6270), .Y(new_n6330));
  nand_5 g05954(.A(new_n6272), .B(new_n6243), .Y(new_n6331));
  nand_5 g05955(.A(new_n6331), .B(new_n6330), .Y(new_n6332));
  nand_5 g05956(.A(new_n6097), .B(new_n6096), .Y(new_n6333));
  nand_5 g05957(.A(new_n6098), .B(new_n6073), .Y(new_n6334));
  nand_5 g05958(.A(new_n6334), .B(new_n6333), .Y(new_n6335));
  not_8  g05959(.A(new_n6145), .Y(new_n6336));
  nor_5  g05960(.A(new_n6149), .B(new_n6336), .Y(new_n6337));
  nor_5  g05961(.A(new_n6150), .B(new_n6142), .Y(new_n6338));
  nor_5  g05962(.A(new_n6338), .B(new_n6337), .Y(new_n6339));
  nand_5 g05963(.A(new_n6147), .B(new_n6146), .Y(new_n6340));
  nand_5 g05964(.A(new_n6148), .B(new_n6047), .Y(new_n6341));
  nand_5 g05965(.A(new_n6341), .B(new_n6340), .Y(new_n6342));
  xor_4  g05966(.A(new_n6342), .B(new_n6339), .Y(new_n6343));
  xor_4  g05967(.A(new_n6343), .B(new_n6335), .Y(new_n6344));
  xor_4  g05968(.A(new_n6344), .B(new_n6332), .Y(new_n6345));
  xor_4  g05969(.A(new_n6345), .B(new_n6329), .Y(new_n6346));
  xor_4  g05970(.A(new_n6346), .B(new_n6222), .Y(new_n6347));
  and_6  g05971(.A(new_n6120), .B(new_n6095), .Y(new_n6348));
  not_8  g05972(.A(new_n6121), .Y(new_n6349));
  nor_5  g05973(.A(new_n6124), .B(new_n6349), .Y(new_n6350));
  nor_5  g05974(.A(new_n6350), .B(new_n6348), .Y(new_n6351));
  nand_5 g05975(.A(new_n6109), .B(new_n6108), .Y(new_n6352));
  nand_5 g05976(.A(new_n6110), .B(new_n6103), .Y(new_n6353));
  nand_5 g05977(.A(new_n6353), .B(new_n6352), .Y(new_n6354));
  xor_4  g05978(.A(new_n6354), .B(new_n6351), .Y(new_n6355));
  nand_5 g05979(.A(pi183), .B(pi004), .Y(new_n6356));
  nand_5 g05980(.A(pi105), .B(pi073), .Y(new_n6357));
  xor_4  g05981(.A(new_n6357), .B(new_n6356), .Y(new_n6358));
  xor_4  g05982(.A(new_n6358), .B(new_n6355), .Y(new_n6359));
  xor_4  g05983(.A(new_n6359), .B(new_n6347), .Y(new_n6360));
  nand_5 g05984(.A(pi172), .B(pi015), .Y(new_n6361));
  nand_5 g05985(.A(pi158), .B(pi018), .Y(new_n6362));
  xor_4  g05986(.A(new_n6362), .B(new_n6361), .Y(new_n6363));
  nand_5 g05987(.A(new_n6279), .B(new_n6278), .Y(new_n6364));
  nand_5 g05988(.A(new_n6280), .B(new_n6236), .Y(new_n6365));
  nand_5 g05989(.A(new_n6365), .B(new_n6364), .Y(new_n6366));
  nand_5 g05990(.A(pi213), .B(pi022), .Y(new_n6367));
  not_8  g05991(.A(new_n6119), .Y(new_n6368));
  nand_5 g05992(.A(new_n6368), .B(new_n6111), .Y(new_n6369));
  nand_5 g05993(.A(new_n6369), .B(new_n6118), .Y(new_n6370));
  xor_4  g05994(.A(new_n6370), .B(new_n6367), .Y(new_n6371));
  xor_4  g05995(.A(new_n6371), .B(new_n6366), .Y(new_n6372));
  nor_5  g05996(.A(new_n6100), .B(new_n6075), .Y(new_n6373));
  nor_5  g05997(.A(new_n6101), .B(new_n6099), .Y(new_n6374));
  or_6   g05998(.A(new_n6374), .B(new_n6373), .Y(new_n6375));
  nand_5 g05999(.A(pi236), .B(pi153), .Y(new_n6376));
  xor_4  g06000(.A(new_n6376), .B(new_n6375), .Y(new_n6377));
  nor_5  g06001(.A(new_n6268), .B(new_n6245), .Y(new_n6378));
  nor_5  g06002(.A(new_n6273), .B(new_n6269), .Y(new_n6379));
  nor_5  g06003(.A(new_n6379), .B(new_n6378), .Y(new_n6380));
  xor_4  g06004(.A(new_n6380), .B(new_n6377), .Y(new_n6381));
  xor_4  g06005(.A(new_n6381), .B(new_n6372), .Y(new_n6382));
  nand_5 g06006(.A(pi170), .B(pi088), .Y(new_n6383));
  nand_5 g06007(.A(new_n6313), .B(new_n6309), .Y(new_n6384));
  nand_5 g06008(.A(new_n6384), .B(new_n6314), .Y(new_n6385));
  xor_4  g06009(.A(new_n6385), .B(new_n6383), .Y(new_n6386));
  nand_5 g06010(.A(new_n6137), .B(new_n6136), .Y(new_n6387));
  nand_5 g06011(.A(new_n6138), .B(new_n6031), .Y(new_n6388));
  nand_5 g06012(.A(new_n6388), .B(new_n6387), .Y(new_n6389));
  nand_5 g06013(.A(pi154), .B(pi090), .Y(new_n6390));
  xnor_4 g06014(.A(new_n6390), .B(new_n6389), .Y(new_n6391));
  nand_5 g06015(.A(pi220), .B(pi131), .Y(new_n6392));
  xor_4  g06016(.A(new_n6392), .B(new_n6391), .Y(new_n6393));
  xor_4  g06017(.A(new_n6393), .B(new_n6386), .Y(new_n6394));
  nand_5 g06018(.A(pi161), .B(pi006), .Y(new_n6395));
  nand_5 g06019(.A(pi089), .B(pi047), .Y(new_n6396));
  nand_5 g06020(.A(pi254), .B(pi128), .Y(new_n6397));
  xor_4  g06021(.A(new_n6397), .B(new_n6396), .Y(new_n6398));
  nand_5 g06022(.A(pi241), .B(pi209), .Y(new_n6399));
  nand_5 g06023(.A(pi190), .B(pi034), .Y(new_n6400));
  xor_4  g06024(.A(new_n6400), .B(new_n6399), .Y(new_n6401));
  nor_5  g06025(.A(new_n6140), .B(new_n6033), .Y(new_n6402));
  nor_5  g06026(.A(new_n6141), .B(new_n6139), .Y(new_n6403));
  or_6   g06027(.A(new_n6403), .B(new_n6402), .Y(new_n6404));
  xor_4  g06028(.A(new_n6404), .B(new_n6401), .Y(new_n6405));
  xor_4  g06029(.A(new_n6405), .B(new_n6398), .Y(new_n6406));
  xor_4  g06030(.A(new_n6406), .B(new_n6395), .Y(new_n6407));
  nor_5  g06031(.A(new_n6134), .B(new_n6048), .Y(new_n6408));
  and_6  g06032(.A(new_n6152), .B(new_n6135), .Y(new_n6409));
  nor_5  g06033(.A(new_n6409), .B(new_n6408), .Y(new_n6410));
  xor_4  g06034(.A(new_n6410), .B(new_n6407), .Y(new_n6411));
  xor_4  g06035(.A(new_n6411), .B(new_n6394), .Y(new_n6412));
  xor_4  g06036(.A(new_n6412), .B(new_n6382), .Y(new_n6413));
  nor_5  g06037(.A(new_n6295), .B(new_n6294), .Y(new_n6414));
  nor_5  g06038(.A(new_n6296), .B(new_n6265), .Y(new_n6415));
  or_6   g06039(.A(new_n6415), .B(new_n6414), .Y(new_n6416));
  nand_5 g06040(.A(pi133), .B(pi053), .Y(new_n6417));
  xor_4  g06041(.A(new_n6417), .B(new_n6416), .Y(new_n6418));
  nand_5 g06042(.A(pi052), .B(pi030), .Y(new_n6419));
  not_8  g06043(.A(new_n6289), .Y(new_n6420));
  nor_5  g06044(.A(new_n6420), .B(new_n6267), .Y(new_n6421));
  nor_5  g06045(.A(new_n6293), .B(new_n6290), .Y(new_n6422));
  nor_5  g06046(.A(new_n6422), .B(new_n6421), .Y(new_n6423));
  xor_4  g06047(.A(new_n6423), .B(new_n6419), .Y(new_n6424));
  xor_4  g06048(.A(new_n6424), .B(new_n6418), .Y(new_n6425));
  xor_4  g06049(.A(new_n6425), .B(new_n6413), .Y(new_n6426));
  nand_5 g06050(.A(new_n6153), .B(new_n6129), .Y(new_n6427));
  not_8  g06051(.A(new_n6157), .Y(new_n6428));
  nand_5 g06052(.A(new_n6428), .B(new_n6154), .Y(new_n6429));
  nand_5 g06053(.A(new_n6429), .B(new_n6427), .Y(new_n6430));
  not_8  g06054(.A(new_n6277), .Y(new_n6431));
  nor_5  g06055(.A(new_n6281), .B(new_n6431), .Y(new_n6432));
  nor_5  g06056(.A(new_n6282), .B(new_n6274), .Y(new_n6433));
  nor_5  g06057(.A(new_n6433), .B(new_n6432), .Y(new_n6434));
  xor_4  g06058(.A(new_n6434), .B(new_n6430), .Y(new_n6435));
  nand_5 g06059(.A(pi124), .B(pi104), .Y(new_n6436));
  nand_5 g06060(.A(pi215), .B(pi212), .Y(new_n6437));
  xor_4  g06061(.A(new_n6437), .B(new_n6436), .Y(new_n6438));
  nand_5 g06062(.A(pi229), .B(pi064), .Y(new_n6439));
  nand_5 g06063(.A(pi112), .B(pi003), .Y(new_n6440));
  xor_4  g06064(.A(new_n6440), .B(new_n6439), .Y(new_n6441));
  xor_4  g06065(.A(new_n6441), .B(new_n6438), .Y(new_n6442));
  xor_4  g06066(.A(new_n6442), .B(new_n6435), .Y(new_n6443));
  nand_5 g06067(.A(pi185), .B(pi077), .Y(new_n6444));
  nand_5 g06068(.A(pi141), .B(pi095), .Y(new_n6445));
  xor_4  g06069(.A(new_n6445), .B(new_n6444), .Y(new_n6446));
  nand_5 g06070(.A(pi092), .B(pi084), .Y(new_n6447));
  xor_4  g06071(.A(new_n6447), .B(new_n6446), .Y(new_n6448));
  nand_5 g06072(.A(pi146), .B(pi062), .Y(new_n6449));
  nand_5 g06073(.A(pi168), .B(pi078), .Y(new_n6450));
  xor_4  g06074(.A(new_n6450), .B(new_n6449), .Y(new_n6451));
  nor_5  g06075(.A(new_n6287), .B(new_n6238), .Y(new_n6452));
  and_6  g06076(.A(new_n6288), .B(new_n6284), .Y(new_n6453));
  nor_5  g06077(.A(new_n6453), .B(new_n6452), .Y(new_n6454));
  nand_5 g06078(.A(pi204), .B(pi120), .Y(new_n6455));
  xor_4  g06079(.A(new_n6455), .B(new_n6454), .Y(new_n6456));
  xor_4  g06080(.A(new_n6456), .B(new_n6451), .Y(new_n6457));
  or_6   g06081(.A(new_n6197), .B(new_n6177), .Y(new_n6458));
  not_8  g06082(.A(new_n6202), .Y(new_n6459));
  nand_5 g06083(.A(new_n6459), .B(new_n6198), .Y(new_n6460));
  nand_5 g06084(.A(new_n6460), .B(new_n6458), .Y(new_n6461));
  nand_5 g06085(.A(new_n6190), .B(new_n6163), .Y(new_n6462));
  nand_5 g06086(.A(new_n6191), .B(new_n6189), .Y(new_n6463));
  nand_5 g06087(.A(new_n6463), .B(new_n6462), .Y(new_n6464));
  nand_5 g06088(.A(pi189), .B(pi067), .Y(new_n6465));
  nand_5 g06089(.A(new_n6195), .B(new_n6192), .Y(new_n6466));
  nand_5 g06090(.A(new_n6203), .B(new_n6196), .Y(new_n6467));
  nand_5 g06091(.A(new_n6467), .B(new_n6466), .Y(new_n6468));
  xnor_4 g06092(.A(new_n6468), .B(new_n6465), .Y(new_n6469));
  xor_4  g06093(.A(new_n6469), .B(new_n6464), .Y(new_n6470));
  xor_4  g06094(.A(new_n6470), .B(new_n6461), .Y(new_n6471));
  xor_4  g06095(.A(new_n6471), .B(new_n6457), .Y(new_n6472));
  xor_4  g06096(.A(new_n6472), .B(new_n6448), .Y(new_n6473));
  xor_4  g06097(.A(new_n6473), .B(new_n6443), .Y(new_n6474));
  xor_4  g06098(.A(new_n6474), .B(new_n6426), .Y(new_n6475));
  xor_4  g06099(.A(new_n6475), .B(new_n6363), .Y(new_n6476));
  xor_4  g06100(.A(new_n6476), .B(new_n6360), .Y(po027));
  nand_5 g06101(.A(new_n4808), .B(new_n4790), .Y(new_n6478));
  nand_5 g06102(.A(pi131), .B(pi036), .Y(new_n6479));
  xor_4  g06103(.A(new_n6479), .B(new_n6478), .Y(new_n6480));
  not_8  g06104(.A(new_n6480), .Y(new_n6481));
  nor_5  g06105(.A(new_n4806), .B(new_n4795), .Y(new_n6482));
  nor_5  g06106(.A(new_n4807), .B(new_n4794), .Y(new_n6483));
  nor_5  g06107(.A(new_n6483), .B(new_n6482), .Y(new_n6484));
  nand_5 g06108(.A(new_n4804), .B(new_n4801), .Y(new_n6485));
  nand_5 g06109(.A(new_n4805), .B(new_n4800), .Y(new_n6486));
  nand_5 g06110(.A(new_n6486), .B(new_n6485), .Y(new_n6487));
  nand_5 g06111(.A(pi085), .B(pi077), .Y(new_n6488));
  nand_5 g06112(.A(pi180), .B(pi052), .Y(new_n6489));
  and_6  g06113(.A(new_n6489), .B(new_n6488), .Y(new_n6490));
  nand_5 g06114(.A(pi180), .B(pi077), .Y(new_n6491));
  nor_5  g06115(.A(new_n6491), .B(new_n4801), .Y(new_n6492));
  or_6   g06116(.A(new_n6492), .B(new_n6490), .Y(new_n6493));
  nand_5 g06117(.A(new_n4798), .B(new_n4797), .Y(new_n6494));
  nand_5 g06118(.A(new_n4799), .B(new_n4796), .Y(new_n6495));
  nand_5 g06119(.A(new_n6495), .B(new_n6494), .Y(new_n6496));
  nand_5 g06120(.A(pi194), .B(pi133), .Y(new_n6497));
  nand_5 g06121(.A(pi143), .B(pi064), .Y(new_n6498));
  nand_5 g06122(.A(pi189), .B(pi057), .Y(new_n6499));
  nand_5 g06123(.A(new_n6499), .B(new_n6498), .Y(new_n6500));
  nand_5 g06124(.A(pi064), .B(pi057), .Y(new_n6501));
  nor_5  g06125(.A(new_n6501), .B(new_n4797), .Y(new_n6502));
  not_8  g06126(.A(new_n6502), .Y(new_n6503));
  nand_5 g06127(.A(new_n6503), .B(new_n6500), .Y(new_n6504));
  xor_4  g06128(.A(new_n6504), .B(new_n6497), .Y(new_n6505));
  xor_4  g06129(.A(new_n6505), .B(new_n6496), .Y(new_n6506));
  xor_4  g06130(.A(new_n6506), .B(new_n6493), .Y(new_n6507));
  xor_4  g06131(.A(new_n6507), .B(new_n6487), .Y(new_n6508));
  xor_4  g06132(.A(new_n6508), .B(new_n6484), .Y(new_n6509));
  xor_4  g06133(.A(new_n6509), .B(new_n6481), .Y(new_n6510));
  nand_5 g06134(.A(new_n4883), .B(new_n4809), .Y(new_n6511));
  nand_5 g06135(.A(new_n4884), .B(new_n4789), .Y(new_n6512));
  nand_5 g06136(.A(new_n6512), .B(new_n6511), .Y(new_n6513));
  xor_4  g06137(.A(new_n6513), .B(new_n6510), .Y(new_n6514));
  or_6   g06138(.A(new_n4881), .B(new_n4878), .Y(new_n6515));
  nand_5 g06139(.A(new_n4882), .B(new_n4857), .Y(new_n6516));
  nand_5 g06140(.A(new_n6516), .B(new_n6515), .Y(new_n6517));
  nand_5 g06141(.A(new_n4877), .B(new_n4858), .Y(new_n6518));
  nand_5 g06142(.A(pi238), .B(pi168), .Y(new_n6519));
  xor_4  g06143(.A(new_n6519), .B(new_n6518), .Y(new_n6520));
  nand_5 g06144(.A(new_n4873), .B(new_n4870), .Y(new_n6521));
  nand_5 g06145(.A(new_n4874), .B(new_n4869), .Y(new_n6522));
  nand_5 g06146(.A(new_n6522), .B(new_n6521), .Y(new_n6523));
  nand_5 g06147(.A(pi139), .B(pi048), .Y(new_n6524));
  nand_5 g06148(.A(pi237), .B(pi208), .Y(new_n6525));
  and_6  g06149(.A(new_n6525), .B(new_n6524), .Y(new_n6526));
  nand_5 g06150(.A(pi237), .B(pi139), .Y(new_n6527));
  nor_5  g06151(.A(new_n6527), .B(new_n4870), .Y(new_n6528));
  or_6   g06152(.A(new_n6528), .B(new_n6526), .Y(new_n6529));
  nand_5 g06153(.A(new_n4867), .B(new_n4866), .Y(new_n6530));
  nand_5 g06154(.A(new_n4868), .B(new_n4865), .Y(new_n6531));
  nand_5 g06155(.A(new_n6531), .B(new_n6530), .Y(new_n6532));
  nand_5 g06156(.A(pi179), .B(pi035), .Y(new_n6533));
  nand_5 g06157(.A(pi033), .B(pi015), .Y(new_n6534));
  nand_5 g06158(.A(pi204), .B(pi162), .Y(new_n6535));
  nand_5 g06159(.A(new_n6535), .B(new_n6534), .Y(new_n6536));
  nand_5 g06160(.A(pi204), .B(pi033), .Y(new_n6537));
  nor_5  g06161(.A(new_n6537), .B(new_n4867), .Y(new_n6538));
  not_8  g06162(.A(new_n6538), .Y(new_n6539));
  nand_5 g06163(.A(new_n6539), .B(new_n6536), .Y(new_n6540));
  xor_4  g06164(.A(new_n6540), .B(new_n6533), .Y(new_n6541));
  xor_4  g06165(.A(new_n6541), .B(new_n6532), .Y(new_n6542));
  xor_4  g06166(.A(new_n6542), .B(new_n6529), .Y(new_n6543));
  not_8  g06167(.A(new_n6543), .Y(new_n6544));
  xor_4  g06168(.A(new_n6544), .B(new_n6523), .Y(new_n6545));
  nor_5  g06169(.A(new_n4863), .B(new_n4859), .Y(new_n6546));
  nand_5 g06170(.A(new_n4876), .B(new_n4864), .Y(new_n6547));
  not_8  g06171(.A(new_n6547), .Y(new_n6548));
  nor_5  g06172(.A(new_n6548), .B(new_n6546), .Y(new_n6549));
  xor_4  g06173(.A(new_n6549), .B(new_n6545), .Y(new_n6550));
  xor_4  g06174(.A(new_n6550), .B(new_n6520), .Y(new_n6551));
  xnor_4 g06175(.A(new_n6551), .B(new_n6517), .Y(new_n6552));
  or_6   g06176(.A(new_n4829), .B(new_n4812), .Y(new_n6553));
  or_6   g06177(.A(new_n4827), .B(new_n4824), .Y(new_n6554));
  not_8  g06178(.A(new_n4828), .Y(new_n6555));
  or_6   g06179(.A(new_n6555), .B(new_n4823), .Y(new_n6556));
  and_6  g06180(.A(new_n6556), .B(new_n6554), .Y(new_n6557));
  nand_5 g06181(.A(new_n4821), .B(new_n4818), .Y(new_n6558));
  nand_5 g06182(.A(new_n4822), .B(new_n4817), .Y(new_n6559));
  nand_5 g06183(.A(new_n6559), .B(new_n6558), .Y(new_n6560));
  nand_5 g06184(.A(pi104), .B(pi012), .Y(new_n6561));
  nand_5 g06185(.A(pi212), .B(pi144), .Y(new_n6562));
  and_6  g06186(.A(new_n6562), .B(new_n6561), .Y(new_n6563));
  nand_5 g06187(.A(pi144), .B(pi104), .Y(new_n6564));
  nor_5  g06188(.A(new_n6564), .B(new_n4818), .Y(new_n6565));
  or_6   g06189(.A(new_n6565), .B(new_n6563), .Y(new_n6566));
  nand_5 g06190(.A(new_n4815), .B(new_n4814), .Y(new_n6567));
  nand_5 g06191(.A(new_n4816), .B(new_n4813), .Y(new_n6568));
  nand_5 g06192(.A(new_n6568), .B(new_n6567), .Y(new_n6569));
  nand_5 g06193(.A(pi061), .B(pi013), .Y(new_n6570));
  nand_5 g06194(.A(pi188), .B(pi105), .Y(new_n6571));
  nand_5 g06195(.A(pi178), .B(pi112), .Y(new_n6572));
  nand_5 g06196(.A(new_n6572), .B(new_n6571), .Y(new_n6573));
  nand_5 g06197(.A(pi178), .B(pi105), .Y(new_n6574));
  nor_5  g06198(.A(new_n6574), .B(new_n4813), .Y(new_n6575));
  not_8  g06199(.A(new_n6575), .Y(new_n6576));
  nand_5 g06200(.A(new_n6576), .B(new_n6573), .Y(new_n6577));
  xor_4  g06201(.A(new_n6577), .B(new_n6570), .Y(new_n6578));
  xor_4  g06202(.A(new_n6578), .B(new_n6569), .Y(new_n6579));
  xor_4  g06203(.A(new_n6579), .B(new_n6566), .Y(new_n6580));
  xor_4  g06204(.A(new_n6580), .B(new_n6560), .Y(new_n6581));
  xnor_4 g06205(.A(new_n6581), .B(new_n6557), .Y(new_n6582));
  nand_5 g06206(.A(pi213), .B(pi098), .Y(new_n6583));
  xor_4  g06207(.A(new_n6583), .B(new_n6582), .Y(new_n6584));
  xnor_4 g06208(.A(new_n6584), .B(new_n6553), .Y(new_n6585));
  nand_5 g06209(.A(new_n4850), .B(new_n4832), .Y(new_n6586));
  nand_5 g06210(.A(pi236), .B(pi113), .Y(new_n6587));
  xor_4  g06211(.A(new_n6587), .B(new_n6586), .Y(new_n6588));
  nand_5 g06212(.A(new_n4846), .B(new_n4843), .Y(new_n6589));
  nand_5 g06213(.A(new_n4847), .B(new_n4842), .Y(new_n6590));
  nand_5 g06214(.A(new_n6590), .B(new_n6589), .Y(new_n6591));
  nand_5 g06215(.A(pi141), .B(pi108), .Y(new_n6592));
  nand_5 g06216(.A(new_n4840), .B(new_n4839), .Y(new_n6593));
  nand_5 g06217(.A(new_n4841), .B(new_n4838), .Y(new_n6594));
  nand_5 g06218(.A(new_n6594), .B(new_n6593), .Y(new_n6595));
  xnor_4 g06219(.A(new_n6595), .B(new_n6592), .Y(new_n6596));
  nand_5 g06220(.A(pi090), .B(pi042), .Y(new_n6597));
  nand_5 g06221(.A(pi051), .B(pi047), .Y(new_n6598));
  nand_5 g06222(.A(new_n6598), .B(new_n6597), .Y(new_n6599));
  nand_5 g06223(.A(pi047), .B(pi042), .Y(new_n6600));
  nor_5  g06224(.A(new_n6600), .B(new_n4840), .Y(new_n6601));
  not_8  g06225(.A(new_n6601), .Y(new_n6602));
  nand_5 g06226(.A(new_n6602), .B(new_n6599), .Y(new_n6603));
  xor_4  g06227(.A(new_n6603), .B(new_n6596), .Y(new_n6604));
  nand_5 g06228(.A(pi161), .B(pi007), .Y(new_n6605));
  nand_5 g06229(.A(pi241), .B(pi118), .Y(new_n6606));
  and_6  g06230(.A(new_n6606), .B(new_n6605), .Y(new_n6607));
  nand_5 g06231(.A(pi161), .B(pi118), .Y(new_n6608));
  nor_5  g06232(.A(new_n6608), .B(new_n4843), .Y(new_n6609));
  or_6   g06233(.A(new_n6609), .B(new_n6607), .Y(new_n6610));
  xor_4  g06234(.A(new_n6610), .B(new_n6604), .Y(new_n6611));
  xor_4  g06235(.A(new_n6611), .B(new_n6591), .Y(new_n6612));
  nor_5  g06236(.A(new_n4836), .B(new_n4833), .Y(new_n6613));
  and_6  g06237(.A(new_n4849), .B(new_n4837), .Y(new_n6614));
  nor_5  g06238(.A(new_n6614), .B(new_n6613), .Y(new_n6615));
  xor_4  g06239(.A(new_n6615), .B(new_n6612), .Y(new_n6616));
  xnor_4 g06240(.A(new_n6616), .B(new_n6588), .Y(new_n6617));
  xor_4  g06241(.A(new_n6617), .B(new_n6585), .Y(new_n6618));
  nand_5 g06242(.A(new_n4851), .B(new_n4830), .Y(new_n6619));
  not_8  g06243(.A(new_n6619), .Y(new_n6620));
  nor_5  g06244(.A(new_n4856), .B(new_n4852), .Y(new_n6621));
  nor_5  g06245(.A(new_n6621), .B(new_n6620), .Y(new_n6622));
  xor_4  g06246(.A(new_n6622), .B(new_n6618), .Y(new_n6623));
  xor_4  g06247(.A(new_n6623), .B(new_n6552), .Y(new_n6624));
  xnor_4 g06248(.A(new_n6624), .B(new_n6514), .Y(po028));
  xnor_4 g06249(.A(new_n884), .B(new_n883), .Y(po029));
  xor_4  g06250(.A(new_n1457), .B(new_n1456), .Y(po030));
  nand_5 g06251(.A(pi217), .B(pi103), .Y(new_n6628));
  nand_5 g06252(.A(pi249), .B(pi175), .Y(new_n6629));
  not_8  g06253(.A(new_n6629), .Y(new_n6630));
  nand_5 g06254(.A(pi242), .B(pi107), .Y(new_n6631));
  nand_5 g06255(.A(pi210), .B(pi163), .Y(new_n6632));
  not_8  g06256(.A(new_n6632), .Y(new_n6633));
  xor_4  g06257(.A(new_n6633), .B(new_n6631), .Y(new_n6634));
  xor_4  g06258(.A(new_n6634), .B(new_n6630), .Y(new_n6635));
  xor_4  g06259(.A(new_n6635), .B(new_n6628), .Y(po031));
  xnor_4 g06260(.A(new_n2579), .B(new_n2578), .Y(po032));
  nor_5  g06261(.A(new_n6634), .B(new_n6629), .Y(new_n6638));
  nand_5 g06262(.A(pi249), .B(pi134), .Y(new_n6639));
  nand_5 g06263(.A(pi222), .B(pi175), .Y(new_n6640));
  xor_4  g06264(.A(new_n6640), .B(new_n6639), .Y(new_n6641));
  or_6   g06265(.A(new_n6641), .B(new_n6638), .Y(new_n6642));
  xor_4  g06266(.A(new_n6641), .B(new_n6638), .Y(new_n6643));
  nand_5 g06267(.A(pi171), .B(pi140), .Y(new_n6644));
  or_6   g06268(.A(new_n6644), .B(new_n6631), .Y(new_n6645));
  nand_5 g06269(.A(pi140), .B(pi107), .Y(new_n6646));
  nand_5 g06270(.A(pi242), .B(pi171), .Y(new_n6647));
  nand_5 g06271(.A(new_n6647), .B(new_n6646), .Y(new_n6648));
  nand_5 g06272(.A(new_n6648), .B(new_n6645), .Y(new_n6649));
  or_6   g06273(.A(new_n6632), .B(new_n6631), .Y(new_n6650));
  nand_5 g06274(.A(pi210), .B(pi148), .Y(new_n6651));
  nand_5 g06275(.A(pi163), .B(pi111), .Y(new_n6652));
  nand_5 g06276(.A(new_n6652), .B(new_n6651), .Y(new_n6653));
  nand_5 g06277(.A(pi148), .B(pi111), .Y(new_n6654));
  or_6   g06278(.A(new_n6654), .B(new_n6632), .Y(new_n6655));
  nand_5 g06279(.A(new_n6655), .B(new_n6653), .Y(new_n6656));
  xnor_4 g06280(.A(new_n6656), .B(new_n6650), .Y(new_n6657));
  xnor_4 g06281(.A(new_n6657), .B(new_n6649), .Y(new_n6658));
  nand_5 g06282(.A(new_n6658), .B(new_n6643), .Y(new_n6659));
  nand_5 g06283(.A(new_n6659), .B(new_n6642), .Y(new_n6660));
  nand_5 g06284(.A(pi222), .B(pi134), .Y(new_n6661));
  nor_5  g06285(.A(new_n6661), .B(new_n6630), .Y(new_n6662));
  nand_5 g06286(.A(pi249), .B(pi240), .Y(new_n6663));
  nand_5 g06287(.A(pi175), .B(pi125), .Y(new_n6664));
  or_6   g06288(.A(new_n6664), .B(new_n6663), .Y(new_n6665));
  nand_5 g06289(.A(new_n6664), .B(new_n6663), .Y(new_n6666));
  and_6  g06290(.A(new_n6666), .B(new_n6665), .Y(new_n6667));
  or_6   g06291(.A(new_n6667), .B(new_n6662), .Y(new_n6668));
  nand_5 g06292(.A(new_n6662), .B(new_n6666), .Y(new_n6669));
  nand_5 g06293(.A(new_n6669), .B(new_n6668), .Y(new_n6670));
  xor_4  g06294(.A(new_n6670), .B(new_n6660), .Y(new_n6671));
  nand_5 g06295(.A(pi242), .B(pi049), .Y(new_n6672));
  nand_5 g06296(.A(pi252), .B(pi107), .Y(new_n6673));
  xor_4  g06297(.A(new_n6673), .B(new_n6644), .Y(new_n6674));
  xor_4  g06298(.A(new_n6674), .B(new_n6672), .Y(new_n6675));
  xnor_4 g06299(.A(new_n6675), .B(new_n6645), .Y(new_n6676));
  nor_5  g06300(.A(new_n6654), .B(new_n6633), .Y(new_n6677));
  nand_5 g06301(.A(pi228), .B(pi210), .Y(new_n6678));
  nand_5 g06302(.A(pi163), .B(pi024), .Y(new_n6679));
  nand_5 g06303(.A(new_n6679), .B(new_n6678), .Y(new_n6680));
  or_6   g06304(.A(new_n6679), .B(new_n6678), .Y(new_n6681));
  and_6  g06305(.A(new_n6681), .B(new_n6680), .Y(new_n6682));
  or_6   g06306(.A(new_n6682), .B(new_n6677), .Y(new_n6683));
  nand_5 g06307(.A(new_n6680), .B(new_n6677), .Y(new_n6684));
  nand_5 g06308(.A(new_n6684), .B(new_n6683), .Y(new_n6685));
  xnor_4 g06309(.A(new_n6685), .B(new_n6676), .Y(new_n6686));
  nor_5  g06310(.A(new_n6656), .B(new_n6650), .Y(new_n6687));
  nor_5  g06311(.A(new_n6657), .B(new_n6649), .Y(new_n6688));
  nor_5  g06312(.A(new_n6688), .B(new_n6687), .Y(new_n6689));
  xnor_4 g06313(.A(new_n6689), .B(new_n6686), .Y(new_n6690));
  xor_4  g06314(.A(new_n6690), .B(new_n6671), .Y(new_n6691));
  or_6   g06315(.A(new_n6635), .B(new_n6628), .Y(new_n6692));
  not_8  g06316(.A(new_n6628), .Y(new_n6693));
  nand_5 g06317(.A(pi117), .B(pi100), .Y(new_n6694));
  not_8  g06318(.A(new_n6694), .Y(new_n6695));
  nand_5 g06319(.A(new_n6695), .B(new_n6693), .Y(new_n6696));
  nand_5 g06320(.A(pi103), .B(pi100), .Y(new_n6697));
  nand_5 g06321(.A(pi217), .B(pi117), .Y(new_n6698));
  nand_5 g06322(.A(new_n6698), .B(new_n6697), .Y(new_n6699));
  nand_5 g06323(.A(new_n6699), .B(new_n6696), .Y(new_n6700));
  nor_5  g06324(.A(new_n6700), .B(new_n6692), .Y(new_n6701));
  xor_4  g06325(.A(new_n6700), .B(new_n6692), .Y(new_n6702));
  xor_4  g06326(.A(new_n6658), .B(new_n6643), .Y(new_n6703));
  not_8  g06327(.A(new_n6703), .Y(new_n6704));
  and_6  g06328(.A(new_n6704), .B(new_n6702), .Y(new_n6705));
  nor_5  g06329(.A(new_n6705), .B(new_n6701), .Y(new_n6706));
  nand_5 g06330(.A(pi227), .B(pi103), .Y(new_n6707));
  nand_5 g06331(.A(pi217), .B(pi016), .Y(new_n6708));
  nor_5  g06332(.A(new_n6708), .B(new_n6707), .Y(new_n6709));
  nand_5 g06333(.A(new_n6708), .B(new_n6707), .Y(new_n6710));
  nor_5  g06334(.A(new_n6694), .B(new_n6693), .Y(new_n6711));
  nor_5  g06335(.A(new_n6711), .B(new_n6710), .Y(new_n6712));
  nor_5  g06336(.A(new_n6712), .B(new_n6709), .Y(new_n6713));
  nand_5 g06337(.A(new_n6711), .B(new_n6710), .Y(new_n6714));
  nand_5 g06338(.A(new_n6714), .B(new_n6713), .Y(new_n6715));
  xor_4  g06339(.A(new_n6715), .B(new_n6706), .Y(new_n6716));
  xnor_4 g06340(.A(new_n6716), .B(new_n6691), .Y(po033));
  xnor_4 g06341(.A(new_n4568), .B(new_n4567), .Y(po034));
  xor_4  g06342(.A(new_n4252), .B(new_n4251), .Y(po035));
  nand_5 g06343(.A(pi233), .B(pi103), .Y(new_n6720));
  nand_5 g06344(.A(pi103), .B(pi081), .Y(new_n6721));
  or_6   g06345(.A(new_n6709), .B(new_n6695), .Y(new_n6722));
  nand_5 g06346(.A(new_n6722), .B(new_n6710), .Y(new_n6723));
  or_6   g06347(.A(new_n6723), .B(new_n6721), .Y(new_n6724));
  xor_4  g06348(.A(new_n6723), .B(new_n6721), .Y(new_n6725));
  nand_5 g06349(.A(pi227), .B(pi117), .Y(new_n6726));
  nand_5 g06350(.A(pi100), .B(pi016), .Y(new_n6727));
  nand_5 g06351(.A(pi217), .B(pi080), .Y(new_n6728));
  xor_4  g06352(.A(new_n6728), .B(new_n6727), .Y(new_n6729));
  xor_4  g06353(.A(new_n6729), .B(new_n6726), .Y(new_n6730));
  not_8  g06354(.A(new_n6730), .Y(new_n6731));
  nand_5 g06355(.A(new_n6731), .B(new_n6725), .Y(new_n6732));
  nand_5 g06356(.A(new_n6732), .B(new_n6724), .Y(new_n6733));
  nand_5 g06357(.A(pi106), .B(pi103), .Y(new_n6734));
  nand_5 g06358(.A(pi247), .B(pi217), .Y(new_n6735));
  nand_5 g06359(.A(pi227), .B(pi016), .Y(new_n6736));
  nand_5 g06360(.A(pi100), .B(pi080), .Y(new_n6737));
  xor_4  g06361(.A(new_n6737), .B(new_n6736), .Y(new_n6738));
  xor_4  g06362(.A(new_n6738), .B(new_n6735), .Y(new_n6739));
  nand_5 g06363(.A(pi117), .B(pi081), .Y(new_n6740));
  nand_5 g06364(.A(new_n6728), .B(new_n6727), .Y(new_n6741));
  nand_5 g06365(.A(new_n6729), .B(new_n6726), .Y(new_n6742));
  nand_5 g06366(.A(new_n6742), .B(new_n6741), .Y(new_n6743));
  xor_4  g06367(.A(new_n6743), .B(new_n6740), .Y(new_n6744));
  xor_4  g06368(.A(new_n6744), .B(new_n6739), .Y(new_n6745));
  xor_4  g06369(.A(new_n6745), .B(new_n6734), .Y(new_n6746));
  xor_4  g06370(.A(new_n6746), .B(new_n6733), .Y(new_n6747));
  nor_5  g06371(.A(new_n6713), .B(new_n6696), .Y(new_n6748));
  xor_4  g06372(.A(new_n6731), .B(new_n6725), .Y(new_n6749));
  nand_5 g06373(.A(new_n6749), .B(new_n6748), .Y(new_n6750));
  not_8  g06374(.A(new_n6750), .Y(new_n6751));
  nand_5 g06375(.A(new_n6751), .B(new_n6747), .Y(new_n6752));
  nand_5 g06376(.A(new_n6752), .B(new_n6720), .Y(new_n6753));
  xor_4  g06377(.A(new_n6752), .B(new_n6720), .Y(new_n6754));
  nor_5  g06378(.A(new_n6745), .B(new_n6734), .Y(new_n6755));
  nand_5 g06379(.A(new_n6746), .B(new_n6733), .Y(new_n6756));
  not_8  g06380(.A(new_n6756), .Y(new_n6757));
  nor_5  g06381(.A(new_n6757), .B(new_n6755), .Y(new_n6758));
  nand_5 g06382(.A(new_n6743), .B(new_n6740), .Y(new_n6759));
  nand_5 g06383(.A(new_n6744), .B(new_n6739), .Y(new_n6760));
  nand_5 g06384(.A(new_n6760), .B(new_n6759), .Y(new_n6761));
  nand_5 g06385(.A(pi081), .B(pi016), .Y(new_n6762));
  nand_5 g06386(.A(pi117), .B(pi106), .Y(new_n6763));
  and_6  g06387(.A(new_n6763), .B(new_n6762), .Y(new_n6764));
  nand_5 g06388(.A(pi106), .B(pi016), .Y(new_n6765));
  nor_5  g06389(.A(new_n6765), .B(new_n6740), .Y(new_n6766));
  or_6   g06390(.A(new_n6766), .B(new_n6764), .Y(new_n6767));
  nand_5 g06391(.A(new_n6737), .B(new_n6736), .Y(new_n6768));
  nand_5 g06392(.A(new_n6738), .B(new_n6735), .Y(new_n6769));
  nand_5 g06393(.A(new_n6769), .B(new_n6768), .Y(new_n6770));
  nand_5 g06394(.A(pi234), .B(pi217), .Y(new_n6771));
  nand_5 g06395(.A(pi247), .B(pi100), .Y(new_n6772));
  nand_5 g06396(.A(new_n6772), .B(new_n6771), .Y(new_n6773));
  nand_5 g06397(.A(pi234), .B(pi100), .Y(new_n6774));
  nor_5  g06398(.A(new_n6774), .B(new_n6735), .Y(new_n6775));
  not_8  g06399(.A(new_n6775), .Y(new_n6776));
  nand_5 g06400(.A(new_n6776), .B(new_n6773), .Y(new_n6777));
  nand_5 g06401(.A(pi227), .B(pi080), .Y(new_n6778));
  xor_4  g06402(.A(new_n6778), .B(new_n6777), .Y(new_n6779));
  xor_4  g06403(.A(new_n6779), .B(new_n6770), .Y(new_n6780));
  xor_4  g06404(.A(new_n6780), .B(new_n6767), .Y(new_n6781));
  xor_4  g06405(.A(new_n6781), .B(new_n6761), .Y(new_n6782));
  xor_4  g06406(.A(new_n6782), .B(new_n6758), .Y(new_n6783));
  not_8  g06407(.A(new_n6783), .Y(new_n6784));
  nand_5 g06408(.A(new_n6784), .B(new_n6754), .Y(new_n6785));
  nand_5 g06409(.A(new_n6785), .B(new_n6753), .Y(new_n6786));
  nor_5  g06410(.A(new_n6782), .B(new_n6758), .Y(new_n6787));
  not_8  g06411(.A(new_n6781), .Y(new_n6788));
  nor_5  g06412(.A(new_n6788), .B(new_n6761), .Y(new_n6789));
  nand_5 g06413(.A(new_n6789), .B(new_n6766), .Y(new_n6790));
  nor_5  g06414(.A(new_n6780), .B(new_n6767), .Y(new_n6791));
  nor_5  g06415(.A(new_n6791), .B(new_n6766), .Y(new_n6792));
  not_8  g06416(.A(new_n6792), .Y(new_n6793));
  nor_5  g06417(.A(new_n6793), .B(new_n6789), .Y(new_n6794));
  not_8  g06418(.A(new_n6794), .Y(new_n6795));
  nand_5 g06419(.A(new_n6795), .B(new_n6790), .Y(new_n6796));
  nand_5 g06420(.A(new_n6778), .B(new_n6777), .Y(new_n6797));
  nand_5 g06421(.A(new_n6779), .B(new_n6770), .Y(new_n6798));
  nand_5 g06422(.A(new_n6798), .B(new_n6797), .Y(new_n6799));
  nand_5 g06423(.A(pi233), .B(pi117), .Y(new_n6800));
  nand_5 g06424(.A(pi187), .B(pi103), .Y(new_n6801));
  xor_4  g06425(.A(new_n6801), .B(new_n6800), .Y(new_n6802));
  xor_4  g06426(.A(new_n6802), .B(new_n6765), .Y(new_n6803));
  xor_4  g06427(.A(new_n6803), .B(new_n6799), .Y(new_n6804));
  nand_5 g06428(.A(pi081), .B(pi080), .Y(new_n6805));
  xor_4  g06429(.A(new_n6805), .B(new_n6775), .Y(new_n6806));
  nand_5 g06430(.A(pi217), .B(pi214), .Y(new_n6807));
  nand_5 g06431(.A(pi247), .B(pi227), .Y(new_n6808));
  xor_4  g06432(.A(new_n6808), .B(new_n6807), .Y(new_n6809));
  xor_4  g06433(.A(new_n6809), .B(new_n6774), .Y(new_n6810));
  xnor_4 g06434(.A(new_n6810), .B(new_n6806), .Y(new_n6811));
  xor_4  g06435(.A(new_n6811), .B(new_n6804), .Y(new_n6812));
  not_8  g06436(.A(new_n6812), .Y(new_n6813));
  xor_4  g06437(.A(new_n6813), .B(new_n6796), .Y(new_n6814));
  xor_4  g06438(.A(new_n6814), .B(new_n6787), .Y(new_n6815));
  xor_4  g06439(.A(new_n6815), .B(new_n6786), .Y(new_n6816));
  xor_4  g06440(.A(new_n6783), .B(new_n6754), .Y(new_n6817));
  nor_5  g06441(.A(new_n6685), .B(new_n6676), .Y(new_n6818));
  nor_5  g06442(.A(new_n6689), .B(new_n6686), .Y(new_n6819));
  nor_5  g06443(.A(new_n6819), .B(new_n6818), .Y(new_n6820));
  nor_5  g06444(.A(new_n6675), .B(new_n6645), .Y(new_n6821));
  nand_5 g06445(.A(pi121), .B(pi107), .Y(new_n6822));
  nand_5 g06446(.A(new_n6673), .B(new_n6644), .Y(new_n6823));
  nand_5 g06447(.A(new_n6674), .B(new_n6672), .Y(new_n6824));
  nand_5 g06448(.A(new_n6824), .B(new_n6823), .Y(new_n6825));
  xor_4  g06449(.A(new_n6825), .B(new_n6822), .Y(new_n6826));
  nand_5 g06450(.A(pi252), .B(pi171), .Y(new_n6827));
  nand_5 g06451(.A(pi245), .B(pi242), .Y(new_n6828));
  nand_5 g06452(.A(pi140), .B(pi049), .Y(new_n6829));
  xor_4  g06453(.A(new_n6829), .B(new_n6828), .Y(new_n6830));
  xor_4  g06454(.A(new_n6830), .B(new_n6827), .Y(new_n6831));
  not_8  g06455(.A(new_n6831), .Y(new_n6832));
  xor_4  g06456(.A(new_n6832), .B(new_n6826), .Y(new_n6833));
  xnor_4 g06457(.A(new_n6833), .B(new_n6821), .Y(new_n6834));
  nand_5 g06458(.A(new_n6834), .B(new_n6820), .Y(new_n6835));
  xor_4  g06459(.A(new_n6834), .B(new_n6820), .Y(new_n6836));
  nand_5 g06460(.A(pi210), .B(pi039), .Y(new_n6837));
  nand_5 g06461(.A(pi228), .B(pi111), .Y(new_n6838));
  nand_5 g06462(.A(pi148), .B(pi024), .Y(new_n6839));
  xor_4  g06463(.A(new_n6839), .B(new_n6838), .Y(new_n6840));
  xor_4  g06464(.A(new_n6840), .B(new_n6837), .Y(new_n6841));
  nand_5 g06465(.A(new_n6681), .B(new_n6654), .Y(new_n6842));
  nand_5 g06466(.A(new_n6842), .B(new_n6680), .Y(new_n6843));
  nand_5 g06467(.A(pi224), .B(pi163), .Y(new_n6844));
  xor_4  g06468(.A(new_n6844), .B(new_n6843), .Y(new_n6845));
  xor_4  g06469(.A(new_n6845), .B(new_n6841), .Y(new_n6846));
  nor_5  g06470(.A(new_n6682), .B(new_n6655), .Y(new_n6847));
  xor_4  g06471(.A(new_n6847), .B(new_n6846), .Y(new_n6848));
  nand_5 g06472(.A(new_n6848), .B(new_n6836), .Y(new_n6849));
  nand_5 g06473(.A(new_n6849), .B(new_n6835), .Y(new_n6850));
  not_8  g06474(.A(new_n6847), .Y(new_n6851));
  nor_5  g06475(.A(new_n6851), .B(new_n6846), .Y(new_n6852));
  nand_5 g06476(.A(pi255), .B(pi163), .Y(new_n6853));
  nand_5 g06477(.A(new_n6844), .B(new_n6843), .Y(new_n6854));
  nand_5 g06478(.A(new_n6845), .B(new_n6841), .Y(new_n6855));
  nand_5 g06479(.A(new_n6855), .B(new_n6854), .Y(new_n6856));
  xor_4  g06480(.A(new_n6856), .B(new_n6853), .Y(new_n6857));
  nand_5 g06481(.A(pi210), .B(pi116), .Y(new_n6858));
  nand_5 g06482(.A(pi228), .B(pi024), .Y(new_n6859));
  nand_5 g06483(.A(pi111), .B(pi039), .Y(new_n6860));
  xor_4  g06484(.A(new_n6860), .B(new_n6859), .Y(new_n6861));
  xor_4  g06485(.A(new_n6861), .B(new_n6858), .Y(new_n6862));
  nand_5 g06486(.A(new_n6839), .B(new_n6838), .Y(new_n6863));
  nand_5 g06487(.A(new_n6840), .B(new_n6837), .Y(new_n6864));
  nand_5 g06488(.A(new_n6864), .B(new_n6863), .Y(new_n6865));
  nand_5 g06489(.A(pi224), .B(pi148), .Y(new_n6866));
  xor_4  g06490(.A(new_n6866), .B(new_n6865), .Y(new_n6867));
  xor_4  g06491(.A(new_n6867), .B(new_n6862), .Y(new_n6868));
  not_8  g06492(.A(new_n6868), .Y(new_n6869));
  xor_4  g06493(.A(new_n6869), .B(new_n6857), .Y(new_n6870));
  xnor_4 g06494(.A(new_n6870), .B(new_n6852), .Y(new_n6871));
  xor_4  g06495(.A(new_n6871), .B(new_n6850), .Y(new_n6872));
  nand_5 g06496(.A(new_n6833), .B(new_n6821), .Y(new_n6873));
  nand_5 g06497(.A(pi252), .B(pi049), .Y(new_n6874));
  nand_5 g06498(.A(pi245), .B(pi140), .Y(new_n6875));
  nand_5 g06499(.A(pi242), .B(pi201), .Y(new_n6876));
  xor_4  g06500(.A(new_n6876), .B(new_n6875), .Y(new_n6877));
  xor_4  g06501(.A(new_n6877), .B(new_n6874), .Y(new_n6878));
  nand_5 g06502(.A(new_n6829), .B(new_n6828), .Y(new_n6879));
  nand_5 g06503(.A(new_n6830), .B(new_n6827), .Y(new_n6880));
  nand_5 g06504(.A(new_n6880), .B(new_n6879), .Y(new_n6881));
  nand_5 g06505(.A(pi171), .B(pi121), .Y(new_n6882));
  xor_4  g06506(.A(new_n6882), .B(new_n6881), .Y(new_n6883));
  xor_4  g06507(.A(new_n6883), .B(new_n6878), .Y(new_n6884));
  nand_5 g06508(.A(pi231), .B(pi107), .Y(new_n6885));
  or_6   g06509(.A(new_n6825), .B(new_n6822), .Y(new_n6886));
  nand_5 g06510(.A(new_n6832), .B(new_n6826), .Y(new_n6887));
  and_6  g06511(.A(new_n6887), .B(new_n6886), .Y(new_n6888));
  xnor_4 g06512(.A(new_n6888), .B(new_n6885), .Y(new_n6889));
  xor_4  g06513(.A(new_n6889), .B(new_n6884), .Y(new_n6890));
  xor_4  g06514(.A(new_n6890), .B(new_n6873), .Y(new_n6891));
  xnor_4 g06515(.A(new_n6891), .B(new_n6872), .Y(new_n6892));
  nand_5 g06516(.A(new_n6661), .B(new_n6665), .Y(new_n6893));
  nand_5 g06517(.A(new_n6893), .B(new_n6666), .Y(new_n6894));
  nand_5 g06518(.A(pi176), .B(pi175), .Y(new_n6895));
  or_6   g06519(.A(new_n6895), .B(new_n6894), .Y(new_n6896));
  xor_4  g06520(.A(new_n6895), .B(new_n6894), .Y(new_n6897));
  nand_5 g06521(.A(pi249), .B(pi149), .Y(new_n6898));
  nand_5 g06522(.A(pi240), .B(pi222), .Y(new_n6899));
  nand_5 g06523(.A(pi134), .B(pi125), .Y(new_n6900));
  xor_4  g06524(.A(new_n6900), .B(new_n6899), .Y(new_n6901));
  xor_4  g06525(.A(new_n6901), .B(new_n6898), .Y(new_n6902));
  not_8  g06526(.A(new_n6902), .Y(new_n6903));
  nand_5 g06527(.A(new_n6903), .B(new_n6897), .Y(new_n6904));
  nand_5 g06528(.A(new_n6904), .B(new_n6896), .Y(new_n6905));
  nand_5 g06529(.A(pi175), .B(pi040), .Y(new_n6906));
  nand_5 g06530(.A(pi249), .B(pi167), .Y(new_n6907));
  nand_5 g06531(.A(pi240), .B(pi125), .Y(new_n6908));
  nand_5 g06532(.A(pi222), .B(pi149), .Y(new_n6909));
  xor_4  g06533(.A(new_n6909), .B(new_n6908), .Y(new_n6910));
  xor_4  g06534(.A(new_n6910), .B(new_n6907), .Y(new_n6911));
  nand_5 g06535(.A(new_n6900), .B(new_n6899), .Y(new_n6912));
  nand_5 g06536(.A(new_n6901), .B(new_n6898), .Y(new_n6913));
  nand_5 g06537(.A(new_n6913), .B(new_n6912), .Y(new_n6914));
  nand_5 g06538(.A(pi176), .B(pi134), .Y(new_n6915));
  xor_4  g06539(.A(new_n6915), .B(new_n6914), .Y(new_n6916));
  xor_4  g06540(.A(new_n6916), .B(new_n6911), .Y(new_n6917));
  xor_4  g06541(.A(new_n6917), .B(new_n6906), .Y(new_n6918));
  xor_4  g06542(.A(new_n6918), .B(new_n6905), .Y(new_n6919));
  xor_4  g06543(.A(new_n6903), .B(new_n6897), .Y(new_n6920));
  nor_5  g06544(.A(new_n6668), .B(new_n6661), .Y(new_n6921));
  and_6  g06545(.A(new_n6921), .B(new_n6920), .Y(new_n6922));
  xor_4  g06546(.A(new_n6922), .B(new_n6919), .Y(new_n6923));
  nor_5  g06547(.A(new_n6923), .B(new_n6892), .Y(new_n6924));
  xor_4  g06548(.A(new_n6923), .B(new_n6892), .Y(new_n6925));
  xor_4  g06549(.A(new_n6921), .B(new_n6920), .Y(new_n6926));
  not_8  g06550(.A(new_n6926), .Y(new_n6927));
  nand_5 g06551(.A(new_n6670), .B(new_n6660), .Y(new_n6928));
  nand_5 g06552(.A(new_n6690), .B(new_n6671), .Y(new_n6929));
  nand_5 g06553(.A(new_n6929), .B(new_n6928), .Y(new_n6930));
  nor_5  g06554(.A(new_n6930), .B(new_n6927), .Y(new_n6931));
  xor_4  g06555(.A(new_n6930), .B(new_n6926), .Y(new_n6932));
  xor_4  g06556(.A(new_n6848), .B(new_n6836), .Y(new_n6933));
  nor_5  g06557(.A(new_n6933), .B(new_n6932), .Y(new_n6934));
  nor_5  g06558(.A(new_n6934), .B(new_n6931), .Y(new_n6935));
  and_6  g06559(.A(new_n6935), .B(new_n6925), .Y(new_n6936));
  nor_5  g06560(.A(new_n6936), .B(new_n6924), .Y(new_n6937));
  nand_5 g06561(.A(new_n6922), .B(new_n6919), .Y(new_n6938));
  nand_5 g06562(.A(pi175), .B(pi174), .Y(new_n6939));
  xor_4  g06563(.A(new_n6939), .B(new_n6938), .Y(new_n6940));
  nor_5  g06564(.A(new_n6917), .B(new_n6906), .Y(new_n6941));
  nand_5 g06565(.A(new_n6918), .B(new_n6905), .Y(new_n6942));
  not_8  g06566(.A(new_n6942), .Y(new_n6943));
  nor_5  g06567(.A(new_n6943), .B(new_n6941), .Y(new_n6944));
  not_8  g06568(.A(new_n6944), .Y(new_n6945));
  nand_5 g06569(.A(new_n6909), .B(new_n6908), .Y(new_n6946));
  nand_5 g06570(.A(new_n6910), .B(new_n6907), .Y(new_n6947));
  nand_5 g06571(.A(new_n6947), .B(new_n6946), .Y(new_n6948));
  nand_5 g06572(.A(pi149), .B(pi125), .Y(new_n6949));
  nand_5 g06573(.A(pi222), .B(pi167), .Y(new_n6950));
  nand_5 g06574(.A(pi249), .B(pi181), .Y(new_n6951));
  nand_5 g06575(.A(new_n6951), .B(new_n6950), .Y(new_n6952));
  nand_5 g06576(.A(pi222), .B(pi181), .Y(new_n6953));
  nor_5  g06577(.A(new_n6953), .B(new_n6907), .Y(new_n6954));
  not_8  g06578(.A(new_n6954), .Y(new_n6955));
  nand_5 g06579(.A(new_n6955), .B(new_n6952), .Y(new_n6956));
  xor_4  g06580(.A(new_n6956), .B(new_n6949), .Y(new_n6957));
  xor_4  g06581(.A(new_n6957), .B(new_n6948), .Y(new_n6958));
  nand_5 g06582(.A(new_n6915), .B(new_n6914), .Y(new_n6959));
  nand_5 g06583(.A(new_n6916), .B(new_n6911), .Y(new_n6960));
  nand_5 g06584(.A(new_n6960), .B(new_n6959), .Y(new_n6961));
  nand_5 g06585(.A(pi240), .B(pi176), .Y(new_n6962));
  nand_5 g06586(.A(pi134), .B(pi040), .Y(new_n6963));
  nand_5 g06587(.A(new_n6963), .B(new_n6962), .Y(new_n6964));
  nand_5 g06588(.A(pi240), .B(pi040), .Y(new_n6965));
  nor_5  g06589(.A(new_n6965), .B(new_n6915), .Y(new_n6966));
  not_8  g06590(.A(new_n6966), .Y(new_n6967));
  nand_5 g06591(.A(new_n6967), .B(new_n6964), .Y(new_n6968));
  xor_4  g06592(.A(new_n6968), .B(new_n6961), .Y(new_n6969));
  xnor_4 g06593(.A(new_n6969), .B(new_n6958), .Y(new_n6970));
  xor_4  g06594(.A(new_n6970), .B(new_n6945), .Y(new_n6971));
  xor_4  g06595(.A(new_n6971), .B(new_n6940), .Y(new_n6972));
  nand_5 g06596(.A(new_n6871), .B(new_n6850), .Y(new_n6973));
  nand_5 g06597(.A(new_n6891), .B(new_n6872), .Y(new_n6974));
  nand_5 g06598(.A(new_n6974), .B(new_n6973), .Y(new_n6975));
  not_8  g06599(.A(new_n6873), .Y(new_n6976));
  nand_5 g06600(.A(new_n6890), .B(new_n6976), .Y(new_n6977));
  nand_5 g06601(.A(pi107), .B(pi005), .Y(new_n6978));
  nand_5 g06602(.A(new_n6882), .B(new_n6881), .Y(new_n6979));
  nand_5 g06603(.A(new_n6883), .B(new_n6878), .Y(new_n6980));
  nand_5 g06604(.A(new_n6980), .B(new_n6979), .Y(new_n6981));
  nand_5 g06605(.A(pi231), .B(pi171), .Y(new_n6982));
  nand_5 g06606(.A(pi121), .B(pi049), .Y(new_n6983));
  and_6  g06607(.A(new_n6983), .B(new_n6982), .Y(new_n6984));
  nand_5 g06608(.A(pi231), .B(pi049), .Y(new_n6985));
  nor_5  g06609(.A(new_n6985), .B(new_n6882), .Y(new_n6986));
  or_6   g06610(.A(new_n6986), .B(new_n6984), .Y(new_n6987));
  nand_5 g06611(.A(pi201), .B(pi140), .Y(new_n6988));
  nand_5 g06612(.A(pi242), .B(pi156), .Y(new_n6989));
  nand_5 g06613(.A(new_n6989), .B(new_n6988), .Y(new_n6990));
  nand_5 g06614(.A(pi156), .B(pi140), .Y(new_n6991));
  nor_5  g06615(.A(new_n6991), .B(new_n6876), .Y(new_n6992));
  not_8  g06616(.A(new_n6992), .Y(new_n6993));
  nand_5 g06617(.A(new_n6993), .B(new_n6990), .Y(new_n6994));
  nand_5 g06618(.A(pi252), .B(pi245), .Y(new_n6995));
  nand_5 g06619(.A(new_n6876), .B(new_n6875), .Y(new_n6996));
  nand_5 g06620(.A(new_n6877), .B(new_n6874), .Y(new_n6997));
  nand_5 g06621(.A(new_n6997), .B(new_n6996), .Y(new_n6998));
  xor_4  g06622(.A(new_n6998), .B(new_n6995), .Y(new_n6999));
  xor_4  g06623(.A(new_n6999), .B(new_n6994), .Y(new_n7000));
  xor_4  g06624(.A(new_n7000), .B(new_n6987), .Y(new_n7001));
  not_8  g06625(.A(new_n7001), .Y(new_n7002));
  xor_4  g06626(.A(new_n7002), .B(new_n6981), .Y(new_n7003));
  nor_5  g06627(.A(new_n6888), .B(new_n6885), .Y(new_n7004));
  nor_5  g06628(.A(new_n6889), .B(new_n6884), .Y(new_n7005));
  nor_5  g06629(.A(new_n7005), .B(new_n7004), .Y(new_n7006));
  xor_4  g06630(.A(new_n7006), .B(new_n7003), .Y(new_n7007));
  xor_4  g06631(.A(new_n7007), .B(new_n6978), .Y(new_n7008));
  xor_4  g06632(.A(new_n7008), .B(new_n6977), .Y(new_n7009));
  nand_5 g06633(.A(new_n6870), .B(new_n6852), .Y(new_n7010));
  nand_5 g06634(.A(pi163), .B(pi127), .Y(new_n7011));
  nor_5  g06635(.A(new_n6856), .B(new_n6853), .Y(new_n7012));
  and_6  g06636(.A(new_n6869), .B(new_n6857), .Y(new_n7013));
  nor_5  g06637(.A(new_n7013), .B(new_n7012), .Y(new_n7014));
  nand_5 g06638(.A(new_n6866), .B(new_n6865), .Y(new_n7015));
  nand_5 g06639(.A(new_n6867), .B(new_n6862), .Y(new_n7016));
  nand_5 g06640(.A(new_n7016), .B(new_n7015), .Y(new_n7017));
  nand_5 g06641(.A(pi228), .B(pi224), .Y(new_n7018));
  nand_5 g06642(.A(pi255), .B(pi148), .Y(new_n7019));
  and_6  g06643(.A(new_n7019), .B(new_n7018), .Y(new_n7020));
  nand_5 g06644(.A(pi255), .B(pi228), .Y(new_n7021));
  nor_5  g06645(.A(new_n7021), .B(new_n6866), .Y(new_n7022));
  or_6   g06646(.A(new_n7022), .B(new_n7020), .Y(new_n7023));
  nand_5 g06647(.A(new_n6860), .B(new_n6859), .Y(new_n7024));
  nand_5 g06648(.A(new_n6861), .B(new_n6858), .Y(new_n7025));
  nand_5 g06649(.A(new_n7025), .B(new_n7024), .Y(new_n7026));
  nand_5 g06650(.A(pi039), .B(pi024), .Y(new_n7027));
  nand_5 g06651(.A(pi116), .B(pi111), .Y(new_n7028));
  nand_5 g06652(.A(pi210), .B(pi070), .Y(new_n7029));
  nand_5 g06653(.A(new_n7029), .B(new_n7028), .Y(new_n7030));
  nand_5 g06654(.A(pi111), .B(pi070), .Y(new_n7031));
  nor_5  g06655(.A(new_n7031), .B(new_n6858), .Y(new_n7032));
  not_8  g06656(.A(new_n7032), .Y(new_n7033));
  nand_5 g06657(.A(new_n7033), .B(new_n7030), .Y(new_n7034));
  xor_4  g06658(.A(new_n7034), .B(new_n7027), .Y(new_n7035));
  xor_4  g06659(.A(new_n7035), .B(new_n7026), .Y(new_n7036));
  xor_4  g06660(.A(new_n7036), .B(new_n7023), .Y(new_n7037));
  not_8  g06661(.A(new_n7037), .Y(new_n7038));
  xor_4  g06662(.A(new_n7038), .B(new_n7017), .Y(new_n7039));
  xor_4  g06663(.A(new_n7039), .B(new_n7014), .Y(new_n7040));
  xor_4  g06664(.A(new_n7040), .B(new_n7011), .Y(new_n7041));
  xor_4  g06665(.A(new_n7041), .B(new_n7010), .Y(new_n7042));
  nand_5 g06666(.A(new_n7042), .B(new_n7009), .Y(new_n7043));
  or_6   g06667(.A(new_n7042), .B(new_n7009), .Y(new_n7044));
  nand_5 g06668(.A(new_n7044), .B(new_n7043), .Y(new_n7045));
  xor_4  g06669(.A(new_n7045), .B(new_n6975), .Y(new_n7046));
  and_6  g06670(.A(new_n7046), .B(new_n6972), .Y(new_n7047));
  nor_5  g06671(.A(new_n7046), .B(new_n6972), .Y(new_n7048));
  nor_5  g06672(.A(new_n7048), .B(new_n7047), .Y(new_n7049));
  xor_4  g06673(.A(new_n7049), .B(new_n6937), .Y(new_n7050));
  nand_5 g06674(.A(new_n7050), .B(new_n6817), .Y(new_n7051));
  xor_4  g06675(.A(new_n6751), .B(new_n6747), .Y(new_n7052));
  not_8  g06676(.A(new_n7052), .Y(new_n7053));
  nand_5 g06677(.A(new_n6715), .B(new_n6706), .Y(new_n7054));
  nand_5 g06678(.A(new_n6716), .B(new_n6691), .Y(new_n7055));
  nand_5 g06679(.A(new_n7055), .B(new_n7054), .Y(new_n7056));
  xor_4  g06680(.A(new_n6749), .B(new_n6748), .Y(new_n7057));
  not_8  g06681(.A(new_n7057), .Y(new_n7058));
  nand_5 g06682(.A(new_n7058), .B(new_n7056), .Y(new_n7059));
  xor_4  g06683(.A(new_n7058), .B(new_n7056), .Y(new_n7060));
  xor_4  g06684(.A(new_n6933), .B(new_n6932), .Y(new_n7061));
  not_8  g06685(.A(new_n7061), .Y(new_n7062));
  nand_5 g06686(.A(new_n7062), .B(new_n7060), .Y(new_n7063));
  nand_5 g06687(.A(new_n7063), .B(new_n7059), .Y(new_n7064));
  nor_5  g06688(.A(new_n7064), .B(new_n7053), .Y(new_n7065));
  xor_4  g06689(.A(new_n6935), .B(new_n6925), .Y(new_n7066));
  xor_4  g06690(.A(new_n7064), .B(new_n7053), .Y(new_n7067));
  not_8  g06691(.A(new_n7067), .Y(new_n7068));
  nor_5  g06692(.A(new_n7068), .B(new_n7066), .Y(new_n7069));
  nor_5  g06693(.A(new_n7069), .B(new_n7065), .Y(new_n7070));
  xnor_4 g06694(.A(new_n7050), .B(new_n6817), .Y(new_n7071));
  or_6   g06695(.A(new_n7071), .B(new_n7070), .Y(new_n7072));
  nand_5 g06696(.A(new_n7072), .B(new_n7051), .Y(new_n7073));
  or_6   g06697(.A(new_n7073), .B(new_n6816), .Y(new_n7074));
  xor_4  g06698(.A(new_n7073), .B(new_n6816), .Y(new_n7075));
  nand_5 g06699(.A(new_n6939), .B(new_n6938), .Y(new_n7076));
  not_8  g06700(.A(new_n6971), .Y(new_n7077));
  nand_5 g06701(.A(new_n7077), .B(new_n6940), .Y(new_n7078));
  nand_5 g06702(.A(new_n7078), .B(new_n7076), .Y(new_n7079));
  nand_5 g06703(.A(new_n6970), .B(new_n6945), .Y(new_n7080));
  nand_5 g06704(.A(new_n6968), .B(new_n6961), .Y(new_n7081));
  nand_5 g06705(.A(new_n6969), .B(new_n6958), .Y(new_n7082));
  nand_5 g06706(.A(new_n7082), .B(new_n7081), .Y(new_n7083));
  xor_4  g06707(.A(new_n7083), .B(new_n6967), .Y(new_n7084));
  nand_5 g06708(.A(pi249), .B(pi200), .Y(new_n7085));
  nand_5 g06709(.A(pi167), .B(pi125), .Y(new_n7086));
  xor_4  g06710(.A(new_n7086), .B(new_n7085), .Y(new_n7087));
  xor_4  g06711(.A(new_n7087), .B(new_n6953), .Y(new_n7088));
  nand_5 g06712(.A(pi176), .B(pi149), .Y(new_n7089));
  xor_4  g06713(.A(new_n7089), .B(new_n6954), .Y(new_n7090));
  xor_4  g06714(.A(new_n7090), .B(new_n7088), .Y(new_n7091));
  nand_5 g06715(.A(new_n6956), .B(new_n6949), .Y(new_n7092));
  nand_5 g06716(.A(new_n6957), .B(new_n6948), .Y(new_n7093));
  nand_5 g06717(.A(new_n7093), .B(new_n7092), .Y(new_n7094));
  nand_5 g06718(.A(pi175), .B(pi157), .Y(new_n7095));
  nand_5 g06719(.A(pi174), .B(pi134), .Y(new_n7096));
  xor_4  g06720(.A(new_n7096), .B(new_n7095), .Y(new_n7097));
  xor_4  g06721(.A(new_n7097), .B(new_n6965), .Y(new_n7098));
  xnor_4 g06722(.A(new_n7098), .B(new_n7094), .Y(new_n7099));
  xor_4  g06723(.A(new_n7099), .B(new_n7091), .Y(new_n7100));
  xor_4  g06724(.A(new_n7100), .B(new_n7084), .Y(new_n7101));
  xnor_4 g06725(.A(new_n7101), .B(new_n7080), .Y(new_n7102));
  xnor_4 g06726(.A(new_n7102), .B(new_n7079), .Y(new_n7103));
  nand_5 g06727(.A(new_n7044), .B(new_n6975), .Y(new_n7104));
  nand_5 g06728(.A(new_n7104), .B(new_n7043), .Y(new_n7105));
  nor_5  g06729(.A(new_n7040), .B(new_n7011), .Y(new_n7106));
  not_8  g06730(.A(new_n7010), .Y(new_n7107));
  and_6  g06731(.A(new_n7041), .B(new_n7107), .Y(new_n7108));
  nor_5  g06732(.A(new_n7108), .B(new_n7106), .Y(new_n7109));
  not_8  g06733(.A(new_n7039), .Y(new_n7110));
  nor_5  g06734(.A(new_n7110), .B(new_n7014), .Y(new_n7111));
  nand_5 g06735(.A(new_n7034), .B(new_n7027), .Y(new_n7112));
  nand_5 g06736(.A(new_n7035), .B(new_n7026), .Y(new_n7113));
  nand_5 g06737(.A(new_n7113), .B(new_n7112), .Y(new_n7114));
  nand_5 g06738(.A(pi232), .B(pi163), .Y(new_n7115));
  nand_5 g06739(.A(pi148), .B(pi127), .Y(new_n7116));
  xor_4  g06740(.A(new_n7116), .B(new_n7115), .Y(new_n7117));
  xor_4  g06741(.A(new_n7117), .B(new_n7021), .Y(new_n7118));
  xnor_4 g06742(.A(new_n7118), .B(new_n7114), .Y(new_n7119));
  nand_5 g06743(.A(pi224), .B(pi039), .Y(new_n7120));
  xor_4  g06744(.A(new_n7120), .B(new_n7033), .Y(new_n7121));
  nand_5 g06745(.A(pi210), .B(pi115), .Y(new_n7122));
  nand_5 g06746(.A(pi116), .B(pi024), .Y(new_n7123));
  xor_4  g06747(.A(new_n7123), .B(new_n7122), .Y(new_n7124));
  xnor_4 g06748(.A(new_n7124), .B(new_n7031), .Y(new_n7125));
  xnor_4 g06749(.A(new_n7125), .B(new_n7121), .Y(new_n7126));
  xor_4  g06750(.A(new_n7126), .B(new_n7119), .Y(new_n7127));
  nor_5  g06751(.A(new_n7038), .B(new_n7017), .Y(new_n7128));
  nand_5 g06752(.A(new_n7128), .B(new_n7022), .Y(new_n7129));
  or_6   g06753(.A(new_n7038), .B(new_n7017), .Y(new_n7130));
  nor_5  g06754(.A(new_n7036), .B(new_n7023), .Y(new_n7131));
  nor_5  g06755(.A(new_n7131), .B(new_n7022), .Y(new_n7132));
  nand_5 g06756(.A(new_n7132), .B(new_n7130), .Y(new_n7133));
  nand_5 g06757(.A(new_n7133), .B(new_n7129), .Y(new_n7134));
  xor_4  g06758(.A(new_n7134), .B(new_n7127), .Y(new_n7135));
  xor_4  g06759(.A(new_n7135), .B(new_n7111), .Y(new_n7136));
  xor_4  g06760(.A(new_n7136), .B(new_n7109), .Y(new_n7137));
  nor_5  g06761(.A(new_n7007), .B(new_n6978), .Y(new_n7138));
  not_8  g06762(.A(new_n6977), .Y(new_n7139));
  and_6  g06763(.A(new_n7008), .B(new_n7139), .Y(new_n7140));
  nor_5  g06764(.A(new_n7140), .B(new_n7138), .Y(new_n7141));
  not_8  g06765(.A(new_n7003), .Y(new_n7142));
  nor_5  g06766(.A(new_n7006), .B(new_n7142), .Y(new_n7143));
  nor_5  g06767(.A(new_n7002), .B(new_n6981), .Y(new_n7144));
  nand_5 g06768(.A(new_n7144), .B(new_n6986), .Y(new_n7145));
  or_6   g06769(.A(new_n7002), .B(new_n6981), .Y(new_n7146));
  nor_5  g06770(.A(new_n7000), .B(new_n6987), .Y(new_n7147));
  nor_5  g06771(.A(new_n7147), .B(new_n6986), .Y(new_n7148));
  nand_5 g06772(.A(new_n7148), .B(new_n7146), .Y(new_n7149));
  nand_5 g06773(.A(new_n7149), .B(new_n7145), .Y(new_n7150));
  nand_5 g06774(.A(pi242), .B(pi063), .Y(new_n7151));
  nand_5 g06775(.A(pi252), .B(pi201), .Y(new_n7152));
  xor_4  g06776(.A(new_n7152), .B(new_n7151), .Y(new_n7153));
  xor_4  g06777(.A(new_n7153), .B(new_n6991), .Y(new_n7154));
  nand_5 g06778(.A(pi245), .B(pi121), .Y(new_n7155));
  xor_4  g06779(.A(new_n7155), .B(new_n6992), .Y(new_n7156));
  xor_4  g06780(.A(new_n7156), .B(new_n7154), .Y(new_n7157));
  nand_5 g06781(.A(new_n6998), .B(new_n6995), .Y(new_n7158));
  nand_5 g06782(.A(new_n6999), .B(new_n6994), .Y(new_n7159));
  nand_5 g06783(.A(new_n7159), .B(new_n7158), .Y(new_n7160));
  nand_5 g06784(.A(pi107), .B(pi021), .Y(new_n7161));
  nand_5 g06785(.A(pi171), .B(pi005), .Y(new_n7162));
  xor_4  g06786(.A(new_n7162), .B(new_n7161), .Y(new_n7163));
  xor_4  g06787(.A(new_n7163), .B(new_n6985), .Y(new_n7164));
  xnor_4 g06788(.A(new_n7164), .B(new_n7160), .Y(new_n7165));
  xor_4  g06789(.A(new_n7165), .B(new_n7157), .Y(new_n7166));
  not_8  g06790(.A(new_n7166), .Y(new_n7167));
  xor_4  g06791(.A(new_n7167), .B(new_n7150), .Y(new_n7168));
  xor_4  g06792(.A(new_n7168), .B(new_n7143), .Y(new_n7169));
  xor_4  g06793(.A(new_n7169), .B(new_n7141), .Y(new_n7170));
  xor_4  g06794(.A(new_n7170), .B(new_n7137), .Y(new_n7171));
  xor_4  g06795(.A(new_n7171), .B(new_n7105), .Y(new_n7172));
  xor_4  g06796(.A(new_n7172), .B(new_n7103), .Y(new_n7173));
  nor_5  g06797(.A(new_n7047), .B(new_n6937), .Y(new_n7174));
  nor_5  g06798(.A(new_n7174), .B(new_n7048), .Y(new_n7175));
  xnor_4 g06799(.A(new_n7175), .B(new_n7173), .Y(new_n7176));
  nand_5 g06800(.A(new_n7176), .B(new_n7075), .Y(new_n7177));
  nand_5 g06801(.A(new_n7177), .B(new_n7074), .Y(new_n7178));
  nand_5 g06802(.A(pi224), .B(pi116), .Y(new_n7179));
  nand_5 g06803(.A(new_n7123), .B(new_n7122), .Y(new_n7180));
  nand_5 g06804(.A(new_n7124), .B(new_n7031), .Y(new_n7181));
  nand_5 g06805(.A(new_n7181), .B(new_n7180), .Y(new_n7182));
  xor_4  g06806(.A(new_n7182), .B(new_n7179), .Y(new_n7183));
  xor_4  g06807(.A(new_n7183), .B(new_n7178), .Y(new_n7184));
  or_6   g06808(.A(new_n6813), .B(new_n6796), .Y(new_n7185));
  nand_5 g06809(.A(new_n7185), .B(new_n6795), .Y(new_n7186));
  or_6   g06810(.A(new_n7167), .B(new_n7150), .Y(new_n7187));
  nand_5 g06811(.A(new_n7187), .B(new_n7149), .Y(new_n7188));
  xor_4  g06812(.A(new_n7188), .B(new_n7186), .Y(new_n7189));
  nor_5  g06813(.A(new_n7164), .B(new_n7160), .Y(new_n7190));
  not_8  g06814(.A(new_n7157), .Y(new_n7191));
  nor_5  g06815(.A(new_n7165), .B(new_n7191), .Y(new_n7192));
  nor_5  g06816(.A(new_n7192), .B(new_n7190), .Y(new_n7193));
  nand_5 g06817(.A(new_n7162), .B(new_n7161), .Y(new_n7194));
  nand_5 g06818(.A(new_n7163), .B(new_n6985), .Y(new_n7195));
  nand_5 g06819(.A(new_n7195), .B(new_n7194), .Y(new_n7196));
  xor_4  g06820(.A(new_n7196), .B(new_n7193), .Y(new_n7197));
  nand_5 g06821(.A(pi181), .B(pi125), .Y(new_n7198));
  nand_5 g06822(.A(new_n7083), .B(new_n6967), .Y(new_n7199));
  nand_5 g06823(.A(new_n7100), .B(new_n7084), .Y(new_n7200));
  nand_5 g06824(.A(new_n7200), .B(new_n7199), .Y(new_n7201));
  nand_5 g06825(.A(pi247), .B(pi081), .Y(new_n7202));
  xnor_4 g06826(.A(new_n7202), .B(new_n7201), .Y(new_n7203));
  xor_4  g06827(.A(new_n7203), .B(new_n7198), .Y(new_n7204));
  nand_5 g06828(.A(pi115), .B(pi111), .Y(new_n7205));
  nand_5 g06829(.A(pi191), .B(pi163), .Y(new_n7206));
  nand_5 g06830(.A(pi106), .B(pi080), .Y(new_n7207));
  nand_5 g06831(.A(new_n6808), .B(new_n6807), .Y(new_n7208));
  nand_5 g06832(.A(new_n6809), .B(new_n6774), .Y(new_n7209));
  nand_5 g06833(.A(new_n7209), .B(new_n7208), .Y(new_n7210));
  xnor_4 g06834(.A(new_n7210), .B(new_n7207), .Y(new_n7211));
  xor_4  g06835(.A(new_n7211), .B(new_n7206), .Y(new_n7212));
  xor_4  g06836(.A(new_n7212), .B(new_n7205), .Y(new_n7213));
  or_6   g06837(.A(new_n7134), .B(new_n7127), .Y(new_n7214));
  nand_5 g06838(.A(new_n7214), .B(new_n7133), .Y(new_n7215));
  nand_5 g06839(.A(new_n7096), .B(new_n7095), .Y(new_n7216));
  nand_5 g06840(.A(new_n7097), .B(new_n6965), .Y(new_n7217));
  nand_5 g06841(.A(new_n7217), .B(new_n7216), .Y(new_n7218));
  nand_5 g06842(.A(pi070), .B(pi024), .Y(new_n7219));
  xnor_4 g06843(.A(new_n7219), .B(new_n7218), .Y(new_n7220));
  xor_4  g06844(.A(new_n7220), .B(new_n7215), .Y(new_n7221));
  xor_4  g06845(.A(new_n7221), .B(new_n7213), .Y(new_n7222));
  xor_4  g06846(.A(new_n7222), .B(new_n7204), .Y(new_n7223));
  xor_4  g06847(.A(new_n7223), .B(new_n7197), .Y(new_n7224));
  nor_5  g06848(.A(new_n7101), .B(new_n7080), .Y(new_n7225));
  nor_5  g06849(.A(new_n7102), .B(new_n7079), .Y(new_n7226));
  nor_5  g06850(.A(new_n7226), .B(new_n7225), .Y(new_n7227));
  nand_5 g06851(.A(pi175), .B(pi017), .Y(new_n7228));
  nand_5 g06852(.A(pi249), .B(pi203), .Y(new_n7229));
  nand_5 g06853(.A(new_n6803), .B(new_n6799), .Y(new_n7230));
  nand_5 g06854(.A(new_n6811), .B(new_n6804), .Y(new_n7231));
  nand_5 g06855(.A(new_n7231), .B(new_n7230), .Y(new_n7232));
  xor_4  g06856(.A(new_n7232), .B(new_n7229), .Y(new_n7233));
  xor_4  g06857(.A(new_n7233), .B(new_n7228), .Y(new_n7234));
  xor_4  g06858(.A(new_n7234), .B(new_n7227), .Y(new_n7235));
  xor_4  g06859(.A(new_n7235), .B(new_n7224), .Y(new_n7236));
  nand_5 g06860(.A(pi171), .B(pi021), .Y(new_n7237));
  nand_5 g06861(.A(pi232), .B(pi148), .Y(new_n7238));
  nand_5 g06862(.A(pi245), .B(pi231), .Y(new_n7239));
  xor_4  g06863(.A(new_n7239), .B(new_n7238), .Y(new_n7240));
  xor_4  g06864(.A(new_n7240), .B(new_n7237), .Y(new_n7241));
  xor_4  g06865(.A(new_n7241), .B(new_n7236), .Y(new_n7242));
  xor_4  g06866(.A(new_n7242), .B(new_n7189), .Y(new_n7243));
  nor_5  g06867(.A(new_n6805), .B(new_n6776), .Y(new_n7244));
  nor_5  g06868(.A(new_n6810), .B(new_n6806), .Y(new_n7245));
  nor_5  g06869(.A(new_n7245), .B(new_n7244), .Y(new_n7246));
  or_6   g06870(.A(new_n7172), .B(new_n7103), .Y(new_n7247));
  nand_5 g06871(.A(new_n7175), .B(new_n7173), .Y(new_n7248));
  nand_5 g06872(.A(new_n7248), .B(new_n7247), .Y(new_n7249));
  nand_5 g06873(.A(pi228), .B(pi127), .Y(new_n7250));
  xor_4  g06874(.A(new_n7250), .B(new_n7249), .Y(new_n7251));
  nand_5 g06875(.A(new_n7152), .B(new_n7151), .Y(new_n7252));
  nand_5 g06876(.A(new_n7153), .B(new_n6991), .Y(new_n7253));
  nand_5 g06877(.A(new_n7253), .B(new_n7252), .Y(new_n7254));
  nand_5 g06878(.A(new_n7116), .B(new_n7115), .Y(new_n7255));
  nand_5 g06879(.A(new_n7117), .B(new_n7021), .Y(new_n7256));
  nand_5 g06880(.A(new_n7256), .B(new_n7255), .Y(new_n7257));
  xor_4  g06881(.A(new_n7257), .B(new_n7254), .Y(new_n7258));
  nand_5 g06882(.A(pi252), .B(pi156), .Y(new_n7259));
  or_6   g06883(.A(new_n7120), .B(new_n7033), .Y(new_n7260));
  nand_5 g06884(.A(new_n7125), .B(new_n7121), .Y(new_n7261));
  nand_5 g06885(.A(new_n7261), .B(new_n7260), .Y(new_n7262));
  nand_5 g06886(.A(pi107), .B(pi082), .Y(new_n7263));
  xor_4  g06887(.A(new_n7263), .B(new_n7262), .Y(new_n7264));
  xor_4  g06888(.A(new_n7264), .B(new_n7259), .Y(new_n7265));
  nand_5 g06889(.A(pi201), .B(pi121), .Y(new_n7266));
  nand_5 g06890(.A(pi255), .B(pi039), .Y(new_n7267));
  xor_4  g06891(.A(new_n7267), .B(new_n7266), .Y(new_n7268));
  xor_4  g06892(.A(new_n7268), .B(new_n7265), .Y(new_n7269));
  xor_4  g06893(.A(new_n7269), .B(new_n7258), .Y(new_n7270));
  xor_4  g06894(.A(new_n7270), .B(new_n7251), .Y(new_n7271));
  xor_4  g06895(.A(new_n7271), .B(new_n7246), .Y(new_n7272));
  nand_5 g06896(.A(pi049), .B(pi005), .Y(new_n7273));
  nor_5  g06897(.A(new_n7155), .B(new_n6993), .Y(new_n7274));
  nor_5  g06898(.A(new_n7156), .B(new_n7154), .Y(new_n7275));
  or_6   g06899(.A(new_n7275), .B(new_n7274), .Y(new_n7276));
  xor_4  g06900(.A(new_n7276), .B(new_n7273), .Y(new_n7277));
  nand_5 g06901(.A(new_n6801), .B(new_n6800), .Y(new_n7278));
  nand_5 g06902(.A(new_n6802), .B(new_n6765), .Y(new_n7279));
  nand_5 g06903(.A(new_n7279), .B(new_n7278), .Y(new_n7280));
  not_8  g06904(.A(new_n7143), .Y(new_n7281));
  nor_5  g06905(.A(new_n7168), .B(new_n7281), .Y(new_n7282));
  nor_5  g06906(.A(new_n7169), .B(new_n7141), .Y(new_n7283));
  nor_5  g06907(.A(new_n7283), .B(new_n7282), .Y(new_n7284));
  xor_4  g06908(.A(new_n7284), .B(new_n7280), .Y(new_n7285));
  nand_5 g06909(.A(pi222), .B(pi200), .Y(new_n7286));
  nand_5 g06910(.A(pi234), .B(pi227), .Y(new_n7287));
  xor_4  g06911(.A(new_n7287), .B(new_n7286), .Y(new_n7288));
  nand_5 g06912(.A(pi157), .B(pi134), .Y(new_n7289));
  nor_5  g06913(.A(new_n7098), .B(new_n7094), .Y(new_n7290));
  not_8  g06914(.A(new_n7091), .Y(new_n7291));
  nor_5  g06915(.A(new_n7099), .B(new_n7291), .Y(new_n7292));
  nor_5  g06916(.A(new_n7292), .B(new_n7290), .Y(new_n7293));
  xor_4  g06917(.A(new_n7293), .B(new_n7289), .Y(new_n7294));
  not_8  g06918(.A(new_n6814), .Y(new_n7295));
  nand_5 g06919(.A(new_n7295), .B(new_n6787), .Y(new_n7296));
  or_6   g06920(.A(new_n6815), .B(new_n6786), .Y(new_n7297));
  nand_5 g06921(.A(new_n7297), .B(new_n7296), .Y(new_n7298));
  nand_5 g06922(.A(pi149), .B(pi040), .Y(new_n7299));
  nor_5  g06923(.A(new_n7089), .B(new_n6955), .Y(new_n7300));
  nor_5  g06924(.A(new_n7090), .B(new_n7088), .Y(new_n7301));
  nor_5  g06925(.A(new_n7301), .B(new_n7300), .Y(new_n7302));
  xor_4  g06926(.A(new_n7302), .B(new_n7299), .Y(new_n7303));
  xor_4  g06927(.A(new_n7303), .B(new_n7298), .Y(new_n7304));
  xor_4  g06928(.A(new_n7304), .B(new_n7294), .Y(new_n7305));
  xor_4  g06929(.A(new_n7305), .B(new_n7288), .Y(new_n7306));
  xor_4  g06930(.A(new_n7306), .B(new_n7285), .Y(new_n7307));
  nand_5 g06931(.A(pi214), .B(pi100), .Y(new_n7308));
  nand_5 g06932(.A(pi187), .B(pi117), .Y(new_n7309));
  xor_4  g06933(.A(new_n7309), .B(new_n7308), .Y(new_n7310));
  nand_5 g06934(.A(new_n7086), .B(new_n7085), .Y(new_n7311));
  nand_5 g06935(.A(new_n7087), .B(new_n6953), .Y(new_n7312));
  nand_5 g06936(.A(new_n7312), .B(new_n7311), .Y(new_n7313));
  nand_5 g06937(.A(pi233), .B(pi016), .Y(new_n7314));
  xor_4  g06938(.A(new_n7314), .B(new_n7313), .Y(new_n7315));
  xor_4  g06939(.A(new_n7315), .B(new_n7310), .Y(new_n7316));
  or_6   g06940(.A(new_n7170), .B(new_n7137), .Y(new_n7317));
  nand_5 g06941(.A(new_n7171), .B(new_n7105), .Y(new_n7318));
  nand_5 g06942(.A(new_n7318), .B(new_n7317), .Y(new_n7319));
  not_8  g06943(.A(new_n7111), .Y(new_n7320));
  nor_5  g06944(.A(new_n7135), .B(new_n7320), .Y(new_n7321));
  nor_5  g06945(.A(new_n7136), .B(new_n7109), .Y(new_n7322));
  nor_5  g06946(.A(new_n7322), .B(new_n7321), .Y(new_n7323));
  xor_4  g06947(.A(new_n7323), .B(new_n7319), .Y(new_n7324));
  xor_4  g06948(.A(new_n7324), .B(new_n7316), .Y(new_n7325));
  nor_5  g06949(.A(new_n7118), .B(new_n7114), .Y(new_n7326));
  nor_5  g06950(.A(new_n7126), .B(new_n7119), .Y(new_n7327));
  nor_5  g06951(.A(new_n7327), .B(new_n7326), .Y(new_n7328));
  nand_5 g06952(.A(pi129), .B(pi103), .Y(new_n7329));
  nand_5 g06953(.A(pi242), .B(pi083), .Y(new_n7330));
  nand_5 g06954(.A(pi140), .B(pi063), .Y(new_n7331));
  xor_4  g06955(.A(new_n7331), .B(new_n7330), .Y(new_n7332));
  nand_5 g06956(.A(pi176), .B(pi167), .Y(new_n7333));
  xor_4  g06957(.A(new_n7333), .B(new_n7332), .Y(new_n7334));
  xor_4  g06958(.A(new_n7334), .B(new_n7329), .Y(new_n7335));
  xor_4  g06959(.A(new_n7335), .B(new_n7328), .Y(new_n7336));
  nand_5 g06960(.A(pi217), .B(pi202), .Y(new_n7337));
  nand_5 g06961(.A(pi240), .B(pi174), .Y(new_n7338));
  nand_5 g06962(.A(pi210), .B(pi000), .Y(new_n7339));
  xor_4  g06963(.A(new_n7339), .B(new_n7338), .Y(new_n7340));
  xor_4  g06964(.A(new_n7340), .B(new_n7337), .Y(new_n7341));
  xor_4  g06965(.A(new_n7341), .B(new_n7336), .Y(new_n7342));
  xor_4  g06966(.A(new_n7342), .B(new_n7325), .Y(new_n7343));
  xor_4  g06967(.A(new_n7343), .B(new_n7307), .Y(new_n7344));
  xor_4  g06968(.A(new_n7344), .B(new_n7277), .Y(new_n7345));
  xor_4  g06969(.A(new_n7345), .B(new_n7272), .Y(new_n7346));
  xor_4  g06970(.A(new_n7346), .B(new_n7243), .Y(new_n7347));
  xor_4  g06971(.A(new_n7347), .B(new_n7184), .Y(po036));
  xor_4  g06972(.A(new_n7071), .B(new_n7070), .Y(po037));
  xnor_4 g06973(.A(new_n3285), .B(new_n3284), .Y(po038));
  nand_5 g06974(.A(pi168), .B(pi075), .Y(new_n7351));
  nand_5 g06975(.A(pi168), .B(pi019), .Y(new_n7352));
  nand_5 g06976(.A(pi147), .B(pi139), .Y(new_n7353));
  nand_5 g06977(.A(new_n7353), .B(new_n7352), .Y(new_n7354));
  nand_5 g06978(.A(pi208), .B(pi151), .Y(new_n7355));
  or_6   g06979(.A(new_n7353), .B(new_n7352), .Y(new_n7356));
  nand_5 g06980(.A(new_n7356), .B(new_n7355), .Y(new_n7357));
  nand_5 g06981(.A(new_n7357), .B(new_n7354), .Y(new_n7358));
  nand_5 g06982(.A(pi168), .B(pi097), .Y(new_n7359));
  nor_5  g06983(.A(new_n7359), .B(new_n7358), .Y(new_n7360));
  nand_5 g06984(.A(pi147), .B(pi035), .Y(new_n7361));
  nand_5 g06985(.A(pi208), .B(pi019), .Y(new_n7362));
  nand_5 g06986(.A(pi151), .B(pi139), .Y(new_n7363));
  xor_4  g06987(.A(new_n7363), .B(new_n7362), .Y(new_n7364));
  xor_4  g06988(.A(new_n7364), .B(new_n7361), .Y(new_n7365));
  not_8  g06989(.A(new_n7365), .Y(new_n7366));
  xor_4  g06990(.A(new_n7359), .B(new_n7358), .Y(new_n7367));
  nand_5 g06991(.A(new_n7367), .B(new_n7366), .Y(new_n7368));
  not_8  g06992(.A(new_n7368), .Y(new_n7369));
  or_6   g06993(.A(new_n7369), .B(new_n7360), .Y(new_n7370));
  not_8  g06994(.A(new_n7370), .Y(new_n7371));
  nor_5  g06995(.A(new_n7371), .B(new_n7351), .Y(new_n7372));
  nand_5 g06996(.A(pi139), .B(pi019), .Y(new_n7373));
  nand_5 g06997(.A(pi147), .B(pi015), .Y(new_n7374));
  nand_5 g06998(.A(pi151), .B(pi035), .Y(new_n7375));
  xor_4  g06999(.A(new_n7375), .B(new_n7374), .Y(new_n7376));
  xor_4  g07000(.A(new_n7376), .B(new_n7373), .Y(new_n7377));
  nand_5 g07001(.A(pi208), .B(pi097), .Y(new_n7378));
  nand_5 g07002(.A(new_n7363), .B(new_n7362), .Y(new_n7379));
  nand_5 g07003(.A(new_n7364), .B(new_n7361), .Y(new_n7380));
  nand_5 g07004(.A(new_n7380), .B(new_n7379), .Y(new_n7381));
  xor_4  g07005(.A(new_n7381), .B(new_n7378), .Y(new_n7382));
  xor_4  g07006(.A(new_n7382), .B(new_n7377), .Y(new_n7383));
  xor_4  g07007(.A(new_n7370), .B(new_n7351), .Y(new_n7384));
  nor_5  g07008(.A(new_n7384), .B(new_n7383), .Y(new_n7385));
  nor_5  g07009(.A(new_n7385), .B(new_n7372), .Y(new_n7386));
  nand_5 g07010(.A(new_n7381), .B(new_n7378), .Y(new_n7387));
  nand_5 g07011(.A(new_n7382), .B(new_n7377), .Y(new_n7388));
  nand_5 g07012(.A(new_n7388), .B(new_n7387), .Y(new_n7389));
  nand_5 g07013(.A(pi139), .B(pi097), .Y(new_n7390));
  nand_5 g07014(.A(pi208), .B(pi075), .Y(new_n7391));
  nand_5 g07015(.A(new_n7391), .B(new_n7390), .Y(new_n7392));
  nand_5 g07016(.A(pi139), .B(pi075), .Y(new_n7393));
  nor_5  g07017(.A(new_n7393), .B(new_n7378), .Y(new_n7394));
  not_8  g07018(.A(new_n7394), .Y(new_n7395));
  nand_5 g07019(.A(new_n7395), .B(new_n7392), .Y(new_n7396));
  nand_5 g07020(.A(pi204), .B(pi147), .Y(new_n7397));
  nand_5 g07021(.A(pi151), .B(pi015), .Y(new_n7398));
  nand_5 g07022(.A(new_n7398), .B(new_n7397), .Y(new_n7399));
  nand_5 g07023(.A(pi204), .B(pi151), .Y(new_n7400));
  nor_5  g07024(.A(new_n7400), .B(new_n7374), .Y(new_n7401));
  not_8  g07025(.A(new_n7401), .Y(new_n7402));
  nand_5 g07026(.A(new_n7402), .B(new_n7399), .Y(new_n7403));
  nand_5 g07027(.A(pi035), .B(pi019), .Y(new_n7404));
  nand_5 g07028(.A(new_n7375), .B(new_n7374), .Y(new_n7405));
  nand_5 g07029(.A(new_n7376), .B(new_n7373), .Y(new_n7406));
  nand_5 g07030(.A(new_n7406), .B(new_n7405), .Y(new_n7407));
  xor_4  g07031(.A(new_n7407), .B(new_n7404), .Y(new_n7408));
  xor_4  g07032(.A(new_n7408), .B(new_n7403), .Y(new_n7409));
  xor_4  g07033(.A(new_n7409), .B(new_n7396), .Y(new_n7410));
  xor_4  g07034(.A(new_n7410), .B(new_n7389), .Y(new_n7411));
  nor_5  g07035(.A(new_n7411), .B(new_n7386), .Y(new_n7412));
  not_8  g07036(.A(new_n7412), .Y(new_n7413));
  nand_5 g07037(.A(new_n7409), .B(new_n7396), .Y(new_n7414));
  nand_5 g07038(.A(new_n7410), .B(new_n7389), .Y(new_n7415));
  nand_5 g07039(.A(new_n7415), .B(new_n7414), .Y(new_n7416));
  xor_4  g07040(.A(new_n7416), .B(new_n7394), .Y(new_n7417));
  nand_5 g07041(.A(pi097), .B(pi035), .Y(new_n7418));
  xor_4  g07042(.A(new_n7418), .B(new_n7401), .Y(new_n7419));
  nand_5 g07043(.A(pi147), .B(pi146), .Y(new_n7420));
  nand_5 g07044(.A(pi019), .B(pi015), .Y(new_n7421));
  xor_4  g07045(.A(new_n7421), .B(new_n7420), .Y(new_n7422));
  xor_4  g07046(.A(new_n7422), .B(new_n7400), .Y(new_n7423));
  xor_4  g07047(.A(new_n7423), .B(new_n7419), .Y(new_n7424));
  nand_5 g07048(.A(new_n7407), .B(new_n7404), .Y(new_n7425));
  nand_5 g07049(.A(new_n7408), .B(new_n7403), .Y(new_n7426));
  nand_5 g07050(.A(new_n7426), .B(new_n7425), .Y(new_n7427));
  nand_5 g07051(.A(pi208), .B(pi093), .Y(new_n7428));
  and_6  g07052(.A(pi168), .B(pi166), .Y(new_n7429));
  xor_4  g07053(.A(new_n7429), .B(new_n7428), .Y(new_n7430));
  xor_4  g07054(.A(new_n7430), .B(new_n7393), .Y(new_n7431));
  xor_4  g07055(.A(new_n7431), .B(new_n7427), .Y(new_n7432));
  xor_4  g07056(.A(new_n7432), .B(new_n7424), .Y(new_n7433));
  xnor_4 g07057(.A(new_n7433), .B(new_n7417), .Y(new_n7434));
  nor_5  g07058(.A(new_n7434), .B(new_n7413), .Y(new_n7435));
  xor_4  g07059(.A(new_n7434), .B(new_n7413), .Y(new_n7436));
  not_8  g07060(.A(new_n7436), .Y(new_n7437));
  nand_5 g07061(.A(pi168), .B(pi093), .Y(new_n7438));
  not_8  g07062(.A(new_n377), .Y(new_n7439));
  nor_5  g07063(.A(new_n7355), .B(new_n7439), .Y(new_n7440));
  and_6  g07064(.A(new_n7356), .B(new_n7354), .Y(new_n7441));
  or_6   g07065(.A(new_n7441), .B(new_n7440), .Y(new_n7442));
  nor_5  g07066(.A(new_n7442), .B(new_n7355), .Y(new_n7443));
  xor_4  g07067(.A(new_n7367), .B(new_n7365), .Y(new_n7444));
  not_8  g07068(.A(new_n7444), .Y(new_n7445));
  nand_5 g07069(.A(new_n7445), .B(new_n7443), .Y(new_n7446));
  xnor_4 g07070(.A(new_n7384), .B(new_n7383), .Y(new_n7447));
  nor_5  g07071(.A(new_n7447), .B(new_n7446), .Y(new_n7448));
  not_8  g07072(.A(new_n7448), .Y(new_n7449));
  nand_5 g07073(.A(new_n7449), .B(new_n7438), .Y(new_n7450));
  xnor_4 g07074(.A(new_n7411), .B(new_n7386), .Y(new_n7451));
  xor_4  g07075(.A(new_n7448), .B(new_n7438), .Y(new_n7452));
  not_8  g07076(.A(new_n7452), .Y(new_n7453));
  nand_5 g07077(.A(new_n7453), .B(new_n7451), .Y(new_n7454));
  nand_5 g07078(.A(new_n7454), .B(new_n7450), .Y(new_n7455));
  nor_5  g07079(.A(new_n7455), .B(new_n7437), .Y(new_n7456));
  nor_5  g07080(.A(new_n7456), .B(new_n7435), .Y(new_n7457));
  nand_5 g07081(.A(pi212), .B(pi145), .Y(new_n7458));
  nand_5 g07082(.A(pi246), .B(pi104), .Y(new_n7459));
  nor_5  g07083(.A(new_n7459), .B(new_n7458), .Y(new_n7460));
  nand_5 g07084(.A(pi206), .B(pi104), .Y(new_n7461));
  nand_5 g07085(.A(pi164), .B(pi013), .Y(new_n7462));
  nand_5 g07086(.A(new_n7462), .B(new_n7461), .Y(new_n7463));
  nand_5 g07087(.A(pi212), .B(pi032), .Y(new_n7464));
  xor_4  g07088(.A(new_n7462), .B(new_n7461), .Y(new_n7465));
  nand_5 g07089(.A(new_n7465), .B(new_n7464), .Y(new_n7466));
  nand_5 g07090(.A(new_n7466), .B(new_n7463), .Y(new_n7467));
  nand_5 g07091(.A(new_n7467), .B(new_n7458), .Y(new_n7468));
  nand_5 g07092(.A(pi164), .B(pi112), .Y(new_n7469));
  nand_5 g07093(.A(pi104), .B(pi032), .Y(new_n7470));
  nand_5 g07094(.A(pi206), .B(pi013), .Y(new_n7471));
  xor_4  g07095(.A(new_n7471), .B(new_n7470), .Y(new_n7472));
  xor_4  g07096(.A(new_n7472), .B(new_n7469), .Y(new_n7473));
  xor_4  g07097(.A(new_n7467), .B(new_n7458), .Y(new_n7474));
  nand_5 g07098(.A(new_n7474), .B(new_n7473), .Y(new_n7475));
  nand_5 g07099(.A(new_n7475), .B(new_n7468), .Y(new_n7476));
  not_8  g07100(.A(new_n7460), .Y(new_n7477));
  nand_5 g07101(.A(pi145), .B(pi104), .Y(new_n7478));
  nand_5 g07102(.A(pi246), .B(pi212), .Y(new_n7479));
  nand_5 g07103(.A(new_n7479), .B(new_n7478), .Y(new_n7480));
  nand_5 g07104(.A(new_n7480), .B(new_n7477), .Y(new_n7481));
  nand_5 g07105(.A(new_n7471), .B(new_n7470), .Y(new_n7482));
  nand_5 g07106(.A(new_n7472), .B(new_n7469), .Y(new_n7483));
  nand_5 g07107(.A(new_n7483), .B(new_n7482), .Y(new_n7484));
  nand_5 g07108(.A(pi032), .B(pi013), .Y(new_n7485));
  nand_5 g07109(.A(pi206), .B(pi112), .Y(new_n7486));
  nand_5 g07110(.A(pi164), .B(pi105), .Y(new_n7487));
  nand_5 g07111(.A(new_n7487), .B(new_n7486), .Y(new_n7488));
  nand_5 g07112(.A(pi206), .B(pi105), .Y(new_n7489));
  nor_5  g07113(.A(new_n7489), .B(new_n7469), .Y(new_n7490));
  not_8  g07114(.A(new_n7490), .Y(new_n7491));
  nand_5 g07115(.A(new_n7491), .B(new_n7488), .Y(new_n7492));
  xor_4  g07116(.A(new_n7492), .B(new_n7485), .Y(new_n7493));
  xor_4  g07117(.A(new_n7493), .B(new_n7484), .Y(new_n7494));
  xnor_4 g07118(.A(new_n7494), .B(new_n7481), .Y(new_n7495));
  nor_5  g07119(.A(new_n7495), .B(new_n7476), .Y(new_n7496));
  nand_5 g07120(.A(new_n7496), .B(new_n7460), .Y(new_n7497));
  nand_5 g07121(.A(pi145), .B(pi013), .Y(new_n7498));
  xor_4  g07122(.A(new_n7498), .B(new_n7491), .Y(new_n7499));
  nand_5 g07123(.A(pi183), .B(pi164), .Y(new_n7500));
  nand_5 g07124(.A(pi112), .B(pi032), .Y(new_n7501));
  xor_4  g07125(.A(new_n7501), .B(new_n7500), .Y(new_n7502));
  xor_4  g07126(.A(new_n7502), .B(new_n7489), .Y(new_n7503));
  not_8  g07127(.A(new_n7503), .Y(new_n7504));
  xor_4  g07128(.A(new_n7504), .B(new_n7499), .Y(new_n7505));
  nand_5 g07129(.A(new_n7492), .B(new_n7485), .Y(new_n7506));
  nand_5 g07130(.A(new_n7493), .B(new_n7484), .Y(new_n7507));
  nand_5 g07131(.A(new_n7507), .B(new_n7506), .Y(new_n7508));
  nand_5 g07132(.A(pi212), .B(pi114), .Y(new_n7509));
  nand_5 g07133(.A(pi213), .B(pi091), .Y(new_n7510));
  xor_4  g07134(.A(new_n7510), .B(new_n7509), .Y(new_n7511));
  xor_4  g07135(.A(new_n7511), .B(new_n7459), .Y(new_n7512));
  xor_4  g07136(.A(new_n7512), .B(new_n7508), .Y(new_n7513));
  xor_4  g07137(.A(new_n7513), .B(new_n7505), .Y(new_n7514));
  not_8  g07138(.A(new_n7514), .Y(new_n7515));
  nor_5  g07139(.A(new_n7494), .B(new_n7481), .Y(new_n7516));
  xor_4  g07140(.A(new_n7496), .B(new_n7477), .Y(new_n7517));
  not_8  g07141(.A(new_n7517), .Y(new_n7518));
  nor_5  g07142(.A(new_n7518), .B(new_n7516), .Y(new_n7519));
  or_6   g07143(.A(new_n7519), .B(new_n7515), .Y(new_n7520));
  nand_5 g07144(.A(new_n7520), .B(new_n7497), .Y(new_n7521));
  nand_5 g07145(.A(pi213), .B(pi031), .Y(new_n7522));
  nand_5 g07146(.A(pi105), .B(pi032), .Y(new_n7523));
  not_8  g07147(.A(new_n7428), .Y(new_n7524));
  nor_5  g07148(.A(new_n7429), .B(new_n7524), .Y(new_n7525));
  not_8  g07149(.A(new_n7393), .Y(new_n7526));
  nor_5  g07150(.A(new_n7430), .B(new_n7526), .Y(new_n7527));
  nor_5  g07151(.A(new_n7527), .B(new_n7525), .Y(new_n7528));
  xor_4  g07152(.A(new_n7528), .B(new_n7523), .Y(new_n7529));
  nand_5 g07153(.A(pi077), .B(pi072), .Y(new_n7530));
  nand_5 g07154(.A(pi208), .B(pi166), .Y(new_n7531));
  xor_4  g07155(.A(new_n7531), .B(new_n7530), .Y(new_n7532));
  xor_4  g07156(.A(new_n7532), .B(new_n7529), .Y(new_n7533));
  xor_4  g07157(.A(new_n7533), .B(new_n7522), .Y(new_n7534));
  xor_4  g07158(.A(new_n7534), .B(new_n7521), .Y(new_n7535));
  nand_5 g07159(.A(pi204), .B(pi019), .Y(new_n7536));
  nand_5 g07160(.A(pi168), .B(pi011), .Y(new_n7537));
  nand_5 g07161(.A(new_n7421), .B(new_n7420), .Y(new_n7538));
  nand_5 g07162(.A(new_n7422), .B(new_n7400), .Y(new_n7539));
  nand_5 g07163(.A(new_n7539), .B(new_n7538), .Y(new_n7540));
  xnor_4 g07164(.A(new_n7540), .B(new_n7537), .Y(new_n7541));
  nand_5 g07165(.A(pi097), .B(pi015), .Y(new_n7542));
  nand_5 g07166(.A(pi164), .B(pi088), .Y(new_n7543));
  xor_4  g07167(.A(new_n7543), .B(new_n7542), .Y(new_n7544));
  xor_4  g07168(.A(new_n7544), .B(new_n7541), .Y(new_n7545));
  xor_4  g07169(.A(new_n7545), .B(new_n7536), .Y(new_n7546));
  xor_4  g07170(.A(new_n7546), .B(new_n7535), .Y(new_n7547));
  xor_4  g07171(.A(new_n7547), .B(new_n7457), .Y(new_n7548));
  nand_5 g07172(.A(pi189), .B(pi044), .Y(new_n7549));
  nand_5 g07173(.A(pi072), .B(pi052), .Y(new_n7550));
  nand_5 g07174(.A(pi248), .B(pi131), .Y(new_n7551));
  nand_5 g07175(.A(new_n7551), .B(new_n7550), .Y(new_n7552));
  nand_5 g07176(.A(pi077), .B(pi054), .Y(new_n7553));
  xor_4  g07177(.A(new_n7551), .B(new_n7550), .Y(new_n7554));
  nand_5 g07178(.A(new_n7554), .B(new_n7553), .Y(new_n7555));
  nand_5 g07179(.A(new_n7555), .B(new_n7552), .Y(new_n7556));
  xor_4  g07180(.A(new_n7554), .B(new_n7553), .Y(new_n7557));
  nand_5 g07181(.A(pi250), .B(pi133), .Y(new_n7558));
  nand_5 g07182(.A(pi189), .B(pi045), .Y(new_n7559));
  nand_5 g07183(.A(pi119), .B(pi064), .Y(new_n7560));
  nand_5 g07184(.A(new_n7560), .B(new_n7559), .Y(new_n7561));
  nand_5 g07185(.A(pi189), .B(pi119), .Y(new_n7562));
  nand_5 g07186(.A(pi064), .B(pi045), .Y(new_n7563));
  or_6   g07187(.A(new_n7563), .B(new_n7562), .Y(new_n7564));
  nand_5 g07188(.A(new_n7564), .B(new_n7561), .Y(new_n7565));
  nand_5 g07189(.A(new_n7565), .B(new_n7558), .Y(new_n7566));
  nand_5 g07190(.A(pi250), .B(pi077), .Y(new_n7567));
  nand_5 g07191(.A(new_n7567), .B(new_n7562), .Y(new_n7568));
  nand_5 g07192(.A(pi133), .B(pi045), .Y(new_n7569));
  xor_4  g07193(.A(new_n7567), .B(new_n7562), .Y(new_n7570));
  nand_5 g07194(.A(new_n7570), .B(new_n7569), .Y(new_n7571));
  nand_5 g07195(.A(new_n7571), .B(new_n7568), .Y(new_n7572));
  xor_4  g07196(.A(new_n7565), .B(new_n7558), .Y(new_n7573));
  nand_5 g07197(.A(new_n7573), .B(new_n7572), .Y(new_n7574));
  nand_5 g07198(.A(new_n7574), .B(new_n7566), .Y(new_n7575));
  xor_4  g07199(.A(new_n7575), .B(new_n7557), .Y(new_n7576));
  nand_5 g07200(.A(pi250), .B(pi189), .Y(new_n7577));
  nand_5 g07201(.A(pi119), .B(pi084), .Y(new_n7578));
  xor_4  g07202(.A(new_n7578), .B(new_n7577), .Y(new_n7579));
  xor_4  g07203(.A(new_n7579), .B(new_n7563), .Y(new_n7580));
  nand_5 g07204(.A(pi133), .B(pi044), .Y(new_n7581));
  xor_4  g07205(.A(new_n7581), .B(new_n7564), .Y(new_n7582));
  xor_4  g07206(.A(new_n7582), .B(new_n7580), .Y(new_n7583));
  xor_4  g07207(.A(new_n7583), .B(new_n7576), .Y(new_n7584));
  nand_5 g07208(.A(pi077), .B(pi044), .Y(new_n7585));
  nand_5 g07209(.A(pi054), .B(pi052), .Y(new_n7586));
  nand_5 g07210(.A(new_n7586), .B(new_n7585), .Y(new_n7587));
  nand_5 g07211(.A(pi052), .B(pi044), .Y(new_n7588));
  nor_5  g07212(.A(new_n7588), .B(new_n7553), .Y(new_n7589));
  not_8  g07213(.A(new_n7589), .Y(new_n7590));
  nand_5 g07214(.A(new_n7590), .B(new_n7587), .Y(new_n7591));
  xor_4  g07215(.A(new_n7573), .B(new_n7572), .Y(new_n7592));
  nor_5  g07216(.A(new_n7592), .B(new_n7591), .Y(new_n7593));
  xor_4  g07217(.A(new_n7592), .B(new_n7591), .Y(new_n7594));
  not_8  g07218(.A(new_n7594), .Y(new_n7595));
  nand_5 g07219(.A(pi133), .B(pi119), .Y(new_n7596));
  nand_5 g07220(.A(pi077), .B(pi045), .Y(new_n7597));
  nand_5 g07221(.A(new_n7597), .B(new_n7596), .Y(new_n7598));
  nand_5 g07222(.A(pi250), .B(pi052), .Y(new_n7599));
  xor_4  g07223(.A(new_n7597), .B(new_n7596), .Y(new_n7600));
  nand_5 g07224(.A(new_n7600), .B(new_n7599), .Y(new_n7601));
  nand_5 g07225(.A(new_n7601), .B(new_n7598), .Y(new_n7602));
  nand_5 g07226(.A(new_n7602), .B(new_n7588), .Y(new_n7603));
  xor_4  g07227(.A(new_n7570), .B(new_n7569), .Y(new_n7604));
  xor_4  g07228(.A(new_n7602), .B(new_n7588), .Y(new_n7605));
  nand_5 g07229(.A(new_n7605), .B(new_n7604), .Y(new_n7606));
  nand_5 g07230(.A(new_n7606), .B(new_n7603), .Y(new_n7607));
  nor_5  g07231(.A(new_n7607), .B(new_n7595), .Y(new_n7608));
  xor_4  g07232(.A(new_n7608), .B(new_n7590), .Y(new_n7609));
  not_8  g07233(.A(new_n7609), .Y(new_n7610));
  nor_5  g07234(.A(new_n7610), .B(new_n7593), .Y(new_n7611));
  xor_4  g07235(.A(new_n7611), .B(new_n7584), .Y(new_n7612));
  nand_5 g07236(.A(pi131), .B(pi054), .Y(new_n7613));
  nand_5 g07237(.A(pi131), .B(pi044), .Y(new_n7614));
  nand_5 g07238(.A(pi250), .B(pi131), .Y(new_n7615));
  nand_5 g07239(.A(pi052), .B(pi045), .Y(new_n7616));
  nand_5 g07240(.A(new_n7616), .B(new_n7615), .Y(new_n7617));
  nand_5 g07241(.A(pi119), .B(pi077), .Y(new_n7618));
  xor_4  g07242(.A(new_n7616), .B(new_n7615), .Y(new_n7619));
  nand_5 g07243(.A(new_n7619), .B(new_n7618), .Y(new_n7620));
  nand_5 g07244(.A(new_n7620), .B(new_n7617), .Y(new_n7621));
  nand_5 g07245(.A(new_n7621), .B(new_n7614), .Y(new_n7622));
  xor_4  g07246(.A(new_n7600), .B(new_n7599), .Y(new_n7623));
  xor_4  g07247(.A(new_n7621), .B(new_n7614), .Y(new_n7624));
  nand_5 g07248(.A(new_n7624), .B(new_n7623), .Y(new_n7625));
  nand_5 g07249(.A(new_n7625), .B(new_n7622), .Y(new_n7626));
  nor_5  g07250(.A(new_n7626), .B(new_n7613), .Y(new_n7627));
  xor_4  g07251(.A(new_n7626), .B(new_n7613), .Y(new_n7628));
  xor_4  g07252(.A(new_n7605), .B(new_n7604), .Y(new_n7629));
  not_8  g07253(.A(new_n7629), .Y(new_n7630));
  nand_5 g07254(.A(new_n7630), .B(new_n7628), .Y(new_n7631));
  not_8  g07255(.A(new_n7631), .Y(new_n7632));
  nor_5  g07256(.A(new_n7632), .B(new_n7627), .Y(new_n7633));
  xor_4  g07257(.A(new_n7607), .B(new_n7594), .Y(new_n7634));
  nor_5  g07258(.A(new_n7634), .B(new_n7633), .Y(new_n7635));
  nor_5  g07259(.A(new_n7635), .B(new_n7612), .Y(new_n7636));
  xor_4  g07260(.A(new_n7635), .B(new_n7612), .Y(new_n7637));
  nand_5 g07261(.A(pi131), .B(pi072), .Y(new_n7638));
  xor_4  g07262(.A(new_n7630), .B(new_n7628), .Y(new_n7639));
  xor_4  g07263(.A(new_n7619), .B(new_n7618), .Y(new_n7640));
  not_8  g07264(.A(new_n7640), .Y(new_n7641));
  nand_5 g07265(.A(pi131), .B(pi045), .Y(new_n7642));
  nand_5 g07266(.A(pi119), .B(pi052), .Y(new_n7643));
  nor_5  g07267(.A(new_n7643), .B(new_n7642), .Y(new_n7644));
  nand_5 g07268(.A(new_n7644), .B(new_n7641), .Y(new_n7645));
  xor_4  g07269(.A(new_n7624), .B(new_n7623), .Y(new_n7646));
  nor_5  g07270(.A(new_n7646), .B(new_n7645), .Y(new_n7647));
  nand_5 g07271(.A(new_n7647), .B(new_n7639), .Y(new_n7648));
  nand_5 g07272(.A(new_n7648), .B(new_n7638), .Y(new_n7649));
  xor_4  g07273(.A(new_n7648), .B(new_n7638), .Y(new_n7650));
  xor_4  g07274(.A(new_n7634), .B(new_n7633), .Y(new_n7651));
  not_8  g07275(.A(new_n7651), .Y(new_n7652));
  nand_5 g07276(.A(new_n7652), .B(new_n7650), .Y(new_n7653));
  nand_5 g07277(.A(new_n7653), .B(new_n7649), .Y(new_n7654));
  and_6  g07278(.A(new_n7654), .B(new_n7637), .Y(new_n7655));
  nor_5  g07279(.A(new_n7655), .B(new_n7636), .Y(new_n7656));
  xor_4  g07280(.A(new_n7656), .B(new_n7556), .Y(new_n7657));
  xor_4  g07281(.A(new_n7657), .B(new_n7549), .Y(new_n7658));
  xor_4  g07282(.A(new_n7658), .B(new_n7548), .Y(new_n7659));
  nand_5 g07283(.A(pi084), .B(pi045), .Y(new_n7660));
  nand_5 g07284(.A(pi236), .B(pi096), .Y(new_n7661));
  nand_5 g07285(.A(pi241), .B(pi026), .Y(new_n7662));
  nand_5 g07286(.A(pi161), .B(pi027), .Y(new_n7663));
  nand_5 g07287(.A(pi236), .B(pi008), .Y(new_n7664));
  nor_5  g07288(.A(new_n7664), .B(new_n7663), .Y(new_n7665));
  nor_5  g07289(.A(new_n7662), .B(new_n378), .Y(new_n7666));
  nand_5 g07290(.A(new_n7664), .B(new_n7663), .Y(new_n7667));
  nor_5  g07291(.A(new_n7667), .B(new_n7666), .Y(new_n7668));
  nor_5  g07292(.A(new_n7668), .B(new_n7665), .Y(new_n7669));
  nor_5  g07293(.A(new_n7669), .B(new_n7662), .Y(new_n7670));
  nand_5 g07294(.A(pi161), .B(pi026), .Y(new_n7671));
  nand_5 g07295(.A(pi141), .B(pi027), .Y(new_n7672));
  nand_5 g07296(.A(pi241), .B(pi008), .Y(new_n7673));
  xor_4  g07297(.A(new_n7673), .B(new_n7672), .Y(new_n7674));
  xor_4  g07298(.A(new_n7674), .B(new_n7671), .Y(new_n7675));
  not_8  g07299(.A(new_n7662), .Y(new_n7676));
  or_6   g07300(.A(new_n7665), .B(new_n7676), .Y(new_n7677));
  nand_5 g07301(.A(new_n7677), .B(new_n7667), .Y(new_n7678));
  nand_5 g07302(.A(pi236), .B(pi056), .Y(new_n7679));
  xnor_4 g07303(.A(new_n7679), .B(new_n7678), .Y(new_n7680));
  xor_4  g07304(.A(new_n7680), .B(new_n7675), .Y(new_n7681));
  nand_5 g07305(.A(new_n7681), .B(new_n7670), .Y(new_n7682));
  not_8  g07306(.A(new_n7682), .Y(new_n7683));
  nor_5  g07307(.A(new_n7679), .B(new_n7678), .Y(new_n7684));
  nor_5  g07308(.A(new_n7680), .B(new_n7675), .Y(new_n7685));
  nor_5  g07309(.A(new_n7685), .B(new_n7684), .Y(new_n7686));
  nand_5 g07310(.A(pi236), .B(pi136), .Y(new_n7687));
  nand_5 g07311(.A(pi161), .B(pi008), .Y(new_n7688));
  nand_5 g07312(.A(pi090), .B(pi027), .Y(new_n7689));
  nand_5 g07313(.A(pi141), .B(pi026), .Y(new_n7690));
  xor_4  g07314(.A(new_n7690), .B(new_n7689), .Y(new_n7691));
  xor_4  g07315(.A(new_n7691), .B(new_n7688), .Y(new_n7692));
  nand_5 g07316(.A(pi241), .B(pi056), .Y(new_n7693));
  nand_5 g07317(.A(new_n7673), .B(new_n7672), .Y(new_n7694));
  nand_5 g07318(.A(new_n7674), .B(new_n7671), .Y(new_n7695));
  nand_5 g07319(.A(new_n7695), .B(new_n7694), .Y(new_n7696));
  xor_4  g07320(.A(new_n7696), .B(new_n7693), .Y(new_n7697));
  xnor_4 g07321(.A(new_n7697), .B(new_n7692), .Y(new_n7698));
  xor_4  g07322(.A(new_n7698), .B(new_n7687), .Y(new_n7699));
  xor_4  g07323(.A(new_n7699), .B(new_n7686), .Y(new_n7700));
  nand_5 g07324(.A(new_n7700), .B(new_n7683), .Y(new_n7701));
  nand_5 g07325(.A(new_n7701), .B(new_n7661), .Y(new_n7702));
  xor_4  g07326(.A(new_n7701), .B(new_n7661), .Y(new_n7703));
  not_8  g07327(.A(new_n7698), .Y(new_n7704));
  nor_5  g07328(.A(new_n7704), .B(new_n7687), .Y(new_n7705));
  nor_5  g07329(.A(new_n7699), .B(new_n7686), .Y(new_n7706));
  or_6   g07330(.A(new_n7706), .B(new_n7705), .Y(new_n7707));
  nand_5 g07331(.A(pi241), .B(pi136), .Y(new_n7708));
  nand_5 g07332(.A(pi161), .B(pi056), .Y(new_n7709));
  and_6  g07333(.A(new_n7709), .B(new_n7708), .Y(new_n7710));
  nand_5 g07334(.A(pi161), .B(pi136), .Y(new_n7711));
  nor_5  g07335(.A(new_n7711), .B(new_n7693), .Y(new_n7712));
  or_6   g07336(.A(new_n7712), .B(new_n7710), .Y(new_n7713));
  nand_5 g07337(.A(new_n7690), .B(new_n7689), .Y(new_n7714));
  nand_5 g07338(.A(new_n7691), .B(new_n7688), .Y(new_n7715));
  nand_5 g07339(.A(new_n7715), .B(new_n7714), .Y(new_n7716));
  nand_5 g07340(.A(pi047), .B(pi026), .Y(new_n7717));
  nor_5  g07341(.A(new_n7717), .B(new_n7689), .Y(new_n7718));
  not_8  g07342(.A(new_n7718), .Y(new_n7719));
  nand_5 g07343(.A(pi047), .B(pi027), .Y(new_n7720));
  nand_5 g07344(.A(pi090), .B(pi026), .Y(new_n7721));
  nand_5 g07345(.A(new_n7721), .B(new_n7720), .Y(new_n7722));
  nand_5 g07346(.A(new_n7722), .B(new_n7719), .Y(new_n7723));
  nand_5 g07347(.A(pi141), .B(pi008), .Y(new_n7724));
  xor_4  g07348(.A(new_n7724), .B(new_n7723), .Y(new_n7725));
  xor_4  g07349(.A(new_n7725), .B(new_n7716), .Y(new_n7726));
  xor_4  g07350(.A(new_n7726), .B(new_n7713), .Y(new_n7727));
  nand_5 g07351(.A(new_n7696), .B(new_n7693), .Y(new_n7728));
  nand_5 g07352(.A(new_n7697), .B(new_n7692), .Y(new_n7729));
  nand_5 g07353(.A(new_n7729), .B(new_n7728), .Y(new_n7730));
  xor_4  g07354(.A(new_n7730), .B(new_n7727), .Y(new_n7731));
  xor_4  g07355(.A(new_n7731), .B(new_n7707), .Y(new_n7732));
  nand_5 g07356(.A(new_n7732), .B(new_n7703), .Y(new_n7733));
  nand_5 g07357(.A(new_n7733), .B(new_n7702), .Y(new_n7734));
  not_8  g07358(.A(new_n7731), .Y(new_n7735));
  nand_5 g07359(.A(new_n7735), .B(new_n7707), .Y(new_n7736));
  nor_5  g07360(.A(new_n7726), .B(new_n7713), .Y(new_n7737));
  not_8  g07361(.A(new_n7727), .Y(new_n7738));
  nor_5  g07362(.A(new_n7730), .B(new_n7738), .Y(new_n7739));
  xor_4  g07363(.A(new_n7739), .B(new_n7712), .Y(new_n7740));
  nor_5  g07364(.A(new_n7740), .B(new_n7737), .Y(new_n7741));
  nand_5 g07365(.A(pi241), .B(pi096), .Y(new_n7742));
  nand_5 g07366(.A(pi236), .B(pi235), .Y(new_n7743));
  xor_4  g07367(.A(new_n7743), .B(new_n7742), .Y(new_n7744));
  xor_4  g07368(.A(new_n7744), .B(new_n7711), .Y(new_n7745));
  nand_5 g07369(.A(new_n7724), .B(new_n7723), .Y(new_n7746));
  nand_5 g07370(.A(new_n7725), .B(new_n7716), .Y(new_n7747));
  nand_5 g07371(.A(new_n7747), .B(new_n7746), .Y(new_n7748));
  xor_4  g07372(.A(new_n7748), .B(new_n7745), .Y(new_n7749));
  nand_5 g07373(.A(pi141), .B(pi056), .Y(new_n7750));
  xor_4  g07374(.A(new_n7750), .B(new_n7718), .Y(new_n7751));
  nand_5 g07375(.A(pi027), .B(pi018), .Y(new_n7752));
  nand_5 g07376(.A(pi090), .B(pi008), .Y(new_n7753));
  xor_4  g07377(.A(new_n7753), .B(new_n7752), .Y(new_n7754));
  xor_4  g07378(.A(new_n7754), .B(new_n7717), .Y(new_n7755));
  xor_4  g07379(.A(new_n7755), .B(new_n7751), .Y(new_n7756));
  not_8  g07380(.A(new_n7756), .Y(new_n7757));
  xor_4  g07381(.A(new_n7757), .B(new_n7749), .Y(new_n7758));
  xor_4  g07382(.A(new_n7758), .B(new_n7741), .Y(new_n7759));
  xor_4  g07383(.A(new_n7759), .B(new_n7736), .Y(new_n7760));
  xnor_4 g07384(.A(new_n7760), .B(new_n7734), .Y(new_n7761));
  nand_5 g07385(.A(pi213), .B(pi114), .Y(new_n7762));
  nand_5 g07386(.A(pi246), .B(pi213), .Y(new_n7763));
  xor_4  g07387(.A(new_n7474), .B(new_n7473), .Y(new_n7764));
  xnor_4 g07388(.A(new_n7764), .B(new_n7763), .Y(new_n7765));
  nand_5 g07389(.A(pi213), .B(pi145), .Y(new_n7766));
  nand_5 g07390(.A(pi213), .B(pi032), .Y(new_n7767));
  nand_5 g07391(.A(pi212), .B(pi206), .Y(new_n7768));
  nand_5 g07392(.A(new_n7768), .B(new_n7767), .Y(new_n7769));
  nand_5 g07393(.A(pi164), .B(pi104), .Y(new_n7770));
  xor_4  g07394(.A(new_n7768), .B(new_n7767), .Y(new_n7771));
  nand_5 g07395(.A(new_n7771), .B(new_n7770), .Y(new_n7772));
  nand_5 g07396(.A(new_n7772), .B(new_n7769), .Y(new_n7773));
  nand_5 g07397(.A(new_n7773), .B(new_n7766), .Y(new_n7774));
  xor_4  g07398(.A(new_n7465), .B(new_n7464), .Y(new_n7775));
  xor_4  g07399(.A(new_n7773), .B(new_n7766), .Y(new_n7776));
  nand_5 g07400(.A(new_n7776), .B(new_n7775), .Y(new_n7777));
  nand_5 g07401(.A(new_n7777), .B(new_n7774), .Y(new_n7778));
  xor_4  g07402(.A(new_n7778), .B(new_n7765), .Y(new_n7779));
  xor_4  g07403(.A(new_n7776), .B(new_n7775), .Y(new_n7780));
  xor_4  g07404(.A(new_n7771), .B(new_n7770), .Y(new_n7781));
  or_6   g07405(.A(new_n7768), .B(new_n380), .Y(new_n7782));
  nor_5  g07406(.A(new_n7782), .B(new_n7781), .Y(new_n7783));
  not_8  g07407(.A(new_n7783), .Y(new_n7784));
  nor_5  g07408(.A(new_n7784), .B(new_n7780), .Y(new_n7785));
  nand_5 g07409(.A(new_n7785), .B(new_n7779), .Y(new_n7786));
  nand_5 g07410(.A(new_n7786), .B(new_n7762), .Y(new_n7787));
  xor_4  g07411(.A(new_n7786), .B(new_n7762), .Y(new_n7788));
  nor_5  g07412(.A(new_n7764), .B(new_n7763), .Y(new_n7789));
  nor_5  g07413(.A(new_n7778), .B(new_n7765), .Y(new_n7790));
  nor_5  g07414(.A(new_n7790), .B(new_n7789), .Y(new_n7791));
  xor_4  g07415(.A(new_n7495), .B(new_n7476), .Y(new_n7792));
  xor_4  g07416(.A(new_n7792), .B(new_n7791), .Y(new_n7793));
  nand_5 g07417(.A(new_n7793), .B(new_n7788), .Y(new_n7794));
  nand_5 g07418(.A(new_n7794), .B(new_n7787), .Y(new_n7795));
  not_8  g07419(.A(new_n7792), .Y(new_n7796));
  nor_5  g07420(.A(new_n7796), .B(new_n7791), .Y(new_n7797));
  xor_4  g07421(.A(new_n7519), .B(new_n7515), .Y(new_n7798));
  or_6   g07422(.A(new_n7798), .B(new_n7797), .Y(new_n7799));
  nand_5 g07423(.A(new_n7798), .B(new_n7797), .Y(new_n7800));
  nand_5 g07424(.A(new_n7800), .B(new_n7799), .Y(new_n7801));
  xnor_4 g07425(.A(new_n7801), .B(new_n7795), .Y(new_n7802));
  nand_5 g07426(.A(new_n7802), .B(new_n7761), .Y(new_n7803));
  xor_4  g07427(.A(new_n7802), .B(new_n7761), .Y(new_n7804));
  xor_4  g07428(.A(new_n7732), .B(new_n7703), .Y(new_n7805));
  not_8  g07429(.A(new_n7805), .Y(new_n7806));
  xnor_4 g07430(.A(new_n7793), .B(new_n7788), .Y(new_n7807));
  nand_5 g07431(.A(new_n7807), .B(new_n7806), .Y(new_n7808));
  xor_4  g07432(.A(new_n7807), .B(new_n7805), .Y(new_n7809));
  not_8  g07433(.A(new_n7809), .Y(new_n7810));
  xnor_4 g07434(.A(new_n7782), .B(new_n7781), .Y(new_n7811));
  nand_5 g07435(.A(new_n7667), .B(new_n7666), .Y(new_n7812));
  nand_5 g07436(.A(new_n7812), .B(new_n7669), .Y(new_n7813));
  nor_5  g07437(.A(new_n7813), .B(new_n7811), .Y(new_n7814));
  or_6   g07438(.A(new_n380), .B(new_n379), .Y(new_n7815));
  nand_5 g07439(.A(pi241), .B(pi027), .Y(new_n7816));
  nor_5  g07440(.A(new_n1063), .B(new_n561), .Y(new_n7817));
  xor_4  g07441(.A(new_n7817), .B(new_n7816), .Y(new_n7818));
  nor_5  g07442(.A(new_n7818), .B(new_n7815), .Y(new_n7819));
  xnor_4 g07443(.A(new_n7818), .B(new_n7815), .Y(new_n7820));
  nand_5 g07444(.A(pi213), .B(pi206), .Y(new_n7821));
  nand_5 g07445(.A(pi212), .B(pi164), .Y(new_n7822));
  nand_5 g07446(.A(new_n7822), .B(new_n7821), .Y(new_n7823));
  nand_5 g07447(.A(new_n7823), .B(new_n7782), .Y(new_n7824));
  nor_5  g07448(.A(new_n7824), .B(new_n7820), .Y(new_n7825));
  nor_5  g07449(.A(new_n7825), .B(new_n7819), .Y(new_n7826));
  xnor_4 g07450(.A(new_n7813), .B(new_n7811), .Y(new_n7827));
  nor_5  g07451(.A(new_n7827), .B(new_n7826), .Y(new_n7828));
  nor_5  g07452(.A(new_n7828), .B(new_n7814), .Y(new_n7829));
  not_8  g07453(.A(new_n7829), .Y(new_n7830));
  xor_4  g07454(.A(new_n7681), .B(new_n7670), .Y(new_n7831));
  nor_5  g07455(.A(new_n7831), .B(new_n7830), .Y(new_n7832));
  xor_4  g07456(.A(new_n7784), .B(new_n7780), .Y(new_n7833));
  xor_4  g07457(.A(new_n7831), .B(new_n7829), .Y(new_n7834));
  nor_5  g07458(.A(new_n7834), .B(new_n7833), .Y(new_n7835));
  or_6   g07459(.A(new_n7835), .B(new_n7832), .Y(new_n7836));
  xor_4  g07460(.A(new_n7700), .B(new_n7682), .Y(new_n7837));
  and_6  g07461(.A(new_n7837), .B(new_n7836), .Y(new_n7838));
  xor_4  g07462(.A(new_n7785), .B(new_n7779), .Y(new_n7839));
  not_8  g07463(.A(new_n7839), .Y(new_n7840));
  xor_4  g07464(.A(new_n7837), .B(new_n7836), .Y(new_n7841));
  and_6  g07465(.A(new_n7841), .B(new_n7840), .Y(new_n7842));
  nor_5  g07466(.A(new_n7842), .B(new_n7838), .Y(new_n7843));
  nand_5 g07467(.A(new_n7843), .B(new_n7810), .Y(new_n7844));
  nand_5 g07468(.A(new_n7844), .B(new_n7808), .Y(new_n7845));
  not_8  g07469(.A(new_n7845), .Y(new_n7846));
  nand_5 g07470(.A(new_n7846), .B(new_n7804), .Y(new_n7847));
  nand_5 g07471(.A(new_n7847), .B(new_n7803), .Y(new_n7848));
  xor_4  g07472(.A(new_n7848), .B(new_n7660), .Y(new_n7849));
  nor_5  g07473(.A(new_n7750), .B(new_n7719), .Y(new_n7850));
  nor_5  g07474(.A(new_n7755), .B(new_n7751), .Y(new_n7851));
  nor_5  g07475(.A(new_n7851), .B(new_n7850), .Y(new_n7852));
  nand_5 g07476(.A(pi161), .B(pi096), .Y(new_n7853));
  nand_5 g07477(.A(pi131), .B(pi009), .Y(new_n7854));
  xor_4  g07478(.A(new_n7854), .B(new_n7853), .Y(new_n7855));
  xor_4  g07479(.A(new_n7855), .B(new_n7852), .Y(new_n7856));
  xor_4  g07480(.A(new_n7856), .B(new_n7849), .Y(new_n7857));
  xor_4  g07481(.A(new_n7857), .B(new_n7659), .Y(new_n7858));
  nor_5  g07482(.A(new_n7416), .B(new_n7395), .Y(new_n7859));
  nor_5  g07483(.A(new_n7433), .B(new_n7417), .Y(new_n7860));
  nor_5  g07484(.A(new_n7860), .B(new_n7859), .Y(new_n7861));
  nand_5 g07485(.A(pi250), .B(pi064), .Y(new_n7862));
  nand_5 g07486(.A(pi151), .B(pi146), .Y(new_n7863));
  xor_4  g07487(.A(new_n7863), .B(new_n7862), .Y(new_n7864));
  xor_4  g07488(.A(new_n7864), .B(new_n7861), .Y(new_n7865));
  nand_5 g07489(.A(pi133), .B(pi054), .Y(new_n7866));
  nand_5 g07490(.A(pi246), .B(pi013), .Y(new_n7867));
  xor_4  g07491(.A(new_n7867), .B(new_n7866), .Y(new_n7868));
  xor_4  g07492(.A(new_n7868), .B(new_n7865), .Y(new_n7869));
  xor_4  g07493(.A(new_n7654), .B(new_n7637), .Y(new_n7870));
  xor_4  g07494(.A(new_n7841), .B(new_n7839), .Y(new_n7871));
  xor_4  g07495(.A(new_n7447), .B(new_n7446), .Y(new_n7872));
  xor_4  g07496(.A(new_n7872), .B(new_n7871), .Y(new_n7873));
  xor_4  g07497(.A(new_n7834), .B(new_n7833), .Y(new_n7874));
  xor_4  g07498(.A(new_n7444), .B(new_n7443), .Y(new_n7875));
  nand_5 g07499(.A(new_n7875), .B(new_n7874), .Y(new_n7876));
  nand_5 g07500(.A(new_n7440), .B(new_n7354), .Y(new_n7877));
  and_6  g07501(.A(new_n7877), .B(new_n7442), .Y(new_n7878));
  xor_4  g07502(.A(new_n7827), .B(new_n7826), .Y(new_n7879));
  nor_5  g07503(.A(new_n7879), .B(new_n7878), .Y(new_n7880));
  xnor_4 g07504(.A(new_n7879), .B(new_n7878), .Y(new_n7881));
  nand_5 g07505(.A(new_n381), .B(new_n7439), .Y(new_n7882));
  not_8  g07506(.A(new_n7882), .Y(new_n7883));
  nand_5 g07507(.A(pi168), .B(pi151), .Y(new_n7884));
  nand_5 g07508(.A(pi208), .B(pi147), .Y(new_n7885));
  xor_4  g07509(.A(new_n7885), .B(new_n7884), .Y(new_n7886));
  nor_5  g07510(.A(new_n7886), .B(new_n7883), .Y(new_n7887));
  xor_4  g07511(.A(new_n7824), .B(new_n7820), .Y(new_n7888));
  xor_4  g07512(.A(new_n7886), .B(new_n7882), .Y(new_n7889));
  nor_5  g07513(.A(new_n7889), .B(new_n7888), .Y(new_n7890));
  nor_5  g07514(.A(new_n7890), .B(new_n7887), .Y(new_n7891));
  nor_5  g07515(.A(new_n7891), .B(new_n7881), .Y(new_n7892));
  nor_5  g07516(.A(new_n7892), .B(new_n7880), .Y(new_n7893));
  xnor_4 g07517(.A(new_n7875), .B(new_n7874), .Y(new_n7894));
  or_6   g07518(.A(new_n7894), .B(new_n7893), .Y(new_n7895));
  nand_5 g07519(.A(new_n7895), .B(new_n7876), .Y(new_n7896));
  xor_4  g07520(.A(new_n7896), .B(new_n7873), .Y(new_n7897));
  xor_4  g07521(.A(new_n7647), .B(new_n7639), .Y(new_n7898));
  not_8  g07522(.A(new_n7898), .Y(new_n7899));
  or_6   g07523(.A(new_n7899), .B(new_n7897), .Y(new_n7900));
  xor_4  g07524(.A(new_n7646), .B(new_n7645), .Y(new_n7901));
  xnor_4 g07525(.A(new_n7894), .B(new_n7893), .Y(new_n7902));
  nand_5 g07526(.A(new_n7902), .B(new_n7901), .Y(new_n7903));
  xor_4  g07527(.A(new_n7902), .B(new_n7901), .Y(new_n7904));
  nor_5  g07528(.A(new_n383), .B(new_n382), .Y(new_n7905));
  xor_4  g07529(.A(new_n7643), .B(new_n7642), .Y(new_n7906));
  nor_5  g07530(.A(new_n7906), .B(new_n7905), .Y(new_n7907));
  xor_4  g07531(.A(new_n7906), .B(new_n7905), .Y(new_n7908));
  not_8  g07532(.A(new_n7908), .Y(new_n7909));
  xnor_4 g07533(.A(new_n7889), .B(new_n7888), .Y(new_n7910));
  nor_5  g07534(.A(new_n7910), .B(new_n7909), .Y(new_n7911));
  nor_5  g07535(.A(new_n7911), .B(new_n7907), .Y(new_n7912));
  not_8  g07536(.A(new_n7912), .Y(new_n7913));
  xor_4  g07537(.A(new_n7891), .B(new_n7881), .Y(new_n7914));
  and_6  g07538(.A(new_n7914), .B(new_n7913), .Y(new_n7915));
  xor_4  g07539(.A(new_n7644), .B(new_n7641), .Y(new_n7916));
  xor_4  g07540(.A(new_n7914), .B(new_n7912), .Y(new_n7917));
  nor_5  g07541(.A(new_n7917), .B(new_n7916), .Y(new_n7918));
  nor_5  g07542(.A(new_n7918), .B(new_n7915), .Y(new_n7919));
  nand_5 g07543(.A(new_n7919), .B(new_n7904), .Y(new_n7920));
  nand_5 g07544(.A(new_n7920), .B(new_n7903), .Y(new_n7921));
  xor_4  g07545(.A(new_n7899), .B(new_n7897), .Y(new_n7922));
  nand_5 g07546(.A(new_n7922), .B(new_n7921), .Y(new_n7923));
  nand_5 g07547(.A(new_n7923), .B(new_n7900), .Y(new_n7924));
  xor_4  g07548(.A(new_n7651), .B(new_n7650), .Y(new_n7925));
  and_6  g07549(.A(new_n7925), .B(new_n7924), .Y(new_n7926));
  xnor_4 g07550(.A(new_n7925), .B(new_n7924), .Y(new_n7927));
  nor_5  g07551(.A(new_n7872), .B(new_n7871), .Y(new_n7928));
  and_6  g07552(.A(new_n7896), .B(new_n7873), .Y(new_n7929));
  nor_5  g07553(.A(new_n7929), .B(new_n7928), .Y(new_n7930));
  xor_4  g07554(.A(new_n7452), .B(new_n7451), .Y(new_n7931));
  xor_4  g07555(.A(new_n7843), .B(new_n7810), .Y(new_n7932));
  xnor_4 g07556(.A(new_n7932), .B(new_n7931), .Y(new_n7933));
  xor_4  g07557(.A(new_n7933), .B(new_n7930), .Y(new_n7934));
  nor_5  g07558(.A(new_n7934), .B(new_n7927), .Y(new_n7935));
  nor_5  g07559(.A(new_n7935), .B(new_n7926), .Y(new_n7936));
  nand_5 g07560(.A(new_n7936), .B(new_n7870), .Y(new_n7937));
  xor_4  g07561(.A(new_n7846), .B(new_n7804), .Y(new_n7938));
  xor_4  g07562(.A(new_n7455), .B(new_n7436), .Y(new_n7939));
  xnor_4 g07563(.A(new_n7939), .B(new_n7938), .Y(new_n7940));
  nor_5  g07564(.A(new_n7932), .B(new_n7931), .Y(new_n7941));
  nor_5  g07565(.A(new_n7933), .B(new_n7930), .Y(new_n7942));
  nor_5  g07566(.A(new_n7942), .B(new_n7941), .Y(new_n7943));
  xor_4  g07567(.A(new_n7943), .B(new_n7940), .Y(new_n7944));
  xor_4  g07568(.A(new_n7936), .B(new_n7870), .Y(new_n7945));
  nand_5 g07569(.A(new_n7945), .B(new_n7944), .Y(new_n7946));
  nand_5 g07570(.A(new_n7946), .B(new_n7937), .Y(new_n7947));
  nand_5 g07571(.A(new_n7578), .B(new_n7577), .Y(new_n7948));
  nand_5 g07572(.A(new_n7579), .B(new_n7563), .Y(new_n7949));
  nand_5 g07573(.A(new_n7949), .B(new_n7948), .Y(new_n7950));
  or_6   g07574(.A(new_n7581), .B(new_n7564), .Y(new_n7951));
  not_8  g07575(.A(new_n7580), .Y(new_n7952));
  nand_5 g07576(.A(new_n7582), .B(new_n7952), .Y(new_n7953));
  nand_5 g07577(.A(new_n7953), .B(new_n7951), .Y(new_n7954));
  nand_5 g07578(.A(pi090), .B(pi056), .Y(new_n7955));
  nand_5 g07579(.A(pi236), .B(pi110), .Y(new_n7956));
  xor_4  g07580(.A(new_n7956), .B(new_n7955), .Y(new_n7957));
  xor_4  g07581(.A(new_n7957), .B(new_n7954), .Y(new_n7958));
  xor_4  g07582(.A(new_n7958), .B(new_n7950), .Y(new_n7959));
  and_6  g07583(.A(new_n7739), .B(new_n7712), .Y(new_n7960));
  nor_5  g07584(.A(new_n7758), .B(new_n7741), .Y(new_n7961));
  nor_5  g07585(.A(new_n7961), .B(new_n7960), .Y(new_n7962));
  not_8  g07586(.A(new_n7759), .Y(new_n7963));
  nor_5  g07587(.A(new_n7963), .B(new_n7736), .Y(new_n7964));
  nor_5  g07588(.A(new_n7760), .B(new_n7734), .Y(new_n7965));
  nor_5  g07589(.A(new_n7965), .B(new_n7964), .Y(new_n7966));
  xor_4  g07590(.A(new_n7966), .B(new_n7962), .Y(new_n7967));
  nand_5 g07591(.A(pi128), .B(pi027), .Y(new_n7968));
  nand_5 g07592(.A(pi026), .B(pi018), .Y(new_n7969));
  xor_4  g07593(.A(new_n7969), .B(new_n7968), .Y(new_n7970));
  nand_5 g07594(.A(pi114), .B(pi104), .Y(new_n7971));
  nand_5 g07595(.A(pi047), .B(pi008), .Y(new_n7972));
  xor_4  g07596(.A(new_n7972), .B(new_n7971), .Y(new_n7973));
  xor_4  g07597(.A(new_n7973), .B(new_n7970), .Y(new_n7974));
  xor_4  g07598(.A(new_n7974), .B(new_n7967), .Y(new_n7975));
  xor_4  g07599(.A(new_n7975), .B(new_n7959), .Y(new_n7976));
  xor_4  g07600(.A(new_n7976), .B(new_n7947), .Y(new_n7977));
  xor_4  g07601(.A(new_n7977), .B(new_n7869), .Y(new_n7978));
  xor_4  g07602(.A(new_n7978), .B(new_n7858), .Y(new_n7979));
  nand_5 g07603(.A(new_n7575), .B(new_n7557), .Y(new_n7980));
  nand_5 g07604(.A(new_n7583), .B(new_n7576), .Y(new_n7981));
  nand_5 g07605(.A(new_n7981), .B(new_n7980), .Y(new_n7982));
  nand_5 g07606(.A(pi206), .B(pi183), .Y(new_n7983));
  nand_5 g07607(.A(pi248), .B(pi052), .Y(new_n7984));
  nand_5 g07608(.A(pi139), .B(pi093), .Y(new_n7985));
  xor_4  g07609(.A(new_n7985), .B(new_n7984), .Y(new_n7986));
  xor_4  g07610(.A(new_n7986), .B(new_n7983), .Y(new_n7987));
  xor_4  g07611(.A(new_n7987), .B(new_n7982), .Y(new_n7988));
  nand_5 g07612(.A(pi241), .B(pi235), .Y(new_n7989));
  nor_5  g07613(.A(new_n7418), .B(new_n7402), .Y(new_n7990));
  nor_5  g07614(.A(new_n7423), .B(new_n7419), .Y(new_n7991));
  nor_5  g07615(.A(new_n7991), .B(new_n7990), .Y(new_n7992));
  not_8  g07616(.A(new_n7427), .Y(new_n7993));
  nor_5  g07617(.A(new_n7431), .B(new_n7993), .Y(new_n7994));
  nor_5  g07618(.A(new_n7432), .B(new_n7424), .Y(new_n7995));
  nor_5  g07619(.A(new_n7995), .B(new_n7994), .Y(new_n7996));
  xor_4  g07620(.A(new_n7996), .B(new_n7992), .Y(new_n7997));
  nand_5 g07621(.A(pi075), .B(pi035), .Y(new_n7998));
  nand_5 g07622(.A(new_n7608), .B(new_n7589), .Y(new_n7999));
  or_6   g07623(.A(new_n7611), .B(new_n7584), .Y(new_n8000));
  nand_5 g07624(.A(new_n8000), .B(new_n7999), .Y(new_n8001));
  nand_5 g07625(.A(new_n7743), .B(new_n7742), .Y(new_n8002));
  nand_5 g07626(.A(new_n7744), .B(new_n7711), .Y(new_n8003));
  nand_5 g07627(.A(new_n8003), .B(new_n8002), .Y(new_n8004));
  or_6   g07628(.A(new_n7498), .B(new_n7491), .Y(new_n8005));
  nand_5 g07629(.A(new_n7504), .B(new_n7499), .Y(new_n8006));
  nand_5 g07630(.A(new_n8006), .B(new_n8005), .Y(new_n8007));
  xor_4  g07631(.A(new_n8007), .B(new_n8004), .Y(new_n8008));
  xor_4  g07632(.A(new_n8008), .B(new_n8001), .Y(new_n8009));
  xor_4  g07633(.A(new_n8009), .B(new_n7998), .Y(new_n8010));
  nand_5 g07634(.A(new_n7800), .B(new_n7795), .Y(new_n8011));
  nand_5 g07635(.A(new_n8011), .B(new_n7799), .Y(new_n8012));
  xor_4  g07636(.A(new_n8012), .B(new_n8010), .Y(new_n8013));
  xor_4  g07637(.A(new_n8013), .B(new_n7997), .Y(new_n8014));
  xor_4  g07638(.A(new_n8014), .B(new_n7989), .Y(new_n8015));
  xor_4  g07639(.A(new_n8015), .B(new_n7988), .Y(new_n8016));
  nand_5 g07640(.A(new_n7753), .B(new_n7752), .Y(new_n8017));
  nand_5 g07641(.A(new_n7754), .B(new_n7717), .Y(new_n8018));
  nand_5 g07642(.A(new_n8018), .B(new_n8017), .Y(new_n8019));
  nand_5 g07643(.A(pi119), .B(pi034), .Y(new_n8020));
  xnor_4 g07644(.A(new_n8020), .B(new_n8019), .Y(new_n8021));
  nand_5 g07645(.A(new_n7748), .B(new_n7745), .Y(new_n8022));
  nand_5 g07646(.A(new_n7757), .B(new_n7749), .Y(new_n8023));
  nand_5 g07647(.A(new_n8023), .B(new_n8022), .Y(new_n8024));
  xor_4  g07648(.A(new_n8024), .B(new_n8021), .Y(new_n8025));
  xor_4  g07649(.A(new_n8025), .B(new_n8016), .Y(new_n8026));
  nand_5 g07650(.A(pi145), .B(pi112), .Y(new_n8027));
  nand_5 g07651(.A(pi212), .B(pi091), .Y(new_n8028));
  nand_5 g07652(.A(pi141), .B(pi136), .Y(new_n8029));
  xor_4  g07653(.A(new_n8029), .B(new_n8028), .Y(new_n8030));
  xor_4  g07654(.A(new_n8030), .B(new_n8027), .Y(new_n8031));
  nand_5 g07655(.A(pi152), .B(pi147), .Y(new_n8032));
  nand_5 g07656(.A(new_n7501), .B(new_n7500), .Y(new_n8033));
  nand_5 g07657(.A(new_n7502), .B(new_n7489), .Y(new_n8034));
  nand_5 g07658(.A(new_n8034), .B(new_n8033), .Y(new_n8035));
  xnor_4 g07659(.A(new_n8035), .B(new_n8032), .Y(new_n8036));
  nand_5 g07660(.A(new_n7510), .B(new_n7509), .Y(new_n8037));
  nand_5 g07661(.A(new_n7511), .B(new_n7459), .Y(new_n8038));
  nand_5 g07662(.A(new_n8038), .B(new_n8037), .Y(new_n8039));
  nand_5 g07663(.A(new_n7512), .B(new_n7508), .Y(new_n8040));
  not_8  g07664(.A(new_n7505), .Y(new_n8041));
  nand_5 g07665(.A(new_n7513), .B(new_n8041), .Y(new_n8042));
  nand_5 g07666(.A(new_n8042), .B(new_n8040), .Y(new_n8043));
  xor_4  g07667(.A(new_n8043), .B(new_n8039), .Y(new_n8044));
  and_6  g07668(.A(new_n7939), .B(new_n7938), .Y(new_n8045));
  nor_5  g07669(.A(new_n7943), .B(new_n7940), .Y(new_n8046));
  nor_5  g07670(.A(new_n8046), .B(new_n8045), .Y(new_n8047));
  xor_4  g07671(.A(new_n8047), .B(new_n8044), .Y(new_n8048));
  xor_4  g07672(.A(new_n8048), .B(new_n8036), .Y(new_n8049));
  xor_4  g07673(.A(new_n8049), .B(new_n8031), .Y(new_n8050));
  xor_4  g07674(.A(new_n8050), .B(new_n8026), .Y(new_n8051));
  xor_4  g07675(.A(new_n8051), .B(new_n7979), .Y(po039));
  xor_4  g07676(.A(new_n7934), .B(new_n7927), .Y(po040));
  nand_5 g07677(.A(pi117), .B(pi069), .Y(new_n8054));
  not_8  g07678(.A(new_n5033), .Y(new_n8055));
  nor_5  g07679(.A(new_n8054), .B(new_n8055), .Y(new_n8056));
  nand_5 g07680(.A(pi244), .B(pi103), .Y(new_n8057));
  nand_5 g07681(.A(pi029), .B(pi016), .Y(new_n8058));
  or_6   g07682(.A(new_n8058), .B(new_n8057), .Y(new_n8059));
  nand_5 g07683(.A(new_n8058), .B(new_n8057), .Y(new_n8060));
  and_6  g07684(.A(new_n8060), .B(new_n8059), .Y(new_n8061));
  or_6   g07685(.A(new_n8061), .B(new_n8056), .Y(new_n8062));
  nor_5  g07686(.A(new_n8062), .B(new_n8054), .Y(new_n8063));
  nand_5 g07687(.A(pi150), .B(pi103), .Y(new_n8064));
  nand_5 g07688(.A(new_n8059), .B(new_n8054), .Y(new_n8065));
  nand_5 g07689(.A(new_n8065), .B(new_n8060), .Y(new_n8066));
  xor_4  g07690(.A(new_n8066), .B(new_n8064), .Y(new_n8067));
  nand_5 g07691(.A(pi069), .B(pi016), .Y(new_n8068));
  nand_5 g07692(.A(pi080), .B(pi029), .Y(new_n8069));
  nand_5 g07693(.A(pi244), .B(pi117), .Y(new_n8070));
  xor_4  g07694(.A(new_n8070), .B(new_n8069), .Y(new_n8071));
  xor_4  g07695(.A(new_n8071), .B(new_n8068), .Y(new_n8072));
  xor_4  g07696(.A(new_n8072), .B(new_n8067), .Y(new_n8073));
  not_8  g07697(.A(new_n8073), .Y(new_n8074));
  nand_5 g07698(.A(new_n8074), .B(new_n8063), .Y(new_n8075));
  nand_5 g07699(.A(pi244), .B(pi016), .Y(new_n8076));
  nand_5 g07700(.A(pi247), .B(pi029), .Y(new_n8077));
  nand_5 g07701(.A(pi080), .B(pi069), .Y(new_n8078));
  xor_4  g07702(.A(new_n8078), .B(new_n8077), .Y(new_n8079));
  xor_4  g07703(.A(new_n8079), .B(new_n8076), .Y(new_n8080));
  nand_5 g07704(.A(pi150), .B(pi117), .Y(new_n8081));
  nand_5 g07705(.A(new_n8070), .B(new_n8069), .Y(new_n8082));
  nand_5 g07706(.A(new_n8071), .B(new_n8068), .Y(new_n8083));
  nand_5 g07707(.A(new_n8083), .B(new_n8082), .Y(new_n8084));
  xor_4  g07708(.A(new_n8084), .B(new_n8081), .Y(new_n8085));
  xor_4  g07709(.A(new_n8085), .B(new_n8080), .Y(new_n8086));
  nand_5 g07710(.A(pi221), .B(pi103), .Y(new_n8087));
  nor_5  g07711(.A(new_n8066), .B(new_n8064), .Y(new_n8088));
  not_8  g07712(.A(new_n8072), .Y(new_n8089));
  nand_5 g07713(.A(new_n8089), .B(new_n8067), .Y(new_n8090));
  not_8  g07714(.A(new_n8090), .Y(new_n8091));
  nor_5  g07715(.A(new_n8091), .B(new_n8088), .Y(new_n8092));
  xor_4  g07716(.A(new_n8092), .B(new_n8087), .Y(new_n8093));
  xor_4  g07717(.A(new_n8093), .B(new_n8086), .Y(new_n8094));
  xor_4  g07718(.A(new_n8094), .B(new_n8075), .Y(new_n8095));
  nand_5 g07719(.A(new_n8056), .B(new_n8060), .Y(new_n8096));
  nand_5 g07720(.A(new_n8096), .B(new_n8062), .Y(new_n8097));
  nand_5 g07721(.A(new_n5042), .B(new_n5039), .Y(new_n8098));
  nand_5 g07722(.A(new_n5069), .B(new_n5043), .Y(new_n8099));
  and_6  g07723(.A(new_n8099), .B(new_n8098), .Y(new_n8100));
  or_6   g07724(.A(new_n8100), .B(new_n8097), .Y(new_n8101));
  nand_5 g07725(.A(new_n5051), .B(new_n5045), .Y(new_n8102));
  nand_5 g07726(.A(new_n5067), .B(new_n5052), .Y(new_n8103));
  nand_5 g07727(.A(new_n8103), .B(new_n8102), .Y(new_n8104));
  nand_5 g07728(.A(pi240), .B(pi132), .Y(new_n8105));
  nand_5 g07729(.A(pi175), .B(pi058), .Y(new_n8106));
  xor_4  g07730(.A(new_n8106), .B(new_n5046), .Y(new_n8107));
  xor_4  g07731(.A(new_n8107), .B(new_n8105), .Y(new_n8108));
  xor_4  g07732(.A(new_n8108), .B(new_n5047), .Y(new_n8109));
  xor_4  g07733(.A(new_n8109), .B(new_n8104), .Y(new_n8110));
  nand_5 g07734(.A(pi109), .B(pi049), .Y(new_n8111));
  nand_5 g07735(.A(pi173), .B(pi107), .Y(new_n8112));
  xor_4  g07736(.A(new_n8112), .B(new_n5053), .Y(new_n8113));
  xor_4  g07737(.A(new_n8113), .B(new_n8111), .Y(new_n8114));
  xnor_4 g07738(.A(new_n8114), .B(new_n5054), .Y(new_n8115));
  nor_5  g07739(.A(new_n5065), .B(new_n5059), .Y(new_n8116));
  nor_5  g07740(.A(new_n5066), .B(new_n5058), .Y(new_n8117));
  nor_5  g07741(.A(new_n8117), .B(new_n8116), .Y(new_n8118));
  xnor_4 g07742(.A(new_n8118), .B(new_n8115), .Y(new_n8119));
  nand_5 g07743(.A(pi163), .B(pi066), .Y(new_n8120));
  xor_4  g07744(.A(new_n8120), .B(new_n5060), .Y(new_n8121));
  nand_5 g07745(.A(pi228), .B(pi226), .Y(new_n8122));
  xor_4  g07746(.A(new_n8122), .B(new_n8121), .Y(new_n8123));
  xor_4  g07747(.A(new_n8123), .B(new_n5061), .Y(new_n8124));
  xnor_4 g07748(.A(new_n8124), .B(new_n8119), .Y(new_n8125));
  xor_4  g07749(.A(new_n8125), .B(new_n8110), .Y(new_n8126));
  xor_4  g07750(.A(new_n8100), .B(new_n8097), .Y(new_n8127));
  nand_5 g07751(.A(new_n8127), .B(new_n8126), .Y(new_n8128));
  nand_5 g07752(.A(new_n8128), .B(new_n8101), .Y(new_n8129));
  xor_4  g07753(.A(new_n8073), .B(new_n8063), .Y(new_n8130));
  not_8  g07754(.A(new_n8130), .Y(new_n8131));
  nor_5  g07755(.A(new_n8131), .B(new_n8129), .Y(new_n8132));
  xor_4  g07756(.A(new_n8130), .B(new_n8129), .Y(new_n8133));
  nor_5  g07757(.A(new_n8109), .B(new_n8104), .Y(new_n8134));
  nand_5 g07758(.A(new_n8125), .B(new_n8110), .Y(new_n8135));
  not_8  g07759(.A(new_n8135), .Y(new_n8136));
  nor_5  g07760(.A(new_n8136), .B(new_n8134), .Y(new_n8137));
  not_8  g07761(.A(new_n8108), .Y(new_n8138));
  nand_5 g07762(.A(new_n8138), .B(new_n5047), .Y(new_n8139));
  nand_5 g07763(.A(pi134), .B(pi058), .Y(new_n8140));
  nand_5 g07764(.A(pi149), .B(pi132), .Y(new_n8141));
  nand_5 g07765(.A(pi240), .B(pi186), .Y(new_n8142));
  xor_4  g07766(.A(new_n8142), .B(new_n8141), .Y(new_n8143));
  xor_4  g07767(.A(new_n8143), .B(new_n8140), .Y(new_n8144));
  nand_5 g07768(.A(pi211), .B(pi175), .Y(new_n8145));
  nand_5 g07769(.A(new_n8106), .B(new_n5046), .Y(new_n8146));
  nand_5 g07770(.A(new_n8107), .B(new_n8105), .Y(new_n8147));
  nand_5 g07771(.A(new_n8147), .B(new_n8146), .Y(new_n8148));
  xor_4  g07772(.A(new_n8148), .B(new_n8145), .Y(new_n8149));
  xor_4  g07773(.A(new_n8149), .B(new_n8144), .Y(new_n8150));
  xor_4  g07774(.A(new_n8150), .B(new_n8139), .Y(new_n8151));
  and_6  g07775(.A(new_n8118), .B(new_n8115), .Y(new_n8152));
  nor_5  g07776(.A(new_n8124), .B(new_n8119), .Y(new_n8153));
  nor_5  g07777(.A(new_n8153), .B(new_n8152), .Y(new_n8154));
  nor_5  g07778(.A(new_n8123), .B(new_n5061), .Y(new_n8155));
  nand_5 g07779(.A(pi228), .B(pi207), .Y(new_n8156));
  nand_5 g07780(.A(pi148), .B(pi066), .Y(new_n8157));
  nand_5 g07781(.A(pi226), .B(pi039), .Y(new_n8158));
  xor_4  g07782(.A(new_n8158), .B(new_n8157), .Y(new_n8159));
  xor_4  g07783(.A(new_n8159), .B(new_n8156), .Y(new_n8160));
  nand_5 g07784(.A(pi163), .B(pi055), .Y(new_n8161));
  nand_5 g07785(.A(new_n8120), .B(new_n5060), .Y(new_n8162));
  nand_5 g07786(.A(new_n8122), .B(new_n8121), .Y(new_n8163));
  nand_5 g07787(.A(new_n8163), .B(new_n8162), .Y(new_n8164));
  xor_4  g07788(.A(new_n8164), .B(new_n8161), .Y(new_n8165));
  xnor_4 g07789(.A(new_n8165), .B(new_n8160), .Y(new_n8166));
  xnor_4 g07790(.A(new_n8166), .B(new_n8155), .Y(new_n8167));
  nor_5  g07791(.A(new_n8114), .B(new_n5054), .Y(new_n8168));
  nand_5 g07792(.A(pi173), .B(pi171), .Y(new_n8169));
  nand_5 g07793(.A(pi245), .B(pi109), .Y(new_n8170));
  nand_5 g07794(.A(pi049), .B(pi014), .Y(new_n8171));
  xor_4  g07795(.A(new_n8171), .B(new_n8170), .Y(new_n8172));
  xor_4  g07796(.A(new_n8172), .B(new_n8169), .Y(new_n8173));
  nand_5 g07797(.A(pi230), .B(pi107), .Y(new_n8174));
  nand_5 g07798(.A(new_n8112), .B(new_n5053), .Y(new_n8175));
  nand_5 g07799(.A(new_n8113), .B(new_n8111), .Y(new_n8176));
  nand_5 g07800(.A(new_n8176), .B(new_n8175), .Y(new_n8177));
  xor_4  g07801(.A(new_n8177), .B(new_n8174), .Y(new_n8178));
  xnor_4 g07802(.A(new_n8178), .B(new_n8173), .Y(new_n8179));
  xnor_4 g07803(.A(new_n8179), .B(new_n8168), .Y(new_n8180));
  nand_5 g07804(.A(new_n8180), .B(new_n8167), .Y(new_n8181));
  not_8  g07805(.A(new_n8181), .Y(new_n8182));
  nor_5  g07806(.A(new_n8180), .B(new_n8167), .Y(new_n8183));
  nor_5  g07807(.A(new_n8183), .B(new_n8182), .Y(new_n8184));
  xor_4  g07808(.A(new_n8184), .B(new_n8154), .Y(new_n8185));
  xnor_4 g07809(.A(new_n8185), .B(new_n8151), .Y(new_n8186));
  xor_4  g07810(.A(new_n8186), .B(new_n8137), .Y(new_n8187));
  nor_5  g07811(.A(new_n8187), .B(new_n8133), .Y(new_n8188));
  nor_5  g07812(.A(new_n8188), .B(new_n8132), .Y(new_n8189));
  xnor_4 g07813(.A(new_n8189), .B(new_n8095), .Y(new_n8190));
  nand_5 g07814(.A(new_n8185), .B(new_n8151), .Y(new_n8191));
  or_6   g07815(.A(new_n8186), .B(new_n8137), .Y(new_n8192));
  and_6  g07816(.A(new_n8192), .B(new_n8191), .Y(new_n8193));
  nor_5  g07817(.A(new_n8150), .B(new_n8139), .Y(new_n8194));
  nand_5 g07818(.A(pi199), .B(pi175), .Y(new_n8195));
  nor_5  g07819(.A(new_n8148), .B(new_n8145), .Y(new_n8196));
  not_8  g07820(.A(new_n8149), .Y(new_n8197));
  nor_5  g07821(.A(new_n8197), .B(new_n8144), .Y(new_n8198));
  nor_5  g07822(.A(new_n8198), .B(new_n8196), .Y(new_n8199));
  xor_4  g07823(.A(new_n8199), .B(new_n8195), .Y(new_n8200));
  nand_5 g07824(.A(pi240), .B(pi058), .Y(new_n8201));
  nand_5 g07825(.A(pi186), .B(pi149), .Y(new_n8202));
  nand_5 g07826(.A(pi167), .B(pi132), .Y(new_n8203));
  xor_4  g07827(.A(new_n8203), .B(new_n8202), .Y(new_n8204));
  xor_4  g07828(.A(new_n8204), .B(new_n8201), .Y(new_n8205));
  nand_5 g07829(.A(pi211), .B(pi134), .Y(new_n8206));
  nand_5 g07830(.A(new_n8142), .B(new_n8141), .Y(new_n8207));
  nand_5 g07831(.A(new_n8143), .B(new_n8140), .Y(new_n8208));
  nand_5 g07832(.A(new_n8208), .B(new_n8207), .Y(new_n8209));
  xor_4  g07833(.A(new_n8209), .B(new_n8206), .Y(new_n8210));
  xnor_4 g07834(.A(new_n8210), .B(new_n8205), .Y(new_n8211));
  xor_4  g07835(.A(new_n8211), .B(new_n8200), .Y(new_n8212));
  xor_4  g07836(.A(new_n8212), .B(new_n8194), .Y(new_n8213));
  or_6   g07837(.A(new_n8183), .B(new_n8154), .Y(new_n8214));
  nand_5 g07838(.A(new_n8214), .B(new_n8181), .Y(new_n8215));
  nand_5 g07839(.A(new_n8166), .B(new_n8155), .Y(new_n8216));
  nand_5 g07840(.A(pi226), .B(pi116), .Y(new_n8217));
  nand_5 g07841(.A(pi228), .B(pi066), .Y(new_n8218));
  nand_5 g07842(.A(pi207), .B(pi039), .Y(new_n8219));
  xor_4  g07843(.A(new_n8219), .B(new_n8218), .Y(new_n8220));
  xor_4  g07844(.A(new_n8220), .B(new_n8217), .Y(new_n8221));
  nand_5 g07845(.A(pi148), .B(pi055), .Y(new_n8222));
  nand_5 g07846(.A(new_n8158), .B(new_n8157), .Y(new_n8223));
  nand_5 g07847(.A(new_n8159), .B(new_n8156), .Y(new_n8224));
  nand_5 g07848(.A(new_n8224), .B(new_n8223), .Y(new_n8225));
  xor_4  g07849(.A(new_n8225), .B(new_n8222), .Y(new_n8226));
  xor_4  g07850(.A(new_n8226), .B(new_n8221), .Y(new_n8227));
  nand_5 g07851(.A(pi163), .B(pi002), .Y(new_n8228));
  nand_5 g07852(.A(new_n8164), .B(new_n8161), .Y(new_n8229));
  nand_5 g07853(.A(new_n8165), .B(new_n8160), .Y(new_n8230));
  nand_5 g07854(.A(new_n8230), .B(new_n8229), .Y(new_n8231));
  xnor_4 g07855(.A(new_n8231), .B(new_n8228), .Y(new_n8232));
  xnor_4 g07856(.A(new_n8232), .B(new_n8227), .Y(new_n8233));
  xor_4  g07857(.A(new_n8233), .B(new_n8216), .Y(new_n8234));
  nand_5 g07858(.A(new_n8179), .B(new_n8168), .Y(new_n8235));
  nand_5 g07859(.A(pi173), .B(pi049), .Y(new_n8236));
  nand_5 g07860(.A(pi245), .B(pi014), .Y(new_n8237));
  nand_5 g07861(.A(pi201), .B(pi109), .Y(new_n8238));
  xor_4  g07862(.A(new_n8238), .B(new_n8237), .Y(new_n8239));
  xor_4  g07863(.A(new_n8239), .B(new_n8236), .Y(new_n8240));
  nand_5 g07864(.A(pi230), .B(pi171), .Y(new_n8241));
  nand_5 g07865(.A(new_n8171), .B(new_n8170), .Y(new_n8242));
  nand_5 g07866(.A(new_n8172), .B(new_n8169), .Y(new_n8243));
  nand_5 g07867(.A(new_n8243), .B(new_n8242), .Y(new_n8244));
  xor_4  g07868(.A(new_n8244), .B(new_n8241), .Y(new_n8245));
  xor_4  g07869(.A(new_n8245), .B(new_n8240), .Y(new_n8246));
  nand_5 g07870(.A(pi107), .B(pi050), .Y(new_n8247));
  nand_5 g07871(.A(new_n8177), .B(new_n8174), .Y(new_n8248));
  nand_5 g07872(.A(new_n8178), .B(new_n8173), .Y(new_n8249));
  nand_5 g07873(.A(new_n8249), .B(new_n8248), .Y(new_n8250));
  xnor_4 g07874(.A(new_n8250), .B(new_n8247), .Y(new_n8251));
  xnor_4 g07875(.A(new_n8251), .B(new_n8246), .Y(new_n8252));
  xor_4  g07876(.A(new_n8252), .B(new_n8235), .Y(new_n8253));
  nand_5 g07877(.A(new_n8253), .B(new_n8234), .Y(new_n8254));
  nor_5  g07878(.A(new_n8253), .B(new_n8234), .Y(new_n8255));
  not_8  g07879(.A(new_n8255), .Y(new_n8256));
  nand_5 g07880(.A(new_n8256), .B(new_n8254), .Y(new_n8257));
  xor_4  g07881(.A(new_n8257), .B(new_n8215), .Y(new_n8258));
  xnor_4 g07882(.A(new_n8258), .B(new_n8213), .Y(new_n8259));
  xor_4  g07883(.A(new_n8259), .B(new_n8193), .Y(new_n8260));
  xnor_4 g07884(.A(new_n8260), .B(new_n8190), .Y(po041));
  xor_4  g07885(.A(new_n7061), .B(new_n7060), .Y(po042));
  xnor_4 g07886(.A(new_n5014), .B(new_n5013), .Y(po043));
  xor_4  g07887(.A(new_n1034), .B(new_n1018), .Y(po044));
  xor_4  g07888(.A(new_n2587), .B(new_n2554), .Y(po045));
  xor_4  g07889(.A(new_n5000), .B(new_n4995), .Y(po046));
  nand_5 g07890(.A(pi175), .B(pi037), .Y(new_n8267));
  nand_5 g07891(.A(pi200), .B(pi186), .Y(new_n8268));
  xor_4  g07892(.A(new_n8268), .B(new_n8267), .Y(new_n8269));
  nand_5 g07893(.A(pi207), .B(pi115), .Y(new_n8270));
  xor_4  g07894(.A(new_n8270), .B(new_n8269), .Y(new_n8271));
  nand_5 g07895(.A(pi171), .B(pi074), .Y(new_n8272));
  nand_5 g07896(.A(pi244), .B(pi080), .Y(new_n8273));
  nand_5 g07897(.A(new_n8078), .B(new_n8077), .Y(new_n8274));
  nand_5 g07898(.A(new_n8079), .B(new_n8076), .Y(new_n8275));
  nand_5 g07899(.A(new_n8275), .B(new_n8274), .Y(new_n8276));
  nand_5 g07900(.A(new_n8276), .B(new_n8273), .Y(new_n8277));
  nand_5 g07901(.A(pi247), .B(pi069), .Y(new_n8278));
  nand_5 g07902(.A(pi234), .B(pi029), .Y(new_n8279));
  nand_5 g07903(.A(new_n8279), .B(new_n8278), .Y(new_n8280));
  nand_5 g07904(.A(pi234), .B(pi069), .Y(new_n8281));
  nor_5  g07905(.A(new_n8281), .B(new_n8077), .Y(new_n8282));
  not_8  g07906(.A(new_n8282), .Y(new_n8283));
  nand_5 g07907(.A(new_n8283), .B(new_n8280), .Y(new_n8284));
  xor_4  g07908(.A(new_n8276), .B(new_n8273), .Y(new_n8285));
  nand_5 g07909(.A(new_n8285), .B(new_n8284), .Y(new_n8286));
  nand_5 g07910(.A(new_n8286), .B(new_n8277), .Y(new_n8287));
  nand_5 g07911(.A(pi221), .B(pi016), .Y(new_n8288));
  nand_5 g07912(.A(pi196), .B(pi117), .Y(new_n8289));
  nand_5 g07913(.A(pi184), .B(pi103), .Y(new_n8290));
  xor_4  g07914(.A(new_n8290), .B(new_n8289), .Y(new_n8291));
  xor_4  g07915(.A(new_n8291), .B(new_n8288), .Y(new_n8292));
  nand_5 g07916(.A(new_n8292), .B(new_n8287), .Y(new_n8293));
  xor_4  g07917(.A(new_n8292), .B(new_n8287), .Y(new_n8294));
  nand_5 g07918(.A(pi150), .B(pi080), .Y(new_n8295));
  xor_4  g07919(.A(new_n8295), .B(new_n8282), .Y(new_n8296));
  nand_5 g07920(.A(pi247), .B(pi244), .Y(new_n8297));
  nand_5 g07921(.A(pi214), .B(pi029), .Y(new_n8298));
  xor_4  g07922(.A(new_n8298), .B(new_n8281), .Y(new_n8299));
  xor_4  g07923(.A(new_n8299), .B(new_n8297), .Y(new_n8300));
  xnor_4 g07924(.A(new_n8300), .B(new_n8296), .Y(new_n8301));
  nand_5 g07925(.A(new_n8301), .B(new_n8294), .Y(new_n8302));
  nand_5 g07926(.A(new_n8302), .B(new_n8293), .Y(new_n8303));
  nand_5 g07927(.A(pi218), .B(pi134), .Y(new_n8304));
  xor_4  g07928(.A(new_n8304), .B(new_n8303), .Y(new_n8305));
  xor_4  g07929(.A(new_n8305), .B(new_n8272), .Y(new_n8306));
  nand_5 g07930(.A(new_n8209), .B(new_n8206), .Y(new_n8307));
  nand_5 g07931(.A(new_n8210), .B(new_n8205), .Y(new_n8308));
  nand_5 g07932(.A(new_n8308), .B(new_n8307), .Y(new_n8309));
  nand_5 g07933(.A(pi240), .B(pi211), .Y(new_n8310));
  nand_5 g07934(.A(pi199), .B(pi134), .Y(new_n8311));
  and_6  g07935(.A(new_n8311), .B(new_n8310), .Y(new_n8312));
  nand_5 g07936(.A(pi240), .B(pi199), .Y(new_n8313));
  nor_5  g07937(.A(new_n8313), .B(new_n8206), .Y(new_n8314));
  or_6   g07938(.A(new_n8314), .B(new_n8312), .Y(new_n8315));
  nand_5 g07939(.A(pi186), .B(pi181), .Y(new_n8316));
  nor_5  g07940(.A(new_n8316), .B(new_n8203), .Y(new_n8317));
  not_8  g07941(.A(new_n8317), .Y(new_n8318));
  nand_5 g07942(.A(pi186), .B(pi167), .Y(new_n8319));
  nand_5 g07943(.A(pi181), .B(pi132), .Y(new_n8320));
  nand_5 g07944(.A(new_n8320), .B(new_n8319), .Y(new_n8321));
  nand_5 g07945(.A(new_n8321), .B(new_n8318), .Y(new_n8322));
  nand_5 g07946(.A(pi149), .B(pi058), .Y(new_n8323));
  nand_5 g07947(.A(new_n8203), .B(new_n8202), .Y(new_n8324));
  nand_5 g07948(.A(new_n8204), .B(new_n8201), .Y(new_n8325));
  nand_5 g07949(.A(new_n8325), .B(new_n8324), .Y(new_n8326));
  xor_4  g07950(.A(new_n8326), .B(new_n8323), .Y(new_n8327));
  xor_4  g07951(.A(new_n8327), .B(new_n8322), .Y(new_n8328));
  xor_4  g07952(.A(new_n8328), .B(new_n8315), .Y(new_n8329));
  not_8  g07953(.A(new_n8329), .Y(new_n8330));
  xor_4  g07954(.A(new_n8330), .B(new_n8309), .Y(new_n8331));
  not_8  g07955(.A(new_n8331), .Y(new_n8332));
  nor_5  g07956(.A(new_n8199), .B(new_n8195), .Y(new_n8333));
  nand_5 g07957(.A(new_n8211), .B(new_n8200), .Y(new_n8334));
  not_8  g07958(.A(new_n8334), .Y(new_n8335));
  nor_5  g07959(.A(new_n8335), .B(new_n8333), .Y(new_n8336));
  nor_5  g07960(.A(new_n8336), .B(new_n8332), .Y(new_n8337));
  nor_5  g07961(.A(new_n8328), .B(new_n8315), .Y(new_n8338));
  nor_5  g07962(.A(new_n8330), .B(new_n8309), .Y(new_n8339));
  xor_4  g07963(.A(new_n8339), .B(new_n8314), .Y(new_n8340));
  nor_5  g07964(.A(new_n8340), .B(new_n8338), .Y(new_n8341));
  nand_5 g07965(.A(pi211), .B(pi149), .Y(new_n8342));
  xor_4  g07966(.A(new_n8342), .B(new_n8317), .Y(new_n8343));
  nand_5 g07967(.A(pi200), .B(pi132), .Y(new_n8344));
  nand_5 g07968(.A(pi167), .B(pi058), .Y(new_n8345));
  xor_4  g07969(.A(new_n8345), .B(new_n8344), .Y(new_n8346));
  xor_4  g07970(.A(new_n8346), .B(new_n8316), .Y(new_n8347));
  xor_4  g07971(.A(new_n8347), .B(new_n8343), .Y(new_n8348));
  nand_5 g07972(.A(new_n8326), .B(new_n8323), .Y(new_n8349));
  nand_5 g07973(.A(new_n8327), .B(new_n8322), .Y(new_n8350));
  nand_5 g07974(.A(new_n8350), .B(new_n8349), .Y(new_n8351));
  nand_5 g07975(.A(pi195), .B(pi134), .Y(new_n8352));
  nand_5 g07976(.A(pi218), .B(pi175), .Y(new_n8353));
  xor_4  g07977(.A(new_n8353), .B(new_n8352), .Y(new_n8354));
  xor_4  g07978(.A(new_n8354), .B(new_n8313), .Y(new_n8355));
  xor_4  g07979(.A(new_n8355), .B(new_n8351), .Y(new_n8356));
  not_8  g07980(.A(new_n8356), .Y(new_n8357));
  xor_4  g07981(.A(new_n8357), .B(new_n8348), .Y(new_n8358));
  xor_4  g07982(.A(new_n8358), .B(new_n8341), .Y(new_n8359));
  or_6   g07983(.A(new_n8359), .B(new_n8337), .Y(new_n8360));
  nand_5 g07984(.A(new_n8212), .B(new_n8194), .Y(new_n8361));
  nand_5 g07985(.A(pi195), .B(pi175), .Y(new_n8362));
  nand_5 g07986(.A(new_n8362), .B(new_n8361), .Y(new_n8363));
  xor_4  g07987(.A(new_n8336), .B(new_n8331), .Y(new_n8364));
  xor_4  g07988(.A(new_n8362), .B(new_n8361), .Y(new_n8365));
  nand_5 g07989(.A(new_n8365), .B(new_n8364), .Y(new_n8366));
  nand_5 g07990(.A(new_n8366), .B(new_n8363), .Y(new_n8367));
  xor_4  g07991(.A(new_n8359), .B(new_n8337), .Y(new_n8368));
  nand_5 g07992(.A(new_n8368), .B(new_n8367), .Y(new_n8369));
  nand_5 g07993(.A(new_n8369), .B(new_n8360), .Y(new_n8370));
  nand_5 g07994(.A(pi253), .B(pi049), .Y(new_n8371));
  nand_5 g07995(.A(pi103), .B(pi010), .Y(new_n8372));
  xor_4  g07996(.A(new_n8372), .B(new_n8371), .Y(new_n8373));
  xor_4  g07997(.A(new_n8373), .B(new_n8370), .Y(new_n8374));
  xor_4  g07998(.A(new_n8374), .B(new_n8306), .Y(new_n8375));
  xor_4  g07999(.A(new_n8375), .B(new_n8271), .Y(new_n8376));
  nand_5 g08000(.A(new_n8258), .B(new_n8213), .Y(new_n8377));
  or_6   g08001(.A(new_n8259), .B(new_n8193), .Y(new_n8378));
  nand_5 g08002(.A(new_n8378), .B(new_n8377), .Y(new_n8379));
  xnor_4 g08003(.A(new_n8365), .B(new_n8364), .Y(new_n8380));
  nand_5 g08004(.A(new_n8380), .B(new_n8379), .Y(new_n8381));
  or_6   g08005(.A(new_n8250), .B(new_n8247), .Y(new_n8382));
  or_6   g08006(.A(new_n8251), .B(new_n8246), .Y(new_n8383));
  and_6  g08007(.A(new_n8383), .B(new_n8382), .Y(new_n8384));
  nand_5 g08008(.A(pi050), .B(pi049), .Y(new_n8385));
  nor_5  g08009(.A(new_n8385), .B(new_n8241), .Y(new_n8386));
  nand_5 g08010(.A(pi230), .B(pi049), .Y(new_n8387));
  nand_5 g08011(.A(pi171), .B(pi050), .Y(new_n8388));
  and_6  g08012(.A(new_n8388), .B(new_n8387), .Y(new_n8389));
  or_6   g08013(.A(new_n8389), .B(new_n8386), .Y(new_n8390));
  nand_5 g08014(.A(new_n8238), .B(new_n8237), .Y(new_n8391));
  nand_5 g08015(.A(new_n8239), .B(new_n8236), .Y(new_n8392));
  nand_5 g08016(.A(new_n8392), .B(new_n8391), .Y(new_n8393));
  nand_5 g08017(.A(pi245), .B(pi173), .Y(new_n8394));
  nand_5 g08018(.A(pi201), .B(pi014), .Y(new_n8395));
  nand_5 g08019(.A(pi156), .B(pi109), .Y(new_n8396));
  nand_5 g08020(.A(new_n8396), .B(new_n8395), .Y(new_n8397));
  nand_5 g08021(.A(pi156), .B(pi014), .Y(new_n8398));
  nor_5  g08022(.A(new_n8398), .B(new_n8238), .Y(new_n8399));
  not_8  g08023(.A(new_n8399), .Y(new_n8400));
  nand_5 g08024(.A(new_n8400), .B(new_n8397), .Y(new_n8401));
  xor_4  g08025(.A(new_n8401), .B(new_n8394), .Y(new_n8402));
  xor_4  g08026(.A(new_n8402), .B(new_n8393), .Y(new_n8403));
  xnor_4 g08027(.A(new_n8403), .B(new_n8390), .Y(new_n8404));
  nand_5 g08028(.A(new_n8244), .B(new_n8241), .Y(new_n8405));
  nand_5 g08029(.A(new_n8245), .B(new_n8240), .Y(new_n8406));
  nand_5 g08030(.A(new_n8406), .B(new_n8405), .Y(new_n8407));
  xnor_4 g08031(.A(new_n8407), .B(new_n8404), .Y(new_n8408));
  xnor_4 g08032(.A(new_n8408), .B(new_n8384), .Y(new_n8409));
  or_6   g08033(.A(new_n8252), .B(new_n8235), .Y(new_n8410));
  nand_5 g08034(.A(pi253), .B(pi107), .Y(new_n8411));
  xor_4  g08035(.A(new_n8411), .B(new_n8410), .Y(new_n8412));
  xor_4  g08036(.A(new_n8412), .B(new_n8409), .Y(new_n8413));
  or_6   g08037(.A(new_n8233), .B(new_n8216), .Y(new_n8414));
  nand_5 g08038(.A(pi163), .B(pi025), .Y(new_n8415));
  xor_4  g08039(.A(new_n8415), .B(new_n8414), .Y(new_n8416));
  nand_5 g08040(.A(new_n8225), .B(new_n8222), .Y(new_n8417));
  nand_5 g08041(.A(new_n8226), .B(new_n8221), .Y(new_n8418));
  nand_5 g08042(.A(new_n8418), .B(new_n8417), .Y(new_n8419));
  nand_5 g08043(.A(pi228), .B(pi055), .Y(new_n8420));
  nand_5 g08044(.A(pi148), .B(pi002), .Y(new_n8421));
  nand_5 g08045(.A(new_n8421), .B(new_n8420), .Y(new_n8422));
  nand_5 g08046(.A(pi228), .B(pi002), .Y(new_n8423));
  or_6   g08047(.A(new_n8423), .B(new_n8222), .Y(new_n8424));
  nand_5 g08048(.A(new_n8424), .B(new_n8422), .Y(new_n8425));
  xor_4  g08049(.A(new_n8425), .B(new_n8419), .Y(new_n8426));
  nand_5 g08050(.A(new_n8219), .B(new_n8218), .Y(new_n8427));
  nand_5 g08051(.A(new_n8220), .B(new_n8217), .Y(new_n8428));
  nand_5 g08052(.A(new_n8428), .B(new_n8427), .Y(new_n8429));
  nand_5 g08053(.A(pi066), .B(pi039), .Y(new_n8430));
  nand_5 g08054(.A(pi207), .B(pi070), .Y(new_n8431));
  nor_5  g08055(.A(new_n8431), .B(new_n8217), .Y(new_n8432));
  not_8  g08056(.A(new_n8432), .Y(new_n8433));
  nand_5 g08057(.A(pi207), .B(pi116), .Y(new_n8434));
  nand_5 g08058(.A(pi226), .B(pi070), .Y(new_n8435));
  nand_5 g08059(.A(new_n8435), .B(new_n8434), .Y(new_n8436));
  nand_5 g08060(.A(new_n8436), .B(new_n8433), .Y(new_n8437));
  xor_4  g08061(.A(new_n8437), .B(new_n8430), .Y(new_n8438));
  xor_4  g08062(.A(new_n8438), .B(new_n8429), .Y(new_n8439));
  xnor_4 g08063(.A(new_n8439), .B(new_n8426), .Y(new_n8440));
  nor_5  g08064(.A(new_n8231), .B(new_n8228), .Y(new_n8441));
  nor_5  g08065(.A(new_n8232), .B(new_n8227), .Y(new_n8442));
  nor_5  g08066(.A(new_n8442), .B(new_n8441), .Y(new_n8443));
  xor_4  g08067(.A(new_n8443), .B(new_n8440), .Y(new_n8444));
  xnor_4 g08068(.A(new_n8444), .B(new_n8416), .Y(new_n8445));
  nand_5 g08069(.A(new_n8254), .B(new_n8215), .Y(new_n8446));
  and_6  g08070(.A(new_n8446), .B(new_n8256), .Y(new_n8447));
  xnor_4 g08071(.A(new_n8447), .B(new_n8445), .Y(new_n8448));
  xor_4  g08072(.A(new_n8448), .B(new_n8413), .Y(new_n8449));
  xor_4  g08073(.A(new_n8380), .B(new_n8379), .Y(new_n8450));
  nand_5 g08074(.A(new_n8450), .B(new_n8449), .Y(new_n8451));
  nand_5 g08075(.A(new_n8451), .B(new_n8381), .Y(new_n8452));
  nand_5 g08076(.A(new_n8411), .B(new_n8410), .Y(new_n8453));
  nand_5 g08077(.A(new_n8412), .B(new_n8409), .Y(new_n8454));
  nand_5 g08078(.A(new_n8454), .B(new_n8453), .Y(new_n8455));
  or_6   g08079(.A(new_n8408), .B(new_n8384), .Y(new_n8456));
  nand_5 g08080(.A(pi245), .B(pi230), .Y(new_n8457));
  xor_4  g08081(.A(new_n8457), .B(new_n8400), .Y(new_n8458));
  nand_5 g08082(.A(pi109), .B(pi063), .Y(new_n8459));
  nand_5 g08083(.A(pi201), .B(pi173), .Y(new_n8460));
  xor_4  g08084(.A(new_n8460), .B(new_n8459), .Y(new_n8461));
  xor_4  g08085(.A(new_n8461), .B(new_n8398), .Y(new_n8462));
  not_8  g08086(.A(new_n8462), .Y(new_n8463));
  xor_4  g08087(.A(new_n8463), .B(new_n8458), .Y(new_n8464));
  nand_5 g08088(.A(new_n8401), .B(new_n8394), .Y(new_n8465));
  nand_5 g08089(.A(new_n8402), .B(new_n8393), .Y(new_n8466));
  nand_5 g08090(.A(new_n8466), .B(new_n8465), .Y(new_n8467));
  nand_5 g08091(.A(pi253), .B(pi171), .Y(new_n8468));
  nand_5 g08092(.A(pi107), .B(pi074), .Y(new_n8469));
  xor_4  g08093(.A(new_n8469), .B(new_n8468), .Y(new_n8470));
  xnor_4 g08094(.A(new_n8470), .B(new_n8385), .Y(new_n8471));
  xor_4  g08095(.A(new_n8471), .B(new_n8467), .Y(new_n8472));
  xor_4  g08096(.A(new_n8472), .B(new_n8464), .Y(new_n8473));
  nor_5  g08097(.A(new_n8403), .B(new_n8390), .Y(new_n8474));
  nor_5  g08098(.A(new_n8407), .B(new_n8404), .Y(new_n8475));
  xor_4  g08099(.A(new_n8475), .B(new_n8386), .Y(new_n8476));
  nor_5  g08100(.A(new_n8476), .B(new_n8474), .Y(new_n8477));
  xor_4  g08101(.A(new_n8477), .B(new_n8473), .Y(new_n8478));
  xor_4  g08102(.A(new_n8478), .B(new_n8456), .Y(new_n8479));
  xor_4  g08103(.A(new_n8479), .B(new_n8455), .Y(new_n8480));
  nand_5 g08104(.A(new_n8415), .B(new_n8414), .Y(new_n8481));
  nand_5 g08105(.A(new_n8444), .B(new_n8416), .Y(new_n8482));
  nand_5 g08106(.A(new_n8482), .B(new_n8481), .Y(new_n8483));
  not_8  g08107(.A(new_n8440), .Y(new_n8484));
  or_6   g08108(.A(new_n8443), .B(new_n8484), .Y(new_n8485));
  nand_5 g08109(.A(new_n8425), .B(new_n8419), .Y(new_n8486));
  nand_5 g08110(.A(new_n8439), .B(new_n8426), .Y(new_n8487));
  nand_5 g08111(.A(new_n8487), .B(new_n8486), .Y(new_n8488));
  xnor_4 g08112(.A(new_n8488), .B(new_n8424), .Y(new_n8489));
  nand_5 g08113(.A(pi055), .B(pi039), .Y(new_n8490));
  xor_4  g08114(.A(new_n8490), .B(new_n8432), .Y(new_n8491));
  nand_5 g08115(.A(pi226), .B(pi115), .Y(new_n8492));
  nand_5 g08116(.A(pi116), .B(pi066), .Y(new_n8493));
  xor_4  g08117(.A(new_n8493), .B(new_n8492), .Y(new_n8494));
  xor_4  g08118(.A(new_n8494), .B(new_n8431), .Y(new_n8495));
  xor_4  g08119(.A(new_n8495), .B(new_n8491), .Y(new_n8496));
  nand_5 g08120(.A(new_n8437), .B(new_n8430), .Y(new_n8497));
  nand_5 g08121(.A(new_n8438), .B(new_n8429), .Y(new_n8498));
  nand_5 g08122(.A(new_n8498), .B(new_n8497), .Y(new_n8499));
  nand_5 g08123(.A(pi239), .B(pi163), .Y(new_n8500));
  nand_5 g08124(.A(pi148), .B(pi025), .Y(new_n8501));
  xor_4  g08125(.A(new_n8501), .B(new_n8500), .Y(new_n8502));
  xor_4  g08126(.A(new_n8502), .B(new_n8423), .Y(new_n8503));
  xor_4  g08127(.A(new_n8503), .B(new_n8499), .Y(new_n8504));
  xor_4  g08128(.A(new_n8504), .B(new_n8496), .Y(new_n8505));
  not_8  g08129(.A(new_n8505), .Y(new_n8506));
  xor_4  g08130(.A(new_n8506), .B(new_n8489), .Y(new_n8507));
  xor_4  g08131(.A(new_n8507), .B(new_n8485), .Y(new_n8508));
  xor_4  g08132(.A(new_n8508), .B(new_n8483), .Y(new_n8509));
  xnor_4 g08133(.A(new_n8509), .B(new_n8480), .Y(new_n8510));
  nand_5 g08134(.A(new_n8447), .B(new_n8445), .Y(new_n8511));
  or_6   g08135(.A(new_n8448), .B(new_n8413), .Y(new_n8512));
  nand_5 g08136(.A(new_n8512), .B(new_n8511), .Y(new_n8513));
  xor_4  g08137(.A(new_n8513), .B(new_n8510), .Y(new_n8514));
  not_8  g08138(.A(new_n8514), .Y(new_n8515));
  xor_4  g08139(.A(new_n8515), .B(new_n8452), .Y(new_n8516));
  xor_4  g08140(.A(new_n8368), .B(new_n8367), .Y(new_n8517));
  xor_4  g08141(.A(new_n8517), .B(new_n8516), .Y(new_n8518));
  nand_5 g08142(.A(new_n8092), .B(new_n8087), .Y(new_n8519));
  nand_5 g08143(.A(new_n8093), .B(new_n8086), .Y(new_n8520));
  nand_5 g08144(.A(new_n8520), .B(new_n8519), .Y(new_n8521));
  nand_5 g08145(.A(new_n8084), .B(new_n8081), .Y(new_n8522));
  nand_5 g08146(.A(new_n8085), .B(new_n8080), .Y(new_n8523));
  nand_5 g08147(.A(new_n8523), .B(new_n8522), .Y(new_n8524));
  nor_5  g08148(.A(new_n8288), .B(new_n8081), .Y(new_n8525));
  not_8  g08149(.A(new_n8525), .Y(new_n8526));
  nand_5 g08150(.A(pi150), .B(pi016), .Y(new_n8527));
  nand_5 g08151(.A(pi221), .B(pi117), .Y(new_n8528));
  nand_5 g08152(.A(new_n8528), .B(new_n8527), .Y(new_n8529));
  nand_5 g08153(.A(new_n8529), .B(new_n8526), .Y(new_n8530));
  xor_4  g08154(.A(new_n8285), .B(new_n8284), .Y(new_n8531));
  xor_4  g08155(.A(new_n8531), .B(new_n8530), .Y(new_n8532));
  xor_4  g08156(.A(new_n8532), .B(new_n8524), .Y(new_n8533));
  nor_5  g08157(.A(new_n8533), .B(new_n8521), .Y(new_n8534));
  xor_4  g08158(.A(new_n8301), .B(new_n8294), .Y(new_n8535));
  nand_5 g08159(.A(new_n8531), .B(new_n8530), .Y(new_n8536));
  nand_5 g08160(.A(new_n8532), .B(new_n8524), .Y(new_n8537));
  nand_5 g08161(.A(new_n8537), .B(new_n8536), .Y(new_n8538));
  xor_4  g08162(.A(new_n8538), .B(new_n8525), .Y(new_n8539));
  xor_4  g08163(.A(new_n8539), .B(new_n8535), .Y(new_n8540));
  xor_4  g08164(.A(new_n8540), .B(new_n8534), .Y(new_n8541));
  nand_5 g08165(.A(pi196), .B(pi103), .Y(new_n8542));
  xnor_4 g08166(.A(new_n8533), .B(new_n8521), .Y(new_n8543));
  nor_5  g08167(.A(new_n8543), .B(new_n8542), .Y(new_n8544));
  not_8  g08168(.A(new_n8544), .Y(new_n8545));
  not_8  g08169(.A(new_n8075), .Y(new_n8546));
  not_8  g08170(.A(new_n8094), .Y(new_n8547));
  nand_5 g08171(.A(new_n8547), .B(new_n8546), .Y(new_n8548));
  not_8  g08172(.A(new_n8548), .Y(new_n8549));
  xor_4  g08173(.A(new_n8543), .B(new_n8542), .Y(new_n8550));
  nand_5 g08174(.A(new_n8550), .B(new_n8549), .Y(new_n8551));
  nand_5 g08175(.A(new_n8551), .B(new_n8545), .Y(new_n8552));
  xor_4  g08176(.A(new_n8552), .B(new_n8541), .Y(new_n8553));
  not_8  g08177(.A(new_n8553), .Y(new_n8554));
  or_6   g08178(.A(new_n8554), .B(new_n8518), .Y(new_n8555));
  nor_5  g08179(.A(new_n8189), .B(new_n8095), .Y(new_n8556));
  nor_5  g08180(.A(new_n8260), .B(new_n8190), .Y(new_n8557));
  nor_5  g08181(.A(new_n8557), .B(new_n8556), .Y(new_n8558));
  xor_4  g08182(.A(new_n8550), .B(new_n8548), .Y(new_n8559));
  not_8  g08183(.A(new_n8559), .Y(new_n8560));
  nor_5  g08184(.A(new_n8560), .B(new_n8558), .Y(new_n8561));
  xor_4  g08185(.A(new_n8450), .B(new_n8449), .Y(new_n8562));
  xor_4  g08186(.A(new_n8559), .B(new_n8558), .Y(new_n8563));
  nor_5  g08187(.A(new_n8563), .B(new_n8562), .Y(new_n8564));
  nor_5  g08188(.A(new_n8564), .B(new_n8561), .Y(new_n8565));
  xor_4  g08189(.A(new_n8554), .B(new_n8518), .Y(new_n8566));
  nand_5 g08190(.A(new_n8566), .B(new_n8565), .Y(new_n8567));
  nand_5 g08191(.A(new_n8567), .B(new_n8555), .Y(new_n8568));
  nand_5 g08192(.A(pi205), .B(pi107), .Y(new_n8569));
  xor_4  g08193(.A(new_n8569), .B(new_n8568), .Y(new_n8570));
  xor_4  g08194(.A(new_n8570), .B(new_n8376), .Y(new_n8571));
  nand_5 g08195(.A(pi196), .B(pi016), .Y(new_n8572));
  nor_5  g08196(.A(new_n8509), .B(new_n8480), .Y(new_n8573));
  nor_5  g08197(.A(new_n8513), .B(new_n8510), .Y(new_n8574));
  nor_5  g08198(.A(new_n8574), .B(new_n8573), .Y(new_n8575));
  xor_4  g08199(.A(new_n8575), .B(new_n8572), .Y(new_n8576));
  not_8  g08200(.A(new_n8507), .Y(new_n8577));
  nand_5 g08201(.A(new_n8577), .B(new_n8485), .Y(new_n8578));
  not_8  g08202(.A(new_n8508), .Y(new_n8579));
  nand_5 g08203(.A(new_n8579), .B(new_n8483), .Y(new_n8580));
  nand_5 g08204(.A(new_n8580), .B(new_n8578), .Y(new_n8581));
  nor_5  g08205(.A(new_n8342), .B(new_n8318), .Y(new_n8582));
  nor_5  g08206(.A(new_n8347), .B(new_n8343), .Y(new_n8583));
  nor_5  g08207(.A(new_n8583), .B(new_n8582), .Y(new_n8584));
  nand_5 g08208(.A(new_n8290), .B(new_n8289), .Y(new_n8585));
  nand_5 g08209(.A(new_n8291), .B(new_n8288), .Y(new_n8586));
  nand_5 g08210(.A(new_n8586), .B(new_n8585), .Y(new_n8587));
  xor_4  g08211(.A(new_n8587), .B(new_n8584), .Y(new_n8588));
  xor_4  g08212(.A(new_n8588), .B(new_n8581), .Y(new_n8589));
  nand_5 g08213(.A(pi243), .B(pi163), .Y(new_n8590));
  nand_5 g08214(.A(new_n8353), .B(new_n8352), .Y(new_n8591));
  nand_5 g08215(.A(new_n8354), .B(new_n8313), .Y(new_n8592));
  nand_5 g08216(.A(new_n8592), .B(new_n8591), .Y(new_n8593));
  xor_4  g08217(.A(new_n8593), .B(new_n8590), .Y(new_n8594));
  xor_4  g08218(.A(new_n8594), .B(new_n8589), .Y(new_n8595));
  xor_4  g08219(.A(new_n8595), .B(new_n8576), .Y(new_n8596));
  nand_5 g08220(.A(pi247), .B(pi150), .Y(new_n8597));
  not_8  g08221(.A(new_n8467), .Y(new_n8598));
  nor_5  g08222(.A(new_n8471), .B(new_n8598), .Y(new_n8599));
  nor_5  g08223(.A(new_n8472), .B(new_n8464), .Y(new_n8600));
  nor_5  g08224(.A(new_n8600), .B(new_n8599), .Y(new_n8601));
  nand_5 g08225(.A(pi203), .B(pi132), .Y(new_n8602));
  xor_4  g08226(.A(new_n8602), .B(new_n8601), .Y(new_n8603));
  xor_4  g08227(.A(new_n8603), .B(new_n8597), .Y(new_n8604));
  nand_5 g08228(.A(new_n8501), .B(new_n8500), .Y(new_n8605));
  nand_5 g08229(.A(new_n8502), .B(new_n8423), .Y(new_n8606));
  nand_5 g08230(.A(new_n8606), .B(new_n8605), .Y(new_n8607));
  nand_5 g08231(.A(new_n8460), .B(new_n8459), .Y(new_n8608));
  nand_5 g08232(.A(new_n8461), .B(new_n8398), .Y(new_n8609));
  nand_5 g08233(.A(new_n8609), .B(new_n8608), .Y(new_n8610));
  nand_5 g08234(.A(new_n8469), .B(new_n8468), .Y(new_n8611));
  nand_5 g08235(.A(new_n8470), .B(new_n8385), .Y(new_n8612));
  nand_5 g08236(.A(new_n8612), .B(new_n8611), .Y(new_n8613));
  xor_4  g08237(.A(new_n8613), .B(new_n8610), .Y(new_n8614));
  nand_5 g08238(.A(pi245), .B(pi050), .Y(new_n8615));
  xor_4  g08239(.A(new_n8615), .B(new_n8614), .Y(new_n8616));
  xor_4  g08240(.A(new_n8616), .B(new_n8607), .Y(new_n8617));
  xor_4  g08241(.A(new_n8617), .B(new_n8604), .Y(new_n8618));
  nor_5  g08242(.A(new_n8538), .B(new_n8526), .Y(new_n8619));
  nor_5  g08243(.A(new_n8539), .B(new_n8535), .Y(new_n8620));
  or_6   g08244(.A(new_n8620), .B(new_n8619), .Y(new_n8621));
  nand_5 g08245(.A(pi214), .B(pi069), .Y(new_n8622));
  xor_4  g08246(.A(new_n8622), .B(new_n8621), .Y(new_n8623));
  nand_5 g08247(.A(new_n8475), .B(new_n8386), .Y(new_n8624));
  or_6   g08248(.A(new_n8477), .B(new_n8473), .Y(new_n8625));
  nand_5 g08249(.A(new_n8625), .B(new_n8624), .Y(new_n8626));
  nand_5 g08250(.A(pi116), .B(pi055), .Y(new_n8627));
  nor_5  g08251(.A(new_n8490), .B(new_n8433), .Y(new_n8628));
  nor_5  g08252(.A(new_n8495), .B(new_n8491), .Y(new_n8629));
  nor_5  g08253(.A(new_n8629), .B(new_n8628), .Y(new_n8630));
  xor_4  g08254(.A(new_n8630), .B(new_n8627), .Y(new_n8631));
  xor_4  g08255(.A(new_n8631), .B(new_n8626), .Y(new_n8632));
  xor_4  g08256(.A(new_n8632), .B(new_n8623), .Y(new_n8633));
  nand_5 g08257(.A(pi181), .B(pi058), .Y(new_n8634));
  nand_5 g08258(.A(new_n8540), .B(new_n8534), .Y(new_n8635));
  nand_5 g08259(.A(new_n8552), .B(new_n8541), .Y(new_n8636));
  nand_5 g08260(.A(new_n8636), .B(new_n8635), .Y(new_n8637));
  xor_4  g08261(.A(new_n8637), .B(new_n8634), .Y(new_n8638));
  nand_5 g08262(.A(pi226), .B(pi000), .Y(new_n8639));
  nand_5 g08263(.A(pi070), .B(pi066), .Y(new_n8640));
  xor_4  g08264(.A(new_n8640), .B(new_n8639), .Y(new_n8641));
  or_6   g08265(.A(new_n8457), .B(new_n8400), .Y(new_n8642));
  nand_5 g08266(.A(new_n8463), .B(new_n8458), .Y(new_n8643));
  nand_5 g08267(.A(new_n8643), .B(new_n8642), .Y(new_n8644));
  not_8  g08268(.A(new_n8478), .Y(new_n8645));
  nor_5  g08269(.A(new_n8645), .B(new_n8456), .Y(new_n8646));
  nor_5  g08270(.A(new_n8479), .B(new_n8455), .Y(new_n8647));
  nor_5  g08271(.A(new_n8647), .B(new_n8646), .Y(new_n8648));
  xor_4  g08272(.A(new_n8648), .B(new_n8644), .Y(new_n8649));
  nand_5 g08273(.A(pi109), .B(pi083), .Y(new_n8650));
  nand_5 g08274(.A(pi039), .B(pi002), .Y(new_n8651));
  xor_4  g08275(.A(new_n8651), .B(new_n8650), .Y(new_n8652));
  xor_4  g08276(.A(new_n8652), .B(new_n8649), .Y(new_n8653));
  xor_4  g08277(.A(new_n8653), .B(new_n8641), .Y(new_n8654));
  xor_4  g08278(.A(new_n8654), .B(new_n8638), .Y(new_n8655));
  xor_4  g08279(.A(new_n8655), .B(new_n8633), .Y(new_n8656));
  nand_5 g08280(.A(pi173), .B(pi156), .Y(new_n8657));
  nand_5 g08281(.A(pi221), .B(pi080), .Y(new_n8658));
  xor_4  g08282(.A(new_n8658), .B(new_n8657), .Y(new_n8659));
  nand_5 g08283(.A(pi202), .B(pi029), .Y(new_n8660));
  nand_5 g08284(.A(pi244), .B(pi234), .Y(new_n8661));
  nand_5 g08285(.A(pi228), .B(pi025), .Y(new_n8662));
  nand_5 g08286(.A(pi239), .B(pi148), .Y(new_n8663));
  xor_4  g08287(.A(new_n8663), .B(new_n8662), .Y(new_n8664));
  xor_4  g08288(.A(new_n8664), .B(new_n8661), .Y(new_n8665));
  xor_4  g08289(.A(new_n8665), .B(new_n8660), .Y(new_n8666));
  xor_4  g08290(.A(new_n8666), .B(new_n8659), .Y(new_n8667));
  nand_5 g08291(.A(new_n8503), .B(new_n8499), .Y(new_n8668));
  not_8  g08292(.A(new_n8496), .Y(new_n8669));
  nand_5 g08293(.A(new_n8504), .B(new_n8669), .Y(new_n8670));
  nand_5 g08294(.A(new_n8670), .B(new_n8668), .Y(new_n8671));
  nand_5 g08295(.A(new_n8493), .B(new_n8492), .Y(new_n8672));
  nand_5 g08296(.A(new_n8494), .B(new_n8431), .Y(new_n8673));
  nand_5 g08297(.A(new_n8673), .B(new_n8672), .Y(new_n8674));
  xor_4  g08298(.A(new_n8674), .B(new_n8671), .Y(new_n8675));
  nand_5 g08299(.A(pi063), .B(pi014), .Y(new_n8676));
  nand_5 g08300(.A(new_n8298), .B(new_n8281), .Y(new_n8677));
  nand_5 g08301(.A(new_n8299), .B(new_n8297), .Y(new_n8678));
  nand_5 g08302(.A(new_n8678), .B(new_n8677), .Y(new_n8679));
  xor_4  g08303(.A(new_n8679), .B(new_n8676), .Y(new_n8680));
  xor_4  g08304(.A(new_n8680), .B(new_n8675), .Y(new_n8681));
  xor_4  g08305(.A(new_n8681), .B(new_n8667), .Y(new_n8682));
  xor_4  g08306(.A(new_n8682), .B(new_n8656), .Y(new_n8683));
  xor_4  g08307(.A(new_n8683), .B(new_n8618), .Y(new_n8684));
  nand_5 g08308(.A(pi199), .B(pi149), .Y(new_n8685));
  nand_5 g08309(.A(pi211), .B(pi167), .Y(new_n8686));
  xor_4  g08310(.A(new_n8686), .B(new_n8685), .Y(new_n8687));
  nand_5 g08311(.A(pi230), .B(pi201), .Y(new_n8688));
  nand_5 g08312(.A(pi184), .B(pi117), .Y(new_n8689));
  xor_4  g08313(.A(new_n8689), .B(new_n8688), .Y(new_n8690));
  nor_5  g08314(.A(new_n8488), .B(new_n8424), .Y(new_n8691));
  nor_5  g08315(.A(new_n8506), .B(new_n8489), .Y(new_n8692));
  nor_5  g08316(.A(new_n8692), .B(new_n8691), .Y(new_n8693));
  xor_4  g08317(.A(new_n8693), .B(new_n8690), .Y(new_n8694));
  xor_4  g08318(.A(new_n8694), .B(new_n8687), .Y(new_n8695));
  xor_4  g08319(.A(new_n8695), .B(new_n8684), .Y(new_n8696));
  xor_4  g08320(.A(new_n8696), .B(new_n8596), .Y(new_n8697));
  and_6  g08321(.A(new_n8339), .B(new_n8314), .Y(new_n8698));
  nor_5  g08322(.A(new_n8358), .B(new_n8341), .Y(new_n8699));
  nor_5  g08323(.A(new_n8699), .B(new_n8698), .Y(new_n8700));
  nor_5  g08324(.A(new_n8295), .B(new_n8283), .Y(new_n8701));
  nor_5  g08325(.A(new_n8300), .B(new_n8296), .Y(new_n8702));
  nor_5  g08326(.A(new_n8702), .B(new_n8701), .Y(new_n8703));
  nand_5 g08327(.A(pi240), .B(pi195), .Y(new_n8704));
  xor_4  g08328(.A(new_n8704), .B(new_n8703), .Y(new_n8705));
  xor_4  g08329(.A(new_n8705), .B(new_n8700), .Y(new_n8706));
  or_6   g08330(.A(new_n8515), .B(new_n8452), .Y(new_n8707));
  nand_5 g08331(.A(new_n8517), .B(new_n8516), .Y(new_n8708));
  nand_5 g08332(.A(new_n8708), .B(new_n8707), .Y(new_n8709));
  nand_5 g08333(.A(new_n8355), .B(new_n8351), .Y(new_n8710));
  or_6   g08334(.A(new_n8357), .B(new_n8348), .Y(new_n8711));
  nand_5 g08335(.A(new_n8711), .B(new_n8710), .Y(new_n8712));
  nand_5 g08336(.A(new_n8345), .B(new_n8344), .Y(new_n8713));
  nand_5 g08337(.A(new_n8346), .B(new_n8316), .Y(new_n8714));
  nand_5 g08338(.A(new_n8714), .B(new_n8713), .Y(new_n8715));
  xor_4  g08339(.A(new_n8715), .B(new_n8712), .Y(new_n8716));
  xor_4  g08340(.A(new_n8716), .B(new_n8709), .Y(new_n8717));
  xor_4  g08341(.A(new_n8717), .B(new_n8706), .Y(new_n8718));
  xor_4  g08342(.A(new_n8718), .B(new_n8697), .Y(new_n8719));
  xor_4  g08343(.A(new_n8719), .B(new_n8571), .Y(po047));
  xnor_4 g08344(.A(new_n4787), .B(new_n4786), .Y(po048));
  xor_4  g08345(.A(new_n2996), .B(new_n2995), .Y(po049));
  not_8  g08346(.A(new_n1160), .Y(new_n8723));
  nand_5 g08347(.A(new_n1161), .B(new_n8723), .Y(new_n8724));
  nand_5 g08348(.A(pi133), .B(pi100), .Y(new_n8725));
  nand_5 g08349(.A(pi217), .B(pi189), .Y(new_n8726));
  nand_5 g08350(.A(pi227), .B(pi077), .Y(new_n8727));
  xor_4  g08351(.A(new_n8727), .B(new_n8726), .Y(new_n8728));
  xor_4  g08352(.A(new_n8728), .B(new_n8725), .Y(new_n8729));
  nand_5 g08353(.A(pi081), .B(pi052), .Y(new_n8730));
  nand_5 g08354(.A(new_n1151), .B(new_n1150), .Y(new_n8731));
  nand_5 g08355(.A(new_n1152), .B(new_n1149), .Y(new_n8732));
  nand_5 g08356(.A(new_n8732), .B(new_n8731), .Y(new_n8733));
  xor_4  g08357(.A(new_n8733), .B(new_n8730), .Y(new_n8734));
  xor_4  g08358(.A(new_n8734), .B(new_n8729), .Y(new_n8735));
  nand_5 g08359(.A(pi131), .B(pi106), .Y(new_n8736));
  nand_5 g08360(.A(new_n1158), .B(new_n1157), .Y(new_n8737));
  not_8  g08361(.A(new_n8737), .Y(new_n8738));
  and_6  g08362(.A(new_n1159), .B(new_n1153), .Y(new_n8739));
  nor_5  g08363(.A(new_n8739), .B(new_n8738), .Y(new_n8740));
  xor_4  g08364(.A(new_n8740), .B(new_n8736), .Y(new_n8741));
  xor_4  g08365(.A(new_n8741), .B(new_n8735), .Y(new_n8742));
  xor_4  g08366(.A(new_n8742), .B(new_n8724), .Y(new_n8743));
  nand_5 g08367(.A(new_n1208), .B(new_n1197), .Y(new_n8744));
  nand_5 g08368(.A(pi236), .B(pi231), .Y(new_n8745));
  nor_5  g08369(.A(new_n1206), .B(new_n1205), .Y(new_n8746));
  and_6  g08370(.A(new_n1207), .B(new_n1202), .Y(new_n8747));
  nor_5  g08371(.A(new_n8747), .B(new_n8746), .Y(new_n8748));
  xor_4  g08372(.A(new_n8748), .B(new_n8745), .Y(new_n8749));
  nand_5 g08373(.A(pi252), .B(pi161), .Y(new_n8750));
  nand_5 g08374(.A(pi242), .B(pi090), .Y(new_n8751));
  nand_5 g08375(.A(pi141), .B(pi140), .Y(new_n8752));
  xor_4  g08376(.A(new_n8752), .B(new_n8751), .Y(new_n8753));
  xor_4  g08377(.A(new_n8753), .B(new_n8750), .Y(new_n8754));
  nand_5 g08378(.A(pi241), .B(pi121), .Y(new_n8755));
  nand_5 g08379(.A(new_n1200), .B(new_n1199), .Y(new_n8756));
  not_8  g08380(.A(new_n1201), .Y(new_n8757));
  nand_5 g08381(.A(new_n8757), .B(new_n1198), .Y(new_n8758));
  nand_5 g08382(.A(new_n8758), .B(new_n8756), .Y(new_n8759));
  xor_4  g08383(.A(new_n8759), .B(new_n8755), .Y(new_n8760));
  xnor_4 g08384(.A(new_n8760), .B(new_n8754), .Y(new_n8761));
  xor_4  g08385(.A(new_n8761), .B(new_n8749), .Y(new_n8762));
  xor_4  g08386(.A(new_n8762), .B(new_n8744), .Y(new_n8763));
  nand_5 g08387(.A(new_n1195), .B(new_n1184), .Y(new_n8764));
  nand_5 g08388(.A(pi104), .B(pi024), .Y(new_n8765));
  nand_5 g08389(.A(pi111), .B(pi013), .Y(new_n8766));
  nand_5 g08390(.A(pi210), .B(pi112), .Y(new_n8767));
  xor_4  g08391(.A(new_n8767), .B(new_n8766), .Y(new_n8768));
  xor_4  g08392(.A(new_n8768), .B(new_n8765), .Y(new_n8769));
  nand_5 g08393(.A(pi224), .B(pi212), .Y(new_n8770));
  nand_5 g08394(.A(new_n1187), .B(new_n1186), .Y(new_n8771));
  nand_5 g08395(.A(new_n1188), .B(new_n1185), .Y(new_n8772));
  nand_5 g08396(.A(new_n8772), .B(new_n8771), .Y(new_n8773));
  xor_4  g08397(.A(new_n8773), .B(new_n8770), .Y(new_n8774));
  xor_4  g08398(.A(new_n8774), .B(new_n8769), .Y(new_n8775));
  nand_5 g08399(.A(pi255), .B(pi213), .Y(new_n8776));
  nand_5 g08400(.A(new_n1193), .B(new_n1192), .Y(new_n8777));
  nand_5 g08401(.A(new_n1194), .B(new_n1189), .Y(new_n8778));
  nand_5 g08402(.A(new_n8778), .B(new_n8777), .Y(new_n8779));
  xor_4  g08403(.A(new_n8779), .B(new_n8776), .Y(new_n8780));
  xor_4  g08404(.A(new_n8780), .B(new_n8775), .Y(new_n8781));
  xnor_4 g08405(.A(new_n8781), .B(new_n8764), .Y(new_n8782));
  nand_5 g08406(.A(new_n1210), .B(new_n1183), .Y(new_n8783));
  nand_5 g08407(.A(new_n8783), .B(new_n1211), .Y(new_n8784));
  xor_4  g08408(.A(new_n8784), .B(new_n8782), .Y(new_n8785));
  xnor_4 g08409(.A(new_n8785), .B(new_n8763), .Y(new_n8786));
  nor_5  g08410(.A(new_n1179), .B(new_n1168), .Y(new_n8787));
  nand_5 g08411(.A(pi222), .B(pi035), .Y(new_n8788));
  nand_5 g08412(.A(pi139), .B(pi125), .Y(new_n8789));
  xor_4  g08413(.A(new_n8789), .B(new_n8788), .Y(new_n8790));
  nand_5 g08414(.A(pi249), .B(pi015), .Y(new_n8791));
  xor_4  g08415(.A(new_n8791), .B(new_n8790), .Y(new_n8792));
  nand_5 g08416(.A(pi208), .B(pi176), .Y(new_n8793));
  nand_5 g08417(.A(new_n1171), .B(new_n1170), .Y(new_n8794));
  nand_5 g08418(.A(new_n1172), .B(new_n1169), .Y(new_n8795));
  nand_5 g08419(.A(new_n8795), .B(new_n8794), .Y(new_n8796));
  xor_4  g08420(.A(new_n8796), .B(new_n8793), .Y(new_n8797));
  xor_4  g08421(.A(new_n8797), .B(new_n8792), .Y(new_n8798));
  nand_5 g08422(.A(pi168), .B(pi040), .Y(new_n8799));
  nand_5 g08423(.A(new_n1177), .B(new_n1174), .Y(new_n8800));
  nand_5 g08424(.A(new_n1178), .B(new_n1173), .Y(new_n8801));
  nand_5 g08425(.A(new_n8801), .B(new_n8800), .Y(new_n8802));
  xor_4  g08426(.A(new_n8802), .B(new_n8799), .Y(new_n8803));
  xor_4  g08427(.A(new_n8803), .B(new_n8798), .Y(new_n8804));
  xor_4  g08428(.A(new_n8804), .B(new_n8787), .Y(new_n8805));
  not_8  g08429(.A(new_n1180), .Y(new_n8806));
  nor_5  g08430(.A(new_n1213), .B(new_n8806), .Y(new_n8807));
  nor_5  g08431(.A(new_n1214), .B(new_n1166), .Y(new_n8808));
  nor_5  g08432(.A(new_n8808), .B(new_n8807), .Y(new_n8809));
  xor_4  g08433(.A(new_n8809), .B(new_n8805), .Y(new_n8810));
  xnor_4 g08434(.A(new_n8810), .B(new_n8786), .Y(new_n8811));
  xnor_4 g08435(.A(new_n8811), .B(new_n8743), .Y(new_n8812));
  and_6  g08436(.A(new_n1162), .B(new_n1148), .Y(new_n8813));
  nor_5  g08437(.A(new_n1215), .B(new_n1163), .Y(new_n8814));
  nor_5  g08438(.A(new_n8814), .B(new_n8813), .Y(new_n8815));
  xnor_4 g08439(.A(new_n8815), .B(new_n8812), .Y(po050));
  nand_5 g08440(.A(pi142), .B(pi127), .Y(new_n8817));
  nand_5 g08441(.A(pi255), .B(pi142), .Y(new_n8818));
  nand_5 g08442(.A(pi111), .B(pi071), .Y(new_n8819));
  not_8  g08443(.A(new_n8819), .Y(new_n8820));
  nand_5 g08444(.A(pi210), .B(pi169), .Y(new_n8821));
  nand_5 g08445(.A(pi142), .B(pi024), .Y(new_n8822));
  nor_5  g08446(.A(new_n8822), .B(new_n8821), .Y(new_n8823));
  nor_5  g08447(.A(new_n8823), .B(new_n8820), .Y(new_n8824));
  nand_5 g08448(.A(new_n8822), .B(new_n8821), .Y(new_n8825));
  not_8  g08449(.A(new_n8825), .Y(new_n8826));
  nor_5  g08450(.A(new_n8826), .B(new_n8824), .Y(new_n8827));
  not_8  g08451(.A(new_n8827), .Y(new_n8828));
  nand_5 g08452(.A(pi224), .B(pi142), .Y(new_n8829));
  nor_5  g08453(.A(new_n8829), .B(new_n8828), .Y(new_n8830));
  nand_5 g08454(.A(pi210), .B(pi123), .Y(new_n8831));
  nand_5 g08455(.A(pi169), .B(pi111), .Y(new_n8832));
  nand_5 g08456(.A(pi071), .B(pi024), .Y(new_n8833));
  xor_4  g08457(.A(new_n8833), .B(new_n8832), .Y(new_n8834));
  xor_4  g08458(.A(new_n8834), .B(new_n8831), .Y(new_n8835));
  xor_4  g08459(.A(new_n8829), .B(new_n8827), .Y(new_n8836));
  nor_5  g08460(.A(new_n8836), .B(new_n8835), .Y(new_n8837));
  nor_5  g08461(.A(new_n8837), .B(new_n8830), .Y(new_n8838));
  xor_4  g08462(.A(new_n8838), .B(new_n8818), .Y(new_n8839));
  nand_5 g08463(.A(pi210), .B(pi099), .Y(new_n8840));
  nand_5 g08464(.A(pi169), .B(pi024), .Y(new_n8841));
  nand_5 g08465(.A(pi123), .B(pi111), .Y(new_n8842));
  xor_4  g08466(.A(new_n8842), .B(new_n8841), .Y(new_n8843));
  xor_4  g08467(.A(new_n8843), .B(new_n8840), .Y(new_n8844));
  nand_5 g08468(.A(pi224), .B(pi071), .Y(new_n8845));
  nand_5 g08469(.A(new_n8833), .B(new_n8832), .Y(new_n8846));
  nand_5 g08470(.A(new_n8834), .B(new_n8831), .Y(new_n8847));
  nand_5 g08471(.A(new_n8847), .B(new_n8846), .Y(new_n8848));
  xor_4  g08472(.A(new_n8848), .B(new_n8845), .Y(new_n8849));
  xnor_4 g08473(.A(new_n8849), .B(new_n8844), .Y(new_n8850));
  xnor_4 g08474(.A(new_n8850), .B(new_n8839), .Y(new_n8851));
  nand_5 g08475(.A(pi210), .B(pi142), .Y(new_n8852));
  and_6  g08476(.A(new_n8852), .B(new_n8820), .Y(new_n8853));
  nor_5  g08477(.A(new_n8853), .B(new_n8825), .Y(new_n8854));
  nor_5  g08478(.A(new_n8854), .B(new_n8823), .Y(new_n8855));
  nor_5  g08479(.A(new_n8855), .B(new_n8819), .Y(new_n8856));
  xor_4  g08480(.A(new_n8836), .B(new_n8835), .Y(new_n8857));
  nand_5 g08481(.A(new_n8857), .B(new_n8856), .Y(new_n8858));
  or_6   g08482(.A(new_n8858), .B(new_n8851), .Y(new_n8859));
  nand_5 g08483(.A(new_n8859), .B(new_n8817), .Y(new_n8860));
  xor_4  g08484(.A(new_n8859), .B(new_n8817), .Y(new_n8861));
  nor_5  g08485(.A(new_n8838), .B(new_n8818), .Y(new_n8862));
  nand_5 g08486(.A(new_n8850), .B(new_n8839), .Y(new_n8863));
  not_8  g08487(.A(new_n8863), .Y(new_n8864));
  nor_5  g08488(.A(new_n8864), .B(new_n8862), .Y(new_n8865));
  nand_5 g08489(.A(new_n8848), .B(new_n8845), .Y(new_n8866));
  nand_5 g08490(.A(new_n8849), .B(new_n8844), .Y(new_n8867));
  nand_5 g08491(.A(new_n8867), .B(new_n8866), .Y(new_n8868));
  nand_5 g08492(.A(pi224), .B(pi169), .Y(new_n8869));
  nand_5 g08493(.A(pi255), .B(pi071), .Y(new_n8870));
  and_6  g08494(.A(new_n8870), .B(new_n8869), .Y(new_n8871));
  nand_5 g08495(.A(pi255), .B(pi169), .Y(new_n8872));
  nor_5  g08496(.A(new_n8872), .B(new_n8845), .Y(new_n8873));
  or_6   g08497(.A(new_n8873), .B(new_n8871), .Y(new_n8874));
  nand_5 g08498(.A(new_n8842), .B(new_n8841), .Y(new_n8875));
  nand_5 g08499(.A(new_n8843), .B(new_n8840), .Y(new_n8876));
  nand_5 g08500(.A(new_n8876), .B(new_n8875), .Y(new_n8877));
  nand_5 g08501(.A(pi123), .B(pi024), .Y(new_n8878));
  nand_5 g08502(.A(pi210), .B(pi023), .Y(new_n8879));
  nand_5 g08503(.A(pi111), .B(pi099), .Y(new_n8880));
  nand_5 g08504(.A(new_n8880), .B(new_n8879), .Y(new_n8881));
  nand_5 g08505(.A(pi111), .B(pi023), .Y(new_n8882));
  nor_5  g08506(.A(new_n8882), .B(new_n8840), .Y(new_n8883));
  not_8  g08507(.A(new_n8883), .Y(new_n8884));
  nand_5 g08508(.A(new_n8884), .B(new_n8881), .Y(new_n8885));
  xor_4  g08509(.A(new_n8885), .B(new_n8878), .Y(new_n8886));
  xor_4  g08510(.A(new_n8886), .B(new_n8877), .Y(new_n8887));
  xor_4  g08511(.A(new_n8887), .B(new_n8874), .Y(new_n8888));
  xor_4  g08512(.A(new_n8888), .B(new_n8868), .Y(new_n8889));
  xnor_4 g08513(.A(new_n8889), .B(new_n8865), .Y(new_n8890));
  nand_5 g08514(.A(new_n8890), .B(new_n8861), .Y(new_n8891));
  nand_5 g08515(.A(new_n8891), .B(new_n8860), .Y(new_n8892));
  nor_5  g08516(.A(new_n8889), .B(new_n8865), .Y(new_n8893));
  not_8  g08517(.A(new_n8888), .Y(new_n8894));
  nor_5  g08518(.A(new_n8894), .B(new_n8868), .Y(new_n8895));
  nand_5 g08519(.A(new_n8895), .B(new_n8873), .Y(new_n8896));
  or_6   g08520(.A(new_n8894), .B(new_n8868), .Y(new_n8897));
  nor_5  g08521(.A(new_n8887), .B(new_n8874), .Y(new_n8898));
  nor_5  g08522(.A(new_n8898), .B(new_n8873), .Y(new_n8899));
  nand_5 g08523(.A(new_n8899), .B(new_n8897), .Y(new_n8900));
  nand_5 g08524(.A(new_n8900), .B(new_n8896), .Y(new_n8901));
  nand_5 g08525(.A(pi099), .B(pi024), .Y(new_n8902));
  nand_5 g08526(.A(pi210), .B(pi155), .Y(new_n8903));
  xor_4  g08527(.A(new_n8903), .B(new_n8882), .Y(new_n8904));
  xor_4  g08528(.A(new_n8904), .B(new_n8902), .Y(new_n8905));
  nand_5 g08529(.A(pi224), .B(pi123), .Y(new_n8906));
  xor_4  g08530(.A(new_n8906), .B(new_n8883), .Y(new_n8907));
  xor_4  g08531(.A(new_n8907), .B(new_n8905), .Y(new_n8908));
  nand_5 g08532(.A(new_n8885), .B(new_n8878), .Y(new_n8909));
  nand_5 g08533(.A(new_n8886), .B(new_n8877), .Y(new_n8910));
  nand_5 g08534(.A(new_n8910), .B(new_n8909), .Y(new_n8911));
  nand_5 g08535(.A(pi127), .B(pi071), .Y(new_n8912));
  nand_5 g08536(.A(pi232), .B(pi142), .Y(new_n8913));
  xor_4  g08537(.A(new_n8913), .B(new_n8912), .Y(new_n8914));
  xor_4  g08538(.A(new_n8914), .B(new_n8872), .Y(new_n8915));
  xor_4  g08539(.A(new_n8915), .B(new_n8911), .Y(new_n8916));
  xor_4  g08540(.A(new_n8916), .B(new_n8908), .Y(new_n8917));
  xor_4  g08541(.A(new_n8917), .B(new_n8901), .Y(new_n8918));
  xor_4  g08542(.A(new_n8918), .B(new_n8893), .Y(new_n8919));
  xor_4  g08543(.A(new_n8919), .B(new_n8892), .Y(new_n8920));
  nand_5 g08544(.A(pi140), .B(pi135), .Y(new_n8921));
  nand_5 g08545(.A(pi252), .B(pi122), .Y(new_n8922));
  nand_5 g08546(.A(pi242), .B(pi059), .Y(new_n8923));
  xor_4  g08547(.A(new_n8923), .B(new_n8922), .Y(new_n8924));
  xor_4  g08548(.A(new_n8924), .B(new_n8921), .Y(new_n8925));
  nand_5 g08549(.A(pi121), .B(pi001), .Y(new_n8926));
  nand_5 g08550(.A(pi242), .B(pi122), .Y(new_n8927));
  nor_5  g08551(.A(new_n8927), .B(new_n8921), .Y(new_n8928));
  xor_4  g08552(.A(new_n8928), .B(new_n8926), .Y(new_n8929));
  xor_4  g08553(.A(new_n8929), .B(new_n8925), .Y(new_n8930));
  not_8  g08554(.A(new_n8928), .Y(new_n8931));
  nand_5 g08555(.A(pi242), .B(pi135), .Y(new_n8932));
  nand_5 g08556(.A(pi140), .B(pi122), .Y(new_n8933));
  nand_5 g08557(.A(new_n8933), .B(new_n8932), .Y(new_n8934));
  nand_5 g08558(.A(new_n8934), .B(new_n8931), .Y(new_n8935));
  nand_5 g08559(.A(pi252), .B(pi001), .Y(new_n8936));
  nand_5 g08560(.A(new_n8936), .B(new_n8935), .Y(new_n8937));
  nand_5 g08561(.A(pi140), .B(pi001), .Y(new_n8938));
  nand_5 g08562(.A(new_n8938), .B(new_n8927), .Y(new_n8939));
  nand_5 g08563(.A(pi252), .B(pi102), .Y(new_n8940));
  xor_4  g08564(.A(new_n8938), .B(new_n8927), .Y(new_n8941));
  nand_5 g08565(.A(new_n8941), .B(new_n8940), .Y(new_n8942));
  nand_5 g08566(.A(new_n8942), .B(new_n8939), .Y(new_n8943));
  xor_4  g08567(.A(new_n8936), .B(new_n8935), .Y(new_n8944));
  nand_5 g08568(.A(new_n8944), .B(new_n8943), .Y(new_n8945));
  nand_5 g08569(.A(new_n8945), .B(new_n8937), .Y(new_n8946));
  nand_5 g08570(.A(pi231), .B(pi102), .Y(new_n8947));
  nand_5 g08571(.A(pi087), .B(pi021), .Y(new_n8948));
  nand_5 g08572(.A(pi219), .B(pi005), .Y(new_n8949));
  xor_4  g08573(.A(new_n8949), .B(new_n8948), .Y(new_n8950));
  xor_4  g08574(.A(new_n8950), .B(new_n8947), .Y(new_n8951));
  xnor_4 g08575(.A(new_n8951), .B(new_n8946), .Y(new_n8952));
  xor_4  g08576(.A(new_n8952), .B(new_n8930), .Y(new_n8953));
  nand_5 g08577(.A(pi219), .B(pi121), .Y(new_n8954));
  or_6   g08578(.A(new_n8954), .B(new_n8947), .Y(new_n8955));
  nand_5 g08579(.A(pi242), .B(pi001), .Y(new_n8956));
  nand_5 g08580(.A(pi252), .B(pi219), .Y(new_n8957));
  and_6  g08581(.A(new_n8957), .B(new_n8956), .Y(new_n8958));
  nand_5 g08582(.A(pi140), .B(pi102), .Y(new_n8959));
  xor_4  g08583(.A(new_n8957), .B(new_n8956), .Y(new_n8960));
  and_6  g08584(.A(new_n8960), .B(new_n8959), .Y(new_n8961));
  or_6   g08585(.A(new_n8961), .B(new_n8958), .Y(new_n8962));
  and_6  g08586(.A(new_n8962), .B(new_n8954), .Y(new_n8963));
  xor_4  g08587(.A(new_n8941), .B(new_n8940), .Y(new_n8964));
  xor_4  g08588(.A(new_n8962), .B(new_n8954), .Y(new_n8965));
  and_6  g08589(.A(new_n8965), .B(new_n8964), .Y(new_n8966));
  or_6   g08590(.A(new_n8966), .B(new_n8963), .Y(new_n8967));
  nand_5 g08591(.A(pi121), .B(pi102), .Y(new_n8968));
  nand_5 g08592(.A(pi231), .B(pi219), .Y(new_n8969));
  nand_5 g08593(.A(new_n8969), .B(new_n8968), .Y(new_n8970));
  nand_5 g08594(.A(new_n8970), .B(new_n8955), .Y(new_n8971));
  nand_5 g08595(.A(new_n8971), .B(new_n8967), .Y(new_n8972));
  xor_4  g08596(.A(new_n8944), .B(new_n8943), .Y(new_n8973));
  xor_4  g08597(.A(new_n8971), .B(new_n8967), .Y(new_n8974));
  nand_5 g08598(.A(new_n8974), .B(new_n8973), .Y(new_n8975));
  nand_5 g08599(.A(new_n8975), .B(new_n8972), .Y(new_n8976));
  xor_4  g08600(.A(new_n8976), .B(new_n8955), .Y(new_n8977));
  xor_4  g08601(.A(new_n8977), .B(new_n8953), .Y(new_n8978));
  not_8  g08602(.A(new_n8978), .Y(new_n8979));
  nand_5 g08603(.A(pi231), .B(pi087), .Y(new_n8980));
  nand_5 g08604(.A(pi219), .B(pi140), .Y(new_n8981));
  not_8  g08605(.A(new_n8981), .Y(new_n8982));
  nand_5 g08606(.A(pi242), .B(pi102), .Y(new_n8983));
  nand_5 g08607(.A(pi252), .B(pi087), .Y(new_n8984));
  nor_5  g08608(.A(new_n8984), .B(new_n8983), .Y(new_n8985));
  or_6   g08609(.A(new_n8985), .B(new_n8982), .Y(new_n8986));
  nand_5 g08610(.A(new_n8984), .B(new_n8983), .Y(new_n8987));
  nand_5 g08611(.A(new_n8987), .B(new_n8986), .Y(new_n8988));
  nand_5 g08612(.A(pi121), .B(pi087), .Y(new_n8989));
  nor_5  g08613(.A(new_n8989), .B(new_n8988), .Y(new_n8990));
  xor_4  g08614(.A(new_n8960), .B(new_n8959), .Y(new_n8991));
  xnor_4 g08615(.A(new_n8989), .B(new_n8988), .Y(new_n8992));
  nor_5  g08616(.A(new_n8992), .B(new_n8991), .Y(new_n8993));
  nor_5  g08617(.A(new_n8993), .B(new_n8990), .Y(new_n8994));
  nor_5  g08618(.A(new_n8994), .B(new_n8980), .Y(new_n8995));
  xnor_4 g08619(.A(new_n8994), .B(new_n8980), .Y(new_n8996));
  xor_4  g08620(.A(new_n8965), .B(new_n8964), .Y(new_n8997));
  nor_5  g08621(.A(new_n8997), .B(new_n8996), .Y(new_n8998));
  nor_5  g08622(.A(new_n8998), .B(new_n8995), .Y(new_n8999));
  xor_4  g08623(.A(new_n8974), .B(new_n8973), .Y(new_n9000));
  nor_5  g08624(.A(new_n9000), .B(new_n8999), .Y(new_n9001));
  nand_5 g08625(.A(pi087), .B(pi005), .Y(new_n9002));
  xnor_4 g08626(.A(new_n9000), .B(new_n8999), .Y(new_n9003));
  xor_4  g08627(.A(new_n9003), .B(new_n9002), .Y(new_n9004));
  nand_5 g08628(.A(pi242), .B(pi087), .Y(new_n9005));
  and_6  g08629(.A(new_n9005), .B(new_n8982), .Y(new_n9006));
  nor_5  g08630(.A(new_n9006), .B(new_n8987), .Y(new_n9007));
  nor_5  g08631(.A(new_n9007), .B(new_n8985), .Y(new_n9008));
  or_6   g08632(.A(new_n9008), .B(new_n8981), .Y(new_n9009));
  xnor_4 g08633(.A(new_n8992), .B(new_n8991), .Y(new_n9010));
  nor_5  g08634(.A(new_n9010), .B(new_n9009), .Y(new_n9011));
  not_8  g08635(.A(new_n9011), .Y(new_n9012));
  xnor_4 g08636(.A(new_n8997), .B(new_n8996), .Y(new_n9013));
  nor_5  g08637(.A(new_n9013), .B(new_n9012), .Y(new_n9014));
  and_6  g08638(.A(new_n9014), .B(new_n9004), .Y(new_n9015));
  nand_5 g08639(.A(new_n9015), .B(new_n9001), .Y(new_n9016));
  nand_5 g08640(.A(new_n9014), .B(new_n9004), .Y(new_n9017));
  nor_5  g08641(.A(new_n9003), .B(new_n9002), .Y(new_n9018));
  nor_5  g08642(.A(new_n9018), .B(new_n9001), .Y(new_n9019));
  nand_5 g08643(.A(new_n9019), .B(new_n9017), .Y(new_n9020));
  nand_5 g08644(.A(new_n9020), .B(new_n9016), .Y(new_n9021));
  xor_4  g08645(.A(new_n9021), .B(new_n8979), .Y(new_n9022));
  xor_4  g08646(.A(new_n9022), .B(new_n8920), .Y(new_n9023));
  xnor_4 g08647(.A(new_n9014), .B(new_n9004), .Y(new_n9024));
  xor_4  g08648(.A(new_n8890), .B(new_n8861), .Y(new_n9025));
  nor_5  g08649(.A(new_n9025), .B(new_n9024), .Y(new_n9026));
  xnor_4 g08650(.A(new_n9025), .B(new_n9024), .Y(new_n9027));
  xor_4  g08651(.A(new_n8858), .B(new_n8851), .Y(new_n9028));
  not_8  g08652(.A(new_n9028), .Y(new_n9029));
  xor_4  g08653(.A(new_n9013), .B(new_n9011), .Y(new_n9030));
  nor_5  g08654(.A(new_n9030), .B(new_n9029), .Y(new_n9031));
  nand_5 g08655(.A(new_n8853), .B(new_n8825), .Y(new_n9032));
  nand_5 g08656(.A(new_n9032), .B(new_n8855), .Y(new_n9033));
  nand_5 g08657(.A(new_n9006), .B(new_n8987), .Y(new_n9034));
  nand_5 g08658(.A(new_n9034), .B(new_n9008), .Y(new_n9035));
  nand_5 g08659(.A(new_n9035), .B(new_n9033), .Y(new_n9036));
  xnor_4 g08660(.A(new_n9035), .B(new_n9033), .Y(new_n9037));
  nand_5 g08661(.A(pi142), .B(pi111), .Y(new_n9038));
  nand_5 g08662(.A(pi210), .B(pi071), .Y(new_n9039));
  xor_4  g08663(.A(new_n9039), .B(new_n9038), .Y(new_n9040));
  nor_5  g08664(.A(new_n9005), .B(new_n8852), .Y(new_n9041));
  nand_5 g08665(.A(new_n9041), .B(new_n9040), .Y(new_n9042));
  nand_5 g08666(.A(pi242), .B(pi219), .Y(new_n9043));
  nand_5 g08667(.A(pi140), .B(pi087), .Y(new_n9044));
  xor_4  g08668(.A(new_n9044), .B(new_n9043), .Y(new_n9045));
  xor_4  g08669(.A(new_n9041), .B(new_n9040), .Y(new_n9046));
  nand_5 g08670(.A(new_n9046), .B(new_n9045), .Y(new_n9047));
  nand_5 g08671(.A(new_n9047), .B(new_n9042), .Y(new_n9048));
  or_6   g08672(.A(new_n9048), .B(new_n9037), .Y(new_n9049));
  nand_5 g08673(.A(new_n9049), .B(new_n9036), .Y(new_n9050));
  xor_4  g08674(.A(new_n9010), .B(new_n9009), .Y(new_n9051));
  not_8  g08675(.A(new_n9051), .Y(new_n9052));
  nand_5 g08676(.A(new_n9052), .B(new_n9050), .Y(new_n9053));
  xor_4  g08677(.A(new_n8857), .B(new_n8856), .Y(new_n9054));
  xor_4  g08678(.A(new_n9051), .B(new_n9050), .Y(new_n9055));
  or_6   g08679(.A(new_n9055), .B(new_n9054), .Y(new_n9056));
  nand_5 g08680(.A(new_n9056), .B(new_n9053), .Y(new_n9057));
  xor_4  g08681(.A(new_n9030), .B(new_n9028), .Y(new_n9058));
  nor_5  g08682(.A(new_n9058), .B(new_n9057), .Y(new_n9059));
  nor_5  g08683(.A(new_n9059), .B(new_n9031), .Y(new_n9060));
  nor_5  g08684(.A(new_n9060), .B(new_n9027), .Y(new_n9061));
  nor_5  g08685(.A(new_n9061), .B(new_n9026), .Y(new_n9062));
  xor_4  g08686(.A(new_n9062), .B(new_n9023), .Y(new_n9063));
  nand_5 g08687(.A(pi174), .B(pi138), .Y(new_n9064));
  nand_5 g08688(.A(pi222), .B(pi182), .Y(new_n9065));
  nand_5 g08689(.A(pi249), .B(pi041), .Y(new_n9066));
  nand_5 g08690(.A(pi138), .B(pi125), .Y(new_n9067));
  or_6   g08691(.A(new_n9067), .B(new_n9066), .Y(new_n9068));
  nand_5 g08692(.A(new_n9068), .B(new_n9065), .Y(new_n9069));
  nand_5 g08693(.A(new_n9067), .B(new_n9066), .Y(new_n9070));
  nand_5 g08694(.A(new_n9070), .B(new_n9069), .Y(new_n9071));
  nand_5 g08695(.A(pi176), .B(pi138), .Y(new_n9072));
  nor_5  g08696(.A(new_n9072), .B(new_n9071), .Y(new_n9073));
  nand_5 g08697(.A(pi182), .B(pi125), .Y(new_n9074));
  nand_5 g08698(.A(pi222), .B(pi041), .Y(new_n9075));
  nand_5 g08699(.A(pi249), .B(pi216), .Y(new_n9076));
  xor_4  g08700(.A(new_n9076), .B(new_n9075), .Y(new_n9077));
  xor_4  g08701(.A(new_n9077), .B(new_n9074), .Y(new_n9078));
  xor_4  g08702(.A(new_n9072), .B(new_n9071), .Y(new_n9079));
  not_8  g08703(.A(new_n9079), .Y(new_n9080));
  nor_5  g08704(.A(new_n9080), .B(new_n9078), .Y(new_n9081));
  nor_5  g08705(.A(new_n9081), .B(new_n9073), .Y(new_n9082));
  nand_5 g08706(.A(pi138), .B(pi040), .Y(new_n9083));
  nand_5 g08707(.A(pi222), .B(pi216), .Y(new_n9084));
  nand_5 g08708(.A(pi125), .B(pi041), .Y(new_n9085));
  nand_5 g08709(.A(pi249), .B(pi076), .Y(new_n9086));
  xor_4  g08710(.A(new_n9086), .B(new_n9085), .Y(new_n9087));
  xor_4  g08711(.A(new_n9087), .B(new_n9084), .Y(new_n9088));
  nand_5 g08712(.A(pi182), .B(pi176), .Y(new_n9089));
  nand_5 g08713(.A(new_n9076), .B(new_n9075), .Y(new_n9090));
  nand_5 g08714(.A(new_n9077), .B(new_n9074), .Y(new_n9091));
  nand_5 g08715(.A(new_n9091), .B(new_n9090), .Y(new_n9092));
  xor_4  g08716(.A(new_n9092), .B(new_n9089), .Y(new_n9093));
  xor_4  g08717(.A(new_n9093), .B(new_n9088), .Y(new_n9094));
  xnor_4 g08718(.A(new_n9094), .B(new_n9083), .Y(new_n9095));
  xor_4  g08719(.A(new_n9095), .B(new_n9082), .Y(new_n9096));
  nand_5 g08720(.A(pi249), .B(pi138), .Y(new_n9097));
  not_8  g08721(.A(new_n9097), .Y(new_n9098));
  nor_5  g08722(.A(new_n9098), .B(new_n9065), .Y(new_n9099));
  or_6   g08723(.A(new_n9099), .B(new_n9070), .Y(new_n9100));
  and_6  g08724(.A(new_n9100), .B(new_n9068), .Y(new_n9101));
  nor_5  g08725(.A(new_n9101), .B(new_n9065), .Y(new_n9102));
  not_8  g08726(.A(new_n9102), .Y(new_n9103));
  xor_4  g08727(.A(new_n9079), .B(new_n9078), .Y(new_n9104));
  nor_5  g08728(.A(new_n9104), .B(new_n9103), .Y(new_n9105));
  nand_5 g08729(.A(new_n9105), .B(new_n9096), .Y(new_n9106));
  nand_5 g08730(.A(new_n9106), .B(new_n9064), .Y(new_n9107));
  xor_4  g08731(.A(new_n9106), .B(new_n9064), .Y(new_n9108));
  nor_5  g08732(.A(new_n9094), .B(new_n9083), .Y(new_n9109));
  nor_5  g08733(.A(new_n9095), .B(new_n9082), .Y(new_n9110));
  nor_5  g08734(.A(new_n9110), .B(new_n9109), .Y(new_n9111));
  nand_5 g08735(.A(new_n9086), .B(new_n9085), .Y(new_n9112));
  nand_5 g08736(.A(new_n9087), .B(new_n9084), .Y(new_n9113));
  nand_5 g08737(.A(new_n9113), .B(new_n9112), .Y(new_n9114));
  nand_5 g08738(.A(pi216), .B(pi125), .Y(new_n9115));
  nand_5 g08739(.A(pi222), .B(pi076), .Y(new_n9116));
  nand_5 g08740(.A(pi249), .B(pi079), .Y(new_n9117));
  nand_5 g08741(.A(new_n9117), .B(new_n9116), .Y(new_n9118));
  nand_5 g08742(.A(pi222), .B(pi079), .Y(new_n9119));
  nor_5  g08743(.A(new_n9119), .B(new_n9086), .Y(new_n9120));
  not_8  g08744(.A(new_n9120), .Y(new_n9121));
  nand_5 g08745(.A(new_n9121), .B(new_n9118), .Y(new_n9122));
  xor_4  g08746(.A(new_n9122), .B(new_n9115), .Y(new_n9123));
  xor_4  g08747(.A(new_n9123), .B(new_n9114), .Y(new_n9124));
  nand_5 g08748(.A(new_n9092), .B(new_n9089), .Y(new_n9125));
  nand_5 g08749(.A(new_n9093), .B(new_n9088), .Y(new_n9126));
  nand_5 g08750(.A(new_n9126), .B(new_n9125), .Y(new_n9127));
  nand_5 g08751(.A(pi176), .B(pi041), .Y(new_n9128));
  nand_5 g08752(.A(pi182), .B(pi040), .Y(new_n9129));
  nand_5 g08753(.A(new_n9129), .B(new_n9128), .Y(new_n9130));
  nand_5 g08754(.A(pi041), .B(pi040), .Y(new_n9131));
  nor_5  g08755(.A(new_n9131), .B(new_n9089), .Y(new_n9132));
  not_8  g08756(.A(new_n9132), .Y(new_n9133));
  nand_5 g08757(.A(new_n9133), .B(new_n9130), .Y(new_n9134));
  xor_4  g08758(.A(new_n9134), .B(new_n9127), .Y(new_n9135));
  xor_4  g08759(.A(new_n9135), .B(new_n9124), .Y(new_n9136));
  xnor_4 g08760(.A(new_n9136), .B(new_n9111), .Y(new_n9137));
  nand_5 g08761(.A(new_n9137), .B(new_n9108), .Y(new_n9138));
  nand_5 g08762(.A(new_n9138), .B(new_n9107), .Y(new_n9139));
  nor_5  g08763(.A(new_n9136), .B(new_n9111), .Y(new_n9140));
  nand_5 g08764(.A(pi125), .B(pi076), .Y(new_n9141));
  nand_5 g08765(.A(pi251), .B(pi249), .Y(new_n9142));
  xor_4  g08766(.A(new_n9142), .B(new_n9141), .Y(new_n9143));
  xor_4  g08767(.A(new_n9143), .B(new_n9119), .Y(new_n9144));
  nand_5 g08768(.A(pi216), .B(pi176), .Y(new_n9145));
  xor_4  g08769(.A(new_n9145), .B(new_n9120), .Y(new_n9146));
  xor_4  g08770(.A(new_n9146), .B(new_n9144), .Y(new_n9147));
  nand_5 g08771(.A(new_n9122), .B(new_n9115), .Y(new_n9148));
  nand_5 g08772(.A(new_n9123), .B(new_n9114), .Y(new_n9149));
  nand_5 g08773(.A(new_n9149), .B(new_n9148), .Y(new_n9150));
  nand_5 g08774(.A(pi182), .B(pi174), .Y(new_n9151));
  and_6  g08775(.A(pi157), .B(pi138), .Y(new_n9152));
  xor_4  g08776(.A(new_n9152), .B(new_n9151), .Y(new_n9153));
  xor_4  g08777(.A(new_n9153), .B(new_n9131), .Y(new_n9154));
  xor_4  g08778(.A(new_n9154), .B(new_n9150), .Y(new_n9155));
  xnor_4 g08779(.A(new_n9155), .B(new_n9147), .Y(new_n9156));
  nand_5 g08780(.A(new_n9134), .B(new_n9127), .Y(new_n9157));
  nand_5 g08781(.A(new_n9135), .B(new_n9124), .Y(new_n9158));
  nand_5 g08782(.A(new_n9158), .B(new_n9157), .Y(new_n9159));
  xor_4  g08783(.A(new_n9159), .B(new_n9132), .Y(new_n9160));
  xor_4  g08784(.A(new_n9160), .B(new_n9156), .Y(new_n9161));
  xor_4  g08785(.A(new_n9161), .B(new_n9140), .Y(new_n9162));
  xor_4  g08786(.A(new_n9162), .B(new_n9139), .Y(new_n9163));
  xor_4  g08787(.A(new_n9163), .B(new_n9063), .Y(new_n9164));
  xor_4  g08788(.A(new_n9137), .B(new_n9108), .Y(new_n9165));
  xnor_4 g08789(.A(new_n9060), .B(new_n9027), .Y(new_n9166));
  nor_5  g08790(.A(new_n9166), .B(new_n9165), .Y(new_n9167));
  xor_4  g08791(.A(new_n9055), .B(new_n9054), .Y(new_n9168));
  xor_4  g08792(.A(new_n9104), .B(new_n9102), .Y(new_n9169));
  nand_5 g08793(.A(new_n9169), .B(new_n9168), .Y(new_n9170));
  xor_4  g08794(.A(new_n9169), .B(new_n9168), .Y(new_n9171));
  xor_4  g08795(.A(new_n9005), .B(new_n8852), .Y(new_n9172));
  and_6  g08796(.A(new_n9172), .B(new_n9098), .Y(new_n9173));
  nand_5 g08797(.A(pi222), .B(pi138), .Y(new_n9174));
  nand_5 g08798(.A(pi249), .B(pi182), .Y(new_n9175));
  xor_4  g08799(.A(new_n9175), .B(new_n9174), .Y(new_n9176));
  nor_5  g08800(.A(new_n9176), .B(new_n9173), .Y(new_n9177));
  xor_4  g08801(.A(new_n9176), .B(new_n9173), .Y(new_n9178));
  xor_4  g08802(.A(new_n9046), .B(new_n9045), .Y(new_n9179));
  not_8  g08803(.A(new_n9179), .Y(new_n9180));
  nand_5 g08804(.A(new_n9180), .B(new_n9178), .Y(new_n9181));
  not_8  g08805(.A(new_n9181), .Y(new_n9182));
  nor_5  g08806(.A(new_n9182), .B(new_n9177), .Y(new_n9183));
  xnor_4 g08807(.A(new_n9048), .B(new_n9037), .Y(new_n9184));
  and_6  g08808(.A(new_n9184), .B(new_n9183), .Y(new_n9185));
  xnor_4 g08809(.A(new_n9184), .B(new_n9183), .Y(new_n9186));
  nand_5 g08810(.A(new_n9099), .B(new_n9070), .Y(new_n9187));
  nand_5 g08811(.A(new_n9187), .B(new_n9101), .Y(new_n9188));
  nor_5  g08812(.A(new_n9188), .B(new_n9186), .Y(new_n9189));
  nor_5  g08813(.A(new_n9189), .B(new_n9185), .Y(new_n9190));
  nand_5 g08814(.A(new_n9190), .B(new_n9171), .Y(new_n9191));
  nand_5 g08815(.A(new_n9191), .B(new_n9170), .Y(new_n9192));
  xor_4  g08816(.A(new_n9105), .B(new_n9096), .Y(new_n9193));
  not_8  g08817(.A(new_n9193), .Y(new_n9194));
  nand_5 g08818(.A(new_n9194), .B(new_n9192), .Y(new_n9195));
  xor_4  g08819(.A(new_n9194), .B(new_n9192), .Y(new_n9196));
  xnor_4 g08820(.A(new_n9058), .B(new_n9057), .Y(new_n9197));
  nand_5 g08821(.A(new_n9197), .B(new_n9196), .Y(new_n9198));
  nand_5 g08822(.A(new_n9198), .B(new_n9195), .Y(new_n9199));
  xnor_4 g08823(.A(new_n9166), .B(new_n9165), .Y(new_n9200));
  nor_5  g08824(.A(new_n9200), .B(new_n9199), .Y(new_n9201));
  nor_5  g08825(.A(new_n9201), .B(new_n9167), .Y(new_n9202));
  xor_4  g08826(.A(new_n9202), .B(new_n9164), .Y(new_n9203));
  nand_5 g08827(.A(pi160), .B(pi081), .Y(new_n9204));
  nand_5 g08828(.A(pi227), .B(pi160), .Y(new_n9205));
  nand_5 g08829(.A(pi100), .B(pi020), .Y(new_n9206));
  nand_5 g08830(.A(new_n9206), .B(new_n9205), .Y(new_n9207));
  nand_5 g08831(.A(pi217), .B(pi060), .Y(new_n9208));
  xor_4  g08832(.A(new_n9206), .B(new_n9205), .Y(new_n9209));
  nand_5 g08833(.A(new_n9209), .B(new_n9208), .Y(new_n9210));
  nand_5 g08834(.A(new_n9210), .B(new_n9207), .Y(new_n9211));
  nor_5  g08835(.A(new_n9211), .B(new_n9204), .Y(new_n9212));
  nand_5 g08836(.A(pi227), .B(pi020), .Y(new_n9213));
  nand_5 g08837(.A(pi223), .B(pi217), .Y(new_n9214));
  nand_5 g08838(.A(pi100), .B(pi060), .Y(new_n9215));
  xor_4  g08839(.A(new_n9215), .B(new_n9214), .Y(new_n9216));
  xor_4  g08840(.A(new_n9216), .B(new_n9213), .Y(new_n9217));
  xor_4  g08841(.A(new_n9211), .B(new_n9204), .Y(new_n9218));
  not_8  g08842(.A(new_n9218), .Y(new_n9219));
  nor_5  g08843(.A(new_n9219), .B(new_n9217), .Y(new_n9220));
  nor_5  g08844(.A(new_n9220), .B(new_n9212), .Y(new_n9221));
  nand_5 g08845(.A(pi160), .B(pi106), .Y(new_n9222));
  nand_5 g08846(.A(pi227), .B(pi060), .Y(new_n9223));
  nand_5 g08847(.A(pi217), .B(pi101), .Y(new_n9224));
  nand_5 g08848(.A(pi223), .B(pi100), .Y(new_n9225));
  xor_4  g08849(.A(new_n9225), .B(new_n9224), .Y(new_n9226));
  xor_4  g08850(.A(new_n9226), .B(new_n9223), .Y(new_n9227));
  nand_5 g08851(.A(pi081), .B(pi020), .Y(new_n9228));
  nand_5 g08852(.A(new_n9215), .B(new_n9214), .Y(new_n9229));
  nand_5 g08853(.A(new_n9216), .B(new_n9213), .Y(new_n9230));
  nand_5 g08854(.A(new_n9230), .B(new_n9229), .Y(new_n9231));
  xor_4  g08855(.A(new_n9231), .B(new_n9228), .Y(new_n9232));
  xor_4  g08856(.A(new_n9232), .B(new_n9227), .Y(new_n9233));
  xnor_4 g08857(.A(new_n9233), .B(new_n9222), .Y(new_n9234));
  xor_4  g08858(.A(new_n9234), .B(new_n9221), .Y(new_n9235));
  xor_4  g08859(.A(new_n9209), .B(new_n9208), .Y(new_n9236));
  not_8  g08860(.A(new_n9236), .Y(new_n9237));
  nand_5 g08861(.A(pi160), .B(pi100), .Y(new_n9238));
  nand_5 g08862(.A(pi217), .B(pi020), .Y(new_n9239));
  nor_5  g08863(.A(new_n9239), .B(new_n9238), .Y(new_n9240));
  nand_5 g08864(.A(new_n9240), .B(new_n9237), .Y(new_n9241));
  xor_4  g08865(.A(new_n9218), .B(new_n9217), .Y(new_n9242));
  nor_5  g08866(.A(new_n9242), .B(new_n9241), .Y(new_n9243));
  nand_5 g08867(.A(new_n9243), .B(new_n9235), .Y(new_n9244));
  nand_5 g08868(.A(pi233), .B(pi160), .Y(new_n9245));
  nand_5 g08869(.A(new_n9245), .B(new_n9244), .Y(new_n9246));
  xor_4  g08870(.A(new_n9245), .B(new_n9244), .Y(new_n9247));
  nor_5  g08871(.A(new_n9233), .B(new_n9222), .Y(new_n9248));
  nor_5  g08872(.A(new_n9234), .B(new_n9221), .Y(new_n9249));
  nor_5  g08873(.A(new_n9249), .B(new_n9248), .Y(new_n9250));
  nand_5 g08874(.A(new_n9231), .B(new_n9228), .Y(new_n9251));
  nand_5 g08875(.A(new_n9232), .B(new_n9227), .Y(new_n9252));
  nand_5 g08876(.A(new_n9252), .B(new_n9251), .Y(new_n9253));
  nand_5 g08877(.A(pi081), .B(pi060), .Y(new_n9254));
  nand_5 g08878(.A(pi106), .B(pi020), .Y(new_n9255));
  nand_5 g08879(.A(new_n9255), .B(new_n9254), .Y(new_n9256));
  nand_5 g08880(.A(pi106), .B(pi060), .Y(new_n9257));
  nor_5  g08881(.A(new_n9257), .B(new_n9228), .Y(new_n9258));
  not_8  g08882(.A(new_n9258), .Y(new_n9259));
  nand_5 g08883(.A(new_n9259), .B(new_n9256), .Y(new_n9260));
  nand_5 g08884(.A(new_n9225), .B(new_n9224), .Y(new_n9261));
  nand_5 g08885(.A(new_n9226), .B(new_n9223), .Y(new_n9262));
  nand_5 g08886(.A(new_n9262), .B(new_n9261), .Y(new_n9263));
  nand_5 g08887(.A(pi227), .B(pi223), .Y(new_n9264));
  nand_5 g08888(.A(pi225), .B(pi100), .Y(new_n9265));
  nor_5  g08889(.A(new_n9265), .B(new_n9224), .Y(new_n9266));
  not_8  g08890(.A(new_n9266), .Y(new_n9267));
  nand_5 g08891(.A(pi101), .B(pi100), .Y(new_n9268));
  nand_5 g08892(.A(pi225), .B(pi217), .Y(new_n9269));
  nand_5 g08893(.A(new_n9269), .B(new_n9268), .Y(new_n9270));
  nand_5 g08894(.A(new_n9270), .B(new_n9267), .Y(new_n9271));
  xor_4  g08895(.A(new_n9271), .B(new_n9264), .Y(new_n9272));
  xor_4  g08896(.A(new_n9272), .B(new_n9263), .Y(new_n9273));
  xor_4  g08897(.A(new_n9273), .B(new_n9260), .Y(new_n9274));
  xor_4  g08898(.A(new_n9274), .B(new_n9253), .Y(new_n9275));
  xor_4  g08899(.A(new_n9275), .B(new_n9250), .Y(new_n9276));
  not_8  g08900(.A(new_n9276), .Y(new_n9277));
  nand_5 g08901(.A(new_n9277), .B(new_n9247), .Y(new_n9278));
  nand_5 g08902(.A(new_n9278), .B(new_n9246), .Y(new_n9279));
  nor_5  g08903(.A(new_n9275), .B(new_n9250), .Y(new_n9280));
  nor_5  g08904(.A(new_n9273), .B(new_n9260), .Y(new_n9281));
  not_8  g08905(.A(new_n9274), .Y(new_n9282));
  nor_5  g08906(.A(new_n9282), .B(new_n9253), .Y(new_n9283));
  xor_4  g08907(.A(new_n9283), .B(new_n9259), .Y(new_n9284));
  not_8  g08908(.A(new_n9284), .Y(new_n9285));
  nor_5  g08909(.A(new_n9285), .B(new_n9281), .Y(new_n9286));
  nand_5 g08910(.A(pi227), .B(pi101), .Y(new_n9287));
  nand_5 g08911(.A(pi217), .B(pi177), .Y(new_n9288));
  xor_4  g08912(.A(new_n9288), .B(new_n9287), .Y(new_n9289));
  xor_4  g08913(.A(new_n9289), .B(new_n9265), .Y(new_n9290));
  nand_5 g08914(.A(pi223), .B(pi081), .Y(new_n9291));
  xor_4  g08915(.A(new_n9291), .B(new_n9266), .Y(new_n9292));
  xnor_4 g08916(.A(new_n9292), .B(new_n9290), .Y(new_n9293));
  nand_5 g08917(.A(new_n9271), .B(new_n9264), .Y(new_n9294));
  nand_5 g08918(.A(new_n9272), .B(new_n9263), .Y(new_n9295));
  nand_5 g08919(.A(new_n9295), .B(new_n9294), .Y(new_n9296));
  nand_5 g08920(.A(pi233), .B(pi020), .Y(new_n9297));
  nand_5 g08921(.A(pi187), .B(pi160), .Y(new_n9298));
  xor_4  g08922(.A(new_n9298), .B(new_n9297), .Y(new_n9299));
  xor_4  g08923(.A(new_n9299), .B(new_n9257), .Y(new_n9300));
  xor_4  g08924(.A(new_n9300), .B(new_n9296), .Y(new_n9301));
  xnor_4 g08925(.A(new_n9301), .B(new_n9293), .Y(new_n9302));
  xor_4  g08926(.A(new_n9302), .B(new_n9286), .Y(new_n9303));
  xor_4  g08927(.A(new_n9303), .B(new_n9280), .Y(new_n9304));
  xor_4  g08928(.A(new_n9304), .B(new_n9279), .Y(new_n9305));
  not_8  g08929(.A(new_n9305), .Y(new_n9306));
  nor_5  g08930(.A(new_n9306), .B(new_n9203), .Y(new_n9307));
  xnor_4 g08931(.A(new_n9200), .B(new_n9199), .Y(new_n9308));
  xor_4  g08932(.A(new_n9276), .B(new_n9247), .Y(new_n9309));
  not_8  g08933(.A(new_n9309), .Y(new_n9310));
  nor_5  g08934(.A(new_n9310), .B(new_n9308), .Y(new_n9311));
  xnor_4 g08935(.A(new_n9190), .B(new_n9171), .Y(new_n9312));
  nand_5 g08936(.A(pi217), .B(pi160), .Y(new_n9313));
  xor_4  g08937(.A(new_n9172), .B(new_n9097), .Y(new_n9314));
  nor_5  g08938(.A(new_n9314), .B(new_n9313), .Y(new_n9315));
  xor_4  g08939(.A(new_n9239), .B(new_n9238), .Y(new_n9316));
  nor_5  g08940(.A(new_n9316), .B(new_n9315), .Y(new_n9317));
  not_8  g08941(.A(new_n9317), .Y(new_n9318));
  xor_4  g08942(.A(new_n9316), .B(new_n9315), .Y(new_n9319));
  xor_4  g08943(.A(new_n9179), .B(new_n9178), .Y(new_n9320));
  not_8  g08944(.A(new_n9320), .Y(new_n9321));
  nand_5 g08945(.A(new_n9321), .B(new_n9319), .Y(new_n9322));
  nand_5 g08946(.A(new_n9322), .B(new_n9318), .Y(new_n9323));
  xor_4  g08947(.A(new_n9240), .B(new_n9236), .Y(new_n9324));
  and_6  g08948(.A(new_n9324), .B(new_n9323), .Y(new_n9325));
  xnor_4 g08949(.A(new_n9188), .B(new_n9186), .Y(new_n9326));
  xor_4  g08950(.A(new_n9324), .B(new_n9323), .Y(new_n9327));
  and_6  g08951(.A(new_n9327), .B(new_n9326), .Y(new_n9328));
  nor_5  g08952(.A(new_n9328), .B(new_n9325), .Y(new_n9329));
  nor_5  g08953(.A(new_n9329), .B(new_n9312), .Y(new_n9330));
  xor_4  g08954(.A(new_n9242), .B(new_n9241), .Y(new_n9331));
  xnor_4 g08955(.A(new_n9329), .B(new_n9312), .Y(new_n9332));
  nor_5  g08956(.A(new_n9332), .B(new_n9331), .Y(new_n9333));
  or_6   g08957(.A(new_n9333), .B(new_n9330), .Y(new_n9334));
  xnor_4 g08958(.A(new_n9243), .B(new_n9235), .Y(new_n9335));
  nor_5  g08959(.A(new_n9335), .B(new_n9334), .Y(new_n9336));
  xor_4  g08960(.A(new_n9197), .B(new_n9196), .Y(new_n9337));
  xnor_4 g08961(.A(new_n9335), .B(new_n9334), .Y(new_n9338));
  nor_5  g08962(.A(new_n9338), .B(new_n9337), .Y(new_n9339));
  nor_5  g08963(.A(new_n9339), .B(new_n9336), .Y(new_n9340));
  xor_4  g08964(.A(new_n9309), .B(new_n9308), .Y(new_n9341));
  nor_5  g08965(.A(new_n9341), .B(new_n9340), .Y(new_n9342));
  nor_5  g08966(.A(new_n9342), .B(new_n9311), .Y(new_n9343));
  xor_4  g08967(.A(new_n9305), .B(new_n9203), .Y(new_n9344));
  nor_5  g08968(.A(new_n9344), .B(new_n9343), .Y(new_n9345));
  nor_5  g08969(.A(new_n9345), .B(new_n9307), .Y(new_n9346));
  or_6   g08970(.A(new_n8917), .B(new_n8901), .Y(new_n9347));
  nand_5 g08971(.A(new_n9347), .B(new_n8900), .Y(new_n9348));
  nor_5  g08972(.A(new_n9291), .B(new_n9267), .Y(new_n9349));
  nor_5  g08973(.A(new_n9292), .B(new_n9290), .Y(new_n9350));
  nor_5  g08974(.A(new_n9350), .B(new_n9349), .Y(new_n9351));
  nand_5 g08975(.A(pi191), .B(pi142), .Y(new_n9352));
  xor_4  g08976(.A(new_n9352), .B(new_n9351), .Y(new_n9353));
  nand_5 g08977(.A(new_n9300), .B(new_n9296), .Y(new_n9354));
  nand_5 g08978(.A(new_n9301), .B(new_n9293), .Y(new_n9355));
  nand_5 g08979(.A(new_n9355), .B(new_n9354), .Y(new_n9356));
  nand_5 g08980(.A(pi138), .B(pi017), .Y(new_n9357));
  not_8  g08981(.A(new_n9151), .Y(new_n9358));
  nor_5  g08982(.A(new_n9152), .B(new_n9358), .Y(new_n9359));
  not_8  g08983(.A(new_n9131), .Y(new_n9360));
  nor_5  g08984(.A(new_n9153), .B(new_n9360), .Y(new_n9361));
  nor_5  g08985(.A(new_n9361), .B(new_n9359), .Y(new_n9362));
  xor_4  g08986(.A(new_n9362), .B(new_n9357), .Y(new_n9363));
  xor_4  g08987(.A(new_n9363), .B(new_n9356), .Y(new_n9364));
  xor_4  g08988(.A(new_n9364), .B(new_n9353), .Y(new_n9365));
  xor_4  g08989(.A(new_n9365), .B(new_n9348), .Y(new_n9366));
  xor_4  g08990(.A(new_n9366), .B(new_n9346), .Y(new_n9367));
  not_8  g08991(.A(new_n9140), .Y(new_n9368));
  nor_5  g08992(.A(new_n9161), .B(new_n9368), .Y(new_n9369));
  nor_5  g08993(.A(new_n9162), .B(new_n9139), .Y(new_n9370));
  nor_5  g08994(.A(new_n9370), .B(new_n9369), .Y(new_n9371));
  nor_5  g08995(.A(new_n9163), .B(new_n9063), .Y(new_n9372));
  and_6  g08996(.A(new_n9202), .B(new_n9164), .Y(new_n9373));
  nor_5  g08997(.A(new_n9373), .B(new_n9372), .Y(new_n9374));
  xor_4  g08998(.A(new_n9374), .B(new_n9371), .Y(new_n9375));
  nand_5 g08999(.A(new_n9288), .B(new_n9287), .Y(new_n9376));
  nand_5 g09000(.A(new_n9289), .B(new_n9265), .Y(new_n9377));
  nand_5 g09001(.A(new_n9377), .B(new_n9376), .Y(new_n9378));
  nand_5 g09002(.A(pi223), .B(pi106), .Y(new_n9379));
  xor_4  g09003(.A(new_n9379), .B(new_n9378), .Y(new_n9380));
  not_8  g09004(.A(new_n9280), .Y(new_n9381));
  nand_5 g09005(.A(new_n9303), .B(new_n9381), .Y(new_n9382));
  not_8  g09006(.A(new_n9304), .Y(new_n9383));
  nand_5 g09007(.A(new_n9383), .B(new_n9279), .Y(new_n9384));
  nand_5 g09008(.A(new_n9384), .B(new_n9382), .Y(new_n9385));
  nand_5 g09009(.A(pi101), .B(pi081), .Y(new_n9386));
  nand_5 g09010(.A(pi177), .B(pi100), .Y(new_n9387));
  xor_4  g09011(.A(new_n9387), .B(new_n9386), .Y(new_n9388));
  nand_5 g09012(.A(pi249), .B(pi192), .Y(new_n9389));
  or_6   g09013(.A(new_n9159), .B(new_n9133), .Y(new_n9390));
  not_8  g09014(.A(new_n9160), .Y(new_n9391));
  nand_5 g09015(.A(new_n9391), .B(new_n9156), .Y(new_n9392));
  nand_5 g09016(.A(new_n9392), .B(new_n9390), .Y(new_n9393));
  nand_5 g09017(.A(pi251), .B(pi222), .Y(new_n9394));
  xor_4  g09018(.A(new_n9394), .B(new_n9393), .Y(new_n9395));
  nand_5 g09019(.A(new_n9298), .B(new_n9297), .Y(new_n9396));
  nand_5 g09020(.A(new_n9299), .B(new_n9257), .Y(new_n9397));
  nand_5 g09021(.A(new_n9397), .B(new_n9396), .Y(new_n9398));
  xor_4  g09022(.A(new_n9398), .B(new_n9395), .Y(new_n9399));
  xor_4  g09023(.A(new_n9399), .B(new_n9389), .Y(new_n9400));
  xnor_4 g09024(.A(new_n9400), .B(new_n9388), .Y(new_n9401));
  xor_4  g09025(.A(new_n9401), .B(new_n9385), .Y(new_n9402));
  xor_4  g09026(.A(new_n9402), .B(new_n9380), .Y(new_n9403));
  xor_4  g09027(.A(new_n9403), .B(new_n9375), .Y(new_n9404));
  xor_4  g09028(.A(new_n9404), .B(new_n9367), .Y(new_n9405));
  nand_5 g09029(.A(pi233), .B(pi060), .Y(new_n9406));
  nand_5 g09030(.A(pi087), .B(pi082), .Y(new_n9407));
  not_8  g09031(.A(new_n8893), .Y(new_n9408));
  nor_5  g09032(.A(new_n8918), .B(new_n9408), .Y(new_n9409));
  nor_5  g09033(.A(new_n8919), .B(new_n8892), .Y(new_n9410));
  nor_5  g09034(.A(new_n9410), .B(new_n9409), .Y(new_n9411));
  xor_4  g09035(.A(new_n9411), .B(new_n9407), .Y(new_n9412));
  xor_4  g09036(.A(new_n9412), .B(new_n9406), .Y(new_n9413));
  nor_5  g09037(.A(new_n8951), .B(new_n8946), .Y(new_n9414));
  not_8  g09038(.A(new_n8930), .Y(new_n9415));
  nor_5  g09039(.A(new_n8952), .B(new_n9415), .Y(new_n9416));
  nor_5  g09040(.A(new_n9416), .B(new_n9414), .Y(new_n9417));
  nand_5 g09041(.A(pi102), .B(pi005), .Y(new_n9418));
  xor_4  g09042(.A(new_n9418), .B(new_n9417), .Y(new_n9419));
  nand_5 g09043(.A(pi232), .B(pi071), .Y(new_n9420));
  xor_4  g09044(.A(new_n9420), .B(new_n9419), .Y(new_n9421));
  xor_4  g09045(.A(new_n9421), .B(new_n9413), .Y(new_n9422));
  xor_4  g09046(.A(new_n9422), .B(new_n9405), .Y(new_n9423));
  nand_5 g09047(.A(pi231), .B(pi001), .Y(new_n9424));
  not_8  g09048(.A(new_n9022), .Y(new_n9425));
  nand_5 g09049(.A(new_n9425), .B(new_n8920), .Y(new_n9426));
  or_6   g09050(.A(new_n9062), .B(new_n9023), .Y(new_n9427));
  nand_5 g09051(.A(new_n9427), .B(new_n9426), .Y(new_n9428));
  nand_5 g09052(.A(new_n9283), .B(new_n9258), .Y(new_n9429));
  not_8  g09053(.A(new_n9286), .Y(new_n9430));
  nand_5 g09054(.A(new_n9302), .B(new_n9430), .Y(new_n9431));
  nand_5 g09055(.A(new_n9431), .B(new_n9429), .Y(new_n9432));
  xor_4  g09056(.A(new_n9432), .B(new_n9428), .Y(new_n9433));
  xor_4  g09057(.A(new_n9433), .B(new_n9424), .Y(new_n9434));
  nand_5 g09058(.A(new_n8923), .B(new_n8922), .Y(new_n9435));
  nand_5 g09059(.A(new_n8924), .B(new_n8921), .Y(new_n9436));
  nand_5 g09060(.A(new_n9436), .B(new_n9435), .Y(new_n9437));
  not_8  g09061(.A(new_n9150), .Y(new_n9438));
  nor_5  g09062(.A(new_n9154), .B(new_n9438), .Y(new_n9439));
  nor_5  g09063(.A(new_n9155), .B(new_n9147), .Y(new_n9440));
  nor_5  g09064(.A(new_n9440), .B(new_n9439), .Y(new_n9441));
  xor_4  g09065(.A(new_n9441), .B(new_n9437), .Y(new_n9442));
  xor_4  g09066(.A(new_n9442), .B(new_n9434), .Y(new_n9443));
  nand_5 g09067(.A(new_n9142), .B(new_n9141), .Y(new_n9444));
  nand_5 g09068(.A(new_n9143), .B(new_n9119), .Y(new_n9445));
  nand_5 g09069(.A(new_n9445), .B(new_n9444), .Y(new_n9446));
  nor_5  g09070(.A(new_n9145), .B(new_n9121), .Y(new_n9447));
  nor_5  g09071(.A(new_n9146), .B(new_n9144), .Y(new_n9448));
  nor_5  g09072(.A(new_n9448), .B(new_n9447), .Y(new_n9449));
  nand_5 g09073(.A(pi174), .B(pi041), .Y(new_n9450));
  nand_5 g09074(.A(pi216), .B(pi040), .Y(new_n9451));
  nand_5 g09075(.A(pi125), .B(pi079), .Y(new_n9452));
  xnor_4 g09076(.A(new_n9452), .B(new_n9451), .Y(new_n9453));
  xor_4  g09077(.A(new_n9453), .B(new_n9450), .Y(new_n9454));
  nand_5 g09078(.A(pi176), .B(pi076), .Y(new_n9455));
  nand_5 g09079(.A(pi182), .B(pi157), .Y(new_n9456));
  nand_5 g09080(.A(pi024), .B(pi023), .Y(new_n9457));
  nand_5 g09081(.A(pi155), .B(pi111), .Y(new_n9458));
  xor_4  g09082(.A(new_n9458), .B(new_n9457), .Y(new_n9459));
  xor_4  g09083(.A(new_n9459), .B(new_n9456), .Y(new_n9460));
  xor_4  g09084(.A(new_n9460), .B(new_n9455), .Y(new_n9461));
  xor_4  g09085(.A(new_n9461), .B(new_n9454), .Y(new_n9462));
  nand_5 g09086(.A(pi255), .B(pi123), .Y(new_n9463));
  nand_5 g09087(.A(new_n8915), .B(new_n8911), .Y(new_n9464));
  not_8  g09088(.A(new_n8908), .Y(new_n9465));
  nand_5 g09089(.A(new_n8916), .B(new_n9465), .Y(new_n9466));
  nand_5 g09090(.A(new_n9466), .B(new_n9464), .Y(new_n9467));
  nand_5 g09091(.A(pi227), .B(pi225), .Y(new_n9468));
  nand_5 g09092(.A(pi187), .B(pi020), .Y(new_n9469));
  xor_4  g09093(.A(new_n9469), .B(new_n9468), .Y(new_n9470));
  xor_4  g09094(.A(new_n9470), .B(new_n9467), .Y(new_n9471));
  xor_4  g09095(.A(new_n9471), .B(new_n9463), .Y(new_n9472));
  xor_4  g09096(.A(new_n9472), .B(new_n9462), .Y(new_n9473));
  xor_4  g09097(.A(new_n9473), .B(new_n9449), .Y(new_n9474));
  xor_4  g09098(.A(new_n9474), .B(new_n9446), .Y(new_n9475));
  xor_4  g09099(.A(new_n9475), .B(new_n9443), .Y(new_n9476));
  nand_5 g09100(.A(pi210), .B(pi086), .Y(new_n9477));
  nor_5  g09101(.A(new_n8906), .B(new_n8884), .Y(new_n9478));
  nor_5  g09102(.A(new_n8907), .B(new_n8905), .Y(new_n9479));
  or_6   g09103(.A(new_n9479), .B(new_n9478), .Y(new_n9480));
  nor_5  g09104(.A(new_n8931), .B(new_n8926), .Y(new_n9481));
  nor_5  g09105(.A(new_n8929), .B(new_n8925), .Y(new_n9482));
  nor_5  g09106(.A(new_n9482), .B(new_n9481), .Y(new_n9483));
  nand_5 g09107(.A(pi122), .B(pi121), .Y(new_n9484));
  nand_5 g09108(.A(pi140), .B(pi059), .Y(new_n9485));
  xor_4  g09109(.A(new_n9485), .B(new_n9484), .Y(new_n9486));
  xor_4  g09110(.A(new_n9486), .B(new_n9483), .Y(new_n9487));
  nand_5 g09111(.A(pi217), .B(pi137), .Y(new_n9488));
  nand_5 g09112(.A(new_n8903), .B(new_n8882), .Y(new_n9489));
  nand_5 g09113(.A(new_n8904), .B(new_n8902), .Y(new_n9490));
  nand_5 g09114(.A(new_n9490), .B(new_n9489), .Y(new_n9491));
  xnor_4 g09115(.A(new_n9491), .B(new_n9488), .Y(new_n9492));
  nand_5 g09116(.A(pi224), .B(pi099), .Y(new_n9493));
  nand_5 g09117(.A(pi219), .B(pi021), .Y(new_n9494));
  xor_4  g09118(.A(new_n9494), .B(new_n9493), .Y(new_n9495));
  xor_4  g09119(.A(new_n9495), .B(new_n9492), .Y(new_n9496));
  or_6   g09120(.A(new_n9021), .B(new_n8979), .Y(new_n9497));
  nand_5 g09121(.A(new_n9497), .B(new_n9020), .Y(new_n9498));
  nand_5 g09122(.A(new_n8913), .B(new_n8912), .Y(new_n9499));
  nand_5 g09123(.A(new_n8914), .B(new_n8872), .Y(new_n9500));
  nand_5 g09124(.A(new_n9500), .B(new_n9499), .Y(new_n9501));
  nand_5 g09125(.A(pi169), .B(pi127), .Y(new_n9502));
  xnor_4 g09126(.A(new_n9502), .B(new_n9501), .Y(new_n9503));
  xor_4  g09127(.A(new_n9503), .B(new_n9498), .Y(new_n9504));
  nand_5 g09128(.A(pi242), .B(pi094), .Y(new_n9505));
  nand_5 g09129(.A(pi160), .B(pi129), .Y(new_n9506));
  xor_4  g09130(.A(new_n9506), .B(new_n9505), .Y(new_n9507));
  nand_5 g09131(.A(new_n8949), .B(new_n8948), .Y(new_n9508));
  nand_5 g09132(.A(new_n8950), .B(new_n8947), .Y(new_n9509));
  nand_5 g09133(.A(new_n9509), .B(new_n9508), .Y(new_n9510));
  nand_5 g09134(.A(pi252), .B(pi135), .Y(new_n9511));
  xor_4  g09135(.A(new_n9511), .B(new_n9510), .Y(new_n9512));
  nand_5 g09136(.A(new_n8976), .B(new_n8955), .Y(new_n9513));
  nand_5 g09137(.A(new_n8977), .B(new_n8953), .Y(new_n9514));
  nand_5 g09138(.A(new_n9514), .B(new_n9513), .Y(new_n9515));
  xor_4  g09139(.A(new_n9515), .B(new_n9512), .Y(new_n9516));
  xor_4  g09140(.A(new_n9516), .B(new_n9507), .Y(new_n9517));
  xor_4  g09141(.A(new_n9517), .B(new_n9504), .Y(new_n9518));
  xor_4  g09142(.A(new_n9518), .B(new_n9496), .Y(new_n9519));
  xor_4  g09143(.A(new_n9519), .B(new_n9487), .Y(new_n9520));
  xor_4  g09144(.A(new_n9520), .B(new_n9480), .Y(new_n9521));
  xor_4  g09145(.A(new_n9521), .B(new_n9477), .Y(new_n9522));
  xor_4  g09146(.A(new_n9522), .B(new_n9476), .Y(new_n9523));
  xor_4  g09147(.A(new_n9523), .B(new_n9423), .Y(po051));
  xor_4  g09148(.A(new_n3277), .B(new_n3272), .Y(po052));
  xor_4  g09149(.A(new_n3530), .B(new_n3521), .Y(po053));
  xor_4  g09150(.A(new_n876), .B(new_n419), .Y(po054));
  xor_4  g09151(.A(new_n7919), .B(new_n7904), .Y(po055));
  xor_4  g09152(.A(new_n4247), .B(new_n4246), .Y(po056));
  xor_4  g09153(.A(new_n1304), .B(new_n1302), .Y(po057));
  xor_4  g09154(.A(new_n4234), .B(new_n4233), .Y(po058));
  xnor_4 g09155(.A(new_n5437), .B(new_n5436), .Y(po059));
  nor_5  g09156(.A(new_n2586), .B(new_n2584), .Y(new_n9533));
  xor_4  g09157(.A(new_n9533), .B(new_n2581), .Y(po060));
  xor_4  g09158(.A(new_n2576), .B(new_n2575), .Y(po061));
  and_6  g09159(.A(new_n8811), .B(new_n8743), .Y(new_n9536));
  nor_5  g09160(.A(new_n8815), .B(new_n8812), .Y(new_n9537));
  nor_5  g09161(.A(new_n9537), .B(new_n9536), .Y(new_n9538));
  not_8  g09162(.A(new_n8724), .Y(new_n9539));
  nand_5 g09163(.A(new_n8742), .B(new_n9539), .Y(new_n9540));
  nand_5 g09164(.A(pi233), .B(pi131), .Y(new_n9541));
  xor_4  g09165(.A(new_n9541), .B(new_n9540), .Y(new_n9542));
  not_8  g09166(.A(new_n8740), .Y(new_n9543));
  nor_5  g09167(.A(new_n9543), .B(new_n8736), .Y(new_n9544));
  nor_5  g09168(.A(new_n8741), .B(new_n8735), .Y(new_n9545));
  nor_5  g09169(.A(new_n9545), .B(new_n9544), .Y(new_n9546));
  nand_5 g09170(.A(new_n8733), .B(new_n8730), .Y(new_n9547));
  nand_5 g09171(.A(new_n8734), .B(new_n8729), .Y(new_n9548));
  nand_5 g09172(.A(new_n9548), .B(new_n9547), .Y(new_n9549));
  nand_5 g09173(.A(pi106), .B(pi077), .Y(new_n9550));
  nor_5  g09174(.A(new_n9550), .B(new_n8730), .Y(new_n9551));
  not_8  g09175(.A(new_n9551), .Y(new_n9552));
  nand_5 g09176(.A(pi081), .B(pi077), .Y(new_n9553));
  nand_5 g09177(.A(pi106), .B(pi052), .Y(new_n9554));
  nand_5 g09178(.A(new_n9554), .B(new_n9553), .Y(new_n9555));
  nand_5 g09179(.A(new_n9555), .B(new_n9552), .Y(new_n9556));
  nand_5 g09180(.A(pi227), .B(pi133), .Y(new_n9557));
  nand_5 g09181(.A(new_n8727), .B(new_n8726), .Y(new_n9558));
  nand_5 g09182(.A(new_n8728), .B(new_n8725), .Y(new_n9559));
  nand_5 g09183(.A(new_n9559), .B(new_n9558), .Y(new_n9560));
  nand_5 g09184(.A(pi100), .B(pi064), .Y(new_n9561));
  nor_5  g09185(.A(new_n9561), .B(new_n8726), .Y(new_n9562));
  not_8  g09186(.A(new_n9562), .Y(new_n9563));
  nand_5 g09187(.A(pi189), .B(pi100), .Y(new_n9564));
  nand_5 g09188(.A(pi217), .B(pi064), .Y(new_n9565));
  nand_5 g09189(.A(new_n9565), .B(new_n9564), .Y(new_n9566));
  nand_5 g09190(.A(new_n9566), .B(new_n9563), .Y(new_n9567));
  xor_4  g09191(.A(new_n9567), .B(new_n9560), .Y(new_n9568));
  xor_4  g09192(.A(new_n9568), .B(new_n9557), .Y(new_n9569));
  xor_4  g09193(.A(new_n9569), .B(new_n9556), .Y(new_n9570));
  xor_4  g09194(.A(new_n9570), .B(new_n9549), .Y(new_n9571));
  not_8  g09195(.A(new_n9571), .Y(new_n9572));
  xor_4  g09196(.A(new_n9572), .B(new_n9546), .Y(new_n9573));
  xor_4  g09197(.A(new_n9573), .B(new_n9542), .Y(new_n9574));
  not_8  g09198(.A(new_n9574), .Y(new_n9575));
  nand_5 g09199(.A(new_n9575), .B(new_n9538), .Y(new_n9576));
  or_6   g09200(.A(new_n8809), .B(new_n8805), .Y(new_n9577));
  nand_5 g09201(.A(new_n8810), .B(new_n8786), .Y(new_n9578));
  nand_5 g09202(.A(new_n9578), .B(new_n9577), .Y(new_n9579));
  not_8  g09203(.A(new_n8787), .Y(new_n9580));
  nor_5  g09204(.A(new_n8804), .B(new_n9580), .Y(new_n9581));
  nand_5 g09205(.A(pi174), .B(pi168), .Y(new_n9582));
  or_6   g09206(.A(new_n8802), .B(new_n8799), .Y(new_n9583));
  not_8  g09207(.A(new_n8798), .Y(new_n9584));
  nand_5 g09208(.A(new_n8803), .B(new_n9584), .Y(new_n9585));
  nand_5 g09209(.A(new_n9585), .B(new_n9583), .Y(new_n9586));
  nand_5 g09210(.A(pi125), .B(pi035), .Y(new_n9587));
  nand_5 g09211(.A(new_n8789), .B(new_n8788), .Y(new_n9588));
  nand_5 g09212(.A(new_n8791), .B(new_n8790), .Y(new_n9589));
  nand_5 g09213(.A(new_n9589), .B(new_n9588), .Y(new_n9590));
  nand_5 g09214(.A(pi249), .B(pi204), .Y(new_n9591));
  nand_5 g09215(.A(pi222), .B(pi015), .Y(new_n9592));
  nand_5 g09216(.A(new_n9592), .B(new_n9591), .Y(new_n9593));
  nand_5 g09217(.A(pi222), .B(pi204), .Y(new_n9594));
  nor_5  g09218(.A(new_n9594), .B(new_n8791), .Y(new_n9595));
  not_8  g09219(.A(new_n9595), .Y(new_n9596));
  nand_5 g09220(.A(new_n9596), .B(new_n9593), .Y(new_n9597));
  xor_4  g09221(.A(new_n9597), .B(new_n9590), .Y(new_n9598));
  xor_4  g09222(.A(new_n9598), .B(new_n9587), .Y(new_n9599));
  nand_5 g09223(.A(new_n8796), .B(new_n8793), .Y(new_n9600));
  nand_5 g09224(.A(new_n8797), .B(new_n8792), .Y(new_n9601));
  nand_5 g09225(.A(new_n9601), .B(new_n9600), .Y(new_n9602));
  xor_4  g09226(.A(new_n9602), .B(new_n9599), .Y(new_n9603));
  nand_5 g09227(.A(pi176), .B(pi139), .Y(new_n9604));
  nand_5 g09228(.A(pi208), .B(pi040), .Y(new_n9605));
  nand_5 g09229(.A(new_n9605), .B(new_n9604), .Y(new_n9606));
  nand_5 g09230(.A(pi139), .B(pi040), .Y(new_n9607));
  nor_5  g09231(.A(new_n9607), .B(new_n8793), .Y(new_n9608));
  not_8  g09232(.A(new_n9608), .Y(new_n9609));
  nand_5 g09233(.A(new_n9609), .B(new_n9606), .Y(new_n9610));
  xor_4  g09234(.A(new_n9610), .B(new_n9603), .Y(new_n9611));
  xor_4  g09235(.A(new_n9611), .B(new_n9586), .Y(new_n9612));
  xor_4  g09236(.A(new_n9612), .B(new_n9582), .Y(new_n9613));
  xnor_4 g09237(.A(new_n9613), .B(new_n9581), .Y(new_n9614));
  xor_4  g09238(.A(new_n9614), .B(new_n9579), .Y(new_n9615));
  nand_5 g09239(.A(new_n8784), .B(new_n8782), .Y(new_n9616));
  nand_5 g09240(.A(new_n8785), .B(new_n8763), .Y(new_n9617));
  and_6  g09241(.A(new_n9617), .B(new_n9616), .Y(new_n9618));
  nand_5 g09242(.A(new_n8773), .B(new_n8770), .Y(new_n9619));
  nand_5 g09243(.A(new_n8774), .B(new_n8769), .Y(new_n9620));
  nand_5 g09244(.A(new_n9620), .B(new_n9619), .Y(new_n9621));
  nand_5 g09245(.A(pi224), .B(pi104), .Y(new_n9622));
  nand_5 g09246(.A(pi255), .B(pi212), .Y(new_n9623));
  nand_5 g09247(.A(new_n9623), .B(new_n9622), .Y(new_n9624));
  nand_5 g09248(.A(pi255), .B(pi104), .Y(new_n9625));
  or_6   g09249(.A(new_n9625), .B(new_n8770), .Y(new_n9626));
  nand_5 g09250(.A(new_n9626), .B(new_n9624), .Y(new_n9627));
  nand_5 g09251(.A(pi024), .B(pi013), .Y(new_n9628));
  nand_5 g09252(.A(new_n8767), .B(new_n8766), .Y(new_n9629));
  nand_5 g09253(.A(new_n8768), .B(new_n8765), .Y(new_n9630));
  nand_5 g09254(.A(new_n9630), .B(new_n9629), .Y(new_n9631));
  nand_5 g09255(.A(pi112), .B(pi111), .Y(new_n9632));
  nand_5 g09256(.A(pi210), .B(pi105), .Y(new_n9633));
  nand_5 g09257(.A(new_n9633), .B(new_n9632), .Y(new_n9634));
  nand_5 g09258(.A(pi111), .B(pi105), .Y(new_n9635));
  nor_5  g09259(.A(new_n9635), .B(new_n8767), .Y(new_n9636));
  not_8  g09260(.A(new_n9636), .Y(new_n9637));
  nand_5 g09261(.A(new_n9637), .B(new_n9634), .Y(new_n9638));
  xor_4  g09262(.A(new_n9638), .B(new_n9631), .Y(new_n9639));
  xor_4  g09263(.A(new_n9639), .B(new_n9628), .Y(new_n9640));
  xor_4  g09264(.A(new_n9640), .B(new_n9627), .Y(new_n9641));
  xor_4  g09265(.A(new_n9641), .B(new_n9621), .Y(new_n9642));
  nor_5  g09266(.A(new_n8779), .B(new_n8776), .Y(new_n9643));
  not_8  g09267(.A(new_n8775), .Y(new_n9644));
  and_6  g09268(.A(new_n8780), .B(new_n9644), .Y(new_n9645));
  nor_5  g09269(.A(new_n9645), .B(new_n9643), .Y(new_n9646));
  xnor_4 g09270(.A(new_n9646), .B(new_n9642), .Y(new_n9647));
  nor_5  g09271(.A(new_n8781), .B(new_n8764), .Y(new_n9648));
  nand_5 g09272(.A(pi213), .B(pi127), .Y(new_n9649));
  xor_4  g09273(.A(new_n9649), .B(new_n9648), .Y(new_n9650));
  xor_4  g09274(.A(new_n9650), .B(new_n9647), .Y(new_n9651));
  not_8  g09275(.A(new_n8762), .Y(new_n9652));
  nor_5  g09276(.A(new_n9652), .B(new_n8744), .Y(new_n9653));
  nand_5 g09277(.A(pi236), .B(pi005), .Y(new_n9654));
  nand_5 g09278(.A(new_n8759), .B(new_n8755), .Y(new_n9655));
  nand_5 g09279(.A(new_n8760), .B(new_n8754), .Y(new_n9656));
  nand_5 g09280(.A(new_n9656), .B(new_n9655), .Y(new_n9657));
  nand_5 g09281(.A(pi161), .B(pi121), .Y(new_n9658));
  nand_5 g09282(.A(pi241), .B(pi231), .Y(new_n9659));
  and_6  g09283(.A(new_n9659), .B(new_n9658), .Y(new_n9660));
  nand_5 g09284(.A(pi231), .B(pi161), .Y(new_n9661));
  nor_5  g09285(.A(new_n9661), .B(new_n8755), .Y(new_n9662));
  or_6   g09286(.A(new_n9662), .B(new_n9660), .Y(new_n9663));
  nand_5 g09287(.A(new_n8752), .B(new_n8751), .Y(new_n9664));
  nand_5 g09288(.A(new_n8753), .B(new_n8750), .Y(new_n9665));
  nand_5 g09289(.A(new_n9665), .B(new_n9664), .Y(new_n9666));
  nand_5 g09290(.A(pi252), .B(pi141), .Y(new_n9667));
  nand_5 g09291(.A(pi140), .B(pi090), .Y(new_n9668));
  nand_5 g09292(.A(pi242), .B(pi047), .Y(new_n9669));
  nand_5 g09293(.A(new_n9669), .B(new_n9668), .Y(new_n9670));
  nand_5 g09294(.A(pi140), .B(pi047), .Y(new_n9671));
  nor_5  g09295(.A(new_n9671), .B(new_n8751), .Y(new_n9672));
  not_8  g09296(.A(new_n9672), .Y(new_n9673));
  nand_5 g09297(.A(new_n9673), .B(new_n9670), .Y(new_n9674));
  xor_4  g09298(.A(new_n9674), .B(new_n9667), .Y(new_n9675));
  xor_4  g09299(.A(new_n9675), .B(new_n9666), .Y(new_n9676));
  xor_4  g09300(.A(new_n9676), .B(new_n9663), .Y(new_n9677));
  xor_4  g09301(.A(new_n9677), .B(new_n9657), .Y(new_n9678));
  nor_5  g09302(.A(new_n8748), .B(new_n8745), .Y(new_n9679));
  and_6  g09303(.A(new_n8761), .B(new_n8749), .Y(new_n9680));
  nor_5  g09304(.A(new_n9680), .B(new_n9679), .Y(new_n9681));
  xnor_4 g09305(.A(new_n9681), .B(new_n9678), .Y(new_n9682));
  xnor_4 g09306(.A(new_n9682), .B(new_n9654), .Y(new_n9683));
  xor_4  g09307(.A(new_n9683), .B(new_n9653), .Y(new_n9684));
  xor_4  g09308(.A(new_n9684), .B(new_n9651), .Y(new_n9685));
  xnor_4 g09309(.A(new_n9685), .B(new_n9618), .Y(new_n9686));
  xnor_4 g09310(.A(new_n9686), .B(new_n9615), .Y(new_n9687));
  xor_4  g09311(.A(new_n9575), .B(new_n9538), .Y(new_n9688));
  nand_5 g09312(.A(new_n9688), .B(new_n9687), .Y(new_n9689));
  nand_5 g09313(.A(new_n9689), .B(new_n9576), .Y(new_n9690));
  nor_5  g09314(.A(new_n9682), .B(new_n9654), .Y(new_n9691));
  not_8  g09315(.A(new_n9691), .Y(new_n9692));
  not_8  g09316(.A(new_n9653), .Y(new_n9693));
  or_6   g09317(.A(new_n9683), .B(new_n9693), .Y(new_n9694));
  nand_5 g09318(.A(new_n9694), .B(new_n9692), .Y(new_n9695));
  or_6   g09319(.A(new_n9681), .B(new_n9678), .Y(new_n9696));
  not_8  g09320(.A(new_n9677), .Y(new_n9697));
  nor_5  g09321(.A(new_n9697), .B(new_n9657), .Y(new_n9698));
  nand_5 g09322(.A(new_n9698), .B(new_n9662), .Y(new_n9699));
  nor_5  g09323(.A(new_n9676), .B(new_n9663), .Y(new_n9700));
  nor_5  g09324(.A(new_n9700), .B(new_n9662), .Y(new_n9701));
  not_8  g09325(.A(new_n9701), .Y(new_n9702));
  nor_5  g09326(.A(new_n9702), .B(new_n9698), .Y(new_n9703));
  not_8  g09327(.A(new_n9703), .Y(new_n9704));
  nand_5 g09328(.A(new_n9704), .B(new_n9699), .Y(new_n9705));
  nand_5 g09329(.A(pi141), .B(pi121), .Y(new_n9706));
  xor_4  g09330(.A(new_n9706), .B(new_n9672), .Y(new_n9707));
  nand_5 g09331(.A(pi242), .B(pi018), .Y(new_n9708));
  nand_5 g09332(.A(pi252), .B(pi090), .Y(new_n9709));
  xor_4  g09333(.A(new_n9709), .B(new_n9708), .Y(new_n9710));
  xor_4  g09334(.A(new_n9710), .B(new_n9671), .Y(new_n9711));
  xor_4  g09335(.A(new_n9711), .B(new_n9707), .Y(new_n9712));
  nand_5 g09336(.A(new_n9674), .B(new_n9667), .Y(new_n9713));
  nand_5 g09337(.A(new_n9675), .B(new_n9666), .Y(new_n9714));
  nand_5 g09338(.A(new_n9714), .B(new_n9713), .Y(new_n9715));
  nand_5 g09339(.A(pi236), .B(pi021), .Y(new_n9716));
  nand_5 g09340(.A(pi241), .B(pi005), .Y(new_n9717));
  xor_4  g09341(.A(new_n9717), .B(new_n9716), .Y(new_n9718));
  xor_4  g09342(.A(new_n9718), .B(new_n9661), .Y(new_n9719));
  xnor_4 g09343(.A(new_n9719), .B(new_n9715), .Y(new_n9720));
  xor_4  g09344(.A(new_n9720), .B(new_n9712), .Y(new_n9721));
  not_8  g09345(.A(new_n9721), .Y(new_n9722));
  xor_4  g09346(.A(new_n9722), .B(new_n9705), .Y(new_n9723));
  xor_4  g09347(.A(new_n9723), .B(new_n9696), .Y(new_n9724));
  xor_4  g09348(.A(new_n9724), .B(new_n9695), .Y(new_n9725));
  not_8  g09349(.A(new_n9649), .Y(new_n9726));
  nor_5  g09350(.A(new_n9726), .B(new_n9648), .Y(new_n9727));
  not_8  g09351(.A(new_n9647), .Y(new_n9728));
  nor_5  g09352(.A(new_n9650), .B(new_n9728), .Y(new_n9729));
  nor_5  g09353(.A(new_n9729), .B(new_n9727), .Y(new_n9730));
  nor_5  g09354(.A(new_n9646), .B(new_n9642), .Y(new_n9731));
  nand_5 g09355(.A(new_n9640), .B(new_n9627), .Y(new_n9732));
  nand_5 g09356(.A(new_n9641), .B(new_n9621), .Y(new_n9733));
  nand_5 g09357(.A(new_n9733), .B(new_n9732), .Y(new_n9734));
  xor_4  g09358(.A(new_n9734), .B(new_n9626), .Y(new_n9735));
  nand_5 g09359(.A(pi224), .B(pi013), .Y(new_n9736));
  xor_4  g09360(.A(new_n9736), .B(new_n9636), .Y(new_n9737));
  nand_5 g09361(.A(pi210), .B(pi183), .Y(new_n9738));
  nand_5 g09362(.A(pi112), .B(pi024), .Y(new_n9739));
  xor_4  g09363(.A(new_n9739), .B(new_n9738), .Y(new_n9740));
  xor_4  g09364(.A(new_n9740), .B(new_n9635), .Y(new_n9741));
  xor_4  g09365(.A(new_n9741), .B(new_n9737), .Y(new_n9742));
  nand_5 g09366(.A(new_n9638), .B(new_n9631), .Y(new_n9743));
  nand_5 g09367(.A(new_n9639), .B(new_n9628), .Y(new_n9744));
  nand_5 g09368(.A(new_n9744), .B(new_n9743), .Y(new_n9745));
  nand_5 g09369(.A(pi212), .B(pi127), .Y(new_n9746));
  nand_5 g09370(.A(pi232), .B(pi213), .Y(new_n9747));
  xor_4  g09371(.A(new_n9747), .B(new_n9746), .Y(new_n9748));
  xor_4  g09372(.A(new_n9748), .B(new_n9625), .Y(new_n9749));
  xor_4  g09373(.A(new_n9749), .B(new_n9745), .Y(new_n9750));
  xor_4  g09374(.A(new_n9750), .B(new_n9742), .Y(new_n9751));
  xor_4  g09375(.A(new_n9751), .B(new_n9735), .Y(new_n9752));
  and_6  g09376(.A(new_n9752), .B(new_n9731), .Y(new_n9753));
  nor_5  g09377(.A(new_n9752), .B(new_n9731), .Y(new_n9754));
  or_6   g09378(.A(new_n9754), .B(new_n9753), .Y(new_n9755));
  xnor_4 g09379(.A(new_n9755), .B(new_n9730), .Y(new_n9756));
  xor_4  g09380(.A(new_n9756), .B(new_n9725), .Y(new_n9757));
  not_8  g09381(.A(new_n9651), .Y(new_n9758));
  nand_5 g09382(.A(new_n9684), .B(new_n9758), .Y(new_n9759));
  or_6   g09383(.A(new_n9685), .B(new_n9618), .Y(new_n9760));
  nand_5 g09384(.A(new_n9760), .B(new_n9759), .Y(new_n9761));
  xor_4  g09385(.A(new_n9761), .B(new_n9757), .Y(new_n9762));
  nor_5  g09386(.A(new_n9612), .B(new_n9582), .Y(new_n9763));
  nand_5 g09387(.A(new_n9613), .B(new_n9581), .Y(new_n9764));
  not_8  g09388(.A(new_n9764), .Y(new_n9765));
  nor_5  g09389(.A(new_n9765), .B(new_n9763), .Y(new_n9766));
  not_8  g09390(.A(new_n9611), .Y(new_n9767));
  nand_5 g09391(.A(new_n9767), .B(new_n9586), .Y(new_n9768));
  nand_5 g09392(.A(pi208), .B(pi174), .Y(new_n9769));
  nand_5 g09393(.A(pi168), .B(pi157), .Y(new_n9770));
  xor_4  g09394(.A(new_n9770), .B(new_n9769), .Y(new_n9771));
  xor_4  g09395(.A(new_n9771), .B(new_n9607), .Y(new_n9772));
  nand_5 g09396(.A(new_n9597), .B(new_n9590), .Y(new_n9773));
  nand_5 g09397(.A(new_n9598), .B(new_n9587), .Y(new_n9774));
  nand_5 g09398(.A(new_n9774), .B(new_n9773), .Y(new_n9775));
  xor_4  g09399(.A(new_n9775), .B(new_n9772), .Y(new_n9776));
  nand_5 g09400(.A(pi176), .B(pi035), .Y(new_n9777));
  xor_4  g09401(.A(new_n9777), .B(new_n9595), .Y(new_n9778));
  nand_5 g09402(.A(pi249), .B(pi146), .Y(new_n9779));
  nand_5 g09403(.A(pi125), .B(pi015), .Y(new_n9780));
  xor_4  g09404(.A(new_n9780), .B(new_n9779), .Y(new_n9781));
  xor_4  g09405(.A(new_n9781), .B(new_n9594), .Y(new_n9782));
  xor_4  g09406(.A(new_n9782), .B(new_n9778), .Y(new_n9783));
  xor_4  g09407(.A(new_n9783), .B(new_n9776), .Y(new_n9784));
  nor_5  g09408(.A(new_n9602), .B(new_n9599), .Y(new_n9785));
  xor_4  g09409(.A(new_n9609), .B(new_n9785), .Y(new_n9786));
  nand_5 g09410(.A(new_n9606), .B(new_n9603), .Y(new_n9787));
  nand_5 g09411(.A(new_n9787), .B(new_n9786), .Y(new_n9788));
  xor_4  g09412(.A(new_n9788), .B(new_n9784), .Y(new_n9789));
  not_8  g09413(.A(new_n9789), .Y(new_n9790));
  xor_4  g09414(.A(new_n9790), .B(new_n9768), .Y(new_n9791));
  xor_4  g09415(.A(new_n9791), .B(new_n9766), .Y(new_n9792));
  not_8  g09416(.A(new_n9614), .Y(new_n9793));
  nor_5  g09417(.A(new_n9793), .B(new_n9579), .Y(new_n9794));
  nor_5  g09418(.A(new_n9686), .B(new_n9615), .Y(new_n9795));
  nor_5  g09419(.A(new_n9795), .B(new_n9794), .Y(new_n9796));
  xor_4  g09420(.A(new_n9796), .B(new_n9792), .Y(new_n9797));
  xnor_4 g09421(.A(new_n9797), .B(new_n9762), .Y(new_n9798));
  not_8  g09422(.A(new_n9546), .Y(new_n9799));
  nand_5 g09423(.A(new_n9572), .B(new_n9799), .Y(new_n9800));
  nand_5 g09424(.A(new_n9541), .B(new_n9540), .Y(new_n9801));
  nand_5 g09425(.A(new_n9573), .B(new_n9542), .Y(new_n9802));
  nand_5 g09426(.A(new_n9802), .B(new_n9801), .Y(new_n9803));
  nand_5 g09427(.A(new_n9569), .B(new_n9556), .Y(new_n9804));
  nand_5 g09428(.A(new_n9570), .B(new_n9549), .Y(new_n9805));
  nand_5 g09429(.A(new_n9805), .B(new_n9804), .Y(new_n9806));
  xor_4  g09430(.A(new_n9806), .B(new_n9552), .Y(new_n9807));
  nand_5 g09431(.A(pi227), .B(pi189), .Y(new_n9808));
  nand_5 g09432(.A(pi217), .B(pi084), .Y(new_n9809));
  xor_4  g09433(.A(new_n9809), .B(new_n9808), .Y(new_n9810));
  xor_4  g09434(.A(new_n9810), .B(new_n9561), .Y(new_n9811));
  nand_5 g09435(.A(pi133), .B(pi081), .Y(new_n9812));
  xor_4  g09436(.A(new_n9812), .B(new_n9562), .Y(new_n9813));
  xor_4  g09437(.A(new_n9813), .B(new_n9811), .Y(new_n9814));
  not_8  g09438(.A(new_n9814), .Y(new_n9815));
  nand_5 g09439(.A(new_n9567), .B(new_n9560), .Y(new_n9816));
  nand_5 g09440(.A(new_n9568), .B(new_n9557), .Y(new_n9817));
  nand_5 g09441(.A(new_n9817), .B(new_n9816), .Y(new_n9818));
  nand_5 g09442(.A(pi187), .B(pi131), .Y(new_n9819));
  nand_5 g09443(.A(pi233), .B(pi052), .Y(new_n9820));
  xor_4  g09444(.A(new_n9820), .B(new_n9819), .Y(new_n9821));
  xor_4  g09445(.A(new_n9821), .B(new_n9550), .Y(new_n9822));
  xor_4  g09446(.A(new_n9822), .B(new_n9818), .Y(new_n9823));
  xor_4  g09447(.A(new_n9823), .B(new_n9815), .Y(new_n9824));
  xor_4  g09448(.A(new_n9824), .B(new_n9807), .Y(new_n9825));
  xor_4  g09449(.A(new_n9825), .B(new_n9803), .Y(new_n9826));
  xor_4  g09450(.A(new_n9826), .B(new_n9800), .Y(new_n9827));
  xor_4  g09451(.A(new_n9827), .B(new_n9798), .Y(new_n9828));
  xor_4  g09452(.A(new_n9828), .B(new_n9690), .Y(po062));
  xor_4  g09453(.A(new_n9314), .B(new_n9313), .Y(po063));
  or_6   g09454(.A(new_n3152), .B(new_n3135), .Y(new_n9831));
  nand_5 g09455(.A(new_n9831), .B(new_n3132), .Y(new_n9832));
  nand_5 g09456(.A(pi095), .B(pi001), .Y(new_n9833));
  nand_5 g09457(.A(new_n3068), .B(new_n2848), .Y(new_n9834));
  nand_5 g09458(.A(new_n3069), .B(new_n3067), .Y(new_n9835));
  nand_5 g09459(.A(new_n9835), .B(new_n9834), .Y(new_n9836));
  xor_4  g09460(.A(new_n9836), .B(new_n9833), .Y(new_n9837));
  xor_4  g09461(.A(new_n9837), .B(new_n9832), .Y(new_n9838));
  nor_5  g09462(.A(new_n3080), .B(new_n3056), .Y(new_n9839));
  not_8  g09463(.A(new_n3081), .Y(new_n9840));
  nor_5  g09464(.A(new_n9840), .B(new_n3055), .Y(new_n9841));
  nor_5  g09465(.A(new_n9841), .B(new_n9839), .Y(new_n9842));
  nand_5 g09466(.A(pi185), .B(pi060), .Y(new_n9843));
  not_8  g09467(.A(new_n3149), .Y(new_n9844));
  nor_5  g09468(.A(new_n9844), .B(new_n3146), .Y(new_n9845));
  nor_5  g09469(.A(new_n3150), .B(new_n3142), .Y(new_n9846));
  nor_5  g09470(.A(new_n9846), .B(new_n9845), .Y(new_n9847));
  nand_5 g09471(.A(pi138), .B(pi078), .Y(new_n9848));
  xor_4  g09472(.A(new_n9848), .B(new_n9847), .Y(new_n9849));
  xor_4  g09473(.A(new_n9849), .B(new_n9843), .Y(new_n9850));
  xor_4  g09474(.A(new_n9850), .B(new_n9842), .Y(new_n9851));
  not_8  g09475(.A(new_n3128), .Y(new_n9852));
  nor_5  g09476(.A(new_n3153), .B(new_n9852), .Y(new_n9853));
  nor_5  g09477(.A(new_n3154), .B(new_n3127), .Y(new_n9854));
  nor_5  g09478(.A(new_n9854), .B(new_n9853), .Y(new_n9855));
  nand_5 g09479(.A(pi135), .B(pi089), .Y(new_n9856));
  xor_4  g09480(.A(new_n9856), .B(new_n9855), .Y(new_n9857));
  xor_4  g09481(.A(new_n9857), .B(new_n9851), .Y(new_n9858));
  xor_4  g09482(.A(new_n9858), .B(new_n9838), .Y(new_n9859));
  or_6   g09483(.A(new_n3114), .B(new_n3097), .Y(new_n9860));
  nand_5 g09484(.A(new_n9860), .B(new_n3095), .Y(new_n9861));
  nand_5 g09485(.A(pi030), .B(pi020), .Y(new_n9862));
  nand_5 g09486(.A(pi251), .B(pi062), .Y(new_n9863));
  nand_5 g09487(.A(pi120), .B(pi079), .Y(new_n9864));
  xor_4  g09488(.A(new_n9864), .B(new_n9863), .Y(new_n9865));
  xor_4  g09489(.A(new_n9865), .B(new_n9862), .Y(new_n9866));
  xor_4  g09490(.A(new_n9866), .B(new_n9861), .Y(new_n9867));
  nand_5 g09491(.A(pi197), .B(pi182), .Y(new_n9868));
  nor_5  g09492(.A(new_n3155), .B(new_n3123), .Y(new_n9869));
  nor_5  g09493(.A(new_n3156), .B(new_n3019), .Y(new_n9870));
  nor_5  g09494(.A(new_n9870), .B(new_n9869), .Y(new_n9871));
  xor_4  g09495(.A(new_n9871), .B(new_n9868), .Y(new_n9872));
  xor_4  g09496(.A(new_n9872), .B(new_n9867), .Y(new_n9873));
  xor_4  g09497(.A(new_n9873), .B(new_n9859), .Y(new_n9874));
  nand_5 g09498(.A(pi220), .B(pi160), .Y(new_n9875));
  nand_5 g09499(.A(new_n3144), .B(new_n3143), .Y(new_n9876));
  nand_5 g09500(.A(new_n3145), .B(new_n2973), .Y(new_n9877));
  nand_5 g09501(.A(new_n9877), .B(new_n9876), .Y(new_n9878));
  xor_4  g09502(.A(new_n9878), .B(new_n9875), .Y(new_n9879));
  nand_5 g09503(.A(pi216), .B(pi198), .Y(new_n9880));
  or_6   g09504(.A(new_n3082), .B(new_n3052), .Y(new_n9881));
  nand_5 g09505(.A(new_n3087), .B(new_n3083), .Y(new_n9882));
  nand_5 g09506(.A(new_n9882), .B(new_n9881), .Y(new_n9883));
  xor_4  g09507(.A(new_n9883), .B(new_n9880), .Y(new_n9884));
  xor_4  g09508(.A(new_n9884), .B(new_n9879), .Y(new_n9885));
  nand_5 g09509(.A(pi177), .B(pi092), .Y(new_n9886));
  nand_5 g09510(.A(new_n3139), .B(new_n3138), .Y(new_n9887));
  nand_5 g09511(.A(new_n3140), .B(new_n2962), .Y(new_n9888));
  nand_5 g09512(.A(new_n9888), .B(new_n9887), .Y(new_n9889));
  xor_4  g09513(.A(new_n9889), .B(new_n9886), .Y(new_n9890));
  nand_5 g09514(.A(pi219), .B(pi209), .Y(new_n9891));
  nand_5 g09515(.A(pi190), .B(pi137), .Y(new_n9892));
  nand_5 g09516(.A(pi170), .B(pi086), .Y(new_n9893));
  xor_4  g09517(.A(new_n9893), .B(new_n9892), .Y(new_n9894));
  nand_5 g09518(.A(pi172), .B(pi076), .Y(new_n9895));
  xor_4  g09519(.A(new_n9895), .B(new_n9894), .Y(new_n9896));
  xor_4  g09520(.A(new_n9896), .B(new_n9891), .Y(new_n9897));
  xor_4  g09521(.A(new_n9897), .B(new_n9890), .Y(new_n9898));
  nor_5  g09522(.A(new_n3115), .B(new_n3089), .Y(new_n9899));
  not_8  g09523(.A(new_n3116), .Y(new_n9900));
  nor_5  g09524(.A(new_n3120), .B(new_n9900), .Y(new_n9901));
  nor_5  g09525(.A(new_n9901), .B(new_n9899), .Y(new_n9902));
  nor_5  g09526(.A(new_n3136), .B(new_n2964), .Y(new_n9903));
  nor_5  g09527(.A(new_n3141), .B(new_n3137), .Y(new_n9904));
  nor_5  g09528(.A(new_n9904), .B(new_n9903), .Y(new_n9905));
  nand_5 g09529(.A(pi192), .B(pi065), .Y(new_n9906));
  nand_5 g09530(.A(pi229), .B(pi225), .Y(new_n9907));
  xor_4  g09531(.A(new_n9907), .B(new_n9906), .Y(new_n9908));
  xor_4  g09532(.A(new_n9908), .B(new_n9905), .Y(new_n9909));
  nand_5 g09533(.A(pi101), .B(pi067), .Y(new_n9910));
  nand_5 g09534(.A(pi223), .B(pi053), .Y(new_n9911));
  xor_4  g09535(.A(new_n9911), .B(new_n9910), .Y(new_n9912));
  nor_5  g09536(.A(new_n3102), .B(new_n2892), .Y(new_n9913));
  nor_5  g09537(.A(new_n3103), .B(new_n3101), .Y(new_n9914));
  nor_5  g09538(.A(new_n9914), .B(new_n9913), .Y(new_n9915));
  nand_5 g09539(.A(pi102), .B(pi006), .Y(new_n9916));
  xor_4  g09540(.A(new_n9916), .B(new_n9915), .Y(new_n9917));
  xor_4  g09541(.A(new_n9917), .B(new_n9912), .Y(new_n9918));
  xor_4  g09542(.A(new_n9918), .B(new_n9909), .Y(new_n9919));
  xor_4  g09543(.A(new_n9919), .B(new_n9902), .Y(new_n9920));
  xor_4  g09544(.A(new_n9920), .B(new_n9898), .Y(new_n9921));
  xor_4  g09545(.A(new_n9921), .B(new_n9885), .Y(new_n9922));
  or_6   g09546(.A(new_n3036), .B(new_n3032), .Y(new_n9923));
  nand_5 g09547(.A(new_n3044), .B(new_n3037), .Y(new_n9924));
  nand_5 g09548(.A(new_n9924), .B(new_n9923), .Y(new_n9925));
  nand_5 g09549(.A(new_n3060), .B(new_n3059), .Y(new_n9926));
  nand_5 g09550(.A(new_n3061), .B(new_n2854), .Y(new_n9927));
  nand_5 g09551(.A(new_n9927), .B(new_n9926), .Y(new_n9928));
  xor_4  g09552(.A(new_n9928), .B(new_n9925), .Y(new_n9929));
  nand_5 g09553(.A(pi153), .B(pi087), .Y(new_n9930));
  nand_5 g09554(.A(new_n3034), .B(new_n3033), .Y(new_n9931));
  nand_5 g09555(.A(new_n3035), .B(new_n2811), .Y(new_n9932));
  nand_5 g09556(.A(new_n9932), .B(new_n9931), .Y(new_n9933));
  xor_4  g09557(.A(new_n9933), .B(new_n9930), .Y(new_n9934));
  nand_5 g09558(.A(new_n3041), .B(new_n3040), .Y(new_n9935));
  nand_5 g09559(.A(new_n3042), .B(new_n2822), .Y(new_n9936));
  nand_5 g09560(.A(new_n9936), .B(new_n9935), .Y(new_n9937));
  nand_5 g09561(.A(pi215), .B(pi071), .Y(new_n9938));
  nand_5 g09562(.A(pi169), .B(pi124), .Y(new_n9939));
  xor_4  g09563(.A(new_n9939), .B(new_n9938), .Y(new_n9940));
  xor_4  g09564(.A(new_n9940), .B(new_n9937), .Y(new_n9941));
  xor_4  g09565(.A(new_n9941), .B(new_n9934), .Y(new_n9942));
  xor_4  g09566(.A(new_n9942), .B(new_n9929), .Y(new_n9943));
  nor_5  g09567(.A(new_n3038), .B(new_n2824), .Y(new_n9944));
  nor_5  g09568(.A(new_n3043), .B(new_n3039), .Y(new_n9945));
  nor_5  g09569(.A(new_n9945), .B(new_n9944), .Y(new_n9946));
  or_6   g09570(.A(new_n3079), .B(new_n3072), .Y(new_n9947));
  nand_5 g09571(.A(new_n9947), .B(new_n3078), .Y(new_n9948));
  xor_4  g09572(.A(new_n9948), .B(new_n9946), .Y(new_n9949));
  nand_5 g09573(.A(pi142), .B(pi022), .Y(new_n9950));
  nand_5 g09574(.A(pi130), .B(pi123), .Y(new_n9951));
  xor_4  g09575(.A(new_n9951), .B(new_n9950), .Y(new_n9952));
  xor_4  g09576(.A(new_n9952), .B(new_n9949), .Y(new_n9953));
  xor_4  g09577(.A(new_n9953), .B(new_n9943), .Y(new_n9954));
  xor_4  g09578(.A(new_n9954), .B(new_n9922), .Y(new_n9955));
  xor_4  g09579(.A(new_n9955), .B(new_n9874), .Y(new_n9956));
  nand_5 g09580(.A(pi155), .B(pi004), .Y(new_n9957));
  nand_5 g09581(.A(pi154), .B(pi122), .Y(new_n9958));
  not_8  g09582(.A(new_n3048), .Y(new_n9959));
  nor_5  g09583(.A(new_n9959), .B(new_n2812), .Y(new_n9960));
  nor_5  g09584(.A(new_n3049), .B(new_n3045), .Y(new_n9961));
  nor_5  g09585(.A(new_n9961), .B(new_n9960), .Y(new_n9962));
  xor_4  g09586(.A(new_n9962), .B(new_n9958), .Y(new_n9963));
  xor_4  g09587(.A(new_n9963), .B(new_n9957), .Y(new_n9964));
  nand_5 g09588(.A(pi165), .B(pi041), .Y(new_n9965));
  xor_4  g09589(.A(new_n9965), .B(new_n9964), .Y(new_n9966));
  nand_5 g09590(.A(new_n3121), .B(new_n3088), .Y(new_n9967));
  not_8  g09591(.A(new_n3022), .Y(new_n9968));
  or_6   g09592(.A(new_n3122), .B(new_n9968), .Y(new_n9969));
  nand_5 g09593(.A(new_n9969), .B(new_n9967), .Y(new_n9970));
  nor_5  g09594(.A(new_n3111), .B(new_n3107), .Y(new_n9971));
  not_8  g09595(.A(new_n3104), .Y(new_n9972));
  nor_5  g09596(.A(new_n3112), .B(new_n9972), .Y(new_n9973));
  nor_5  g09597(.A(new_n9973), .B(new_n9971), .Y(new_n9974));
  xor_4  g09598(.A(new_n9974), .B(new_n9970), .Y(new_n9975));
  or_6   g09599(.A(new_n3070), .B(new_n3066), .Y(new_n9976));
  nand_5 g09600(.A(new_n3071), .B(new_n3063), .Y(new_n9977));
  nand_5 g09601(.A(new_n9977), .B(new_n9976), .Y(new_n9978));
  nand_5 g09602(.A(new_n3109), .B(new_n3108), .Y(new_n9979));
  nand_5 g09603(.A(new_n3110), .B(new_n2880), .Y(new_n9980));
  nand_5 g09604(.A(new_n9980), .B(new_n9979), .Y(new_n9981));
  nand_5 g09605(.A(pi073), .B(pi023), .Y(new_n9982));
  xor_4  g09606(.A(new_n9982), .B(new_n9981), .Y(new_n9983));
  xor_4  g09607(.A(new_n9983), .B(new_n9978), .Y(new_n9984));
  nor_5  g09608(.A(new_n3057), .B(new_n2856), .Y(new_n9985));
  nor_5  g09609(.A(new_n3062), .B(new_n3058), .Y(new_n9986));
  nor_5  g09610(.A(new_n9986), .B(new_n9985), .Y(new_n9987));
  nand_5 g09611(.A(pi254), .B(pi094), .Y(new_n9988));
  nand_5 g09612(.A(pi158), .B(pi059), .Y(new_n9989));
  xor_4  g09613(.A(new_n9989), .B(new_n9988), .Y(new_n9990));
  xor_4  g09614(.A(new_n9990), .B(new_n9987), .Y(new_n9991));
  xor_4  g09615(.A(new_n9991), .B(new_n9984), .Y(new_n9992));
  xor_4  g09616(.A(new_n9992), .B(new_n9975), .Y(new_n9993));
  nand_5 g09617(.A(new_n3099), .B(new_n3098), .Y(new_n9994));
  nand_5 g09618(.A(new_n3100), .B(new_n2890), .Y(new_n9995));
  nand_5 g09619(.A(new_n9995), .B(new_n9994), .Y(new_n9996));
  nand_5 g09620(.A(pi099), .B(pi003), .Y(new_n9997));
  xor_4  g09621(.A(new_n9997), .B(new_n9996), .Y(new_n9998));
  nor_5  g09622(.A(new_n3050), .B(new_n3029), .Y(new_n9999));
  not_8  g09623(.A(new_n3051), .Y(new_n10000));
  nor_5  g09624(.A(new_n10000), .B(new_n3027), .Y(new_n10001));
  or_6   g09625(.A(new_n10001), .B(new_n9999), .Y(new_n10002));
  xor_4  g09626(.A(new_n10002), .B(new_n9998), .Y(new_n10003));
  xor_4  g09627(.A(new_n10003), .B(new_n9993), .Y(new_n10004));
  xor_4  g09628(.A(new_n10004), .B(new_n9966), .Y(new_n10005));
  xor_4  g09629(.A(new_n10005), .B(new_n9956), .Y(po064));
  xnor_4 g09630(.A(new_n9327), .B(new_n9326), .Y(po065));
  xnor_4 g09631(.A(new_n3003), .B(new_n3002), .Y(po066));
  xor_4  g09632(.A(new_n5038), .B(new_n5033), .Y(po067));
  xor_4  g09633(.A(new_n7068), .B(new_n7066), .Y(po068));
  xnor_4 g09634(.A(new_n4241), .B(new_n4240), .Y(po069));
  xnor_4 g09635(.A(new_n1146), .B(new_n1111), .Y(po070));
  xnor_4 g09636(.A(new_n9332), .B(new_n9331), .Y(po071));
  nand_5 g09637(.A(new_n6587), .B(new_n6586), .Y(new_n10014));
  nand_5 g09638(.A(new_n6616), .B(new_n6588), .Y(new_n10015));
  nand_5 g09639(.A(new_n10015), .B(new_n10014), .Y(new_n10016));
  not_8  g09640(.A(new_n6612), .Y(new_n10017));
  nor_5  g09641(.A(new_n6615), .B(new_n10017), .Y(new_n10018));
  not_8  g09642(.A(new_n6604), .Y(new_n10019));
  nor_5  g09643(.A(new_n6610), .B(new_n10019), .Y(new_n10020));
  nor_5  g09644(.A(new_n6611), .B(new_n6591), .Y(new_n10021));
  xor_4  g09645(.A(new_n10021), .B(new_n6609), .Y(new_n10022));
  nor_5  g09646(.A(new_n10022), .B(new_n10020), .Y(new_n10023));
  nor_5  g09647(.A(new_n6595), .B(new_n6592), .Y(new_n10024));
  nor_5  g09648(.A(new_n6603), .B(new_n6596), .Y(new_n10025));
  nor_5  g09649(.A(new_n10025), .B(new_n10024), .Y(new_n10026));
  nand_5 g09650(.A(pi241), .B(pi113), .Y(new_n10027));
  nand_5 g09651(.A(pi236), .B(pi038), .Y(new_n10028));
  xor_4  g09652(.A(new_n10028), .B(new_n10027), .Y(new_n10029));
  xor_4  g09653(.A(new_n10029), .B(new_n6608), .Y(new_n10030));
  xor_4  g09654(.A(new_n10030), .B(new_n10026), .Y(new_n10031));
  nand_5 g09655(.A(pi051), .B(pi018), .Y(new_n10032));
  nand_5 g09656(.A(pi108), .B(pi090), .Y(new_n10033));
  xor_4  g09657(.A(new_n10033), .B(new_n10032), .Y(new_n10034));
  xor_4  g09658(.A(new_n10034), .B(new_n6600), .Y(new_n10035));
  nand_5 g09659(.A(pi141), .B(pi007), .Y(new_n10036));
  xor_4  g09660(.A(new_n10036), .B(new_n6601), .Y(new_n10037));
  xor_4  g09661(.A(new_n10037), .B(new_n10035), .Y(new_n10038));
  not_8  g09662(.A(new_n10038), .Y(new_n10039));
  xor_4  g09663(.A(new_n10039), .B(new_n10031), .Y(new_n10040));
  xor_4  g09664(.A(new_n10040), .B(new_n10023), .Y(new_n10041));
  xor_4  g09665(.A(new_n10041), .B(new_n10018), .Y(new_n10042));
  xor_4  g09666(.A(new_n10042), .B(new_n10016), .Y(new_n10043));
  nand_5 g09667(.A(new_n6583), .B(new_n6582), .Y(new_n10044));
  nand_5 g09668(.A(new_n6584), .B(new_n6553), .Y(new_n10045));
  nand_5 g09669(.A(new_n10045), .B(new_n10044), .Y(new_n10046));
  nor_5  g09670(.A(new_n6581), .B(new_n6557), .Y(new_n10047));
  nand_5 g09671(.A(new_n6577), .B(new_n6570), .Y(new_n10048));
  nand_5 g09672(.A(new_n6578), .B(new_n6569), .Y(new_n10049));
  nand_5 g09673(.A(new_n10049), .B(new_n10048), .Y(new_n10050));
  nand_5 g09674(.A(pi212), .B(pi098), .Y(new_n10051));
  nand_5 g09675(.A(pi213), .B(pi043), .Y(new_n10052));
  xor_4  g09676(.A(new_n10052), .B(new_n10051), .Y(new_n10053));
  xor_4  g09677(.A(new_n10053), .B(new_n6564), .Y(new_n10054));
  xor_4  g09678(.A(new_n10054), .B(new_n10050), .Y(new_n10055));
  not_8  g09679(.A(new_n10055), .Y(new_n10056));
  nand_5 g09680(.A(pi013), .B(pi012), .Y(new_n10057));
  xor_4  g09681(.A(new_n10057), .B(new_n6575), .Y(new_n10058));
  nand_5 g09682(.A(pi188), .B(pi183), .Y(new_n10059));
  nand_5 g09683(.A(pi112), .B(pi061), .Y(new_n10060));
  xor_4  g09684(.A(new_n10060), .B(new_n10059), .Y(new_n10061));
  xor_4  g09685(.A(new_n10061), .B(new_n6574), .Y(new_n10062));
  xor_4  g09686(.A(new_n10062), .B(new_n10058), .Y(new_n10063));
  xor_4  g09687(.A(new_n10063), .B(new_n10056), .Y(new_n10064));
  nor_5  g09688(.A(new_n6579), .B(new_n6566), .Y(new_n10065));
  not_8  g09689(.A(new_n6580), .Y(new_n10066));
  nor_5  g09690(.A(new_n10066), .B(new_n6560), .Y(new_n10067));
  xor_4  g09691(.A(new_n10067), .B(new_n6565), .Y(new_n10068));
  nor_5  g09692(.A(new_n10068), .B(new_n10065), .Y(new_n10069));
  xor_4  g09693(.A(new_n10069), .B(new_n10064), .Y(new_n10070));
  nand_5 g09694(.A(new_n10070), .B(new_n10047), .Y(new_n10071));
  or_6   g09695(.A(new_n10070), .B(new_n10047), .Y(new_n10072));
  and_6  g09696(.A(new_n10072), .B(new_n10071), .Y(new_n10073));
  xor_4  g09697(.A(new_n10073), .B(new_n10046), .Y(new_n10074));
  xor_4  g09698(.A(new_n10074), .B(new_n10043), .Y(new_n10075));
  or_6   g09699(.A(new_n6617), .B(new_n6585), .Y(new_n10076));
  nand_5 g09700(.A(new_n6622), .B(new_n6618), .Y(new_n10077));
  and_6  g09701(.A(new_n10077), .B(new_n10076), .Y(new_n10078));
  xnor_4 g09702(.A(new_n10078), .B(new_n10075), .Y(new_n10079));
  nand_5 g09703(.A(new_n6519), .B(new_n6518), .Y(new_n10080));
  nand_5 g09704(.A(new_n6550), .B(new_n6520), .Y(new_n10081));
  nand_5 g09705(.A(new_n10081), .B(new_n10080), .Y(new_n10082));
  not_8  g09706(.A(new_n6545), .Y(new_n10083));
  nor_5  g09707(.A(new_n6549), .B(new_n10083), .Y(new_n10084));
  nand_5 g09708(.A(pi048), .B(pi035), .Y(new_n10085));
  xor_4  g09709(.A(new_n10085), .B(new_n6538), .Y(new_n10086));
  nand_5 g09710(.A(pi179), .B(pi015), .Y(new_n10087));
  nand_5 g09711(.A(pi162), .B(pi146), .Y(new_n10088));
  xor_4  g09712(.A(new_n10088), .B(new_n10087), .Y(new_n10089));
  xor_4  g09713(.A(new_n10089), .B(new_n6537), .Y(new_n10090));
  xor_4  g09714(.A(new_n10090), .B(new_n10086), .Y(new_n10091));
  nand_5 g09715(.A(new_n6540), .B(new_n6533), .Y(new_n10092));
  nand_5 g09716(.A(new_n6541), .B(new_n6532), .Y(new_n10093));
  nand_5 g09717(.A(new_n10093), .B(new_n10092), .Y(new_n10094));
  nand_5 g09718(.A(pi193), .B(pi168), .Y(new_n10095));
  nand_5 g09719(.A(pi238), .B(pi208), .Y(new_n10096));
  xor_4  g09720(.A(new_n10096), .B(new_n10095), .Y(new_n10097));
  xor_4  g09721(.A(new_n10097), .B(new_n6527), .Y(new_n10098));
  xor_4  g09722(.A(new_n10098), .B(new_n10094), .Y(new_n10099));
  xor_4  g09723(.A(new_n10099), .B(new_n10091), .Y(new_n10100));
  nor_5  g09724(.A(new_n6544), .B(new_n6523), .Y(new_n10101));
  and_6  g09725(.A(new_n10101), .B(new_n6528), .Y(new_n10102));
  nor_5  g09726(.A(new_n6542), .B(new_n6529), .Y(new_n10103));
  nor_5  g09727(.A(new_n10103), .B(new_n6528), .Y(new_n10104));
  not_8  g09728(.A(new_n10104), .Y(new_n10105));
  nor_5  g09729(.A(new_n10105), .B(new_n10101), .Y(new_n10106));
  or_6   g09730(.A(new_n10106), .B(new_n10102), .Y(new_n10107));
  xor_4  g09731(.A(new_n10107), .B(new_n10100), .Y(new_n10108));
  xor_4  g09732(.A(new_n10108), .B(new_n10084), .Y(new_n10109));
  xnor_4 g09733(.A(new_n10109), .B(new_n10082), .Y(new_n10110));
  xor_4  g09734(.A(new_n10110), .B(new_n10079), .Y(new_n10111));
  nor_5  g09735(.A(new_n6551), .B(new_n6517), .Y(new_n10112));
  nor_5  g09736(.A(new_n6623), .B(new_n6552), .Y(new_n10113));
  nor_5  g09737(.A(new_n10113), .B(new_n10112), .Y(new_n10114));
  xor_4  g09738(.A(new_n10114), .B(new_n10111), .Y(new_n10115));
  nand_5 g09739(.A(new_n6479), .B(new_n6478), .Y(new_n10116));
  not_8  g09740(.A(new_n10116), .Y(new_n10117));
  nor_5  g09741(.A(new_n6509), .B(new_n6481), .Y(new_n10118));
  nor_5  g09742(.A(new_n10118), .B(new_n10117), .Y(new_n10119));
  nor_5  g09743(.A(new_n6508), .B(new_n6484), .Y(new_n10120));
  not_8  g09744(.A(new_n6507), .Y(new_n10121));
  nor_5  g09745(.A(new_n10121), .B(new_n6487), .Y(new_n10122));
  and_6  g09746(.A(new_n10122), .B(new_n6492), .Y(new_n10123));
  nor_5  g09747(.A(new_n6506), .B(new_n6493), .Y(new_n10124));
  nor_5  g09748(.A(new_n10124), .B(new_n6492), .Y(new_n10125));
  not_8  g09749(.A(new_n10125), .Y(new_n10126));
  nor_5  g09750(.A(new_n10126), .B(new_n10122), .Y(new_n10127));
  or_6   g09751(.A(new_n10127), .B(new_n10123), .Y(new_n10128));
  nand_5 g09752(.A(new_n6504), .B(new_n6497), .Y(new_n10129));
  nand_5 g09753(.A(new_n6505), .B(new_n6496), .Y(new_n10130));
  nand_5 g09754(.A(new_n10130), .B(new_n10129), .Y(new_n10131));
  nand_5 g09755(.A(pi131), .B(pi068), .Y(new_n10132));
  nand_5 g09756(.A(pi052), .B(pi036), .Y(new_n10133));
  xor_4  g09757(.A(new_n10133), .B(new_n10132), .Y(new_n10134));
  xor_4  g09758(.A(new_n10134), .B(new_n6491), .Y(new_n10135));
  xnor_4 g09759(.A(new_n10135), .B(new_n10131), .Y(new_n10136));
  nand_5 g09760(.A(pi133), .B(pi085), .Y(new_n10137));
  xor_4  g09761(.A(new_n10137), .B(new_n6503), .Y(new_n10138));
  nand_5 g09762(.A(pi194), .B(pi189), .Y(new_n10139));
  nand_5 g09763(.A(pi143), .B(pi084), .Y(new_n10140));
  xor_4  g09764(.A(new_n10140), .B(new_n10139), .Y(new_n10141));
  xnor_4 g09765(.A(new_n10141), .B(new_n6501), .Y(new_n10142));
  xnor_4 g09766(.A(new_n10142), .B(new_n10138), .Y(new_n10143));
  xor_4  g09767(.A(new_n10143), .B(new_n10136), .Y(new_n10144));
  xor_4  g09768(.A(new_n10144), .B(new_n10128), .Y(new_n10145));
  xor_4  g09769(.A(new_n10145), .B(new_n10120), .Y(new_n10146));
  xor_4  g09770(.A(new_n10146), .B(new_n10119), .Y(new_n10147));
  or_6   g09771(.A(new_n10147), .B(new_n10115), .Y(new_n10148));
  not_8  g09772(.A(new_n6510), .Y(new_n10149));
  nor_5  g09773(.A(new_n6513), .B(new_n10149), .Y(new_n10150));
  nor_5  g09774(.A(new_n6624), .B(new_n6514), .Y(new_n10151));
  nor_5  g09775(.A(new_n10151), .B(new_n10150), .Y(new_n10152));
  xor_4  g09776(.A(new_n10147), .B(new_n10115), .Y(new_n10153));
  nand_5 g09777(.A(new_n10153), .B(new_n10152), .Y(new_n10154));
  nand_5 g09778(.A(new_n10154), .B(new_n10148), .Y(new_n10155));
  nand_5 g09779(.A(pi112), .B(pi012), .Y(new_n10156));
  xor_4  g09780(.A(new_n10156), .B(new_n10155), .Y(new_n10157));
  nand_5 g09781(.A(new_n10033), .B(new_n10032), .Y(new_n10158));
  nand_5 g09782(.A(new_n10034), .B(new_n6600), .Y(new_n10159));
  nand_5 g09783(.A(new_n10159), .B(new_n10158), .Y(new_n10160));
  nand_5 g09784(.A(pi084), .B(pi057), .Y(new_n10161));
  xor_4  g09785(.A(new_n10161), .B(new_n10160), .Y(new_n10162));
  nand_5 g09786(.A(new_n10071), .B(new_n10046), .Y(new_n10163));
  nand_5 g09787(.A(new_n10163), .B(new_n10072), .Y(new_n10164));
  nand_5 g09788(.A(pi204), .B(pi179), .Y(new_n10165));
  nor_5  g09789(.A(new_n10098), .B(new_n10094), .Y(new_n10166));
  and_6  g09790(.A(new_n10099), .B(new_n10091), .Y(new_n10167));
  nor_5  g09791(.A(new_n10167), .B(new_n10166), .Y(new_n10168));
  xor_4  g09792(.A(new_n10168), .B(new_n10165), .Y(new_n10169));
  xor_4  g09793(.A(new_n10169), .B(new_n10164), .Y(new_n10170));
  nand_5 g09794(.A(pi183), .B(pi178), .Y(new_n10171));
  nand_5 g09795(.A(new_n10096), .B(new_n10095), .Y(new_n10172));
  nand_5 g09796(.A(new_n10097), .B(new_n6527), .Y(new_n10173));
  nand_5 g09797(.A(new_n10173), .B(new_n10172), .Y(new_n10174));
  nand_5 g09798(.A(pi237), .B(pi035), .Y(new_n10175));
  xnor_4 g09799(.A(new_n10175), .B(new_n10174), .Y(new_n10176));
  xor_4  g09800(.A(new_n10176), .B(new_n10171), .Y(new_n10177));
  xor_4  g09801(.A(new_n10177), .B(new_n10170), .Y(new_n10178));
  nand_5 g09802(.A(pi161), .B(pi113), .Y(new_n10179));
  nand_5 g09803(.A(pi194), .B(pi064), .Y(new_n10180));
  nand_5 g09804(.A(pi068), .B(pi052), .Y(new_n10181));
  nand_5 g09805(.A(pi162), .B(pi152), .Y(new_n10182));
  xor_4  g09806(.A(new_n10182), .B(new_n10181), .Y(new_n10183));
  xor_4  g09807(.A(new_n10183), .B(new_n10180), .Y(new_n10184));
  xor_4  g09808(.A(new_n10184), .B(new_n10179), .Y(new_n10185));
  nand_5 g09809(.A(new_n10110), .B(new_n10079), .Y(new_n10186));
  nand_5 g09810(.A(new_n10114), .B(new_n10111), .Y(new_n10187));
  nand_5 g09811(.A(new_n10187), .B(new_n10186), .Y(new_n10188));
  nand_5 g09812(.A(pi180), .B(pi133), .Y(new_n10189));
  nor_5  g09813(.A(new_n10135), .B(new_n10131), .Y(new_n10190));
  nor_5  g09814(.A(new_n10143), .B(new_n10136), .Y(new_n10191));
  nor_5  g09815(.A(new_n10191), .B(new_n10190), .Y(new_n10192));
  xor_4  g09816(.A(new_n10192), .B(new_n10189), .Y(new_n10193));
  nor_5  g09817(.A(new_n10036), .B(new_n6602), .Y(new_n10194));
  nor_5  g09818(.A(new_n10037), .B(new_n10035), .Y(new_n10195));
  or_6   g09819(.A(new_n10195), .B(new_n10194), .Y(new_n10196));
  nand_5 g09820(.A(pi108), .B(pi047), .Y(new_n10197));
  nand_5 g09821(.A(pi212), .B(pi043), .Y(new_n10198));
  nand_5 g09822(.A(pi104), .B(pi098), .Y(new_n10199));
  xor_4  g09823(.A(new_n10199), .B(new_n10198), .Y(new_n10200));
  xor_4  g09824(.A(new_n10200), .B(new_n10197), .Y(new_n10201));
  xor_4  g09825(.A(new_n10201), .B(new_n10196), .Y(new_n10202));
  nand_5 g09826(.A(pi189), .B(pi085), .Y(new_n10203));
  nor_5  g09827(.A(new_n10107), .B(new_n10100), .Y(new_n10204));
  nor_5  g09828(.A(new_n10204), .B(new_n10106), .Y(new_n10205));
  nand_5 g09829(.A(pi168), .B(pi159), .Y(new_n10206));
  xor_4  g09830(.A(new_n10206), .B(new_n10205), .Y(new_n10207));
  xor_4  g09831(.A(new_n10207), .B(new_n10203), .Y(new_n10208));
  xor_4  g09832(.A(new_n10208), .B(new_n10202), .Y(new_n10209));
  xor_4  g09833(.A(new_n10209), .B(new_n10193), .Y(new_n10210));
  nand_5 g09834(.A(pi141), .B(pi118), .Y(new_n10211));
  nand_5 g09835(.A(new_n10052), .B(new_n10051), .Y(new_n10212));
  nand_5 g09836(.A(new_n10053), .B(new_n6564), .Y(new_n10213));
  nand_5 g09837(.A(new_n10213), .B(new_n10212), .Y(new_n10214));
  xor_4  g09838(.A(new_n10214), .B(new_n10211), .Y(new_n10215));
  or_6   g09839(.A(new_n10041), .B(new_n10018), .Y(new_n10216));
  nand_5 g09840(.A(new_n10042), .B(new_n10016), .Y(new_n10217));
  nand_5 g09841(.A(new_n10217), .B(new_n10216), .Y(new_n10218));
  and_6  g09842(.A(new_n10021), .B(new_n6609), .Y(new_n10219));
  nor_5  g09843(.A(new_n10040), .B(new_n10023), .Y(new_n10220));
  nor_5  g09844(.A(new_n10220), .B(new_n10219), .Y(new_n10221));
  xor_4  g09845(.A(new_n10221), .B(new_n10218), .Y(new_n10222));
  xor_4  g09846(.A(new_n10222), .B(new_n10215), .Y(new_n10223));
  and_6  g09847(.A(new_n10054), .B(new_n10050), .Y(new_n10224));
  nor_5  g09848(.A(new_n10063), .B(new_n10056), .Y(new_n10225));
  nor_5  g09849(.A(new_n10225), .B(new_n10224), .Y(new_n10226));
  nand_5 g09850(.A(pi144), .B(pi013), .Y(new_n10227));
  xor_4  g09851(.A(new_n10227), .B(new_n10226), .Y(new_n10228));
  nand_5 g09852(.A(pi077), .B(pi036), .Y(new_n10229));
  xor_4  g09853(.A(new_n10229), .B(new_n10228), .Y(new_n10230));
  xor_4  g09854(.A(new_n10230), .B(new_n10223), .Y(new_n10231));
  xor_4  g09855(.A(new_n10231), .B(new_n10210), .Y(new_n10232));
  xor_4  g09856(.A(new_n10232), .B(new_n10188), .Y(new_n10233));
  xor_4  g09857(.A(new_n10233), .B(new_n10185), .Y(new_n10234));
  xor_4  g09858(.A(new_n10234), .B(new_n10178), .Y(new_n10235));
  xor_4  g09859(.A(new_n10235), .B(new_n10162), .Y(new_n10236));
  xor_4  g09860(.A(new_n10236), .B(new_n10157), .Y(new_n10237));
  or_6   g09861(.A(new_n10137), .B(new_n6503), .Y(new_n10238));
  nand_5 g09862(.A(new_n10142), .B(new_n10138), .Y(new_n10239));
  nand_5 g09863(.A(new_n10239), .B(new_n10238), .Y(new_n10240));
  nand_5 g09864(.A(pi188), .B(pi088), .Y(new_n10241));
  xor_4  g09865(.A(new_n10241), .B(new_n10240), .Y(new_n10242));
  nor_5  g09866(.A(new_n10144), .B(new_n10128), .Y(new_n10243));
  nor_5  g09867(.A(new_n10243), .B(new_n10127), .Y(new_n10244));
  xor_4  g09868(.A(new_n10244), .B(new_n10242), .Y(new_n10245));
  nand_5 g09869(.A(pi090), .B(pi007), .Y(new_n10246));
  nand_5 g09870(.A(pi146), .B(pi033), .Y(new_n10247));
  nand_5 g09871(.A(pi236), .B(pi028), .Y(new_n10248));
  xor_4  g09872(.A(new_n10248), .B(new_n10247), .Y(new_n10249));
  xor_4  g09873(.A(new_n10249), .B(new_n10246), .Y(new_n10250));
  xor_4  g09874(.A(new_n10250), .B(new_n10245), .Y(new_n10251));
  nand_5 g09875(.A(new_n10030), .B(new_n10026), .Y(new_n10252));
  nand_5 g09876(.A(new_n10039), .B(new_n10031), .Y(new_n10253));
  nand_5 g09877(.A(new_n10253), .B(new_n10252), .Y(new_n10254));
  nand_5 g09878(.A(pi131), .B(pi046), .Y(new_n10255));
  xnor_4 g09879(.A(new_n10255), .B(new_n10254), .Y(new_n10256));
  or_6   g09880(.A(new_n10074), .B(new_n10043), .Y(new_n10257));
  nand_5 g09881(.A(new_n10078), .B(new_n10075), .Y(new_n10258));
  nand_5 g09882(.A(new_n10258), .B(new_n10257), .Y(new_n10259));
  nand_5 g09883(.A(new_n10067), .B(new_n6565), .Y(new_n10260));
  or_6   g09884(.A(new_n10069), .B(new_n10064), .Y(new_n10261));
  nand_5 g09885(.A(new_n10261), .B(new_n10260), .Y(new_n10262));
  xor_4  g09886(.A(new_n10262), .B(new_n10259), .Y(new_n10263));
  nand_5 g09887(.A(pi128), .B(pi051), .Y(new_n10264));
  not_8  g09888(.A(new_n10084), .Y(new_n10265));
  nor_5  g09889(.A(new_n10108), .B(new_n10265), .Y(new_n10266));
  nor_5  g09890(.A(new_n10109), .B(new_n10082), .Y(new_n10267));
  nor_5  g09891(.A(new_n10267), .B(new_n10266), .Y(new_n10268));
  xor_4  g09892(.A(new_n10268), .B(new_n10264), .Y(new_n10269));
  nor_5  g09893(.A(new_n10085), .B(new_n6539), .Y(new_n10270));
  nor_5  g09894(.A(new_n10090), .B(new_n10086), .Y(new_n10271));
  nor_5  g09895(.A(new_n10271), .B(new_n10270), .Y(new_n10272));
  xor_4  g09896(.A(new_n10272), .B(new_n10269), .Y(new_n10273));
  xor_4  g09897(.A(new_n10273), .B(new_n10263), .Y(new_n10274));
  xor_4  g09898(.A(new_n10274), .B(new_n10256), .Y(new_n10275));
  nand_5 g09899(.A(new_n10133), .B(new_n10132), .Y(new_n10276));
  nand_5 g09900(.A(new_n10134), .B(new_n6491), .Y(new_n10277));
  nand_5 g09901(.A(new_n10277), .B(new_n10276), .Y(new_n10278));
  nand_5 g09902(.A(pi042), .B(pi018), .Y(new_n10279));
  nand_5 g09903(.A(new_n10028), .B(new_n10027), .Y(new_n10280));
  nand_5 g09904(.A(new_n10029), .B(new_n6608), .Y(new_n10281));
  nand_5 g09905(.A(new_n10281), .B(new_n10280), .Y(new_n10282));
  nand_5 g09906(.A(pi213), .B(pi126), .Y(new_n10283));
  xor_4  g09907(.A(new_n10283), .B(new_n10282), .Y(new_n10284));
  nand_5 g09908(.A(pi143), .B(pi034), .Y(new_n10285));
  nand_5 g09909(.A(new_n10088), .B(new_n10087), .Y(new_n10286));
  nand_5 g09910(.A(new_n10089), .B(new_n6537), .Y(new_n10287));
  nand_5 g09911(.A(new_n10287), .B(new_n10286), .Y(new_n10288));
  xnor_4 g09912(.A(new_n10288), .B(new_n10285), .Y(new_n10289));
  xor_4  g09913(.A(new_n10289), .B(new_n10284), .Y(new_n10290));
  xor_4  g09914(.A(new_n10290), .B(new_n10279), .Y(new_n10291));
  not_8  g09915(.A(new_n10145), .Y(new_n10292));
  nand_5 g09916(.A(new_n10292), .B(new_n10120), .Y(new_n10293));
  not_8  g09917(.A(new_n10146), .Y(new_n10294));
  nand_5 g09918(.A(new_n10294), .B(new_n10119), .Y(new_n10295));
  nand_5 g09919(.A(new_n10295), .B(new_n10293), .Y(new_n10296));
  nand_5 g09920(.A(pi241), .B(pi038), .Y(new_n10297));
  nand_5 g09921(.A(pi208), .B(pi193), .Y(new_n10298));
  nor_5  g09922(.A(new_n10057), .B(new_n6576), .Y(new_n10299));
  nor_5  g09923(.A(new_n10062), .B(new_n10058), .Y(new_n10300));
  nor_5  g09924(.A(new_n10300), .B(new_n10299), .Y(new_n10301));
  xor_4  g09925(.A(new_n10301), .B(new_n10298), .Y(new_n10302));
  xor_4  g09926(.A(new_n10302), .B(new_n10297), .Y(new_n10303));
  xor_4  g09927(.A(new_n10303), .B(new_n10296), .Y(new_n10304));
  nand_5 g09928(.A(new_n10140), .B(new_n10139), .Y(new_n10305));
  nand_5 g09929(.A(new_n10141), .B(new_n6501), .Y(new_n10306));
  nand_5 g09930(.A(new_n10306), .B(new_n10305), .Y(new_n10307));
  nand_5 g09931(.A(pi105), .B(pi061), .Y(new_n10308));
  xor_4  g09932(.A(new_n10308), .B(new_n10307), .Y(new_n10309));
  nand_5 g09933(.A(pi238), .B(pi139), .Y(new_n10310));
  nand_5 g09934(.A(pi048), .B(pi015), .Y(new_n10311));
  nand_5 g09935(.A(new_n10060), .B(new_n10059), .Y(new_n10312));
  nand_5 g09936(.A(new_n10061), .B(new_n6574), .Y(new_n10313));
  nand_5 g09937(.A(new_n10313), .B(new_n10312), .Y(new_n10314));
  xnor_4 g09938(.A(new_n10314), .B(new_n10311), .Y(new_n10315));
  xor_4  g09939(.A(new_n10315), .B(new_n10310), .Y(new_n10316));
  xor_4  g09940(.A(new_n10316), .B(new_n10309), .Y(new_n10317));
  xor_4  g09941(.A(new_n10317), .B(new_n10304), .Y(new_n10318));
  xor_4  g09942(.A(new_n10318), .B(new_n10291), .Y(new_n10319));
  xor_4  g09943(.A(new_n10319), .B(new_n10278), .Y(new_n10320));
  xor_4  g09944(.A(new_n10320), .B(new_n10275), .Y(new_n10321));
  xor_4  g09945(.A(new_n10321), .B(new_n10251), .Y(new_n10322));
  xor_4  g09946(.A(new_n10322), .B(new_n10237), .Y(po072));
  xor_4  g09947(.A(new_n898), .B(new_n897), .Y(po073));
  xor_4  g09948(.A(new_n6325), .B(new_n6322), .Y(po074));
  xor_4  g09949(.A(new_n7922), .B(new_n7921), .Y(po075));
  xor_4  g09950(.A(new_n6704), .B(new_n6702), .Y(po076));
  xor_4  g09951(.A(new_n1070), .B(new_n1061), .Y(po077));
  xor_4  g09952(.A(new_n1744), .B(new_n1743), .Y(po078));
  xnor_4 g09953(.A(new_n5953), .B(new_n5952), .Y(po079));
  xor_4  g09954(.A(new_n9320), .B(new_n9319), .Y(po080));
  xnor_4 g09955(.A(new_n7917), .B(new_n7916), .Y(po081));
  xor_4  g09956(.A(new_n6327), .B(new_n6318), .Y(po082));
  xnor_4 g09957(.A(new_n1095), .B(new_n1094), .Y(po083));
  nand_5 g09958(.A(pi110), .B(pi107), .Y(new_n10335));
  nand_5 g09959(.A(new_n784), .B(new_n783), .Y(new_n10336));
  nand_5 g09960(.A(new_n785), .B(new_n694), .Y(new_n10337));
  nand_5 g09961(.A(new_n10337), .B(new_n10336), .Y(new_n10338));
  nand_5 g09962(.A(pi063), .B(pi026), .Y(new_n10339));
  not_8  g09963(.A(new_n484), .Y(new_n10340));
  nor_5  g09964(.A(new_n10340), .B(new_n459), .Y(new_n10341));
  nor_5  g09965(.A(new_n485), .B(new_n457), .Y(new_n10342));
  nor_5  g09966(.A(new_n10342), .B(new_n10341), .Y(new_n10343));
  xor_4  g09967(.A(new_n10343), .B(new_n10339), .Y(new_n10344));
  xor_4  g09968(.A(new_n10344), .B(new_n10338), .Y(new_n10345));
  xor_4  g09969(.A(new_n10345), .B(new_n10335), .Y(new_n10346));
  nand_5 g09970(.A(new_n471), .B(new_n470), .Y(new_n10347));
  nand_5 g09971(.A(new_n472), .B(new_n443), .Y(new_n10348));
  nand_5 g09972(.A(new_n10348), .B(new_n10347), .Y(new_n10349));
  nor_5  g09973(.A(new_n481), .B(new_n477), .Y(new_n10350));
  not_8  g09974(.A(new_n474), .Y(new_n10351));
  nor_5  g09975(.A(new_n482), .B(new_n10351), .Y(new_n10352));
  nor_5  g09976(.A(new_n10352), .B(new_n10350), .Y(new_n10353));
  xor_4  g09977(.A(new_n10353), .B(new_n10349), .Y(new_n10354));
  nand_5 g09978(.A(pi200), .B(pi151), .Y(new_n10355));
  nand_5 g09979(.A(pi164), .B(pi000), .Y(new_n10356));
  nand_5 g09980(.A(pi070), .B(pi032), .Y(new_n10357));
  xor_4  g09981(.A(new_n10357), .B(new_n10356), .Y(new_n10358));
  xor_4  g09982(.A(new_n10358), .B(new_n10355), .Y(new_n10359));
  xor_4  g09983(.A(new_n10359), .B(new_n10354), .Y(new_n10360));
  xor_4  g09984(.A(new_n10360), .B(new_n10346), .Y(new_n10361));
  nand_5 g09985(.A(new_n868), .B(new_n486), .Y(new_n10362));
  nand_5 g09986(.A(new_n906), .B(new_n869), .Y(new_n10363));
  nand_5 g09987(.A(new_n10363), .B(new_n10362), .Y(new_n10364));
  nand_5 g09988(.A(pi149), .B(pi075), .Y(new_n10365));
  nand_5 g09989(.A(new_n833), .B(new_n802), .Y(new_n10366));
  nand_5 g09990(.A(new_n838), .B(new_n834), .Y(new_n10367));
  nand_5 g09991(.A(new_n10367), .B(new_n10366), .Y(new_n10368));
  xor_4  g09992(.A(new_n10368), .B(new_n10365), .Y(new_n10369));
  nand_5 g09993(.A(pi166), .B(pi134), .Y(new_n10370));
  nand_5 g09994(.A(pi167), .B(pi097), .Y(new_n10371));
  xor_4  g09995(.A(new_n10371), .B(new_n10370), .Y(new_n10372));
  xor_4  g09996(.A(new_n10372), .B(new_n10369), .Y(new_n10373));
  or_6   g09997(.A(new_n853), .B(new_n546), .Y(new_n10374));
  nand_5 g09998(.A(new_n858), .B(new_n854), .Y(new_n10375));
  nand_5 g09999(.A(new_n10375), .B(new_n10374), .Y(new_n10376));
  nand_5 g10000(.A(new_n856), .B(new_n855), .Y(new_n10377));
  nand_5 g10001(.A(new_n857), .B(new_n544), .Y(new_n10378));
  nand_5 g10002(.A(new_n10378), .B(new_n10377), .Y(new_n10379));
  xor_4  g10003(.A(new_n10379), .B(new_n10376), .Y(new_n10380));
  nand_5 g10004(.A(pi214), .B(pi045), .Y(new_n10381));
  nand_5 g10005(.A(new_n791), .B(new_n790), .Y(new_n10382));
  nand_5 g10006(.A(new_n792), .B(new_n682), .Y(new_n10383));
  nand_5 g10007(.A(new_n10383), .B(new_n10382), .Y(new_n10384));
  not_8  g10008(.A(new_n483), .Y(new_n10385));
  nor_5  g10009(.A(new_n10385), .B(new_n467), .Y(new_n10386));
  nor_5  g10010(.A(new_n10386), .B(new_n466), .Y(new_n10387));
  xor_4  g10011(.A(new_n10387), .B(new_n10384), .Y(new_n10388));
  nor_5  g10012(.A(new_n820), .B(new_n714), .Y(new_n10389));
  nor_5  g10013(.A(new_n821), .B(new_n819), .Y(new_n10390));
  nor_5  g10014(.A(new_n10390), .B(new_n10389), .Y(new_n10391));
  nand_5 g10015(.A(new_n786), .B(new_n782), .Y(new_n10392));
  nand_5 g10016(.A(new_n794), .B(new_n787), .Y(new_n10393));
  nand_5 g10017(.A(new_n10393), .B(new_n10392), .Y(new_n10394));
  xor_4  g10018(.A(new_n10394), .B(new_n10391), .Y(new_n10395));
  xor_4  g10019(.A(new_n10395), .B(new_n10388), .Y(new_n10396));
  xor_4  g10020(.A(new_n10396), .B(new_n10381), .Y(new_n10397));
  nand_5 g10021(.A(pi247), .B(pi044), .Y(new_n10398));
  not_8  g10022(.A(new_n861), .Y(new_n10399));
  nor_5  g10023(.A(new_n10399), .B(new_n840), .Y(new_n10400));
  nor_5  g10024(.A(new_n865), .B(new_n862), .Y(new_n10401));
  nor_5  g10025(.A(new_n10401), .B(new_n10400), .Y(new_n10402));
  xor_4  g10026(.A(new_n10402), .B(new_n10398), .Y(new_n10403));
  nand_5 g10027(.A(new_n479), .B(new_n437), .Y(new_n10404));
  nand_5 g10028(.A(new_n480), .B(new_n478), .Y(new_n10405));
  nand_5 g10029(.A(new_n10405), .B(new_n10404), .Y(new_n10406));
  nand_5 g10030(.A(pi080), .B(pi054), .Y(new_n10407));
  xor_4  g10031(.A(new_n10407), .B(new_n10406), .Y(new_n10408));
  xor_4  g10032(.A(new_n10408), .B(new_n10403), .Y(new_n10409));
  xor_4  g10033(.A(new_n10409), .B(new_n10397), .Y(new_n10410));
  xor_4  g10034(.A(new_n10410), .B(new_n10380), .Y(new_n10411));
  xor_4  g10035(.A(new_n10411), .B(new_n10373), .Y(new_n10412));
  xor_4  g10036(.A(new_n10412), .B(new_n10364), .Y(new_n10413));
  nor_5  g10037(.A(new_n866), .B(new_n839), .Y(new_n10414));
  nor_5  g10038(.A(new_n867), .B(new_n775), .Y(new_n10415));
  or_6   g10039(.A(new_n10415), .B(new_n10414), .Y(new_n10416));
  nand_5 g10040(.A(pi083), .B(pi027), .Y(new_n10417));
  nand_5 g10041(.A(pi228), .B(pi114), .Y(new_n10418));
  nand_5 g10042(.A(new_n809), .B(new_n808), .Y(new_n10419));
  nand_5 g10043(.A(new_n810), .B(new_n724), .Y(new_n10420));
  nand_5 g10044(.A(new_n10420), .B(new_n10419), .Y(new_n10421));
  nand_5 g10045(.A(pi096), .B(pi049), .Y(new_n10422));
  nand_5 g10046(.A(pi246), .B(pi039), .Y(new_n10423));
  xor_4  g10047(.A(new_n10423), .B(new_n10422), .Y(new_n10424));
  xor_4  g10048(.A(new_n10424), .B(new_n10421), .Y(new_n10425));
  xor_4  g10049(.A(new_n10425), .B(new_n10418), .Y(new_n10426));
  xor_4  g10050(.A(new_n10426), .B(new_n10417), .Y(new_n10427));
  or_6   g10051(.A(new_n788), .B(new_n684), .Y(new_n10428));
  not_8  g10052(.A(new_n793), .Y(new_n10429));
  nand_5 g10053(.A(new_n10429), .B(new_n789), .Y(new_n10430));
  nand_5 g10054(.A(new_n10430), .B(new_n10428), .Y(new_n10431));
  nand_5 g10055(.A(pi245), .B(pi136), .Y(new_n10432));
  xor_4  g10056(.A(new_n10432), .B(new_n10431), .Y(new_n10433));
  nand_5 g10057(.A(pi103), .B(pi009), .Y(new_n10434));
  nand_5 g10058(.A(new_n817), .B(new_n816), .Y(new_n10435));
  nand_5 g10059(.A(new_n818), .B(new_n712), .Y(new_n10436));
  nand_5 g10060(.A(new_n10436), .B(new_n10435), .Y(new_n10437));
  nand_5 g10061(.A(pi201), .B(pi056), .Y(new_n10438));
  xnor_4 g10062(.A(new_n10438), .B(new_n10437), .Y(new_n10439));
  xor_4  g10063(.A(new_n10439), .B(new_n10434), .Y(new_n10440));
  xor_4  g10064(.A(new_n10440), .B(new_n10433), .Y(new_n10441));
  xor_4  g10065(.A(new_n10441), .B(new_n10427), .Y(new_n10442));
  xor_4  g10066(.A(new_n10442), .B(new_n10416), .Y(new_n10443));
  xor_4  g10067(.A(new_n10443), .B(new_n10413), .Y(new_n10444));
  nand_5 g10068(.A(new_n851), .B(new_n847), .Y(new_n10445));
  nand_5 g10069(.A(new_n859), .B(new_n852), .Y(new_n10446));
  nand_5 g10070(.A(new_n10446), .B(new_n10445), .Y(new_n10447));
  nand_5 g10071(.A(pi202), .B(pi119), .Y(new_n10448));
  xor_4  g10072(.A(new_n10448), .B(new_n10447), .Y(new_n10449));
  nand_5 g10073(.A(pi181), .B(pi019), .Y(new_n10450));
  nor_5  g10074(.A(new_n468), .B(new_n445), .Y(new_n10451));
  nor_5  g10075(.A(new_n473), .B(new_n469), .Y(new_n10452));
  nor_5  g10076(.A(new_n10452), .B(new_n10451), .Y(new_n10453));
  xor_4  g10077(.A(new_n10453), .B(new_n10450), .Y(new_n10454));
  nand_5 g10078(.A(pi072), .B(pi016), .Y(new_n10455));
  nand_5 g10079(.A(pi248), .B(pi117), .Y(new_n10456));
  xor_4  g10080(.A(new_n10456), .B(new_n10455), .Y(new_n10457));
  nand_5 g10081(.A(new_n825), .B(new_n725), .Y(new_n10458));
  nand_5 g10082(.A(new_n828), .B(new_n823), .Y(new_n10459));
  nand_5 g10083(.A(new_n10459), .B(new_n10458), .Y(new_n10460));
  xor_4  g10084(.A(new_n10460), .B(new_n10457), .Y(new_n10461));
  xor_4  g10085(.A(new_n10461), .B(new_n10454), .Y(new_n10462));
  xor_4  g10086(.A(new_n10462), .B(new_n10449), .Y(new_n10463));
  xor_4  g10087(.A(new_n10463), .B(new_n10444), .Y(new_n10464));
  nand_5 g10088(.A(pi240), .B(pi093), .Y(new_n10465));
  nand_5 g10089(.A(pi250), .B(pi234), .Y(new_n10466));
  xor_4  g10090(.A(new_n10466), .B(new_n10465), .Y(new_n10467));
  nand_5 g10091(.A(new_n800), .B(new_n779), .Y(new_n10468));
  or_6   g10092(.A(new_n801), .B(new_n778), .Y(new_n10469));
  nand_5 g10093(.A(new_n10469), .B(new_n10468), .Y(new_n10470));
  nand_5 g10094(.A(pi175), .B(pi011), .Y(new_n10471));
  xor_4  g10095(.A(new_n10471), .B(new_n10470), .Y(new_n10472));
  nand_5 g10096(.A(new_n842), .B(new_n538), .Y(new_n10473));
  or_6   g10097(.A(new_n860), .B(new_n844), .Y(new_n10474));
  nand_5 g10098(.A(new_n10474), .B(new_n10473), .Y(new_n10475));
  xor_4  g10099(.A(new_n10475), .B(new_n10472), .Y(new_n10476));
  nand_5 g10100(.A(new_n814), .B(new_n811), .Y(new_n10477));
  nand_5 g10101(.A(new_n822), .B(new_n815), .Y(new_n10478));
  nand_5 g10102(.A(new_n10478), .B(new_n10477), .Y(new_n10479));
  nand_5 g10103(.A(pi203), .B(pi147), .Y(new_n10480));
  xor_4  g10104(.A(new_n10480), .B(new_n10479), .Y(new_n10481));
  xor_4  g10105(.A(new_n10481), .B(new_n10476), .Y(new_n10482));
  nand_5 g10106(.A(pi148), .B(pi091), .Y(new_n10483));
  nand_5 g10107(.A(pi145), .B(pi116), .Y(new_n10484));
  xor_4  g10108(.A(new_n10484), .B(new_n10483), .Y(new_n10485));
  xor_4  g10109(.A(new_n10485), .B(new_n10482), .Y(new_n10486));
  nand_5 g10110(.A(pi206), .B(pi115), .Y(new_n10487));
  nand_5 g10111(.A(pi156), .B(pi008), .Y(new_n10488));
  nand_5 g10112(.A(new_n831), .B(new_n805), .Y(new_n10489));
  nand_5 g10113(.A(new_n10489), .B(new_n830), .Y(new_n10490));
  or_6   g10114(.A(new_n798), .B(new_n696), .Y(new_n10491));
  nand_5 g10115(.A(new_n799), .B(new_n795), .Y(new_n10492));
  nand_5 g10116(.A(new_n10492), .B(new_n10491), .Y(new_n10493));
  nand_5 g10117(.A(pi235), .B(pi171), .Y(new_n10494));
  xor_4  g10118(.A(new_n10494), .B(new_n10493), .Y(new_n10495));
  xor_4  g10119(.A(new_n10495), .B(new_n10490), .Y(new_n10496));
  xor_4  g10120(.A(new_n10496), .B(new_n10488), .Y(new_n10497));
  xor_4  g10121(.A(new_n10497), .B(new_n10487), .Y(new_n10498));
  xor_4  g10122(.A(new_n10498), .B(new_n10486), .Y(new_n10499));
  nand_5 g10123(.A(new_n849), .B(new_n848), .Y(new_n10500));
  nand_5 g10124(.A(new_n850), .B(new_n537), .Y(new_n10501));
  nand_5 g10125(.A(new_n10501), .B(new_n10500), .Y(new_n10502));
  nand_5 g10126(.A(pi163), .B(pi031), .Y(new_n10503));
  xor_4  g10127(.A(new_n10503), .B(new_n10502), .Y(new_n10504));
  xor_4  g10128(.A(new_n10504), .B(new_n10499), .Y(new_n10505));
  xor_4  g10129(.A(new_n10505), .B(new_n10467), .Y(new_n10506));
  xor_4  g10130(.A(new_n10506), .B(new_n10464), .Y(new_n10507));
  xor_4  g10131(.A(new_n10507), .B(new_n10361), .Y(po084));
  xor_4  g10132(.A(new_n10153), .B(new_n10152), .Y(po085));
  not_8  g10133(.A(new_n9792), .Y(new_n10510));
  nand_5 g10134(.A(new_n9796), .B(new_n10510), .Y(new_n10511));
  or_6   g10135(.A(new_n9797), .B(new_n9762), .Y(new_n10512));
  nand_5 g10136(.A(new_n10512), .B(new_n10511), .Y(new_n10513));
  nand_5 g10137(.A(pi241), .B(pi021), .Y(new_n10514));
  nand_5 g10138(.A(pi217), .B(pi034), .Y(new_n10515));
  xor_4  g10139(.A(new_n10515), .B(new_n10514), .Y(new_n10516));
  xor_4  g10140(.A(new_n10516), .B(new_n10513), .Y(new_n10517));
  nand_5 g10141(.A(new_n9749), .B(new_n9745), .Y(new_n10518));
  not_8  g10142(.A(new_n9742), .Y(new_n10519));
  nand_5 g10143(.A(new_n9750), .B(new_n10519), .Y(new_n10520));
  nand_5 g10144(.A(new_n10520), .B(new_n10518), .Y(new_n10521));
  nand_5 g10145(.A(pi232), .B(pi212), .Y(new_n10522));
  xor_4  g10146(.A(new_n10522), .B(new_n10521), .Y(new_n10523));
  nand_5 g10147(.A(new_n9747), .B(new_n9746), .Y(new_n10524));
  nand_5 g10148(.A(new_n9748), .B(new_n9625), .Y(new_n10525));
  nand_5 g10149(.A(new_n10525), .B(new_n10524), .Y(new_n10526));
  nand_5 g10150(.A(pi127), .B(pi104), .Y(new_n10527));
  xor_4  g10151(.A(new_n10527), .B(new_n10526), .Y(new_n10528));
  nand_5 g10152(.A(new_n9739), .B(new_n9738), .Y(new_n10529));
  nand_5 g10153(.A(new_n9740), .B(new_n9635), .Y(new_n10530));
  nand_5 g10154(.A(new_n10530), .B(new_n10529), .Y(new_n10531));
  nand_5 g10155(.A(pi224), .B(pi112), .Y(new_n10532));
  xor_4  g10156(.A(new_n10532), .B(new_n10531), .Y(new_n10533));
  xor_4  g10157(.A(new_n10533), .B(new_n10528), .Y(new_n10534));
  xor_4  g10158(.A(new_n10534), .B(new_n10523), .Y(new_n10535));
  xor_4  g10159(.A(new_n10535), .B(new_n10517), .Y(new_n10536));
  nand_5 g10160(.A(pi255), .B(pi013), .Y(new_n10537));
  nand_5 g10161(.A(pi252), .B(pi047), .Y(new_n10538));
  nand_5 g10162(.A(pi131), .B(pi129), .Y(new_n10539));
  nand_5 g10163(.A(pi236), .B(pi082), .Y(new_n10540));
  xor_4  g10164(.A(new_n10540), .B(new_n10539), .Y(new_n10541));
  nand_5 g10165(.A(pi161), .B(pi005), .Y(new_n10542));
  xor_4  g10166(.A(new_n10542), .B(new_n10541), .Y(new_n10543));
  xor_4  g10167(.A(new_n10543), .B(new_n10538), .Y(new_n10544));
  xor_4  g10168(.A(new_n10544), .B(new_n10537), .Y(new_n10545));
  nor_5  g10169(.A(new_n9719), .B(new_n9715), .Y(new_n10546));
  not_8  g10170(.A(new_n9712), .Y(new_n10547));
  nor_5  g10171(.A(new_n9720), .B(new_n10547), .Y(new_n10548));
  nor_5  g10172(.A(new_n10548), .B(new_n10546), .Y(new_n10549));
  nor_5  g10173(.A(new_n9723), .B(new_n9696), .Y(new_n10550));
  and_6  g10174(.A(new_n9724), .B(new_n9695), .Y(new_n10551));
  nor_5  g10175(.A(new_n10551), .B(new_n10550), .Y(new_n10552));
  xor_4  g10176(.A(new_n10552), .B(new_n10549), .Y(new_n10553));
  xor_4  g10177(.A(new_n10553), .B(new_n10545), .Y(new_n10554));
  xor_4  g10178(.A(new_n10554), .B(new_n10536), .Y(new_n10555));
  or_6   g10179(.A(new_n9722), .B(new_n9705), .Y(new_n10556));
  nand_5 g10180(.A(new_n10556), .B(new_n9704), .Y(new_n10557));
  nand_5 g10181(.A(pi227), .B(pi064), .Y(new_n10558));
  nand_5 g10182(.A(pi105), .B(pi024), .Y(new_n10559));
  xor_4  g10183(.A(new_n10559), .B(new_n10558), .Y(new_n10560));
  xor_4  g10184(.A(new_n10560), .B(new_n10557), .Y(new_n10561));
  xor_4  g10185(.A(new_n10561), .B(new_n10555), .Y(new_n10562));
  nor_5  g10186(.A(new_n9736), .B(new_n9637), .Y(new_n10563));
  nor_5  g10187(.A(new_n9741), .B(new_n9737), .Y(new_n10564));
  nor_5  g10188(.A(new_n10564), .B(new_n10563), .Y(new_n10565));
  or_6   g10189(.A(new_n9827), .B(new_n9798), .Y(new_n10566));
  nand_5 g10190(.A(new_n9828), .B(new_n9690), .Y(new_n10567));
  nand_5 g10191(.A(new_n10567), .B(new_n10566), .Y(new_n10568));
  xor_4  g10192(.A(new_n10568), .B(new_n10565), .Y(new_n10569));
  nand_5 g10193(.A(pi121), .B(pi090), .Y(new_n10570));
  nand_5 g10194(.A(new_n9709), .B(new_n9708), .Y(new_n10571));
  nand_5 g10195(.A(new_n9710), .B(new_n9671), .Y(new_n10572));
  nand_5 g10196(.A(new_n10572), .B(new_n10571), .Y(new_n10573));
  nand_5 g10197(.A(new_n9809), .B(new_n9808), .Y(new_n10574));
  nand_5 g10198(.A(new_n9810), .B(new_n9561), .Y(new_n10575));
  nand_5 g10199(.A(new_n10575), .B(new_n10574), .Y(new_n10576));
  xnor_4 g10200(.A(new_n10576), .B(new_n10573), .Y(new_n10577));
  xor_4  g10201(.A(new_n10577), .B(new_n10570), .Y(new_n10578));
  xor_4  g10202(.A(new_n10578), .B(new_n10569), .Y(new_n10579));
  nand_5 g10203(.A(new_n9806), .B(new_n9552), .Y(new_n10580));
  nand_5 g10204(.A(new_n9824), .B(new_n9807), .Y(new_n10581));
  nand_5 g10205(.A(new_n10581), .B(new_n10580), .Y(new_n10582));
  nand_5 g10206(.A(new_n9770), .B(new_n9769), .Y(new_n10583));
  nand_5 g10207(.A(new_n9771), .B(new_n9607), .Y(new_n10584));
  nand_5 g10208(.A(new_n10584), .B(new_n10583), .Y(new_n10585));
  nand_5 g10209(.A(pi249), .B(pi152), .Y(new_n10586));
  xnor_4 g10210(.A(new_n10586), .B(new_n10585), .Y(new_n10587));
  xor_4  g10211(.A(new_n10587), .B(new_n10582), .Y(new_n10588));
  nand_5 g10212(.A(new_n9608), .B(new_n9785), .Y(new_n10589));
  nand_5 g10213(.A(new_n9788), .B(new_n9784), .Y(new_n10590));
  nand_5 g10214(.A(new_n10590), .B(new_n10589), .Y(new_n10591));
  nand_5 g10215(.A(pi231), .B(pi141), .Y(new_n10592));
  nand_5 g10216(.A(pi183), .B(pi111), .Y(new_n10593));
  xor_4  g10217(.A(new_n10593), .B(new_n10592), .Y(new_n10594));
  nand_5 g10218(.A(pi189), .B(pi081), .Y(new_n10595));
  xor_4  g10219(.A(new_n10595), .B(new_n10594), .Y(new_n10596));
  xor_4  g10220(.A(new_n10596), .B(new_n10591), .Y(new_n10597));
  xor_4  g10221(.A(new_n10597), .B(new_n10588), .Y(new_n10598));
  nand_5 g10222(.A(pi233), .B(pi077), .Y(new_n10599));
  or_6   g10223(.A(new_n9825), .B(new_n9803), .Y(new_n10600));
  not_8  g10224(.A(new_n9800), .Y(new_n10601));
  nand_5 g10225(.A(new_n9826), .B(new_n10601), .Y(new_n10602));
  nand_5 g10226(.A(new_n10602), .B(new_n10600), .Y(new_n10603));
  nand_5 g10227(.A(new_n9775), .B(new_n9772), .Y(new_n10604));
  not_8  g10228(.A(new_n9783), .Y(new_n10605));
  nand_5 g10229(.A(new_n10605), .B(new_n9776), .Y(new_n10606));
  nand_5 g10230(.A(new_n10606), .B(new_n10604), .Y(new_n10607));
  nor_5  g10231(.A(new_n9777), .B(new_n9596), .Y(new_n10608));
  nor_5  g10232(.A(new_n9782), .B(new_n9778), .Y(new_n10609));
  nor_5  g10233(.A(new_n10609), .B(new_n10608), .Y(new_n10610));
  xor_4  g10234(.A(new_n10610), .B(new_n10607), .Y(new_n10611));
  xor_4  g10235(.A(new_n10611), .B(new_n10603), .Y(new_n10612));
  nand_5 g10236(.A(pi222), .B(pi146), .Y(new_n10613));
  nand_5 g10237(.A(pi204), .B(pi125), .Y(new_n10614));
  nor_5  g10238(.A(new_n9753), .B(new_n9730), .Y(new_n10615));
  nor_5  g10239(.A(new_n10615), .B(new_n9754), .Y(new_n10616));
  xor_4  g10240(.A(new_n10616), .B(new_n10614), .Y(new_n10617));
  xor_4  g10241(.A(new_n10617), .B(new_n10613), .Y(new_n10618));
  xor_4  g10242(.A(new_n10618), .B(new_n10612), .Y(new_n10619));
  xor_4  g10243(.A(new_n10619), .B(new_n10599), .Y(new_n10620));
  xor_4  g10244(.A(new_n10620), .B(new_n10598), .Y(new_n10621));
  nand_5 g10245(.A(pi208), .B(pi157), .Y(new_n10622));
  nand_5 g10246(.A(new_n9780), .B(new_n9779), .Y(new_n10623));
  nand_5 g10247(.A(new_n9781), .B(new_n9594), .Y(new_n10624));
  nand_5 g10248(.A(new_n10624), .B(new_n10623), .Y(new_n10625));
  xor_4  g10249(.A(new_n10625), .B(new_n10622), .Y(new_n10626));
  nand_5 g10250(.A(pi168), .B(pi017), .Y(new_n10627));
  nand_5 g10251(.A(pi213), .B(pi191), .Y(new_n10628));
  xor_4  g10252(.A(new_n10628), .B(new_n10627), .Y(new_n10629));
  nand_5 g10253(.A(pi140), .B(pi018), .Y(new_n10630));
  nand_5 g10254(.A(pi187), .B(pi052), .Y(new_n10631));
  nand_5 g10255(.A(pi100), .B(pi084), .Y(new_n10632));
  xor_4  g10256(.A(new_n10632), .B(new_n10631), .Y(new_n10633));
  nor_5  g10257(.A(new_n9734), .B(new_n9626), .Y(new_n10634));
  and_6  g10258(.A(new_n9751), .B(new_n9735), .Y(new_n10635));
  nor_5  g10259(.A(new_n10635), .B(new_n10634), .Y(new_n10636));
  nand_5 g10260(.A(pi176), .B(pi015), .Y(new_n10637));
  xor_4  g10261(.A(new_n10637), .B(new_n10636), .Y(new_n10638));
  xor_4  g10262(.A(new_n10638), .B(new_n10633), .Y(new_n10639));
  xor_4  g10263(.A(new_n10639), .B(new_n10630), .Y(new_n10640));
  xor_4  g10264(.A(new_n10640), .B(new_n10629), .Y(new_n10641));
  nand_5 g10265(.A(new_n9822), .B(new_n9818), .Y(new_n10642));
  nand_5 g10266(.A(new_n9823), .B(new_n9815), .Y(new_n10643));
  nand_5 g10267(.A(new_n10643), .B(new_n10642), .Y(new_n10644));
  nand_5 g10268(.A(pi040), .B(pi035), .Y(new_n10645));
  nor_5  g10269(.A(new_n9812), .B(new_n9563), .Y(new_n10646));
  nor_5  g10270(.A(new_n9813), .B(new_n9811), .Y(new_n10647));
  or_6   g10271(.A(new_n10647), .B(new_n10646), .Y(new_n10648));
  xor_4  g10272(.A(new_n10648), .B(new_n10645), .Y(new_n10649));
  xor_4  g10273(.A(new_n10649), .B(new_n10644), .Y(new_n10650));
  xor_4  g10274(.A(new_n10650), .B(new_n10641), .Y(new_n10651));
  xor_4  g10275(.A(new_n10651), .B(new_n10626), .Y(new_n10652));
  nand_5 g10276(.A(pi174), .B(pi139), .Y(new_n10653));
  nand_5 g10277(.A(pi133), .B(pi106), .Y(new_n10654));
  xor_4  g10278(.A(new_n10654), .B(new_n10653), .Y(new_n10655));
  nand_5 g10279(.A(pi242), .B(pi128), .Y(new_n10656));
  nand_5 g10280(.A(new_n9717), .B(new_n9716), .Y(new_n10657));
  nand_5 g10281(.A(new_n9718), .B(new_n9661), .Y(new_n10658));
  nand_5 g10282(.A(new_n10658), .B(new_n10657), .Y(new_n10659));
  nand_5 g10283(.A(new_n9820), .B(new_n9819), .Y(new_n10660));
  nand_5 g10284(.A(new_n9821), .B(new_n9550), .Y(new_n10661));
  nand_5 g10285(.A(new_n10661), .B(new_n10660), .Y(new_n10662));
  xnor_4 g10286(.A(new_n10662), .B(new_n10659), .Y(new_n10663));
  xor_4  g10287(.A(new_n10663), .B(new_n10656), .Y(new_n10664));
  xor_4  g10288(.A(new_n10664), .B(new_n10655), .Y(new_n10665));
  or_6   g10289(.A(new_n9756), .B(new_n9725), .Y(new_n10666));
  nand_5 g10290(.A(new_n9761), .B(new_n9757), .Y(new_n10667));
  nand_5 g10291(.A(new_n10667), .B(new_n10666), .Y(new_n10668));
  nor_5  g10292(.A(new_n9706), .B(new_n9673), .Y(new_n10669));
  nor_5  g10293(.A(new_n9711), .B(new_n9707), .Y(new_n10670));
  nor_5  g10294(.A(new_n10670), .B(new_n10669), .Y(new_n10671));
  nand_5 g10295(.A(pi210), .B(pi088), .Y(new_n10672));
  xor_4  g10296(.A(new_n10672), .B(new_n10671), .Y(new_n10673));
  xor_4  g10297(.A(new_n10673), .B(new_n10668), .Y(new_n10674));
  xor_4  g10298(.A(new_n10674), .B(new_n10665), .Y(new_n10675));
  xor_4  g10299(.A(new_n10675), .B(new_n10652), .Y(new_n10676));
  xor_4  g10300(.A(new_n10676), .B(new_n10621), .Y(new_n10677));
  nor_5  g10301(.A(new_n9790), .B(new_n9768), .Y(new_n10678));
  not_8  g10302(.A(new_n9791), .Y(new_n10679));
  nor_5  g10303(.A(new_n10679), .B(new_n9766), .Y(new_n10680));
  nor_5  g10304(.A(new_n10680), .B(new_n10678), .Y(new_n10681));
  xor_4  g10305(.A(new_n10681), .B(new_n10677), .Y(new_n10682));
  xor_4  g10306(.A(new_n10682), .B(new_n10579), .Y(new_n10683));
  xor_4  g10307(.A(new_n10683), .B(new_n10562), .Y(po086));
  xor_4  g10308(.A(new_n7910), .B(new_n7908), .Y(po087));
  xor_4  g10309(.A(new_n4780), .B(new_n4778), .Y(po088));
  xor_4  g10310(.A(new_n2989), .B(new_n2925), .Y(po089));
  xor_4  g10311(.A(new_n2568), .B(new_n2566), .Y(po090));
  xor_4  g10312(.A(new_n3540), .B(new_n3538), .Y(po091));
  xnor_4 g10313(.A(new_n5956), .B(new_n5955), .Y(po092));
  xor_4  g10314(.A(new_n9341), .B(new_n9340), .Y(po093));
  xnor_4 g10315(.A(new_n904), .B(new_n903), .Y(po094));
  xor_4  g10316(.A(new_n1049), .B(new_n1048), .Y(po095));
  xor_4  g10317(.A(new_n3547), .B(new_n3546), .Y(po096));
  nand_5 g10318(.A(pi173), .B(pi047), .Y(new_n10695));
  nand_5 g10319(.A(pi189), .B(pi150), .Y(new_n10696));
  nand_5 g10320(.A(pi211), .B(pi015), .Y(new_n10697));
  xor_4  g10321(.A(new_n10697), .B(new_n10696), .Y(new_n10698));
  nand_5 g10322(.A(pi196), .B(pi077), .Y(new_n10699));
  nand_5 g10323(.A(pi018), .B(pi014), .Y(new_n10700));
  xnor_4 g10324(.A(new_n10700), .B(new_n10699), .Y(new_n10701));
  xor_4  g10325(.A(new_n10701), .B(new_n10698), .Y(new_n10702));
  xor_4  g10326(.A(new_n10702), .B(new_n10695), .Y(new_n10703));
  or_6   g10327(.A(new_n5397), .B(new_n5368), .Y(new_n10704));
  not_8  g10328(.A(new_n5402), .Y(new_n10705));
  nand_5 g10329(.A(new_n10705), .B(new_n5398), .Y(new_n10706));
  nand_5 g10330(.A(new_n10706), .B(new_n10704), .Y(new_n10707));
  nand_5 g10331(.A(pi084), .B(pi069), .Y(new_n10708));
  nand_5 g10332(.A(pi236), .B(pi205), .Y(new_n10709));
  xor_4  g10333(.A(new_n10709), .B(new_n10708), .Y(new_n10710));
  xor_4  g10334(.A(new_n10710), .B(new_n10707), .Y(new_n10711));
  nand_5 g10335(.A(pi239), .B(pi212), .Y(new_n10712));
  nand_5 g10336(.A(pi104), .B(pi025), .Y(new_n10713));
  xor_4  g10337(.A(new_n10713), .B(new_n10712), .Y(new_n10714));
  xor_4  g10338(.A(new_n10714), .B(new_n10711), .Y(new_n10715));
  xor_4  g10339(.A(new_n10715), .B(new_n10703), .Y(new_n10716));
  nor_5  g10340(.A(new_n5128), .B(new_n5110), .Y(new_n10717));
  nor_5  g10341(.A(new_n5133), .B(new_n5129), .Y(new_n10718));
  nor_5  g10342(.A(new_n10718), .B(new_n10717), .Y(new_n10719));
  nor_5  g10343(.A(new_n5330), .B(new_n5307), .Y(new_n10720));
  and_6  g10344(.A(new_n5331), .B(new_n5296), .Y(new_n10721));
  nor_5  g10345(.A(new_n10721), .B(new_n10720), .Y(new_n10722));
  xor_4  g10346(.A(new_n10722), .B(new_n10719), .Y(new_n10723));
  nand_5 g10347(.A(pi244), .B(pi064), .Y(new_n10724));
  nand_5 g10348(.A(new_n5310), .B(new_n5275), .Y(new_n10725));
  not_8  g10349(.A(new_n5312), .Y(new_n10726));
  nand_5 g10350(.A(new_n5328), .B(new_n10726), .Y(new_n10727));
  nand_5 g10351(.A(new_n10727), .B(new_n10725), .Y(new_n10728));
  nand_5 g10352(.A(new_n5395), .B(new_n5392), .Y(new_n10729));
  nand_5 g10353(.A(new_n5403), .B(new_n5396), .Y(new_n10730));
  nand_5 g10354(.A(new_n10730), .B(new_n10729), .Y(new_n10731));
  nand_5 g10355(.A(pi186), .B(pi146), .Y(new_n10732));
  nand_5 g10356(.A(new_n5390), .B(new_n5389), .Y(new_n10733));
  nand_5 g10357(.A(new_n5391), .B(new_n5353), .Y(new_n10734));
  nand_5 g10358(.A(new_n10734), .B(new_n10733), .Y(new_n10735));
  xor_4  g10359(.A(new_n10735), .B(new_n10732), .Y(new_n10736));
  xor_4  g10360(.A(new_n10736), .B(new_n10731), .Y(new_n10737));
  xor_4  g10361(.A(new_n10737), .B(new_n10728), .Y(new_n10738));
  nand_5 g10362(.A(pi168), .B(pi037), .Y(new_n10739));
  nand_5 g10363(.A(pi152), .B(pi132), .Y(new_n10740));
  xor_4  g10364(.A(new_n10740), .B(new_n10739), .Y(new_n10741));
  xor_4  g10365(.A(new_n10741), .B(new_n10738), .Y(new_n10742));
  xor_4  g10366(.A(new_n10742), .B(new_n10724), .Y(new_n10743));
  nand_5 g10367(.A(pi199), .B(pi035), .Y(new_n10744));
  not_8  g10368(.A(new_n5315), .Y(new_n10745));
  nor_5  g10369(.A(new_n5319), .B(new_n10745), .Y(new_n10746));
  nor_5  g10370(.A(new_n5327), .B(new_n5320), .Y(new_n10747));
  nor_5  g10371(.A(new_n10747), .B(new_n10746), .Y(new_n10748));
  xor_4  g10372(.A(new_n10748), .B(new_n10744), .Y(new_n10749));
  nand_5 g10373(.A(pi184), .B(pi052), .Y(new_n10750));
  xor_4  g10374(.A(new_n10750), .B(new_n10749), .Y(new_n10751));
  xor_4  g10375(.A(new_n10751), .B(new_n10743), .Y(new_n10752));
  xor_4  g10376(.A(new_n10752), .B(new_n10723), .Y(new_n10753));
  or_6   g10377(.A(new_n5233), .B(new_n5207), .Y(new_n10754));
  nand_5 g10378(.A(new_n5234), .B(new_n5206), .Y(new_n10755));
  nand_5 g10379(.A(new_n10755), .B(new_n10754), .Y(new_n10756));
  nand_5 g10380(.A(pi112), .B(pi055), .Y(new_n10757));
  not_8  g10381(.A(new_n5225), .Y(new_n10758));
  nor_5  g10382(.A(new_n5229), .B(new_n10758), .Y(new_n10759));
  nor_5  g10383(.A(new_n5230), .B(new_n5222), .Y(new_n10760));
  nor_5  g10384(.A(new_n10760), .B(new_n10759), .Y(new_n10761));
  nand_5 g10385(.A(new_n5227), .B(new_n5226), .Y(new_n10762));
  nand_5 g10386(.A(new_n5228), .B(new_n5179), .Y(new_n10763));
  nand_5 g10387(.A(new_n10763), .B(new_n10762), .Y(new_n10764));
  xor_4  g10388(.A(new_n10764), .B(new_n10761), .Y(new_n10765));
  xor_4  g10389(.A(new_n10765), .B(new_n10757), .Y(new_n10766));
  xor_4  g10390(.A(new_n10766), .B(new_n10756), .Y(new_n10767));
  nor_5  g10391(.A(new_n5429), .B(new_n5349), .Y(new_n10768));
  nor_5  g10392(.A(new_n5446), .B(new_n5430), .Y(new_n10769));
  nor_5  g10393(.A(new_n10769), .B(new_n10768), .Y(new_n10770));
  xor_4  g10394(.A(new_n10770), .B(new_n10767), .Y(new_n10771));
  xor_4  g10395(.A(new_n10771), .B(new_n10753), .Y(new_n10772));
  xor_4  g10396(.A(new_n10772), .B(new_n10716), .Y(new_n10773));
  nand_5 g10397(.A(pi195), .B(pi139), .Y(new_n10774));
  nand_5 g10398(.A(new_n5400), .B(new_n5399), .Y(new_n10775));
  nand_5 g10399(.A(new_n5401), .B(new_n5366), .Y(new_n10776));
  nand_5 g10400(.A(new_n10776), .B(new_n10775), .Y(new_n10777));
  xor_4  g10401(.A(new_n10777), .B(new_n10774), .Y(new_n10778));
  nand_5 g10402(.A(pi226), .B(pi088), .Y(new_n10779));
  or_6   g10403(.A(new_n5232), .B(new_n5214), .Y(new_n10780));
  nand_5 g10404(.A(new_n10780), .B(new_n5213), .Y(new_n10781));
  nand_5 g10405(.A(new_n5131), .B(new_n5130), .Y(new_n10782));
  nand_5 g10406(.A(new_n5132), .B(new_n5108), .Y(new_n10783));
  nand_5 g10407(.A(new_n10783), .B(new_n10782), .Y(new_n10784));
  xor_4  g10408(.A(new_n10784), .B(new_n10781), .Y(new_n10785));
  nor_5  g10409(.A(new_n5235), .B(new_n5152), .Y(new_n10786));
  nor_5  g10410(.A(new_n5250), .B(new_n5236), .Y(new_n10787));
  nor_5  g10411(.A(new_n10787), .B(new_n10786), .Y(new_n10788));
  xor_4  g10412(.A(new_n10788), .B(new_n10785), .Y(new_n10789));
  xor_4  g10413(.A(new_n10789), .B(new_n10779), .Y(new_n10790));
  xor_4  g10414(.A(new_n10790), .B(new_n10778), .Y(new_n10791));
  nand_5 g10415(.A(new_n5141), .B(new_n5137), .Y(new_n10792));
  or_6   g10416(.A(new_n5143), .B(new_n5134), .Y(new_n10793));
  nand_5 g10417(.A(new_n10793), .B(new_n10792), .Y(new_n10794));
  nand_5 g10418(.A(pi243), .B(pi213), .Y(new_n10795));
  xor_4  g10419(.A(new_n10795), .B(new_n10794), .Y(new_n10796));
  nand_5 g10420(.A(new_n5385), .B(new_n5355), .Y(new_n10797));
  or_6   g10421(.A(new_n5404), .B(new_n5388), .Y(new_n10798));
  nand_5 g10422(.A(new_n10798), .B(new_n10797), .Y(new_n10799));
  nand_5 g10423(.A(pi218), .B(pi208), .Y(new_n10800));
  nor_5  g10424(.A(new_n5321), .B(new_n5286), .Y(new_n10801));
  nor_5  g10425(.A(new_n5326), .B(new_n5322), .Y(new_n10802));
  nor_5  g10426(.A(new_n10802), .B(new_n10801), .Y(new_n10803));
  xor_4  g10427(.A(new_n10803), .B(new_n10800), .Y(new_n10804));
  xor_4  g10428(.A(new_n10804), .B(new_n10799), .Y(new_n10805));
  nand_5 g10429(.A(new_n5417), .B(new_n5405), .Y(new_n10806));
  nand_5 g10430(.A(new_n5428), .B(new_n5418), .Y(new_n10807));
  nand_5 g10431(.A(new_n10807), .B(new_n10806), .Y(new_n10808));
  and_6  g10432(.A(new_n5147), .B(new_n5102), .Y(new_n10809));
  nor_5  g10433(.A(new_n5149), .B(new_n5144), .Y(new_n10810));
  nor_5  g10434(.A(new_n10810), .B(new_n10809), .Y(new_n10811));
  nand_5 g10435(.A(pi034), .B(pi029), .Y(new_n10812));
  nand_5 g10436(.A(pi253), .B(pi161), .Y(new_n10813));
  xor_4  g10437(.A(new_n10813), .B(new_n10812), .Y(new_n10814));
  xor_4  g10438(.A(new_n10814), .B(new_n10811), .Y(new_n10815));
  xor_4  g10439(.A(new_n10815), .B(new_n10808), .Y(new_n10816));
  nand_5 g10440(.A(pi241), .B(pi074), .Y(new_n10817));
  nand_5 g10441(.A(pi207), .B(pi183), .Y(new_n10818));
  xor_4  g10442(.A(new_n10818), .B(new_n10817), .Y(new_n10819));
  nand_5 g10443(.A(pi105), .B(pi066), .Y(new_n10820));
  xor_4  g10444(.A(new_n10820), .B(new_n10819), .Y(new_n10821));
  xor_4  g10445(.A(new_n10821), .B(new_n10816), .Y(new_n10822));
  xor_4  g10446(.A(new_n10822), .B(new_n10805), .Y(new_n10823));
  xor_4  g10447(.A(new_n10823), .B(new_n10796), .Y(new_n10824));
  xor_4  g10448(.A(new_n10824), .B(new_n10791), .Y(new_n10825));
  not_8  g10449(.A(new_n5127), .Y(new_n10826));
  nand_5 g10450(.A(new_n5150), .B(new_n10826), .Y(new_n10827));
  or_6   g10451(.A(new_n5151), .B(new_n5126), .Y(new_n10828));
  nand_5 g10452(.A(new_n10828), .B(new_n10827), .Y(new_n10829));
  nand_5 g10453(.A(pi128), .B(pi109), .Y(new_n10830));
  xor_4  g10454(.A(new_n10830), .B(new_n10829), .Y(new_n10831));
  nand_5 g10455(.A(pi013), .B(pi002), .Y(new_n10832));
  or_6   g10456(.A(new_n5215), .B(new_n5188), .Y(new_n10833));
  nand_5 g10457(.A(new_n5221), .B(new_n5216), .Y(new_n10834));
  nand_5 g10458(.A(new_n10834), .B(new_n10833), .Y(new_n10835));
  nand_5 g10459(.A(new_n5218), .B(new_n5217), .Y(new_n10836));
  nand_5 g10460(.A(new_n5219), .B(new_n5186), .Y(new_n10837));
  nand_5 g10461(.A(new_n10837), .B(new_n10836), .Y(new_n10838));
  nand_5 g10462(.A(pi230), .B(pi090), .Y(new_n10839));
  nand_5 g10463(.A(pi141), .B(pi050), .Y(new_n10840));
  xor_4  g10464(.A(new_n10840), .B(new_n10839), .Y(new_n10841));
  xor_4  g10465(.A(new_n10841), .B(new_n10838), .Y(new_n10842));
  xor_4  g10466(.A(new_n10842), .B(new_n10835), .Y(new_n10843));
  xor_4  g10467(.A(new_n10843), .B(new_n10832), .Y(new_n10844));
  xor_4  g10468(.A(new_n10844), .B(new_n10831), .Y(new_n10845));
  nand_5 g10469(.A(new_n5332), .B(new_n5251), .Y(new_n10846));
  nand_5 g10470(.A(new_n5348), .B(new_n5333), .Y(new_n10847));
  nand_5 g10471(.A(new_n10847), .B(new_n10846), .Y(new_n10848));
  nand_5 g10472(.A(pi221), .B(pi133), .Y(new_n10849));
  xor_4  g10473(.A(new_n10849), .B(new_n10848), .Y(new_n10850));
  nand_5 g10474(.A(new_n5324), .B(new_n5323), .Y(new_n10851));
  nand_5 g10475(.A(new_n5325), .B(new_n5284), .Y(new_n10852));
  nand_5 g10476(.A(new_n10852), .B(new_n10851), .Y(new_n10853));
  nand_5 g10477(.A(pi204), .B(pi058), .Y(new_n10854));
  nand_5 g10478(.A(new_n5139), .B(new_n5138), .Y(new_n10855));
  nand_5 g10479(.A(new_n5140), .B(new_n5101), .Y(new_n10856));
  nand_5 g10480(.A(new_n10856), .B(new_n10855), .Y(new_n10857));
  nand_5 g10481(.A(new_n5317), .B(new_n5316), .Y(new_n10858));
  nand_5 g10482(.A(new_n5318), .B(new_n5274), .Y(new_n10859));
  nand_5 g10483(.A(new_n10859), .B(new_n10858), .Y(new_n10860));
  nand_5 g10484(.A(pi131), .B(pi010), .Y(new_n10861));
  xor_4  g10485(.A(new_n10861), .B(new_n10860), .Y(new_n10862));
  xor_4  g10486(.A(new_n10862), .B(new_n10857), .Y(new_n10863));
  xor_4  g10487(.A(new_n10863), .B(new_n10854), .Y(new_n10864));
  xor_4  g10488(.A(new_n10864), .B(new_n10853), .Y(new_n10865));
  xor_4  g10489(.A(new_n10865), .B(new_n10850), .Y(new_n10866));
  xor_4  g10490(.A(new_n10866), .B(new_n10845), .Y(new_n10867));
  xor_4  g10491(.A(new_n10867), .B(new_n10825), .Y(new_n10868));
  xor_4  g10492(.A(new_n10868), .B(new_n10773), .Y(po097));
  xnor_4 g10493(.A(new_n1267), .B(new_n1266), .Y(po098));
  xnor_4 g10494(.A(new_n7945), .B(new_n7944), .Y(po099));
  xnor_4 g10495(.A(new_n891), .B(new_n873), .Y(po100));
  xnor_4 g10496(.A(new_n889), .B(new_n888), .Y(po101));
  xnor_4 g10497(.A(new_n1042), .B(new_n1041), .Y(po102));
  xor_4  g10498(.A(new_n3017), .B(new_n3016), .Y(po103));
  xor_4  g10499(.A(new_n2559), .B(new_n2497), .Y(po104));
  xnor_4 g10500(.A(new_n4228), .B(new_n4227), .Y(po105));
  xnor_4 g10501(.A(new_n5962), .B(new_n5961), .Y(po106));
  xor_4  g10502(.A(new_n9344), .B(new_n9343), .Y(po107));
  xor_4  g10503(.A(new_n4217), .B(new_n4193), .Y(po108));
  nand_5 g10504(.A(pi103), .B(pi046), .Y(new_n10881));
  nor_5  g10505(.A(new_n4643), .B(new_n4610), .Y(new_n10882));
  nor_5  g10506(.A(new_n4644), .B(new_n4541), .Y(new_n10883));
  nor_5  g10507(.A(new_n10883), .B(new_n10882), .Y(new_n10884));
  xor_4  g10508(.A(new_n10884), .B(new_n10881), .Y(new_n10885));
  nand_5 g10509(.A(new_n4462), .B(new_n4461), .Y(new_n10886));
  nand_5 g10510(.A(new_n4463), .B(new_n4418), .Y(new_n10887));
  nand_5 g10511(.A(new_n10887), .B(new_n10886), .Y(new_n10888));
  nand_5 g10512(.A(pi175), .B(pi159), .Y(new_n10889));
  nand_5 g10513(.A(new_n4620), .B(new_n4619), .Y(new_n10890));
  nand_5 g10514(.A(new_n4621), .B(new_n4582), .Y(new_n10891));
  nand_5 g10515(.A(new_n10891), .B(new_n10890), .Y(new_n10892));
  xor_4  g10516(.A(new_n10892), .B(new_n10889), .Y(new_n10893));
  nand_5 g10517(.A(new_n4626), .B(new_n4622), .Y(new_n10894));
  nand_5 g10518(.A(new_n4634), .B(new_n4627), .Y(new_n10895));
  nand_5 g10519(.A(new_n10895), .B(new_n10894), .Y(new_n10896));
  nand_5 g10520(.A(pi117), .B(pi068), .Y(new_n10897));
  xor_4  g10521(.A(new_n10897), .B(new_n10896), .Y(new_n10898));
  xor_4  g10522(.A(new_n10898), .B(new_n10893), .Y(new_n10899));
  xor_4  g10523(.A(new_n10899), .B(new_n10888), .Y(new_n10900));
  xor_4  g10524(.A(new_n10900), .B(new_n10885), .Y(new_n10901));
  nand_5 g10525(.A(new_n4642), .B(new_n4637), .Y(new_n10902));
  nand_5 g10526(.A(new_n10902), .B(new_n4638), .Y(new_n10903));
  nand_5 g10527(.A(new_n4526), .B(new_n4525), .Y(new_n10904));
  nand_5 g10528(.A(new_n4527), .B(new_n4348), .Y(new_n10905));
  nand_5 g10529(.A(new_n10905), .B(new_n10904), .Y(new_n10906));
  not_8  g10530(.A(new_n4507), .Y(new_n10907));
  nor_5  g10531(.A(new_n10907), .B(new_n4479), .Y(new_n10908));
  nor_5  g10532(.A(new_n4508), .B(new_n4451), .Y(new_n10909));
  nor_5  g10533(.A(new_n10909), .B(new_n10908), .Y(new_n10910));
  xor_4  g10534(.A(new_n10910), .B(new_n10906), .Y(new_n10911));
  nor_5  g10535(.A(new_n4465), .B(new_n4420), .Y(new_n10912));
  nor_5  g10536(.A(new_n4466), .B(new_n4464), .Y(new_n10913));
  or_6   g10537(.A(new_n10913), .B(new_n10912), .Y(new_n10914));
  nand_5 g10538(.A(pi180), .B(pi080), .Y(new_n10915));
  and_6  g10539(.A(new_n4534), .B(new_n4362), .Y(new_n10916));
  nor_5  g10540(.A(new_n4536), .B(new_n4531), .Y(new_n10917));
  nor_5  g10541(.A(new_n10917), .B(new_n10916), .Y(new_n10918));
  nand_5 g10542(.A(pi200), .B(pi033), .Y(new_n10919));
  xor_4  g10543(.A(new_n10919), .B(new_n10918), .Y(new_n10920));
  xor_4  g10544(.A(new_n10920), .B(new_n10915), .Y(new_n10921));
  and_6  g10545(.A(new_n4502), .B(new_n4390), .Y(new_n10922));
  nor_5  g10546(.A(new_n4504), .B(new_n4500), .Y(new_n10923));
  nor_5  g10547(.A(new_n10923), .B(new_n10922), .Y(new_n10924));
  nand_5 g10548(.A(pi193), .B(pi134), .Y(new_n10925));
  nand_5 g10549(.A(pi181), .B(pi179), .Y(new_n10926));
  xor_4  g10550(.A(new_n10926), .B(new_n10925), .Y(new_n10927));
  nand_5 g10551(.A(pi240), .B(pi238), .Y(new_n10928));
  nand_5 g10552(.A(pi237), .B(pi149), .Y(new_n10929));
  xor_4  g10553(.A(new_n10929), .B(new_n10928), .Y(new_n10930));
  xor_4  g10554(.A(new_n10930), .B(new_n10927), .Y(new_n10931));
  xor_4  g10555(.A(new_n10931), .B(new_n10924), .Y(new_n10932));
  xor_4  g10556(.A(new_n10932), .B(new_n10921), .Y(new_n10933));
  nand_5 g10557(.A(pi247), .B(pi085), .Y(new_n10934));
  nand_5 g10558(.A(pi203), .B(pi162), .Y(new_n10935));
  xor_4  g10559(.A(new_n10935), .B(new_n10934), .Y(new_n10936));
  nand_5 g10560(.A(pi070), .B(pi061), .Y(new_n10937));
  xor_4  g10561(.A(new_n10937), .B(new_n10936), .Y(new_n10938));
  xor_4  g10562(.A(new_n10938), .B(new_n10933), .Y(new_n10939));
  xor_4  g10563(.A(new_n10939), .B(new_n10914), .Y(new_n10940));
  xor_4  g10564(.A(new_n10940), .B(new_n10911), .Y(new_n10941));
  xor_4  g10565(.A(new_n10941), .B(new_n10903), .Y(new_n10942));
  nand_5 g10566(.A(new_n4519), .B(new_n4518), .Y(new_n10943));
  nand_5 g10567(.A(new_n4520), .B(new_n4361), .Y(new_n10944));
  nand_5 g10568(.A(new_n10944), .B(new_n10943), .Y(new_n10945));
  nand_5 g10569(.A(new_n4521), .B(new_n4517), .Y(new_n10946));
  nand_5 g10570(.A(new_n4530), .B(new_n4522), .Y(new_n10947));
  nand_5 g10571(.A(new_n10947), .B(new_n10946), .Y(new_n10948));
  xnor_4 g10572(.A(new_n10948), .B(new_n10945), .Y(new_n10949));
  nand_5 g10573(.A(pi178), .B(pi115), .Y(new_n10950));
  nand_5 g10574(.A(pi202), .B(pi143), .Y(new_n10951));
  xor_4  g10575(.A(new_n10951), .B(new_n10950), .Y(new_n10952));
  xor_4  g10576(.A(new_n10952), .B(new_n10949), .Y(new_n10953));
  xor_4  g10577(.A(new_n10953), .B(new_n10942), .Y(new_n10954));
  xor_4  g10578(.A(new_n10954), .B(new_n10901), .Y(new_n10955));
  nand_5 g10579(.A(pi234), .B(pi194), .Y(new_n10956));
  nand_5 g10580(.A(pi148), .B(pi043), .Y(new_n10957));
  nand_5 g10581(.A(pi228), .B(pi098), .Y(new_n10958));
  xnor_4 g10582(.A(new_n10958), .B(new_n10957), .Y(new_n10959));
  nand_5 g10583(.A(new_n4472), .B(new_n4471), .Y(new_n10960));
  nand_5 g10584(.A(new_n4473), .B(new_n4430), .Y(new_n10961));
  nand_5 g10585(.A(new_n10961), .B(new_n10960), .Y(new_n10962));
  xor_4  g10586(.A(new_n10962), .B(new_n10959), .Y(new_n10963));
  xor_4  g10587(.A(new_n10963), .B(new_n10956), .Y(new_n10964));
  nand_5 g10588(.A(new_n4537), .B(new_n4514), .Y(new_n10965));
  or_6   g10589(.A(new_n4538), .B(new_n4512), .Y(new_n10966));
  nand_5 g10590(.A(new_n10966), .B(new_n10965), .Y(new_n10967));
  xor_4  g10591(.A(new_n10967), .B(new_n10964), .Y(new_n10968));
  nand_5 g10592(.A(new_n4615), .B(new_n4583), .Y(new_n10969));
  not_8  g10593(.A(new_n4618), .Y(new_n10970));
  nand_5 g10594(.A(new_n4635), .B(new_n10970), .Y(new_n10971));
  nand_5 g10595(.A(new_n10971), .B(new_n10969), .Y(new_n10972));
  or_6   g10596(.A(new_n4505), .B(new_n4484), .Y(new_n10973));
  nand_5 g10597(.A(new_n4505), .B(new_n4484), .Y(new_n10974));
  nand_5 g10598(.A(new_n10974), .B(new_n4482), .Y(new_n10975));
  nand_5 g10599(.A(new_n10975), .B(new_n10973), .Y(new_n10976));
  nand_5 g10600(.A(pi116), .B(pi012), .Y(new_n10977));
  xor_4  g10601(.A(new_n10977), .B(new_n10976), .Y(new_n10978));
  xor_4  g10602(.A(new_n10978), .B(new_n10972), .Y(new_n10979));
  nand_5 g10603(.A(pi163), .B(pi126), .Y(new_n10980));
  nand_5 g10604(.A(pi036), .B(pi016), .Y(new_n10981));
  xor_4  g10605(.A(new_n10981), .B(new_n10980), .Y(new_n10982));
  or_6   g10606(.A(new_n4474), .B(new_n4470), .Y(new_n10983));
  nand_5 g10607(.A(new_n4475), .B(new_n4467), .Y(new_n10984));
  nand_5 g10608(.A(new_n10984), .B(new_n10983), .Y(new_n10985));
  xor_4  g10609(.A(new_n10985), .B(new_n10982), .Y(new_n10986));
  xor_4  g10610(.A(new_n10986), .B(new_n10979), .Y(new_n10987));
  xor_4  g10611(.A(new_n10987), .B(new_n10968), .Y(new_n10988));
  nand_5 g10612(.A(new_n4539), .B(new_n4509), .Y(new_n10989));
  nand_5 g10613(.A(new_n4540), .B(new_n4448), .Y(new_n10990));
  nand_5 g10614(.A(new_n10990), .B(new_n10989), .Y(new_n10991));
  nand_5 g10615(.A(pi167), .B(pi048), .Y(new_n10992));
  xor_4  g10616(.A(new_n10992), .B(new_n10991), .Y(new_n10993));
  nand_5 g10617(.A(pi201), .B(pi007), .Y(new_n10994));
  and_6  g10618(.A(new_n4458), .B(new_n4431), .Y(new_n10995));
  nor_5  g10619(.A(new_n4476), .B(new_n4460), .Y(new_n10996));
  nor_5  g10620(.A(new_n10996), .B(new_n10995), .Y(new_n10997));
  xor_4  g10621(.A(new_n10997), .B(new_n10994), .Y(new_n10998));
  not_8  g10622(.A(new_n4494), .Y(new_n10999));
  nor_5  g10623(.A(new_n4498), .B(new_n10999), .Y(new_n11000));
  nor_5  g10624(.A(new_n4499), .B(new_n4491), .Y(new_n11001));
  nor_5  g10625(.A(new_n11001), .B(new_n11000), .Y(new_n11002));
  nand_5 g10626(.A(pi113), .B(pi049), .Y(new_n11003));
  xor_4  g10627(.A(new_n11003), .B(new_n11002), .Y(new_n11004));
  xor_4  g10628(.A(new_n11004), .B(new_n10998), .Y(new_n11005));
  nand_5 g10629(.A(pi083), .B(pi051), .Y(new_n11006));
  nor_5  g10630(.A(new_n4489), .B(new_n4401), .Y(new_n11007));
  nor_5  g10631(.A(new_n4490), .B(new_n4488), .Y(new_n11008));
  nor_5  g10632(.A(new_n11008), .B(new_n11007), .Y(new_n11009));
  xor_4  g10633(.A(new_n11009), .B(new_n11006), .Y(new_n11010));
  nor_5  g10634(.A(new_n4523), .B(new_n4350), .Y(new_n11011));
  nor_5  g10635(.A(new_n4528), .B(new_n4524), .Y(new_n11012));
  nor_5  g10636(.A(new_n11012), .B(new_n11011), .Y(new_n11013));
  xor_4  g10637(.A(new_n11013), .B(new_n11010), .Y(new_n11014));
  or_6   g10638(.A(new_n4628), .B(new_n4596), .Y(new_n11015));
  not_8  g10639(.A(new_n4633), .Y(new_n11016));
  nand_5 g10640(.A(new_n11016), .B(new_n4629), .Y(new_n11017));
  nand_5 g10641(.A(new_n11017), .B(new_n11015), .Y(new_n11018));
  nand_5 g10642(.A(pi214), .B(pi057), .Y(new_n11019));
  nand_5 g10643(.A(new_n4631), .B(new_n4630), .Y(new_n11020));
  nand_5 g10644(.A(new_n4632), .B(new_n4594), .Y(new_n11021));
  nand_5 g10645(.A(new_n11021), .B(new_n11020), .Y(new_n11022));
  xor_4  g10646(.A(new_n11022), .B(new_n11019), .Y(new_n11023));
  nand_5 g10647(.A(pi188), .B(pi000), .Y(new_n11024));
  nand_5 g10648(.A(pi171), .B(pi038), .Y(new_n11025));
  xor_4  g10649(.A(new_n11025), .B(new_n11024), .Y(new_n11026));
  xor_4  g10650(.A(new_n11026), .B(new_n11023), .Y(new_n11027));
  xor_4  g10651(.A(new_n11027), .B(new_n11018), .Y(new_n11028));
  xor_4  g10652(.A(new_n11028), .B(new_n11014), .Y(new_n11029));
  nand_5 g10653(.A(pi144), .B(pi039), .Y(new_n11030));
  nand_5 g10654(.A(pi063), .B(pi042), .Y(new_n11031));
  xor_4  g10655(.A(new_n11031), .B(new_n11030), .Y(new_n11032));
  or_6   g10656(.A(new_n4477), .B(new_n4456), .Y(new_n11033));
  nand_5 g10657(.A(new_n4478), .B(new_n4454), .Y(new_n11034));
  nand_5 g10658(.A(new_n11034), .B(new_n11033), .Y(new_n11035));
  nand_5 g10659(.A(new_n4486), .B(new_n4485), .Y(new_n11036));
  nand_5 g10660(.A(new_n4487), .B(new_n4399), .Y(new_n11037));
  nand_5 g10661(.A(new_n11037), .B(new_n11036), .Y(new_n11038));
  nand_5 g10662(.A(new_n4496), .B(new_n4495), .Y(new_n11039));
  nand_5 g10663(.A(new_n4497), .B(new_n4389), .Y(new_n11040));
  nand_5 g10664(.A(new_n11040), .B(new_n11039), .Y(new_n11041));
  nand_5 g10665(.A(pi245), .B(pi118), .Y(new_n11042));
  nand_5 g10666(.A(pi156), .B(pi108), .Y(new_n11043));
  nand_5 g10667(.A(pi107), .B(pi028), .Y(new_n11044));
  xor_4  g10668(.A(new_n11044), .B(new_n11043), .Y(new_n11045));
  xor_4  g10669(.A(new_n11045), .B(new_n11042), .Y(new_n11046));
  xor_4  g10670(.A(new_n11046), .B(new_n11041), .Y(new_n11047));
  xor_4  g10671(.A(new_n11047), .B(new_n11038), .Y(new_n11048));
  xor_4  g10672(.A(new_n11048), .B(new_n11035), .Y(new_n11049));
  xor_4  g10673(.A(new_n11049), .B(new_n11032), .Y(new_n11050));
  xor_4  g10674(.A(new_n11050), .B(new_n11029), .Y(new_n11051));
  xor_4  g10675(.A(new_n11051), .B(new_n11005), .Y(new_n11052));
  xor_4  g10676(.A(new_n11052), .B(new_n10993), .Y(new_n11053));
  xor_4  g10677(.A(new_n11053), .B(new_n10988), .Y(new_n11054));
  xor_4  g10678(.A(new_n11054), .B(new_n10955), .Y(po109));
  xor_4  g10679(.A(new_n5009), .B(new_n5008), .Y(po110));
  xor_4  g10680(.A(new_n3008), .B(new_n3007), .Y(po111));
  xor_4  g10681(.A(new_n8127), .B(new_n8126), .Y(po112));
  xnor_4 g10682(.A(new_n8187), .B(new_n8133), .Y(po113));
  xnor_4 g10683(.A(new_n8563), .B(new_n8562), .Y(po114));
  xnor_4 g10684(.A(new_n7176), .B(new_n7075), .Y(po115));
  xor_4  g10685(.A(new_n9338), .B(new_n9337), .Y(po116));
  xor_4  g10686(.A(new_n9688), .B(new_n9687), .Y(po117));
  xor_4  g10687(.A(new_n8566), .B(new_n8565), .Y(po118));
  xnor_4 g10688(.A(new_n4608), .B(new_n4607), .Y(po119));
endmodule


