// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Mon Aug 12 17:50:58 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119;
  wire new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n384,
    new_n385, new_n386, new_n387, new_n388, new_n389, new_n390, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1875, new_n1876, new_n1877, new_n1878, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1890, new_n1891, new_n1892,
    new_n1893, new_n1894, new_n1895, new_n1896, new_n1897, new_n1898,
    new_n1899, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019,
    new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025,
    new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031,
    new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055,
    new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061,
    new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067,
    new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896,
    new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914,
    new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944,
    new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956,
    new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962,
    new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046,
    new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052,
    new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058,
    new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064,
    new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070,
    new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076,
    new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088,
    new_n3089, new_n3090, new_n3091, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3101, new_n3102, new_n3103, new_n3104, new_n3105, new_n3106,
    new_n3107, new_n3108, new_n3109, new_n3110, new_n3111, new_n3112,
    new_n3113, new_n3114, new_n3115, new_n3116, new_n3117, new_n3118,
    new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125,
    new_n3126, new_n3127, new_n3128, new_n3129, new_n3130, new_n3131,
    new_n3132, new_n3133, new_n3134, new_n3135, new_n3136, new_n3137,
    new_n3138, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143,
    new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149,
    new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3155,
    new_n3156, new_n3157, new_n3158, new_n3159, new_n3160, new_n3161,
    new_n3162, new_n3163, new_n3164, new_n3165, new_n3166, new_n3167,
    new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173,
    new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179,
    new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185,
    new_n3186, new_n3187, new_n3188, new_n3189, new_n3190, new_n3191,
    new_n3192, new_n3193, new_n3194, new_n3195, new_n3196, new_n3197,
    new_n3198, new_n3199, new_n3200, new_n3201, new_n3202, new_n3203,
    new_n3204, new_n3205, new_n3206, new_n3207, new_n3208, new_n3209,
    new_n3210, new_n3211, new_n3212, new_n3213, new_n3214, new_n3215,
    new_n3216, new_n3217, new_n3218, new_n3219, new_n3220, new_n3221,
    new_n3222, new_n3223, new_n3224, new_n3225, new_n3226, new_n3227,
    new_n3228, new_n3229, new_n3230, new_n3231, new_n3232, new_n3233,
    new_n3234, new_n3235, new_n3236, new_n3237, new_n3238, new_n3239,
    new_n3240, new_n3241, new_n3242, new_n3243, new_n3244, new_n3245,
    new_n3246, new_n3247, new_n3248, new_n3249, new_n3250, new_n3251,
    new_n3252, new_n3253, new_n3254, new_n3255, new_n3256, new_n3257,
    new_n3258, new_n3259, new_n3260, new_n3261, new_n3262, new_n3263,
    new_n3264, new_n3265, new_n3266, new_n3267, new_n3268, new_n3269,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3513, new_n3514, new_n3515, new_n3516, new_n3517,
    new_n3518, new_n3522, new_n3523, new_n3524, new_n3525, new_n3526,
    new_n3527, new_n3528, new_n3529, new_n3530, new_n3531, new_n3532,
    new_n3533, new_n3534, new_n3535, new_n3536, new_n3537, new_n3538,
    new_n3539, new_n3540, new_n3541, new_n3542, new_n3543, new_n3544,
    new_n3545, new_n3546, new_n3547, new_n3548, new_n3549, new_n3550,
    new_n3551, new_n3552, new_n3553, new_n3554, new_n3555, new_n3556,
    new_n3557, new_n3558, new_n3559, new_n3560, new_n3561, new_n3562,
    new_n3563, new_n3564, new_n3565, new_n3566, new_n3567, new_n3568,
    new_n3569, new_n3570, new_n3571, new_n3572, new_n3573, new_n3574,
    new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4214, new_n4215, new_n4216, new_n4217,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226, new_n4227, new_n4228, new_n4229,
    new_n4230, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4812, new_n4813,
    new_n4814, new_n4815, new_n4816, new_n4817, new_n4818, new_n4819,
    new_n4820, new_n4821, new_n4822, new_n4823, new_n4824, new_n4825,
    new_n4826, new_n4827, new_n4828, new_n4829, new_n4830, new_n4831,
    new_n4832, new_n4833, new_n4834, new_n4835, new_n4836, new_n4837,
    new_n4838, new_n4839, new_n4840, new_n4841, new_n4842, new_n4843,
    new_n4844, new_n4845, new_n4846, new_n4847, new_n4848, new_n4849,
    new_n4850, new_n4851, new_n4852, new_n4853, new_n4854, new_n4855,
    new_n4856, new_n4857, new_n4858, new_n4859, new_n4860, new_n4861,
    new_n4862, new_n4863, new_n4864, new_n4865, new_n4866, new_n4867,
    new_n4868, new_n4869, new_n4870, new_n4871, new_n4872, new_n4873,
    new_n4874, new_n4875, new_n4876, new_n4877, new_n4878, new_n4879,
    new_n4880, new_n4881, new_n4882, new_n4883, new_n4884, new_n4885,
    new_n4886, new_n4887, new_n4888, new_n4889, new_n4890, new_n4891,
    new_n4892, new_n4893, new_n4894, new_n4895, new_n4896, new_n4897,
    new_n4898, new_n4899, new_n4900, new_n4901, new_n4902, new_n4903,
    new_n4904, new_n4905, new_n4906, new_n4907, new_n4908, new_n4909,
    new_n4910, new_n4911, new_n4912, new_n4913, new_n4914, new_n4915,
    new_n4916, new_n4917, new_n4918, new_n4919, new_n4920, new_n4921,
    new_n4922, new_n4923, new_n4924, new_n4925, new_n4926, new_n4927,
    new_n4928, new_n4929, new_n4930, new_n4931, new_n4932, new_n4933,
    new_n4934, new_n4935, new_n4936, new_n4937, new_n4938, new_n4939,
    new_n4940, new_n4941, new_n4942, new_n4943, new_n4944, new_n4945,
    new_n4946, new_n4947, new_n4948, new_n4949, new_n4950, new_n4951,
    new_n4952, new_n4953, new_n4954, new_n4955, new_n4956, new_n4957,
    new_n4958, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970,
    new_n4971, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020,
    new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026,
    new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6377, new_n6378, new_n6379,
    new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385,
    new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391,
    new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397,
    new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429, new_n6430, new_n6431, new_n6432, new_n6433,
    new_n6434, new_n6435, new_n6436, new_n6437, new_n6438, new_n6439,
    new_n6440, new_n6441, new_n6442, new_n6443, new_n6444, new_n6445,
    new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451,
    new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457,
    new_n6458, new_n6459, new_n6460, new_n6461, new_n6462, new_n6463,
    new_n6464, new_n6465, new_n6466, new_n6467, new_n6468, new_n6469,
    new_n6470, new_n6471, new_n6472, new_n6473, new_n6474, new_n6475,
    new_n6476, new_n6477, new_n6478, new_n6479, new_n6480, new_n6481,
    new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487,
    new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493,
    new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558,
    new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6567, new_n6568, new_n6569, new_n6570,
    new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576,
    new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582,
    new_n6583, new_n6584, new_n6585, new_n6586, new_n6587, new_n6588,
    new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611, new_n6612,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687,
    new_n6688, new_n6689, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254,
    new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278,
    new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7917, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922,
    new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959, new_n7960, new_n7961, new_n7962, new_n7963, new_n7964,
    new_n7965, new_n7966, new_n7967, new_n7968, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637, new_n8638, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663,
    new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9652, new_n9653, new_n9654, new_n9655,
    new_n9656, new_n9657, new_n9658, new_n9659, new_n9660, new_n9661,
    new_n9662, new_n9663, new_n9664, new_n9665, new_n9666, new_n9667,
    new_n9668, new_n9669, new_n9670, new_n9671, new_n9672, new_n9673,
    new_n9674, new_n9675, new_n9676, new_n9677, new_n9678, new_n9679,
    new_n9680, new_n9681, new_n9682, new_n9683, new_n9684, new_n9685,
    new_n9686, new_n9687, new_n9688, new_n9689, new_n9690, new_n9691,
    new_n9692, new_n9693, new_n9694, new_n9695, new_n9696, new_n9697,
    new_n9698, new_n9699, new_n9700, new_n9701, new_n9702, new_n9703,
    new_n9704, new_n9705, new_n9706, new_n9707, new_n9708, new_n9709,
    new_n9710, new_n9711, new_n9712, new_n9713, new_n9714, new_n9715,
    new_n9716, new_n9717, new_n9718, new_n9719, new_n9720, new_n9721,
    new_n9722, new_n9723, new_n9724, new_n9725, new_n9726, new_n9727,
    new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733,
    new_n9734, new_n9735, new_n9736, new_n9737, new_n9738, new_n9739,
    new_n9740, new_n9741, new_n9742, new_n9743, new_n9744, new_n9745,
    new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751,
    new_n9752, new_n9753, new_n9754, new_n9755, new_n9756, new_n9757,
    new_n9758, new_n9759, new_n9760, new_n9761, new_n9762, new_n9763,
    new_n9764, new_n9765, new_n9766, new_n9767, new_n9768, new_n9769,
    new_n9770, new_n9771, new_n9772, new_n9773, new_n9774, new_n9775,
    new_n9776, new_n9777, new_n9778, new_n9779, new_n9780, new_n9781,
    new_n9782, new_n9783, new_n9784, new_n9785, new_n9786, new_n9787,
    new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793,
    new_n9794, new_n9795, new_n9796, new_n9797, new_n9798, new_n9799,
    new_n9800, new_n9801, new_n9802, new_n9803, new_n9804, new_n9805,
    new_n9806, new_n9807, new_n9808, new_n9809, new_n9810, new_n9811,
    new_n9812, new_n9813, new_n9814, new_n9815, new_n9816, new_n9817,
    new_n9818, new_n9819, new_n9820, new_n9829, new_n9830, new_n9831,
    new_n9832, new_n9833, new_n9834, new_n9835, new_n9836, new_n9837,
    new_n9838, new_n9839, new_n9840, new_n9841, new_n9842, new_n9843,
    new_n9844, new_n9845, new_n9846, new_n9847, new_n9848, new_n9849,
    new_n9850, new_n9851, new_n9852, new_n9853, new_n9854, new_n9855,
    new_n9856, new_n9857, new_n9858, new_n9859, new_n9860, new_n9861,
    new_n9862, new_n9863, new_n9864, new_n9865, new_n9866, new_n9867,
    new_n9868, new_n9869, new_n9870, new_n9871, new_n9872, new_n9873,
    new_n9874, new_n9875, new_n9876, new_n9877, new_n9878, new_n9879,
    new_n9880, new_n9881, new_n9882, new_n9883, new_n9884, new_n9885,
    new_n9886, new_n9887, new_n9888, new_n9889, new_n9890, new_n9891,
    new_n9892, new_n9893, new_n9894, new_n9895, new_n9896, new_n9897,
    new_n9898, new_n9899, new_n9900, new_n9901, new_n9902, new_n9903,
    new_n9904, new_n9905, new_n9906, new_n9907, new_n9908, new_n9909,
    new_n9910, new_n9911, new_n9912, new_n9913, new_n9914, new_n9915,
    new_n9916, new_n9917, new_n9918, new_n9919, new_n9920, new_n9921,
    new_n9922, new_n9923, new_n9924, new_n9925, new_n9926, new_n9927,
    new_n9928, new_n9929, new_n9930, new_n9931, new_n9932, new_n9933,
    new_n9934, new_n9935, new_n9936, new_n9937, new_n9938, new_n9939,
    new_n9940, new_n9941, new_n9942, new_n9943, new_n9944, new_n9945,
    new_n9946, new_n9947, new_n9948, new_n9949, new_n9950, new_n9951,
    new_n9952, new_n9953, new_n9954, new_n9955, new_n9956, new_n9957,
    new_n9958, new_n9959, new_n9960, new_n9961, new_n9962, new_n9963,
    new_n9964, new_n9965, new_n9966, new_n9967, new_n9968, new_n9969,
    new_n9970, new_n9971, new_n9972, new_n9973, new_n9974, new_n9975,
    new_n9976, new_n9977, new_n9978, new_n9979, new_n9980, new_n9981,
    new_n9982, new_n9983, new_n9984, new_n9985, new_n9986, new_n9987,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009, new_n10010, new_n10011,
    new_n10012, new_n10013, new_n10014, new_n10015, new_n10016, new_n10017,
    new_n10018, new_n10019, new_n10020, new_n10021, new_n10022, new_n10023,
    new_n10024, new_n10025, new_n10026, new_n10027, new_n10028, new_n10029,
    new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035,
    new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041,
    new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047,
    new_n10048, new_n10049, new_n10050, new_n10051, new_n10052, new_n10053,
    new_n10054, new_n10055, new_n10056, new_n10057, new_n10058, new_n10059,
    new_n10060, new_n10061, new_n10062, new_n10063, new_n10064, new_n10065,
    new_n10066, new_n10067, new_n10068, new_n10069, new_n10070, new_n10071,
    new_n10072, new_n10073, new_n10074, new_n10075, new_n10076, new_n10077,
    new_n10078, new_n10079, new_n10080, new_n10081, new_n10082, new_n10083,
    new_n10084, new_n10085, new_n10086, new_n10087, new_n10088, new_n10089,
    new_n10090, new_n10091, new_n10092, new_n10093, new_n10094, new_n10095,
    new_n10096, new_n10097, new_n10098, new_n10099, new_n10100, new_n10101,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111, new_n10112, new_n10113,
    new_n10114, new_n10115, new_n10116, new_n10117, new_n10118, new_n10119,
    new_n10120, new_n10121, new_n10122, new_n10123, new_n10124, new_n10125,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158, new_n10159, new_n10160, new_n10161,
    new_n10162, new_n10163, new_n10164, new_n10165, new_n10166, new_n10167,
    new_n10168, new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174, new_n10175, new_n10176, new_n10177, new_n10178, new_n10179,
    new_n10180, new_n10181, new_n10182, new_n10183, new_n10184, new_n10185,
    new_n10186, new_n10187, new_n10188, new_n10189, new_n10190, new_n10191,
    new_n10192, new_n10193, new_n10194, new_n10195, new_n10196, new_n10197,
    new_n10198, new_n10199, new_n10200, new_n10201, new_n10202, new_n10203,
    new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209,
    new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215,
    new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236, new_n10237, new_n10238, new_n10239,
    new_n10240, new_n10241, new_n10242, new_n10243, new_n10244, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250, new_n10251,
    new_n10252, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10263,
    new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274, new_n10275,
    new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283, new_n10284, new_n10285, new_n10286, new_n10287,
    new_n10288, new_n10289, new_n10290, new_n10291, new_n10292, new_n10293,
    new_n10294, new_n10295, new_n10296, new_n10297, new_n10298, new_n10299,
    new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305,
    new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311,
    new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317,
    new_n10318, new_n10319, new_n10320, new_n10323, new_n10324, new_n10325,
    new_n10326, new_n10327, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361,
    new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367,
    new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385,
    new_n10386, new_n10387, new_n10388, new_n10389, new_n10390, new_n10391,
    new_n10392, new_n10393, new_n10394, new_n10395, new_n10396, new_n10397,
    new_n10398, new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404, new_n10405, new_n10406, new_n10407, new_n10408, new_n10409,
    new_n10410, new_n10411, new_n10412, new_n10413, new_n10414, new_n10415,
    new_n10416, new_n10417, new_n10418, new_n10419, new_n10420, new_n10421,
    new_n10422, new_n10423, new_n10424, new_n10425, new_n10426, new_n10427,
    new_n10428, new_n10429, new_n10430, new_n10431, new_n10432, new_n10433,
    new_n10434, new_n10435, new_n10436, new_n10437, new_n10438, new_n10439,
    new_n10440, new_n10441, new_n10442, new_n10443, new_n10444, new_n10445,
    new_n10446, new_n10447, new_n10448, new_n10449, new_n10450, new_n10451,
    new_n10452, new_n10453, new_n10454, new_n10455, new_n10456, new_n10457,
    new_n10458, new_n10459, new_n10460, new_n10461, new_n10462, new_n10463,
    new_n10464, new_n10465, new_n10466, new_n10467, new_n10468, new_n10469,
    new_n10470, new_n10471, new_n10472, new_n10473, new_n10474, new_n10475,
    new_n10476, new_n10477, new_n10478, new_n10479, new_n10480, new_n10481,
    new_n10482, new_n10483, new_n10484, new_n10485, new_n10486, new_n10487,
    new_n10488, new_n10489, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10505, new_n10506, new_n10507, new_n10508, new_n10509, new_n10510,
    new_n10511, new_n10512, new_n10513, new_n10514, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525, new_n10526, new_n10527, new_n10528,
    new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534,
    new_n10535, new_n10536, new_n10537, new_n10538, new_n10539, new_n10540,
    new_n10541, new_n10542, new_n10543, new_n10544, new_n10545, new_n10546,
    new_n10547, new_n10548, new_n10549, new_n10550, new_n10551, new_n10552,
    new_n10553, new_n10554, new_n10555, new_n10556, new_n10557, new_n10558,
    new_n10559, new_n10560, new_n10561, new_n10562, new_n10563, new_n10564,
    new_n10565, new_n10566, new_n10567, new_n10568, new_n10569, new_n10570,
    new_n10571, new_n10572, new_n10573, new_n10574, new_n10575, new_n10576,
    new_n10577, new_n10578, new_n10579, new_n10580, new_n10581, new_n10582,
    new_n10583, new_n10584, new_n10585, new_n10586, new_n10587, new_n10588,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593, new_n10594,
    new_n10595, new_n10596, new_n10597, new_n10598, new_n10599, new_n10600,
    new_n10601, new_n10602, new_n10603, new_n10604, new_n10605, new_n10606,
    new_n10607, new_n10608, new_n10609, new_n10610, new_n10611, new_n10612,
    new_n10613, new_n10614, new_n10615, new_n10616, new_n10617, new_n10618,
    new_n10619, new_n10620, new_n10621, new_n10622, new_n10623, new_n10624,
    new_n10625, new_n10626, new_n10627, new_n10628, new_n10629, new_n10630,
    new_n10631, new_n10632, new_n10633, new_n10634, new_n10635, new_n10636,
    new_n10637, new_n10638, new_n10639, new_n10640, new_n10641, new_n10642,
    new_n10643, new_n10644, new_n10645, new_n10646, new_n10647, new_n10648,
    new_n10649, new_n10650, new_n10651, new_n10652, new_n10653, new_n10654,
    new_n10655, new_n10656, new_n10657, new_n10658, new_n10659, new_n10660,
    new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666,
    new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10675, new_n10676, new_n10677, new_n10678,
    new_n10679, new_n10680, new_n10681, new_n10682, new_n10683, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874;
  nand_5 g00000(.A(pi236), .B(pi027), .Y(new_n377));
  nand_5 g00001(.A(pi213), .B(pi164), .Y(new_n378));
  xor_4  g00002(.A(new_n378), .B(new_n377), .Y(new_n379));
  nand_5 g00003(.A(pi168), .B(pi147), .Y(new_n380));
  xor_4  g00004(.A(new_n380), .B(new_n379), .Y(new_n381));
  nand_5 g00005(.A(pi131), .B(pi119), .Y(new_n382));
  xor_4  g00006(.A(new_n382), .B(new_n381), .Y(po000));
  nand_5 g00007(.A(pi245), .B(pi008), .Y(new_n384));
  nand_5 g00008(.A(pi156), .B(pi027), .Y(new_n385));
  nand_5 g00009(.A(pi201), .B(pi026), .Y(new_n386));
  nand_5 g00010(.A(new_n386), .B(new_n385), .Y(new_n387));
  nand_5 g00011(.A(pi201), .B(pi027), .Y(new_n388));
  nand_5 g00012(.A(pi156), .B(pi026), .Y(new_n389));
  or_6   g00013(.A(new_n389), .B(new_n388), .Y(new_n390));
  nand_5 g00014(.A(new_n390), .B(new_n387), .Y(new_n391));
  xor_4  g00015(.A(new_n391), .B(new_n384), .Y(new_n392));
  nand_5 g00016(.A(pi245), .B(pi026), .Y(new_n393));
  nand_5 g00017(.A(pi049), .B(pi008), .Y(new_n394));
  nand_5 g00018(.A(new_n394), .B(new_n393), .Y(new_n395));
  xor_4  g00019(.A(new_n394), .B(new_n393), .Y(new_n396));
  nand_5 g00020(.A(new_n396), .B(new_n388), .Y(new_n397));
  nand_5 g00021(.A(new_n397), .B(new_n395), .Y(new_n398));
  xor_4  g00022(.A(new_n398), .B(new_n392), .Y(new_n399));
  nand_5 g00023(.A(pi171), .B(pi056), .Y(new_n400));
  nand_5 g00024(.A(pi049), .B(pi026), .Y(new_n401));
  nand_5 g00025(.A(pi171), .B(pi008), .Y(new_n402));
  nand_5 g00026(.A(new_n402), .B(new_n401), .Y(new_n403));
  nand_5 g00027(.A(pi245), .B(pi027), .Y(new_n404));
  xor_4  g00028(.A(new_n402), .B(new_n401), .Y(new_n405));
  nand_5 g00029(.A(new_n405), .B(new_n404), .Y(new_n406));
  nand_5 g00030(.A(new_n406), .B(new_n403), .Y(new_n407));
  nand_5 g00031(.A(new_n407), .B(new_n400), .Y(new_n408));
  xor_4  g00032(.A(new_n396), .B(new_n388), .Y(new_n409));
  xor_4  g00033(.A(new_n407), .B(new_n400), .Y(new_n410));
  nand_5 g00034(.A(new_n410), .B(new_n409), .Y(new_n411));
  nand_5 g00035(.A(new_n411), .B(new_n408), .Y(new_n412));
  nand_5 g00036(.A(pi056), .B(pi049), .Y(new_n413));
  nand_5 g00037(.A(pi171), .B(pi136), .Y(new_n414));
  nand_5 g00038(.A(new_n414), .B(new_n413), .Y(new_n415));
  nand_5 g00039(.A(pi136), .B(pi049), .Y(new_n416));
  or_6   g00040(.A(new_n416), .B(new_n400), .Y(new_n417));
  nand_5 g00041(.A(new_n417), .B(new_n415), .Y(new_n418));
  xor_4  g00042(.A(new_n418), .B(new_n412), .Y(new_n419));
  xor_4  g00043(.A(new_n419), .B(new_n399), .Y(new_n420));
  not_8  g00044(.A(new_n420), .Y(new_n421));
  nand_5 g00045(.A(pi136), .B(pi107), .Y(new_n422));
  not_8  g00046(.A(new_n422), .Y(new_n423));
  nand_5 g00047(.A(pi049), .B(pi027), .Y(new_n424));
  nand_5 g00048(.A(pi107), .B(pi008), .Y(new_n425));
  nand_5 g00049(.A(new_n425), .B(new_n424), .Y(new_n426));
  nand_5 g00050(.A(pi171), .B(pi026), .Y(new_n427));
  or_6   g00051(.A(new_n425), .B(new_n424), .Y(new_n428));
  nand_5 g00052(.A(new_n428), .B(new_n427), .Y(new_n429));
  nand_5 g00053(.A(new_n429), .B(new_n426), .Y(new_n430));
  nand_5 g00054(.A(pi107), .B(pi056), .Y(new_n431));
  or_6   g00055(.A(new_n431), .B(new_n430), .Y(new_n432));
  xnor_4 g00056(.A(new_n405), .B(new_n404), .Y(new_n433));
  xor_4  g00057(.A(new_n431), .B(new_n430), .Y(new_n434));
  nand_5 g00058(.A(new_n434), .B(new_n433), .Y(new_n435));
  nand_5 g00059(.A(new_n435), .B(new_n432), .Y(new_n436));
  nand_5 g00060(.A(new_n436), .B(new_n423), .Y(new_n437));
  xor_4  g00061(.A(new_n410), .B(new_n409), .Y(new_n438));
  xor_4  g00062(.A(new_n436), .B(new_n422), .Y(new_n439));
  or_6   g00063(.A(new_n439), .B(new_n438), .Y(new_n440));
  nand_5 g00064(.A(new_n440), .B(new_n437), .Y(new_n441));
  nand_5 g00065(.A(new_n441), .B(new_n421), .Y(new_n442));
  nand_5 g00066(.A(pi201), .B(pi008), .Y(new_n443));
  nand_5 g00067(.A(pi063), .B(pi027), .Y(new_n444));
  xor_4  g00068(.A(new_n444), .B(new_n443), .Y(new_n445));
  xor_4  g00069(.A(new_n445), .B(new_n389), .Y(new_n446));
  not_8  g00070(.A(new_n446), .Y(new_n447));
  nand_5 g00071(.A(pi245), .B(pi056), .Y(new_n448));
  xor_4  g00072(.A(new_n448), .B(new_n390), .Y(new_n449));
  xor_4  g00073(.A(new_n449), .B(new_n447), .Y(new_n450));
  nand_5 g00074(.A(pi171), .B(pi096), .Y(new_n451));
  nand_5 g00075(.A(pi235), .B(pi107), .Y(new_n452));
  xor_4  g00076(.A(new_n452), .B(new_n451), .Y(new_n453));
  xor_4  g00077(.A(new_n453), .B(new_n416), .Y(new_n454));
  nand_5 g00078(.A(new_n391), .B(new_n384), .Y(new_n455));
  nand_5 g00079(.A(new_n398), .B(new_n392), .Y(new_n456));
  nand_5 g00080(.A(new_n456), .B(new_n455), .Y(new_n457));
  xor_4  g00081(.A(new_n457), .B(new_n454), .Y(new_n458));
  xor_4  g00082(.A(new_n458), .B(new_n450), .Y(new_n459));
  nand_5 g00083(.A(new_n418), .B(new_n412), .Y(new_n460));
  nand_5 g00084(.A(new_n419), .B(new_n399), .Y(new_n461));
  nand_5 g00085(.A(new_n461), .B(new_n460), .Y(new_n462));
  xor_4  g00086(.A(new_n462), .B(new_n417), .Y(new_n463));
  xnor_4 g00087(.A(new_n463), .B(new_n459), .Y(new_n464));
  xnor_4 g00088(.A(new_n464), .B(new_n442), .Y(new_n465));
  nand_5 g00089(.A(pi107), .B(pi096), .Y(new_n466));
  xnor_4 g00090(.A(new_n434), .B(new_n433), .Y(new_n467));
  not_8  g00091(.A(new_n427), .Y(new_n468));
  not_8  g00092(.A(new_n426), .Y(new_n469));
  nand_5 g00093(.A(pi107), .B(pi027), .Y(new_n470));
  nand_5 g00094(.A(new_n470), .B(new_n468), .Y(new_n471));
  nand_5 g00095(.A(new_n471), .B(new_n469), .Y(new_n472));
  nand_5 g00096(.A(new_n472), .B(new_n428), .Y(new_n473));
  nand_5 g00097(.A(new_n473), .B(new_n468), .Y(new_n474));
  nor_5  g00098(.A(new_n474), .B(new_n467), .Y(new_n475));
  xor_4  g00099(.A(new_n439), .B(new_n438), .Y(new_n476));
  nand_5 g00100(.A(new_n476), .B(new_n475), .Y(new_n477));
  nand_5 g00101(.A(new_n477), .B(new_n466), .Y(new_n478));
  xor_4  g00102(.A(new_n441), .B(new_n420), .Y(new_n479));
  xor_4  g00103(.A(new_n477), .B(new_n466), .Y(new_n480));
  nand_5 g00104(.A(new_n480), .B(new_n479), .Y(new_n481));
  nand_5 g00105(.A(new_n481), .B(new_n478), .Y(new_n482));
  xor_4  g00106(.A(new_n482), .B(new_n465), .Y(new_n483));
  nand_5 g00107(.A(pi039), .B(pi032), .Y(new_n484));
  nand_5 g00108(.A(pi206), .B(pi116), .Y(new_n485));
  nand_5 g00109(.A(pi164), .B(pi070), .Y(new_n486));
  nand_5 g00110(.A(new_n486), .B(new_n485), .Y(new_n487));
  nand_5 g00111(.A(pi164), .B(pi116), .Y(new_n488));
  nand_5 g00112(.A(pi206), .B(pi070), .Y(new_n489));
  or_6   g00113(.A(new_n489), .B(new_n488), .Y(new_n490));
  nand_5 g00114(.A(new_n490), .B(new_n487), .Y(new_n491));
  xor_4  g00115(.A(new_n491), .B(new_n484), .Y(new_n492));
  nand_5 g00116(.A(pi228), .B(pi032), .Y(new_n493));
  nand_5 g00117(.A(pi206), .B(pi039), .Y(new_n494));
  nand_5 g00118(.A(new_n494), .B(new_n493), .Y(new_n495));
  xor_4  g00119(.A(new_n494), .B(new_n493), .Y(new_n496));
  nand_5 g00120(.A(new_n496), .B(new_n488), .Y(new_n497));
  nand_5 g00121(.A(new_n497), .B(new_n495), .Y(new_n498));
  xor_4  g00122(.A(new_n498), .B(new_n492), .Y(new_n499));
  nand_5 g00123(.A(pi228), .B(pi145), .Y(new_n500));
  nand_5 g00124(.A(pi246), .B(pi148), .Y(new_n501));
  and_6  g00125(.A(new_n501), .B(new_n500), .Y(new_n502));
  nand_5 g00126(.A(pi148), .B(pi145), .Y(new_n503));
  nand_5 g00127(.A(pi246), .B(pi228), .Y(new_n504));
  nor_5  g00128(.A(new_n504), .B(new_n503), .Y(new_n505));
  or_6   g00129(.A(new_n505), .B(new_n502), .Y(new_n506));
  xnor_4 g00130(.A(new_n506), .B(new_n499), .Y(new_n507));
  nand_5 g00131(.A(pi148), .B(pi032), .Y(new_n508));
  nand_5 g00132(.A(pi164), .B(pi039), .Y(new_n509));
  nand_5 g00133(.A(new_n509), .B(new_n508), .Y(new_n510));
  nand_5 g00134(.A(pi228), .B(pi206), .Y(new_n511));
  xor_4  g00135(.A(new_n509), .B(new_n508), .Y(new_n512));
  nand_5 g00136(.A(new_n512), .B(new_n511), .Y(new_n513));
  nand_5 g00137(.A(new_n513), .B(new_n510), .Y(new_n514));
  nand_5 g00138(.A(new_n514), .B(new_n503), .Y(new_n515));
  xor_4  g00139(.A(new_n496), .B(new_n488), .Y(new_n516));
  xor_4  g00140(.A(new_n514), .B(new_n503), .Y(new_n517));
  nand_5 g00141(.A(new_n517), .B(new_n516), .Y(new_n518));
  nand_5 g00142(.A(new_n518), .B(new_n515), .Y(new_n519));
  xor_4  g00143(.A(new_n519), .B(new_n507), .Y(new_n520));
  nand_5 g00144(.A(pi246), .B(pi163), .Y(new_n521));
  nand_5 g00145(.A(pi163), .B(pi145), .Y(new_n522));
  nand_5 g00146(.A(pi206), .B(pi148), .Y(new_n523));
  nand_5 g00147(.A(pi163), .B(pi032), .Y(new_n524));
  nand_5 g00148(.A(new_n524), .B(new_n523), .Y(new_n525));
  nand_5 g00149(.A(pi228), .B(pi164), .Y(new_n526));
  xor_4  g00150(.A(new_n524), .B(new_n523), .Y(new_n527));
  nand_5 g00151(.A(new_n527), .B(new_n526), .Y(new_n528));
  nand_5 g00152(.A(new_n528), .B(new_n525), .Y(new_n529));
  nand_5 g00153(.A(new_n529), .B(new_n522), .Y(new_n530));
  xor_4  g00154(.A(new_n512), .B(new_n511), .Y(new_n531));
  xor_4  g00155(.A(new_n529), .B(new_n522), .Y(new_n532));
  nand_5 g00156(.A(new_n532), .B(new_n531), .Y(new_n533));
  nand_5 g00157(.A(new_n533), .B(new_n530), .Y(new_n534));
  or_6   g00158(.A(new_n534), .B(new_n521), .Y(new_n535));
  xnor_4 g00159(.A(new_n517), .B(new_n516), .Y(new_n536));
  xor_4  g00160(.A(new_n534), .B(new_n521), .Y(new_n537));
  nand_5 g00161(.A(new_n537), .B(new_n536), .Y(new_n538));
  nand_5 g00162(.A(new_n538), .B(new_n535), .Y(new_n539));
  nand_5 g00163(.A(new_n539), .B(new_n520), .Y(new_n540));
  nand_5 g00164(.A(pi164), .B(pi115), .Y(new_n541));
  nand_5 g00165(.A(pi116), .B(pi032), .Y(new_n542));
  xor_4  g00166(.A(new_n542), .B(new_n541), .Y(new_n543));
  xor_4  g00167(.A(new_n543), .B(new_n489), .Y(new_n544));
  nand_5 g00168(.A(pi145), .B(pi039), .Y(new_n545));
  xor_4  g00169(.A(new_n545), .B(new_n490), .Y(new_n546));
  xor_4  g00170(.A(new_n546), .B(new_n544), .Y(new_n547));
  nand_5 g00171(.A(pi148), .B(pi114), .Y(new_n548));
  nand_5 g00172(.A(pi163), .B(pi091), .Y(new_n549));
  xor_4  g00173(.A(new_n549), .B(new_n548), .Y(new_n550));
  xor_4  g00174(.A(new_n550), .B(new_n504), .Y(new_n551));
  nand_5 g00175(.A(new_n491), .B(new_n484), .Y(new_n552));
  nand_5 g00176(.A(new_n498), .B(new_n492), .Y(new_n553));
  nand_5 g00177(.A(new_n553), .B(new_n552), .Y(new_n554));
  xor_4  g00178(.A(new_n554), .B(new_n551), .Y(new_n555));
  xnor_4 g00179(.A(new_n555), .B(new_n547), .Y(new_n556));
  nor_5  g00180(.A(new_n506), .B(new_n499), .Y(new_n557));
  nor_5  g00181(.A(new_n519), .B(new_n507), .Y(new_n558));
  xor_4  g00182(.A(new_n558), .B(new_n505), .Y(new_n559));
  nor_5  g00183(.A(new_n559), .B(new_n557), .Y(new_n560));
  not_8  g00184(.A(new_n560), .Y(new_n561));
  xor_4  g00185(.A(new_n561), .B(new_n556), .Y(new_n562));
  xor_4  g00186(.A(new_n562), .B(new_n540), .Y(new_n563));
  nand_5 g00187(.A(pi163), .B(pi114), .Y(new_n564));
  xor_4  g00188(.A(new_n527), .B(new_n526), .Y(new_n565));
  nand_5 g00189(.A(pi164), .B(pi163), .Y(new_n566));
  nor_5  g00190(.A(new_n566), .B(new_n523), .Y(new_n567));
  not_8  g00191(.A(new_n567), .Y(new_n568));
  nor_5  g00192(.A(new_n568), .B(new_n565), .Y(new_n569));
  not_8  g00193(.A(new_n569), .Y(new_n570));
  xor_4  g00194(.A(new_n532), .B(new_n531), .Y(new_n571));
  nor_5  g00195(.A(new_n571), .B(new_n570), .Y(new_n572));
  xor_4  g00196(.A(new_n537), .B(new_n536), .Y(new_n573));
  nand_5 g00197(.A(new_n573), .B(new_n572), .Y(new_n574));
  nand_5 g00198(.A(new_n574), .B(new_n564), .Y(new_n575));
  xnor_4 g00199(.A(new_n539), .B(new_n520), .Y(new_n576));
  xor_4  g00200(.A(new_n574), .B(new_n564), .Y(new_n577));
  nand_5 g00201(.A(new_n577), .B(new_n576), .Y(new_n578));
  nand_5 g00202(.A(new_n578), .B(new_n575), .Y(new_n579));
  xor_4  g00203(.A(new_n579), .B(new_n563), .Y(new_n580));
  xor_4  g00204(.A(new_n580), .B(new_n483), .Y(new_n581));
  xor_4  g00205(.A(new_n480), .B(new_n479), .Y(new_n582));
  xor_4  g00206(.A(new_n577), .B(new_n576), .Y(new_n583));
  nor_5  g00207(.A(new_n583), .B(new_n582), .Y(new_n584));
  xnor_4 g00208(.A(new_n583), .B(new_n582), .Y(new_n585));
  xnor_4 g00209(.A(new_n476), .B(new_n475), .Y(new_n586));
  xnor_4 g00210(.A(new_n474), .B(new_n467), .Y(new_n587));
  nand_5 g00211(.A(pi107), .B(pi026), .Y(new_n588));
  nand_5 g00212(.A(pi171), .B(pi027), .Y(new_n589));
  xor_4  g00213(.A(new_n589), .B(new_n588), .Y(new_n590));
  not_8  g00214(.A(new_n590), .Y(new_n591));
  nand_5 g00215(.A(pi164), .B(pi148), .Y(new_n592));
  nand_5 g00216(.A(pi206), .B(pi163), .Y(new_n593));
  nand_5 g00217(.A(new_n593), .B(new_n592), .Y(new_n594));
  nand_5 g00218(.A(new_n594), .B(new_n568), .Y(new_n595));
  nand_5 g00219(.A(new_n595), .B(new_n591), .Y(new_n596));
  nor_5  g00220(.A(new_n566), .B(new_n470), .Y(new_n597));
  xor_4  g00221(.A(new_n595), .B(new_n590), .Y(new_n598));
  or_6   g00222(.A(new_n598), .B(new_n597), .Y(new_n599));
  nand_5 g00223(.A(new_n599), .B(new_n596), .Y(new_n600));
  nor_5  g00224(.A(new_n471), .B(new_n469), .Y(new_n601));
  nor_5  g00225(.A(new_n601), .B(new_n473), .Y(new_n602));
  not_8  g00226(.A(new_n602), .Y(new_n603));
  nand_5 g00227(.A(new_n603), .B(new_n600), .Y(new_n604));
  xor_4  g00228(.A(new_n567), .B(new_n565), .Y(new_n605));
  xor_4  g00229(.A(new_n603), .B(new_n600), .Y(new_n606));
  nand_5 g00230(.A(new_n606), .B(new_n605), .Y(new_n607));
  nand_5 g00231(.A(new_n607), .B(new_n604), .Y(new_n608));
  nand_5 g00232(.A(new_n608), .B(new_n587), .Y(new_n609));
  xor_4  g00233(.A(new_n571), .B(new_n569), .Y(new_n610));
  xor_4  g00234(.A(new_n608), .B(new_n587), .Y(new_n611));
  nand_5 g00235(.A(new_n611), .B(new_n610), .Y(new_n612));
  nand_5 g00236(.A(new_n612), .B(new_n609), .Y(new_n613));
  nand_5 g00237(.A(new_n613), .B(new_n586), .Y(new_n614));
  xor_4  g00238(.A(new_n573), .B(new_n572), .Y(new_n615));
  not_8  g00239(.A(new_n615), .Y(new_n616));
  xor_4  g00240(.A(new_n613), .B(new_n586), .Y(new_n617));
  nand_5 g00241(.A(new_n617), .B(new_n616), .Y(new_n618));
  nand_5 g00242(.A(new_n618), .B(new_n614), .Y(new_n619));
  nor_5  g00243(.A(new_n619), .B(new_n585), .Y(new_n620));
  nor_5  g00244(.A(new_n620), .B(new_n584), .Y(new_n621));
  xor_4  g00245(.A(new_n621), .B(new_n581), .Y(new_n622));
  nand_5 g00246(.A(pi149), .B(pi019), .Y(new_n623));
  nand_5 g00247(.A(pi167), .B(pi151), .Y(new_n624));
  nand_5 g00248(.A(pi181), .B(pi147), .Y(new_n625));
  nand_5 g00249(.A(new_n625), .B(new_n624), .Y(new_n626));
  nand_5 g00250(.A(pi167), .B(pi147), .Y(new_n627));
  nand_5 g00251(.A(pi181), .B(pi151), .Y(new_n628));
  or_6   g00252(.A(new_n628), .B(new_n627), .Y(new_n629));
  nand_5 g00253(.A(new_n629), .B(new_n626), .Y(new_n630));
  xor_4  g00254(.A(new_n630), .B(new_n623), .Y(new_n631));
  nand_5 g00255(.A(pi151), .B(pi149), .Y(new_n632));
  nand_5 g00256(.A(new_n632), .B(new_n627), .Y(new_n633));
  nand_5 g00257(.A(pi240), .B(pi019), .Y(new_n634));
  xor_4  g00258(.A(new_n632), .B(new_n627), .Y(new_n635));
  nand_5 g00259(.A(new_n635), .B(new_n634), .Y(new_n636));
  nand_5 g00260(.A(new_n636), .B(new_n633), .Y(new_n637));
  xor_4  g00261(.A(new_n637), .B(new_n631), .Y(new_n638));
  nand_5 g00262(.A(pi240), .B(pi097), .Y(new_n639));
  nand_5 g00263(.A(pi134), .B(pi075), .Y(new_n640));
  and_6  g00264(.A(new_n640), .B(new_n639), .Y(new_n641));
  nand_5 g00265(.A(pi134), .B(pi097), .Y(new_n642));
  nand_5 g00266(.A(pi240), .B(pi075), .Y(new_n643));
  nor_5  g00267(.A(new_n643), .B(new_n642), .Y(new_n644));
  or_6   g00268(.A(new_n644), .B(new_n641), .Y(new_n645));
  xnor_4 g00269(.A(new_n645), .B(new_n638), .Y(new_n646));
  nand_5 g00270(.A(pi134), .B(pi019), .Y(new_n647));
  nand_5 g00271(.A(pi240), .B(pi151), .Y(new_n648));
  nand_5 g00272(.A(new_n648), .B(new_n647), .Y(new_n649));
  nand_5 g00273(.A(pi149), .B(pi147), .Y(new_n650));
  xor_4  g00274(.A(new_n648), .B(new_n647), .Y(new_n651));
  nand_5 g00275(.A(new_n651), .B(new_n650), .Y(new_n652));
  nand_5 g00276(.A(new_n652), .B(new_n649), .Y(new_n653));
  nand_5 g00277(.A(new_n653), .B(new_n642), .Y(new_n654));
  xor_4  g00278(.A(new_n635), .B(new_n634), .Y(new_n655));
  xor_4  g00279(.A(new_n653), .B(new_n642), .Y(new_n656));
  nand_5 g00280(.A(new_n656), .B(new_n655), .Y(new_n657));
  nand_5 g00281(.A(new_n657), .B(new_n654), .Y(new_n658));
  xor_4  g00282(.A(new_n658), .B(new_n646), .Y(new_n659));
  nand_5 g00283(.A(pi175), .B(pi075), .Y(new_n660));
  not_8  g00284(.A(new_n660), .Y(new_n661));
  nand_5 g00285(.A(pi240), .B(pi147), .Y(new_n662));
  nand_5 g00286(.A(pi175), .B(pi019), .Y(new_n663));
  nand_5 g00287(.A(new_n663), .B(new_n662), .Y(new_n664));
  nand_5 g00288(.A(pi151), .B(pi134), .Y(new_n665));
  or_6   g00289(.A(new_n663), .B(new_n662), .Y(new_n666));
  nand_5 g00290(.A(new_n666), .B(new_n665), .Y(new_n667));
  nand_5 g00291(.A(new_n667), .B(new_n664), .Y(new_n668));
  nand_5 g00292(.A(pi175), .B(pi097), .Y(new_n669));
  or_6   g00293(.A(new_n669), .B(new_n668), .Y(new_n670));
  xor_4  g00294(.A(new_n651), .B(new_n650), .Y(new_n671));
  not_8  g00295(.A(new_n671), .Y(new_n672));
  xor_4  g00296(.A(new_n669), .B(new_n668), .Y(new_n673));
  nand_5 g00297(.A(new_n673), .B(new_n672), .Y(new_n674));
  nand_5 g00298(.A(new_n674), .B(new_n670), .Y(new_n675));
  nand_5 g00299(.A(new_n675), .B(new_n661), .Y(new_n676));
  xor_4  g00300(.A(new_n656), .B(new_n655), .Y(new_n677));
  xor_4  g00301(.A(new_n675), .B(new_n660), .Y(new_n678));
  or_6   g00302(.A(new_n678), .B(new_n677), .Y(new_n679));
  nand_5 g00303(.A(new_n679), .B(new_n676), .Y(new_n680));
  nand_5 g00304(.A(new_n680), .B(new_n659), .Y(new_n681));
  nand_5 g00305(.A(pi167), .B(pi019), .Y(new_n682));
  nand_5 g00306(.A(pi200), .B(pi147), .Y(new_n683));
  xor_4  g00307(.A(new_n683), .B(new_n682), .Y(new_n684));
  xor_4  g00308(.A(new_n684), .B(new_n628), .Y(new_n685));
  nand_5 g00309(.A(pi149), .B(pi097), .Y(new_n686));
  xor_4  g00310(.A(new_n686), .B(new_n629), .Y(new_n687));
  xor_4  g00311(.A(new_n687), .B(new_n685), .Y(new_n688));
  nand_5 g00312(.A(pi134), .B(pi093), .Y(new_n689));
  nand_5 g00313(.A(pi175), .B(pi166), .Y(new_n690));
  xor_4  g00314(.A(new_n690), .B(new_n689), .Y(new_n691));
  xor_4  g00315(.A(new_n691), .B(new_n643), .Y(new_n692));
  nand_5 g00316(.A(new_n630), .B(new_n623), .Y(new_n693));
  nand_5 g00317(.A(new_n637), .B(new_n631), .Y(new_n694));
  nand_5 g00318(.A(new_n694), .B(new_n693), .Y(new_n695));
  xor_4  g00319(.A(new_n695), .B(new_n692), .Y(new_n696));
  xnor_4 g00320(.A(new_n696), .B(new_n688), .Y(new_n697));
  nor_5  g00321(.A(new_n645), .B(new_n638), .Y(new_n698));
  nor_5  g00322(.A(new_n658), .B(new_n646), .Y(new_n699));
  xor_4  g00323(.A(new_n699), .B(new_n644), .Y(new_n700));
  nor_5  g00324(.A(new_n700), .B(new_n698), .Y(new_n701));
  xor_4  g00325(.A(new_n701), .B(new_n697), .Y(new_n702));
  xor_4  g00326(.A(new_n702), .B(new_n681), .Y(new_n703));
  nand_5 g00327(.A(pi175), .B(pi093), .Y(new_n704));
  xnor_4 g00328(.A(new_n680), .B(new_n659), .Y(new_n705));
  nor_5  g00329(.A(new_n705), .B(new_n704), .Y(new_n706));
  xor_4  g00330(.A(new_n673), .B(new_n671), .Y(new_n707));
  not_8  g00331(.A(new_n665), .Y(new_n708));
  not_8  g00332(.A(new_n664), .Y(new_n709));
  nand_5 g00333(.A(pi175), .B(pi147), .Y(new_n710));
  nand_5 g00334(.A(new_n710), .B(new_n708), .Y(new_n711));
  nand_5 g00335(.A(new_n711), .B(new_n709), .Y(new_n712));
  nand_5 g00336(.A(new_n712), .B(new_n666), .Y(new_n713));
  nand_5 g00337(.A(new_n713), .B(new_n708), .Y(new_n714));
  nor_5  g00338(.A(new_n714), .B(new_n707), .Y(new_n715));
  xor_4  g00339(.A(new_n678), .B(new_n677), .Y(new_n716));
  nand_5 g00340(.A(new_n716), .B(new_n715), .Y(new_n717));
  xor_4  g00341(.A(new_n705), .B(new_n704), .Y(new_n718));
  not_8  g00342(.A(new_n718), .Y(new_n719));
  nor_5  g00343(.A(new_n719), .B(new_n717), .Y(new_n720));
  or_6   g00344(.A(new_n720), .B(new_n706), .Y(new_n721));
  xor_4  g00345(.A(new_n721), .B(new_n703), .Y(new_n722));
  xor_4  g00346(.A(new_n722), .B(new_n622), .Y(new_n723));
  xor_4  g00347(.A(new_n619), .B(new_n585), .Y(new_n724));
  xor_4  g00348(.A(new_n719), .B(new_n717), .Y(new_n725));
  nand_5 g00349(.A(new_n725), .B(new_n724), .Y(new_n726));
  xor_4  g00350(.A(new_n716), .B(new_n715), .Y(new_n727));
  xor_4  g00351(.A(new_n714), .B(new_n707), .Y(new_n728));
  xnor_4 g00352(.A(new_n606), .B(new_n605), .Y(new_n729));
  nor_5  g00353(.A(new_n711), .B(new_n709), .Y(new_n730));
  nor_5  g00354(.A(new_n730), .B(new_n713), .Y(new_n731));
  nand_5 g00355(.A(new_n731), .B(new_n729), .Y(new_n732));
  xor_4  g00356(.A(new_n731), .B(new_n729), .Y(new_n733));
  xor_4  g00357(.A(new_n566), .B(new_n470), .Y(new_n734));
  not_8  g00358(.A(new_n734), .Y(new_n735));
  nor_5  g00359(.A(new_n735), .B(new_n710), .Y(new_n736));
  nand_5 g00360(.A(pi175), .B(pi151), .Y(new_n737));
  nand_5 g00361(.A(pi147), .B(pi134), .Y(new_n738));
  xor_4  g00362(.A(new_n738), .B(new_n737), .Y(new_n739));
  nand_5 g00363(.A(new_n739), .B(new_n736), .Y(new_n740));
  xor_4  g00364(.A(new_n598), .B(new_n597), .Y(new_n741));
  not_8  g00365(.A(new_n741), .Y(new_n742));
  xor_4  g00366(.A(new_n739), .B(new_n736), .Y(new_n743));
  nand_5 g00367(.A(new_n743), .B(new_n742), .Y(new_n744));
  nand_5 g00368(.A(new_n744), .B(new_n740), .Y(new_n745));
  nand_5 g00369(.A(new_n745), .B(new_n733), .Y(new_n746));
  nand_5 g00370(.A(new_n746), .B(new_n732), .Y(new_n747));
  nand_5 g00371(.A(new_n747), .B(new_n728), .Y(new_n748));
  xnor_4 g00372(.A(new_n611), .B(new_n610), .Y(new_n749));
  xor_4  g00373(.A(new_n747), .B(new_n728), .Y(new_n750));
  nand_5 g00374(.A(new_n750), .B(new_n749), .Y(new_n751));
  nand_5 g00375(.A(new_n751), .B(new_n748), .Y(new_n752));
  nand_5 g00376(.A(new_n752), .B(new_n727), .Y(new_n753));
  xor_4  g00377(.A(new_n617), .B(new_n615), .Y(new_n754));
  xor_4  g00378(.A(new_n752), .B(new_n727), .Y(new_n755));
  nand_5 g00379(.A(new_n755), .B(new_n754), .Y(new_n756));
  nand_5 g00380(.A(new_n756), .B(new_n753), .Y(new_n757));
  xor_4  g00381(.A(new_n725), .B(new_n724), .Y(new_n758));
  nand_5 g00382(.A(new_n758), .B(new_n757), .Y(new_n759));
  nand_5 g00383(.A(new_n759), .B(new_n726), .Y(new_n760));
  xor_4  g00384(.A(new_n760), .B(new_n723), .Y(new_n761));
  nand_5 g00385(.A(pi250), .B(pi080), .Y(new_n762));
  nand_5 g00386(.A(pi080), .B(pi045), .Y(new_n763));
  nand_5 g00387(.A(pi247), .B(pi119), .Y(new_n764));
  nand_5 g00388(.A(new_n764), .B(new_n763), .Y(new_n765));
  nand_5 g00389(.A(pi250), .B(pi016), .Y(new_n766));
  xor_4  g00390(.A(new_n764), .B(new_n763), .Y(new_n767));
  nand_5 g00391(.A(new_n767), .B(new_n766), .Y(new_n768));
  nand_5 g00392(.A(new_n768), .B(new_n765), .Y(new_n769));
  xor_4  g00393(.A(new_n769), .B(new_n762), .Y(new_n770));
  nand_5 g00394(.A(pi247), .B(pi045), .Y(new_n771));
  nand_5 g00395(.A(pi234), .B(pi119), .Y(new_n772));
  nand_5 g00396(.A(new_n772), .B(new_n771), .Y(new_n773));
  nand_5 g00397(.A(pi234), .B(pi045), .Y(new_n774));
  nor_5  g00398(.A(new_n774), .B(new_n764), .Y(new_n775));
  not_8  g00399(.A(new_n775), .Y(new_n776));
  nand_5 g00400(.A(new_n776), .B(new_n773), .Y(new_n777));
  xor_4  g00401(.A(new_n777), .B(new_n770), .Y(new_n778));
  nand_5 g00402(.A(pi117), .B(pi054), .Y(new_n779));
  nand_5 g00403(.A(pi044), .B(pi016), .Y(new_n780));
  and_6  g00404(.A(new_n780), .B(new_n779), .Y(new_n781));
  nand_5 g00405(.A(pi117), .B(pi044), .Y(new_n782));
  nand_5 g00406(.A(pi054), .B(pi016), .Y(new_n783));
  nor_5  g00407(.A(new_n783), .B(new_n782), .Y(new_n784));
  or_6   g00408(.A(new_n784), .B(new_n781), .Y(new_n785));
  xnor_4 g00409(.A(new_n785), .B(new_n778), .Y(new_n786));
  nand_5 g00410(.A(pi119), .B(pi080), .Y(new_n787));
  nand_5 g00411(.A(pi045), .B(pi016), .Y(new_n788));
  nand_5 g00412(.A(new_n788), .B(new_n787), .Y(new_n789));
  nand_5 g00413(.A(pi250), .B(pi117), .Y(new_n790));
  xor_4  g00414(.A(new_n788), .B(new_n787), .Y(new_n791));
  nand_5 g00415(.A(new_n791), .B(new_n790), .Y(new_n792));
  nand_5 g00416(.A(new_n792), .B(new_n789), .Y(new_n793));
  nand_5 g00417(.A(new_n793), .B(new_n782), .Y(new_n794));
  xor_4  g00418(.A(new_n767), .B(new_n766), .Y(new_n795));
  xor_4  g00419(.A(new_n793), .B(new_n782), .Y(new_n796));
  nand_5 g00420(.A(new_n796), .B(new_n795), .Y(new_n797));
  nand_5 g00421(.A(new_n797), .B(new_n794), .Y(new_n798));
  xor_4  g00422(.A(new_n798), .B(new_n786), .Y(new_n799));
  xor_4  g00423(.A(new_n796), .B(new_n795), .Y(new_n800));
  nand_5 g00424(.A(pi103), .B(pi054), .Y(new_n801));
  or_6   g00425(.A(new_n801), .B(new_n800), .Y(new_n802));
  xor_4  g00426(.A(new_n801), .B(new_n800), .Y(new_n803));
  nand_5 g00427(.A(pi103), .B(pi044), .Y(new_n804));
  nand_5 g00428(.A(pi117), .B(pi045), .Y(new_n805));
  nand_5 g00429(.A(pi250), .B(pi103), .Y(new_n806));
  nand_5 g00430(.A(new_n806), .B(new_n805), .Y(new_n807));
  nand_5 g00431(.A(pi119), .B(pi016), .Y(new_n808));
  xor_4  g00432(.A(new_n806), .B(new_n805), .Y(new_n809));
  nand_5 g00433(.A(new_n809), .B(new_n808), .Y(new_n810));
  nand_5 g00434(.A(new_n810), .B(new_n807), .Y(new_n811));
  or_6   g00435(.A(new_n811), .B(new_n804), .Y(new_n812));
  xor_4  g00436(.A(new_n811), .B(new_n804), .Y(new_n813));
  xnor_4 g00437(.A(new_n791), .B(new_n790), .Y(new_n814));
  nand_5 g00438(.A(new_n814), .B(new_n813), .Y(new_n815));
  nand_5 g00439(.A(new_n815), .B(new_n812), .Y(new_n816));
  nand_5 g00440(.A(new_n816), .B(new_n803), .Y(new_n817));
  nand_5 g00441(.A(new_n817), .B(new_n802), .Y(new_n818));
  nand_5 g00442(.A(new_n818), .B(new_n799), .Y(new_n819));
  nand_5 g00443(.A(pi250), .B(pi247), .Y(new_n820));
  nand_5 g00444(.A(pi214), .B(pi119), .Y(new_n821));
  xor_4  g00445(.A(new_n821), .B(new_n820), .Y(new_n822));
  xor_4  g00446(.A(new_n822), .B(new_n774), .Y(new_n823));
  nand_5 g00447(.A(pi080), .B(pi044), .Y(new_n824));
  xor_4  g00448(.A(new_n824), .B(new_n776), .Y(new_n825));
  not_8  g00449(.A(new_n825), .Y(new_n826));
  xor_4  g00450(.A(new_n826), .B(new_n823), .Y(new_n827));
  nand_5 g00451(.A(pi248), .B(pi103), .Y(new_n828));
  nand_5 g00452(.A(pi117), .B(pi072), .Y(new_n829));
  xor_4  g00453(.A(new_n829), .B(new_n783), .Y(new_n830));
  xor_4  g00454(.A(new_n830), .B(new_n828), .Y(new_n831));
  nand_5 g00455(.A(new_n769), .B(new_n762), .Y(new_n832));
  nand_5 g00456(.A(new_n777), .B(new_n770), .Y(new_n833));
  nand_5 g00457(.A(new_n833), .B(new_n832), .Y(new_n834));
  xor_4  g00458(.A(new_n834), .B(new_n831), .Y(new_n835));
  xor_4  g00459(.A(new_n835), .B(new_n827), .Y(new_n836));
  nor_5  g00460(.A(new_n798), .B(new_n786), .Y(new_n837));
  nand_5 g00461(.A(new_n837), .B(new_n784), .Y(new_n838));
  nor_5  g00462(.A(new_n785), .B(new_n778), .Y(new_n839));
  or_6   g00463(.A(new_n839), .B(new_n784), .Y(new_n840));
  or_6   g00464(.A(new_n840), .B(new_n837), .Y(new_n841));
  nand_5 g00465(.A(new_n841), .B(new_n838), .Y(new_n842));
  xor_4  g00466(.A(new_n842), .B(new_n836), .Y(new_n843));
  xnor_4 g00467(.A(new_n843), .B(new_n819), .Y(new_n844));
  xor_4  g00468(.A(new_n809), .B(new_n808), .Y(new_n845));
  nand_5 g00469(.A(pi119), .B(pi103), .Y(new_n846));
  nor_5  g00470(.A(new_n846), .B(new_n805), .Y(new_n847));
  not_8  g00471(.A(new_n847), .Y(new_n848));
  nor_5  g00472(.A(new_n848), .B(new_n845), .Y(new_n849));
  not_8  g00473(.A(new_n849), .Y(new_n850));
  xnor_4 g00474(.A(new_n814), .B(new_n813), .Y(new_n851));
  nor_5  g00475(.A(new_n851), .B(new_n850), .Y(new_n852));
  xor_4  g00476(.A(new_n816), .B(new_n803), .Y(new_n853));
  nand_5 g00477(.A(new_n853), .B(new_n852), .Y(new_n854));
  nand_5 g00478(.A(pi103), .B(pi072), .Y(new_n855));
  nand_5 g00479(.A(new_n855), .B(new_n854), .Y(new_n856));
  xor_4  g00480(.A(new_n818), .B(new_n799), .Y(new_n857));
  not_8  g00481(.A(new_n857), .Y(new_n858));
  xor_4  g00482(.A(new_n855), .B(new_n854), .Y(new_n859));
  nand_5 g00483(.A(new_n859), .B(new_n858), .Y(new_n860));
  nand_5 g00484(.A(new_n860), .B(new_n856), .Y(new_n861));
  xor_4  g00485(.A(new_n861), .B(new_n844), .Y(new_n862));
  not_8  g00486(.A(new_n862), .Y(new_n863));
  xor_4  g00487(.A(new_n863), .B(new_n761), .Y(new_n864));
  xor_4  g00488(.A(new_n859), .B(new_n857), .Y(new_n865));
  xnor_4 g00489(.A(new_n853), .B(new_n852), .Y(new_n866));
  xnor_4 g00490(.A(new_n750), .B(new_n749), .Y(new_n867));
  xor_4  g00491(.A(new_n851), .B(new_n850), .Y(new_n868));
  not_8  g00492(.A(new_n868), .Y(new_n869));
  nand_5 g00493(.A(new_n869), .B(new_n867), .Y(new_n870));
  xor_4  g00494(.A(new_n847), .B(new_n845), .Y(new_n871));
  xor_4  g00495(.A(new_n734), .B(new_n710), .Y(new_n872));
  nor_5  g00496(.A(new_n872), .B(new_n846), .Y(new_n873));
  not_8  g00497(.A(new_n873), .Y(new_n874));
  nand_5 g00498(.A(pi103), .B(pi045), .Y(new_n875));
  nand_5 g00499(.A(pi119), .B(pi117), .Y(new_n876));
  nand_5 g00500(.A(new_n876), .B(new_n875), .Y(new_n877));
  nand_5 g00501(.A(new_n877), .B(new_n848), .Y(new_n878));
  nand_5 g00502(.A(new_n878), .B(new_n874), .Y(new_n879));
  xor_4  g00503(.A(new_n743), .B(new_n741), .Y(new_n880));
  xor_4  g00504(.A(new_n878), .B(new_n874), .Y(new_n881));
  nand_5 g00505(.A(new_n881), .B(new_n880), .Y(new_n882));
  nand_5 g00506(.A(new_n882), .B(new_n879), .Y(new_n883));
  nand_5 g00507(.A(new_n883), .B(new_n871), .Y(new_n884));
  xor_4  g00508(.A(new_n745), .B(new_n733), .Y(new_n885));
  not_8  g00509(.A(new_n885), .Y(new_n886));
  xor_4  g00510(.A(new_n883), .B(new_n871), .Y(new_n887));
  nand_5 g00511(.A(new_n887), .B(new_n886), .Y(new_n888));
  nand_5 g00512(.A(new_n888), .B(new_n884), .Y(new_n889));
  xor_4  g00513(.A(new_n869), .B(new_n867), .Y(new_n890));
  nand_5 g00514(.A(new_n890), .B(new_n889), .Y(new_n891));
  nand_5 g00515(.A(new_n891), .B(new_n870), .Y(new_n892));
  or_6   g00516(.A(new_n892), .B(new_n866), .Y(new_n893));
  xor_4  g00517(.A(new_n755), .B(new_n754), .Y(new_n894));
  xor_4  g00518(.A(new_n892), .B(new_n866), .Y(new_n895));
  nand_5 g00519(.A(new_n895), .B(new_n894), .Y(new_n896));
  nand_5 g00520(.A(new_n896), .B(new_n893), .Y(new_n897));
  or_6   g00521(.A(new_n897), .B(new_n865), .Y(new_n898));
  xor_4  g00522(.A(new_n758), .B(new_n757), .Y(new_n899));
  not_8  g00523(.A(new_n899), .Y(new_n900));
  xor_4  g00524(.A(new_n897), .B(new_n865), .Y(new_n901));
  nand_5 g00525(.A(new_n901), .B(new_n900), .Y(new_n902));
  nand_5 g00526(.A(new_n902), .B(new_n898), .Y(new_n903));
  xnor_4 g00527(.A(new_n903), .B(new_n864), .Y(po001));
  nand_5 g00528(.A(pi171), .B(pi042), .Y(new_n905));
  nand_5 g00529(.A(pi108), .B(pi107), .Y(new_n906));
  xor_4  g00530(.A(new_n906), .B(new_n905), .Y(new_n907));
  nand_5 g00531(.A(pi051), .B(pi049), .Y(new_n908));
  xor_4  g00532(.A(new_n908), .B(new_n907), .Y(new_n909));
  nand_5 g00533(.A(pi107), .B(pi051), .Y(new_n910));
  nor_5  g00534(.A(new_n910), .B(new_n905), .Y(new_n911));
  not_8  g00535(.A(new_n911), .Y(new_n912));
  or_6   g00536(.A(new_n912), .B(new_n909), .Y(new_n913));
  nand_5 g00537(.A(pi107), .B(pi007), .Y(new_n914));
  nand_5 g00538(.A(new_n906), .B(new_n905), .Y(new_n915));
  nand_5 g00539(.A(new_n908), .B(new_n907), .Y(new_n916));
  nand_5 g00540(.A(new_n916), .B(new_n915), .Y(new_n917));
  xor_4  g00541(.A(new_n917), .B(new_n914), .Y(new_n918));
  nand_5 g00542(.A(pi171), .B(pi108), .Y(new_n919));
  nand_5 g00543(.A(pi245), .B(pi051), .Y(new_n920));
  nand_5 g00544(.A(pi049), .B(pi042), .Y(new_n921));
  xor_4  g00545(.A(new_n921), .B(new_n920), .Y(new_n922));
  xor_4  g00546(.A(new_n922), .B(new_n919), .Y(new_n923));
  xor_4  g00547(.A(new_n923), .B(new_n918), .Y(new_n924));
  xor_4  g00548(.A(new_n924), .B(new_n913), .Y(new_n925));
  nand_5 g00549(.A(pi178), .B(pi148), .Y(new_n926));
  nand_5 g00550(.A(pi163), .B(pi061), .Y(new_n927));
  xor_4  g00551(.A(new_n927), .B(new_n926), .Y(new_n928));
  nand_5 g00552(.A(pi228), .B(pi188), .Y(new_n929));
  xor_4  g00553(.A(new_n929), .B(new_n928), .Y(new_n930));
  nand_5 g00554(.A(pi188), .B(pi163), .Y(new_n931));
  nor_5  g00555(.A(new_n931), .B(new_n926), .Y(new_n932));
  not_8  g00556(.A(new_n932), .Y(new_n933));
  or_6   g00557(.A(new_n933), .B(new_n930), .Y(new_n934));
  nand_5 g00558(.A(pi148), .B(pi061), .Y(new_n935));
  nand_5 g00559(.A(pi188), .B(pi039), .Y(new_n936));
  nand_5 g00560(.A(pi228), .B(pi178), .Y(new_n937));
  xor_4  g00561(.A(new_n937), .B(new_n936), .Y(new_n938));
  xor_4  g00562(.A(new_n938), .B(new_n935), .Y(new_n939));
  nand_5 g00563(.A(pi163), .B(pi012), .Y(new_n940));
  nand_5 g00564(.A(new_n927), .B(new_n926), .Y(new_n941));
  nand_5 g00565(.A(new_n929), .B(new_n928), .Y(new_n942));
  nand_5 g00566(.A(new_n942), .B(new_n941), .Y(new_n943));
  xor_4  g00567(.A(new_n943), .B(new_n940), .Y(new_n944));
  xor_4  g00568(.A(new_n944), .B(new_n939), .Y(new_n945));
  xor_4  g00569(.A(new_n945), .B(new_n934), .Y(new_n946));
  xor_4  g00570(.A(new_n946), .B(new_n925), .Y(new_n947));
  xor_4  g00571(.A(new_n932), .B(new_n930), .Y(new_n948));
  xor_4  g00572(.A(new_n912), .B(new_n909), .Y(new_n949));
  not_8  g00573(.A(new_n949), .Y(new_n950));
  nor_5  g00574(.A(new_n950), .B(new_n948), .Y(new_n951));
  xor_4  g00575(.A(new_n949), .B(new_n948), .Y(new_n952));
  nand_5 g00576(.A(pi107), .B(pi042), .Y(new_n953));
  nand_5 g00577(.A(pi171), .B(pi051), .Y(new_n954));
  nand_5 g00578(.A(new_n954), .B(new_n953), .Y(new_n955));
  nand_5 g00579(.A(new_n955), .B(new_n912), .Y(new_n956));
  nand_5 g00580(.A(pi178), .B(pi163), .Y(new_n957));
  nand_5 g00581(.A(pi188), .B(pi148), .Y(new_n958));
  nand_5 g00582(.A(new_n958), .B(new_n957), .Y(new_n959));
  nand_5 g00583(.A(new_n959), .B(new_n933), .Y(new_n960));
  nand_5 g00584(.A(new_n960), .B(new_n956), .Y(new_n961));
  nor_5  g00585(.A(new_n931), .B(new_n910), .Y(new_n962));
  not_8  g00586(.A(new_n962), .Y(new_n963));
  xor_4  g00587(.A(new_n960), .B(new_n956), .Y(new_n964));
  nand_5 g00588(.A(new_n964), .B(new_n963), .Y(new_n965));
  nand_5 g00589(.A(new_n965), .B(new_n961), .Y(new_n966));
  nor_5  g00590(.A(new_n966), .B(new_n952), .Y(new_n967));
  nor_5  g00591(.A(new_n967), .B(new_n951), .Y(new_n968));
  not_8  g00592(.A(new_n968), .Y(new_n969));
  xor_4  g00593(.A(new_n969), .B(new_n947), .Y(new_n970));
  nand_5 g00594(.A(pi240), .B(pi162), .Y(new_n971));
  nand_5 g00595(.A(pi179), .B(pi175), .Y(new_n972));
  nand_5 g00596(.A(new_n972), .B(new_n971), .Y(new_n973));
  nand_5 g00597(.A(pi134), .B(pi033), .Y(new_n974));
  or_6   g00598(.A(new_n972), .B(new_n971), .Y(new_n975));
  nand_5 g00599(.A(new_n975), .B(new_n974), .Y(new_n976));
  nand_5 g00600(.A(new_n976), .B(new_n973), .Y(new_n977));
  nand_5 g00601(.A(pi175), .B(pi048), .Y(new_n978));
  xor_4  g00602(.A(new_n978), .B(new_n977), .Y(new_n979));
  nand_5 g00603(.A(pi179), .B(pi134), .Y(new_n980));
  nand_5 g00604(.A(pi162), .B(pi149), .Y(new_n981));
  nand_5 g00605(.A(pi240), .B(pi033), .Y(new_n982));
  xor_4  g00606(.A(new_n982), .B(new_n981), .Y(new_n983));
  xnor_4 g00607(.A(new_n983), .B(new_n980), .Y(new_n984));
  xnor_4 g00608(.A(new_n984), .B(new_n979), .Y(new_n985));
  not_8  g00609(.A(new_n974), .Y(new_n986));
  not_8  g00610(.A(new_n973), .Y(new_n987));
  nand_5 g00611(.A(pi175), .B(pi162), .Y(new_n988));
  nand_5 g00612(.A(new_n988), .B(new_n986), .Y(new_n989));
  nand_5 g00613(.A(new_n989), .B(new_n987), .Y(new_n990));
  nand_5 g00614(.A(new_n990), .B(new_n975), .Y(new_n991));
  nand_5 g00615(.A(new_n991), .B(new_n986), .Y(new_n992));
  xor_4  g00616(.A(new_n992), .B(new_n985), .Y(new_n993));
  xor_4  g00617(.A(new_n966), .B(new_n952), .Y(new_n994));
  nor_5  g00618(.A(new_n989), .B(new_n987), .Y(new_n995));
  nor_5  g00619(.A(new_n995), .B(new_n991), .Y(new_n996));
  nor_5  g00620(.A(new_n996), .B(new_n994), .Y(new_n997));
  xnor_4 g00621(.A(new_n996), .B(new_n994), .Y(new_n998));
  xor_4  g00622(.A(new_n931), .B(new_n910), .Y(new_n999));
  not_8  g00623(.A(new_n999), .Y(new_n1000));
  nor_5  g00624(.A(new_n1000), .B(new_n988), .Y(new_n1001));
  nand_5 g00625(.A(pi162), .B(pi134), .Y(new_n1002));
  nand_5 g00626(.A(pi175), .B(pi033), .Y(new_n1003));
  xor_4  g00627(.A(new_n1003), .B(new_n1002), .Y(new_n1004));
  nand_5 g00628(.A(new_n1004), .B(new_n1001), .Y(new_n1005));
  xor_4  g00629(.A(new_n964), .B(new_n962), .Y(new_n1006));
  xor_4  g00630(.A(new_n1004), .B(new_n1001), .Y(new_n1007));
  nand_5 g00631(.A(new_n1007), .B(new_n1006), .Y(new_n1008));
  nand_5 g00632(.A(new_n1008), .B(new_n1005), .Y(new_n1009));
  nor_5  g00633(.A(new_n1009), .B(new_n998), .Y(new_n1010));
  nor_5  g00634(.A(new_n1010), .B(new_n997), .Y(new_n1011));
  xor_4  g00635(.A(new_n1011), .B(new_n993), .Y(new_n1012));
  xor_4  g00636(.A(new_n1012), .B(new_n970), .Y(new_n1013));
  nand_5 g00637(.A(pi117), .B(pi057), .Y(new_n1014));
  nand_5 g00638(.A(pi194), .B(pi103), .Y(new_n1015));
  xor_4  g00639(.A(new_n1015), .B(new_n1014), .Y(new_n1016));
  nand_5 g00640(.A(pi143), .B(pi016), .Y(new_n1017));
  xor_4  g00641(.A(new_n1017), .B(new_n1016), .Y(new_n1018));
  nand_5 g00642(.A(pi143), .B(pi103), .Y(new_n1019));
  nor_5  g00643(.A(new_n1019), .B(new_n1014), .Y(new_n1020));
  not_8  g00644(.A(new_n1020), .Y(new_n1021));
  or_6   g00645(.A(new_n1021), .B(new_n1018), .Y(new_n1022));
  nand_5 g00646(.A(pi143), .B(pi080), .Y(new_n1023));
  nand_5 g00647(.A(pi194), .B(pi117), .Y(new_n1024));
  nand_5 g00648(.A(pi057), .B(pi016), .Y(new_n1025));
  xor_4  g00649(.A(new_n1025), .B(new_n1024), .Y(new_n1026));
  xor_4  g00650(.A(new_n1026), .B(new_n1023), .Y(new_n1027));
  nand_5 g00651(.A(pi103), .B(pi085), .Y(new_n1028));
  nand_5 g00652(.A(new_n1015), .B(new_n1014), .Y(new_n1029));
  nand_5 g00653(.A(new_n1017), .B(new_n1016), .Y(new_n1030));
  nand_5 g00654(.A(new_n1030), .B(new_n1029), .Y(new_n1031));
  xor_4  g00655(.A(new_n1031), .B(new_n1028), .Y(new_n1032));
  xor_4  g00656(.A(new_n1032), .B(new_n1027), .Y(new_n1033));
  xor_4  g00657(.A(new_n1033), .B(new_n1022), .Y(new_n1034));
  xor_4  g00658(.A(new_n1020), .B(new_n1018), .Y(new_n1035));
  xor_4  g00659(.A(new_n999), .B(new_n988), .Y(new_n1036));
  or_6   g00660(.A(new_n1036), .B(new_n1019), .Y(new_n1037));
  nand_5 g00661(.A(pi103), .B(pi057), .Y(new_n1038));
  nand_5 g00662(.A(pi143), .B(pi117), .Y(new_n1039));
  nand_5 g00663(.A(new_n1039), .B(new_n1038), .Y(new_n1040));
  nand_5 g00664(.A(new_n1040), .B(new_n1021), .Y(new_n1041));
  nand_5 g00665(.A(new_n1041), .B(new_n1037), .Y(new_n1042));
  xor_4  g00666(.A(new_n1007), .B(new_n1006), .Y(new_n1043));
  not_8  g00667(.A(new_n1043), .Y(new_n1044));
  xor_4  g00668(.A(new_n1041), .B(new_n1037), .Y(new_n1045));
  nand_5 g00669(.A(new_n1045), .B(new_n1044), .Y(new_n1046));
  nand_5 g00670(.A(new_n1046), .B(new_n1042), .Y(new_n1047));
  or_6   g00671(.A(new_n1047), .B(new_n1035), .Y(new_n1048));
  xnor_4 g00672(.A(new_n1009), .B(new_n998), .Y(new_n1049));
  xor_4  g00673(.A(new_n1047), .B(new_n1035), .Y(new_n1050));
  nand_5 g00674(.A(new_n1050), .B(new_n1049), .Y(new_n1051));
  nand_5 g00675(.A(new_n1051), .B(new_n1048), .Y(new_n1052));
  xor_4  g00676(.A(new_n1052), .B(new_n1034), .Y(new_n1053));
  xor_4  g00677(.A(new_n1053), .B(new_n1013), .Y(po002));
  nand_5 g00678(.A(pi164), .B(pi142), .Y(new_n1055));
  nand_5 g00679(.A(pi087), .B(pi027), .Y(new_n1056));
  xor_4  g00680(.A(new_n1056), .B(new_n1055), .Y(new_n1057));
  nand_5 g00681(.A(pi147), .B(pi138), .Y(new_n1058));
  xor_4  g00682(.A(new_n1058), .B(new_n1057), .Y(new_n1059));
  nand_5 g00683(.A(pi160), .B(pi119), .Y(new_n1060));
  xor_4  g00684(.A(new_n1060), .B(new_n1059), .Y(po003));
  nand_5 g00685(.A(pi222), .B(pi208), .Y(new_n1062));
  nand_5 g00686(.A(pi168), .B(pi125), .Y(new_n1063));
  xor_4  g00687(.A(new_n1063), .B(new_n1062), .Y(new_n1064));
  nand_5 g00688(.A(pi249), .B(pi139), .Y(new_n1065));
  xor_4  g00689(.A(new_n1065), .B(new_n1064), .Y(new_n1066));
  nand_5 g00690(.A(pi249), .B(pi168), .Y(new_n1067));
  nor_5  g00691(.A(new_n1067), .B(new_n1062), .Y(new_n1068));
  not_8  g00692(.A(new_n1068), .Y(new_n1069));
  or_6   g00693(.A(new_n1069), .B(new_n1066), .Y(new_n1070));
  nand_5 g00694(.A(pi208), .B(pi125), .Y(new_n1071));
  nand_5 g00695(.A(pi249), .B(pi035), .Y(new_n1072));
  nand_5 g00696(.A(pi222), .B(pi139), .Y(new_n1073));
  xor_4  g00697(.A(new_n1073), .B(new_n1072), .Y(new_n1074));
  xor_4  g00698(.A(new_n1074), .B(new_n1071), .Y(new_n1075));
  nand_5 g00699(.A(pi176), .B(pi168), .Y(new_n1076));
  nand_5 g00700(.A(new_n1063), .B(new_n1062), .Y(new_n1077));
  nand_5 g00701(.A(new_n1065), .B(new_n1064), .Y(new_n1078));
  nand_5 g00702(.A(new_n1078), .B(new_n1077), .Y(new_n1079));
  xor_4  g00703(.A(new_n1079), .B(new_n1076), .Y(new_n1080));
  xor_4  g00704(.A(new_n1080), .B(new_n1075), .Y(new_n1081));
  xor_4  g00705(.A(new_n1081), .B(new_n1070), .Y(new_n1082));
  nand_5 g00706(.A(pi242), .B(pi161), .Y(new_n1083));
  nand_5 g00707(.A(pi252), .B(pi236), .Y(new_n1084));
  nand_5 g00708(.A(new_n1084), .B(new_n1083), .Y(new_n1085));
  nand_5 g00709(.A(pi241), .B(pi140), .Y(new_n1086));
  or_6   g00710(.A(new_n1084), .B(new_n1083), .Y(new_n1087));
  nand_5 g00711(.A(new_n1087), .B(new_n1086), .Y(new_n1088));
  nand_5 g00712(.A(new_n1088), .B(new_n1085), .Y(new_n1089));
  nand_5 g00713(.A(pi236), .B(pi121), .Y(new_n1090));
  xor_4  g00714(.A(new_n1090), .B(new_n1089), .Y(new_n1091));
  nand_5 g00715(.A(pi161), .B(pi140), .Y(new_n1092));
  nand_5 g00716(.A(pi242), .B(pi141), .Y(new_n1093));
  nand_5 g00717(.A(pi252), .B(pi241), .Y(new_n1094));
  xor_4  g00718(.A(new_n1094), .B(new_n1093), .Y(new_n1095));
  xnor_4 g00719(.A(new_n1095), .B(new_n1092), .Y(new_n1096));
  xnor_4 g00720(.A(new_n1096), .B(new_n1091), .Y(new_n1097));
  not_8  g00721(.A(new_n1086), .Y(new_n1098));
  not_8  g00722(.A(new_n1085), .Y(new_n1099));
  nand_5 g00723(.A(pi242), .B(pi236), .Y(new_n1100));
  nand_5 g00724(.A(new_n1100), .B(new_n1098), .Y(new_n1101));
  nand_5 g00725(.A(new_n1101), .B(new_n1099), .Y(new_n1102));
  nand_5 g00726(.A(new_n1102), .B(new_n1087), .Y(new_n1103));
  nand_5 g00727(.A(new_n1103), .B(new_n1098), .Y(new_n1104));
  xnor_4 g00728(.A(new_n1104), .B(new_n1097), .Y(new_n1105));
  nand_5 g00729(.A(pi111), .B(pi104), .Y(new_n1106));
  nand_5 g00730(.A(pi210), .B(pi013), .Y(new_n1107));
  nand_5 g00731(.A(pi212), .B(pi024), .Y(new_n1108));
  xor_4  g00732(.A(new_n1108), .B(new_n1107), .Y(new_n1109));
  xor_4  g00733(.A(new_n1109), .B(new_n1106), .Y(new_n1110));
  nand_5 g00734(.A(pi210), .B(pi104), .Y(new_n1111));
  nand_5 g00735(.A(pi213), .B(pi024), .Y(new_n1112));
  nand_5 g00736(.A(new_n1112), .B(new_n1111), .Y(new_n1113));
  nand_5 g00737(.A(pi212), .B(pi111), .Y(new_n1114));
  or_6   g00738(.A(new_n1112), .B(new_n1111), .Y(new_n1115));
  nand_5 g00739(.A(new_n1115), .B(new_n1114), .Y(new_n1116));
  nand_5 g00740(.A(new_n1116), .B(new_n1113), .Y(new_n1117));
  nand_5 g00741(.A(pi224), .B(pi213), .Y(new_n1118));
  xor_4  g00742(.A(new_n1118), .B(new_n1117), .Y(new_n1119));
  xor_4  g00743(.A(new_n1119), .B(new_n1110), .Y(new_n1120));
  not_8  g00744(.A(new_n1114), .Y(new_n1121));
  not_8  g00745(.A(new_n1113), .Y(new_n1122));
  nand_5 g00746(.A(pi213), .B(pi210), .Y(new_n1123));
  nand_5 g00747(.A(new_n1123), .B(new_n1121), .Y(new_n1124));
  nand_5 g00748(.A(new_n1124), .B(new_n1122), .Y(new_n1125));
  nand_5 g00749(.A(new_n1125), .B(new_n1115), .Y(new_n1126));
  nand_5 g00750(.A(new_n1126), .B(new_n1121), .Y(new_n1127));
  xor_4  g00751(.A(new_n1127), .B(new_n1120), .Y(new_n1128));
  xor_4  g00752(.A(new_n1128), .B(new_n1105), .Y(new_n1129));
  nor_5  g00753(.A(new_n1101), .B(new_n1099), .Y(new_n1130));
  or_6   g00754(.A(new_n1130), .B(new_n1103), .Y(new_n1131));
  nor_5  g00755(.A(new_n1124), .B(new_n1122), .Y(new_n1132));
  nor_5  g00756(.A(new_n1132), .B(new_n1126), .Y(new_n1133));
  not_8  g00757(.A(new_n1133), .Y(new_n1134));
  nand_5 g00758(.A(new_n1134), .B(new_n1131), .Y(new_n1135));
  nand_5 g00759(.A(pi212), .B(pi210), .Y(new_n1136));
  nand_5 g00760(.A(pi213), .B(pi111), .Y(new_n1137));
  xor_4  g00761(.A(new_n1137), .B(new_n1136), .Y(new_n1138));
  nand_5 g00762(.A(pi242), .B(pi241), .Y(new_n1139));
  nand_5 g00763(.A(pi236), .B(pi140), .Y(new_n1140));
  xor_4  g00764(.A(new_n1140), .B(new_n1139), .Y(new_n1141));
  or_6   g00765(.A(new_n1141), .B(new_n1138), .Y(new_n1142));
  nor_5  g00766(.A(new_n1123), .B(new_n1100), .Y(new_n1143));
  not_8  g00767(.A(new_n1143), .Y(new_n1144));
  xor_4  g00768(.A(new_n1141), .B(new_n1138), .Y(new_n1145));
  nand_5 g00769(.A(new_n1145), .B(new_n1144), .Y(new_n1146));
  nand_5 g00770(.A(new_n1146), .B(new_n1142), .Y(new_n1147));
  xor_4  g00771(.A(new_n1134), .B(new_n1131), .Y(new_n1148));
  nand_5 g00772(.A(new_n1148), .B(new_n1147), .Y(new_n1149));
  nand_5 g00773(.A(new_n1149), .B(new_n1135), .Y(new_n1150));
  xor_4  g00774(.A(new_n1150), .B(new_n1129), .Y(new_n1151));
  xor_4  g00775(.A(new_n1151), .B(new_n1082), .Y(new_n1152));
  xor_4  g00776(.A(new_n1148), .B(new_n1147), .Y(new_n1153));
  xor_4  g00777(.A(new_n1069), .B(new_n1066), .Y(new_n1154));
  not_8  g00778(.A(new_n1154), .Y(new_n1155));
  or_6   g00779(.A(new_n1155), .B(new_n1153), .Y(new_n1156));
  xor_4  g00780(.A(new_n1155), .B(new_n1153), .Y(new_n1157));
  xor_4  g00781(.A(new_n1123), .B(new_n1100), .Y(new_n1158));
  not_8  g00782(.A(new_n1158), .Y(new_n1159));
  or_6   g00783(.A(new_n1159), .B(new_n1067), .Y(new_n1160));
  nand_5 g00784(.A(pi222), .B(pi168), .Y(new_n1161));
  nand_5 g00785(.A(pi249), .B(pi208), .Y(new_n1162));
  nand_5 g00786(.A(new_n1162), .B(new_n1161), .Y(new_n1163));
  nand_5 g00787(.A(new_n1163), .B(new_n1069), .Y(new_n1164));
  or_6   g00788(.A(new_n1164), .B(new_n1160), .Y(new_n1165));
  xor_4  g00789(.A(new_n1145), .B(new_n1143), .Y(new_n1166));
  xor_4  g00790(.A(new_n1164), .B(new_n1160), .Y(new_n1167));
  nand_5 g00791(.A(new_n1167), .B(new_n1166), .Y(new_n1168));
  nand_5 g00792(.A(new_n1168), .B(new_n1165), .Y(new_n1169));
  nand_5 g00793(.A(new_n1169), .B(new_n1157), .Y(new_n1170));
  nand_5 g00794(.A(new_n1170), .B(new_n1156), .Y(new_n1171));
  xor_4  g00795(.A(new_n1171), .B(new_n1152), .Y(new_n1172));
  nand_5 g00796(.A(pi100), .B(pi077), .Y(new_n1173));
  nand_5 g00797(.A(pi217), .B(pi133), .Y(new_n1174));
  nand_5 g00798(.A(pi227), .B(pi052), .Y(new_n1175));
  xor_4  g00799(.A(new_n1175), .B(new_n1174), .Y(new_n1176));
  xor_4  g00800(.A(new_n1176), .B(new_n1173), .Y(new_n1177));
  nand_5 g00801(.A(pi217), .B(pi077), .Y(new_n1178));
  nand_5 g00802(.A(pi227), .B(pi131), .Y(new_n1179));
  nand_5 g00803(.A(new_n1179), .B(new_n1178), .Y(new_n1180));
  nand_5 g00804(.A(pi100), .B(pi052), .Y(new_n1181));
  or_6   g00805(.A(new_n1179), .B(new_n1178), .Y(new_n1182));
  nand_5 g00806(.A(new_n1182), .B(new_n1181), .Y(new_n1183));
  nand_5 g00807(.A(new_n1183), .B(new_n1180), .Y(new_n1184));
  nand_5 g00808(.A(pi131), .B(pi081), .Y(new_n1185));
  xor_4  g00809(.A(new_n1185), .B(new_n1184), .Y(new_n1186));
  xor_4  g00810(.A(new_n1186), .B(new_n1177), .Y(new_n1187));
  not_8  g00811(.A(new_n1181), .Y(new_n1188));
  not_8  g00812(.A(new_n1180), .Y(new_n1189));
  nand_5 g00813(.A(pi217), .B(pi131), .Y(new_n1190));
  nand_5 g00814(.A(new_n1190), .B(new_n1188), .Y(new_n1191));
  nand_5 g00815(.A(new_n1191), .B(new_n1189), .Y(new_n1192));
  nand_5 g00816(.A(new_n1192), .B(new_n1182), .Y(new_n1193));
  nand_5 g00817(.A(new_n1193), .B(new_n1188), .Y(new_n1194));
  xnor_4 g00818(.A(new_n1194), .B(new_n1187), .Y(new_n1195));
  xor_4  g00819(.A(new_n1158), .B(new_n1067), .Y(new_n1196));
  nor_5  g00820(.A(new_n1196), .B(new_n1190), .Y(new_n1197));
  nand_5 g00821(.A(pi217), .B(pi052), .Y(new_n1198));
  nand_5 g00822(.A(pi131), .B(pi100), .Y(new_n1199));
  xor_4  g00823(.A(new_n1199), .B(new_n1198), .Y(new_n1200));
  or_6   g00824(.A(new_n1200), .B(new_n1197), .Y(new_n1201));
  xor_4  g00825(.A(new_n1167), .B(new_n1166), .Y(new_n1202));
  not_8  g00826(.A(new_n1202), .Y(new_n1203));
  xor_4  g00827(.A(new_n1200), .B(new_n1197), .Y(new_n1204));
  nand_5 g00828(.A(new_n1204), .B(new_n1203), .Y(new_n1205));
  nand_5 g00829(.A(new_n1205), .B(new_n1201), .Y(new_n1206));
  nor_5  g00830(.A(new_n1191), .B(new_n1189), .Y(new_n1207));
  or_6   g00831(.A(new_n1207), .B(new_n1193), .Y(new_n1208));
  nand_5 g00832(.A(new_n1208), .B(new_n1206), .Y(new_n1209));
  xnor_4 g00833(.A(new_n1169), .B(new_n1157), .Y(new_n1210));
  xor_4  g00834(.A(new_n1208), .B(new_n1206), .Y(new_n1211));
  nand_5 g00835(.A(new_n1211), .B(new_n1210), .Y(new_n1212));
  nand_5 g00836(.A(new_n1212), .B(new_n1209), .Y(new_n1213));
  xor_4  g00837(.A(new_n1213), .B(new_n1195), .Y(new_n1214));
  xor_4  g00838(.A(new_n1214), .B(new_n1172), .Y(po004));
  nand_5 g00839(.A(pi192), .B(pi147), .Y(new_n1216));
  nand_5 g00840(.A(pi216), .B(pi019), .Y(new_n1217));
  nand_5 g00841(.A(pi041), .B(pi019), .Y(new_n1218));
  nand_5 g00842(.A(pi147), .B(pi076), .Y(new_n1219));
  nand_5 g00843(.A(new_n1219), .B(new_n1218), .Y(new_n1220));
  nand_5 g00844(.A(pi216), .B(pi151), .Y(new_n1221));
  xor_4  g00845(.A(new_n1219), .B(new_n1218), .Y(new_n1222));
  nand_5 g00846(.A(new_n1222), .B(new_n1221), .Y(new_n1223));
  nand_5 g00847(.A(new_n1223), .B(new_n1220), .Y(new_n1224));
  nand_5 g00848(.A(pi147), .B(pi079), .Y(new_n1225));
  nand_5 g00849(.A(pi151), .B(pi076), .Y(new_n1226));
  nand_5 g00850(.A(new_n1226), .B(new_n1225), .Y(new_n1227));
  nand_5 g00851(.A(pi151), .B(pi079), .Y(new_n1228));
  or_6   g00852(.A(new_n1228), .B(new_n1219), .Y(new_n1229));
  nand_5 g00853(.A(new_n1229), .B(new_n1227), .Y(new_n1230));
  xor_4  g00854(.A(new_n1230), .B(new_n1224), .Y(new_n1231));
  xor_4  g00855(.A(new_n1231), .B(new_n1217), .Y(new_n1232));
  nand_5 g00856(.A(pi097), .B(pi041), .Y(new_n1233));
  nand_5 g00857(.A(pi182), .B(pi075), .Y(new_n1234));
  nand_5 g00858(.A(new_n1234), .B(new_n1233), .Y(new_n1235));
  nand_5 g00859(.A(pi182), .B(pi097), .Y(new_n1236));
  nand_5 g00860(.A(pi075), .B(pi041), .Y(new_n1237));
  nor_5  g00861(.A(new_n1237), .B(new_n1236), .Y(new_n1238));
  not_8  g00862(.A(new_n1238), .Y(new_n1239));
  nand_5 g00863(.A(new_n1239), .B(new_n1235), .Y(new_n1240));
  xnor_4 g00864(.A(new_n1240), .B(new_n1232), .Y(new_n1241));
  nand_5 g00865(.A(pi216), .B(pi147), .Y(new_n1242));
  nand_5 g00866(.A(pi151), .B(pi041), .Y(new_n1243));
  nand_5 g00867(.A(new_n1243), .B(new_n1242), .Y(new_n1244));
  nand_5 g00868(.A(pi182), .B(pi019), .Y(new_n1245));
  xor_4  g00869(.A(new_n1243), .B(new_n1242), .Y(new_n1246));
  nand_5 g00870(.A(new_n1246), .B(new_n1245), .Y(new_n1247));
  nand_5 g00871(.A(new_n1247), .B(new_n1244), .Y(new_n1248));
  nand_5 g00872(.A(new_n1248), .B(new_n1236), .Y(new_n1249));
  xor_4  g00873(.A(new_n1222), .B(new_n1221), .Y(new_n1250));
  xor_4  g00874(.A(new_n1248), .B(new_n1236), .Y(new_n1251));
  nand_5 g00875(.A(new_n1251), .B(new_n1250), .Y(new_n1252));
  nand_5 g00876(.A(new_n1252), .B(new_n1249), .Y(new_n1253));
  xor_4  g00877(.A(new_n1253), .B(new_n1241), .Y(new_n1254));
  nand_5 g00878(.A(pi138), .B(pi075), .Y(new_n1255));
  not_8  g00879(.A(new_n1255), .Y(new_n1256));
  nand_5 g00880(.A(pi138), .B(pi097), .Y(new_n1257));
  nand_5 g00881(.A(pi182), .B(pi151), .Y(new_n1258));
  nand_5 g00882(.A(pi138), .B(pi019), .Y(new_n1259));
  nand_5 g00883(.A(new_n1259), .B(new_n1258), .Y(new_n1260));
  nand_5 g00884(.A(pi147), .B(pi041), .Y(new_n1261));
  xor_4  g00885(.A(new_n1259), .B(new_n1258), .Y(new_n1262));
  nand_5 g00886(.A(new_n1262), .B(new_n1261), .Y(new_n1263));
  nand_5 g00887(.A(new_n1263), .B(new_n1260), .Y(new_n1264));
  or_6   g00888(.A(new_n1264), .B(new_n1257), .Y(new_n1265));
  xnor_4 g00889(.A(new_n1246), .B(new_n1245), .Y(new_n1266));
  xor_4  g00890(.A(new_n1264), .B(new_n1257), .Y(new_n1267));
  nand_5 g00891(.A(new_n1267), .B(new_n1266), .Y(new_n1268));
  nand_5 g00892(.A(new_n1268), .B(new_n1265), .Y(new_n1269));
  nand_5 g00893(.A(new_n1269), .B(new_n1256), .Y(new_n1270));
  xor_4  g00894(.A(new_n1251), .B(new_n1250), .Y(new_n1271));
  xor_4  g00895(.A(new_n1269), .B(new_n1255), .Y(new_n1272));
  or_6   g00896(.A(new_n1272), .B(new_n1271), .Y(new_n1273));
  nand_5 g00897(.A(new_n1273), .B(new_n1270), .Y(new_n1274));
  nand_5 g00898(.A(new_n1274), .B(new_n1254), .Y(new_n1275));
  nand_5 g00899(.A(pi076), .B(pi019), .Y(new_n1276));
  nand_5 g00900(.A(pi251), .B(pi147), .Y(new_n1277));
  xor_4  g00901(.A(new_n1277), .B(new_n1276), .Y(new_n1278));
  xor_4  g00902(.A(new_n1278), .B(new_n1228), .Y(new_n1279));
  nand_5 g00903(.A(pi216), .B(pi097), .Y(new_n1280));
  xor_4  g00904(.A(new_n1280), .B(new_n1229), .Y(new_n1281));
  xor_4  g00905(.A(new_n1281), .B(new_n1279), .Y(new_n1282));
  nand_5 g00906(.A(pi166), .B(pi138), .Y(new_n1283));
  nand_5 g00907(.A(pi182), .B(pi093), .Y(new_n1284));
  xor_4  g00908(.A(new_n1284), .B(new_n1283), .Y(new_n1285));
  xor_4  g00909(.A(new_n1285), .B(new_n1237), .Y(new_n1286));
  nand_5 g00910(.A(new_n1230), .B(new_n1224), .Y(new_n1287));
  nand_5 g00911(.A(new_n1231), .B(new_n1217), .Y(new_n1288));
  nand_5 g00912(.A(new_n1288), .B(new_n1287), .Y(new_n1289));
  xor_4  g00913(.A(new_n1289), .B(new_n1286), .Y(new_n1290));
  xnor_4 g00914(.A(new_n1290), .B(new_n1282), .Y(new_n1291));
  nor_5  g00915(.A(new_n1253), .B(new_n1241), .Y(new_n1292));
  and_6  g00916(.A(new_n1292), .B(new_n1238), .Y(new_n1293));
  or_6   g00917(.A(new_n1240), .B(new_n1232), .Y(new_n1294));
  nand_5 g00918(.A(new_n1294), .B(new_n1239), .Y(new_n1295));
  nor_5  g00919(.A(new_n1295), .B(new_n1292), .Y(new_n1296));
  or_6   g00920(.A(new_n1296), .B(new_n1293), .Y(new_n1297));
  xor_4  g00921(.A(new_n1297), .B(new_n1291), .Y(new_n1298));
  xnor_4 g00922(.A(new_n1298), .B(new_n1275), .Y(new_n1299));
  xor_4  g00923(.A(new_n1262), .B(new_n1261), .Y(new_n1300));
  or_6   g00924(.A(new_n1258), .B(new_n1058), .Y(new_n1301));
  or_6   g00925(.A(new_n1301), .B(new_n1300), .Y(new_n1302));
  xnor_4 g00926(.A(new_n1267), .B(new_n1266), .Y(new_n1303));
  nor_5  g00927(.A(new_n1303), .B(new_n1302), .Y(new_n1304));
  xor_4  g00928(.A(new_n1272), .B(new_n1271), .Y(new_n1305));
  nand_5 g00929(.A(new_n1305), .B(new_n1304), .Y(new_n1306));
  nand_5 g00930(.A(pi138), .B(pi093), .Y(new_n1307));
  nand_5 g00931(.A(new_n1307), .B(new_n1306), .Y(new_n1308));
  xnor_4 g00932(.A(new_n1274), .B(new_n1254), .Y(new_n1309));
  xor_4  g00933(.A(new_n1307), .B(new_n1306), .Y(new_n1310));
  nand_5 g00934(.A(new_n1310), .B(new_n1309), .Y(new_n1311));
  nand_5 g00935(.A(new_n1311), .B(new_n1308), .Y(new_n1312));
  xor_4  g00936(.A(new_n1312), .B(new_n1299), .Y(new_n1313));
  nand_5 g00937(.A(pi145), .B(pi071), .Y(new_n1314));
  nand_5 g00938(.A(pi164), .B(pi123), .Y(new_n1315));
  nand_5 g00939(.A(pi206), .B(pi169), .Y(new_n1316));
  nand_5 g00940(.A(new_n1316), .B(new_n1315), .Y(new_n1317));
  nand_5 g00941(.A(pi071), .B(pi032), .Y(new_n1318));
  xor_4  g00942(.A(new_n1316), .B(new_n1315), .Y(new_n1319));
  nand_5 g00943(.A(new_n1319), .B(new_n1318), .Y(new_n1320));
  nand_5 g00944(.A(new_n1320), .B(new_n1317), .Y(new_n1321));
  nand_5 g00945(.A(new_n1321), .B(new_n1314), .Y(new_n1322));
  nand_5 g00946(.A(pi169), .B(pi032), .Y(new_n1323));
  nand_5 g00947(.A(pi206), .B(pi123), .Y(new_n1324));
  nand_5 g00948(.A(pi164), .B(pi099), .Y(new_n1325));
  xor_4  g00949(.A(new_n1325), .B(new_n1324), .Y(new_n1326));
  xor_4  g00950(.A(new_n1326), .B(new_n1323), .Y(new_n1327));
  xor_4  g00951(.A(new_n1321), .B(new_n1314), .Y(new_n1328));
  nand_5 g00952(.A(new_n1328), .B(new_n1327), .Y(new_n1329));
  nand_5 g00953(.A(new_n1329), .B(new_n1322), .Y(new_n1330));
  nand_5 g00954(.A(pi123), .B(pi032), .Y(new_n1331));
  nand_5 g00955(.A(new_n1325), .B(new_n1324), .Y(new_n1332));
  nand_5 g00956(.A(new_n1326), .B(new_n1323), .Y(new_n1333));
  nand_5 g00957(.A(new_n1333), .B(new_n1332), .Y(new_n1334));
  xor_4  g00958(.A(new_n1334), .B(new_n1331), .Y(new_n1335));
  nand_5 g00959(.A(pi206), .B(pi099), .Y(new_n1336));
  nand_5 g00960(.A(pi164), .B(pi023), .Y(new_n1337));
  nand_5 g00961(.A(new_n1337), .B(new_n1336), .Y(new_n1338));
  nand_5 g00962(.A(pi206), .B(pi023), .Y(new_n1339));
  nor_5  g00963(.A(new_n1339), .B(new_n1325), .Y(new_n1340));
  not_8  g00964(.A(new_n1340), .Y(new_n1341));
  nand_5 g00965(.A(new_n1341), .B(new_n1338), .Y(new_n1342));
  xor_4  g00966(.A(new_n1342), .B(new_n1335), .Y(new_n1343));
  nand_5 g00967(.A(pi246), .B(pi071), .Y(new_n1344));
  nand_5 g00968(.A(pi169), .B(pi145), .Y(new_n1345));
  nand_5 g00969(.A(new_n1345), .B(new_n1344), .Y(new_n1346));
  nand_5 g00970(.A(pi246), .B(pi169), .Y(new_n1347));
  or_6   g00971(.A(new_n1347), .B(new_n1314), .Y(new_n1348));
  nand_5 g00972(.A(new_n1348), .B(new_n1346), .Y(new_n1349));
  xor_4  g00973(.A(new_n1349), .B(new_n1343), .Y(new_n1350));
  xnor_4 g00974(.A(new_n1350), .B(new_n1330), .Y(new_n1351));
  nand_5 g00975(.A(pi246), .B(pi142), .Y(new_n1352));
  nand_5 g00976(.A(pi169), .B(pi164), .Y(new_n1353));
  nand_5 g00977(.A(pi142), .B(pi032), .Y(new_n1354));
  nand_5 g00978(.A(new_n1354), .B(new_n1353), .Y(new_n1355));
  nand_5 g00979(.A(pi206), .B(pi071), .Y(new_n1356));
  or_6   g00980(.A(new_n1354), .B(new_n1353), .Y(new_n1357));
  nand_5 g00981(.A(new_n1357), .B(new_n1356), .Y(new_n1358));
  nand_5 g00982(.A(new_n1358), .B(new_n1355), .Y(new_n1359));
  nand_5 g00983(.A(pi145), .B(pi142), .Y(new_n1360));
  nand_5 g00984(.A(new_n1360), .B(new_n1359), .Y(new_n1361));
  xor_4  g00985(.A(new_n1319), .B(new_n1318), .Y(new_n1362));
  xor_4  g00986(.A(new_n1360), .B(new_n1359), .Y(new_n1363));
  nand_5 g00987(.A(new_n1363), .B(new_n1362), .Y(new_n1364));
  nand_5 g00988(.A(new_n1364), .B(new_n1361), .Y(new_n1365));
  or_6   g00989(.A(new_n1365), .B(new_n1352), .Y(new_n1366));
  xnor_4 g00990(.A(new_n1328), .B(new_n1327), .Y(new_n1367));
  xor_4  g00991(.A(new_n1365), .B(new_n1352), .Y(new_n1368));
  nand_5 g00992(.A(new_n1368), .B(new_n1367), .Y(new_n1369));
  nand_5 g00993(.A(new_n1369), .B(new_n1366), .Y(new_n1370));
  xnor_4 g00994(.A(new_n1370), .B(new_n1351), .Y(new_n1371));
  xor_4  g00995(.A(new_n1363), .B(new_n1362), .Y(new_n1372));
  not_8  g00996(.A(new_n1356), .Y(new_n1373));
  not_8  g00997(.A(new_n1355), .Y(new_n1374));
  nand_5 g00998(.A(new_n1373), .B(new_n1055), .Y(new_n1375));
  nand_5 g00999(.A(new_n1375), .B(new_n1374), .Y(new_n1376));
  nand_5 g01000(.A(new_n1376), .B(new_n1357), .Y(new_n1377));
  nand_5 g01001(.A(new_n1377), .B(new_n1373), .Y(new_n1378));
  nor_5  g01002(.A(new_n1378), .B(new_n1372), .Y(new_n1379));
  xor_4  g01003(.A(new_n1368), .B(new_n1367), .Y(new_n1380));
  nand_5 g01004(.A(new_n1380), .B(new_n1379), .Y(new_n1381));
  nand_5 g01005(.A(pi142), .B(pi114), .Y(new_n1382));
  xor_4  g01006(.A(new_n1382), .B(new_n1381), .Y(new_n1383));
  xor_4  g01007(.A(new_n1383), .B(new_n1371), .Y(new_n1384));
  xnor_4 g01008(.A(new_n1380), .B(new_n1379), .Y(new_n1385));
  nand_5 g01009(.A(pi219), .B(pi026), .Y(new_n1386));
  nand_5 g01010(.A(pi087), .B(pi008), .Y(new_n1387));
  xor_4  g01011(.A(new_n1387), .B(new_n1386), .Y(new_n1388));
  nand_5 g01012(.A(pi102), .B(pi027), .Y(new_n1389));
  xor_4  g01013(.A(new_n1389), .B(new_n1388), .Y(new_n1390));
  nor_5  g01014(.A(new_n1386), .B(new_n1056), .Y(new_n1391));
  not_8  g01015(.A(new_n1391), .Y(new_n1392));
  nor_5  g01016(.A(new_n1392), .B(new_n1390), .Y(new_n1393));
  nand_5 g01017(.A(pi087), .B(pi056), .Y(new_n1394));
  nand_5 g01018(.A(new_n1387), .B(new_n1386), .Y(new_n1395));
  nand_5 g01019(.A(new_n1389), .B(new_n1388), .Y(new_n1396));
  nand_5 g01020(.A(new_n1396), .B(new_n1395), .Y(new_n1397));
  xor_4  g01021(.A(new_n1397), .B(new_n1394), .Y(new_n1398));
  nand_5 g01022(.A(pi219), .B(pi008), .Y(new_n1399));
  nand_5 g01023(.A(pi102), .B(pi026), .Y(new_n1400));
  nand_5 g01024(.A(pi027), .B(pi001), .Y(new_n1401));
  xor_4  g01025(.A(new_n1401), .B(new_n1400), .Y(new_n1402));
  xnor_4 g01026(.A(new_n1402), .B(new_n1399), .Y(new_n1403));
  xnor_4 g01027(.A(new_n1403), .B(new_n1398), .Y(new_n1404));
  xor_4  g01028(.A(new_n1404), .B(new_n1393), .Y(new_n1405));
  nand_5 g01029(.A(pi164), .B(pi071), .Y(new_n1406));
  nand_5 g01030(.A(pi206), .B(pi142), .Y(new_n1407));
  xor_4  g01031(.A(new_n1407), .B(new_n1406), .Y(new_n1408));
  not_8  g01032(.A(new_n1408), .Y(new_n1409));
  nand_5 g01033(.A(pi087), .B(pi026), .Y(new_n1410));
  nand_5 g01034(.A(pi219), .B(pi027), .Y(new_n1411));
  nand_5 g01035(.A(new_n1411), .B(new_n1410), .Y(new_n1412));
  nand_5 g01036(.A(new_n1412), .B(new_n1392), .Y(new_n1413));
  nand_5 g01037(.A(new_n1413), .B(new_n1409), .Y(new_n1414));
  nor_5  g01038(.A(new_n1056), .B(new_n1055), .Y(new_n1415));
  xor_4  g01039(.A(new_n1413), .B(new_n1408), .Y(new_n1416));
  or_6   g01040(.A(new_n1416), .B(new_n1415), .Y(new_n1417));
  nand_5 g01041(.A(new_n1417), .B(new_n1414), .Y(new_n1418));
  nor_5  g01042(.A(new_n1375), .B(new_n1374), .Y(new_n1419));
  nor_5  g01043(.A(new_n1419), .B(new_n1377), .Y(new_n1420));
  not_8  g01044(.A(new_n1420), .Y(new_n1421));
  nand_5 g01045(.A(new_n1421), .B(new_n1418), .Y(new_n1422));
  xor_4  g01046(.A(new_n1391), .B(new_n1390), .Y(new_n1423));
  xor_4  g01047(.A(new_n1421), .B(new_n1418), .Y(new_n1424));
  nand_5 g01048(.A(new_n1424), .B(new_n1423), .Y(new_n1425));
  nand_5 g01049(.A(new_n1425), .B(new_n1422), .Y(new_n1426));
  nand_5 g01050(.A(new_n1426), .B(new_n1405), .Y(new_n1427));
  xor_4  g01051(.A(new_n1378), .B(new_n1372), .Y(new_n1428));
  not_8  g01052(.A(new_n1428), .Y(new_n1429));
  xor_4  g01053(.A(new_n1426), .B(new_n1405), .Y(new_n1430));
  nand_5 g01054(.A(new_n1430), .B(new_n1429), .Y(new_n1431));
  nand_5 g01055(.A(new_n1431), .B(new_n1427), .Y(new_n1432));
  nand_5 g01056(.A(new_n1432), .B(new_n1385), .Y(new_n1433));
  not_8  g01057(.A(new_n1393), .Y(new_n1434));
  nor_5  g01058(.A(new_n1404), .B(new_n1434), .Y(new_n1435));
  nand_5 g01059(.A(pi102), .B(pi008), .Y(new_n1436));
  nand_5 g01060(.A(pi026), .B(pi001), .Y(new_n1437));
  nand_5 g01061(.A(pi122), .B(pi027), .Y(new_n1438));
  xor_4  g01062(.A(new_n1438), .B(new_n1437), .Y(new_n1439));
  xor_4  g01063(.A(new_n1439), .B(new_n1436), .Y(new_n1440));
  nand_5 g01064(.A(pi219), .B(pi056), .Y(new_n1441));
  nand_5 g01065(.A(new_n1401), .B(new_n1400), .Y(new_n1442));
  nand_5 g01066(.A(new_n1402), .B(new_n1399), .Y(new_n1443));
  nand_5 g01067(.A(new_n1443), .B(new_n1442), .Y(new_n1444));
  xor_4  g01068(.A(new_n1444), .B(new_n1441), .Y(new_n1445));
  xor_4  g01069(.A(new_n1445), .B(new_n1440), .Y(new_n1446));
  nand_5 g01070(.A(pi136), .B(pi087), .Y(new_n1447));
  xor_4  g01071(.A(new_n1447), .B(new_n1446), .Y(new_n1448));
  or_6   g01072(.A(new_n1397), .B(new_n1394), .Y(new_n1449));
  nand_5 g01073(.A(new_n1403), .B(new_n1398), .Y(new_n1450));
  nand_5 g01074(.A(new_n1450), .B(new_n1449), .Y(new_n1451));
  xor_4  g01075(.A(new_n1451), .B(new_n1448), .Y(new_n1452));
  xnor_4 g01076(.A(new_n1452), .B(new_n1435), .Y(new_n1453));
  xor_4  g01077(.A(new_n1432), .B(new_n1385), .Y(new_n1454));
  nand_5 g01078(.A(new_n1454), .B(new_n1453), .Y(new_n1455));
  nand_5 g01079(.A(new_n1455), .B(new_n1433), .Y(new_n1456));
  nand_5 g01080(.A(pi008), .B(pi001), .Y(new_n1457));
  nand_5 g01081(.A(pi122), .B(pi026), .Y(new_n1458));
  nand_5 g01082(.A(pi135), .B(pi027), .Y(new_n1459));
  nand_5 g01083(.A(new_n1459), .B(new_n1458), .Y(new_n1460));
  nand_5 g01084(.A(pi135), .B(pi026), .Y(new_n1461));
  or_6   g01085(.A(new_n1461), .B(new_n1438), .Y(new_n1462));
  nand_5 g01086(.A(new_n1462), .B(new_n1460), .Y(new_n1463));
  xor_4  g01087(.A(new_n1463), .B(new_n1457), .Y(new_n1464));
  nand_5 g01088(.A(new_n1438), .B(new_n1437), .Y(new_n1465));
  nand_5 g01089(.A(new_n1439), .B(new_n1436), .Y(new_n1466));
  nand_5 g01090(.A(new_n1466), .B(new_n1465), .Y(new_n1467));
  xor_4  g01091(.A(new_n1467), .B(new_n1464), .Y(new_n1468));
  nand_5 g01092(.A(pi102), .B(pi056), .Y(new_n1469));
  nand_5 g01093(.A(pi219), .B(pi136), .Y(new_n1470));
  and_6  g01094(.A(new_n1470), .B(new_n1469), .Y(new_n1471));
  nand_5 g01095(.A(pi136), .B(pi102), .Y(new_n1472));
  nor_5  g01096(.A(new_n1472), .B(new_n1441), .Y(new_n1473));
  or_6   g01097(.A(new_n1473), .B(new_n1471), .Y(new_n1474));
  xnor_4 g01098(.A(new_n1474), .B(new_n1468), .Y(new_n1475));
  nand_5 g01099(.A(new_n1444), .B(new_n1441), .Y(new_n1476));
  nand_5 g01100(.A(new_n1445), .B(new_n1440), .Y(new_n1477));
  nand_5 g01101(.A(new_n1477), .B(new_n1476), .Y(new_n1478));
  xor_4  g01102(.A(new_n1478), .B(new_n1475), .Y(new_n1479));
  or_6   g01103(.A(new_n1447), .B(new_n1446), .Y(new_n1480));
  nand_5 g01104(.A(new_n1451), .B(new_n1448), .Y(new_n1481));
  nand_5 g01105(.A(new_n1481), .B(new_n1480), .Y(new_n1482));
  xnor_4 g01106(.A(new_n1482), .B(new_n1479), .Y(new_n1483));
  nand_5 g01107(.A(new_n1452), .B(new_n1435), .Y(new_n1484));
  nand_5 g01108(.A(pi096), .B(pi087), .Y(new_n1485));
  xor_4  g01109(.A(new_n1485), .B(new_n1484), .Y(new_n1486));
  xor_4  g01110(.A(new_n1486), .B(new_n1483), .Y(new_n1487));
  xor_4  g01111(.A(new_n1487), .B(new_n1456), .Y(new_n1488));
  xor_4  g01112(.A(new_n1488), .B(new_n1384), .Y(new_n1489));
  xor_4  g01113(.A(new_n1310), .B(new_n1309), .Y(new_n1490));
  or_6   g01114(.A(new_n1490), .B(new_n1489), .Y(new_n1491));
  xor_4  g01115(.A(new_n1454), .B(new_n1453), .Y(new_n1492));
  not_8  g01116(.A(new_n1492), .Y(new_n1493));
  xor_4  g01117(.A(new_n1305), .B(new_n1304), .Y(new_n1494));
  nor_5  g01118(.A(new_n1494), .B(new_n1493), .Y(new_n1495));
  xor_4  g01119(.A(new_n1494), .B(new_n1492), .Y(new_n1496));
  xor_4  g01120(.A(new_n1303), .B(new_n1302), .Y(new_n1497));
  xor_4  g01121(.A(new_n1301), .B(new_n1300), .Y(new_n1498));
  not_8  g01122(.A(new_n1057), .Y(new_n1499));
  or_6   g01123(.A(new_n1058), .B(new_n1499), .Y(new_n1500));
  nand_5 g01124(.A(pi151), .B(pi138), .Y(new_n1501));
  nand_5 g01125(.A(pi182), .B(pi147), .Y(new_n1502));
  nand_5 g01126(.A(new_n1502), .B(new_n1501), .Y(new_n1503));
  nand_5 g01127(.A(new_n1503), .B(new_n1301), .Y(new_n1504));
  or_6   g01128(.A(new_n1504), .B(new_n1500), .Y(new_n1505));
  xor_4  g01129(.A(new_n1416), .B(new_n1415), .Y(new_n1506));
  not_8  g01130(.A(new_n1506), .Y(new_n1507));
  xor_4  g01131(.A(new_n1504), .B(new_n1500), .Y(new_n1508));
  nand_5 g01132(.A(new_n1508), .B(new_n1507), .Y(new_n1509));
  nand_5 g01133(.A(new_n1509), .B(new_n1505), .Y(new_n1510));
  nand_5 g01134(.A(new_n1510), .B(new_n1498), .Y(new_n1511));
  xnor_4 g01135(.A(new_n1424), .B(new_n1423), .Y(new_n1512));
  xor_4  g01136(.A(new_n1510), .B(new_n1498), .Y(new_n1513));
  nand_5 g01137(.A(new_n1513), .B(new_n1512), .Y(new_n1514));
  nand_5 g01138(.A(new_n1514), .B(new_n1511), .Y(new_n1515));
  nand_5 g01139(.A(new_n1515), .B(new_n1497), .Y(new_n1516));
  xor_4  g01140(.A(new_n1430), .B(new_n1428), .Y(new_n1517));
  xor_4  g01141(.A(new_n1515), .B(new_n1497), .Y(new_n1518));
  nand_5 g01142(.A(new_n1518), .B(new_n1517), .Y(new_n1519));
  nand_5 g01143(.A(new_n1519), .B(new_n1516), .Y(new_n1520));
  nor_5  g01144(.A(new_n1520), .B(new_n1496), .Y(new_n1521));
  nor_5  g01145(.A(new_n1521), .B(new_n1495), .Y(new_n1522));
  xor_4  g01146(.A(new_n1490), .B(new_n1489), .Y(new_n1523));
  nand_5 g01147(.A(new_n1523), .B(new_n1522), .Y(new_n1524));
  nand_5 g01148(.A(new_n1524), .B(new_n1491), .Y(new_n1525));
  or_6   g01149(.A(new_n1525), .B(new_n1313), .Y(new_n1526));
  nand_5 g01150(.A(new_n1382), .B(new_n1381), .Y(new_n1527));
  nand_5 g01151(.A(new_n1383), .B(new_n1371), .Y(new_n1528));
  nand_5 g01152(.A(new_n1528), .B(new_n1527), .Y(new_n1529));
  nand_5 g01153(.A(new_n1370), .B(new_n1351), .Y(new_n1530));
  nand_5 g01154(.A(pi099), .B(pi032), .Y(new_n1531));
  nand_5 g01155(.A(pi164), .B(pi155), .Y(new_n1532));
  xor_4  g01156(.A(new_n1532), .B(new_n1339), .Y(new_n1533));
  xor_4  g01157(.A(new_n1533), .B(new_n1531), .Y(new_n1534));
  nand_5 g01158(.A(pi145), .B(pi123), .Y(new_n1535));
  xor_4  g01159(.A(new_n1535), .B(new_n1341), .Y(new_n1536));
  not_8  g01160(.A(new_n1536), .Y(new_n1537));
  xor_4  g01161(.A(new_n1537), .B(new_n1534), .Y(new_n1538));
  nand_5 g01162(.A(pi114), .B(pi071), .Y(new_n1539));
  nand_5 g01163(.A(pi142), .B(pi091), .Y(new_n1540));
  xor_4  g01164(.A(new_n1540), .B(new_n1539), .Y(new_n1541));
  xor_4  g01165(.A(new_n1541), .B(new_n1347), .Y(new_n1542));
  nand_5 g01166(.A(new_n1334), .B(new_n1331), .Y(new_n1543));
  nand_5 g01167(.A(new_n1342), .B(new_n1335), .Y(new_n1544));
  nand_5 g01168(.A(new_n1544), .B(new_n1543), .Y(new_n1545));
  xor_4  g01169(.A(new_n1545), .B(new_n1542), .Y(new_n1546));
  xor_4  g01170(.A(new_n1546), .B(new_n1538), .Y(new_n1547));
  nand_5 g01171(.A(new_n1349), .B(new_n1343), .Y(new_n1548));
  nand_5 g01172(.A(new_n1350), .B(new_n1330), .Y(new_n1549));
  nand_5 g01173(.A(new_n1549), .B(new_n1548), .Y(new_n1550));
  xor_4  g01174(.A(new_n1550), .B(new_n1348), .Y(new_n1551));
  xnor_4 g01175(.A(new_n1551), .B(new_n1547), .Y(new_n1552));
  xnor_4 g01176(.A(new_n1552), .B(new_n1530), .Y(new_n1553));
  xor_4  g01177(.A(new_n1553), .B(new_n1529), .Y(new_n1554));
  nand_5 g01178(.A(new_n1485), .B(new_n1484), .Y(new_n1555));
  nand_5 g01179(.A(new_n1486), .B(new_n1483), .Y(new_n1556));
  nand_5 g01180(.A(new_n1556), .B(new_n1555), .Y(new_n1557));
  nand_5 g01181(.A(new_n1482), .B(new_n1479), .Y(new_n1558));
  nand_5 g01182(.A(pi122), .B(pi008), .Y(new_n1559));
  nand_5 g01183(.A(pi059), .B(pi027), .Y(new_n1560));
  xor_4  g01184(.A(new_n1560), .B(new_n1559), .Y(new_n1561));
  xor_4  g01185(.A(new_n1561), .B(new_n1461), .Y(new_n1562));
  not_8  g01186(.A(new_n1562), .Y(new_n1563));
  nand_5 g01187(.A(pi056), .B(pi001), .Y(new_n1564));
  xor_4  g01188(.A(new_n1564), .B(new_n1462), .Y(new_n1565));
  xor_4  g01189(.A(new_n1565), .B(new_n1563), .Y(new_n1566));
  nand_5 g01190(.A(pi235), .B(pi087), .Y(new_n1567));
  nand_5 g01191(.A(pi219), .B(pi096), .Y(new_n1568));
  xor_4  g01192(.A(new_n1568), .B(new_n1472), .Y(new_n1569));
  xor_4  g01193(.A(new_n1569), .B(new_n1567), .Y(new_n1570));
  nand_5 g01194(.A(new_n1463), .B(new_n1457), .Y(new_n1571));
  nand_5 g01195(.A(new_n1467), .B(new_n1464), .Y(new_n1572));
  nand_5 g01196(.A(new_n1572), .B(new_n1571), .Y(new_n1573));
  xor_4  g01197(.A(new_n1573), .B(new_n1570), .Y(new_n1574));
  xor_4  g01198(.A(new_n1574), .B(new_n1566), .Y(new_n1575));
  nor_5  g01199(.A(new_n1474), .B(new_n1468), .Y(new_n1576));
  nor_5  g01200(.A(new_n1478), .B(new_n1475), .Y(new_n1577));
  xor_4  g01201(.A(new_n1577), .B(new_n1473), .Y(new_n1578));
  nor_5  g01202(.A(new_n1578), .B(new_n1576), .Y(new_n1579));
  xor_4  g01203(.A(new_n1579), .B(new_n1575), .Y(new_n1580));
  xor_4  g01204(.A(new_n1580), .B(new_n1558), .Y(new_n1581));
  xor_4  g01205(.A(new_n1581), .B(new_n1557), .Y(new_n1582));
  nand_5 g01206(.A(new_n1487), .B(new_n1456), .Y(new_n1583));
  nand_5 g01207(.A(new_n1488), .B(new_n1384), .Y(new_n1584));
  nand_5 g01208(.A(new_n1584), .B(new_n1583), .Y(new_n1585));
  xor_4  g01209(.A(new_n1585), .B(new_n1582), .Y(new_n1586));
  xor_4  g01210(.A(new_n1586), .B(new_n1554), .Y(new_n1587));
  not_8  g01211(.A(new_n1587), .Y(new_n1588));
  xor_4  g01212(.A(new_n1525), .B(new_n1313), .Y(new_n1589));
  nand_5 g01213(.A(new_n1589), .B(new_n1588), .Y(new_n1590));
  nand_5 g01214(.A(new_n1590), .B(new_n1526), .Y(new_n1591));
  xor_4  g01215(.A(new_n1591), .B(new_n1216), .Y(new_n1592));
  nor_5  g01216(.A(new_n1298), .B(new_n1275), .Y(new_n1593));
  nor_5  g01217(.A(new_n1312), .B(new_n1299), .Y(new_n1594));
  nor_5  g01218(.A(new_n1594), .B(new_n1593), .Y(new_n1595));
  nand_5 g01219(.A(pi137), .B(pi119), .Y(new_n1596));
  nand_5 g01220(.A(pi160), .B(pi009), .Y(new_n1597));
  xor_4  g01221(.A(new_n1597), .B(new_n1596), .Y(new_n1598));
  nand_5 g01222(.A(pi044), .B(pi020), .Y(new_n1599));
  nand_5 g01223(.A(pi060), .B(pi054), .Y(new_n1600));
  or_6   g01224(.A(new_n1600), .B(new_n1599), .Y(new_n1601));
  nand_5 g01225(.A(pi060), .B(pi045), .Y(new_n1602));
  nand_5 g01226(.A(pi223), .B(pi119), .Y(new_n1603));
  nand_5 g01227(.A(new_n1603), .B(new_n1602), .Y(new_n1604));
  nand_5 g01228(.A(pi250), .B(pi020), .Y(new_n1605));
  xor_4  g01229(.A(new_n1603), .B(new_n1602), .Y(new_n1606));
  nand_5 g01230(.A(new_n1606), .B(new_n1605), .Y(new_n1607));
  nand_5 g01231(.A(new_n1607), .B(new_n1604), .Y(new_n1608));
  nand_5 g01232(.A(new_n1608), .B(new_n1599), .Y(new_n1609));
  nand_5 g01233(.A(pi223), .B(pi045), .Y(new_n1610));
  nand_5 g01234(.A(pi250), .B(pi060), .Y(new_n1611));
  nand_5 g01235(.A(pi119), .B(pi101), .Y(new_n1612));
  xor_4  g01236(.A(new_n1612), .B(new_n1611), .Y(new_n1613));
  xor_4  g01237(.A(new_n1613), .B(new_n1610), .Y(new_n1614));
  xor_4  g01238(.A(new_n1608), .B(new_n1599), .Y(new_n1615));
  nand_5 g01239(.A(new_n1615), .B(new_n1614), .Y(new_n1616));
  nand_5 g01240(.A(new_n1616), .B(new_n1609), .Y(new_n1617));
  nand_5 g01241(.A(pi060), .B(pi044), .Y(new_n1618));
  nand_5 g01242(.A(pi054), .B(pi020), .Y(new_n1619));
  nand_5 g01243(.A(new_n1619), .B(new_n1618), .Y(new_n1620));
  nand_5 g01244(.A(new_n1620), .B(new_n1601), .Y(new_n1621));
  nand_5 g01245(.A(new_n1621), .B(new_n1617), .Y(new_n1622));
  nand_5 g01246(.A(pi250), .B(pi223), .Y(new_n1623));
  nand_5 g01247(.A(new_n1612), .B(new_n1611), .Y(new_n1624));
  nand_5 g01248(.A(new_n1613), .B(new_n1610), .Y(new_n1625));
  nand_5 g01249(.A(new_n1625), .B(new_n1624), .Y(new_n1626));
  nand_5 g01250(.A(pi225), .B(pi119), .Y(new_n1627));
  nand_5 g01251(.A(pi101), .B(pi045), .Y(new_n1628));
  nand_5 g01252(.A(new_n1628), .B(new_n1627), .Y(new_n1629));
  nand_5 g01253(.A(pi225), .B(pi045), .Y(new_n1630));
  or_6   g01254(.A(new_n1630), .B(new_n1612), .Y(new_n1631));
  nand_5 g01255(.A(new_n1631), .B(new_n1629), .Y(new_n1632));
  xor_4  g01256(.A(new_n1632), .B(new_n1626), .Y(new_n1633));
  xor_4  g01257(.A(new_n1633), .B(new_n1623), .Y(new_n1634));
  xor_4  g01258(.A(new_n1621), .B(new_n1617), .Y(new_n1635));
  nand_5 g01259(.A(new_n1635), .B(new_n1634), .Y(new_n1636));
  nand_5 g01260(.A(new_n1636), .B(new_n1622), .Y(new_n1637));
  or_6   g01261(.A(new_n1637), .B(new_n1601), .Y(new_n1638));
  xor_4  g01262(.A(new_n1637), .B(new_n1601), .Y(new_n1639));
  nand_5 g01263(.A(pi250), .B(pi101), .Y(new_n1640));
  nand_5 g01264(.A(pi177), .B(pi119), .Y(new_n1641));
  xor_4  g01265(.A(new_n1641), .B(new_n1630), .Y(new_n1642));
  xor_4  g01266(.A(new_n1642), .B(new_n1640), .Y(new_n1643));
  nand_5 g01267(.A(pi223), .B(pi044), .Y(new_n1644));
  xor_4  g01268(.A(new_n1644), .B(new_n1631), .Y(new_n1645));
  not_8  g01269(.A(new_n1645), .Y(new_n1646));
  xor_4  g01270(.A(new_n1646), .B(new_n1643), .Y(new_n1647));
  nand_5 g01271(.A(pi248), .B(pi160), .Y(new_n1648));
  nand_5 g01272(.A(pi072), .B(pi020), .Y(new_n1649));
  xor_4  g01273(.A(new_n1649), .B(new_n1648), .Y(new_n1650));
  xor_4  g01274(.A(new_n1650), .B(new_n1600), .Y(new_n1651));
  nand_5 g01275(.A(new_n1632), .B(new_n1626), .Y(new_n1652));
  nand_5 g01276(.A(new_n1633), .B(new_n1623), .Y(new_n1653));
  nand_5 g01277(.A(new_n1653), .B(new_n1652), .Y(new_n1654));
  xor_4  g01278(.A(new_n1654), .B(new_n1651), .Y(new_n1655));
  xor_4  g01279(.A(new_n1655), .B(new_n1647), .Y(new_n1656));
  nand_5 g01280(.A(new_n1656), .B(new_n1639), .Y(new_n1657));
  nand_5 g01281(.A(new_n1657), .B(new_n1638), .Y(new_n1658));
  xor_4  g01282(.A(new_n1635), .B(new_n1634), .Y(new_n1659));
  not_8  g01283(.A(new_n1659), .Y(new_n1660));
  xor_4  g01284(.A(new_n1615), .B(new_n1614), .Y(new_n1661));
  nand_5 g01285(.A(pi160), .B(pi054), .Y(new_n1662));
  or_6   g01286(.A(new_n1662), .B(new_n1661), .Y(new_n1663));
  xor_4  g01287(.A(new_n1662), .B(new_n1661), .Y(new_n1664));
  nand_5 g01288(.A(pi119), .B(pi060), .Y(new_n1665));
  nand_5 g01289(.A(pi250), .B(pi160), .Y(new_n1666));
  nand_5 g01290(.A(new_n1666), .B(new_n1665), .Y(new_n1667));
  nand_5 g01291(.A(pi045), .B(pi020), .Y(new_n1668));
  or_6   g01292(.A(new_n1666), .B(new_n1665), .Y(new_n1669));
  nand_5 g01293(.A(new_n1669), .B(new_n1668), .Y(new_n1670));
  nand_5 g01294(.A(new_n1670), .B(new_n1667), .Y(new_n1671));
  nand_5 g01295(.A(pi160), .B(pi044), .Y(new_n1672));
  or_6   g01296(.A(new_n1672), .B(new_n1671), .Y(new_n1673));
  xor_4  g01297(.A(new_n1606), .B(new_n1605), .Y(new_n1674));
  not_8  g01298(.A(new_n1674), .Y(new_n1675));
  xor_4  g01299(.A(new_n1672), .B(new_n1671), .Y(new_n1676));
  nand_5 g01300(.A(new_n1676), .B(new_n1675), .Y(new_n1677));
  nand_5 g01301(.A(new_n1677), .B(new_n1673), .Y(new_n1678));
  nand_5 g01302(.A(new_n1678), .B(new_n1664), .Y(new_n1679));
  nand_5 g01303(.A(new_n1679), .B(new_n1663), .Y(new_n1680));
  nand_5 g01304(.A(new_n1680), .B(new_n1660), .Y(new_n1681));
  xnor_4 g01305(.A(new_n1656), .B(new_n1639), .Y(new_n1682));
  nor_5  g01306(.A(new_n1682), .B(new_n1681), .Y(new_n1683));
  xor_4  g01307(.A(new_n1676), .B(new_n1674), .Y(new_n1684));
  not_8  g01308(.A(new_n1668), .Y(new_n1685));
  not_8  g01309(.A(new_n1667), .Y(new_n1686));
  nand_5 g01310(.A(new_n1685), .B(new_n1060), .Y(new_n1687));
  nand_5 g01311(.A(new_n1687), .B(new_n1686), .Y(new_n1688));
  nand_5 g01312(.A(new_n1688), .B(new_n1669), .Y(new_n1689));
  nand_5 g01313(.A(new_n1689), .B(new_n1685), .Y(new_n1690));
  nor_5  g01314(.A(new_n1690), .B(new_n1684), .Y(new_n1691));
  xor_4  g01315(.A(new_n1678), .B(new_n1664), .Y(new_n1692));
  nand_5 g01316(.A(new_n1692), .B(new_n1691), .Y(new_n1693));
  nand_5 g01317(.A(pi160), .B(pi072), .Y(new_n1694));
  nand_5 g01318(.A(new_n1694), .B(new_n1693), .Y(new_n1695));
  xor_4  g01319(.A(new_n1680), .B(new_n1659), .Y(new_n1696));
  xor_4  g01320(.A(new_n1694), .B(new_n1693), .Y(new_n1697));
  nand_5 g01321(.A(new_n1697), .B(new_n1696), .Y(new_n1698));
  nand_5 g01322(.A(new_n1698), .B(new_n1695), .Y(new_n1699));
  xor_4  g01323(.A(new_n1682), .B(new_n1681), .Y(new_n1700));
  not_8  g01324(.A(new_n1700), .Y(new_n1701));
  nor_5  g01325(.A(new_n1701), .B(new_n1699), .Y(new_n1702));
  or_6   g01326(.A(new_n1702), .B(new_n1683), .Y(new_n1703));
  xor_4  g01327(.A(new_n1703), .B(new_n1658), .Y(new_n1704));
  xor_4  g01328(.A(new_n1704), .B(new_n1598), .Y(new_n1705));
  nand_5 g01329(.A(pi102), .B(pi096), .Y(new_n1706));
  nand_5 g01330(.A(pi235), .B(pi219), .Y(new_n1707));
  or_6   g01331(.A(new_n1564), .B(new_n1462), .Y(new_n1708));
  nand_5 g01332(.A(new_n1565), .B(new_n1563), .Y(new_n1709));
  nand_5 g01333(.A(new_n1709), .B(new_n1708), .Y(new_n1710));
  xor_4  g01334(.A(new_n1710), .B(new_n1707), .Y(new_n1711));
  xor_4  g01335(.A(new_n1711), .B(new_n1706), .Y(new_n1712));
  xor_4  g01336(.A(new_n1712), .B(new_n1705), .Y(new_n1713));
  nand_5 g01337(.A(pi110), .B(pi087), .Y(new_n1714));
  nand_5 g01338(.A(pi094), .B(pi027), .Y(new_n1715));
  nand_5 g01339(.A(pi059), .B(pi026), .Y(new_n1716));
  nand_5 g01340(.A(pi135), .B(pi008), .Y(new_n1717));
  xor_4  g01341(.A(new_n1717), .B(new_n1716), .Y(new_n1718));
  nand_5 g01342(.A(new_n1577), .B(new_n1473), .Y(new_n1719));
  not_8  g01343(.A(new_n1579), .Y(new_n1720));
  nand_5 g01344(.A(new_n1720), .B(new_n1575), .Y(new_n1721));
  nand_5 g01345(.A(new_n1721), .B(new_n1719), .Y(new_n1722));
  nand_5 g01346(.A(new_n1540), .B(new_n1539), .Y(new_n1723));
  nand_5 g01347(.A(new_n1541), .B(new_n1347), .Y(new_n1724));
  nand_5 g01348(.A(new_n1724), .B(new_n1723), .Y(new_n1725));
  xor_4  g01349(.A(new_n1725), .B(new_n1722), .Y(new_n1726));
  nand_5 g01350(.A(pi091), .B(pi071), .Y(new_n1727));
  nand_5 g01351(.A(pi169), .B(pi114), .Y(new_n1728));
  xnor_4 g01352(.A(new_n1728), .B(new_n1727), .Y(new_n1729));
  nand_5 g01353(.A(pi145), .B(pi099), .Y(new_n1730));
  xor_4  g01354(.A(new_n1730), .B(new_n1729), .Y(new_n1731));
  nand_5 g01355(.A(new_n1545), .B(new_n1542), .Y(new_n1732));
  not_8  g01356(.A(new_n1538), .Y(new_n1733));
  nand_5 g01357(.A(new_n1546), .B(new_n1733), .Y(new_n1734));
  nand_5 g01358(.A(new_n1734), .B(new_n1732), .Y(new_n1735));
  nand_5 g01359(.A(pi246), .B(pi123), .Y(new_n1736));
  xor_4  g01360(.A(new_n1736), .B(new_n1735), .Y(new_n1737));
  xor_4  g01361(.A(new_n1737), .B(new_n1731), .Y(new_n1738));
  nand_5 g01362(.A(new_n1532), .B(new_n1339), .Y(new_n1739));
  nand_5 g01363(.A(new_n1533), .B(new_n1531), .Y(new_n1740));
  nand_5 g01364(.A(new_n1740), .B(new_n1739), .Y(new_n1741));
  nor_5  g01365(.A(new_n1535), .B(new_n1341), .Y(new_n1742));
  nor_5  g01366(.A(new_n1537), .B(new_n1534), .Y(new_n1743));
  or_6   g01367(.A(new_n1743), .B(new_n1742), .Y(new_n1744));
  xor_4  g01368(.A(new_n1744), .B(new_n1741), .Y(new_n1745));
  xor_4  g01369(.A(new_n1745), .B(new_n1738), .Y(new_n1746));
  xor_4  g01370(.A(new_n1746), .B(new_n1726), .Y(new_n1747));
  xor_4  g01371(.A(new_n1747), .B(new_n1718), .Y(new_n1748));
  xor_4  g01372(.A(new_n1748), .B(new_n1715), .Y(new_n1749));
  xor_4  g01373(.A(new_n1749), .B(new_n1714), .Y(new_n1750));
  nand_5 g01374(.A(new_n1568), .B(new_n1472), .Y(new_n1751));
  nand_5 g01375(.A(new_n1569), .B(new_n1567), .Y(new_n1752));
  nand_5 g01376(.A(new_n1752), .B(new_n1751), .Y(new_n1753));
  nand_5 g01377(.A(new_n1580), .B(new_n1558), .Y(new_n1754));
  nand_5 g01378(.A(new_n1581), .B(new_n1557), .Y(new_n1755));
  nand_5 g01379(.A(new_n1755), .B(new_n1754), .Y(new_n1756));
  nand_5 g01380(.A(pi122), .B(pi056), .Y(new_n1757));
  nand_5 g01381(.A(pi136), .B(pi001), .Y(new_n1758));
  xor_4  g01382(.A(new_n1758), .B(new_n1757), .Y(new_n1759));
  xor_4  g01383(.A(new_n1759), .B(new_n1756), .Y(new_n1760));
  xor_4  g01384(.A(new_n1760), .B(new_n1753), .Y(new_n1761));
  xor_4  g01385(.A(new_n1761), .B(new_n1750), .Y(new_n1762));
  nand_5 g01386(.A(new_n1573), .B(new_n1570), .Y(new_n1763));
  not_8  g01387(.A(new_n1566), .Y(new_n1764));
  nand_5 g01388(.A(new_n1574), .B(new_n1764), .Y(new_n1765));
  nand_5 g01389(.A(new_n1765), .B(new_n1763), .Y(new_n1766));
  nand_5 g01390(.A(new_n1560), .B(new_n1559), .Y(new_n1767));
  nand_5 g01391(.A(new_n1561), .B(new_n1461), .Y(new_n1768));
  nand_5 g01392(.A(new_n1768), .B(new_n1767), .Y(new_n1769));
  xor_4  g01393(.A(new_n1769), .B(new_n1766), .Y(new_n1770));
  xor_4  g01394(.A(new_n1770), .B(new_n1762), .Y(new_n1771));
  xor_4  g01395(.A(new_n1771), .B(new_n1713), .Y(new_n1772));
  nand_5 g01396(.A(new_n1641), .B(new_n1630), .Y(new_n1773));
  nand_5 g01397(.A(new_n1642), .B(new_n1640), .Y(new_n1774));
  nand_5 g01398(.A(new_n1774), .B(new_n1773), .Y(new_n1775));
  nor_5  g01399(.A(new_n1644), .B(new_n1631), .Y(new_n1776));
  nor_5  g01400(.A(new_n1646), .B(new_n1643), .Y(new_n1777));
  or_6   g01401(.A(new_n1777), .B(new_n1776), .Y(new_n1778));
  xor_4  g01402(.A(new_n1778), .B(new_n1775), .Y(new_n1779));
  xor_4  g01403(.A(new_n1779), .B(new_n1772), .Y(new_n1780));
  xor_4  g01404(.A(new_n1780), .B(new_n1595), .Y(new_n1781));
  xor_4  g01405(.A(new_n1781), .B(new_n1592), .Y(new_n1782));
  nand_5 g01406(.A(pi251), .B(pi151), .Y(new_n1783));
  nand_5 g01407(.A(new_n1649), .B(new_n1648), .Y(new_n1784));
  nand_5 g01408(.A(new_n1650), .B(new_n1600), .Y(new_n1785));
  nand_5 g01409(.A(new_n1785), .B(new_n1784), .Y(new_n1786));
  or_6   g01410(.A(new_n1654), .B(new_n1651), .Y(new_n1787));
  nand_5 g01411(.A(new_n1655), .B(new_n1647), .Y(new_n1788));
  nand_5 g01412(.A(new_n1788), .B(new_n1787), .Y(new_n1789));
  xor_4  g01413(.A(new_n1789), .B(new_n1786), .Y(new_n1790));
  xor_4  g01414(.A(new_n1790), .B(new_n1783), .Y(new_n1791));
  xor_4  g01415(.A(new_n1700), .B(new_n1699), .Y(new_n1792));
  xnor_4 g01416(.A(new_n1692), .B(new_n1691), .Y(new_n1793));
  xor_4  g01417(.A(new_n1690), .B(new_n1684), .Y(new_n1794));
  xnor_4 g01418(.A(new_n1513), .B(new_n1512), .Y(new_n1795));
  nor_5  g01419(.A(new_n1060), .B(new_n1059), .Y(new_n1796));
  nand_5 g01420(.A(pi160), .B(pi045), .Y(new_n1797));
  nand_5 g01421(.A(pi119), .B(pi020), .Y(new_n1798));
  xor_4  g01422(.A(new_n1798), .B(new_n1797), .Y(new_n1799));
  or_6   g01423(.A(new_n1799), .B(new_n1796), .Y(new_n1800));
  xor_4  g01424(.A(new_n1508), .B(new_n1507), .Y(new_n1801));
  not_8  g01425(.A(new_n1801), .Y(new_n1802));
  xor_4  g01426(.A(new_n1799), .B(new_n1796), .Y(new_n1803));
  nand_5 g01427(.A(new_n1803), .B(new_n1802), .Y(new_n1804));
  nand_5 g01428(.A(new_n1804), .B(new_n1800), .Y(new_n1805));
  or_6   g01429(.A(new_n1805), .B(new_n1795), .Y(new_n1806));
  xor_4  g01430(.A(new_n1805), .B(new_n1795), .Y(new_n1807));
  nor_5  g01431(.A(new_n1687), .B(new_n1686), .Y(new_n1808));
  nor_5  g01432(.A(new_n1808), .B(new_n1689), .Y(new_n1809));
  nand_5 g01433(.A(new_n1809), .B(new_n1807), .Y(new_n1810));
  nand_5 g01434(.A(new_n1810), .B(new_n1806), .Y(new_n1811));
  or_6   g01435(.A(new_n1811), .B(new_n1794), .Y(new_n1812));
  xor_4  g01436(.A(new_n1518), .B(new_n1517), .Y(new_n1813));
  not_8  g01437(.A(new_n1813), .Y(new_n1814));
  xor_4  g01438(.A(new_n1811), .B(new_n1794), .Y(new_n1815));
  nand_5 g01439(.A(new_n1815), .B(new_n1814), .Y(new_n1816));
  nand_5 g01440(.A(new_n1816), .B(new_n1812), .Y(new_n1817));
  or_6   g01441(.A(new_n1817), .B(new_n1793), .Y(new_n1818));
  xnor_4 g01442(.A(new_n1520), .B(new_n1496), .Y(new_n1819));
  xor_4  g01443(.A(new_n1817), .B(new_n1793), .Y(new_n1820));
  nand_5 g01444(.A(new_n1820), .B(new_n1819), .Y(new_n1821));
  nand_5 g01445(.A(new_n1821), .B(new_n1818), .Y(new_n1822));
  xnor_4 g01446(.A(new_n1697), .B(new_n1696), .Y(new_n1823));
  or_6   g01447(.A(new_n1823), .B(new_n1822), .Y(new_n1824));
  xor_4  g01448(.A(new_n1523), .B(new_n1522), .Y(new_n1825));
  not_8  g01449(.A(new_n1825), .Y(new_n1826));
  xor_4  g01450(.A(new_n1823), .B(new_n1822), .Y(new_n1827));
  nand_5 g01451(.A(new_n1827), .B(new_n1826), .Y(new_n1828));
  nand_5 g01452(.A(new_n1828), .B(new_n1824), .Y(new_n1829));
  or_6   g01453(.A(new_n1829), .B(new_n1792), .Y(new_n1830));
  xor_4  g01454(.A(new_n1589), .B(new_n1587), .Y(new_n1831));
  xor_4  g01455(.A(new_n1829), .B(new_n1792), .Y(new_n1832));
  nand_5 g01456(.A(new_n1832), .B(new_n1831), .Y(new_n1833));
  nand_5 g01457(.A(new_n1833), .B(new_n1830), .Y(new_n1834));
  nand_5 g01458(.A(pi138), .B(pi011), .Y(new_n1835));
  xor_4  g01459(.A(new_n1835), .B(new_n1834), .Y(new_n1836));
  xor_4  g01460(.A(new_n1836), .B(new_n1791), .Y(new_n1837));
  nor_5  g01461(.A(new_n1297), .B(new_n1291), .Y(new_n1838));
  nor_5  g01462(.A(new_n1838), .B(new_n1296), .Y(new_n1839));
  nand_5 g01463(.A(pi177), .B(pi045), .Y(new_n1840));
  nand_5 g01464(.A(pi101), .B(pi044), .Y(new_n1841));
  xor_4  g01465(.A(new_n1841), .B(new_n1840), .Y(new_n1842));
  nand_5 g01466(.A(pi223), .B(pi054), .Y(new_n1843));
  or_6   g01467(.A(new_n1585), .B(new_n1582), .Y(new_n1844));
  nand_5 g01468(.A(new_n1586), .B(new_n1554), .Y(new_n1845));
  nand_5 g01469(.A(new_n1845), .B(new_n1844), .Y(new_n1846));
  nand_5 g01470(.A(pi216), .B(pi075), .Y(new_n1847));
  nand_5 g01471(.A(pi093), .B(pi041), .Y(new_n1848));
  xor_4  g01472(.A(new_n1848), .B(new_n1847), .Y(new_n1849));
  nand_5 g01473(.A(pi097), .B(pi076), .Y(new_n1850));
  nand_5 g01474(.A(new_n1289), .B(new_n1286), .Y(new_n1851));
  nand_5 g01475(.A(new_n1290), .B(new_n1282), .Y(new_n1852));
  nand_5 g01476(.A(new_n1852), .B(new_n1851), .Y(new_n1853));
  xor_4  g01477(.A(new_n1853), .B(new_n1850), .Y(new_n1854));
  xor_4  g01478(.A(new_n1854), .B(new_n1849), .Y(new_n1855));
  xor_4  g01479(.A(new_n1855), .B(new_n1846), .Y(new_n1856));
  or_6   g01480(.A(new_n1550), .B(new_n1348), .Y(new_n1857));
  nand_5 g01481(.A(new_n1551), .B(new_n1547), .Y(new_n1858));
  nand_5 g01482(.A(new_n1858), .B(new_n1857), .Y(new_n1859));
  nand_5 g01483(.A(pi164), .B(pi086), .Y(new_n1860));
  nand_5 g01484(.A(new_n1284), .B(new_n1283), .Y(new_n1861));
  nand_5 g01485(.A(new_n1285), .B(new_n1237), .Y(new_n1862));
  nand_5 g01486(.A(new_n1862), .B(new_n1861), .Y(new_n1863));
  nand_5 g01487(.A(pi206), .B(pi155), .Y(new_n1864));
  nand_5 g01488(.A(pi032), .B(pi023), .Y(new_n1865));
  xor_4  g01489(.A(new_n1865), .B(new_n1864), .Y(new_n1866));
  xor_4  g01490(.A(new_n1866), .B(new_n1863), .Y(new_n1867));
  xor_4  g01491(.A(new_n1867), .B(new_n1860), .Y(new_n1868));
  xor_4  g01492(.A(new_n1868), .B(new_n1859), .Y(new_n1869));
  nand_5 g01493(.A(new_n1277), .B(new_n1276), .Y(new_n1870));
  nand_5 g01494(.A(new_n1278), .B(new_n1228), .Y(new_n1871));
  nand_5 g01495(.A(new_n1871), .B(new_n1870), .Y(new_n1872));
  or_6   g01496(.A(new_n1280), .B(new_n1229), .Y(new_n1873));
  not_8  g01497(.A(new_n1279), .Y(new_n1874));
  nand_5 g01498(.A(new_n1281), .B(new_n1874), .Y(new_n1875));
  nand_5 g01499(.A(new_n1875), .B(new_n1873), .Y(new_n1876));
  xor_4  g01500(.A(new_n1876), .B(new_n1872), .Y(new_n1877));
  nor_5  g01501(.A(new_n1552), .B(new_n1530), .Y(new_n1878));
  nor_5  g01502(.A(new_n1553), .B(new_n1529), .Y(new_n1879));
  nor_5  g01503(.A(new_n1879), .B(new_n1878), .Y(new_n1880));
  nand_5 g01504(.A(pi142), .B(pi031), .Y(new_n1881));
  xor_4  g01505(.A(new_n1881), .B(new_n1880), .Y(new_n1882));
  xor_4  g01506(.A(new_n1882), .B(new_n1877), .Y(new_n1883));
  xor_4  g01507(.A(new_n1883), .B(new_n1869), .Y(new_n1884));
  nand_5 g01508(.A(pi182), .B(pi166), .Y(new_n1885));
  nand_5 g01509(.A(pi079), .B(pi019), .Y(new_n1886));
  xor_4  g01510(.A(new_n1886), .B(new_n1885), .Y(new_n1887));
  xor_4  g01511(.A(new_n1887), .B(new_n1884), .Y(new_n1888));
  xor_4  g01512(.A(new_n1888), .B(new_n1856), .Y(new_n1889));
  xor_4  g01513(.A(new_n1889), .B(new_n1843), .Y(new_n1890));
  xor_4  g01514(.A(new_n1890), .B(new_n1842), .Y(new_n1891));
  nand_5 g01515(.A(pi250), .B(pi225), .Y(new_n1892));
  nand_5 g01516(.A(pi248), .B(pi020), .Y(new_n1893));
  nand_5 g01517(.A(pi072), .B(pi060), .Y(new_n1894));
  xor_4  g01518(.A(new_n1894), .B(new_n1893), .Y(new_n1895));
  xor_4  g01519(.A(new_n1895), .B(new_n1892), .Y(new_n1896));
  xor_4  g01520(.A(new_n1896), .B(new_n1891), .Y(new_n1897));
  xor_4  g01521(.A(new_n1897), .B(new_n1839), .Y(new_n1898));
  xor_4  g01522(.A(new_n1898), .B(new_n1837), .Y(new_n1899));
  xor_4  g01523(.A(new_n1899), .B(new_n1782), .Y(po005));
  nand_5 g01524(.A(pi117), .B(pi067), .Y(new_n1901));
  nand_5 g01525(.A(pi053), .B(pi016), .Y(new_n1902));
  nor_5  g01526(.A(new_n1902), .B(new_n1901), .Y(new_n1903));
  nand_5 g01527(.A(pi229), .B(pi080), .Y(new_n1904));
  nand_5 g01528(.A(pi092), .B(pi080), .Y(new_n1905));
  nand_5 g01529(.A(pi229), .B(pi016), .Y(new_n1906));
  nand_5 g01530(.A(new_n1906), .B(new_n1905), .Y(new_n1907));
  nand_5 g01531(.A(pi247), .B(pi190), .Y(new_n1908));
  xor_4  g01532(.A(new_n1906), .B(new_n1905), .Y(new_n1909));
  nand_5 g01533(.A(new_n1909), .B(new_n1908), .Y(new_n1910));
  nand_5 g01534(.A(new_n1910), .B(new_n1907), .Y(new_n1911));
  xor_4  g01535(.A(new_n1911), .B(new_n1904), .Y(new_n1912));
  nand_5 g01536(.A(pi234), .B(pi190), .Y(new_n1913));
  nand_5 g01537(.A(pi247), .B(pi092), .Y(new_n1914));
  nand_5 g01538(.A(new_n1914), .B(new_n1913), .Y(new_n1915));
  nand_5 g01539(.A(pi234), .B(pi092), .Y(new_n1916));
  or_6   g01540(.A(new_n1916), .B(new_n1908), .Y(new_n1917));
  nand_5 g01541(.A(new_n1917), .B(new_n1915), .Y(new_n1918));
  xor_4  g01542(.A(new_n1918), .B(new_n1912), .Y(new_n1919));
  nand_5 g01543(.A(pi067), .B(pi016), .Y(new_n1920));
  nand_5 g01544(.A(pi117), .B(pi053), .Y(new_n1921));
  and_6  g01545(.A(new_n1921), .B(new_n1920), .Y(new_n1922));
  or_6   g01546(.A(new_n1922), .B(new_n1903), .Y(new_n1923));
  xnor_4 g01547(.A(new_n1923), .B(new_n1919), .Y(new_n1924));
  nand_5 g01548(.A(pi092), .B(pi016), .Y(new_n1925));
  nand_5 g01549(.A(pi190), .B(pi080), .Y(new_n1926));
  nand_5 g01550(.A(new_n1926), .B(new_n1925), .Y(new_n1927));
  nand_5 g01551(.A(pi229), .B(pi117), .Y(new_n1928));
  xor_4  g01552(.A(new_n1926), .B(new_n1925), .Y(new_n1929));
  nand_5 g01553(.A(new_n1929), .B(new_n1928), .Y(new_n1930));
  nand_5 g01554(.A(new_n1930), .B(new_n1927), .Y(new_n1931));
  nand_5 g01555(.A(new_n1931), .B(new_n1901), .Y(new_n1932));
  xor_4  g01556(.A(new_n1909), .B(new_n1908), .Y(new_n1933));
  xor_4  g01557(.A(new_n1931), .B(new_n1901), .Y(new_n1934));
  nand_5 g01558(.A(new_n1934), .B(new_n1933), .Y(new_n1935));
  nand_5 g01559(.A(new_n1935), .B(new_n1932), .Y(new_n1936));
  nor_5  g01560(.A(new_n1936), .B(new_n1924), .Y(new_n1937));
  nand_5 g01561(.A(new_n1937), .B(new_n1903), .Y(new_n1938));
  nand_5 g01562(.A(pi214), .B(pi190), .Y(new_n1939));
  nand_5 g01563(.A(pi247), .B(pi229), .Y(new_n1940));
  xor_4  g01564(.A(new_n1940), .B(new_n1939), .Y(new_n1941));
  xor_4  g01565(.A(new_n1941), .B(new_n1916), .Y(new_n1942));
  nand_5 g01566(.A(pi080), .B(pi067), .Y(new_n1943));
  xor_4  g01567(.A(new_n1943), .B(new_n1917), .Y(new_n1944));
  xor_4  g01568(.A(new_n1944), .B(new_n1942), .Y(new_n1945));
  nand_5 g01569(.A(pi103), .B(pi030), .Y(new_n1946));
  nand_5 g01570(.A(pi185), .B(pi117), .Y(new_n1947));
  xor_4  g01571(.A(new_n1947), .B(new_n1946), .Y(new_n1948));
  xor_4  g01572(.A(new_n1948), .B(new_n1902), .Y(new_n1949));
  nand_5 g01573(.A(new_n1911), .B(new_n1904), .Y(new_n1950));
  nand_5 g01574(.A(new_n1918), .B(new_n1912), .Y(new_n1951));
  nand_5 g01575(.A(new_n1951), .B(new_n1950), .Y(new_n1952));
  xor_4  g01576(.A(new_n1952), .B(new_n1949), .Y(new_n1953));
  xnor_4 g01577(.A(new_n1953), .B(new_n1945), .Y(new_n1954));
  nor_5  g01578(.A(new_n1923), .B(new_n1919), .Y(new_n1955));
  xor_4  g01579(.A(new_n1937), .B(new_n1903), .Y(new_n1956));
  nor_5  g01580(.A(new_n1956), .B(new_n1955), .Y(new_n1957));
  not_8  g01581(.A(new_n1957), .Y(new_n1958));
  nand_5 g01582(.A(new_n1958), .B(new_n1954), .Y(new_n1959));
  nand_5 g01583(.A(new_n1959), .B(new_n1938), .Y(new_n1960));
  xor_4  g01584(.A(new_n1936), .B(new_n1924), .Y(new_n1961));
  xor_4  g01585(.A(new_n1934), .B(new_n1933), .Y(new_n1962));
  nand_5 g01586(.A(pi103), .B(pi053), .Y(new_n1963));
  or_6   g01587(.A(new_n1963), .B(new_n1962), .Y(new_n1964));
  xor_4  g01588(.A(new_n1963), .B(new_n1962), .Y(new_n1965));
  nand_5 g01589(.A(pi103), .B(pi067), .Y(new_n1966));
  nand_5 g01590(.A(pi117), .B(pi092), .Y(new_n1967));
  nand_5 g01591(.A(pi229), .B(pi103), .Y(new_n1968));
  nand_5 g01592(.A(new_n1968), .B(new_n1967), .Y(new_n1969));
  xor_4  g01593(.A(new_n1968), .B(new_n1967), .Y(new_n1970));
  nand_5 g01594(.A(pi190), .B(pi016), .Y(new_n1971));
  nand_5 g01595(.A(new_n1971), .B(new_n1970), .Y(new_n1972));
  nand_5 g01596(.A(new_n1972), .B(new_n1969), .Y(new_n1973));
  or_6   g01597(.A(new_n1973), .B(new_n1966), .Y(new_n1974));
  xor_4  g01598(.A(new_n1973), .B(new_n1966), .Y(new_n1975));
  xor_4  g01599(.A(new_n1929), .B(new_n1928), .Y(new_n1976));
  not_8  g01600(.A(new_n1976), .Y(new_n1977));
  nand_5 g01601(.A(new_n1977), .B(new_n1975), .Y(new_n1978));
  nand_5 g01602(.A(new_n1978), .B(new_n1974), .Y(new_n1979));
  nand_5 g01603(.A(new_n1979), .B(new_n1965), .Y(new_n1980));
  nand_5 g01604(.A(new_n1980), .B(new_n1964), .Y(new_n1981));
  nand_5 g01605(.A(new_n1981), .B(new_n1961), .Y(new_n1982));
  xor_4  g01606(.A(new_n1957), .B(new_n1954), .Y(new_n1983));
  nand_5 g01607(.A(new_n1983), .B(new_n1982), .Y(new_n1984));
  xor_4  g01608(.A(new_n1971), .B(new_n1970), .Y(new_n1985));
  nand_5 g01609(.A(pi190), .B(pi103), .Y(new_n1986));
  nor_5  g01610(.A(new_n1986), .B(new_n1967), .Y(new_n1987));
  not_8  g01611(.A(new_n1987), .Y(new_n1988));
  or_6   g01612(.A(new_n1988), .B(new_n1985), .Y(new_n1989));
  xor_4  g01613(.A(new_n1976), .B(new_n1975), .Y(new_n1990));
  nor_5  g01614(.A(new_n1990), .B(new_n1989), .Y(new_n1991));
  xor_4  g01615(.A(new_n1979), .B(new_n1965), .Y(new_n1992));
  nand_5 g01616(.A(new_n1992), .B(new_n1991), .Y(new_n1993));
  nand_5 g01617(.A(pi185), .B(pi103), .Y(new_n1994));
  nand_5 g01618(.A(new_n1994), .B(new_n1993), .Y(new_n1995));
  xnor_4 g01619(.A(new_n1981), .B(new_n1961), .Y(new_n1996));
  xor_4  g01620(.A(new_n1994), .B(new_n1993), .Y(new_n1997));
  nand_5 g01621(.A(new_n1997), .B(new_n1996), .Y(new_n1998));
  nand_5 g01622(.A(new_n1998), .B(new_n1995), .Y(new_n1999));
  xor_4  g01623(.A(new_n1983), .B(new_n1982), .Y(new_n2000));
  nand_5 g01624(.A(new_n2000), .B(new_n1999), .Y(new_n2001));
  nand_5 g01625(.A(new_n2001), .B(new_n1984), .Y(new_n2002));
  xor_4  g01626(.A(new_n2002), .B(new_n1960), .Y(new_n2003));
  nand_5 g01627(.A(pi107), .B(pi006), .Y(new_n2004));
  nand_5 g01628(.A(pi158), .B(pi049), .Y(new_n2005));
  nand_5 g01629(.A(pi254), .B(pi245), .Y(new_n2006));
  nand_5 g01630(.A(pi171), .B(pi089), .Y(new_n2007));
  xor_4  g01631(.A(new_n2007), .B(new_n2006), .Y(new_n2008));
  xnor_4 g01632(.A(new_n2008), .B(new_n2005), .Y(new_n2009));
  nand_5 g01633(.A(pi254), .B(pi049), .Y(new_n2010));
  nand_5 g01634(.A(pi107), .B(pi089), .Y(new_n2011));
  nand_5 g01635(.A(new_n2011), .B(new_n2010), .Y(new_n2012));
  nand_5 g01636(.A(pi171), .B(pi158), .Y(new_n2013));
  or_6   g01637(.A(new_n2011), .B(new_n2010), .Y(new_n2014));
  nand_5 g01638(.A(new_n2014), .B(new_n2013), .Y(new_n2015));
  nand_5 g01639(.A(new_n2015), .B(new_n2012), .Y(new_n2016));
  nand_5 g01640(.A(pi154), .B(pi107), .Y(new_n2017));
  xor_4  g01641(.A(new_n2017), .B(new_n2016), .Y(new_n2018));
  xnor_4 g01642(.A(new_n2018), .B(new_n2009), .Y(new_n2019));
  not_8  g01643(.A(new_n2013), .Y(new_n2020));
  nand_5 g01644(.A(pi254), .B(pi107), .Y(new_n2021));
  nand_5 g01645(.A(new_n2021), .B(new_n2020), .Y(new_n2022));
  not_8  g01646(.A(new_n2022), .Y(new_n2023));
  or_6   g01647(.A(new_n2023), .B(new_n2012), .Y(new_n2024));
  nand_5 g01648(.A(new_n2024), .B(new_n2014), .Y(new_n2025));
  nand_5 g01649(.A(new_n2025), .B(new_n2020), .Y(new_n2026));
  nor_5  g01650(.A(new_n2026), .B(new_n2019), .Y(new_n2027));
  nand_5 g01651(.A(pi089), .B(pi049), .Y(new_n2028));
  nand_5 g01652(.A(pi245), .B(pi158), .Y(new_n2029));
  nand_5 g01653(.A(pi254), .B(pi201), .Y(new_n2030));
  xor_4  g01654(.A(new_n2030), .B(new_n2029), .Y(new_n2031));
  xor_4  g01655(.A(new_n2031), .B(new_n2028), .Y(new_n2032));
  nand_5 g01656(.A(pi171), .B(pi154), .Y(new_n2033));
  nand_5 g01657(.A(new_n2007), .B(new_n2006), .Y(new_n2034));
  nand_5 g01658(.A(new_n2008), .B(new_n2005), .Y(new_n2035));
  nand_5 g01659(.A(new_n2035), .B(new_n2034), .Y(new_n2036));
  xor_4  g01660(.A(new_n2036), .B(new_n2033), .Y(new_n2037));
  xor_4  g01661(.A(new_n2037), .B(new_n2032), .Y(new_n2038));
  nand_5 g01662(.A(pi107), .B(pi095), .Y(new_n2039));
  or_6   g01663(.A(new_n2017), .B(new_n2016), .Y(new_n2040));
  nand_5 g01664(.A(new_n2018), .B(new_n2009), .Y(new_n2041));
  nand_5 g01665(.A(new_n2041), .B(new_n2040), .Y(new_n2042));
  xor_4  g01666(.A(new_n2042), .B(new_n2039), .Y(new_n2043));
  xor_4  g01667(.A(new_n2043), .B(new_n2038), .Y(new_n2044));
  nand_5 g01668(.A(new_n2044), .B(new_n2027), .Y(new_n2045));
  nand_5 g01669(.A(new_n2045), .B(new_n2004), .Y(new_n2046));
  nand_5 g01670(.A(new_n2036), .B(new_n2033), .Y(new_n2047));
  nand_5 g01671(.A(new_n2037), .B(new_n2032), .Y(new_n2048));
  nand_5 g01672(.A(new_n2048), .B(new_n2047), .Y(new_n2049));
  nand_5 g01673(.A(pi245), .B(pi089), .Y(new_n2050));
  nand_5 g01674(.A(pi254), .B(pi156), .Y(new_n2051));
  nand_5 g01675(.A(pi201), .B(pi158), .Y(new_n2052));
  nand_5 g01676(.A(new_n2052), .B(new_n2051), .Y(new_n2053));
  nand_5 g01677(.A(pi158), .B(pi156), .Y(new_n2054));
  or_6   g01678(.A(new_n2054), .B(new_n2030), .Y(new_n2055));
  nand_5 g01679(.A(new_n2055), .B(new_n2053), .Y(new_n2056));
  xor_4  g01680(.A(new_n2056), .B(new_n2050), .Y(new_n2057));
  nand_5 g01681(.A(new_n2030), .B(new_n2029), .Y(new_n2058));
  nand_5 g01682(.A(new_n2031), .B(new_n2028), .Y(new_n2059));
  nand_5 g01683(.A(new_n2059), .B(new_n2058), .Y(new_n2060));
  xor_4  g01684(.A(new_n2060), .B(new_n2057), .Y(new_n2061));
  nand_5 g01685(.A(pi154), .B(pi049), .Y(new_n2062));
  nand_5 g01686(.A(pi171), .B(pi095), .Y(new_n2063));
  nand_5 g01687(.A(new_n2063), .B(new_n2062), .Y(new_n2064));
  nand_5 g01688(.A(pi095), .B(pi049), .Y(new_n2065));
  or_6   g01689(.A(new_n2065), .B(new_n2033), .Y(new_n2066));
  nand_5 g01690(.A(new_n2066), .B(new_n2064), .Y(new_n2067));
  xor_4  g01691(.A(new_n2067), .B(new_n2061), .Y(new_n2068));
  xor_4  g01692(.A(new_n2068), .B(new_n2049), .Y(new_n2069));
  not_8  g01693(.A(new_n2039), .Y(new_n2070));
  nand_5 g01694(.A(new_n2042), .B(new_n2070), .Y(new_n2071));
  or_6   g01695(.A(new_n2043), .B(new_n2038), .Y(new_n2072));
  nand_5 g01696(.A(new_n2072), .B(new_n2071), .Y(new_n2073));
  xor_4  g01697(.A(new_n2073), .B(new_n2069), .Y(new_n2074));
  xor_4  g01698(.A(new_n2045), .B(new_n2004), .Y(new_n2075));
  nand_5 g01699(.A(new_n2075), .B(new_n2074), .Y(new_n2076));
  nand_5 g01700(.A(new_n2076), .B(new_n2046), .Y(new_n2077));
  not_8  g01701(.A(new_n2069), .Y(new_n2078));
  nand_5 g01702(.A(new_n2073), .B(new_n2078), .Y(new_n2079));
  nand_5 g01703(.A(pi201), .B(pi089), .Y(new_n2080));
  nand_5 g01704(.A(pi254), .B(pi063), .Y(new_n2081));
  xor_4  g01705(.A(new_n2081), .B(new_n2080), .Y(new_n2082));
  xor_4  g01706(.A(new_n2082), .B(new_n2054), .Y(new_n2083));
  not_8  g01707(.A(new_n2083), .Y(new_n2084));
  nand_5 g01708(.A(pi245), .B(pi154), .Y(new_n2085));
  xor_4  g01709(.A(new_n2085), .B(new_n2055), .Y(new_n2086));
  xor_4  g01710(.A(new_n2086), .B(new_n2084), .Y(new_n2087));
  nand_5 g01711(.A(pi171), .B(pi006), .Y(new_n2088));
  nand_5 g01712(.A(pi209), .B(pi107), .Y(new_n2089));
  xor_4  g01713(.A(new_n2089), .B(new_n2088), .Y(new_n2090));
  xor_4  g01714(.A(new_n2090), .B(new_n2065), .Y(new_n2091));
  nand_5 g01715(.A(new_n2056), .B(new_n2050), .Y(new_n2092));
  nand_5 g01716(.A(new_n2060), .B(new_n2057), .Y(new_n2093));
  nand_5 g01717(.A(new_n2093), .B(new_n2092), .Y(new_n2094));
  xor_4  g01718(.A(new_n2094), .B(new_n2091), .Y(new_n2095));
  xor_4  g01719(.A(new_n2095), .B(new_n2087), .Y(new_n2096));
  nand_5 g01720(.A(new_n2067), .B(new_n2061), .Y(new_n2097));
  nand_5 g01721(.A(new_n2068), .B(new_n2049), .Y(new_n2098));
  nand_5 g01722(.A(new_n2098), .B(new_n2097), .Y(new_n2099));
  xor_4  g01723(.A(new_n2099), .B(new_n2066), .Y(new_n2100));
  xnor_4 g01724(.A(new_n2100), .B(new_n2096), .Y(new_n2101));
  xor_4  g01725(.A(new_n2101), .B(new_n2079), .Y(new_n2102));
  xnor_4 g01726(.A(new_n2102), .B(new_n2077), .Y(new_n2103));
  nand_5 g01727(.A(pi073), .B(pi039), .Y(new_n2104));
  nand_5 g01728(.A(pi228), .B(pi073), .Y(new_n2105));
  nand_5 g01729(.A(pi170), .B(pi116), .Y(new_n2106));
  nand_5 g01730(.A(new_n2106), .B(new_n2105), .Y(new_n2107));
  nand_5 g01731(.A(pi039), .B(pi004), .Y(new_n2108));
  xor_4  g01732(.A(new_n2106), .B(new_n2105), .Y(new_n2109));
  nand_5 g01733(.A(new_n2109), .B(new_n2108), .Y(new_n2110));
  nand_5 g01734(.A(new_n2110), .B(new_n2107), .Y(new_n2111));
  xor_4  g01735(.A(new_n2111), .B(new_n2104), .Y(new_n2112));
  nand_5 g01736(.A(pi170), .B(pi070), .Y(new_n2113));
  nand_5 g01737(.A(pi116), .B(pi004), .Y(new_n2114));
  nand_5 g01738(.A(new_n2114), .B(new_n2113), .Y(new_n2115));
  nand_5 g01739(.A(pi070), .B(pi004), .Y(new_n2116));
  nor_5  g01740(.A(new_n2116), .B(new_n2106), .Y(new_n2117));
  not_8  g01741(.A(new_n2117), .Y(new_n2118));
  nand_5 g01742(.A(new_n2118), .B(new_n2115), .Y(new_n2119));
  xor_4  g01743(.A(new_n2119), .B(new_n2112), .Y(new_n2120));
  nand_5 g01744(.A(pi148), .B(pi130), .Y(new_n2121));
  nand_5 g01745(.A(pi228), .B(pi003), .Y(new_n2122));
  and_6  g01746(.A(new_n2122), .B(new_n2121), .Y(new_n2123));
  nand_5 g01747(.A(pi228), .B(pi130), .Y(new_n2124));
  nand_5 g01748(.A(pi148), .B(pi003), .Y(new_n2125));
  nor_5  g01749(.A(new_n2125), .B(new_n2124), .Y(new_n2126));
  or_6   g01750(.A(new_n2126), .B(new_n2123), .Y(new_n2127));
  xnor_4 g01751(.A(new_n2127), .B(new_n2120), .Y(new_n2128));
  nand_5 g01752(.A(pi228), .B(pi004), .Y(new_n2129));
  nand_5 g01753(.A(pi148), .B(pi073), .Y(new_n2130));
  nand_5 g01754(.A(new_n2130), .B(new_n2129), .Y(new_n2131));
  nand_5 g01755(.A(pi170), .B(pi039), .Y(new_n2132));
  xor_4  g01756(.A(new_n2130), .B(new_n2129), .Y(new_n2133));
  nand_5 g01757(.A(new_n2133), .B(new_n2132), .Y(new_n2134));
  nand_5 g01758(.A(new_n2134), .B(new_n2131), .Y(new_n2135));
  nand_5 g01759(.A(new_n2135), .B(new_n2125), .Y(new_n2136));
  xor_4  g01760(.A(new_n2109), .B(new_n2108), .Y(new_n2137));
  xor_4  g01761(.A(new_n2135), .B(new_n2125), .Y(new_n2138));
  nand_5 g01762(.A(new_n2138), .B(new_n2137), .Y(new_n2139));
  nand_5 g01763(.A(new_n2139), .B(new_n2136), .Y(new_n2140));
  xor_4  g01764(.A(new_n2140), .B(new_n2128), .Y(new_n2141));
  nand_5 g01765(.A(pi163), .B(pi130), .Y(new_n2142));
  nand_5 g01766(.A(pi228), .B(pi170), .Y(new_n2143));
  nand_5 g01767(.A(pi163), .B(pi073), .Y(new_n2144));
  nand_5 g01768(.A(new_n2144), .B(new_n2143), .Y(new_n2145));
  nand_5 g01769(.A(pi148), .B(pi004), .Y(new_n2146));
  or_6   g01770(.A(new_n2144), .B(new_n2143), .Y(new_n2147));
  nand_5 g01771(.A(new_n2147), .B(new_n2146), .Y(new_n2148));
  nand_5 g01772(.A(new_n2148), .B(new_n2145), .Y(new_n2149));
  nand_5 g01773(.A(pi163), .B(pi003), .Y(new_n2150));
  nand_5 g01774(.A(new_n2150), .B(new_n2149), .Y(new_n2151));
  xor_4  g01775(.A(new_n2133), .B(new_n2132), .Y(new_n2152));
  xor_4  g01776(.A(new_n2150), .B(new_n2149), .Y(new_n2153));
  nand_5 g01777(.A(new_n2153), .B(new_n2152), .Y(new_n2154));
  nand_5 g01778(.A(new_n2154), .B(new_n2151), .Y(new_n2155));
  or_6   g01779(.A(new_n2155), .B(new_n2142), .Y(new_n2156));
  xnor_4 g01780(.A(new_n2138), .B(new_n2137), .Y(new_n2157));
  xor_4  g01781(.A(new_n2155), .B(new_n2142), .Y(new_n2158));
  nand_5 g01782(.A(new_n2158), .B(new_n2157), .Y(new_n2159));
  nand_5 g01783(.A(new_n2159), .B(new_n2156), .Y(new_n2160));
  nand_5 g01784(.A(new_n2160), .B(new_n2141), .Y(new_n2161));
  nand_5 g01785(.A(pi116), .B(pi073), .Y(new_n2162));
  nand_5 g01786(.A(pi170), .B(pi115), .Y(new_n2163));
  xor_4  g01787(.A(new_n2163), .B(new_n2162), .Y(new_n2164));
  xor_4  g01788(.A(new_n2164), .B(new_n2116), .Y(new_n2165));
  nand_5 g01789(.A(pi039), .B(pi003), .Y(new_n2166));
  xor_4  g01790(.A(new_n2166), .B(new_n2118), .Y(new_n2167));
  not_8  g01791(.A(new_n2167), .Y(new_n2168));
  xor_4  g01792(.A(new_n2168), .B(new_n2165), .Y(new_n2169));
  nand_5 g01793(.A(pi148), .B(pi124), .Y(new_n2170));
  nand_5 g01794(.A(pi215), .B(pi163), .Y(new_n2171));
  xor_4  g01795(.A(new_n2171), .B(new_n2124), .Y(new_n2172));
  xor_4  g01796(.A(new_n2172), .B(new_n2170), .Y(new_n2173));
  nand_5 g01797(.A(new_n2111), .B(new_n2104), .Y(new_n2174));
  nand_5 g01798(.A(new_n2119), .B(new_n2112), .Y(new_n2175));
  nand_5 g01799(.A(new_n2175), .B(new_n2174), .Y(new_n2176));
  xor_4  g01800(.A(new_n2176), .B(new_n2173), .Y(new_n2177));
  xor_4  g01801(.A(new_n2177), .B(new_n2169), .Y(new_n2178));
  nor_5  g01802(.A(new_n2140), .B(new_n2128), .Y(new_n2179));
  nand_5 g01803(.A(new_n2179), .B(new_n2126), .Y(new_n2180));
  nor_5  g01804(.A(new_n2127), .B(new_n2120), .Y(new_n2181));
  or_6   g01805(.A(new_n2181), .B(new_n2126), .Y(new_n2182));
  or_6   g01806(.A(new_n2182), .B(new_n2179), .Y(new_n2183));
  nand_5 g01807(.A(new_n2183), .B(new_n2180), .Y(new_n2184));
  xor_4  g01808(.A(new_n2184), .B(new_n2178), .Y(new_n2185));
  xor_4  g01809(.A(new_n2185), .B(new_n2161), .Y(new_n2186));
  xnor_4 g01810(.A(new_n2160), .B(new_n2141), .Y(new_n2187));
  nand_5 g01811(.A(pi163), .B(pi124), .Y(new_n2188));
  or_6   g01812(.A(new_n2188), .B(new_n2187), .Y(new_n2189));
  xor_4  g01813(.A(new_n2153), .B(new_n2152), .Y(new_n2190));
  not_8  g01814(.A(new_n2146), .Y(new_n2191));
  not_8  g01815(.A(new_n2145), .Y(new_n2192));
  nand_5 g01816(.A(pi170), .B(pi163), .Y(new_n2193));
  nand_5 g01817(.A(new_n2193), .B(new_n2191), .Y(new_n2194));
  nand_5 g01818(.A(new_n2194), .B(new_n2192), .Y(new_n2195));
  nand_5 g01819(.A(new_n2195), .B(new_n2147), .Y(new_n2196));
  nand_5 g01820(.A(new_n2196), .B(new_n2191), .Y(new_n2197));
  nor_5  g01821(.A(new_n2197), .B(new_n2190), .Y(new_n2198));
  not_8  g01822(.A(new_n2198), .Y(new_n2199));
  xnor_4 g01823(.A(new_n2158), .B(new_n2157), .Y(new_n2200));
  nor_5  g01824(.A(new_n2200), .B(new_n2199), .Y(new_n2201));
  xor_4  g01825(.A(new_n2188), .B(new_n2187), .Y(new_n2202));
  nand_5 g01826(.A(new_n2202), .B(new_n2201), .Y(new_n2203));
  nand_5 g01827(.A(new_n2203), .B(new_n2189), .Y(new_n2204));
  xor_4  g01828(.A(new_n2204), .B(new_n2186), .Y(new_n2205));
  xor_4  g01829(.A(new_n2205), .B(new_n2103), .Y(new_n2206));
  xor_4  g01830(.A(new_n2075), .B(new_n2074), .Y(new_n2207));
  not_8  g01831(.A(new_n2207), .Y(new_n2208));
  xor_4  g01832(.A(new_n2202), .B(new_n2201), .Y(new_n2209));
  nand_5 g01833(.A(new_n2209), .B(new_n2208), .Y(new_n2210));
  not_8  g01834(.A(new_n2210), .Y(new_n2211));
  xnor_4 g01835(.A(new_n2044), .B(new_n2027), .Y(new_n2212));
  xnor_4 g01836(.A(new_n2026), .B(new_n2019), .Y(new_n2213));
  and_6  g01837(.A(new_n2023), .B(new_n2012), .Y(new_n2214));
  or_6   g01838(.A(new_n2214), .B(new_n2025), .Y(new_n2215));
  nor_5  g01839(.A(new_n2194), .B(new_n2192), .Y(new_n2216));
  nor_5  g01840(.A(new_n2216), .B(new_n2196), .Y(new_n2217));
  not_8  g01841(.A(new_n2217), .Y(new_n2218));
  nand_5 g01842(.A(new_n2218), .B(new_n2215), .Y(new_n2219));
  xor_4  g01843(.A(new_n2217), .B(new_n2215), .Y(new_n2220));
  nor_5  g01844(.A(new_n2193), .B(new_n2021), .Y(new_n2221));
  nand_5 g01845(.A(pi254), .B(pi171), .Y(new_n2222));
  nand_5 g01846(.A(pi158), .B(pi107), .Y(new_n2223));
  xor_4  g01847(.A(new_n2223), .B(new_n2222), .Y(new_n2224));
  nand_5 g01848(.A(new_n2224), .B(new_n2221), .Y(new_n2225));
  nand_5 g01849(.A(pi163), .B(pi004), .Y(new_n2226));
  nand_5 g01850(.A(pi170), .B(pi148), .Y(new_n2227));
  xor_4  g01851(.A(new_n2227), .B(new_n2226), .Y(new_n2228));
  xor_4  g01852(.A(new_n2224), .B(new_n2221), .Y(new_n2229));
  nand_5 g01853(.A(new_n2229), .B(new_n2228), .Y(new_n2230));
  nand_5 g01854(.A(new_n2230), .B(new_n2225), .Y(new_n2231));
  or_6   g01855(.A(new_n2231), .B(new_n2220), .Y(new_n2232));
  nand_5 g01856(.A(new_n2232), .B(new_n2219), .Y(new_n2233));
  nand_5 g01857(.A(new_n2233), .B(new_n2213), .Y(new_n2234));
  xor_4  g01858(.A(new_n2197), .B(new_n2190), .Y(new_n2235));
  not_8  g01859(.A(new_n2235), .Y(new_n2236));
  xor_4  g01860(.A(new_n2233), .B(new_n2213), .Y(new_n2237));
  nand_5 g01861(.A(new_n2237), .B(new_n2236), .Y(new_n2238));
  nand_5 g01862(.A(new_n2238), .B(new_n2234), .Y(new_n2239));
  nand_5 g01863(.A(new_n2239), .B(new_n2212), .Y(new_n2240));
  xor_4  g01864(.A(new_n2200), .B(new_n2198), .Y(new_n2241));
  xor_4  g01865(.A(new_n2239), .B(new_n2212), .Y(new_n2242));
  nand_5 g01866(.A(new_n2242), .B(new_n2241), .Y(new_n2243));
  nand_5 g01867(.A(new_n2243), .B(new_n2240), .Y(new_n2244));
  xor_4  g01868(.A(new_n2209), .B(new_n2207), .Y(new_n2245));
  nor_5  g01869(.A(new_n2245), .B(new_n2244), .Y(new_n2246));
  nor_5  g01870(.A(new_n2246), .B(new_n2211), .Y(new_n2247));
  xor_4  g01871(.A(new_n2247), .B(new_n2206), .Y(new_n2248));
  nand_5 g01872(.A(pi172), .B(pi134), .Y(new_n2249));
  nand_5 g01873(.A(pi240), .B(pi062), .Y(new_n2250));
  nand_5 g01874(.A(pi149), .B(pi065), .Y(new_n2251));
  nand_5 g01875(.A(new_n2251), .B(new_n2250), .Y(new_n2252));
  nand_5 g01876(.A(pi134), .B(pi120), .Y(new_n2253));
  xor_4  g01877(.A(new_n2251), .B(new_n2250), .Y(new_n2254));
  nand_5 g01878(.A(new_n2254), .B(new_n2253), .Y(new_n2255));
  nand_5 g01879(.A(new_n2255), .B(new_n2252), .Y(new_n2256));
  nand_5 g01880(.A(new_n2256), .B(new_n2249), .Y(new_n2257));
  nand_5 g01881(.A(pi167), .B(pi065), .Y(new_n2258));
  nand_5 g01882(.A(pi240), .B(pi120), .Y(new_n2259));
  nand_5 g01883(.A(pi149), .B(pi062), .Y(new_n2260));
  xor_4  g01884(.A(new_n2260), .B(new_n2259), .Y(new_n2261));
  xor_4  g01885(.A(new_n2261), .B(new_n2258), .Y(new_n2262));
  xor_4  g01886(.A(new_n2256), .B(new_n2249), .Y(new_n2263));
  nand_5 g01887(.A(new_n2263), .B(new_n2262), .Y(new_n2264));
  nand_5 g01888(.A(new_n2264), .B(new_n2257), .Y(new_n2265));
  nand_5 g01889(.A(pi149), .B(pi120), .Y(new_n2266));
  nand_5 g01890(.A(pi167), .B(pi062), .Y(new_n2267));
  nand_5 g01891(.A(pi181), .B(pi065), .Y(new_n2268));
  nand_5 g01892(.A(new_n2268), .B(new_n2267), .Y(new_n2269));
  nand_5 g01893(.A(pi181), .B(pi062), .Y(new_n2270));
  or_6   g01894(.A(new_n2270), .B(new_n2258), .Y(new_n2271));
  nand_5 g01895(.A(new_n2271), .B(new_n2269), .Y(new_n2272));
  xor_4  g01896(.A(new_n2272), .B(new_n2266), .Y(new_n2273));
  nand_5 g01897(.A(new_n2260), .B(new_n2259), .Y(new_n2274));
  nand_5 g01898(.A(new_n2261), .B(new_n2258), .Y(new_n2275));
  nand_5 g01899(.A(new_n2275), .B(new_n2274), .Y(new_n2276));
  xor_4  g01900(.A(new_n2276), .B(new_n2273), .Y(new_n2277));
  nand_5 g01901(.A(pi240), .B(pi172), .Y(new_n2278));
  nand_5 g01902(.A(pi198), .B(pi134), .Y(new_n2279));
  nand_5 g01903(.A(new_n2279), .B(new_n2278), .Y(new_n2280));
  nand_5 g01904(.A(pi240), .B(pi198), .Y(new_n2281));
  or_6   g01905(.A(new_n2281), .B(new_n2249), .Y(new_n2282));
  nand_5 g01906(.A(new_n2282), .B(new_n2280), .Y(new_n2283));
  xor_4  g01907(.A(new_n2283), .B(new_n2277), .Y(new_n2284));
  xor_4  g01908(.A(new_n2284), .B(new_n2265), .Y(new_n2285));
  xor_4  g01909(.A(new_n2263), .B(new_n2262), .Y(new_n2286));
  nand_5 g01910(.A(pi198), .B(pi175), .Y(new_n2287));
  or_6   g01911(.A(new_n2287), .B(new_n2286), .Y(new_n2288));
  xor_4  g01912(.A(new_n2287), .B(new_n2286), .Y(new_n2289));
  nand_5 g01913(.A(pi175), .B(pi120), .Y(new_n2290));
  nand_5 g01914(.A(pi240), .B(pi065), .Y(new_n2291));
  nand_5 g01915(.A(new_n2291), .B(new_n2290), .Y(new_n2292));
  nand_5 g01916(.A(pi134), .B(pi062), .Y(new_n2293));
  or_6   g01917(.A(new_n2291), .B(new_n2290), .Y(new_n2294));
  nand_5 g01918(.A(new_n2294), .B(new_n2293), .Y(new_n2295));
  nand_5 g01919(.A(new_n2295), .B(new_n2292), .Y(new_n2296));
  nand_5 g01920(.A(pi175), .B(pi172), .Y(new_n2297));
  or_6   g01921(.A(new_n2297), .B(new_n2296), .Y(new_n2298));
  xor_4  g01922(.A(new_n2297), .B(new_n2296), .Y(new_n2299));
  xnor_4 g01923(.A(new_n2254), .B(new_n2253), .Y(new_n2300));
  nand_5 g01924(.A(new_n2300), .B(new_n2299), .Y(new_n2301));
  nand_5 g01925(.A(new_n2301), .B(new_n2298), .Y(new_n2302));
  nand_5 g01926(.A(new_n2302), .B(new_n2289), .Y(new_n2303));
  nand_5 g01927(.A(new_n2303), .B(new_n2288), .Y(new_n2304));
  xor_4  g01928(.A(new_n2304), .B(new_n2285), .Y(new_n2305));
  xnor_4 g01929(.A(new_n2300), .B(new_n2299), .Y(new_n2306));
  not_8  g01930(.A(new_n2293), .Y(new_n2307));
  not_8  g01931(.A(new_n2292), .Y(new_n2308));
  nand_5 g01932(.A(pi175), .B(pi065), .Y(new_n2309));
  nand_5 g01933(.A(new_n2309), .B(new_n2307), .Y(new_n2310));
  nand_5 g01934(.A(new_n2310), .B(new_n2308), .Y(new_n2311));
  nand_5 g01935(.A(new_n2311), .B(new_n2294), .Y(new_n2312));
  nand_5 g01936(.A(new_n2312), .B(new_n2307), .Y(new_n2313));
  nor_5  g01937(.A(new_n2313), .B(new_n2306), .Y(new_n2314));
  xor_4  g01938(.A(new_n2302), .B(new_n2289), .Y(new_n2315));
  nand_5 g01939(.A(new_n2315), .B(new_n2314), .Y(new_n2316));
  nand_5 g01940(.A(pi175), .B(pi165), .Y(new_n2317));
  xor_4  g01941(.A(new_n2317), .B(new_n2316), .Y(new_n2318));
  xor_4  g01942(.A(new_n2318), .B(new_n2305), .Y(new_n2319));
  xor_4  g01943(.A(new_n2242), .B(new_n2241), .Y(new_n2320));
  xor_4  g01944(.A(new_n2315), .B(new_n2314), .Y(new_n2321));
  not_8  g01945(.A(new_n2321), .Y(new_n2322));
  nor_5  g01946(.A(new_n2322), .B(new_n2320), .Y(new_n2323));
  xor_4  g01947(.A(new_n2321), .B(new_n2320), .Y(new_n2324));
  xor_4  g01948(.A(new_n2237), .B(new_n2236), .Y(new_n2325));
  xor_4  g01949(.A(new_n2313), .B(new_n2306), .Y(new_n2326));
  not_8  g01950(.A(new_n2326), .Y(new_n2327));
  nand_5 g01951(.A(new_n2327), .B(new_n2325), .Y(new_n2328));
  xor_4  g01952(.A(new_n2327), .B(new_n2325), .Y(new_n2329));
  xor_4  g01953(.A(new_n2231), .B(new_n2220), .Y(new_n2330));
  nor_5  g01954(.A(new_n2310), .B(new_n2308), .Y(new_n2331));
  nor_5  g01955(.A(new_n2331), .B(new_n2312), .Y(new_n2332));
  not_8  g01956(.A(new_n2332), .Y(new_n2333));
  nor_5  g01957(.A(new_n2333), .B(new_n2330), .Y(new_n2334));
  xor_4  g01958(.A(new_n2332), .B(new_n2330), .Y(new_n2335));
  xor_4  g01959(.A(new_n2193), .B(new_n2021), .Y(new_n2336));
  not_8  g01960(.A(new_n2336), .Y(new_n2337));
  nor_5  g01961(.A(new_n2337), .B(new_n2309), .Y(new_n2338));
  nand_5 g01962(.A(pi175), .B(pi062), .Y(new_n2339));
  nand_5 g01963(.A(pi134), .B(pi065), .Y(new_n2340));
  xor_4  g01964(.A(new_n2340), .B(new_n2339), .Y(new_n2341));
  or_6   g01965(.A(new_n2341), .B(new_n2338), .Y(new_n2342));
  xor_4  g01966(.A(new_n2229), .B(new_n2228), .Y(new_n2343));
  not_8  g01967(.A(new_n2343), .Y(new_n2344));
  xor_4  g01968(.A(new_n2341), .B(new_n2338), .Y(new_n2345));
  nand_5 g01969(.A(new_n2345), .B(new_n2344), .Y(new_n2346));
  nand_5 g01970(.A(new_n2346), .B(new_n2342), .Y(new_n2347));
  nor_5  g01971(.A(new_n2347), .B(new_n2335), .Y(new_n2348));
  nor_5  g01972(.A(new_n2348), .B(new_n2334), .Y(new_n2349));
  nand_5 g01973(.A(new_n2349), .B(new_n2329), .Y(new_n2350));
  nand_5 g01974(.A(new_n2350), .B(new_n2328), .Y(new_n2351));
  nor_5  g01975(.A(new_n2351), .B(new_n2324), .Y(new_n2352));
  nor_5  g01976(.A(new_n2352), .B(new_n2323), .Y(new_n2353));
  nand_5 g01977(.A(new_n2353), .B(new_n2319), .Y(new_n2354));
  xnor_4 g01978(.A(new_n2245), .B(new_n2244), .Y(new_n2355));
  xor_4  g01979(.A(new_n2353), .B(new_n2319), .Y(new_n2356));
  nand_5 g01980(.A(new_n2356), .B(new_n2355), .Y(new_n2357));
  nand_5 g01981(.A(new_n2357), .B(new_n2354), .Y(new_n2358));
  nand_5 g01982(.A(new_n2358), .B(new_n2248), .Y(new_n2359));
  nand_5 g01983(.A(new_n2317), .B(new_n2316), .Y(new_n2360));
  nand_5 g01984(.A(new_n2318), .B(new_n2305), .Y(new_n2361));
  nand_5 g01985(.A(new_n2361), .B(new_n2360), .Y(new_n2362));
  not_8  g01986(.A(new_n2285), .Y(new_n2363));
  nand_5 g01987(.A(new_n2304), .B(new_n2363), .Y(new_n2364));
  nand_5 g01988(.A(pi200), .B(pi065), .Y(new_n2365));
  nand_5 g01989(.A(pi167), .B(pi120), .Y(new_n2366));
  xor_4  g01990(.A(new_n2366), .B(new_n2365), .Y(new_n2367));
  xor_4  g01991(.A(new_n2367), .B(new_n2270), .Y(new_n2368));
  not_8  g01992(.A(new_n2368), .Y(new_n2369));
  nand_5 g01993(.A(pi172), .B(pi149), .Y(new_n2370));
  xor_4  g01994(.A(new_n2370), .B(new_n2271), .Y(new_n2371));
  xor_4  g01995(.A(new_n2371), .B(new_n2369), .Y(new_n2372));
  nand_5 g01996(.A(pi165), .B(pi134), .Y(new_n2373));
  nand_5 g01997(.A(pi197), .B(pi175), .Y(new_n2374));
  xor_4  g01998(.A(new_n2374), .B(new_n2373), .Y(new_n2375));
  xor_4  g01999(.A(new_n2375), .B(new_n2281), .Y(new_n2376));
  nand_5 g02000(.A(new_n2272), .B(new_n2266), .Y(new_n2377));
  nand_5 g02001(.A(new_n2276), .B(new_n2273), .Y(new_n2378));
  nand_5 g02002(.A(new_n2378), .B(new_n2377), .Y(new_n2379));
  xor_4  g02003(.A(new_n2379), .B(new_n2376), .Y(new_n2380));
  xor_4  g02004(.A(new_n2380), .B(new_n2372), .Y(new_n2381));
  nand_5 g02005(.A(new_n2283), .B(new_n2277), .Y(new_n2382));
  nand_5 g02006(.A(new_n2284), .B(new_n2265), .Y(new_n2383));
  nand_5 g02007(.A(new_n2383), .B(new_n2382), .Y(new_n2384));
  xor_4  g02008(.A(new_n2384), .B(new_n2282), .Y(new_n2385));
  xnor_4 g02009(.A(new_n2385), .B(new_n2381), .Y(new_n2386));
  xor_4  g02010(.A(new_n2386), .B(new_n2364), .Y(new_n2387));
  xor_4  g02011(.A(new_n2387), .B(new_n2362), .Y(new_n2388));
  xor_4  g02012(.A(new_n2358), .B(new_n2248), .Y(new_n2389));
  nand_5 g02013(.A(new_n2389), .B(new_n2388), .Y(new_n2390));
  nand_5 g02014(.A(new_n2390), .B(new_n2359), .Y(new_n2391));
  nand_5 g02015(.A(pi234), .B(pi229), .Y(new_n2392));
  nand_5 g02016(.A(new_n1940), .B(new_n1939), .Y(new_n2393));
  nand_5 g02017(.A(new_n1941), .B(new_n1916), .Y(new_n2394));
  nand_5 g02018(.A(new_n2394), .B(new_n2393), .Y(new_n2395));
  xor_4  g02019(.A(new_n2395), .B(new_n2392), .Y(new_n2396));
  xor_4  g02020(.A(new_n2396), .B(new_n2391), .Y(new_n2397));
  nand_5 g02021(.A(new_n1947), .B(new_n1946), .Y(new_n2398));
  nand_5 g02022(.A(new_n1948), .B(new_n1902), .Y(new_n2399));
  nand_5 g02023(.A(new_n2399), .B(new_n2398), .Y(new_n2400));
  nand_5 g02024(.A(pi247), .B(pi067), .Y(new_n2401));
  nand_5 g02025(.A(pi080), .B(pi053), .Y(new_n2402));
  xor_4  g02026(.A(new_n2402), .B(new_n2401), .Y(new_n2403));
  xor_4  g02027(.A(new_n2403), .B(new_n2400), .Y(new_n2404));
  nand_5 g02028(.A(new_n2386), .B(new_n2364), .Y(new_n2405));
  nand_5 g02029(.A(new_n2387), .B(new_n2362), .Y(new_n2406));
  nand_5 g02030(.A(new_n2406), .B(new_n2405), .Y(new_n2407));
  nand_5 g02031(.A(pi214), .B(pi092), .Y(new_n2408));
  xor_4  g02032(.A(new_n2408), .B(new_n2407), .Y(new_n2409));
  xor_4  g02033(.A(new_n2409), .B(new_n2404), .Y(new_n2410));
  nand_5 g02034(.A(pi200), .B(pi062), .Y(new_n2411));
  nand_5 g02035(.A(pi203), .B(pi065), .Y(new_n2412));
  or_6   g02036(.A(new_n2384), .B(new_n2282), .Y(new_n2413));
  nand_5 g02037(.A(new_n2385), .B(new_n2381), .Y(new_n2414));
  nand_5 g02038(.A(new_n2414), .B(new_n2413), .Y(new_n2415));
  xnor_4 g02039(.A(new_n2415), .B(new_n2412), .Y(new_n2416));
  xor_4  g02040(.A(new_n2416), .B(new_n2411), .Y(new_n2417));
  nand_5 g02041(.A(pi175), .B(pi078), .Y(new_n2418));
  nand_5 g02042(.A(new_n1952), .B(new_n1949), .Y(new_n2419));
  nand_5 g02043(.A(new_n1953), .B(new_n1945), .Y(new_n2420));
  nand_5 g02044(.A(new_n2420), .B(new_n2419), .Y(new_n2421));
  xor_4  g02045(.A(new_n2421), .B(new_n2418), .Y(new_n2422));
  xor_4  g02046(.A(new_n2422), .B(new_n2417), .Y(new_n2423));
  nand_5 g02047(.A(pi117), .B(pi030), .Y(new_n2424));
  nand_5 g02048(.A(pi185), .B(pi016), .Y(new_n2425));
  or_6   g02049(.A(new_n1943), .B(new_n1917), .Y(new_n2426));
  not_8  g02050(.A(new_n1942), .Y(new_n2427));
  nand_5 g02051(.A(new_n1944), .B(new_n2427), .Y(new_n2428));
  nand_5 g02052(.A(new_n2428), .B(new_n2426), .Y(new_n2429));
  xor_4  g02053(.A(new_n2429), .B(new_n2425), .Y(new_n2430));
  xor_4  g02054(.A(new_n2430), .B(new_n2424), .Y(new_n2431));
  xor_4  g02055(.A(new_n2431), .B(new_n2423), .Y(new_n2432));
  xor_4  g02056(.A(new_n2432), .B(new_n2410), .Y(new_n2433));
  xor_4  g02057(.A(new_n2433), .B(new_n2397), .Y(new_n2434));
  nand_5 g02058(.A(pi197), .B(pi134), .Y(new_n2435));
  nand_5 g02059(.A(new_n2366), .B(new_n2365), .Y(new_n2436));
  nand_5 g02060(.A(new_n2367), .B(new_n2270), .Y(new_n2437));
  nand_5 g02061(.A(new_n2437), .B(new_n2436), .Y(new_n2438));
  xor_4  g02062(.A(new_n2438), .B(new_n2435), .Y(new_n2439));
  nand_5 g02063(.A(pi170), .B(pi000), .Y(new_n2440));
  nand_5 g02064(.A(pi115), .B(pi004), .Y(new_n2441));
  nand_5 g02065(.A(pi073), .B(pi070), .Y(new_n2442));
  xor_4  g02066(.A(new_n2442), .B(new_n2441), .Y(new_n2443));
  nand_5 g02067(.A(pi163), .B(pi022), .Y(new_n2444));
  nand_5 g02068(.A(new_n2379), .B(new_n2376), .Y(new_n2445));
  not_8  g02069(.A(new_n2372), .Y(new_n2446));
  nand_5 g02070(.A(new_n2380), .B(new_n2446), .Y(new_n2447));
  nand_5 g02071(.A(new_n2447), .B(new_n2445), .Y(new_n2448));
  xor_4  g02072(.A(new_n2448), .B(new_n2444), .Y(new_n2449));
  xor_4  g02073(.A(new_n2449), .B(new_n2443), .Y(new_n2450));
  xor_4  g02074(.A(new_n2450), .B(new_n2440), .Y(new_n2451));
  xor_4  g02075(.A(new_n2451), .B(new_n2439), .Y(new_n2452));
  xor_4  g02076(.A(new_n2452), .B(new_n2434), .Y(new_n2453));
  xor_4  g02077(.A(new_n2453), .B(new_n2003), .Y(new_n2454));
  nand_5 g02078(.A(pi202), .B(pi190), .Y(new_n2455));
  nand_5 g02079(.A(pi220), .B(pi103), .Y(new_n2456));
  xor_4  g02080(.A(new_n2456), .B(new_n2455), .Y(new_n2457));
  nand_5 g02081(.A(pi209), .B(pi171), .Y(new_n2458));
  nand_5 g02082(.A(new_n2094), .B(new_n2091), .Y(new_n2459));
  not_8  g02083(.A(new_n2087), .Y(new_n2460));
  nand_5 g02084(.A(new_n2095), .B(new_n2460), .Y(new_n2461));
  nand_5 g02085(.A(new_n2461), .B(new_n2459), .Y(new_n2462));
  xor_4  g02086(.A(new_n2462), .B(new_n2458), .Y(new_n2463));
  xor_4  g02087(.A(new_n2463), .B(new_n2457), .Y(new_n2464));
  nand_5 g02088(.A(new_n2176), .B(new_n2173), .Y(new_n2465));
  not_8  g02089(.A(new_n2169), .Y(new_n2466));
  nand_5 g02090(.A(new_n2177), .B(new_n2466), .Y(new_n2467));
  nand_5 g02091(.A(new_n2467), .B(new_n2465), .Y(new_n2468));
  nand_5 g02092(.A(new_n2101), .B(new_n2079), .Y(new_n2469));
  nand_5 g02093(.A(new_n2102), .B(new_n2077), .Y(new_n2470));
  nand_5 g02094(.A(new_n2470), .B(new_n2469), .Y(new_n2471));
  xor_4  g02095(.A(new_n2471), .B(new_n2468), .Y(new_n2472));
  nand_5 g02096(.A(new_n2171), .B(new_n2124), .Y(new_n2473));
  nand_5 g02097(.A(new_n2172), .B(new_n2170), .Y(new_n2474));
  nand_5 g02098(.A(new_n2474), .B(new_n2473), .Y(new_n2475));
  xor_4  g02099(.A(new_n2475), .B(new_n2472), .Y(new_n2476));
  nor_5  g02100(.A(new_n2166), .B(new_n2118), .Y(new_n2477));
  nor_5  g02101(.A(new_n2168), .B(new_n2165), .Y(new_n2478));
  or_6   g02102(.A(new_n2478), .B(new_n2477), .Y(new_n2479));
  nand_5 g02103(.A(new_n2163), .B(new_n2162), .Y(new_n2480));
  nand_5 g02104(.A(new_n2164), .B(new_n2116), .Y(new_n2481));
  nand_5 g02105(.A(new_n2481), .B(new_n2480), .Y(new_n2482));
  nand_5 g02106(.A(pi116), .B(pi003), .Y(new_n2483));
  xor_4  g02107(.A(new_n2483), .B(new_n2482), .Y(new_n2484));
  or_6   g02108(.A(new_n2099), .B(new_n2066), .Y(new_n2485));
  nand_5 g02109(.A(new_n2100), .B(new_n2096), .Y(new_n2486));
  nand_5 g02110(.A(new_n2486), .B(new_n2485), .Y(new_n2487));
  nand_5 g02111(.A(pi201), .B(pi154), .Y(new_n2488));
  nand_5 g02112(.A(pi245), .B(pi095), .Y(new_n2489));
  xor_4  g02113(.A(new_n2489), .B(new_n2488), .Y(new_n2490));
  xor_4  g02114(.A(new_n2490), .B(new_n2487), .Y(new_n2491));
  nand_5 g02115(.A(pi158), .B(pi063), .Y(new_n2492));
  nand_5 g02116(.A(pi153), .B(pi107), .Y(new_n2493));
  nand_5 g02117(.A(pi156), .B(pi089), .Y(new_n2494));
  nand_5 g02118(.A(pi254), .B(pi083), .Y(new_n2495));
  xor_4  g02119(.A(new_n2495), .B(new_n2494), .Y(new_n2496));
  xor_4  g02120(.A(new_n2496), .B(new_n2493), .Y(new_n2497));
  xor_4  g02121(.A(new_n2497), .B(new_n2492), .Y(new_n2498));
  xor_4  g02122(.A(new_n2498), .B(new_n2491), .Y(new_n2499));
  nand_5 g02123(.A(pi130), .B(pi039), .Y(new_n2500));
  nand_5 g02124(.A(pi228), .B(pi124), .Y(new_n2501));
  nand_5 g02125(.A(pi215), .B(pi148), .Y(new_n2502));
  xor_4  g02126(.A(new_n2502), .B(new_n2501), .Y(new_n2503));
  xor_4  g02127(.A(new_n2503), .B(new_n2500), .Y(new_n2504));
  xor_4  g02128(.A(new_n2504), .B(new_n2499), .Y(new_n2505));
  xor_4  g02129(.A(new_n2505), .B(new_n2484), .Y(new_n2506));
  xor_4  g02130(.A(new_n2506), .B(new_n2479), .Y(new_n2507));
  xor_4  g02131(.A(new_n2507), .B(new_n2476), .Y(new_n2508));
  nand_5 g02132(.A(new_n2081), .B(new_n2080), .Y(new_n2509));
  nand_5 g02133(.A(new_n2082), .B(new_n2054), .Y(new_n2510));
  nand_5 g02134(.A(new_n2510), .B(new_n2509), .Y(new_n2511));
  or_6   g02135(.A(new_n2085), .B(new_n2055), .Y(new_n2512));
  nand_5 g02136(.A(new_n2086), .B(new_n2084), .Y(new_n2513));
  nand_5 g02137(.A(new_n2513), .B(new_n2512), .Y(new_n2514));
  nand_5 g02138(.A(new_n2089), .B(new_n2088), .Y(new_n2515));
  nand_5 g02139(.A(new_n2090), .B(new_n2065), .Y(new_n2516));
  nand_5 g02140(.A(new_n2516), .B(new_n2515), .Y(new_n2517));
  nand_5 g02141(.A(pi049), .B(pi006), .Y(new_n2518));
  xor_4  g02142(.A(new_n2518), .B(new_n2517), .Y(new_n2519));
  xor_4  g02143(.A(new_n2519), .B(new_n2514), .Y(new_n2520));
  xor_4  g02144(.A(new_n2520), .B(new_n2511), .Y(new_n2521));
  xor_4  g02145(.A(new_n2521), .B(new_n2508), .Y(new_n2522));
  xor_4  g02146(.A(new_n2522), .B(new_n2464), .Y(new_n2523));
  nand_5 g02147(.A(pi181), .B(pi120), .Y(new_n2524));
  nand_5 g02148(.A(new_n2374), .B(new_n2373), .Y(new_n2525));
  nand_5 g02149(.A(new_n2375), .B(new_n2281), .Y(new_n2526));
  nand_5 g02150(.A(new_n2526), .B(new_n2525), .Y(new_n2527));
  or_6   g02151(.A(new_n2184), .B(new_n2178), .Y(new_n2528));
  nand_5 g02152(.A(new_n2528), .B(new_n2183), .Y(new_n2529));
  xor_4  g02153(.A(new_n2529), .B(new_n2527), .Y(new_n2530));
  or_6   g02154(.A(new_n2185), .B(new_n2161), .Y(new_n2531));
  nand_5 g02155(.A(new_n2204), .B(new_n2186), .Y(new_n2532));
  nand_5 g02156(.A(new_n2532), .B(new_n2531), .Y(new_n2533));
  xor_4  g02157(.A(new_n2533), .B(new_n2530), .Y(new_n2534));
  xor_4  g02158(.A(new_n2534), .B(new_n2524), .Y(new_n2535));
  xor_4  g02159(.A(new_n2000), .B(new_n1999), .Y(new_n2536));
  xor_4  g02160(.A(new_n2389), .B(new_n2388), .Y(new_n2537));
  or_6   g02161(.A(new_n2537), .B(new_n2536), .Y(new_n2538));
  xor_4  g02162(.A(new_n2537), .B(new_n2536), .Y(new_n2539));
  xor_4  g02163(.A(new_n2356), .B(new_n2355), .Y(new_n2540));
  xor_4  g02164(.A(new_n1997), .B(new_n1996), .Y(new_n2541));
  or_6   g02165(.A(new_n2541), .B(new_n2540), .Y(new_n2542));
  xor_4  g02166(.A(new_n2541), .B(new_n2540), .Y(new_n2543));
  xor_4  g02167(.A(new_n2351), .B(new_n2324), .Y(new_n2544));
  xor_4  g02168(.A(new_n1992), .B(new_n1991), .Y(new_n2545));
  nand_5 g02169(.A(new_n2545), .B(new_n2544), .Y(new_n2546));
  xor_4  g02170(.A(new_n2545), .B(new_n2544), .Y(new_n2547));
  xnor_4 g02171(.A(new_n2349), .B(new_n2329), .Y(new_n2548));
  xor_4  g02172(.A(new_n1990), .B(new_n1989), .Y(new_n2549));
  nor_5  g02173(.A(new_n2549), .B(new_n2548), .Y(new_n2550));
  xor_4  g02174(.A(new_n2549), .B(new_n2548), .Y(new_n2551));
  not_8  g02175(.A(new_n2551), .Y(new_n2552));
  xor_4  g02176(.A(new_n1988), .B(new_n1985), .Y(new_n2553));
  xor_4  g02177(.A(new_n2336), .B(new_n2309), .Y(new_n2554));
  or_6   g02178(.A(new_n2554), .B(new_n1986), .Y(new_n2555));
  nand_5 g02179(.A(pi103), .B(pi092), .Y(new_n2556));
  nand_5 g02180(.A(pi190), .B(pi117), .Y(new_n2557));
  nand_5 g02181(.A(new_n2557), .B(new_n2556), .Y(new_n2558));
  nand_5 g02182(.A(new_n2558), .B(new_n1988), .Y(new_n2559));
  or_6   g02183(.A(new_n2559), .B(new_n2555), .Y(new_n2560));
  xor_4  g02184(.A(new_n2345), .B(new_n2343), .Y(new_n2561));
  xor_4  g02185(.A(new_n2559), .B(new_n2555), .Y(new_n2562));
  nand_5 g02186(.A(new_n2562), .B(new_n2561), .Y(new_n2563));
  nand_5 g02187(.A(new_n2563), .B(new_n2560), .Y(new_n2564));
  nand_5 g02188(.A(new_n2564), .B(new_n2553), .Y(new_n2565));
  xor_4  g02189(.A(new_n2347), .B(new_n2335), .Y(new_n2566));
  xor_4  g02190(.A(new_n2564), .B(new_n2553), .Y(new_n2567));
  nand_5 g02191(.A(new_n2567), .B(new_n2566), .Y(new_n2568));
  nand_5 g02192(.A(new_n2568), .B(new_n2565), .Y(new_n2569));
  nor_5  g02193(.A(new_n2569), .B(new_n2552), .Y(new_n2570));
  nor_5  g02194(.A(new_n2570), .B(new_n2550), .Y(new_n2571));
  nand_5 g02195(.A(new_n2571), .B(new_n2547), .Y(new_n2572));
  nand_5 g02196(.A(new_n2572), .B(new_n2546), .Y(new_n2573));
  nand_5 g02197(.A(new_n2573), .B(new_n2543), .Y(new_n2574));
  nand_5 g02198(.A(new_n2574), .B(new_n2542), .Y(new_n2575));
  nand_5 g02199(.A(new_n2575), .B(new_n2539), .Y(new_n2576));
  nand_5 g02200(.A(new_n2576), .B(new_n2538), .Y(new_n2577));
  or_6   g02201(.A(new_n2370), .B(new_n2271), .Y(new_n2578));
  nand_5 g02202(.A(new_n2371), .B(new_n2369), .Y(new_n2579));
  nand_5 g02203(.A(new_n2579), .B(new_n2578), .Y(new_n2580));
  nand_5 g02204(.A(pi198), .B(pi149), .Y(new_n2581));
  nand_5 g02205(.A(pi240), .B(pi165), .Y(new_n2582));
  xor_4  g02206(.A(new_n2582), .B(new_n2581), .Y(new_n2583));
  xor_4  g02207(.A(new_n2583), .B(new_n2580), .Y(new_n2584));
  xor_4  g02208(.A(new_n2584), .B(new_n2577), .Y(new_n2585));
  xor_4  g02209(.A(new_n2585), .B(new_n2535), .Y(new_n2586));
  nand_5 g02210(.A(new_n2205), .B(new_n2103), .Y(new_n2587));
  not_8  g02211(.A(new_n2247), .Y(new_n2588));
  nand_5 g02212(.A(new_n2588), .B(new_n2206), .Y(new_n2589));
  nand_5 g02213(.A(new_n2589), .B(new_n2587), .Y(new_n2590));
  nand_5 g02214(.A(pi172), .B(pi167), .Y(new_n2591));
  xor_4  g02215(.A(new_n2591), .B(new_n2590), .Y(new_n2592));
  xor_4  g02216(.A(new_n2592), .B(new_n2586), .Y(new_n2593));
  xor_4  g02217(.A(new_n2593), .B(new_n2523), .Y(new_n2594));
  xor_4  g02218(.A(new_n2594), .B(new_n2454), .Y(po006));
  nand_5 g02219(.A(pi216), .B(pi120), .Y(new_n2596));
  nand_5 g02220(.A(pi076), .B(pi062), .Y(new_n2597));
  nand_5 g02221(.A(pi079), .B(pi065), .Y(new_n2598));
  nand_5 g02222(.A(new_n2598), .B(new_n2597), .Y(new_n2599));
  nand_5 g02223(.A(pi076), .B(pi065), .Y(new_n2600));
  nand_5 g02224(.A(pi079), .B(pi062), .Y(new_n2601));
  or_6   g02225(.A(new_n2601), .B(new_n2600), .Y(new_n2602));
  nand_5 g02226(.A(new_n2602), .B(new_n2599), .Y(new_n2603));
  xor_4  g02227(.A(new_n2603), .B(new_n2596), .Y(new_n2604));
  nand_5 g02228(.A(pi120), .B(pi041), .Y(new_n2605));
  nand_5 g02229(.A(new_n2605), .B(new_n2600), .Y(new_n2606));
  nand_5 g02230(.A(pi216), .B(pi062), .Y(new_n2607));
  xor_4  g02231(.A(new_n2605), .B(new_n2600), .Y(new_n2608));
  nand_5 g02232(.A(new_n2608), .B(new_n2607), .Y(new_n2609));
  nand_5 g02233(.A(new_n2609), .B(new_n2606), .Y(new_n2610));
  xor_4  g02234(.A(new_n2610), .B(new_n2604), .Y(new_n2611));
  nand_5 g02235(.A(pi172), .B(pi041), .Y(new_n2612));
  nand_5 g02236(.A(pi198), .B(pi182), .Y(new_n2613));
  and_6  g02237(.A(new_n2613), .B(new_n2612), .Y(new_n2614));
  nand_5 g02238(.A(pi182), .B(pi172), .Y(new_n2615));
  nand_5 g02239(.A(pi198), .B(pi041), .Y(new_n2616));
  nor_5  g02240(.A(new_n2616), .B(new_n2615), .Y(new_n2617));
  or_6   g02241(.A(new_n2617), .B(new_n2614), .Y(new_n2618));
  xnor_4 g02242(.A(new_n2618), .B(new_n2611), .Y(new_n2619));
  nand_5 g02243(.A(pi062), .B(pi041), .Y(new_n2620));
  nand_5 g02244(.A(pi216), .B(pi065), .Y(new_n2621));
  nand_5 g02245(.A(new_n2621), .B(new_n2620), .Y(new_n2622));
  nand_5 g02246(.A(pi182), .B(pi120), .Y(new_n2623));
  xor_4  g02247(.A(new_n2621), .B(new_n2620), .Y(new_n2624));
  nand_5 g02248(.A(new_n2624), .B(new_n2623), .Y(new_n2625));
  nand_5 g02249(.A(new_n2625), .B(new_n2622), .Y(new_n2626));
  nand_5 g02250(.A(new_n2626), .B(new_n2615), .Y(new_n2627));
  xor_4  g02251(.A(new_n2608), .B(new_n2607), .Y(new_n2628));
  xor_4  g02252(.A(new_n2626), .B(new_n2615), .Y(new_n2629));
  nand_5 g02253(.A(new_n2629), .B(new_n2628), .Y(new_n2630));
  nand_5 g02254(.A(new_n2630), .B(new_n2627), .Y(new_n2631));
  xor_4  g02255(.A(new_n2631), .B(new_n2619), .Y(new_n2632));
  xor_4  g02256(.A(new_n2629), .B(new_n2628), .Y(new_n2633));
  nand_5 g02257(.A(pi198), .B(pi138), .Y(new_n2634));
  or_6   g02258(.A(new_n2634), .B(new_n2633), .Y(new_n2635));
  xor_4  g02259(.A(new_n2634), .B(new_n2633), .Y(new_n2636));
  nand_5 g02260(.A(pi172), .B(pi138), .Y(new_n2637));
  nand_5 g02261(.A(pi182), .B(pi062), .Y(new_n2638));
  nand_5 g02262(.A(pi138), .B(pi120), .Y(new_n2639));
  nand_5 g02263(.A(new_n2639), .B(new_n2638), .Y(new_n2640));
  nand_5 g02264(.A(pi065), .B(pi041), .Y(new_n2641));
  xor_4  g02265(.A(new_n2639), .B(new_n2638), .Y(new_n2642));
  nand_5 g02266(.A(new_n2642), .B(new_n2641), .Y(new_n2643));
  nand_5 g02267(.A(new_n2643), .B(new_n2640), .Y(new_n2644));
  or_6   g02268(.A(new_n2644), .B(new_n2637), .Y(new_n2645));
  xnor_4 g02269(.A(new_n2624), .B(new_n2623), .Y(new_n2646));
  xor_4  g02270(.A(new_n2644), .B(new_n2637), .Y(new_n2647));
  nand_5 g02271(.A(new_n2647), .B(new_n2646), .Y(new_n2648));
  nand_5 g02272(.A(new_n2648), .B(new_n2645), .Y(new_n2649));
  nand_5 g02273(.A(new_n2649), .B(new_n2636), .Y(new_n2650));
  nand_5 g02274(.A(new_n2650), .B(new_n2635), .Y(new_n2651));
  nand_5 g02275(.A(new_n2651), .B(new_n2632), .Y(new_n2652));
  nand_5 g02276(.A(pi120), .B(pi076), .Y(new_n2653));
  nand_5 g02277(.A(pi251), .B(pi065), .Y(new_n2654));
  xor_4  g02278(.A(new_n2654), .B(new_n2653), .Y(new_n2655));
  xor_4  g02279(.A(new_n2655), .B(new_n2601), .Y(new_n2656));
  not_8  g02280(.A(new_n2656), .Y(new_n2657));
  nand_5 g02281(.A(pi216), .B(pi172), .Y(new_n2658));
  xor_4  g02282(.A(new_n2658), .B(new_n2602), .Y(new_n2659));
  xor_4  g02283(.A(new_n2659), .B(new_n2657), .Y(new_n2660));
  nand_5 g02284(.A(pi197), .B(pi138), .Y(new_n2661));
  nand_5 g02285(.A(pi182), .B(pi165), .Y(new_n2662));
  xor_4  g02286(.A(new_n2662), .B(new_n2661), .Y(new_n2663));
  xor_4  g02287(.A(new_n2663), .B(new_n2616), .Y(new_n2664));
  nand_5 g02288(.A(new_n2603), .B(new_n2596), .Y(new_n2665));
  nand_5 g02289(.A(new_n2610), .B(new_n2604), .Y(new_n2666));
  nand_5 g02290(.A(new_n2666), .B(new_n2665), .Y(new_n2667));
  xor_4  g02291(.A(new_n2667), .B(new_n2664), .Y(new_n2668));
  xor_4  g02292(.A(new_n2668), .B(new_n2660), .Y(new_n2669));
  nor_5  g02293(.A(new_n2631), .B(new_n2619), .Y(new_n2670));
  nand_5 g02294(.A(new_n2670), .B(new_n2617), .Y(new_n2671));
  nor_5  g02295(.A(new_n2618), .B(new_n2611), .Y(new_n2672));
  or_6   g02296(.A(new_n2672), .B(new_n2617), .Y(new_n2673));
  or_6   g02297(.A(new_n2673), .B(new_n2670), .Y(new_n2674));
  nand_5 g02298(.A(new_n2674), .B(new_n2671), .Y(new_n2675));
  xor_4  g02299(.A(new_n2675), .B(new_n2669), .Y(new_n2676));
  xnor_4 g02300(.A(new_n2676), .B(new_n2652), .Y(new_n2677));
  nand_5 g02301(.A(pi165), .B(pi138), .Y(new_n2678));
  xor_4  g02302(.A(new_n2642), .B(new_n2641), .Y(new_n2679));
  nand_5 g02303(.A(pi138), .B(pi065), .Y(new_n2680));
  nor_5  g02304(.A(new_n2680), .B(new_n2638), .Y(new_n2681));
  not_8  g02305(.A(new_n2681), .Y(new_n2682));
  or_6   g02306(.A(new_n2682), .B(new_n2679), .Y(new_n2683));
  xnor_4 g02307(.A(new_n2647), .B(new_n2646), .Y(new_n2684));
  nor_5  g02308(.A(new_n2684), .B(new_n2683), .Y(new_n2685));
  xor_4  g02309(.A(new_n2649), .B(new_n2636), .Y(new_n2686));
  nand_5 g02310(.A(new_n2686), .B(new_n2685), .Y(new_n2687));
  nand_5 g02311(.A(new_n2687), .B(new_n2678), .Y(new_n2688));
  xnor_4 g02312(.A(new_n2651), .B(new_n2632), .Y(new_n2689));
  xor_4  g02313(.A(new_n2687), .B(new_n2678), .Y(new_n2690));
  nand_5 g02314(.A(new_n2690), .B(new_n2689), .Y(new_n2691));
  nand_5 g02315(.A(new_n2691), .B(new_n2688), .Y(new_n2692));
  xor_4  g02316(.A(new_n2692), .B(new_n2677), .Y(new_n2693));
  nand_5 g02317(.A(pi089), .B(pi001), .Y(new_n2694));
  nand_5 g02318(.A(pi158), .B(pi001), .Y(new_n2695));
  nand_5 g02319(.A(pi254), .B(pi122), .Y(new_n2696));
  nand_5 g02320(.A(new_n2696), .B(new_n2695), .Y(new_n2697));
  nand_5 g02321(.A(pi102), .B(pi089), .Y(new_n2698));
  xor_4  g02322(.A(new_n2696), .B(new_n2695), .Y(new_n2699));
  nand_5 g02323(.A(new_n2699), .B(new_n2698), .Y(new_n2700));
  nand_5 g02324(.A(new_n2700), .B(new_n2697), .Y(new_n2701));
  xor_4  g02325(.A(new_n2701), .B(new_n2694), .Y(new_n2702));
  nand_5 g02326(.A(pi158), .B(pi122), .Y(new_n2703));
  nand_5 g02327(.A(pi254), .B(pi135), .Y(new_n2704));
  nand_5 g02328(.A(new_n2704), .B(new_n2703), .Y(new_n2705));
  nand_5 g02329(.A(pi158), .B(pi135), .Y(new_n2706));
  nor_5  g02330(.A(new_n2706), .B(new_n2696), .Y(new_n2707));
  not_8  g02331(.A(new_n2707), .Y(new_n2708));
  nand_5 g02332(.A(new_n2708), .B(new_n2705), .Y(new_n2709));
  xor_4  g02333(.A(new_n2709), .B(new_n2702), .Y(new_n2710));
  nand_5 g02334(.A(pi219), .B(pi095), .Y(new_n2711));
  nand_5 g02335(.A(pi154), .B(pi102), .Y(new_n2712));
  and_6  g02336(.A(new_n2712), .B(new_n2711), .Y(new_n2713));
  nand_5 g02337(.A(pi219), .B(pi154), .Y(new_n2714));
  nand_5 g02338(.A(pi102), .B(pi095), .Y(new_n2715));
  nor_5  g02339(.A(new_n2715), .B(new_n2714), .Y(new_n2716));
  or_6   g02340(.A(new_n2716), .B(new_n2713), .Y(new_n2717));
  xnor_4 g02341(.A(new_n2717), .B(new_n2710), .Y(new_n2718));
  nand_5 g02342(.A(pi158), .B(pi102), .Y(new_n2719));
  nand_5 g02343(.A(pi219), .B(pi089), .Y(new_n2720));
  nand_5 g02344(.A(new_n2720), .B(new_n2719), .Y(new_n2721));
  nand_5 g02345(.A(pi254), .B(pi001), .Y(new_n2722));
  xor_4  g02346(.A(new_n2720), .B(new_n2719), .Y(new_n2723));
  nand_5 g02347(.A(new_n2723), .B(new_n2722), .Y(new_n2724));
  nand_5 g02348(.A(new_n2724), .B(new_n2721), .Y(new_n2725));
  nand_5 g02349(.A(new_n2725), .B(new_n2714), .Y(new_n2726));
  xor_4  g02350(.A(new_n2699), .B(new_n2698), .Y(new_n2727));
  xor_4  g02351(.A(new_n2725), .B(new_n2714), .Y(new_n2728));
  nand_5 g02352(.A(new_n2728), .B(new_n2727), .Y(new_n2729));
  nand_5 g02353(.A(new_n2729), .B(new_n2726), .Y(new_n2730));
  xor_4  g02354(.A(new_n2730), .B(new_n2718), .Y(new_n2731));
  xor_4  g02355(.A(new_n2728), .B(new_n2727), .Y(new_n2732));
  nand_5 g02356(.A(pi095), .B(pi087), .Y(new_n2733));
  or_6   g02357(.A(new_n2733), .B(new_n2732), .Y(new_n2734));
  xor_4  g02358(.A(new_n2733), .B(new_n2732), .Y(new_n2735));
  nand_5 g02359(.A(pi254), .B(pi102), .Y(new_n2736));
  nand_5 g02360(.A(pi089), .B(pi087), .Y(new_n2737));
  nand_5 g02361(.A(new_n2737), .B(new_n2736), .Y(new_n2738));
  nand_5 g02362(.A(pi219), .B(pi158), .Y(new_n2739));
  or_6   g02363(.A(new_n2737), .B(new_n2736), .Y(new_n2740));
  nand_5 g02364(.A(new_n2740), .B(new_n2739), .Y(new_n2741));
  nand_5 g02365(.A(new_n2741), .B(new_n2738), .Y(new_n2742));
  nand_5 g02366(.A(pi154), .B(pi087), .Y(new_n2743));
  or_6   g02367(.A(new_n2743), .B(new_n2742), .Y(new_n2744));
  xor_4  g02368(.A(new_n2743), .B(new_n2742), .Y(new_n2745));
  xnor_4 g02369(.A(new_n2723), .B(new_n2722), .Y(new_n2746));
  nand_5 g02370(.A(new_n2746), .B(new_n2745), .Y(new_n2747));
  nand_5 g02371(.A(new_n2747), .B(new_n2744), .Y(new_n2748));
  nand_5 g02372(.A(new_n2748), .B(new_n2735), .Y(new_n2749));
  nand_5 g02373(.A(new_n2749), .B(new_n2734), .Y(new_n2750));
  nand_5 g02374(.A(new_n2750), .B(new_n2731), .Y(new_n2751));
  nand_5 g02375(.A(pi122), .B(pi089), .Y(new_n2752));
  nand_5 g02376(.A(pi254), .B(pi059), .Y(new_n2753));
  xor_4  g02377(.A(new_n2753), .B(new_n2752), .Y(new_n2754));
  xor_4  g02378(.A(new_n2754), .B(new_n2706), .Y(new_n2755));
  nand_5 g02379(.A(pi154), .B(pi001), .Y(new_n2756));
  xor_4  g02380(.A(new_n2756), .B(new_n2708), .Y(new_n2757));
  not_8  g02381(.A(new_n2757), .Y(new_n2758));
  xor_4  g02382(.A(new_n2758), .B(new_n2755), .Y(new_n2759));
  nand_5 g02383(.A(pi209), .B(pi087), .Y(new_n2760));
  nand_5 g02384(.A(pi219), .B(pi006), .Y(new_n2761));
  xor_4  g02385(.A(new_n2761), .B(new_n2715), .Y(new_n2762));
  xor_4  g02386(.A(new_n2762), .B(new_n2760), .Y(new_n2763));
  nand_5 g02387(.A(new_n2701), .B(new_n2694), .Y(new_n2764));
  nand_5 g02388(.A(new_n2709), .B(new_n2702), .Y(new_n2765));
  nand_5 g02389(.A(new_n2765), .B(new_n2764), .Y(new_n2766));
  xor_4  g02390(.A(new_n2766), .B(new_n2763), .Y(new_n2767));
  xor_4  g02391(.A(new_n2767), .B(new_n2759), .Y(new_n2768));
  nor_5  g02392(.A(new_n2730), .B(new_n2718), .Y(new_n2769));
  nand_5 g02393(.A(new_n2769), .B(new_n2716), .Y(new_n2770));
  nor_5  g02394(.A(new_n2717), .B(new_n2710), .Y(new_n2771));
  or_6   g02395(.A(new_n2771), .B(new_n2716), .Y(new_n2772));
  or_6   g02396(.A(new_n2772), .B(new_n2769), .Y(new_n2773));
  nand_5 g02397(.A(new_n2773), .B(new_n2770), .Y(new_n2774));
  xor_4  g02398(.A(new_n2774), .B(new_n2768), .Y(new_n2775));
  xnor_4 g02399(.A(new_n2775), .B(new_n2751), .Y(new_n2776));
  xnor_4 g02400(.A(new_n2746), .B(new_n2745), .Y(new_n2777));
  not_8  g02401(.A(new_n2739), .Y(new_n2778));
  not_8  g02402(.A(new_n2738), .Y(new_n2779));
  nand_5 g02403(.A(pi254), .B(pi087), .Y(new_n2780));
  nand_5 g02404(.A(new_n2780), .B(new_n2778), .Y(new_n2781));
  nand_5 g02405(.A(new_n2781), .B(new_n2779), .Y(new_n2782));
  nand_5 g02406(.A(new_n2782), .B(new_n2740), .Y(new_n2783));
  nand_5 g02407(.A(new_n2783), .B(new_n2778), .Y(new_n2784));
  nor_5  g02408(.A(new_n2784), .B(new_n2777), .Y(new_n2785));
  xor_4  g02409(.A(new_n2748), .B(new_n2735), .Y(new_n2786));
  nand_5 g02410(.A(new_n2786), .B(new_n2785), .Y(new_n2787));
  nand_5 g02411(.A(pi087), .B(pi006), .Y(new_n2788));
  nand_5 g02412(.A(new_n2788), .B(new_n2787), .Y(new_n2789));
  xnor_4 g02413(.A(new_n2750), .B(new_n2731), .Y(new_n2790));
  xor_4  g02414(.A(new_n2788), .B(new_n2787), .Y(new_n2791));
  nand_5 g02415(.A(new_n2791), .B(new_n2790), .Y(new_n2792));
  nand_5 g02416(.A(new_n2792), .B(new_n2789), .Y(new_n2793));
  xor_4  g02417(.A(new_n2793), .B(new_n2776), .Y(new_n2794));
  nand_5 g02418(.A(pi071), .B(pi003), .Y(new_n2795));
  nand_5 g02419(.A(pi169), .B(pi004), .Y(new_n2796));
  nand_5 g02420(.A(pi073), .B(pi071), .Y(new_n2797));
  nand_5 g02421(.A(new_n2797), .B(new_n2796), .Y(new_n2798));
  nand_5 g02422(.A(pi170), .B(pi123), .Y(new_n2799));
  xor_4  g02423(.A(new_n2797), .B(new_n2796), .Y(new_n2800));
  nand_5 g02424(.A(new_n2800), .B(new_n2799), .Y(new_n2801));
  nand_5 g02425(.A(new_n2801), .B(new_n2798), .Y(new_n2802));
  nand_5 g02426(.A(new_n2802), .B(new_n2795), .Y(new_n2803));
  nand_5 g02427(.A(pi170), .B(pi099), .Y(new_n2804));
  nand_5 g02428(.A(pi169), .B(pi073), .Y(new_n2805));
  nand_5 g02429(.A(pi123), .B(pi004), .Y(new_n2806));
  xor_4  g02430(.A(new_n2806), .B(new_n2805), .Y(new_n2807));
  xor_4  g02431(.A(new_n2807), .B(new_n2804), .Y(new_n2808));
  xor_4  g02432(.A(new_n2802), .B(new_n2795), .Y(new_n2809));
  nand_5 g02433(.A(new_n2809), .B(new_n2808), .Y(new_n2810));
  nand_5 g02434(.A(new_n2810), .B(new_n2803), .Y(new_n2811));
  nand_5 g02435(.A(pi123), .B(pi073), .Y(new_n2812));
  nand_5 g02436(.A(new_n2806), .B(new_n2805), .Y(new_n2813));
  nand_5 g02437(.A(new_n2807), .B(new_n2804), .Y(new_n2814));
  nand_5 g02438(.A(new_n2814), .B(new_n2813), .Y(new_n2815));
  xor_4  g02439(.A(new_n2815), .B(new_n2812), .Y(new_n2816));
  nand_5 g02440(.A(pi099), .B(pi004), .Y(new_n2817));
  nand_5 g02441(.A(pi170), .B(pi023), .Y(new_n2818));
  nand_5 g02442(.A(new_n2818), .B(new_n2817), .Y(new_n2819));
  nand_5 g02443(.A(pi023), .B(pi004), .Y(new_n2820));
  nor_5  g02444(.A(new_n2820), .B(new_n2804), .Y(new_n2821));
  not_8  g02445(.A(new_n2821), .Y(new_n2822));
  nand_5 g02446(.A(new_n2822), .B(new_n2819), .Y(new_n2823));
  xor_4  g02447(.A(new_n2823), .B(new_n2816), .Y(new_n2824));
  nand_5 g02448(.A(pi130), .B(pi071), .Y(new_n2825));
  nand_5 g02449(.A(pi169), .B(pi003), .Y(new_n2826));
  nand_5 g02450(.A(new_n2826), .B(new_n2825), .Y(new_n2827));
  nand_5 g02451(.A(pi169), .B(pi130), .Y(new_n2828));
  or_6   g02452(.A(new_n2828), .B(new_n2795), .Y(new_n2829));
  nand_5 g02453(.A(new_n2829), .B(new_n2827), .Y(new_n2830));
  xor_4  g02454(.A(new_n2830), .B(new_n2824), .Y(new_n2831));
  xnor_4 g02455(.A(new_n2831), .B(new_n2811), .Y(new_n2832));
  xor_4  g02456(.A(new_n2809), .B(new_n2808), .Y(new_n2833));
  nand_5 g02457(.A(pi142), .B(pi130), .Y(new_n2834));
  or_6   g02458(.A(new_n2834), .B(new_n2833), .Y(new_n2835));
  xor_4  g02459(.A(new_n2834), .B(new_n2833), .Y(new_n2836));
  nand_5 g02460(.A(pi170), .B(pi169), .Y(new_n2837));
  nand_5 g02461(.A(pi142), .B(pi073), .Y(new_n2838));
  nand_5 g02462(.A(new_n2838), .B(new_n2837), .Y(new_n2839));
  nand_5 g02463(.A(pi071), .B(pi004), .Y(new_n2840));
  or_6   g02464(.A(new_n2838), .B(new_n2837), .Y(new_n2841));
  nand_5 g02465(.A(new_n2841), .B(new_n2840), .Y(new_n2842));
  nand_5 g02466(.A(new_n2842), .B(new_n2839), .Y(new_n2843));
  nand_5 g02467(.A(pi142), .B(pi003), .Y(new_n2844));
  or_6   g02468(.A(new_n2844), .B(new_n2843), .Y(new_n2845));
  xor_4  g02469(.A(new_n2844), .B(new_n2843), .Y(new_n2846));
  xnor_4 g02470(.A(new_n2800), .B(new_n2799), .Y(new_n2847));
  nand_5 g02471(.A(new_n2847), .B(new_n2846), .Y(new_n2848));
  nand_5 g02472(.A(new_n2848), .B(new_n2845), .Y(new_n2849));
  nand_5 g02473(.A(new_n2849), .B(new_n2836), .Y(new_n2850));
  nand_5 g02474(.A(new_n2850), .B(new_n2835), .Y(new_n2851));
  nand_5 g02475(.A(new_n2851), .B(new_n2832), .Y(new_n2852));
  nand_5 g02476(.A(pi099), .B(pi073), .Y(new_n2853));
  nand_5 g02477(.A(pi170), .B(pi155), .Y(new_n2854));
  xor_4  g02478(.A(new_n2854), .B(new_n2853), .Y(new_n2855));
  xor_4  g02479(.A(new_n2855), .B(new_n2820), .Y(new_n2856));
  nand_5 g02480(.A(pi123), .B(pi003), .Y(new_n2857));
  xor_4  g02481(.A(new_n2857), .B(new_n2822), .Y(new_n2858));
  not_8  g02482(.A(new_n2858), .Y(new_n2859));
  xor_4  g02483(.A(new_n2859), .B(new_n2856), .Y(new_n2860));
  nand_5 g02484(.A(pi215), .B(pi142), .Y(new_n2861));
  nand_5 g02485(.A(pi124), .B(pi071), .Y(new_n2862));
  xor_4  g02486(.A(new_n2862), .B(new_n2861), .Y(new_n2863));
  xor_4  g02487(.A(new_n2863), .B(new_n2828), .Y(new_n2864));
  nand_5 g02488(.A(new_n2815), .B(new_n2812), .Y(new_n2865));
  nand_5 g02489(.A(new_n2823), .B(new_n2816), .Y(new_n2866));
  nand_5 g02490(.A(new_n2866), .B(new_n2865), .Y(new_n2867));
  xor_4  g02491(.A(new_n2867), .B(new_n2864), .Y(new_n2868));
  xor_4  g02492(.A(new_n2868), .B(new_n2860), .Y(new_n2869));
  not_8  g02493(.A(new_n2869), .Y(new_n2870));
  nand_5 g02494(.A(new_n2830), .B(new_n2824), .Y(new_n2871));
  nand_5 g02495(.A(new_n2831), .B(new_n2811), .Y(new_n2872));
  nand_5 g02496(.A(new_n2872), .B(new_n2871), .Y(new_n2873));
  xor_4  g02497(.A(new_n2873), .B(new_n2829), .Y(new_n2874));
  xor_4  g02498(.A(new_n2874), .B(new_n2870), .Y(new_n2875));
  xnor_4 g02499(.A(new_n2875), .B(new_n2852), .Y(new_n2876));
  nand_5 g02500(.A(pi142), .B(pi124), .Y(new_n2877));
  xnor_4 g02501(.A(new_n2847), .B(new_n2846), .Y(new_n2878));
  not_8  g02502(.A(new_n2840), .Y(new_n2879));
  not_8  g02503(.A(new_n2839), .Y(new_n2880));
  nand_5 g02504(.A(pi170), .B(pi142), .Y(new_n2881));
  nand_5 g02505(.A(new_n2881), .B(new_n2879), .Y(new_n2882));
  nand_5 g02506(.A(new_n2882), .B(new_n2880), .Y(new_n2883));
  nand_5 g02507(.A(new_n2883), .B(new_n2841), .Y(new_n2884));
  nand_5 g02508(.A(new_n2884), .B(new_n2879), .Y(new_n2885));
  nor_5  g02509(.A(new_n2885), .B(new_n2878), .Y(new_n2886));
  xor_4  g02510(.A(new_n2849), .B(new_n2836), .Y(new_n2887));
  nand_5 g02511(.A(new_n2887), .B(new_n2886), .Y(new_n2888));
  nand_5 g02512(.A(new_n2888), .B(new_n2877), .Y(new_n2889));
  xnor_4 g02513(.A(new_n2851), .B(new_n2832), .Y(new_n2890));
  xor_4  g02514(.A(new_n2888), .B(new_n2877), .Y(new_n2891));
  nand_5 g02515(.A(new_n2891), .B(new_n2890), .Y(new_n2892));
  nand_5 g02516(.A(new_n2892), .B(new_n2889), .Y(new_n2893));
  xor_4  g02517(.A(new_n2893), .B(new_n2876), .Y(new_n2894));
  xor_4  g02518(.A(new_n2894), .B(new_n2794), .Y(new_n2895));
  xor_4  g02519(.A(new_n2791), .B(new_n2790), .Y(new_n2896));
  xor_4  g02520(.A(new_n2891), .B(new_n2890), .Y(new_n2897));
  or_6   g02521(.A(new_n2897), .B(new_n2896), .Y(new_n2898));
  xor_4  g02522(.A(new_n2897), .B(new_n2896), .Y(new_n2899));
  xor_4  g02523(.A(new_n2786), .B(new_n2785), .Y(new_n2900));
  xor_4  g02524(.A(new_n2887), .B(new_n2886), .Y(new_n2901));
  nand_5 g02525(.A(new_n2901), .B(new_n2900), .Y(new_n2902));
  not_8  g02526(.A(new_n2902), .Y(new_n2903));
  xnor_4 g02527(.A(new_n2901), .B(new_n2900), .Y(new_n2904));
  xnor_4 g02528(.A(new_n2784), .B(new_n2777), .Y(new_n2905));
  nor_5  g02529(.A(new_n2882), .B(new_n2880), .Y(new_n2906));
  or_6   g02530(.A(new_n2906), .B(new_n2884), .Y(new_n2907));
  nor_5  g02531(.A(new_n2781), .B(new_n2779), .Y(new_n2908));
  nor_5  g02532(.A(new_n2908), .B(new_n2783), .Y(new_n2909));
  not_8  g02533(.A(new_n2909), .Y(new_n2910));
  nand_5 g02534(.A(new_n2910), .B(new_n2907), .Y(new_n2911));
  xor_4  g02535(.A(new_n2909), .B(new_n2907), .Y(new_n2912));
  nor_5  g02536(.A(new_n2881), .B(new_n2780), .Y(new_n2913));
  nand_5 g02537(.A(pi158), .B(pi087), .Y(new_n2914));
  nand_5 g02538(.A(pi254), .B(pi219), .Y(new_n2915));
  xor_4  g02539(.A(new_n2915), .B(new_n2914), .Y(new_n2916));
  nand_5 g02540(.A(new_n2916), .B(new_n2913), .Y(new_n2917));
  nand_5 g02541(.A(pi142), .B(pi004), .Y(new_n2918));
  nand_5 g02542(.A(pi170), .B(pi071), .Y(new_n2919));
  xor_4  g02543(.A(new_n2919), .B(new_n2918), .Y(new_n2920));
  xor_4  g02544(.A(new_n2916), .B(new_n2913), .Y(new_n2921));
  nand_5 g02545(.A(new_n2921), .B(new_n2920), .Y(new_n2922));
  nand_5 g02546(.A(new_n2922), .B(new_n2917), .Y(new_n2923));
  or_6   g02547(.A(new_n2923), .B(new_n2912), .Y(new_n2924));
  nand_5 g02548(.A(new_n2924), .B(new_n2911), .Y(new_n2925));
  nand_5 g02549(.A(new_n2925), .B(new_n2905), .Y(new_n2926));
  xor_4  g02550(.A(new_n2885), .B(new_n2878), .Y(new_n2927));
  not_8  g02551(.A(new_n2927), .Y(new_n2928));
  xor_4  g02552(.A(new_n2925), .B(new_n2905), .Y(new_n2929));
  nand_5 g02553(.A(new_n2929), .B(new_n2928), .Y(new_n2930));
  nand_5 g02554(.A(new_n2930), .B(new_n2926), .Y(new_n2931));
  nor_5  g02555(.A(new_n2931), .B(new_n2904), .Y(new_n2932));
  nor_5  g02556(.A(new_n2932), .B(new_n2903), .Y(new_n2933));
  not_8  g02557(.A(new_n2933), .Y(new_n2934));
  nand_5 g02558(.A(new_n2934), .B(new_n2899), .Y(new_n2935));
  nand_5 g02559(.A(new_n2935), .B(new_n2898), .Y(new_n2936));
  xor_4  g02560(.A(new_n2936), .B(new_n2895), .Y(new_n2937));
  xor_4  g02561(.A(new_n2937), .B(new_n2693), .Y(new_n2938));
  xor_4  g02562(.A(new_n2933), .B(new_n2899), .Y(new_n2939));
  xor_4  g02563(.A(new_n2690), .B(new_n2689), .Y(new_n2940));
  nor_5  g02564(.A(new_n2940), .B(new_n2939), .Y(new_n2941));
  xnor_4 g02565(.A(new_n2940), .B(new_n2939), .Y(new_n2942));
  xor_4  g02566(.A(new_n2686), .B(new_n2685), .Y(new_n2943));
  xor_4  g02567(.A(new_n2929), .B(new_n2928), .Y(new_n2944));
  not_8  g02568(.A(new_n2944), .Y(new_n2945));
  xor_4  g02569(.A(new_n2684), .B(new_n2683), .Y(new_n2946));
  nor_5  g02570(.A(new_n2946), .B(new_n2945), .Y(new_n2947));
  xor_4  g02571(.A(new_n2946), .B(new_n2944), .Y(new_n2948));
  xor_4  g02572(.A(new_n2681), .B(new_n2679), .Y(new_n2949));
  xor_4  g02573(.A(new_n2881), .B(new_n2780), .Y(new_n2950));
  not_8  g02574(.A(new_n2950), .Y(new_n2951));
  or_6   g02575(.A(new_n2951), .B(new_n2680), .Y(new_n2952));
  nand_5 g02576(.A(pi138), .B(pi062), .Y(new_n2953));
  nand_5 g02577(.A(pi182), .B(pi065), .Y(new_n2954));
  nand_5 g02578(.A(new_n2954), .B(new_n2953), .Y(new_n2955));
  nand_5 g02579(.A(new_n2955), .B(new_n2682), .Y(new_n2956));
  nand_5 g02580(.A(new_n2956), .B(new_n2952), .Y(new_n2957));
  xor_4  g02581(.A(new_n2921), .B(new_n2920), .Y(new_n2958));
  not_8  g02582(.A(new_n2958), .Y(new_n2959));
  xor_4  g02583(.A(new_n2956), .B(new_n2952), .Y(new_n2960));
  nand_5 g02584(.A(new_n2960), .B(new_n2959), .Y(new_n2961));
  nand_5 g02585(.A(new_n2961), .B(new_n2957), .Y(new_n2962));
  or_6   g02586(.A(new_n2962), .B(new_n2949), .Y(new_n2963));
  xnor_4 g02587(.A(new_n2923), .B(new_n2912), .Y(new_n2964));
  xor_4  g02588(.A(new_n2962), .B(new_n2949), .Y(new_n2965));
  nand_5 g02589(.A(new_n2965), .B(new_n2964), .Y(new_n2966));
  nand_5 g02590(.A(new_n2966), .B(new_n2963), .Y(new_n2967));
  nor_5  g02591(.A(new_n2967), .B(new_n2948), .Y(new_n2968));
  nor_5  g02592(.A(new_n2968), .B(new_n2947), .Y(new_n2969));
  or_6   g02593(.A(new_n2969), .B(new_n2943), .Y(new_n2970));
  xor_4  g02594(.A(new_n2931), .B(new_n2904), .Y(new_n2971));
  not_8  g02595(.A(new_n2971), .Y(new_n2972));
  xor_4  g02596(.A(new_n2969), .B(new_n2943), .Y(new_n2973));
  nand_5 g02597(.A(new_n2973), .B(new_n2972), .Y(new_n2974));
  nand_5 g02598(.A(new_n2974), .B(new_n2970), .Y(new_n2975));
  nor_5  g02599(.A(new_n2975), .B(new_n2942), .Y(new_n2976));
  nor_5  g02600(.A(new_n2976), .B(new_n2941), .Y(new_n2977));
  xnor_4 g02601(.A(new_n2977), .B(new_n2938), .Y(new_n2978));
  nand_5 g02602(.A(pi190), .B(pi101), .Y(new_n2979));
  nand_5 g02603(.A(pi229), .B(pi060), .Y(new_n2980));
  nand_5 g02604(.A(pi223), .B(pi092), .Y(new_n2981));
  xor_4  g02605(.A(new_n2981), .B(new_n2980), .Y(new_n2982));
  xor_4  g02606(.A(new_n2982), .B(new_n2979), .Y(new_n2983));
  nand_5 g02607(.A(pi067), .B(pi020), .Y(new_n2984));
  nand_5 g02608(.A(pi092), .B(pi060), .Y(new_n2985));
  nand_5 g02609(.A(pi229), .B(pi020), .Y(new_n2986));
  nand_5 g02610(.A(new_n2986), .B(new_n2985), .Y(new_n2987));
  nand_5 g02611(.A(pi223), .B(pi190), .Y(new_n2988));
  xor_4  g02612(.A(new_n2986), .B(new_n2985), .Y(new_n2989));
  nand_5 g02613(.A(new_n2989), .B(new_n2988), .Y(new_n2990));
  nand_5 g02614(.A(new_n2990), .B(new_n2987), .Y(new_n2991));
  xor_4  g02615(.A(new_n2991), .B(new_n2984), .Y(new_n2992));
  xor_4  g02616(.A(new_n2992), .B(new_n2983), .Y(new_n2993));
  nand_5 g02617(.A(pi160), .B(pi053), .Y(new_n2994));
  or_6   g02618(.A(new_n2994), .B(new_n2993), .Y(new_n2995));
  xor_4  g02619(.A(new_n2994), .B(new_n2993), .Y(new_n2996));
  nand_5 g02620(.A(pi190), .B(pi060), .Y(new_n2997));
  nand_5 g02621(.A(pi229), .B(pi160), .Y(new_n2998));
  nand_5 g02622(.A(new_n2998), .B(new_n2997), .Y(new_n2999));
  nand_5 g02623(.A(pi092), .B(pi020), .Y(new_n3000));
  or_6   g02624(.A(new_n2998), .B(new_n2997), .Y(new_n3001));
  nand_5 g02625(.A(new_n3001), .B(new_n3000), .Y(new_n3002));
  nand_5 g02626(.A(new_n3002), .B(new_n2999), .Y(new_n3003));
  nand_5 g02627(.A(pi160), .B(pi067), .Y(new_n3004));
  or_6   g02628(.A(new_n3004), .B(new_n3003), .Y(new_n3005));
  xnor_4 g02629(.A(new_n2989), .B(new_n2988), .Y(new_n3006));
  xor_4  g02630(.A(new_n3004), .B(new_n3003), .Y(new_n3007));
  nand_5 g02631(.A(new_n3007), .B(new_n3006), .Y(new_n3008));
  nand_5 g02632(.A(new_n3008), .B(new_n3005), .Y(new_n3009));
  nand_5 g02633(.A(new_n3009), .B(new_n2996), .Y(new_n3010));
  nand_5 g02634(.A(new_n3010), .B(new_n2995), .Y(new_n3011));
  nand_5 g02635(.A(pi229), .B(pi223), .Y(new_n3012));
  nand_5 g02636(.A(new_n2981), .B(new_n2980), .Y(new_n3013));
  nand_5 g02637(.A(new_n2982), .B(new_n2979), .Y(new_n3014));
  nand_5 g02638(.A(new_n3014), .B(new_n3013), .Y(new_n3015));
  nand_5 g02639(.A(pi225), .B(pi190), .Y(new_n3016));
  nand_5 g02640(.A(pi101), .B(pi092), .Y(new_n3017));
  nand_5 g02641(.A(new_n3017), .B(new_n3016), .Y(new_n3018));
  nand_5 g02642(.A(pi225), .B(pi092), .Y(new_n3019));
  or_6   g02643(.A(new_n3019), .B(new_n2979), .Y(new_n3020));
  nand_5 g02644(.A(new_n3020), .B(new_n3018), .Y(new_n3021));
  xnor_4 g02645(.A(new_n3021), .B(new_n3015), .Y(new_n3022));
  xnor_4 g02646(.A(new_n3022), .B(new_n3012), .Y(new_n3023));
  nand_5 g02647(.A(new_n2991), .B(new_n2984), .Y(new_n3024));
  nand_5 g02648(.A(new_n2992), .B(new_n2983), .Y(new_n3025));
  nand_5 g02649(.A(new_n3025), .B(new_n3024), .Y(new_n3026));
  xor_4  g02650(.A(new_n3026), .B(new_n3023), .Y(new_n3027));
  nand_5 g02651(.A(pi067), .B(pi060), .Y(new_n3028));
  nand_5 g02652(.A(pi053), .B(pi020), .Y(new_n3029));
  nand_5 g02653(.A(new_n3029), .B(new_n3028), .Y(new_n3030));
  nand_5 g02654(.A(pi060), .B(pi053), .Y(new_n3031));
  nor_5  g02655(.A(new_n3031), .B(new_n2984), .Y(new_n3032));
  not_8  g02656(.A(new_n3032), .Y(new_n3033));
  nand_5 g02657(.A(new_n3033), .B(new_n3030), .Y(new_n3034));
  xnor_4 g02658(.A(new_n3034), .B(new_n3027), .Y(new_n3035));
  nand_5 g02659(.A(new_n3035), .B(new_n3011), .Y(new_n3036));
  nand_5 g02660(.A(new_n3026), .B(new_n3023), .Y(new_n3037));
  nand_5 g02661(.A(new_n3034), .B(new_n3027), .Y(new_n3038));
  nand_5 g02662(.A(new_n3038), .B(new_n3037), .Y(new_n3039));
  nand_5 g02663(.A(new_n3039), .B(new_n3033), .Y(new_n3040));
  nor_5  g02664(.A(new_n3026), .B(new_n3023), .Y(new_n3041));
  nand_5 g02665(.A(new_n3032), .B(new_n3041), .Y(new_n3042));
  nand_5 g02666(.A(new_n3042), .B(new_n3040), .Y(new_n3043));
  nand_5 g02667(.A(pi190), .B(pi177), .Y(new_n3044));
  nand_5 g02668(.A(pi229), .B(pi101), .Y(new_n3045));
  xor_4  g02669(.A(new_n3045), .B(new_n3044), .Y(new_n3046));
  xor_4  g02670(.A(new_n3046), .B(new_n3019), .Y(new_n3047));
  nand_5 g02671(.A(pi223), .B(pi067), .Y(new_n3048));
  xor_4  g02672(.A(new_n3048), .B(new_n3020), .Y(new_n3049));
  xor_4  g02673(.A(new_n3049), .B(new_n3047), .Y(new_n3050));
  nand_5 g02674(.A(pi160), .B(pi030), .Y(new_n3051));
  nand_5 g02675(.A(pi185), .B(pi020), .Y(new_n3052));
  xor_4  g02676(.A(new_n3052), .B(new_n3051), .Y(new_n3053));
  xor_4  g02677(.A(new_n3053), .B(new_n3031), .Y(new_n3054));
  nor_5  g02678(.A(new_n3021), .B(new_n3015), .Y(new_n3055));
  nor_5  g02679(.A(new_n3022), .B(new_n3012), .Y(new_n3056));
  nor_5  g02680(.A(new_n3056), .B(new_n3055), .Y(new_n3057));
  xor_4  g02681(.A(new_n3057), .B(new_n3054), .Y(new_n3058));
  xnor_4 g02682(.A(new_n3058), .B(new_n3050), .Y(new_n3059));
  xor_4  g02683(.A(new_n3059), .B(new_n3043), .Y(new_n3060));
  xnor_4 g02684(.A(new_n3060), .B(new_n3036), .Y(new_n3061));
  nand_5 g02685(.A(pi185), .B(pi160), .Y(new_n3062));
  xor_4  g02686(.A(new_n3007), .B(new_n3006), .Y(new_n3063));
  not_8  g02687(.A(new_n3063), .Y(new_n3064));
  not_8  g02688(.A(new_n3000), .Y(new_n3065));
  not_8  g02689(.A(new_n2999), .Y(new_n3066));
  nand_5 g02690(.A(pi190), .B(pi160), .Y(new_n3067));
  nand_5 g02691(.A(new_n3067), .B(new_n3065), .Y(new_n3068));
  nand_5 g02692(.A(new_n3068), .B(new_n3066), .Y(new_n3069));
  nand_5 g02693(.A(new_n3069), .B(new_n3001), .Y(new_n3070));
  nand_5 g02694(.A(new_n3070), .B(new_n3065), .Y(new_n3071));
  nor_5  g02695(.A(new_n3071), .B(new_n3064), .Y(new_n3072));
  xor_4  g02696(.A(new_n3009), .B(new_n2996), .Y(new_n3073));
  nand_5 g02697(.A(new_n3073), .B(new_n3072), .Y(new_n3074));
  nand_5 g02698(.A(new_n3074), .B(new_n3062), .Y(new_n3075));
  xnor_4 g02699(.A(new_n3035), .B(new_n3011), .Y(new_n3076));
  xor_4  g02700(.A(new_n3074), .B(new_n3062), .Y(new_n3077));
  nand_5 g02701(.A(new_n3077), .B(new_n3076), .Y(new_n3078));
  nand_5 g02702(.A(new_n3078), .B(new_n3075), .Y(new_n3079));
  xor_4  g02703(.A(new_n3079), .B(new_n3061), .Y(new_n3080));
  xor_4  g02704(.A(new_n3080), .B(new_n2978), .Y(new_n3081));
  xor_4  g02705(.A(new_n2975), .B(new_n2942), .Y(new_n3082));
  not_8  g02706(.A(new_n3082), .Y(new_n3083));
  xor_4  g02707(.A(new_n3077), .B(new_n3076), .Y(new_n3084));
  or_6   g02708(.A(new_n3084), .B(new_n3083), .Y(new_n3085));
  xor_4  g02709(.A(new_n3073), .B(new_n3072), .Y(new_n3086));
  xor_4  g02710(.A(new_n3071), .B(new_n3063), .Y(new_n3087));
  xor_4  g02711(.A(new_n2950), .B(new_n2680), .Y(new_n3088));
  nor_5  g02712(.A(new_n3088), .B(new_n3067), .Y(new_n3089));
  nand_5 g02713(.A(pi160), .B(pi092), .Y(new_n3090));
  nand_5 g02714(.A(pi190), .B(pi020), .Y(new_n3091));
  xor_4  g02715(.A(new_n3091), .B(new_n3090), .Y(new_n3092));
  nand_5 g02716(.A(new_n3092), .B(new_n3089), .Y(new_n3093));
  xor_4  g02717(.A(new_n2960), .B(new_n2958), .Y(new_n3094));
  xor_4  g02718(.A(new_n3092), .B(new_n3089), .Y(new_n3095));
  nand_5 g02719(.A(new_n3095), .B(new_n3094), .Y(new_n3096));
  nand_5 g02720(.A(new_n3096), .B(new_n3093), .Y(new_n3097));
  nor_5  g02721(.A(new_n3068), .B(new_n3066), .Y(new_n3098));
  nor_5  g02722(.A(new_n3098), .B(new_n3070), .Y(new_n3099));
  or_6   g02723(.A(new_n3099), .B(new_n3097), .Y(new_n3100));
  xor_4  g02724(.A(new_n2965), .B(new_n2964), .Y(new_n3101));
  not_8  g02725(.A(new_n3101), .Y(new_n3102));
  xor_4  g02726(.A(new_n3099), .B(new_n3097), .Y(new_n3103));
  nand_5 g02727(.A(new_n3103), .B(new_n3102), .Y(new_n3104));
  nand_5 g02728(.A(new_n3104), .B(new_n3100), .Y(new_n3105));
  or_6   g02729(.A(new_n3105), .B(new_n3087), .Y(new_n3106));
  xnor_4 g02730(.A(new_n2967), .B(new_n2948), .Y(new_n3107));
  xor_4  g02731(.A(new_n3105), .B(new_n3087), .Y(new_n3108));
  nand_5 g02732(.A(new_n3108), .B(new_n3107), .Y(new_n3109));
  nand_5 g02733(.A(new_n3109), .B(new_n3106), .Y(new_n3110));
  nand_5 g02734(.A(new_n3110), .B(new_n3086), .Y(new_n3111));
  xor_4  g02735(.A(new_n2973), .B(new_n2971), .Y(new_n3112));
  xor_4  g02736(.A(new_n3110), .B(new_n3086), .Y(new_n3113));
  nand_5 g02737(.A(new_n3113), .B(new_n3112), .Y(new_n3114));
  nand_5 g02738(.A(new_n3114), .B(new_n3111), .Y(new_n3115));
  xor_4  g02739(.A(new_n3084), .B(new_n3083), .Y(new_n3116));
  nand_5 g02740(.A(new_n3116), .B(new_n3115), .Y(new_n3117));
  nand_5 g02741(.A(new_n3117), .B(new_n3085), .Y(new_n3118));
  xor_4  g02742(.A(new_n3118), .B(new_n3081), .Y(po007));
  nand_5 g02743(.A(pi236), .B(pi230), .Y(new_n3120));
  nand_5 g02744(.A(pi236), .B(pi173), .Y(new_n3121));
  nand_5 g02745(.A(pi161), .B(pi109), .Y(new_n3122));
  nand_5 g02746(.A(new_n3122), .B(new_n3121), .Y(new_n3123));
  nand_5 g02747(.A(pi241), .B(pi014), .Y(new_n3124));
  xor_4  g02748(.A(new_n3122), .B(new_n3121), .Y(new_n3125));
  nand_5 g02749(.A(new_n3125), .B(new_n3124), .Y(new_n3126));
  nand_5 g02750(.A(new_n3126), .B(new_n3123), .Y(new_n3127));
  xor_4  g02751(.A(new_n3127), .B(new_n3120), .Y(new_n3128));
  nand_5 g02752(.A(pi161), .B(pi014), .Y(new_n3129));
  nand_5 g02753(.A(pi141), .B(pi109), .Y(new_n3130));
  nand_5 g02754(.A(pi241), .B(pi173), .Y(new_n3131));
  xor_4  g02755(.A(new_n3131), .B(new_n3130), .Y(new_n3132));
  xnor_4 g02756(.A(new_n3132), .B(new_n3129), .Y(new_n3133));
  xnor_4 g02757(.A(new_n3133), .B(new_n3128), .Y(new_n3134));
  nand_5 g02758(.A(pi236), .B(pi109), .Y(new_n3135));
  nor_5  g02759(.A(new_n3125), .B(new_n3124), .Y(new_n3136));
  not_8  g02760(.A(new_n3136), .Y(new_n3137));
  nor_5  g02761(.A(new_n3137), .B(new_n3135), .Y(new_n3138));
  xor_4  g02762(.A(new_n3138), .B(new_n3134), .Y(new_n3139));
  nand_5 g02763(.A(pi212), .B(pi207), .Y(new_n3140));
  nand_5 g02764(.A(pi213), .B(pi066), .Y(new_n3141));
  xor_4  g02765(.A(new_n3141), .B(new_n3140), .Y(new_n3142));
  nand_5 g02766(.A(pi226), .B(pi104), .Y(new_n3143));
  xor_4  g02767(.A(new_n3143), .B(new_n3142), .Y(new_n3144));
  nand_5 g02768(.A(pi226), .B(pi213), .Y(new_n3145));
  nor_5  g02769(.A(new_n3145), .B(new_n3140), .Y(new_n3146));
  not_8  g02770(.A(new_n3146), .Y(new_n3147));
  nor_5  g02771(.A(new_n3147), .B(new_n3144), .Y(new_n3148));
  nand_5 g02772(.A(pi212), .B(pi066), .Y(new_n3149));
  nand_5 g02773(.A(pi207), .B(pi104), .Y(new_n3150));
  nand_5 g02774(.A(pi226), .B(pi013), .Y(new_n3151));
  xor_4  g02775(.A(new_n3151), .B(new_n3150), .Y(new_n3152));
  xor_4  g02776(.A(new_n3152), .B(new_n3149), .Y(new_n3153));
  nand_5 g02777(.A(pi213), .B(pi055), .Y(new_n3154));
  nand_5 g02778(.A(new_n3141), .B(new_n3140), .Y(new_n3155));
  nand_5 g02779(.A(new_n3143), .B(new_n3142), .Y(new_n3156));
  nand_5 g02780(.A(new_n3156), .B(new_n3155), .Y(new_n3157));
  xor_4  g02781(.A(new_n3157), .B(new_n3154), .Y(new_n3158));
  xor_4  g02782(.A(new_n3158), .B(new_n3153), .Y(new_n3159));
  not_8  g02783(.A(new_n3159), .Y(new_n3160));
  xor_4  g02784(.A(new_n3160), .B(new_n3148), .Y(new_n3161));
  xor_4  g02785(.A(new_n3161), .B(new_n3139), .Y(new_n3162));
  xor_4  g02786(.A(new_n3146), .B(new_n3144), .Y(new_n3163));
  nand_5 g02787(.A(pi213), .B(pi207), .Y(new_n3164));
  nand_5 g02788(.A(pi226), .B(pi212), .Y(new_n3165));
  nand_5 g02789(.A(new_n3165), .B(new_n3164), .Y(new_n3166));
  nand_5 g02790(.A(new_n3166), .B(new_n3147), .Y(new_n3167));
  nand_5 g02791(.A(pi241), .B(pi109), .Y(new_n3168));
  nand_5 g02792(.A(pi236), .B(pi014), .Y(new_n3169));
  nand_5 g02793(.A(new_n3169), .B(new_n3168), .Y(new_n3170));
  or_6   g02794(.A(new_n3135), .B(new_n3124), .Y(new_n3171));
  nand_5 g02795(.A(new_n3171), .B(new_n3170), .Y(new_n3172));
  nand_5 g02796(.A(new_n3172), .B(new_n3167), .Y(new_n3173));
  nor_5  g02797(.A(new_n3145), .B(new_n3135), .Y(new_n3174));
  not_8  g02798(.A(new_n3174), .Y(new_n3175));
  xor_4  g02799(.A(new_n3172), .B(new_n3167), .Y(new_n3176));
  nand_5 g02800(.A(new_n3176), .B(new_n3175), .Y(new_n3177));
  nand_5 g02801(.A(new_n3177), .B(new_n3173), .Y(new_n3178));
  nand_5 g02802(.A(new_n3178), .B(new_n3163), .Y(new_n3179));
  xor_4  g02803(.A(new_n3178), .B(new_n3163), .Y(new_n3180));
  not_8  g02804(.A(new_n3138), .Y(new_n3181));
  nand_5 g02805(.A(new_n3171), .B(new_n3126), .Y(new_n3182));
  or_6   g02806(.A(new_n3182), .B(new_n3136), .Y(new_n3183));
  nand_5 g02807(.A(new_n3183), .B(new_n3181), .Y(new_n3184));
  nand_5 g02808(.A(new_n3184), .B(new_n3180), .Y(new_n3185));
  nand_5 g02809(.A(new_n3185), .B(new_n3179), .Y(new_n3186));
  xor_4  g02810(.A(new_n3186), .B(new_n3162), .Y(new_n3187));
  nand_5 g02811(.A(pi208), .B(pi186), .Y(new_n3188));
  nand_5 g02812(.A(pi168), .B(pi058), .Y(new_n3189));
  xor_4  g02813(.A(new_n3189), .B(new_n3188), .Y(new_n3190));
  nand_5 g02814(.A(pi139), .B(pi132), .Y(new_n3191));
  xor_4  g02815(.A(new_n3191), .B(new_n3190), .Y(new_n3192));
  nand_5 g02816(.A(pi168), .B(pi132), .Y(new_n3193));
  or_6   g02817(.A(new_n3193), .B(new_n3188), .Y(new_n3194));
  or_6   g02818(.A(new_n3194), .B(new_n3192), .Y(new_n3195));
  nand_5 g02819(.A(pi211), .B(pi168), .Y(new_n3196));
  nand_5 g02820(.A(new_n3189), .B(new_n3188), .Y(new_n3197));
  nand_5 g02821(.A(new_n3191), .B(new_n3190), .Y(new_n3198));
  nand_5 g02822(.A(new_n3198), .B(new_n3197), .Y(new_n3199));
  xor_4  g02823(.A(new_n3199), .B(new_n3196), .Y(new_n3200));
  nand_5 g02824(.A(pi132), .B(pi035), .Y(new_n3201));
  nand_5 g02825(.A(pi208), .B(pi058), .Y(new_n3202));
  nand_5 g02826(.A(pi186), .B(pi139), .Y(new_n3203));
  xor_4  g02827(.A(new_n3203), .B(new_n3202), .Y(new_n3204));
  xnor_4 g02828(.A(new_n3204), .B(new_n3201), .Y(new_n3205));
  xnor_4 g02829(.A(new_n3205), .B(new_n3200), .Y(new_n3206));
  xor_4  g02830(.A(new_n3206), .B(new_n3195), .Y(new_n3207));
  xor_4  g02831(.A(new_n3194), .B(new_n3192), .Y(new_n3208));
  xor_4  g02832(.A(new_n3145), .B(new_n3135), .Y(new_n3209));
  not_8  g02833(.A(new_n3209), .Y(new_n3210));
  nor_5  g02834(.A(new_n3210), .B(new_n3193), .Y(new_n3211));
  not_8  g02835(.A(new_n3211), .Y(new_n3212));
  nand_5 g02836(.A(pi186), .B(pi168), .Y(new_n3213));
  nand_5 g02837(.A(pi208), .B(pi132), .Y(new_n3214));
  nand_5 g02838(.A(new_n3214), .B(new_n3213), .Y(new_n3215));
  nand_5 g02839(.A(new_n3215), .B(new_n3194), .Y(new_n3216));
  or_6   g02840(.A(new_n3216), .B(new_n3212), .Y(new_n3217));
  xor_4  g02841(.A(new_n3176), .B(new_n3174), .Y(new_n3218));
  xor_4  g02842(.A(new_n3216), .B(new_n3212), .Y(new_n3219));
  nand_5 g02843(.A(new_n3219), .B(new_n3218), .Y(new_n3220));
  nand_5 g02844(.A(new_n3220), .B(new_n3217), .Y(new_n3221));
  nand_5 g02845(.A(new_n3221), .B(new_n3208), .Y(new_n3222));
  xnor_4 g02846(.A(new_n3184), .B(new_n3180), .Y(new_n3223));
  xor_4  g02847(.A(new_n3221), .B(new_n3208), .Y(new_n3224));
  nand_5 g02848(.A(new_n3224), .B(new_n3223), .Y(new_n3225));
  nand_5 g02849(.A(new_n3225), .B(new_n3222), .Y(new_n3226));
  xor_4  g02850(.A(new_n3226), .B(new_n3207), .Y(new_n3227));
  xor_4  g02851(.A(new_n3227), .B(new_n3187), .Y(new_n3228));
  nand_5 g02852(.A(pi069), .B(pi052), .Y(new_n3229));
  nand_5 g02853(.A(pi244), .B(pi131), .Y(new_n3230));
  xor_4  g02854(.A(new_n3230), .B(new_n3229), .Y(new_n3231));
  nand_5 g02855(.A(pi077), .B(pi029), .Y(new_n3232));
  xor_4  g02856(.A(new_n3232), .B(new_n3231), .Y(new_n3233));
  nand_5 g02857(.A(pi131), .B(pi029), .Y(new_n3234));
  nor_5  g02858(.A(new_n3234), .B(new_n3229), .Y(new_n3235));
  not_8  g02859(.A(new_n3235), .Y(new_n3236));
  nor_5  g02860(.A(new_n3236), .B(new_n3233), .Y(new_n3237));
  nand_5 g02861(.A(pi133), .B(pi029), .Y(new_n3238));
  nand_5 g02862(.A(pi244), .B(pi052), .Y(new_n3239));
  nand_5 g02863(.A(pi077), .B(pi069), .Y(new_n3240));
  xor_4  g02864(.A(new_n3240), .B(new_n3239), .Y(new_n3241));
  xor_4  g02865(.A(new_n3241), .B(new_n3238), .Y(new_n3242));
  nand_5 g02866(.A(pi150), .B(pi131), .Y(new_n3243));
  nand_5 g02867(.A(new_n3230), .B(new_n3229), .Y(new_n3244));
  nand_5 g02868(.A(new_n3232), .B(new_n3231), .Y(new_n3245));
  nand_5 g02869(.A(new_n3245), .B(new_n3244), .Y(new_n3246));
  xor_4  g02870(.A(new_n3246), .B(new_n3243), .Y(new_n3247));
  xor_4  g02871(.A(new_n3247), .B(new_n3242), .Y(new_n3248));
  xor_4  g02872(.A(new_n3248), .B(new_n3237), .Y(new_n3249));
  xor_4  g02873(.A(new_n3235), .B(new_n3233), .Y(new_n3250));
  xor_4  g02874(.A(new_n3209), .B(new_n3193), .Y(new_n3251));
  nor_5  g02875(.A(new_n3251), .B(new_n3234), .Y(new_n3252));
  not_8  g02876(.A(new_n3252), .Y(new_n3253));
  nand_5 g02877(.A(pi131), .B(pi069), .Y(new_n3254));
  nand_5 g02878(.A(pi052), .B(pi029), .Y(new_n3255));
  nand_5 g02879(.A(new_n3255), .B(new_n3254), .Y(new_n3256));
  nand_5 g02880(.A(new_n3256), .B(new_n3236), .Y(new_n3257));
  nand_5 g02881(.A(new_n3257), .B(new_n3253), .Y(new_n3258));
  xnor_4 g02882(.A(new_n3219), .B(new_n3218), .Y(new_n3259));
  xor_4  g02883(.A(new_n3257), .B(new_n3253), .Y(new_n3260));
  nand_5 g02884(.A(new_n3260), .B(new_n3259), .Y(new_n3261));
  nand_5 g02885(.A(new_n3261), .B(new_n3258), .Y(new_n3262));
  nand_5 g02886(.A(new_n3262), .B(new_n3250), .Y(new_n3263));
  xor_4  g02887(.A(new_n3224), .B(new_n3223), .Y(new_n3264));
  not_8  g02888(.A(new_n3264), .Y(new_n3265));
  xor_4  g02889(.A(new_n3262), .B(new_n3250), .Y(new_n3266));
  nand_5 g02890(.A(new_n3266), .B(new_n3265), .Y(new_n3267));
  nand_5 g02891(.A(new_n3267), .B(new_n3263), .Y(new_n3268));
  xor_4  g02892(.A(new_n3268), .B(new_n3249), .Y(new_n3269));
  xor_4  g02893(.A(new_n3269), .B(new_n3228), .Y(po008));
  nand_5 g02894(.A(pi170), .B(pi013), .Y(new_n3271));
  nand_5 g02895(.A(pi212), .B(pi073), .Y(new_n3272));
  nand_5 g02896(.A(pi104), .B(pi004), .Y(new_n3273));
  xor_4  g02897(.A(new_n3273), .B(new_n3272), .Y(new_n3274));
  xor_4  g02898(.A(new_n3274), .B(new_n3271), .Y(new_n3275));
  nand_5 g02899(.A(pi213), .B(pi003), .Y(new_n3276));
  nand_5 g02900(.A(pi170), .B(pi104), .Y(new_n3277));
  nand_5 g02901(.A(pi213), .B(pi073), .Y(new_n3278));
  nand_5 g02902(.A(new_n3278), .B(new_n3277), .Y(new_n3279));
  nand_5 g02903(.A(pi212), .B(pi004), .Y(new_n3280));
  or_6   g02904(.A(new_n3278), .B(new_n3277), .Y(new_n3281));
  nand_5 g02905(.A(new_n3281), .B(new_n3280), .Y(new_n3282));
  nand_5 g02906(.A(new_n3282), .B(new_n3279), .Y(new_n3283));
  xor_4  g02907(.A(new_n3283), .B(new_n3276), .Y(new_n3284));
  xor_4  g02908(.A(new_n3284), .B(new_n3275), .Y(new_n3285));
  not_8  g02909(.A(new_n3280), .Y(new_n3286));
  not_8  g02910(.A(new_n3279), .Y(new_n3287));
  nand_5 g02911(.A(pi213), .B(pi170), .Y(new_n3288));
  nand_5 g02912(.A(new_n3288), .B(new_n3286), .Y(new_n3289));
  nand_5 g02913(.A(new_n3289), .B(new_n3287), .Y(new_n3290));
  nand_5 g02914(.A(new_n3290), .B(new_n3281), .Y(new_n3291));
  nand_5 g02915(.A(new_n3291), .B(new_n3286), .Y(new_n3292));
  nor_5  g02916(.A(new_n3292), .B(new_n3285), .Y(new_n3293));
  nand_5 g02917(.A(pi104), .B(pi073), .Y(new_n3294));
  nand_5 g02918(.A(pi170), .B(pi112), .Y(new_n3295));
  nand_5 g02919(.A(pi013), .B(pi004), .Y(new_n3296));
  xor_4  g02920(.A(new_n3296), .B(new_n3295), .Y(new_n3297));
  xor_4  g02921(.A(new_n3297), .B(new_n3294), .Y(new_n3298));
  nand_5 g02922(.A(pi212), .B(pi003), .Y(new_n3299));
  nand_5 g02923(.A(new_n3273), .B(new_n3272), .Y(new_n3300));
  nand_5 g02924(.A(new_n3274), .B(new_n3271), .Y(new_n3301));
  nand_5 g02925(.A(new_n3301), .B(new_n3300), .Y(new_n3302));
  xor_4  g02926(.A(new_n3302), .B(new_n3299), .Y(new_n3303));
  xnor_4 g02927(.A(new_n3303), .B(new_n3298), .Y(new_n3304));
  nand_5 g02928(.A(pi213), .B(pi130), .Y(new_n3305));
  or_6   g02929(.A(new_n3283), .B(new_n3276), .Y(new_n3306));
  not_8  g02930(.A(new_n3275), .Y(new_n3307));
  nand_5 g02931(.A(new_n3284), .B(new_n3307), .Y(new_n3308));
  nand_5 g02932(.A(new_n3308), .B(new_n3306), .Y(new_n3309));
  xor_4  g02933(.A(new_n3309), .B(new_n3305), .Y(new_n3310));
  xor_4  g02934(.A(new_n3310), .B(new_n3304), .Y(new_n3311));
  xor_4  g02935(.A(new_n3311), .B(new_n3293), .Y(new_n3312));
  nand_5 g02936(.A(pi241), .B(pi158), .Y(new_n3313));
  nand_5 g02937(.A(pi236), .B(pi089), .Y(new_n3314));
  xor_4  g02938(.A(new_n3314), .B(new_n3313), .Y(new_n3315));
  nand_5 g02939(.A(pi254), .B(pi161), .Y(new_n3316));
  xor_4  g02940(.A(new_n3316), .B(new_n3315), .Y(new_n3317));
  nand_5 g02941(.A(pi254), .B(pi236), .Y(new_n3318));
  or_6   g02942(.A(new_n3318), .B(new_n3313), .Y(new_n3319));
  or_6   g02943(.A(new_n3319), .B(new_n3317), .Y(new_n3320));
  nand_5 g02944(.A(pi236), .B(pi154), .Y(new_n3321));
  nand_5 g02945(.A(new_n3314), .B(new_n3313), .Y(new_n3322));
  nand_5 g02946(.A(new_n3316), .B(new_n3315), .Y(new_n3323));
  nand_5 g02947(.A(new_n3323), .B(new_n3322), .Y(new_n3324));
  xor_4  g02948(.A(new_n3324), .B(new_n3321), .Y(new_n3325));
  nand_5 g02949(.A(pi161), .B(pi158), .Y(new_n3326));
  nand_5 g02950(.A(pi241), .B(pi089), .Y(new_n3327));
  nand_5 g02951(.A(pi254), .B(pi141), .Y(new_n3328));
  xor_4  g02952(.A(new_n3328), .B(new_n3327), .Y(new_n3329));
  xnor_4 g02953(.A(new_n3329), .B(new_n3326), .Y(new_n3330));
  xnor_4 g02954(.A(new_n3330), .B(new_n3325), .Y(new_n3331));
  nor_5  g02955(.A(new_n3331), .B(new_n3320), .Y(new_n3332));
  nand_5 g02956(.A(pi158), .B(pi141), .Y(new_n3333));
  nand_5 g02957(.A(pi161), .B(pi089), .Y(new_n3334));
  nand_5 g02958(.A(pi254), .B(pi090), .Y(new_n3335));
  xor_4  g02959(.A(new_n3335), .B(new_n3334), .Y(new_n3336));
  xor_4  g02960(.A(new_n3336), .B(new_n3333), .Y(new_n3337));
  nand_5 g02961(.A(pi241), .B(pi154), .Y(new_n3338));
  nand_5 g02962(.A(new_n3328), .B(new_n3327), .Y(new_n3339));
  nand_5 g02963(.A(new_n3329), .B(new_n3326), .Y(new_n3340));
  nand_5 g02964(.A(new_n3340), .B(new_n3339), .Y(new_n3341));
  xor_4  g02965(.A(new_n3341), .B(new_n3338), .Y(new_n3342));
  xor_4  g02966(.A(new_n3342), .B(new_n3337), .Y(new_n3343));
  nand_5 g02967(.A(pi236), .B(pi095), .Y(new_n3344));
  or_6   g02968(.A(new_n3324), .B(new_n3321), .Y(new_n3345));
  nand_5 g02969(.A(new_n3330), .B(new_n3325), .Y(new_n3346));
  nand_5 g02970(.A(new_n3346), .B(new_n3345), .Y(new_n3347));
  xor_4  g02971(.A(new_n3347), .B(new_n3344), .Y(new_n3348));
  xor_4  g02972(.A(new_n3348), .B(new_n3343), .Y(new_n3349));
  xor_4  g02973(.A(new_n3349), .B(new_n3332), .Y(new_n3350));
  xor_4  g02974(.A(new_n3331), .B(new_n3320), .Y(new_n3351));
  xor_4  g02975(.A(new_n3292), .B(new_n3285), .Y(new_n3352));
  nand_5 g02976(.A(new_n3352), .B(new_n3351), .Y(new_n3353));
  xor_4  g02977(.A(new_n3352), .B(new_n3351), .Y(new_n3354));
  xor_4  g02978(.A(new_n3319), .B(new_n3317), .Y(new_n3355));
  nor_5  g02979(.A(new_n3289), .B(new_n3287), .Y(new_n3356));
  nor_5  g02980(.A(new_n3356), .B(new_n3291), .Y(new_n3357));
  nand_5 g02981(.A(new_n3357), .B(new_n3355), .Y(new_n3358));
  nand_5 g02982(.A(pi213), .B(pi004), .Y(new_n3359));
  nand_5 g02983(.A(pi212), .B(pi170), .Y(new_n3360));
  xor_4  g02984(.A(new_n3360), .B(new_n3359), .Y(new_n3361));
  not_8  g02985(.A(new_n3361), .Y(new_n3362));
  nand_5 g02986(.A(pi236), .B(pi158), .Y(new_n3363));
  nand_5 g02987(.A(pi254), .B(pi241), .Y(new_n3364));
  nand_5 g02988(.A(new_n3364), .B(new_n3363), .Y(new_n3365));
  nand_5 g02989(.A(new_n3365), .B(new_n3319), .Y(new_n3366));
  nand_5 g02990(.A(new_n3366), .B(new_n3362), .Y(new_n3367));
  not_8  g02991(.A(new_n3367), .Y(new_n3368));
  nor_5  g02992(.A(new_n3318), .B(new_n3288), .Y(new_n3369));
  xor_4  g02993(.A(new_n3366), .B(new_n3361), .Y(new_n3370));
  nor_5  g02994(.A(new_n3370), .B(new_n3369), .Y(new_n3371));
  nor_5  g02995(.A(new_n3371), .B(new_n3368), .Y(new_n3372));
  xor_4  g02996(.A(new_n3357), .B(new_n3355), .Y(new_n3373));
  nand_5 g02997(.A(new_n3373), .B(new_n3372), .Y(new_n3374));
  nand_5 g02998(.A(new_n3374), .B(new_n3358), .Y(new_n3375));
  nand_5 g02999(.A(new_n3375), .B(new_n3354), .Y(new_n3376));
  nand_5 g03000(.A(new_n3376), .B(new_n3353), .Y(new_n3377));
  xor_4  g03001(.A(new_n3377), .B(new_n3350), .Y(new_n3378));
  xnor_4 g03002(.A(new_n3378), .B(new_n3312), .Y(new_n3379));
  nand_5 g03003(.A(pi208), .B(pi062), .Y(new_n3380));
  nand_5 g03004(.A(pi168), .B(pi120), .Y(new_n3381));
  xor_4  g03005(.A(new_n3381), .B(new_n3380), .Y(new_n3382));
  nand_5 g03006(.A(pi139), .B(pi065), .Y(new_n3383));
  xor_4  g03007(.A(new_n3383), .B(new_n3382), .Y(new_n3384));
  nand_5 g03008(.A(pi168), .B(pi065), .Y(new_n3385));
  nor_5  g03009(.A(new_n3385), .B(new_n3380), .Y(new_n3386));
  not_8  g03010(.A(new_n3386), .Y(new_n3387));
  nor_5  g03011(.A(new_n3387), .B(new_n3384), .Y(new_n3388));
  not_8  g03012(.A(new_n3388), .Y(new_n3389));
  nand_5 g03013(.A(pi172), .B(pi168), .Y(new_n3390));
  nand_5 g03014(.A(new_n3381), .B(new_n3380), .Y(new_n3391));
  nand_5 g03015(.A(new_n3383), .B(new_n3382), .Y(new_n3392));
  nand_5 g03016(.A(new_n3392), .B(new_n3391), .Y(new_n3393));
  xor_4  g03017(.A(new_n3393), .B(new_n3390), .Y(new_n3394));
  nand_5 g03018(.A(pi208), .B(pi120), .Y(new_n3395));
  nand_5 g03019(.A(pi065), .B(pi035), .Y(new_n3396));
  nand_5 g03020(.A(pi139), .B(pi062), .Y(new_n3397));
  xor_4  g03021(.A(new_n3397), .B(new_n3396), .Y(new_n3398));
  xnor_4 g03022(.A(new_n3398), .B(new_n3395), .Y(new_n3399));
  xnor_4 g03023(.A(new_n3399), .B(new_n3394), .Y(new_n3400));
  nor_5  g03024(.A(new_n3400), .B(new_n3389), .Y(new_n3401));
  nand_5 g03025(.A(pi139), .B(pi120), .Y(new_n3402));
  nand_5 g03026(.A(pi062), .B(pi035), .Y(new_n3403));
  nand_5 g03027(.A(pi065), .B(pi015), .Y(new_n3404));
  xor_4  g03028(.A(new_n3404), .B(new_n3403), .Y(new_n3405));
  xor_4  g03029(.A(new_n3405), .B(new_n3402), .Y(new_n3406));
  nand_5 g03030(.A(pi208), .B(pi172), .Y(new_n3407));
  nand_5 g03031(.A(new_n3397), .B(new_n3396), .Y(new_n3408));
  nand_5 g03032(.A(new_n3398), .B(new_n3395), .Y(new_n3409));
  nand_5 g03033(.A(new_n3409), .B(new_n3408), .Y(new_n3410));
  xor_4  g03034(.A(new_n3410), .B(new_n3407), .Y(new_n3411));
  xor_4  g03035(.A(new_n3411), .B(new_n3406), .Y(new_n3412));
  nand_5 g03036(.A(pi198), .B(pi168), .Y(new_n3413));
  or_6   g03037(.A(new_n3393), .B(new_n3390), .Y(new_n3414));
  nand_5 g03038(.A(new_n3399), .B(new_n3394), .Y(new_n3415));
  nand_5 g03039(.A(new_n3415), .B(new_n3414), .Y(new_n3416));
  xor_4  g03040(.A(new_n3416), .B(new_n3413), .Y(new_n3417));
  xor_4  g03041(.A(new_n3417), .B(new_n3412), .Y(new_n3418));
  xnor_4 g03042(.A(new_n3418), .B(new_n3401), .Y(new_n3419));
  xor_4  g03043(.A(new_n3400), .B(new_n3389), .Y(new_n3420));
  xor_4  g03044(.A(new_n3375), .B(new_n3354), .Y(new_n3421));
  or_6   g03045(.A(new_n3421), .B(new_n3420), .Y(new_n3422));
  xor_4  g03046(.A(new_n3373), .B(new_n3372), .Y(new_n3423));
  xor_4  g03047(.A(new_n3387), .B(new_n3384), .Y(new_n3424));
  nor_5  g03048(.A(new_n3424), .B(new_n3423), .Y(new_n3425));
  xnor_4 g03049(.A(new_n3424), .B(new_n3423), .Y(new_n3426));
  xor_4  g03050(.A(new_n3318), .B(new_n3288), .Y(new_n3427));
  not_8  g03051(.A(new_n3427), .Y(new_n3428));
  or_6   g03052(.A(new_n3428), .B(new_n3385), .Y(new_n3429));
  nand_5 g03053(.A(pi168), .B(pi062), .Y(new_n3430));
  nand_5 g03054(.A(pi208), .B(pi065), .Y(new_n3431));
  nand_5 g03055(.A(new_n3431), .B(new_n3430), .Y(new_n3432));
  nand_5 g03056(.A(new_n3432), .B(new_n3387), .Y(new_n3433));
  or_6   g03057(.A(new_n3433), .B(new_n3429), .Y(new_n3434));
  xor_4  g03058(.A(new_n3370), .B(new_n3369), .Y(new_n3435));
  not_8  g03059(.A(new_n3435), .Y(new_n3436));
  xor_4  g03060(.A(new_n3433), .B(new_n3429), .Y(new_n3437));
  nand_5 g03061(.A(new_n3437), .B(new_n3436), .Y(new_n3438));
  nand_5 g03062(.A(new_n3438), .B(new_n3434), .Y(new_n3439));
  nor_5  g03063(.A(new_n3439), .B(new_n3426), .Y(new_n3440));
  or_6   g03064(.A(new_n3440), .B(new_n3425), .Y(new_n3441));
  xor_4  g03065(.A(new_n3421), .B(new_n3420), .Y(new_n3442));
  nand_5 g03066(.A(new_n3442), .B(new_n3441), .Y(new_n3443));
  nand_5 g03067(.A(new_n3443), .B(new_n3422), .Y(new_n3444));
  xor_4  g03068(.A(new_n3444), .B(new_n3419), .Y(new_n3445));
  xor_4  g03069(.A(new_n3445), .B(new_n3379), .Y(new_n3446));
  nand_5 g03070(.A(pi092), .B(pi052), .Y(new_n3447));
  nand_5 g03071(.A(pi229), .B(pi131), .Y(new_n3448));
  xor_4  g03072(.A(new_n3448), .B(new_n3447), .Y(new_n3449));
  nand_5 g03073(.A(pi190), .B(pi077), .Y(new_n3450));
  xor_4  g03074(.A(new_n3450), .B(new_n3449), .Y(new_n3451));
  nand_5 g03075(.A(pi190), .B(pi131), .Y(new_n3452));
  nor_5  g03076(.A(new_n3452), .B(new_n3447), .Y(new_n3453));
  not_8  g03077(.A(new_n3453), .Y(new_n3454));
  or_6   g03078(.A(new_n3454), .B(new_n3451), .Y(new_n3455));
  nand_5 g03079(.A(pi131), .B(pi067), .Y(new_n3456));
  nand_5 g03080(.A(new_n3448), .B(new_n3447), .Y(new_n3457));
  nand_5 g03081(.A(new_n3450), .B(new_n3449), .Y(new_n3458));
  nand_5 g03082(.A(new_n3458), .B(new_n3457), .Y(new_n3459));
  xor_4  g03083(.A(new_n3459), .B(new_n3456), .Y(new_n3460));
  nand_5 g03084(.A(pi229), .B(pi052), .Y(new_n3461));
  nand_5 g03085(.A(pi190), .B(pi133), .Y(new_n3462));
  nand_5 g03086(.A(pi092), .B(pi077), .Y(new_n3463));
  xor_4  g03087(.A(new_n3463), .B(new_n3462), .Y(new_n3464));
  xnor_4 g03088(.A(new_n3464), .B(new_n3461), .Y(new_n3465));
  xnor_4 g03089(.A(new_n3465), .B(new_n3460), .Y(new_n3466));
  nor_5  g03090(.A(new_n3466), .B(new_n3455), .Y(new_n3467));
  nand_5 g03091(.A(pi229), .B(pi077), .Y(new_n3468));
  nand_5 g03092(.A(pi133), .B(pi092), .Y(new_n3469));
  nand_5 g03093(.A(pi190), .B(pi189), .Y(new_n3470));
  xor_4  g03094(.A(new_n3470), .B(new_n3469), .Y(new_n3471));
  xor_4  g03095(.A(new_n3471), .B(new_n3468), .Y(new_n3472));
  nand_5 g03096(.A(pi067), .B(pi052), .Y(new_n3473));
  nand_5 g03097(.A(new_n3463), .B(new_n3462), .Y(new_n3474));
  nand_5 g03098(.A(new_n3464), .B(new_n3461), .Y(new_n3475));
  nand_5 g03099(.A(new_n3475), .B(new_n3474), .Y(new_n3476));
  xor_4  g03100(.A(new_n3476), .B(new_n3473), .Y(new_n3477));
  xor_4  g03101(.A(new_n3477), .B(new_n3472), .Y(new_n3478));
  nand_5 g03102(.A(pi131), .B(pi053), .Y(new_n3479));
  or_6   g03103(.A(new_n3459), .B(new_n3456), .Y(new_n3480));
  nand_5 g03104(.A(new_n3465), .B(new_n3460), .Y(new_n3481));
  nand_5 g03105(.A(new_n3481), .B(new_n3480), .Y(new_n3482));
  xor_4  g03106(.A(new_n3482), .B(new_n3479), .Y(new_n3483));
  xor_4  g03107(.A(new_n3483), .B(new_n3478), .Y(new_n3484));
  xor_4  g03108(.A(new_n3484), .B(new_n3467), .Y(new_n3485));
  xor_4  g03109(.A(new_n3442), .B(new_n3441), .Y(new_n3486));
  not_8  g03110(.A(new_n3486), .Y(new_n3487));
  xor_4  g03111(.A(new_n3466), .B(new_n3455), .Y(new_n3488));
  nor_5  g03112(.A(new_n3488), .B(new_n3487), .Y(new_n3489));
  xor_4  g03113(.A(new_n3488), .B(new_n3486), .Y(new_n3490));
  xor_4  g03114(.A(new_n3453), .B(new_n3451), .Y(new_n3491));
  xor_4  g03115(.A(new_n3427), .B(new_n3385), .Y(new_n3492));
  or_6   g03116(.A(new_n3492), .B(new_n3452), .Y(new_n3493));
  nand_5 g03117(.A(pi131), .B(pi092), .Y(new_n3494));
  nand_5 g03118(.A(pi190), .B(pi052), .Y(new_n3495));
  nand_5 g03119(.A(new_n3495), .B(new_n3494), .Y(new_n3496));
  nand_5 g03120(.A(new_n3496), .B(new_n3454), .Y(new_n3497));
  nand_5 g03121(.A(new_n3497), .B(new_n3493), .Y(new_n3498));
  xor_4  g03122(.A(new_n3437), .B(new_n3436), .Y(new_n3499));
  not_8  g03123(.A(new_n3499), .Y(new_n3500));
  xor_4  g03124(.A(new_n3497), .B(new_n3493), .Y(new_n3501));
  nand_5 g03125(.A(new_n3501), .B(new_n3500), .Y(new_n3502));
  nand_5 g03126(.A(new_n3502), .B(new_n3498), .Y(new_n3503));
  or_6   g03127(.A(new_n3503), .B(new_n3491), .Y(new_n3504));
  xnor_4 g03128(.A(new_n3439), .B(new_n3426), .Y(new_n3505));
  xor_4  g03129(.A(new_n3503), .B(new_n3491), .Y(new_n3506));
  nand_5 g03130(.A(new_n3506), .B(new_n3505), .Y(new_n3507));
  nand_5 g03131(.A(new_n3507), .B(new_n3504), .Y(new_n3508));
  nor_5  g03132(.A(new_n3508), .B(new_n3490), .Y(new_n3509));
  nor_5  g03133(.A(new_n3509), .B(new_n3489), .Y(new_n3510));
  xor_4  g03134(.A(new_n3510), .B(new_n3485), .Y(new_n3511));
  xor_4  g03135(.A(new_n3511), .B(new_n3446), .Y(po009));
  nand_5 g03136(.A(pi236), .B(pi051), .Y(new_n3513));
  nand_5 g03137(.A(pi213), .B(pi188), .Y(new_n3514));
  xor_4  g03138(.A(new_n3514), .B(new_n3513), .Y(new_n3515));
  nand_5 g03139(.A(pi168), .B(pi162), .Y(new_n3516));
  xor_4  g03140(.A(new_n3516), .B(new_n3515), .Y(new_n3517));
  nand_5 g03141(.A(pi143), .B(pi131), .Y(new_n3518));
  xor_4  g03142(.A(new_n3518), .B(new_n3517), .Y(po010));
  xor_4  g03143(.A(new_n1827), .B(new_n1825), .Y(po011));
  xnor_4 g03144(.A(new_n3508), .B(new_n3490), .Y(po012));
  nand_5 g03145(.A(pi244), .B(pi223), .Y(new_n3522));
  nand_5 g03146(.A(pi101), .B(pi069), .Y(new_n3523));
  nand_5 g03147(.A(pi225), .B(pi029), .Y(new_n3524));
  nand_5 g03148(.A(new_n3524), .B(new_n3523), .Y(new_n3525));
  nand_5 g03149(.A(pi101), .B(pi029), .Y(new_n3526));
  nand_5 g03150(.A(pi225), .B(pi069), .Y(new_n3527));
  or_6   g03151(.A(new_n3527), .B(new_n3526), .Y(new_n3528));
  nand_5 g03152(.A(new_n3528), .B(new_n3525), .Y(new_n3529));
  xor_4  g03153(.A(new_n3529), .B(new_n3522), .Y(new_n3530));
  nand_5 g03154(.A(pi223), .B(pi069), .Y(new_n3531));
  nand_5 g03155(.A(new_n3531), .B(new_n3526), .Y(new_n3532));
  nand_5 g03156(.A(pi244), .B(pi060), .Y(new_n3533));
  xor_4  g03157(.A(new_n3531), .B(new_n3526), .Y(new_n3534));
  nand_5 g03158(.A(new_n3534), .B(new_n3533), .Y(new_n3535));
  nand_5 g03159(.A(new_n3535), .B(new_n3532), .Y(new_n3536));
  xor_4  g03160(.A(new_n3536), .B(new_n3530), .Y(new_n3537));
  nand_5 g03161(.A(pi150), .B(pi060), .Y(new_n3538));
  nand_5 g03162(.A(pi221), .B(pi020), .Y(new_n3539));
  nand_5 g03163(.A(new_n3539), .B(new_n3538), .Y(new_n3540));
  nand_5 g03164(.A(pi150), .B(pi020), .Y(new_n3541));
  nand_5 g03165(.A(pi221), .B(pi060), .Y(new_n3542));
  nor_5  g03166(.A(new_n3542), .B(new_n3541), .Y(new_n3543));
  not_8  g03167(.A(new_n3543), .Y(new_n3544));
  nand_5 g03168(.A(new_n3544), .B(new_n3540), .Y(new_n3545));
  xnor_4 g03169(.A(new_n3545), .B(new_n3537), .Y(new_n3546));
  nand_5 g03170(.A(pi223), .B(pi029), .Y(new_n3547));
  nand_5 g03171(.A(pi244), .B(pi020), .Y(new_n3548));
  nand_5 g03172(.A(new_n3548), .B(new_n3547), .Y(new_n3549));
  nand_5 g03173(.A(pi069), .B(pi060), .Y(new_n3550));
  xor_4  g03174(.A(new_n3548), .B(new_n3547), .Y(new_n3551));
  nand_5 g03175(.A(new_n3551), .B(new_n3550), .Y(new_n3552));
  nand_5 g03176(.A(new_n3552), .B(new_n3549), .Y(new_n3553));
  nand_5 g03177(.A(new_n3553), .B(new_n3541), .Y(new_n3554));
  xor_4  g03178(.A(new_n3534), .B(new_n3533), .Y(new_n3555));
  xor_4  g03179(.A(new_n3553), .B(new_n3541), .Y(new_n3556));
  nand_5 g03180(.A(new_n3556), .B(new_n3555), .Y(new_n3557));
  nand_5 g03181(.A(new_n3557), .B(new_n3554), .Y(new_n3558));
  xor_4  g03182(.A(new_n3558), .B(new_n3546), .Y(new_n3559));
  xor_4  g03183(.A(new_n3556), .B(new_n3555), .Y(new_n3560));
  nand_5 g03184(.A(pi221), .B(pi160), .Y(new_n3561));
  nor_5  g03185(.A(new_n3561), .B(new_n3560), .Y(new_n3562));
  xnor_4 g03186(.A(new_n3561), .B(new_n3560), .Y(new_n3563));
  nand_5 g03187(.A(pi160), .B(pi150), .Y(new_n3564));
  nand_5 g03188(.A(pi069), .B(pi020), .Y(new_n3565));
  nand_5 g03189(.A(pi244), .B(pi160), .Y(new_n3566));
  nand_5 g03190(.A(new_n3566), .B(new_n3565), .Y(new_n3567));
  nand_5 g03191(.A(pi060), .B(pi029), .Y(new_n3568));
  xor_4  g03192(.A(new_n3566), .B(new_n3565), .Y(new_n3569));
  nand_5 g03193(.A(new_n3569), .B(new_n3568), .Y(new_n3570));
  nand_5 g03194(.A(new_n3570), .B(new_n3567), .Y(new_n3571));
  nand_5 g03195(.A(new_n3571), .B(new_n3564), .Y(new_n3572));
  xor_4  g03196(.A(new_n3551), .B(new_n3550), .Y(new_n3573));
  xor_4  g03197(.A(new_n3571), .B(new_n3564), .Y(new_n3574));
  nand_5 g03198(.A(new_n3574), .B(new_n3573), .Y(new_n3575));
  nand_5 g03199(.A(new_n3575), .B(new_n3572), .Y(new_n3576));
  nor_5  g03200(.A(new_n3576), .B(new_n3563), .Y(new_n3577));
  nor_5  g03201(.A(new_n3577), .B(new_n3562), .Y(new_n3578));
  not_8  g03202(.A(new_n3578), .Y(new_n3579));
  nand_5 g03203(.A(new_n3579), .B(new_n3559), .Y(new_n3580));
  nand_5 g03204(.A(pi177), .B(pi029), .Y(new_n3581));
  nand_5 g03205(.A(pi244), .B(pi101), .Y(new_n3582));
  xor_4  g03206(.A(new_n3582), .B(new_n3581), .Y(new_n3583));
  xor_4  g03207(.A(new_n3583), .B(new_n3527), .Y(new_n3584));
  nand_5 g03208(.A(pi223), .B(pi150), .Y(new_n3585));
  xor_4  g03209(.A(new_n3585), .B(new_n3528), .Y(new_n3586));
  xor_4  g03210(.A(new_n3586), .B(new_n3584), .Y(new_n3587));
  nand_5 g03211(.A(pi196), .B(pi020), .Y(new_n3588));
  nand_5 g03212(.A(pi184), .B(pi160), .Y(new_n3589));
  xor_4  g03213(.A(new_n3589), .B(new_n3588), .Y(new_n3590));
  xor_4  g03214(.A(new_n3590), .B(new_n3542), .Y(new_n3591));
  nand_5 g03215(.A(new_n3529), .B(new_n3522), .Y(new_n3592));
  nand_5 g03216(.A(new_n3536), .B(new_n3530), .Y(new_n3593));
  nand_5 g03217(.A(new_n3593), .B(new_n3592), .Y(new_n3594));
  xor_4  g03218(.A(new_n3594), .B(new_n3591), .Y(new_n3595));
  xnor_4 g03219(.A(new_n3595), .B(new_n3587), .Y(new_n3596));
  nor_5  g03220(.A(new_n3558), .B(new_n3546), .Y(new_n3597));
  and_6  g03221(.A(new_n3597), .B(new_n3543), .Y(new_n3598));
  or_6   g03222(.A(new_n3545), .B(new_n3537), .Y(new_n3599));
  nand_5 g03223(.A(new_n3599), .B(new_n3544), .Y(new_n3600));
  nor_5  g03224(.A(new_n3600), .B(new_n3597), .Y(new_n3601));
  or_6   g03225(.A(new_n3601), .B(new_n3598), .Y(new_n3602));
  xor_4  g03226(.A(new_n3602), .B(new_n3596), .Y(new_n3603));
  xnor_4 g03227(.A(new_n3603), .B(new_n3580), .Y(new_n3604));
  nand_5 g03228(.A(pi196), .B(pi160), .Y(new_n3605));
  xor_4  g03229(.A(new_n3569), .B(new_n3568), .Y(new_n3606));
  nand_5 g03230(.A(pi160), .B(pi029), .Y(new_n3607));
  nor_5  g03231(.A(new_n3607), .B(new_n3565), .Y(new_n3608));
  not_8  g03232(.A(new_n3608), .Y(new_n3609));
  nor_5  g03233(.A(new_n3609), .B(new_n3606), .Y(new_n3610));
  not_8  g03234(.A(new_n3610), .Y(new_n3611));
  xor_4  g03235(.A(new_n3574), .B(new_n3573), .Y(new_n3612));
  nor_5  g03236(.A(new_n3612), .B(new_n3611), .Y(new_n3613));
  xor_4  g03237(.A(new_n3576), .B(new_n3563), .Y(new_n3614));
  nand_5 g03238(.A(new_n3614), .B(new_n3613), .Y(new_n3615));
  nand_5 g03239(.A(new_n3615), .B(new_n3605), .Y(new_n3616));
  xor_4  g03240(.A(new_n3578), .B(new_n3559), .Y(new_n3617));
  xor_4  g03241(.A(new_n3615), .B(new_n3605), .Y(new_n3618));
  nand_5 g03242(.A(new_n3618), .B(new_n3617), .Y(new_n3619));
  nand_5 g03243(.A(new_n3619), .B(new_n3616), .Y(new_n3620));
  xor_4  g03244(.A(new_n3620), .B(new_n3604), .Y(new_n3621));
  xor_4  g03245(.A(new_n3614), .B(new_n3613), .Y(new_n3622));
  xor_4  g03246(.A(new_n3612), .B(new_n3610), .Y(new_n3623));
  xor_4  g03247(.A(new_n3608), .B(new_n3606), .Y(new_n3624));
  nand_5 g03248(.A(pi226), .B(pi169), .Y(new_n3625));
  nand_5 g03249(.A(pi207), .B(pi071), .Y(new_n3626));
  nand_5 g03250(.A(pi142), .B(pi066), .Y(new_n3627));
  xor_4  g03251(.A(new_n3627), .B(new_n3626), .Y(new_n3628));
  xor_4  g03252(.A(new_n3628), .B(new_n3625), .Y(new_n3629));
  nand_5 g03253(.A(pi207), .B(pi142), .Y(new_n3630));
  nand_5 g03254(.A(pi226), .B(pi071), .Y(new_n3631));
  nor_5  g03255(.A(new_n3631), .B(new_n3630), .Y(new_n3632));
  xor_4  g03256(.A(new_n3632), .B(new_n3629), .Y(new_n3633));
  xor_4  g03257(.A(new_n3631), .B(new_n3630), .Y(new_n3634));
  nand_5 g03258(.A(pi226), .B(pi142), .Y(new_n3635));
  nand_5 g03259(.A(pi109), .B(pi087), .Y(new_n3636));
  nor_5  g03260(.A(new_n3636), .B(new_n3635), .Y(new_n3637));
  nor_5  g03261(.A(new_n3637), .B(new_n3634), .Y(new_n3638));
  nand_5 g03262(.A(pi219), .B(pi109), .Y(new_n3639));
  nand_5 g03263(.A(pi087), .B(pi014), .Y(new_n3640));
  xor_4  g03264(.A(new_n3640), .B(new_n3639), .Y(new_n3641));
  xnor_4 g03265(.A(new_n3637), .B(new_n3634), .Y(new_n3642));
  nor_5  g03266(.A(new_n3642), .B(new_n3641), .Y(new_n3643));
  nor_5  g03267(.A(new_n3643), .B(new_n3638), .Y(new_n3644));
  nand_5 g03268(.A(pi173), .B(pi087), .Y(new_n3645));
  nand_5 g03269(.A(pi109), .B(pi102), .Y(new_n3646));
  nand_5 g03270(.A(new_n3646), .B(new_n3645), .Y(new_n3647));
  not_8  g03271(.A(new_n3647), .Y(new_n3648));
  nand_5 g03272(.A(pi219), .B(pi014), .Y(new_n3649));
  not_8  g03273(.A(new_n3649), .Y(new_n3650));
  nand_5 g03274(.A(new_n3650), .B(new_n3636), .Y(new_n3651));
  nor_5  g03275(.A(new_n3651), .B(new_n3648), .Y(new_n3652));
  nand_5 g03276(.A(new_n3651), .B(new_n3648), .Y(new_n3653));
  or_6   g03277(.A(new_n3646), .B(new_n3645), .Y(new_n3654));
  nand_5 g03278(.A(new_n3654), .B(new_n3653), .Y(new_n3655));
  nor_5  g03279(.A(new_n3655), .B(new_n3652), .Y(new_n3656));
  xor_4  g03280(.A(new_n3656), .B(new_n3644), .Y(new_n3657));
  xnor_4 g03281(.A(new_n3657), .B(new_n3633), .Y(new_n3658));
  nand_5 g03282(.A(pi132), .B(pi041), .Y(new_n3659));
  nand_5 g03283(.A(pi186), .B(pi182), .Y(new_n3660));
  nand_5 g03284(.A(pi138), .B(pi058), .Y(new_n3661));
  xor_4  g03285(.A(new_n3661), .B(new_n3660), .Y(new_n3662));
  xor_4  g03286(.A(new_n3662), .B(new_n3659), .Y(new_n3663));
  nand_5 g03287(.A(pi138), .B(pi132), .Y(new_n3664));
  or_6   g03288(.A(new_n3664), .B(new_n3660), .Y(new_n3665));
  xor_4  g03289(.A(new_n3665), .B(new_n3663), .Y(new_n3666));
  xor_4  g03290(.A(new_n3636), .B(new_n3635), .Y(new_n3667));
  not_8  g03291(.A(new_n3667), .Y(new_n3668));
  nor_5  g03292(.A(new_n3668), .B(new_n3664), .Y(new_n3669));
  not_8  g03293(.A(new_n3669), .Y(new_n3670));
  nand_5 g03294(.A(pi186), .B(pi138), .Y(new_n3671));
  nand_5 g03295(.A(pi182), .B(pi132), .Y(new_n3672));
  nand_5 g03296(.A(new_n3672), .B(new_n3671), .Y(new_n3673));
  nand_5 g03297(.A(new_n3673), .B(new_n3665), .Y(new_n3674));
  or_6   g03298(.A(new_n3674), .B(new_n3670), .Y(new_n3675));
  xnor_4 g03299(.A(new_n3642), .B(new_n3641), .Y(new_n3676));
  xor_4  g03300(.A(new_n3674), .B(new_n3670), .Y(new_n3677));
  nand_5 g03301(.A(new_n3677), .B(new_n3676), .Y(new_n3678));
  nand_5 g03302(.A(new_n3678), .B(new_n3675), .Y(new_n3679));
  xor_4  g03303(.A(new_n3679), .B(new_n3666), .Y(new_n3680));
  xnor_4 g03304(.A(new_n3680), .B(new_n3658), .Y(new_n3681));
  nand_5 g03305(.A(new_n3681), .B(new_n3624), .Y(new_n3682));
  xor_4  g03306(.A(new_n3667), .B(new_n3664), .Y(new_n3683));
  nor_5  g03307(.A(new_n3683), .B(new_n3607), .Y(new_n3684));
  not_8  g03308(.A(new_n3684), .Y(new_n3685));
  nand_5 g03309(.A(pi029), .B(pi020), .Y(new_n3686));
  nand_5 g03310(.A(pi160), .B(pi069), .Y(new_n3687));
  nand_5 g03311(.A(new_n3687), .B(new_n3686), .Y(new_n3688));
  nand_5 g03312(.A(new_n3688), .B(new_n3609), .Y(new_n3689));
  nand_5 g03313(.A(new_n3689), .B(new_n3685), .Y(new_n3690));
  xnor_4 g03314(.A(new_n3677), .B(new_n3676), .Y(new_n3691));
  xor_4  g03315(.A(new_n3689), .B(new_n3685), .Y(new_n3692));
  nand_5 g03316(.A(new_n3692), .B(new_n3691), .Y(new_n3693));
  nand_5 g03317(.A(new_n3693), .B(new_n3690), .Y(new_n3694));
  xor_4  g03318(.A(new_n3681), .B(new_n3624), .Y(new_n3695));
  nand_5 g03319(.A(new_n3695), .B(new_n3694), .Y(new_n3696));
  nand_5 g03320(.A(new_n3696), .B(new_n3682), .Y(new_n3697));
  or_6   g03321(.A(new_n3697), .B(new_n3623), .Y(new_n3698));
  or_6   g03322(.A(new_n3665), .B(new_n3663), .Y(new_n3699));
  nand_5 g03323(.A(pi182), .B(pi058), .Y(new_n3700));
  nand_5 g03324(.A(pi216), .B(pi132), .Y(new_n3701));
  nand_5 g03325(.A(pi186), .B(pi041), .Y(new_n3702));
  xor_4  g03326(.A(new_n3702), .B(new_n3701), .Y(new_n3703));
  xnor_4 g03327(.A(new_n3703), .B(new_n3700), .Y(new_n3704));
  nand_5 g03328(.A(pi211), .B(pi138), .Y(new_n3705));
  nand_5 g03329(.A(new_n3661), .B(new_n3660), .Y(new_n3706));
  nand_5 g03330(.A(new_n3662), .B(new_n3659), .Y(new_n3707));
  nand_5 g03331(.A(new_n3707), .B(new_n3706), .Y(new_n3708));
  xor_4  g03332(.A(new_n3708), .B(new_n3705), .Y(new_n3709));
  xnor_4 g03333(.A(new_n3709), .B(new_n3704), .Y(new_n3710));
  xor_4  g03334(.A(new_n3710), .B(new_n3699), .Y(new_n3711));
  nand_5 g03335(.A(new_n3654), .B(new_n3649), .Y(new_n3712));
  nand_5 g03336(.A(new_n3712), .B(new_n3647), .Y(new_n3713));
  nand_5 g03337(.A(pi230), .B(pi087), .Y(new_n3714));
  xor_4  g03338(.A(new_n3714), .B(new_n3713), .Y(new_n3715));
  nand_5 g03339(.A(pi109), .B(pi001), .Y(new_n3716));
  nand_5 g03340(.A(pi219), .B(pi173), .Y(new_n3717));
  nand_5 g03341(.A(pi102), .B(pi014), .Y(new_n3718));
  xor_4  g03342(.A(new_n3718), .B(new_n3717), .Y(new_n3719));
  xnor_4 g03343(.A(new_n3719), .B(new_n3716), .Y(new_n3720));
  xnor_4 g03344(.A(new_n3720), .B(new_n3715), .Y(new_n3721));
  nand_5 g03345(.A(new_n3655), .B(new_n3650), .Y(new_n3722));
  xor_4  g03346(.A(new_n3722), .B(new_n3721), .Y(new_n3723));
  not_8  g03347(.A(new_n3723), .Y(new_n3724));
  not_8  g03348(.A(new_n3632), .Y(new_n3725));
  nor_5  g03349(.A(new_n3725), .B(new_n3629), .Y(new_n3726));
  nand_5 g03350(.A(pi207), .B(pi169), .Y(new_n3727));
  nand_5 g03351(.A(pi071), .B(pi066), .Y(new_n3728));
  nand_5 g03352(.A(pi226), .B(pi123), .Y(new_n3729));
  xor_4  g03353(.A(new_n3729), .B(new_n3728), .Y(new_n3730));
  xnor_4 g03354(.A(new_n3730), .B(new_n3727), .Y(new_n3731));
  nand_5 g03355(.A(pi142), .B(pi055), .Y(new_n3732));
  nand_5 g03356(.A(new_n3627), .B(new_n3626), .Y(new_n3733));
  nand_5 g03357(.A(new_n3628), .B(new_n3625), .Y(new_n3734));
  nand_5 g03358(.A(new_n3734), .B(new_n3733), .Y(new_n3735));
  xor_4  g03359(.A(new_n3735), .B(new_n3732), .Y(new_n3736));
  xnor_4 g03360(.A(new_n3736), .B(new_n3731), .Y(new_n3737));
  xor_4  g03361(.A(new_n3737), .B(new_n3726), .Y(new_n3738));
  or_6   g03362(.A(new_n3656), .B(new_n3644), .Y(new_n3739));
  nand_5 g03363(.A(new_n3657), .B(new_n3633), .Y(new_n3740));
  nand_5 g03364(.A(new_n3740), .B(new_n3739), .Y(new_n3741));
  xor_4  g03365(.A(new_n3741), .B(new_n3738), .Y(new_n3742));
  xor_4  g03366(.A(new_n3742), .B(new_n3724), .Y(new_n3743));
  not_8  g03367(.A(new_n3743), .Y(new_n3744));
  xor_4  g03368(.A(new_n3744), .B(new_n3711), .Y(new_n3745));
  nand_5 g03369(.A(new_n3679), .B(new_n3666), .Y(new_n3746));
  nand_5 g03370(.A(new_n3680), .B(new_n3658), .Y(new_n3747));
  nand_5 g03371(.A(new_n3747), .B(new_n3746), .Y(new_n3748));
  xor_4  g03372(.A(new_n3748), .B(new_n3745), .Y(new_n3749));
  xor_4  g03373(.A(new_n3697), .B(new_n3623), .Y(new_n3750));
  nand_5 g03374(.A(new_n3750), .B(new_n3749), .Y(new_n3751));
  nand_5 g03375(.A(new_n3751), .B(new_n3698), .Y(new_n3752));
  or_6   g03376(.A(new_n3752), .B(new_n3622), .Y(new_n3753));
  not_8  g03377(.A(new_n3726), .Y(new_n3754));
  nor_5  g03378(.A(new_n3737), .B(new_n3754), .Y(new_n3755));
  nand_5 g03379(.A(pi207), .B(pi123), .Y(new_n3756));
  nand_5 g03380(.A(pi226), .B(pi099), .Y(new_n3757));
  nand_5 g03381(.A(pi169), .B(pi066), .Y(new_n3758));
  xor_4  g03382(.A(new_n3758), .B(new_n3757), .Y(new_n3759));
  xor_4  g03383(.A(new_n3759), .B(new_n3756), .Y(new_n3760));
  nand_5 g03384(.A(pi071), .B(pi055), .Y(new_n3761));
  nand_5 g03385(.A(new_n3729), .B(new_n3728), .Y(new_n3762));
  nand_5 g03386(.A(new_n3730), .B(new_n3727), .Y(new_n3763));
  nand_5 g03387(.A(new_n3763), .B(new_n3762), .Y(new_n3764));
  xor_4  g03388(.A(new_n3764), .B(new_n3761), .Y(new_n3765));
  xor_4  g03389(.A(new_n3765), .B(new_n3760), .Y(new_n3766));
  nand_5 g03390(.A(pi142), .B(pi002), .Y(new_n3767));
  or_6   g03391(.A(new_n3735), .B(new_n3732), .Y(new_n3768));
  nand_5 g03392(.A(new_n3736), .B(new_n3731), .Y(new_n3769));
  nand_5 g03393(.A(new_n3769), .B(new_n3768), .Y(new_n3770));
  xor_4  g03394(.A(new_n3770), .B(new_n3767), .Y(new_n3771));
  xor_4  g03395(.A(new_n3771), .B(new_n3766), .Y(new_n3772));
  xnor_4 g03396(.A(new_n3772), .B(new_n3755), .Y(new_n3773));
  nor_5  g03397(.A(new_n3722), .B(new_n3721), .Y(new_n3774));
  nand_5 g03398(.A(pi087), .B(pi050), .Y(new_n3775));
  or_6   g03399(.A(new_n3714), .B(new_n3713), .Y(new_n3776));
  nand_5 g03400(.A(new_n3720), .B(new_n3715), .Y(new_n3777));
  nand_5 g03401(.A(new_n3777), .B(new_n3776), .Y(new_n3778));
  xor_4  g03402(.A(new_n3778), .B(new_n3775), .Y(new_n3779));
  nand_5 g03403(.A(pi173), .B(pi102), .Y(new_n3780));
  nand_5 g03404(.A(pi014), .B(pi001), .Y(new_n3781));
  nand_5 g03405(.A(pi122), .B(pi109), .Y(new_n3782));
  xor_4  g03406(.A(new_n3782), .B(new_n3781), .Y(new_n3783));
  xor_4  g03407(.A(new_n3783), .B(new_n3780), .Y(new_n3784));
  nand_5 g03408(.A(pi230), .B(pi219), .Y(new_n3785));
  nand_5 g03409(.A(new_n3718), .B(new_n3717), .Y(new_n3786));
  nand_5 g03410(.A(new_n3719), .B(new_n3716), .Y(new_n3787));
  nand_5 g03411(.A(new_n3787), .B(new_n3786), .Y(new_n3788));
  xor_4  g03412(.A(new_n3788), .B(new_n3785), .Y(new_n3789));
  xor_4  g03413(.A(new_n3789), .B(new_n3784), .Y(new_n3790));
  xor_4  g03414(.A(new_n3790), .B(new_n3779), .Y(new_n3791));
  xnor_4 g03415(.A(new_n3791), .B(new_n3774), .Y(new_n3792));
  nand_5 g03416(.A(new_n3741), .B(new_n3738), .Y(new_n3793));
  nand_5 g03417(.A(new_n3742), .B(new_n3724), .Y(new_n3794));
  nand_5 g03418(.A(new_n3794), .B(new_n3793), .Y(new_n3795));
  xor_4  g03419(.A(new_n3795), .B(new_n3792), .Y(new_n3796));
  xnor_4 g03420(.A(new_n3796), .B(new_n3773), .Y(new_n3797));
  nor_5  g03421(.A(new_n3710), .B(new_n3699), .Y(new_n3798));
  nand_5 g03422(.A(pi132), .B(pi076), .Y(new_n3799));
  nand_5 g03423(.A(pi216), .B(pi186), .Y(new_n3800));
  nand_5 g03424(.A(pi058), .B(pi041), .Y(new_n3801));
  xor_4  g03425(.A(new_n3801), .B(new_n3800), .Y(new_n3802));
  xor_4  g03426(.A(new_n3802), .B(new_n3799), .Y(new_n3803));
  nand_5 g03427(.A(pi211), .B(pi182), .Y(new_n3804));
  nand_5 g03428(.A(new_n3702), .B(new_n3701), .Y(new_n3805));
  nand_5 g03429(.A(new_n3703), .B(new_n3700), .Y(new_n3806));
  nand_5 g03430(.A(new_n3806), .B(new_n3805), .Y(new_n3807));
  xor_4  g03431(.A(new_n3807), .B(new_n3804), .Y(new_n3808));
  xor_4  g03432(.A(new_n3808), .B(new_n3803), .Y(new_n3809));
  nand_5 g03433(.A(pi199), .B(pi138), .Y(new_n3810));
  or_6   g03434(.A(new_n3708), .B(new_n3705), .Y(new_n3811));
  nand_5 g03435(.A(new_n3709), .B(new_n3704), .Y(new_n3812));
  nand_5 g03436(.A(new_n3812), .B(new_n3811), .Y(new_n3813));
  xor_4  g03437(.A(new_n3813), .B(new_n3810), .Y(new_n3814));
  xor_4  g03438(.A(new_n3814), .B(new_n3809), .Y(new_n3815));
  xor_4  g03439(.A(new_n3815), .B(new_n3798), .Y(new_n3816));
  nor_5  g03440(.A(new_n3744), .B(new_n3711), .Y(new_n3817));
  not_8  g03441(.A(new_n3745), .Y(new_n3818));
  nor_5  g03442(.A(new_n3748), .B(new_n3818), .Y(new_n3819));
  nor_5  g03443(.A(new_n3819), .B(new_n3817), .Y(new_n3820));
  xor_4  g03444(.A(new_n3820), .B(new_n3816), .Y(new_n3821));
  xor_4  g03445(.A(new_n3821), .B(new_n3797), .Y(new_n3822));
  not_8  g03446(.A(new_n3822), .Y(new_n3823));
  xor_4  g03447(.A(new_n3752), .B(new_n3622), .Y(new_n3824));
  nand_5 g03448(.A(new_n3824), .B(new_n3823), .Y(new_n3825));
  nand_5 g03449(.A(new_n3825), .B(new_n3753), .Y(new_n3826));
  xor_4  g03450(.A(new_n3618), .B(new_n3617), .Y(new_n3827));
  or_6   g03451(.A(new_n3827), .B(new_n3826), .Y(new_n3828));
  nand_5 g03452(.A(new_n3795), .B(new_n3792), .Y(new_n3829));
  nand_5 g03453(.A(new_n3796), .B(new_n3773), .Y(new_n3830));
  nand_5 g03454(.A(new_n3830), .B(new_n3829), .Y(new_n3831));
  and_6  g03455(.A(new_n3772), .B(new_n3755), .Y(new_n3832));
  nand_5 g03456(.A(pi142), .B(pi025), .Y(new_n3833));
  nand_5 g03457(.A(pi123), .B(pi066), .Y(new_n3834));
  nand_5 g03458(.A(pi226), .B(pi023), .Y(new_n3835));
  nand_5 g03459(.A(pi207), .B(pi099), .Y(new_n3836));
  nand_5 g03460(.A(new_n3836), .B(new_n3835), .Y(new_n3837));
  nand_5 g03461(.A(pi207), .B(pi023), .Y(new_n3838));
  or_6   g03462(.A(new_n3838), .B(new_n3757), .Y(new_n3839));
  nand_5 g03463(.A(new_n3839), .B(new_n3837), .Y(new_n3840));
  xor_4  g03464(.A(new_n3840), .B(new_n3834), .Y(new_n3841));
  nand_5 g03465(.A(new_n3758), .B(new_n3757), .Y(new_n3842));
  nand_5 g03466(.A(new_n3759), .B(new_n3756), .Y(new_n3843));
  nand_5 g03467(.A(new_n3843), .B(new_n3842), .Y(new_n3844));
  xor_4  g03468(.A(new_n3844), .B(new_n3841), .Y(new_n3845));
  nand_5 g03469(.A(new_n3764), .B(new_n3761), .Y(new_n3846));
  nand_5 g03470(.A(new_n3765), .B(new_n3760), .Y(new_n3847));
  nand_5 g03471(.A(new_n3847), .B(new_n3846), .Y(new_n3848));
  nand_5 g03472(.A(pi071), .B(pi002), .Y(new_n3849));
  nand_5 g03473(.A(pi169), .B(pi055), .Y(new_n3850));
  nand_5 g03474(.A(new_n3850), .B(new_n3849), .Y(new_n3851));
  nand_5 g03475(.A(pi169), .B(pi002), .Y(new_n3852));
  or_6   g03476(.A(new_n3852), .B(new_n3761), .Y(new_n3853));
  nand_5 g03477(.A(new_n3853), .B(new_n3851), .Y(new_n3854));
  xor_4  g03478(.A(new_n3854), .B(new_n3848), .Y(new_n3855));
  xor_4  g03479(.A(new_n3855), .B(new_n3845), .Y(new_n3856));
  not_8  g03480(.A(new_n3767), .Y(new_n3857));
  nand_5 g03481(.A(new_n3770), .B(new_n3857), .Y(new_n3858));
  or_6   g03482(.A(new_n3771), .B(new_n3766), .Y(new_n3859));
  nand_5 g03483(.A(new_n3859), .B(new_n3858), .Y(new_n3860));
  xor_4  g03484(.A(new_n3860), .B(new_n3856), .Y(new_n3861));
  xor_4  g03485(.A(new_n3861), .B(new_n3833), .Y(new_n3862));
  xor_4  g03486(.A(new_n3862), .B(new_n3832), .Y(new_n3863));
  nand_5 g03487(.A(pi173), .B(pi001), .Y(new_n3864));
  nand_5 g03488(.A(new_n3782), .B(new_n3781), .Y(new_n3865));
  nand_5 g03489(.A(new_n3783), .B(new_n3780), .Y(new_n3866));
  nand_5 g03490(.A(new_n3866), .B(new_n3865), .Y(new_n3867));
  xor_4  g03491(.A(new_n3867), .B(new_n3864), .Y(new_n3868));
  nand_5 g03492(.A(pi122), .B(pi014), .Y(new_n3869));
  nand_5 g03493(.A(pi135), .B(pi109), .Y(new_n3870));
  nand_5 g03494(.A(new_n3870), .B(new_n3869), .Y(new_n3871));
  nand_5 g03495(.A(pi135), .B(pi014), .Y(new_n3872));
  nor_5  g03496(.A(new_n3872), .B(new_n3782), .Y(new_n3873));
  not_8  g03497(.A(new_n3873), .Y(new_n3874));
  nand_5 g03498(.A(new_n3874), .B(new_n3871), .Y(new_n3875));
  xor_4  g03499(.A(new_n3875), .B(new_n3868), .Y(new_n3876));
  nand_5 g03500(.A(pi230), .B(pi102), .Y(new_n3877));
  nand_5 g03501(.A(pi219), .B(pi050), .Y(new_n3878));
  and_6  g03502(.A(new_n3878), .B(new_n3877), .Y(new_n3879));
  nand_5 g03503(.A(pi102), .B(pi050), .Y(new_n3880));
  nor_5  g03504(.A(new_n3880), .B(new_n3785), .Y(new_n3881));
  or_6   g03505(.A(new_n3881), .B(new_n3879), .Y(new_n3882));
  xnor_4 g03506(.A(new_n3882), .B(new_n3876), .Y(new_n3883));
  nand_5 g03507(.A(new_n3788), .B(new_n3785), .Y(new_n3884));
  nand_5 g03508(.A(new_n3789), .B(new_n3784), .Y(new_n3885));
  nand_5 g03509(.A(new_n3885), .B(new_n3884), .Y(new_n3886));
  xor_4  g03510(.A(new_n3886), .B(new_n3883), .Y(new_n3887));
  not_8  g03511(.A(new_n3775), .Y(new_n3888));
  nand_5 g03512(.A(new_n3778), .B(new_n3888), .Y(new_n3889));
  or_6   g03513(.A(new_n3790), .B(new_n3779), .Y(new_n3890));
  nand_5 g03514(.A(new_n3890), .B(new_n3889), .Y(new_n3891));
  xnor_4 g03515(.A(new_n3891), .B(new_n3887), .Y(new_n3892));
  nand_5 g03516(.A(new_n3791), .B(new_n3774), .Y(new_n3893));
  nand_5 g03517(.A(pi253), .B(pi087), .Y(new_n3894));
  xor_4  g03518(.A(new_n3894), .B(new_n3893), .Y(new_n3895));
  xor_4  g03519(.A(new_n3895), .B(new_n3892), .Y(new_n3896));
  xor_4  g03520(.A(new_n3896), .B(new_n3863), .Y(new_n3897));
  xor_4  g03521(.A(new_n3897), .B(new_n3831), .Y(new_n3898));
  nand_5 g03522(.A(new_n3815), .B(new_n3798), .Y(new_n3899));
  nand_5 g03523(.A(pi195), .B(pi138), .Y(new_n3900));
  nand_5 g03524(.A(pi216), .B(pi058), .Y(new_n3901));
  nand_5 g03525(.A(pi186), .B(pi076), .Y(new_n3902));
  nand_5 g03526(.A(pi132), .B(pi079), .Y(new_n3903));
  nand_5 g03527(.A(new_n3903), .B(new_n3902), .Y(new_n3904));
  nand_5 g03528(.A(pi186), .B(pi079), .Y(new_n3905));
  or_6   g03529(.A(new_n3905), .B(new_n3799), .Y(new_n3906));
  nand_5 g03530(.A(new_n3906), .B(new_n3904), .Y(new_n3907));
  xor_4  g03531(.A(new_n3907), .B(new_n3901), .Y(new_n3908));
  nand_5 g03532(.A(new_n3801), .B(new_n3800), .Y(new_n3909));
  nand_5 g03533(.A(new_n3802), .B(new_n3799), .Y(new_n3910));
  nand_5 g03534(.A(new_n3910), .B(new_n3909), .Y(new_n3911));
  xor_4  g03535(.A(new_n3911), .B(new_n3908), .Y(new_n3912));
  nand_5 g03536(.A(pi211), .B(pi041), .Y(new_n3913));
  nand_5 g03537(.A(pi199), .B(pi182), .Y(new_n3914));
  nand_5 g03538(.A(new_n3914), .B(new_n3913), .Y(new_n3915));
  nand_5 g03539(.A(pi199), .B(pi041), .Y(new_n3916));
  nor_5  g03540(.A(new_n3916), .B(new_n3804), .Y(new_n3917));
  not_8  g03541(.A(new_n3917), .Y(new_n3918));
  nand_5 g03542(.A(new_n3918), .B(new_n3915), .Y(new_n3919));
  xnor_4 g03543(.A(new_n3919), .B(new_n3912), .Y(new_n3920));
  nand_5 g03544(.A(new_n3807), .B(new_n3804), .Y(new_n3921));
  nand_5 g03545(.A(new_n3808), .B(new_n3803), .Y(new_n3922));
  nand_5 g03546(.A(new_n3922), .B(new_n3921), .Y(new_n3923));
  xor_4  g03547(.A(new_n3923), .B(new_n3920), .Y(new_n3924));
  not_8  g03548(.A(new_n3810), .Y(new_n3925));
  nand_5 g03549(.A(new_n3813), .B(new_n3925), .Y(new_n3926));
  or_6   g03550(.A(new_n3814), .B(new_n3809), .Y(new_n3927));
  nand_5 g03551(.A(new_n3927), .B(new_n3926), .Y(new_n3928));
  xnor_4 g03552(.A(new_n3928), .B(new_n3924), .Y(new_n3929));
  xor_4  g03553(.A(new_n3929), .B(new_n3900), .Y(new_n3930));
  not_8  g03554(.A(new_n3930), .Y(new_n3931));
  xor_4  g03555(.A(new_n3931), .B(new_n3899), .Y(new_n3932));
  nand_5 g03556(.A(new_n3820), .B(new_n3816), .Y(new_n3933));
  nand_5 g03557(.A(new_n3821), .B(new_n3797), .Y(new_n3934));
  nand_5 g03558(.A(new_n3934), .B(new_n3933), .Y(new_n3935));
  xor_4  g03559(.A(new_n3935), .B(new_n3932), .Y(new_n3936));
  xor_4  g03560(.A(new_n3936), .B(new_n3898), .Y(new_n3937));
  xor_4  g03561(.A(new_n3827), .B(new_n3826), .Y(new_n3938));
  nand_5 g03562(.A(new_n3938), .B(new_n3937), .Y(new_n3939));
  nand_5 g03563(.A(new_n3939), .B(new_n3828), .Y(new_n3940));
  nand_5 g03564(.A(new_n3940), .B(new_n3621), .Y(new_n3941));
  not_8  g03565(.A(new_n3856), .Y(new_n3942));
  nand_5 g03566(.A(new_n3860), .B(new_n3942), .Y(new_n3943));
  nand_5 g03567(.A(pi099), .B(pi066), .Y(new_n3944));
  nand_5 g03568(.A(pi226), .B(pi155), .Y(new_n3945));
  xor_4  g03569(.A(new_n3945), .B(new_n3838), .Y(new_n3946));
  xor_4  g03570(.A(new_n3946), .B(new_n3944), .Y(new_n3947));
  nand_5 g03571(.A(pi123), .B(pi055), .Y(new_n3948));
  xor_4  g03572(.A(new_n3948), .B(new_n3839), .Y(new_n3949));
  xor_4  g03573(.A(new_n3949), .B(new_n3947), .Y(new_n3950));
  nand_5 g03574(.A(pi071), .B(pi025), .Y(new_n3951));
  nand_5 g03575(.A(pi239), .B(pi142), .Y(new_n3952));
  xor_4  g03576(.A(new_n3952), .B(new_n3951), .Y(new_n3953));
  xor_4  g03577(.A(new_n3953), .B(new_n3852), .Y(new_n3954));
  nand_5 g03578(.A(new_n3840), .B(new_n3834), .Y(new_n3955));
  nand_5 g03579(.A(new_n3844), .B(new_n3841), .Y(new_n3956));
  nand_5 g03580(.A(new_n3956), .B(new_n3955), .Y(new_n3957));
  xor_4  g03581(.A(new_n3957), .B(new_n3954), .Y(new_n3958));
  xor_4  g03582(.A(new_n3958), .B(new_n3950), .Y(new_n3959));
  nand_5 g03583(.A(new_n3854), .B(new_n3848), .Y(new_n3960));
  nand_5 g03584(.A(new_n3855), .B(new_n3845), .Y(new_n3961));
  nand_5 g03585(.A(new_n3961), .B(new_n3960), .Y(new_n3962));
  xor_4  g03586(.A(new_n3962), .B(new_n3853), .Y(new_n3963));
  xor_4  g03587(.A(new_n3963), .B(new_n3959), .Y(new_n3964));
  xor_4  g03588(.A(new_n3964), .B(new_n3943), .Y(new_n3965));
  or_6   g03589(.A(new_n3861), .B(new_n3833), .Y(new_n3966));
  nand_5 g03590(.A(new_n3862), .B(new_n3832), .Y(new_n3967));
  nand_5 g03591(.A(new_n3967), .B(new_n3966), .Y(new_n3968));
  xor_4  g03592(.A(new_n3968), .B(new_n3965), .Y(new_n3969));
  nand_5 g03593(.A(new_n3891), .B(new_n3887), .Y(new_n3970));
  nand_5 g03594(.A(pi173), .B(pi122), .Y(new_n3971));
  nand_5 g03595(.A(pi109), .B(pi059), .Y(new_n3972));
  xor_4  g03596(.A(new_n3972), .B(new_n3971), .Y(new_n3973));
  xor_4  g03597(.A(new_n3973), .B(new_n3872), .Y(new_n3974));
  nand_5 g03598(.A(pi230), .B(pi001), .Y(new_n3975));
  xor_4  g03599(.A(new_n3975), .B(new_n3874), .Y(new_n3976));
  not_8  g03600(.A(new_n3976), .Y(new_n3977));
  xor_4  g03601(.A(new_n3977), .B(new_n3974), .Y(new_n3978));
  nand_5 g03602(.A(pi087), .B(pi074), .Y(new_n3979));
  nand_5 g03603(.A(pi253), .B(pi219), .Y(new_n3980));
  xor_4  g03604(.A(new_n3980), .B(new_n3979), .Y(new_n3981));
  xor_4  g03605(.A(new_n3981), .B(new_n3880), .Y(new_n3982));
  nand_5 g03606(.A(new_n3867), .B(new_n3864), .Y(new_n3983));
  nand_5 g03607(.A(new_n3875), .B(new_n3868), .Y(new_n3984));
  nand_5 g03608(.A(new_n3984), .B(new_n3983), .Y(new_n3985));
  xor_4  g03609(.A(new_n3985), .B(new_n3982), .Y(new_n3986));
  xor_4  g03610(.A(new_n3986), .B(new_n3978), .Y(new_n3987));
  nor_5  g03611(.A(new_n3882), .B(new_n3876), .Y(new_n3988));
  nor_5  g03612(.A(new_n3886), .B(new_n3883), .Y(new_n3989));
  xor_4  g03613(.A(new_n3989), .B(new_n3881), .Y(new_n3990));
  nor_5  g03614(.A(new_n3990), .B(new_n3988), .Y(new_n3991));
  not_8  g03615(.A(new_n3991), .Y(new_n3992));
  xor_4  g03616(.A(new_n3992), .B(new_n3987), .Y(new_n3993));
  xor_4  g03617(.A(new_n3993), .B(new_n3970), .Y(new_n3994));
  nand_5 g03618(.A(new_n3894), .B(new_n3893), .Y(new_n3995));
  nand_5 g03619(.A(new_n3895), .B(new_n3892), .Y(new_n3996));
  nand_5 g03620(.A(new_n3996), .B(new_n3995), .Y(new_n3997));
  xor_4  g03621(.A(new_n3997), .B(new_n3994), .Y(new_n3998));
  xor_4  g03622(.A(new_n3998), .B(new_n3969), .Y(new_n3999));
  not_8  g03623(.A(new_n3863), .Y(new_n4000));
  nor_5  g03624(.A(new_n3896), .B(new_n4000), .Y(new_n4001));
  nor_5  g03625(.A(new_n3897), .B(new_n3831), .Y(new_n4002));
  nor_5  g03626(.A(new_n4002), .B(new_n4001), .Y(new_n4003));
  not_8  g03627(.A(new_n4003), .Y(new_n4004));
  xor_4  g03628(.A(new_n4004), .B(new_n3999), .Y(new_n4005));
  nand_5 g03629(.A(new_n3928), .B(new_n3924), .Y(new_n4006));
  nand_5 g03630(.A(pi251), .B(pi132), .Y(new_n4007));
  nand_5 g03631(.A(pi076), .B(pi058), .Y(new_n4008));
  xor_4  g03632(.A(new_n4008), .B(new_n3905), .Y(new_n4009));
  xor_4  g03633(.A(new_n4009), .B(new_n4007), .Y(new_n4010));
  nand_5 g03634(.A(pi216), .B(pi211), .Y(new_n4011));
  xor_4  g03635(.A(new_n4011), .B(new_n3906), .Y(new_n4012));
  not_8  g03636(.A(new_n4012), .Y(new_n4013));
  xor_4  g03637(.A(new_n4013), .B(new_n4010), .Y(new_n4014));
  nand_5 g03638(.A(pi218), .B(pi138), .Y(new_n4015));
  nand_5 g03639(.A(pi195), .B(pi182), .Y(new_n4016));
  xor_4  g03640(.A(new_n4016), .B(new_n4015), .Y(new_n4017));
  xor_4  g03641(.A(new_n4017), .B(new_n3916), .Y(new_n4018));
  nand_5 g03642(.A(new_n3907), .B(new_n3901), .Y(new_n4019));
  nand_5 g03643(.A(new_n3911), .B(new_n3908), .Y(new_n4020));
  nand_5 g03644(.A(new_n4020), .B(new_n4019), .Y(new_n4021));
  xor_4  g03645(.A(new_n4021), .B(new_n4018), .Y(new_n4022));
  xor_4  g03646(.A(new_n4022), .B(new_n4014), .Y(new_n4023));
  nor_5  g03647(.A(new_n3923), .B(new_n3920), .Y(new_n4024));
  and_6  g03648(.A(new_n4024), .B(new_n3917), .Y(new_n4025));
  or_6   g03649(.A(new_n3919), .B(new_n3912), .Y(new_n4026));
  nand_5 g03650(.A(new_n4026), .B(new_n3918), .Y(new_n4027));
  nor_5  g03651(.A(new_n4027), .B(new_n4024), .Y(new_n4028));
  or_6   g03652(.A(new_n4028), .B(new_n4025), .Y(new_n4029));
  xor_4  g03653(.A(new_n4029), .B(new_n4023), .Y(new_n4030));
  xor_4  g03654(.A(new_n4030), .B(new_n4006), .Y(new_n4031));
  nor_5  g03655(.A(new_n3929), .B(new_n3900), .Y(new_n4032));
  nor_5  g03656(.A(new_n3931), .B(new_n3899), .Y(new_n4033));
  or_6   g03657(.A(new_n4033), .B(new_n4032), .Y(new_n4034));
  xor_4  g03658(.A(new_n4034), .B(new_n4031), .Y(new_n4035));
  nand_5 g03659(.A(new_n3935), .B(new_n3932), .Y(new_n4036));
  nand_5 g03660(.A(new_n3936), .B(new_n3898), .Y(new_n4037));
  nand_5 g03661(.A(new_n4037), .B(new_n4036), .Y(new_n4038));
  xor_4  g03662(.A(new_n4038), .B(new_n4035), .Y(new_n4039));
  xor_4  g03663(.A(new_n4039), .B(new_n4005), .Y(new_n4040));
  xor_4  g03664(.A(new_n3940), .B(new_n3621), .Y(new_n4041));
  nand_5 g03665(.A(new_n4041), .B(new_n4040), .Y(new_n4042));
  nand_5 g03666(.A(new_n4042), .B(new_n3941), .Y(new_n4043));
  or_6   g03667(.A(new_n4038), .B(new_n4035), .Y(new_n4044));
  not_8  g03668(.A(new_n4005), .Y(new_n4045));
  nand_5 g03669(.A(new_n4039), .B(new_n4045), .Y(new_n4046));
  nand_5 g03670(.A(new_n4046), .B(new_n4044), .Y(new_n4047));
  nand_5 g03671(.A(new_n3998), .B(new_n3969), .Y(new_n4048));
  nand_5 g03672(.A(new_n4004), .B(new_n3999), .Y(new_n4049));
  nand_5 g03673(.A(new_n4049), .B(new_n4048), .Y(new_n4050));
  nor_5  g03674(.A(new_n4029), .B(new_n4023), .Y(new_n4051));
  nor_5  g03675(.A(new_n4051), .B(new_n4028), .Y(new_n4052));
  nand_5 g03676(.A(pi138), .B(pi037), .Y(new_n4053));
  xor_4  g03677(.A(new_n4053), .B(new_n4052), .Y(new_n4054));
  xor_4  g03678(.A(new_n4054), .B(new_n4050), .Y(new_n4055));
  nand_5 g03679(.A(new_n3594), .B(new_n3591), .Y(new_n4056));
  nand_5 g03680(.A(new_n3595), .B(new_n3587), .Y(new_n4057));
  nand_5 g03681(.A(new_n4057), .B(new_n4056), .Y(new_n4058));
  nand_5 g03682(.A(new_n3589), .B(new_n3588), .Y(new_n4059));
  nand_5 g03683(.A(new_n3590), .B(new_n3542), .Y(new_n4060));
  nand_5 g03684(.A(new_n4060), .B(new_n4059), .Y(new_n4061));
  xor_4  g03685(.A(new_n4061), .B(new_n4058), .Y(new_n4062));
  nand_5 g03686(.A(pi177), .B(pi069), .Y(new_n4063));
  nand_5 g03687(.A(pi150), .B(pi101), .Y(new_n4064));
  nand_5 g03688(.A(pi223), .B(pi221), .Y(new_n4065));
  xor_4  g03689(.A(new_n4065), .B(new_n4064), .Y(new_n4066));
  xor_4  g03690(.A(new_n4066), .B(new_n4063), .Y(new_n4067));
  xor_4  g03691(.A(new_n4067), .B(new_n4062), .Y(new_n4068));
  or_6   g03692(.A(new_n4030), .B(new_n4006), .Y(new_n4069));
  nand_5 g03693(.A(new_n4034), .B(new_n4031), .Y(new_n4070));
  nand_5 g03694(.A(new_n4070), .B(new_n4069), .Y(new_n4071));
  nand_5 g03695(.A(pi196), .B(pi060), .Y(new_n4072));
  nand_5 g03696(.A(pi244), .B(pi225), .Y(new_n4073));
  xor_4  g03697(.A(new_n4073), .B(new_n4072), .Y(new_n4074));
  xor_4  g03698(.A(new_n4074), .B(new_n4071), .Y(new_n4075));
  xor_4  g03699(.A(new_n4075), .B(new_n4068), .Y(new_n4076));
  nand_5 g03700(.A(pi184), .B(pi020), .Y(new_n4077));
  nand_5 g03701(.A(new_n3582), .B(new_n3581), .Y(new_n4078));
  nand_5 g03702(.A(new_n3583), .B(new_n3527), .Y(new_n4079));
  nand_5 g03703(.A(new_n4079), .B(new_n4078), .Y(new_n4080));
  xor_4  g03704(.A(new_n4080), .B(new_n4077), .Y(new_n4081));
  nand_5 g03705(.A(pi192), .B(pi132), .Y(new_n4082));
  nand_5 g03706(.A(pi251), .B(pi186), .Y(new_n4083));
  xor_4  g03707(.A(new_n4083), .B(new_n4082), .Y(new_n4084));
  xor_4  g03708(.A(new_n4084), .B(new_n4081), .Y(new_n4085));
  xor_4  g03709(.A(new_n4085), .B(new_n4076), .Y(new_n4086));
  xor_4  g03710(.A(new_n4086), .B(new_n4055), .Y(new_n4087));
  nand_5 g03711(.A(pi195), .B(pi041), .Y(new_n4088));
  nand_5 g03712(.A(pi211), .B(pi076), .Y(new_n4089));
  or_6   g03713(.A(new_n4021), .B(new_n4018), .Y(new_n4090));
  nand_5 g03714(.A(new_n4022), .B(new_n4014), .Y(new_n4091));
  nand_5 g03715(.A(new_n4091), .B(new_n4090), .Y(new_n4092));
  xor_4  g03716(.A(new_n4092), .B(new_n4089), .Y(new_n4093));
  xor_4  g03717(.A(new_n4093), .B(new_n4088), .Y(new_n4094));
  xor_4  g03718(.A(new_n4094), .B(new_n4087), .Y(new_n4095));
  nand_5 g03719(.A(new_n3962), .B(new_n3853), .Y(new_n4096));
  nand_5 g03720(.A(new_n3963), .B(new_n3959), .Y(new_n4097));
  nand_5 g03721(.A(new_n4097), .B(new_n4096), .Y(new_n4098));
  nand_5 g03722(.A(pi226), .B(pi086), .Y(new_n4099));
  nand_5 g03723(.A(new_n4016), .B(new_n4015), .Y(new_n4100));
  nand_5 g03724(.A(new_n4017), .B(new_n3916), .Y(new_n4101));
  nand_5 g03725(.A(new_n4101), .B(new_n4100), .Y(new_n4102));
  nand_5 g03726(.A(pi207), .B(pi155), .Y(new_n4103));
  nand_5 g03727(.A(pi066), .B(pi023), .Y(new_n4104));
  xnor_4 g03728(.A(new_n4104), .B(new_n4103), .Y(new_n4105));
  xor_4  g03729(.A(new_n4105), .B(new_n4102), .Y(new_n4106));
  xor_4  g03730(.A(new_n4106), .B(new_n4099), .Y(new_n4107));
  xor_4  g03731(.A(new_n4107), .B(new_n4098), .Y(new_n4108));
  nor_5  g03732(.A(new_n4011), .B(new_n3906), .Y(new_n4109));
  nor_5  g03733(.A(new_n4013), .B(new_n4010), .Y(new_n4110));
  or_6   g03734(.A(new_n4110), .B(new_n4109), .Y(new_n4111));
  or_6   g03735(.A(new_n3964), .B(new_n3943), .Y(new_n4112));
  nand_5 g03736(.A(new_n3968), .B(new_n3965), .Y(new_n4113));
  nand_5 g03737(.A(new_n4113), .B(new_n4112), .Y(new_n4114));
  nand_5 g03738(.A(pi243), .B(pi142), .Y(new_n4115));
  xor_4  g03739(.A(new_n4115), .B(new_n4114), .Y(new_n4116));
  xor_4  g03740(.A(new_n4116), .B(new_n4111), .Y(new_n4117));
  xor_4  g03741(.A(new_n4117), .B(new_n4108), .Y(new_n4118));
  nand_5 g03742(.A(pi218), .B(pi182), .Y(new_n4119));
  nand_5 g03743(.A(new_n4008), .B(new_n3905), .Y(new_n4120));
  nand_5 g03744(.A(new_n4009), .B(new_n4007), .Y(new_n4121));
  nand_5 g03745(.A(new_n4121), .B(new_n4120), .Y(new_n4122));
  xor_4  g03746(.A(new_n4122), .B(new_n4119), .Y(new_n4123));
  nand_5 g03747(.A(pi079), .B(pi058), .Y(new_n4124));
  nand_5 g03748(.A(pi216), .B(pi199), .Y(new_n4125));
  xor_4  g03749(.A(new_n4125), .B(new_n4124), .Y(new_n4126));
  xor_4  g03750(.A(new_n4126), .B(new_n4123), .Y(new_n4127));
  xor_4  g03751(.A(new_n4127), .B(new_n4118), .Y(new_n4128));
  xor_4  g03752(.A(new_n4128), .B(new_n4095), .Y(new_n4129));
  nand_5 g03753(.A(new_n3989), .B(new_n3881), .Y(new_n4130));
  nand_5 g03754(.A(new_n3992), .B(new_n3987), .Y(new_n4131));
  nand_5 g03755(.A(new_n4131), .B(new_n4130), .Y(new_n4132));
  nand_5 g03756(.A(pi059), .B(pi014), .Y(new_n4133));
  nand_5 g03757(.A(pi173), .B(pi135), .Y(new_n4134));
  xor_4  g03758(.A(new_n4134), .B(new_n4133), .Y(new_n4135));
  xor_4  g03759(.A(new_n4135), .B(new_n4132), .Y(new_n4136));
  xor_4  g03760(.A(new_n4136), .B(new_n4129), .Y(new_n4137));
  xor_4  g03761(.A(new_n4137), .B(new_n4047), .Y(new_n4138));
  xor_4  g03762(.A(new_n4138), .B(new_n4043), .Y(new_n4139));
  nor_5  g03763(.A(new_n3603), .B(new_n3580), .Y(new_n4140));
  nor_5  g03764(.A(new_n3620), .B(new_n3604), .Y(new_n4141));
  nor_5  g03765(.A(new_n4141), .B(new_n4140), .Y(new_n4142));
  or_6   g03766(.A(new_n3585), .B(new_n3528), .Y(new_n4143));
  not_8  g03767(.A(new_n3584), .Y(new_n4144));
  nand_5 g03768(.A(new_n3586), .B(new_n4144), .Y(new_n4145));
  nand_5 g03769(.A(new_n4145), .B(new_n4143), .Y(new_n4146));
  nand_5 g03770(.A(pi230), .B(pi122), .Y(new_n4147));
  nand_5 g03771(.A(pi050), .B(pi001), .Y(new_n4148));
  xor_4  g03772(.A(new_n4148), .B(new_n4147), .Y(new_n4149));
  nand_5 g03773(.A(new_n3945), .B(new_n3838), .Y(new_n4150));
  nand_5 g03774(.A(new_n3946), .B(new_n3944), .Y(new_n4151));
  nand_5 g03775(.A(new_n4151), .B(new_n4150), .Y(new_n4152));
  nand_5 g03776(.A(pi099), .B(pi055), .Y(new_n4153));
  nand_5 g03777(.A(pi123), .B(pi002), .Y(new_n4154));
  xor_4  g03778(.A(new_n4154), .B(new_n4153), .Y(new_n4155));
  xor_4  g03779(.A(new_n4155), .B(new_n4152), .Y(new_n4156));
  nand_5 g03780(.A(pi239), .B(pi071), .Y(new_n4157));
  nand_5 g03781(.A(pi169), .B(pi025), .Y(new_n4158));
  xnor_4 g03782(.A(new_n4158), .B(new_n4157), .Y(new_n4159));
  or_6   g03783(.A(new_n3948), .B(new_n3839), .Y(new_n4160));
  not_8  g03784(.A(new_n3947), .Y(new_n4161));
  nand_5 g03785(.A(new_n3949), .B(new_n4161), .Y(new_n4162));
  nand_5 g03786(.A(new_n4162), .B(new_n4160), .Y(new_n4163));
  xor_4  g03787(.A(new_n4163), .B(new_n4159), .Y(new_n4164));
  nand_5 g03788(.A(new_n3952), .B(new_n3951), .Y(new_n4165));
  nand_5 g03789(.A(new_n3953), .B(new_n3852), .Y(new_n4166));
  nand_5 g03790(.A(new_n4166), .B(new_n4165), .Y(new_n4167));
  nand_5 g03791(.A(new_n3957), .B(new_n3954), .Y(new_n4168));
  nand_5 g03792(.A(new_n3958), .B(new_n3950), .Y(new_n4169));
  nand_5 g03793(.A(new_n4169), .B(new_n4168), .Y(new_n4170));
  xor_4  g03794(.A(new_n4170), .B(new_n4167), .Y(new_n4171));
  xor_4  g03795(.A(new_n4171), .B(new_n4164), .Y(new_n4172));
  xor_4  g03796(.A(new_n4172), .B(new_n4156), .Y(new_n4173));
  xor_4  g03797(.A(new_n4173), .B(new_n4149), .Y(new_n4174));
  not_8  g03798(.A(new_n3993), .Y(new_n4175));
  nor_5  g03799(.A(new_n4175), .B(new_n3970), .Y(new_n4176));
  nor_5  g03800(.A(new_n3997), .B(new_n3994), .Y(new_n4177));
  nor_5  g03801(.A(new_n4177), .B(new_n4176), .Y(new_n4178));
  nand_5 g03802(.A(pi205), .B(pi087), .Y(new_n4179));
  xor_4  g03803(.A(new_n4179), .B(new_n4178), .Y(new_n4180));
  xor_4  g03804(.A(new_n4180), .B(new_n4174), .Y(new_n4181));
  nand_5 g03805(.A(pi109), .B(pi094), .Y(new_n4182));
  nand_5 g03806(.A(pi137), .B(pi029), .Y(new_n4183));
  nand_5 g03807(.A(pi160), .B(pi010), .Y(new_n4184));
  xor_4  g03808(.A(new_n4184), .B(new_n4183), .Y(new_n4185));
  nand_5 g03809(.A(new_n3980), .B(new_n3979), .Y(new_n4186));
  nand_5 g03810(.A(new_n3981), .B(new_n3880), .Y(new_n4187));
  nand_5 g03811(.A(new_n4187), .B(new_n4186), .Y(new_n4188));
  nor_5  g03812(.A(new_n3975), .B(new_n3874), .Y(new_n4189));
  nor_5  g03813(.A(new_n3977), .B(new_n3974), .Y(new_n4190));
  or_6   g03814(.A(new_n4190), .B(new_n4189), .Y(new_n4191));
  xor_4  g03815(.A(new_n4191), .B(new_n4188), .Y(new_n4192));
  xor_4  g03816(.A(new_n4192), .B(new_n4185), .Y(new_n4193));
  nor_5  g03817(.A(new_n3602), .B(new_n3596), .Y(new_n4194));
  nor_5  g03818(.A(new_n4194), .B(new_n3601), .Y(new_n4195));
  nand_5 g03819(.A(new_n3972), .B(new_n3971), .Y(new_n4196));
  nand_5 g03820(.A(new_n3973), .B(new_n3872), .Y(new_n4197));
  nand_5 g03821(.A(new_n4197), .B(new_n4196), .Y(new_n4198));
  nand_5 g03822(.A(pi219), .B(pi074), .Y(new_n4199));
  nand_5 g03823(.A(pi253), .B(pi102), .Y(new_n4200));
  xor_4  g03824(.A(new_n4200), .B(new_n4199), .Y(new_n4201));
  or_6   g03825(.A(new_n3985), .B(new_n3982), .Y(new_n4202));
  nand_5 g03826(.A(new_n3986), .B(new_n3978), .Y(new_n4203));
  nand_5 g03827(.A(new_n4203), .B(new_n4202), .Y(new_n4204));
  xor_4  g03828(.A(new_n4204), .B(new_n4201), .Y(new_n4205));
  xor_4  g03829(.A(new_n4205), .B(new_n4198), .Y(new_n4206));
  xor_4  g03830(.A(new_n4206), .B(new_n4195), .Y(new_n4207));
  xor_4  g03831(.A(new_n4207), .B(new_n4193), .Y(new_n4208));
  xor_4  g03832(.A(new_n4208), .B(new_n4182), .Y(new_n4209));
  xor_4  g03833(.A(new_n4209), .B(new_n4181), .Y(new_n4210));
  xor_4  g03834(.A(new_n4210), .B(new_n4146), .Y(new_n4211));
  xor_4  g03835(.A(new_n4211), .B(new_n4142), .Y(new_n4212));
  xor_4  g03836(.A(new_n4212), .B(new_n4139), .Y(po013));
  nor_5  g03837(.A(new_n924), .B(new_n913), .Y(new_n4214));
  nand_5 g03838(.A(pi108), .B(pi049), .Y(new_n4215));
  nand_5 g03839(.A(pi245), .B(pi042), .Y(new_n4216));
  nand_5 g03840(.A(pi201), .B(pi051), .Y(new_n4217));
  xor_4  g03841(.A(new_n4217), .B(new_n4216), .Y(new_n4218));
  xor_4  g03842(.A(new_n4218), .B(new_n4215), .Y(new_n4219));
  nand_5 g03843(.A(pi171), .B(pi007), .Y(new_n4220));
  nand_5 g03844(.A(new_n921), .B(new_n920), .Y(new_n4221));
  nand_5 g03845(.A(new_n922), .B(new_n919), .Y(new_n4222));
  nand_5 g03846(.A(new_n4222), .B(new_n4221), .Y(new_n4223));
  xor_4  g03847(.A(new_n4223), .B(new_n4220), .Y(new_n4224));
  xor_4  g03848(.A(new_n4224), .B(new_n4219), .Y(new_n4225));
  nand_5 g03849(.A(pi118), .B(pi107), .Y(new_n4226));
  or_6   g03850(.A(new_n917), .B(new_n914), .Y(new_n4227));
  not_8  g03851(.A(new_n923), .Y(new_n4228));
  nand_5 g03852(.A(new_n4228), .B(new_n918), .Y(new_n4229));
  nand_5 g03853(.A(new_n4229), .B(new_n4227), .Y(new_n4230));
  xor_4  g03854(.A(new_n4230), .B(new_n4226), .Y(new_n4231));
  xor_4  g03855(.A(new_n4231), .B(new_n4225), .Y(new_n4232));
  nand_5 g03856(.A(new_n4232), .B(new_n4214), .Y(new_n4233));
  nand_5 g03857(.A(pi113), .B(pi107), .Y(new_n4234));
  nand_5 g03858(.A(new_n4234), .B(new_n4233), .Y(new_n4235));
  nand_5 g03859(.A(pi245), .B(pi108), .Y(new_n4236));
  nand_5 g03860(.A(pi201), .B(pi042), .Y(new_n4237));
  nand_5 g03861(.A(pi156), .B(pi051), .Y(new_n4238));
  nand_5 g03862(.A(new_n4238), .B(new_n4237), .Y(new_n4239));
  nand_5 g03863(.A(pi156), .B(pi042), .Y(new_n4240));
  or_6   g03864(.A(new_n4240), .B(new_n4217), .Y(new_n4241));
  nand_5 g03865(.A(new_n4241), .B(new_n4239), .Y(new_n4242));
  xor_4  g03866(.A(new_n4242), .B(new_n4236), .Y(new_n4243));
  nand_5 g03867(.A(new_n4217), .B(new_n4216), .Y(new_n4244));
  nand_5 g03868(.A(new_n4218), .B(new_n4215), .Y(new_n4245));
  nand_5 g03869(.A(new_n4245), .B(new_n4244), .Y(new_n4246));
  xor_4  g03870(.A(new_n4246), .B(new_n4243), .Y(new_n4247));
  nand_5 g03871(.A(pi049), .B(pi007), .Y(new_n4248));
  nand_5 g03872(.A(pi171), .B(pi118), .Y(new_n4249));
  and_6  g03873(.A(new_n4249), .B(new_n4248), .Y(new_n4250));
  nand_5 g03874(.A(pi118), .B(pi049), .Y(new_n4251));
  nor_5  g03875(.A(new_n4251), .B(new_n4220), .Y(new_n4252));
  or_6   g03876(.A(new_n4252), .B(new_n4250), .Y(new_n4253));
  xnor_4 g03877(.A(new_n4253), .B(new_n4247), .Y(new_n4254));
  nand_5 g03878(.A(new_n4223), .B(new_n4220), .Y(new_n4255));
  nand_5 g03879(.A(new_n4224), .B(new_n4219), .Y(new_n4256));
  nand_5 g03880(.A(new_n4256), .B(new_n4255), .Y(new_n4257));
  xor_4  g03881(.A(new_n4257), .B(new_n4254), .Y(new_n4258));
  not_8  g03882(.A(new_n4226), .Y(new_n4259));
  nand_5 g03883(.A(new_n4230), .B(new_n4259), .Y(new_n4260));
  or_6   g03884(.A(new_n4231), .B(new_n4225), .Y(new_n4261));
  nand_5 g03885(.A(new_n4261), .B(new_n4260), .Y(new_n4262));
  xnor_4 g03886(.A(new_n4262), .B(new_n4258), .Y(new_n4263));
  xor_4  g03887(.A(new_n4234), .B(new_n4233), .Y(new_n4264));
  nand_5 g03888(.A(new_n4264), .B(new_n4263), .Y(new_n4265));
  nand_5 g03889(.A(new_n4265), .B(new_n4235), .Y(new_n4266));
  nand_5 g03890(.A(new_n4262), .B(new_n4258), .Y(new_n4267));
  nand_5 g03891(.A(pi063), .B(pi051), .Y(new_n4268));
  nand_5 g03892(.A(pi201), .B(pi108), .Y(new_n4269));
  xor_4  g03893(.A(new_n4269), .B(new_n4268), .Y(new_n4270));
  xor_4  g03894(.A(new_n4270), .B(new_n4240), .Y(new_n4271));
  not_8  g03895(.A(new_n4271), .Y(new_n4272));
  nand_5 g03896(.A(pi245), .B(pi007), .Y(new_n4273));
  xor_4  g03897(.A(new_n4273), .B(new_n4241), .Y(new_n4274));
  xor_4  g03898(.A(new_n4274), .B(new_n4272), .Y(new_n4275));
  nand_5 g03899(.A(pi107), .B(pi038), .Y(new_n4276));
  nand_5 g03900(.A(pi171), .B(pi113), .Y(new_n4277));
  xor_4  g03901(.A(new_n4277), .B(new_n4276), .Y(new_n4278));
  xor_4  g03902(.A(new_n4278), .B(new_n4251), .Y(new_n4279));
  nand_5 g03903(.A(new_n4242), .B(new_n4236), .Y(new_n4280));
  nand_5 g03904(.A(new_n4246), .B(new_n4243), .Y(new_n4281));
  nand_5 g03905(.A(new_n4281), .B(new_n4280), .Y(new_n4282));
  xor_4  g03906(.A(new_n4282), .B(new_n4279), .Y(new_n4283));
  xor_4  g03907(.A(new_n4283), .B(new_n4275), .Y(new_n4284));
  nor_5  g03908(.A(new_n4253), .B(new_n4247), .Y(new_n4285));
  nor_5  g03909(.A(new_n4257), .B(new_n4254), .Y(new_n4286));
  xor_4  g03910(.A(new_n4286), .B(new_n4252), .Y(new_n4287));
  nor_5  g03911(.A(new_n4287), .B(new_n4285), .Y(new_n4288));
  xor_4  g03912(.A(new_n4288), .B(new_n4284), .Y(new_n4289));
  xor_4  g03913(.A(new_n4289), .B(new_n4267), .Y(new_n4290));
  xor_4  g03914(.A(new_n4290), .B(new_n4266), .Y(new_n4291));
  nand_5 g03915(.A(pi061), .B(pi039), .Y(new_n4292));
  nand_5 g03916(.A(pi178), .B(pi116), .Y(new_n4293));
  nand_5 g03917(.A(pi188), .B(pi070), .Y(new_n4294));
  nand_5 g03918(.A(new_n4294), .B(new_n4293), .Y(new_n4295));
  nand_5 g03919(.A(pi188), .B(pi116), .Y(new_n4296));
  nand_5 g03920(.A(pi178), .B(pi070), .Y(new_n4297));
  or_6   g03921(.A(new_n4297), .B(new_n4296), .Y(new_n4298));
  nand_5 g03922(.A(new_n4298), .B(new_n4295), .Y(new_n4299));
  xor_4  g03923(.A(new_n4299), .B(new_n4292), .Y(new_n4300));
  nand_5 g03924(.A(pi178), .B(pi039), .Y(new_n4301));
  nand_5 g03925(.A(new_n4301), .B(new_n4296), .Y(new_n4302));
  nand_5 g03926(.A(pi228), .B(pi061), .Y(new_n4303));
  xor_4  g03927(.A(new_n4301), .B(new_n4296), .Y(new_n4304));
  nand_5 g03928(.A(new_n4304), .B(new_n4303), .Y(new_n4305));
  nand_5 g03929(.A(new_n4305), .B(new_n4302), .Y(new_n4306));
  xor_4  g03930(.A(new_n4306), .B(new_n4300), .Y(new_n4307));
  nand_5 g03931(.A(pi228), .B(pi012), .Y(new_n4308));
  nand_5 g03932(.A(pi148), .B(pi144), .Y(new_n4309));
  and_6  g03933(.A(new_n4309), .B(new_n4308), .Y(new_n4310));
  nand_5 g03934(.A(pi148), .B(pi012), .Y(new_n4311));
  nand_5 g03935(.A(pi228), .B(pi144), .Y(new_n4312));
  nor_5  g03936(.A(new_n4312), .B(new_n4311), .Y(new_n4313));
  or_6   g03937(.A(new_n4313), .B(new_n4310), .Y(new_n4314));
  xnor_4 g03938(.A(new_n4314), .B(new_n4307), .Y(new_n4315));
  nand_5 g03939(.A(new_n937), .B(new_n936), .Y(new_n4316));
  nand_5 g03940(.A(new_n938), .B(new_n935), .Y(new_n4317));
  nand_5 g03941(.A(new_n4317), .B(new_n4316), .Y(new_n4318));
  nand_5 g03942(.A(new_n4318), .B(new_n4311), .Y(new_n4319));
  xor_4  g03943(.A(new_n4304), .B(new_n4303), .Y(new_n4320));
  xor_4  g03944(.A(new_n4318), .B(new_n4311), .Y(new_n4321));
  nand_5 g03945(.A(new_n4321), .B(new_n4320), .Y(new_n4322));
  nand_5 g03946(.A(new_n4322), .B(new_n4319), .Y(new_n4323));
  xor_4  g03947(.A(new_n4323), .B(new_n4315), .Y(new_n4324));
  xor_4  g03948(.A(new_n4321), .B(new_n4320), .Y(new_n4325));
  nand_5 g03949(.A(pi163), .B(pi144), .Y(new_n4326));
  nor_5  g03950(.A(new_n4326), .B(new_n4325), .Y(new_n4327));
  xnor_4 g03951(.A(new_n4326), .B(new_n4325), .Y(new_n4328));
  nand_5 g03952(.A(new_n943), .B(new_n940), .Y(new_n4329));
  nand_5 g03953(.A(new_n944), .B(new_n939), .Y(new_n4330));
  nand_5 g03954(.A(new_n4330), .B(new_n4329), .Y(new_n4331));
  nor_5  g03955(.A(new_n4331), .B(new_n4328), .Y(new_n4332));
  nor_5  g03956(.A(new_n4332), .B(new_n4327), .Y(new_n4333));
  not_8  g03957(.A(new_n4333), .Y(new_n4334));
  nand_5 g03958(.A(new_n4334), .B(new_n4324), .Y(new_n4335));
  nand_5 g03959(.A(pi188), .B(pi115), .Y(new_n4336));
  nand_5 g03960(.A(pi116), .B(pi061), .Y(new_n4337));
  xor_4  g03961(.A(new_n4337), .B(new_n4336), .Y(new_n4338));
  xor_4  g03962(.A(new_n4338), .B(new_n4297), .Y(new_n4339));
  nand_5 g03963(.A(pi039), .B(pi012), .Y(new_n4340));
  xor_4  g03964(.A(new_n4340), .B(new_n4298), .Y(new_n4341));
  xor_4  g03965(.A(new_n4341), .B(new_n4339), .Y(new_n4342));
  nand_5 g03966(.A(pi148), .B(pi098), .Y(new_n4343));
  nand_5 g03967(.A(pi163), .B(pi043), .Y(new_n4344));
  xor_4  g03968(.A(new_n4344), .B(new_n4343), .Y(new_n4345));
  xor_4  g03969(.A(new_n4345), .B(new_n4312), .Y(new_n4346));
  nand_5 g03970(.A(new_n4299), .B(new_n4292), .Y(new_n4347));
  nand_5 g03971(.A(new_n4306), .B(new_n4300), .Y(new_n4348));
  nand_5 g03972(.A(new_n4348), .B(new_n4347), .Y(new_n4349));
  xor_4  g03973(.A(new_n4349), .B(new_n4346), .Y(new_n4350));
  xnor_4 g03974(.A(new_n4350), .B(new_n4342), .Y(new_n4351));
  nor_5  g03975(.A(new_n4314), .B(new_n4307), .Y(new_n4352));
  nor_5  g03976(.A(new_n4323), .B(new_n4315), .Y(new_n4353));
  xor_4  g03977(.A(new_n4353), .B(new_n4313), .Y(new_n4354));
  nor_5  g03978(.A(new_n4354), .B(new_n4352), .Y(new_n4355));
  not_8  g03979(.A(new_n4355), .Y(new_n4356));
  xor_4  g03980(.A(new_n4356), .B(new_n4351), .Y(new_n4357));
  xor_4  g03981(.A(new_n4357), .B(new_n4335), .Y(new_n4358));
  nand_5 g03982(.A(pi163), .B(pi098), .Y(new_n4359));
  xor_4  g03983(.A(new_n4333), .B(new_n4324), .Y(new_n4360));
  nand_5 g03984(.A(new_n4360), .B(new_n4359), .Y(new_n4361));
  nor_5  g03985(.A(new_n945), .B(new_n934), .Y(new_n4362));
  xor_4  g03986(.A(new_n4331), .B(new_n4328), .Y(new_n4363));
  nand_5 g03987(.A(new_n4363), .B(new_n4362), .Y(new_n4364));
  xor_4  g03988(.A(new_n4360), .B(new_n4359), .Y(new_n4365));
  nand_5 g03989(.A(new_n4365), .B(new_n4364), .Y(new_n4366));
  nand_5 g03990(.A(new_n4366), .B(new_n4361), .Y(new_n4367));
  xor_4  g03991(.A(new_n4367), .B(new_n4358), .Y(new_n4368));
  not_8  g03992(.A(new_n4368), .Y(new_n4369));
  xor_4  g03993(.A(new_n4369), .B(new_n4291), .Y(new_n4370));
  xor_4  g03994(.A(new_n4264), .B(new_n4263), .Y(new_n4371));
  xor_4  g03995(.A(new_n4365), .B(new_n4364), .Y(new_n4372));
  nor_5  g03996(.A(new_n4372), .B(new_n4371), .Y(new_n4373));
  xnor_4 g03997(.A(new_n4372), .B(new_n4371), .Y(new_n4374));
  xor_4  g03998(.A(new_n4232), .B(new_n4214), .Y(new_n4375));
  nand_5 g03999(.A(new_n946), .B(new_n925), .Y(new_n4376));
  nand_5 g04000(.A(new_n969), .B(new_n947), .Y(new_n4377));
  nand_5 g04001(.A(new_n4377), .B(new_n4376), .Y(new_n4378));
  or_6   g04002(.A(new_n4378), .B(new_n4375), .Y(new_n4379));
  xnor_4 g04003(.A(new_n4363), .B(new_n4362), .Y(new_n4380));
  xor_4  g04004(.A(new_n4378), .B(new_n4375), .Y(new_n4381));
  nand_5 g04005(.A(new_n4381), .B(new_n4380), .Y(new_n4382));
  nand_5 g04006(.A(new_n4382), .B(new_n4379), .Y(new_n4383));
  nor_5  g04007(.A(new_n4383), .B(new_n4374), .Y(new_n4384));
  nor_5  g04008(.A(new_n4384), .B(new_n4373), .Y(new_n4385));
  xnor_4 g04009(.A(new_n4385), .B(new_n4370), .Y(new_n4386));
  nand_5 g04010(.A(pi179), .B(pi149), .Y(new_n4387));
  nand_5 g04011(.A(pi240), .B(pi179), .Y(new_n4388));
  nand_5 g04012(.A(pi149), .B(pi033), .Y(new_n4389));
  nand_5 g04013(.A(new_n4389), .B(new_n4388), .Y(new_n4390));
  nand_5 g04014(.A(pi167), .B(pi162), .Y(new_n4391));
  xor_4  g04015(.A(new_n4389), .B(new_n4388), .Y(new_n4392));
  nand_5 g04016(.A(new_n4392), .B(new_n4391), .Y(new_n4393));
  nand_5 g04017(.A(new_n4393), .B(new_n4390), .Y(new_n4394));
  xnor_4 g04018(.A(new_n4394), .B(new_n4387), .Y(new_n4395));
  nand_5 g04019(.A(pi167), .B(pi033), .Y(new_n4396));
  nand_5 g04020(.A(pi181), .B(pi162), .Y(new_n4397));
  nand_5 g04021(.A(new_n4397), .B(new_n4396), .Y(new_n4398));
  nand_5 g04022(.A(pi181), .B(pi033), .Y(new_n4399));
  or_6   g04023(.A(new_n4399), .B(new_n4391), .Y(new_n4400));
  nand_5 g04024(.A(new_n4400), .B(new_n4398), .Y(new_n4401));
  xnor_4 g04025(.A(new_n4401), .B(new_n4395), .Y(new_n4402));
  nand_5 g04026(.A(pi240), .B(pi048), .Y(new_n4403));
  nand_5 g04027(.A(pi237), .B(pi134), .Y(new_n4404));
  and_6  g04028(.A(new_n4404), .B(new_n4403), .Y(new_n4405));
  nand_5 g04029(.A(pi134), .B(pi048), .Y(new_n4406));
  nand_5 g04030(.A(pi240), .B(pi237), .Y(new_n4407));
  nor_5  g04031(.A(new_n4407), .B(new_n4406), .Y(new_n4408));
  or_6   g04032(.A(new_n4408), .B(new_n4405), .Y(new_n4409));
  xnor_4 g04033(.A(new_n4409), .B(new_n4402), .Y(new_n4410));
  nand_5 g04034(.A(new_n982), .B(new_n981), .Y(new_n4411));
  nand_5 g04035(.A(new_n983), .B(new_n980), .Y(new_n4412));
  nand_5 g04036(.A(new_n4412), .B(new_n4411), .Y(new_n4413));
  nand_5 g04037(.A(new_n4413), .B(new_n4406), .Y(new_n4414));
  xor_4  g04038(.A(new_n4392), .B(new_n4391), .Y(new_n4415));
  xor_4  g04039(.A(new_n4413), .B(new_n4406), .Y(new_n4416));
  nand_5 g04040(.A(new_n4416), .B(new_n4415), .Y(new_n4417));
  nand_5 g04041(.A(new_n4417), .B(new_n4414), .Y(new_n4418));
  xor_4  g04042(.A(new_n4418), .B(new_n4410), .Y(new_n4419));
  nand_5 g04043(.A(pi237), .B(pi175), .Y(new_n4420));
  not_8  g04044(.A(new_n4420), .Y(new_n4421));
  or_6   g04045(.A(new_n978), .B(new_n977), .Y(new_n4422));
  nand_5 g04046(.A(new_n984), .B(new_n979), .Y(new_n4423));
  nand_5 g04047(.A(new_n4423), .B(new_n4422), .Y(new_n4424));
  nand_5 g04048(.A(new_n4424), .B(new_n4421), .Y(new_n4425));
  xor_4  g04049(.A(new_n4424), .B(new_n4420), .Y(new_n4426));
  xor_4  g04050(.A(new_n4416), .B(new_n4415), .Y(new_n4427));
  or_6   g04051(.A(new_n4427), .B(new_n4426), .Y(new_n4428));
  nand_5 g04052(.A(new_n4428), .B(new_n4425), .Y(new_n4429));
  nand_5 g04053(.A(new_n4429), .B(new_n4419), .Y(new_n4430));
  nand_5 g04054(.A(pi200), .B(pi162), .Y(new_n4431));
  nand_5 g04055(.A(pi179), .B(pi167), .Y(new_n4432));
  xor_4  g04056(.A(new_n4432), .B(new_n4431), .Y(new_n4433));
  xor_4  g04057(.A(new_n4433), .B(new_n4399), .Y(new_n4434));
  nand_5 g04058(.A(pi149), .B(pi048), .Y(new_n4435));
  xor_4  g04059(.A(new_n4435), .B(new_n4400), .Y(new_n4436));
  xor_4  g04060(.A(new_n4436), .B(new_n4434), .Y(new_n4437));
  nand_5 g04061(.A(pi238), .B(pi134), .Y(new_n4438));
  nand_5 g04062(.A(pi193), .B(pi175), .Y(new_n4439));
  xor_4  g04063(.A(new_n4439), .B(new_n4438), .Y(new_n4440));
  xor_4  g04064(.A(new_n4440), .B(new_n4407), .Y(new_n4441));
  nor_5  g04065(.A(new_n4394), .B(new_n4387), .Y(new_n4442));
  nor_5  g04066(.A(new_n4401), .B(new_n4395), .Y(new_n4443));
  nor_5  g04067(.A(new_n4443), .B(new_n4442), .Y(new_n4444));
  xor_4  g04068(.A(new_n4444), .B(new_n4441), .Y(new_n4445));
  xnor_4 g04069(.A(new_n4445), .B(new_n4437), .Y(new_n4446));
  nor_5  g04070(.A(new_n4409), .B(new_n4402), .Y(new_n4447));
  nor_5  g04071(.A(new_n4418), .B(new_n4410), .Y(new_n4448));
  xor_4  g04072(.A(new_n4448), .B(new_n4408), .Y(new_n4449));
  nor_5  g04073(.A(new_n4449), .B(new_n4447), .Y(new_n4450));
  not_8  g04074(.A(new_n4450), .Y(new_n4451));
  xor_4  g04075(.A(new_n4451), .B(new_n4446), .Y(new_n4452));
  xor_4  g04076(.A(new_n4452), .B(new_n4430), .Y(new_n4453));
  nand_5 g04077(.A(pi238), .B(pi175), .Y(new_n4454));
  nor_5  g04078(.A(new_n992), .B(new_n985), .Y(new_n4455));
  xor_4  g04079(.A(new_n4427), .B(new_n4426), .Y(new_n4456));
  nand_5 g04080(.A(new_n4456), .B(new_n4455), .Y(new_n4457));
  nand_5 g04081(.A(new_n4457), .B(new_n4454), .Y(new_n4458));
  xor_4  g04082(.A(new_n4429), .B(new_n4419), .Y(new_n4459));
  not_8  g04083(.A(new_n4459), .Y(new_n4460));
  xor_4  g04084(.A(new_n4457), .B(new_n4454), .Y(new_n4461));
  nand_5 g04085(.A(new_n4461), .B(new_n4460), .Y(new_n4462));
  nand_5 g04086(.A(new_n4462), .B(new_n4458), .Y(new_n4463));
  xor_4  g04087(.A(new_n4463), .B(new_n4453), .Y(new_n4464));
  xor_4  g04088(.A(new_n4464), .B(new_n4386), .Y(new_n4465));
  xor_4  g04089(.A(new_n4461), .B(new_n4459), .Y(new_n4466));
  xnor_4 g04090(.A(new_n4456), .B(new_n4455), .Y(new_n4467));
  or_6   g04091(.A(new_n1011), .B(new_n993), .Y(new_n4468));
  not_8  g04092(.A(new_n970), .Y(new_n4469));
  nand_5 g04093(.A(new_n1012), .B(new_n4469), .Y(new_n4470));
  nand_5 g04094(.A(new_n4470), .B(new_n4468), .Y(new_n4471));
  or_6   g04095(.A(new_n4471), .B(new_n4467), .Y(new_n4472));
  xnor_4 g04096(.A(new_n4381), .B(new_n4380), .Y(new_n4473));
  xor_4  g04097(.A(new_n4471), .B(new_n4467), .Y(new_n4474));
  nand_5 g04098(.A(new_n4474), .B(new_n4473), .Y(new_n4475));
  nand_5 g04099(.A(new_n4475), .B(new_n4472), .Y(new_n4476));
  nand_5 g04100(.A(new_n4476), .B(new_n4466), .Y(new_n4477));
  xor_4  g04101(.A(new_n4383), .B(new_n4374), .Y(new_n4478));
  xor_4  g04102(.A(new_n4476), .B(new_n4466), .Y(new_n4479));
  nand_5 g04103(.A(new_n4479), .B(new_n4478), .Y(new_n4480));
  nand_5 g04104(.A(new_n4480), .B(new_n4477), .Y(new_n4481));
  xor_4  g04105(.A(new_n4481), .B(new_n4465), .Y(new_n4482));
  nand_5 g04106(.A(pi194), .B(pi080), .Y(new_n4483));
  nand_5 g04107(.A(pi247), .B(pi143), .Y(new_n4484));
  nand_5 g04108(.A(pi080), .B(pi057), .Y(new_n4485));
  nand_5 g04109(.A(new_n4485), .B(new_n4484), .Y(new_n4486));
  nand_5 g04110(.A(pi194), .B(pi016), .Y(new_n4487));
  xor_4  g04111(.A(new_n4485), .B(new_n4484), .Y(new_n4488));
  nand_5 g04112(.A(new_n4488), .B(new_n4487), .Y(new_n4489));
  nand_5 g04113(.A(new_n4489), .B(new_n4486), .Y(new_n4490));
  xnor_4 g04114(.A(new_n4490), .B(new_n4483), .Y(new_n4491));
  nand_5 g04115(.A(pi247), .B(pi057), .Y(new_n4492));
  nand_5 g04116(.A(pi234), .B(pi143), .Y(new_n4493));
  nand_5 g04117(.A(new_n4493), .B(new_n4492), .Y(new_n4494));
  nand_5 g04118(.A(pi234), .B(pi057), .Y(new_n4495));
  or_6   g04119(.A(new_n4495), .B(new_n4484), .Y(new_n4496));
  nand_5 g04120(.A(new_n4496), .B(new_n4494), .Y(new_n4497));
  xnor_4 g04121(.A(new_n4497), .B(new_n4491), .Y(new_n4498));
  nand_5 g04122(.A(pi085), .B(pi016), .Y(new_n4499));
  nand_5 g04123(.A(pi180), .B(pi117), .Y(new_n4500));
  and_6  g04124(.A(new_n4500), .B(new_n4499), .Y(new_n4501));
  nand_5 g04125(.A(pi117), .B(pi085), .Y(new_n4502));
  nand_5 g04126(.A(pi180), .B(pi016), .Y(new_n4503));
  nor_5  g04127(.A(new_n4503), .B(new_n4502), .Y(new_n4504));
  or_6   g04128(.A(new_n4504), .B(new_n4501), .Y(new_n4505));
  xnor_4 g04129(.A(new_n4505), .B(new_n4498), .Y(new_n4506));
  nand_5 g04130(.A(new_n1025), .B(new_n1024), .Y(new_n4507));
  nand_5 g04131(.A(new_n1026), .B(new_n1023), .Y(new_n4508));
  nand_5 g04132(.A(new_n4508), .B(new_n4507), .Y(new_n4509));
  nand_5 g04133(.A(new_n4509), .B(new_n4502), .Y(new_n4510));
  xor_4  g04134(.A(new_n4488), .B(new_n4487), .Y(new_n4511));
  xor_4  g04135(.A(new_n4509), .B(new_n4502), .Y(new_n4512));
  nand_5 g04136(.A(new_n4512), .B(new_n4511), .Y(new_n4513));
  nand_5 g04137(.A(new_n4513), .B(new_n4510), .Y(new_n4514));
  xor_4  g04138(.A(new_n4514), .B(new_n4506), .Y(new_n4515));
  nand_5 g04139(.A(pi180), .B(pi103), .Y(new_n4516));
  nand_5 g04140(.A(new_n1031), .B(new_n1028), .Y(new_n4517));
  nand_5 g04141(.A(new_n1032), .B(new_n1027), .Y(new_n4518));
  nand_5 g04142(.A(new_n4518), .B(new_n4517), .Y(new_n4519));
  or_6   g04143(.A(new_n4519), .B(new_n4516), .Y(new_n4520));
  xnor_4 g04144(.A(new_n4512), .B(new_n4511), .Y(new_n4521));
  xor_4  g04145(.A(new_n4519), .B(new_n4516), .Y(new_n4522));
  nand_5 g04146(.A(new_n4522), .B(new_n4521), .Y(new_n4523));
  nand_5 g04147(.A(new_n4523), .B(new_n4520), .Y(new_n4524));
  nand_5 g04148(.A(new_n4524), .B(new_n4515), .Y(new_n4525));
  nand_5 g04149(.A(pi214), .B(pi143), .Y(new_n4526));
  nand_5 g04150(.A(pi247), .B(pi194), .Y(new_n4527));
  xor_4  g04151(.A(new_n4527), .B(new_n4526), .Y(new_n4528));
  xor_4  g04152(.A(new_n4528), .B(new_n4495), .Y(new_n4529));
  nand_5 g04153(.A(pi085), .B(pi080), .Y(new_n4530));
  xor_4  g04154(.A(new_n4530), .B(new_n4496), .Y(new_n4531));
  xor_4  g04155(.A(new_n4531), .B(new_n4529), .Y(new_n4532));
  nand_5 g04156(.A(pi117), .B(pi036), .Y(new_n4533));
  nand_5 g04157(.A(pi103), .B(pi068), .Y(new_n4534));
  xor_4  g04158(.A(new_n4534), .B(new_n4533), .Y(new_n4535));
  xor_4  g04159(.A(new_n4535), .B(new_n4503), .Y(new_n4536));
  nor_5  g04160(.A(new_n4490), .B(new_n4483), .Y(new_n4537));
  nor_5  g04161(.A(new_n4497), .B(new_n4491), .Y(new_n4538));
  nor_5  g04162(.A(new_n4538), .B(new_n4537), .Y(new_n4539));
  xor_4  g04163(.A(new_n4539), .B(new_n4536), .Y(new_n4540));
  xnor_4 g04164(.A(new_n4540), .B(new_n4532), .Y(new_n4541));
  nor_5  g04165(.A(new_n4505), .B(new_n4498), .Y(new_n4542));
  nor_5  g04166(.A(new_n4514), .B(new_n4506), .Y(new_n4543));
  xor_4  g04167(.A(new_n4543), .B(new_n4504), .Y(new_n4544));
  nor_5  g04168(.A(new_n4544), .B(new_n4542), .Y(new_n4545));
  xor_4  g04169(.A(new_n4545), .B(new_n4541), .Y(new_n4546));
  xor_4  g04170(.A(new_n4546), .B(new_n4525), .Y(new_n4547));
  nand_5 g04171(.A(pi103), .B(pi036), .Y(new_n4548));
  nor_5  g04172(.A(new_n1033), .B(new_n1022), .Y(new_n4549));
  xor_4  g04173(.A(new_n4522), .B(new_n4521), .Y(new_n4550));
  nand_5 g04174(.A(new_n4550), .B(new_n4549), .Y(new_n4551));
  nand_5 g04175(.A(new_n4551), .B(new_n4548), .Y(new_n4552));
  xnor_4 g04176(.A(new_n4524), .B(new_n4515), .Y(new_n4553));
  xor_4  g04177(.A(new_n4551), .B(new_n4548), .Y(new_n4554));
  nand_5 g04178(.A(new_n4554), .B(new_n4553), .Y(new_n4555));
  nand_5 g04179(.A(new_n4555), .B(new_n4552), .Y(new_n4556));
  xor_4  g04180(.A(new_n4556), .B(new_n4547), .Y(new_n4557));
  xor_4  g04181(.A(new_n4554), .B(new_n4553), .Y(new_n4558));
  xor_4  g04182(.A(new_n4550), .B(new_n4549), .Y(new_n4559));
  nand_5 g04183(.A(new_n1052), .B(new_n1034), .Y(new_n4560));
  nand_5 g04184(.A(new_n1053), .B(new_n1013), .Y(new_n4561));
  nand_5 g04185(.A(new_n4561), .B(new_n4560), .Y(new_n4562));
  or_6   g04186(.A(new_n4562), .B(new_n4559), .Y(new_n4563));
  xor_4  g04187(.A(new_n4474), .B(new_n4473), .Y(new_n4564));
  not_8  g04188(.A(new_n4564), .Y(new_n4565));
  xor_4  g04189(.A(new_n4562), .B(new_n4559), .Y(new_n4566));
  nand_5 g04190(.A(new_n4566), .B(new_n4565), .Y(new_n4567));
  nand_5 g04191(.A(new_n4567), .B(new_n4563), .Y(new_n4568));
  nand_5 g04192(.A(new_n4568), .B(new_n4558), .Y(new_n4569));
  xor_4  g04193(.A(new_n4479), .B(new_n4478), .Y(new_n4570));
  not_8  g04194(.A(new_n4570), .Y(new_n4571));
  xor_4  g04195(.A(new_n4568), .B(new_n4558), .Y(new_n4572));
  nand_5 g04196(.A(new_n4572), .B(new_n4571), .Y(new_n4573));
  nand_5 g04197(.A(new_n4573), .B(new_n4569), .Y(new_n4574));
  xor_4  g04198(.A(new_n4574), .B(new_n4557), .Y(new_n4575));
  xor_4  g04199(.A(new_n4575), .B(new_n4482), .Y(po014));
  nand_5 g04200(.A(pi241), .B(pi042), .Y(new_n4577));
  nand_5 g04201(.A(pi236), .B(pi108), .Y(new_n4578));
  xor_4  g04202(.A(new_n4578), .B(new_n4577), .Y(new_n4579));
  nand_5 g04203(.A(pi161), .B(pi051), .Y(new_n4580));
  xor_4  g04204(.A(new_n4580), .B(new_n4579), .Y(new_n4581));
  nor_5  g04205(.A(new_n4577), .B(new_n3513), .Y(new_n4582));
  not_8  g04206(.A(new_n4582), .Y(new_n4583));
  or_6   g04207(.A(new_n4583), .B(new_n4581), .Y(new_n4584));
  nand_5 g04208(.A(pi236), .B(pi007), .Y(new_n4585));
  nand_5 g04209(.A(new_n4578), .B(new_n4577), .Y(new_n4586));
  nand_5 g04210(.A(new_n4580), .B(new_n4579), .Y(new_n4587));
  nand_5 g04211(.A(new_n4587), .B(new_n4586), .Y(new_n4588));
  xor_4  g04212(.A(new_n4588), .B(new_n4585), .Y(new_n4589));
  nand_5 g04213(.A(pi141), .B(pi051), .Y(new_n4590));
  nand_5 g04214(.A(pi241), .B(pi108), .Y(new_n4591));
  nand_5 g04215(.A(pi161), .B(pi042), .Y(new_n4592));
  xor_4  g04216(.A(new_n4592), .B(new_n4591), .Y(new_n4593));
  xor_4  g04217(.A(new_n4593), .B(new_n4590), .Y(new_n4594));
  xor_4  g04218(.A(new_n4594), .B(new_n4589), .Y(new_n4595));
  nor_5  g04219(.A(new_n4595), .B(new_n4584), .Y(new_n4596));
  nand_5 g04220(.A(pi161), .B(pi108), .Y(new_n4597));
  nand_5 g04221(.A(pi090), .B(pi051), .Y(new_n4598));
  nand_5 g04222(.A(pi141), .B(pi042), .Y(new_n4599));
  xor_4  g04223(.A(new_n4599), .B(new_n4598), .Y(new_n4600));
  xor_4  g04224(.A(new_n4600), .B(new_n4597), .Y(new_n4601));
  nand_5 g04225(.A(pi241), .B(pi007), .Y(new_n4602));
  nand_5 g04226(.A(new_n4592), .B(new_n4591), .Y(new_n4603));
  nand_5 g04227(.A(new_n4593), .B(new_n4590), .Y(new_n4604));
  nand_5 g04228(.A(new_n4604), .B(new_n4603), .Y(new_n4605));
  xor_4  g04229(.A(new_n4605), .B(new_n4602), .Y(new_n4606));
  xor_4  g04230(.A(new_n4606), .B(new_n4601), .Y(new_n4607));
  nand_5 g04231(.A(pi236), .B(pi118), .Y(new_n4608));
  or_6   g04232(.A(new_n4588), .B(new_n4585), .Y(new_n4609));
  not_8  g04233(.A(new_n4594), .Y(new_n4610));
  nand_5 g04234(.A(new_n4610), .B(new_n4589), .Y(new_n4611));
  nand_5 g04235(.A(new_n4611), .B(new_n4609), .Y(new_n4612));
  xor_4  g04236(.A(new_n4612), .B(new_n4608), .Y(new_n4613));
  xor_4  g04237(.A(new_n4613), .B(new_n4607), .Y(new_n4614));
  xor_4  g04238(.A(new_n4614), .B(new_n4596), .Y(new_n4615));
  nand_5 g04239(.A(pi212), .B(pi178), .Y(new_n4616));
  nand_5 g04240(.A(pi213), .B(pi061), .Y(new_n4617));
  xor_4  g04241(.A(new_n4617), .B(new_n4616), .Y(new_n4618));
  nand_5 g04242(.A(pi188), .B(pi104), .Y(new_n4619));
  xor_4  g04243(.A(new_n4619), .B(new_n4618), .Y(new_n4620));
  nor_5  g04244(.A(new_n4616), .B(new_n3514), .Y(new_n4621));
  not_8  g04245(.A(new_n4621), .Y(new_n4622));
  or_6   g04246(.A(new_n4622), .B(new_n4620), .Y(new_n4623));
  nand_5 g04247(.A(pi188), .B(pi013), .Y(new_n4624));
  nand_5 g04248(.A(pi212), .B(pi061), .Y(new_n4625));
  nand_5 g04249(.A(pi178), .B(pi104), .Y(new_n4626));
  xor_4  g04250(.A(new_n4626), .B(new_n4625), .Y(new_n4627));
  xor_4  g04251(.A(new_n4627), .B(new_n4624), .Y(new_n4628));
  nand_5 g04252(.A(pi213), .B(pi012), .Y(new_n4629));
  nand_5 g04253(.A(new_n4617), .B(new_n4616), .Y(new_n4630));
  nand_5 g04254(.A(new_n4619), .B(new_n4618), .Y(new_n4631));
  nand_5 g04255(.A(new_n4631), .B(new_n4630), .Y(new_n4632));
  xor_4  g04256(.A(new_n4632), .B(new_n4629), .Y(new_n4633));
  xor_4  g04257(.A(new_n4633), .B(new_n4628), .Y(new_n4634));
  or_6   g04258(.A(new_n4634), .B(new_n4623), .Y(new_n4635));
  nand_5 g04259(.A(pi188), .B(pi112), .Y(new_n4636));
  nand_5 g04260(.A(pi104), .B(pi061), .Y(new_n4637));
  nand_5 g04261(.A(pi178), .B(pi013), .Y(new_n4638));
  xor_4  g04262(.A(new_n4638), .B(new_n4637), .Y(new_n4639));
  xor_4  g04263(.A(new_n4639), .B(new_n4636), .Y(new_n4640));
  nand_5 g04264(.A(pi212), .B(pi012), .Y(new_n4641));
  nand_5 g04265(.A(new_n4626), .B(new_n4625), .Y(new_n4642));
  nand_5 g04266(.A(new_n4627), .B(new_n4624), .Y(new_n4643));
  nand_5 g04267(.A(new_n4643), .B(new_n4642), .Y(new_n4644));
  xor_4  g04268(.A(new_n4644), .B(new_n4641), .Y(new_n4645));
  xnor_4 g04269(.A(new_n4645), .B(new_n4640), .Y(new_n4646));
  nand_5 g04270(.A(pi213), .B(pi144), .Y(new_n4647));
  nand_5 g04271(.A(new_n4632), .B(new_n4629), .Y(new_n4648));
  nand_5 g04272(.A(new_n4633), .B(new_n4628), .Y(new_n4649));
  nand_5 g04273(.A(new_n4649), .B(new_n4648), .Y(new_n4650));
  xor_4  g04274(.A(new_n4650), .B(new_n4647), .Y(new_n4651));
  xnor_4 g04275(.A(new_n4651), .B(new_n4646), .Y(new_n4652));
  xor_4  g04276(.A(new_n4652), .B(new_n4635), .Y(new_n4653));
  xor_4  g04277(.A(new_n4653), .B(new_n4615), .Y(new_n4654));
  xor_4  g04278(.A(new_n4595), .B(new_n4584), .Y(new_n4655));
  xor_4  g04279(.A(new_n4634), .B(new_n4623), .Y(new_n4656));
  nand_5 g04280(.A(new_n4656), .B(new_n4655), .Y(new_n4657));
  not_8  g04281(.A(new_n4657), .Y(new_n4658));
  xnor_4 g04282(.A(new_n4656), .B(new_n4655), .Y(new_n4659));
  xor_4  g04283(.A(new_n4621), .B(new_n4620), .Y(new_n4660));
  nor_5  g04284(.A(new_n3514), .B(new_n3513), .Y(new_n4661));
  not_8  g04285(.A(new_n4661), .Y(new_n4662));
  nand_5 g04286(.A(pi236), .B(pi042), .Y(new_n4663));
  nand_5 g04287(.A(pi241), .B(pi051), .Y(new_n4664));
  nand_5 g04288(.A(new_n4664), .B(new_n4663), .Y(new_n4665));
  nand_5 g04289(.A(new_n4665), .B(new_n4583), .Y(new_n4666));
  nor_5  g04290(.A(new_n4666), .B(new_n4662), .Y(new_n4667));
  xor_4  g04291(.A(new_n4666), .B(new_n4661), .Y(new_n4668));
  nand_5 g04292(.A(pi213), .B(pi178), .Y(new_n4669));
  nand_5 g04293(.A(pi212), .B(pi188), .Y(new_n4670));
  nand_5 g04294(.A(new_n4670), .B(new_n4669), .Y(new_n4671));
  nand_5 g04295(.A(new_n4671), .B(new_n4622), .Y(new_n4672));
  nor_5  g04296(.A(new_n4672), .B(new_n4668), .Y(new_n4673));
  nor_5  g04297(.A(new_n4673), .B(new_n4667), .Y(new_n4674));
  nand_5 g04298(.A(new_n4674), .B(new_n4660), .Y(new_n4675));
  xor_4  g04299(.A(new_n4582), .B(new_n4581), .Y(new_n4676));
  xor_4  g04300(.A(new_n4674), .B(new_n4660), .Y(new_n4677));
  nand_5 g04301(.A(new_n4677), .B(new_n4676), .Y(new_n4678));
  nand_5 g04302(.A(new_n4678), .B(new_n4675), .Y(new_n4679));
  nor_5  g04303(.A(new_n4679), .B(new_n4659), .Y(new_n4680));
  nor_5  g04304(.A(new_n4680), .B(new_n4658), .Y(new_n4681));
  xor_4  g04305(.A(new_n4681), .B(new_n4654), .Y(new_n4682));
  nand_5 g04306(.A(pi208), .B(pi033), .Y(new_n4683));
  nand_5 g04307(.A(pi179), .B(pi168), .Y(new_n4684));
  xor_4  g04308(.A(new_n4684), .B(new_n4683), .Y(new_n4685));
  nand_5 g04309(.A(pi162), .B(pi139), .Y(new_n4686));
  xor_4  g04310(.A(new_n4686), .B(new_n4685), .Y(new_n4687));
  nor_5  g04311(.A(new_n4683), .B(new_n3516), .Y(new_n4688));
  not_8  g04312(.A(new_n4688), .Y(new_n4689));
  or_6   g04313(.A(new_n4689), .B(new_n4687), .Y(new_n4690));
  nand_5 g04314(.A(pi168), .B(pi048), .Y(new_n4691));
  nand_5 g04315(.A(new_n4684), .B(new_n4683), .Y(new_n4692));
  nand_5 g04316(.A(new_n4686), .B(new_n4685), .Y(new_n4693));
  nand_5 g04317(.A(new_n4693), .B(new_n4692), .Y(new_n4694));
  xor_4  g04318(.A(new_n4694), .B(new_n4691), .Y(new_n4695));
  nand_5 g04319(.A(pi208), .B(pi179), .Y(new_n4696));
  nand_5 g04320(.A(pi162), .B(pi035), .Y(new_n4697));
  nand_5 g04321(.A(pi139), .B(pi033), .Y(new_n4698));
  xor_4  g04322(.A(new_n4698), .B(new_n4697), .Y(new_n4699));
  xnor_4 g04323(.A(new_n4699), .B(new_n4696), .Y(new_n4700));
  xnor_4 g04324(.A(new_n4700), .B(new_n4695), .Y(new_n4701));
  nor_5  g04325(.A(new_n4701), .B(new_n4690), .Y(new_n4702));
  nand_5 g04326(.A(pi179), .B(pi139), .Y(new_n4703));
  nand_5 g04327(.A(pi035), .B(pi033), .Y(new_n4704));
  nand_5 g04328(.A(pi162), .B(pi015), .Y(new_n4705));
  xor_4  g04329(.A(new_n4705), .B(new_n4704), .Y(new_n4706));
  xor_4  g04330(.A(new_n4706), .B(new_n4703), .Y(new_n4707));
  nand_5 g04331(.A(pi208), .B(pi048), .Y(new_n4708));
  nand_5 g04332(.A(new_n4698), .B(new_n4697), .Y(new_n4709));
  nand_5 g04333(.A(new_n4699), .B(new_n4696), .Y(new_n4710));
  nand_5 g04334(.A(new_n4710), .B(new_n4709), .Y(new_n4711));
  xor_4  g04335(.A(new_n4711), .B(new_n4708), .Y(new_n4712));
  xor_4  g04336(.A(new_n4712), .B(new_n4707), .Y(new_n4713));
  nand_5 g04337(.A(pi237), .B(pi168), .Y(new_n4714));
  or_6   g04338(.A(new_n4694), .B(new_n4691), .Y(new_n4715));
  nand_5 g04339(.A(new_n4700), .B(new_n4695), .Y(new_n4716));
  nand_5 g04340(.A(new_n4716), .B(new_n4715), .Y(new_n4717));
  xor_4  g04341(.A(new_n4717), .B(new_n4714), .Y(new_n4718));
  xor_4  g04342(.A(new_n4718), .B(new_n4713), .Y(new_n4719));
  xor_4  g04343(.A(new_n4719), .B(new_n4702), .Y(new_n4720));
  xor_4  g04344(.A(new_n4679), .B(new_n4659), .Y(new_n4721));
  xor_4  g04345(.A(new_n4701), .B(new_n4690), .Y(new_n4722));
  nor_5  g04346(.A(new_n4722), .B(new_n4721), .Y(new_n4723));
  xnor_4 g04347(.A(new_n4722), .B(new_n4721), .Y(new_n4724));
  xor_4  g04348(.A(new_n4688), .B(new_n4687), .Y(new_n4725));
  not_8  g04349(.A(new_n3515), .Y(new_n4726));
  or_6   g04350(.A(new_n3516), .B(new_n4726), .Y(new_n4727));
  nand_5 g04351(.A(pi168), .B(pi033), .Y(new_n4728));
  nand_5 g04352(.A(pi208), .B(pi162), .Y(new_n4729));
  nand_5 g04353(.A(new_n4729), .B(new_n4728), .Y(new_n4730));
  nand_5 g04354(.A(new_n4730), .B(new_n4689), .Y(new_n4731));
  nand_5 g04355(.A(new_n4731), .B(new_n4727), .Y(new_n4732));
  xor_4  g04356(.A(new_n4672), .B(new_n4668), .Y(new_n4733));
  not_8  g04357(.A(new_n4733), .Y(new_n4734));
  xor_4  g04358(.A(new_n4731), .B(new_n4727), .Y(new_n4735));
  nand_5 g04359(.A(new_n4735), .B(new_n4734), .Y(new_n4736));
  nand_5 g04360(.A(new_n4736), .B(new_n4732), .Y(new_n4737));
  or_6   g04361(.A(new_n4737), .B(new_n4725), .Y(new_n4738));
  xor_4  g04362(.A(new_n4677), .B(new_n4676), .Y(new_n4739));
  not_8  g04363(.A(new_n4739), .Y(new_n4740));
  xor_4  g04364(.A(new_n4737), .B(new_n4725), .Y(new_n4741));
  nand_5 g04365(.A(new_n4741), .B(new_n4740), .Y(new_n4742));
  nand_5 g04366(.A(new_n4742), .B(new_n4738), .Y(new_n4743));
  nor_5  g04367(.A(new_n4743), .B(new_n4724), .Y(new_n4744));
  nor_5  g04368(.A(new_n4744), .B(new_n4723), .Y(new_n4745));
  xor_4  g04369(.A(new_n4745), .B(new_n4720), .Y(new_n4746));
  xor_4  g04370(.A(new_n4746), .B(new_n4682), .Y(new_n4747));
  nand_5 g04371(.A(pi057), .B(pi052), .Y(new_n4748));
  nand_5 g04372(.A(pi194), .B(pi131), .Y(new_n4749));
  xor_4  g04373(.A(new_n4749), .B(new_n4748), .Y(new_n4750));
  nand_5 g04374(.A(pi143), .B(pi077), .Y(new_n4751));
  xor_4  g04375(.A(new_n4751), .B(new_n4750), .Y(new_n4752));
  nand_5 g04376(.A(pi131), .B(pi057), .Y(new_n4753));
  nand_5 g04377(.A(pi143), .B(pi052), .Y(new_n4754));
  nor_5  g04378(.A(new_n4754), .B(new_n4753), .Y(new_n4755));
  not_8  g04379(.A(new_n4755), .Y(new_n4756));
  nor_5  g04380(.A(new_n4756), .B(new_n4752), .Y(new_n4757));
  not_8  g04381(.A(new_n4757), .Y(new_n4758));
  nand_5 g04382(.A(pi131), .B(pi085), .Y(new_n4759));
  nand_5 g04383(.A(new_n4749), .B(new_n4748), .Y(new_n4760));
  nand_5 g04384(.A(new_n4751), .B(new_n4750), .Y(new_n4761));
  nand_5 g04385(.A(new_n4761), .B(new_n4760), .Y(new_n4762));
  xor_4  g04386(.A(new_n4762), .B(new_n4759), .Y(new_n4763));
  nand_5 g04387(.A(pi077), .B(pi057), .Y(new_n4764));
  nand_5 g04388(.A(pi194), .B(pi052), .Y(new_n4765));
  nand_5 g04389(.A(pi143), .B(pi133), .Y(new_n4766));
  xor_4  g04390(.A(new_n4766), .B(new_n4765), .Y(new_n4767));
  xnor_4 g04391(.A(new_n4767), .B(new_n4764), .Y(new_n4768));
  xnor_4 g04392(.A(new_n4768), .B(new_n4763), .Y(new_n4769));
  nor_5  g04393(.A(new_n4769), .B(new_n4758), .Y(new_n4770));
  nand_5 g04394(.A(pi133), .B(pi057), .Y(new_n4771));
  nand_5 g04395(.A(pi189), .B(pi143), .Y(new_n4772));
  nand_5 g04396(.A(pi194), .B(pi077), .Y(new_n4773));
  xor_4  g04397(.A(new_n4773), .B(new_n4772), .Y(new_n4774));
  xor_4  g04398(.A(new_n4774), .B(new_n4771), .Y(new_n4775));
  nand_5 g04399(.A(pi085), .B(pi052), .Y(new_n4776));
  nand_5 g04400(.A(new_n4766), .B(new_n4765), .Y(new_n4777));
  nand_5 g04401(.A(new_n4767), .B(new_n4764), .Y(new_n4778));
  nand_5 g04402(.A(new_n4778), .B(new_n4777), .Y(new_n4779));
  xor_4  g04403(.A(new_n4779), .B(new_n4776), .Y(new_n4780));
  xor_4  g04404(.A(new_n4780), .B(new_n4775), .Y(new_n4781));
  nand_5 g04405(.A(pi180), .B(pi131), .Y(new_n4782));
  xor_4  g04406(.A(new_n4782), .B(new_n4781), .Y(new_n4783));
  or_6   g04407(.A(new_n4762), .B(new_n4759), .Y(new_n4784));
  nand_5 g04408(.A(new_n4768), .B(new_n4763), .Y(new_n4785));
  nand_5 g04409(.A(new_n4785), .B(new_n4784), .Y(new_n4786));
  xor_4  g04410(.A(new_n4786), .B(new_n4783), .Y(new_n4787));
  xor_4  g04411(.A(new_n4787), .B(new_n4770), .Y(new_n4788));
  xor_4  g04412(.A(new_n4788), .B(new_n4747), .Y(new_n4789));
  xor_4  g04413(.A(new_n4743), .B(new_n4724), .Y(new_n4790));
  xor_4  g04414(.A(new_n4769), .B(new_n4758), .Y(new_n4791));
  not_8  g04415(.A(new_n4791), .Y(new_n4792));
  nand_5 g04416(.A(new_n4792), .B(new_n4790), .Y(new_n4793));
  xor_4  g04417(.A(new_n4792), .B(new_n4790), .Y(new_n4794));
  xor_4  g04418(.A(new_n4741), .B(new_n4739), .Y(new_n4795));
  xor_4  g04419(.A(new_n4756), .B(new_n4752), .Y(new_n4796));
  not_8  g04420(.A(new_n4796), .Y(new_n4797));
  nor_5  g04421(.A(new_n4797), .B(new_n4795), .Y(new_n4798));
  xor_4  g04422(.A(new_n4796), .B(new_n4795), .Y(new_n4799));
  nor_5  g04423(.A(new_n3518), .B(new_n3517), .Y(new_n4800));
  xor_4  g04424(.A(new_n4754), .B(new_n4753), .Y(new_n4801));
  or_6   g04425(.A(new_n4801), .B(new_n4800), .Y(new_n4802));
  xor_4  g04426(.A(new_n4735), .B(new_n4734), .Y(new_n4803));
  xor_4  g04427(.A(new_n4801), .B(new_n4800), .Y(new_n4804));
  nand_5 g04428(.A(new_n4804), .B(new_n4803), .Y(new_n4805));
  nand_5 g04429(.A(new_n4805), .B(new_n4802), .Y(new_n4806));
  nor_5  g04430(.A(new_n4806), .B(new_n4799), .Y(new_n4807));
  nor_5  g04431(.A(new_n4807), .B(new_n4798), .Y(new_n4808));
  nand_5 g04432(.A(new_n4808), .B(new_n4794), .Y(new_n4809));
  nand_5 g04433(.A(new_n4809), .B(new_n4793), .Y(new_n4810));
  xor_4  g04434(.A(new_n4810), .B(new_n4789), .Y(po015));
  nand_5 g04435(.A(pi087), .B(pi007), .Y(new_n4812));
  nand_5 g04436(.A(pi108), .B(pi087), .Y(new_n4813));
  nand_5 g04437(.A(pi102), .B(pi051), .Y(new_n4814));
  nand_5 g04438(.A(new_n4814), .B(new_n4813), .Y(new_n4815));
  nand_5 g04439(.A(pi219), .B(pi042), .Y(new_n4816));
  or_6   g04440(.A(new_n4814), .B(new_n4813), .Y(new_n4817));
  nand_5 g04441(.A(new_n4817), .B(new_n4816), .Y(new_n4818));
  nand_5 g04442(.A(new_n4818), .B(new_n4815), .Y(new_n4819));
  xor_4  g04443(.A(new_n4819), .B(new_n4812), .Y(new_n4820));
  nand_5 g04444(.A(pi051), .B(pi001), .Y(new_n4821));
  nand_5 g04445(.A(pi219), .B(pi108), .Y(new_n4822));
  nand_5 g04446(.A(pi102), .B(pi042), .Y(new_n4823));
  xor_4  g04447(.A(new_n4823), .B(new_n4822), .Y(new_n4824));
  xnor_4 g04448(.A(new_n4824), .B(new_n4821), .Y(new_n4825));
  xnor_4 g04449(.A(new_n4825), .B(new_n4820), .Y(new_n4826));
  not_8  g04450(.A(new_n4816), .Y(new_n4827));
  not_8  g04451(.A(new_n4815), .Y(new_n4828));
  nand_5 g04452(.A(pi087), .B(pi051), .Y(new_n4829));
  nand_5 g04453(.A(new_n4829), .B(new_n4827), .Y(new_n4830));
  nand_5 g04454(.A(new_n4830), .B(new_n4828), .Y(new_n4831));
  nand_5 g04455(.A(new_n4831), .B(new_n4817), .Y(new_n4832));
  nand_5 g04456(.A(new_n4832), .B(new_n4827), .Y(new_n4833));
  xor_4  g04457(.A(new_n4833), .B(new_n4826), .Y(new_n4834));
  nand_5 g04458(.A(pi188), .B(pi169), .Y(new_n4835));
  nand_5 g04459(.A(pi142), .B(pi061), .Y(new_n4836));
  nand_5 g04460(.A(new_n4836), .B(new_n4835), .Y(new_n4837));
  nand_5 g04461(.A(pi178), .B(pi071), .Y(new_n4838));
  or_6   g04462(.A(new_n4836), .B(new_n4835), .Y(new_n4839));
  nand_5 g04463(.A(new_n4839), .B(new_n4838), .Y(new_n4840));
  nand_5 g04464(.A(new_n4840), .B(new_n4837), .Y(new_n4841));
  nand_5 g04465(.A(pi142), .B(pi012), .Y(new_n4842));
  xor_4  g04466(.A(new_n4842), .B(new_n4841), .Y(new_n4843));
  nand_5 g04467(.A(pi188), .B(pi123), .Y(new_n4844));
  nand_5 g04468(.A(pi071), .B(pi061), .Y(new_n4845));
  nand_5 g04469(.A(pi178), .B(pi169), .Y(new_n4846));
  xor_4  g04470(.A(new_n4846), .B(new_n4845), .Y(new_n4847));
  xor_4  g04471(.A(new_n4847), .B(new_n4844), .Y(new_n4848));
  xor_4  g04472(.A(new_n4848), .B(new_n4843), .Y(new_n4849));
  not_8  g04473(.A(new_n4838), .Y(new_n4850));
  not_8  g04474(.A(new_n4837), .Y(new_n4851));
  nand_5 g04475(.A(pi188), .B(pi142), .Y(new_n4852));
  nand_5 g04476(.A(new_n4852), .B(new_n4850), .Y(new_n4853));
  nand_5 g04477(.A(new_n4853), .B(new_n4851), .Y(new_n4854));
  nand_5 g04478(.A(new_n4854), .B(new_n4839), .Y(new_n4855));
  nand_5 g04479(.A(new_n4855), .B(new_n4850), .Y(new_n4856));
  xor_4  g04480(.A(new_n4856), .B(new_n4849), .Y(new_n4857));
  xor_4  g04481(.A(new_n4857), .B(new_n4834), .Y(new_n4858));
  nand_5 g04482(.A(pi087), .B(pi042), .Y(new_n4859));
  nand_5 g04483(.A(pi219), .B(pi051), .Y(new_n4860));
  xor_4  g04484(.A(new_n4860), .B(new_n4859), .Y(new_n4861));
  nand_5 g04485(.A(pi178), .B(pi142), .Y(new_n4862));
  nand_5 g04486(.A(pi188), .B(pi071), .Y(new_n4863));
  xor_4  g04487(.A(new_n4863), .B(new_n4862), .Y(new_n4864));
  or_6   g04488(.A(new_n4864), .B(new_n4861), .Y(new_n4865));
  nor_5  g04489(.A(new_n4852), .B(new_n4829), .Y(new_n4866));
  not_8  g04490(.A(new_n4866), .Y(new_n4867));
  xor_4  g04491(.A(new_n4864), .B(new_n4861), .Y(new_n4868));
  nand_5 g04492(.A(new_n4868), .B(new_n4867), .Y(new_n4869));
  nand_5 g04493(.A(new_n4869), .B(new_n4865), .Y(new_n4870));
  nor_5  g04494(.A(new_n4853), .B(new_n4851), .Y(new_n4871));
  or_6   g04495(.A(new_n4871), .B(new_n4855), .Y(new_n4872));
  or_6   g04496(.A(new_n4872), .B(new_n4870), .Y(new_n4873));
  xor_4  g04497(.A(new_n4872), .B(new_n4870), .Y(new_n4874));
  nor_5  g04498(.A(new_n4830), .B(new_n4828), .Y(new_n4875));
  nor_5  g04499(.A(new_n4875), .B(new_n4832), .Y(new_n4876));
  nand_5 g04500(.A(new_n4876), .B(new_n4874), .Y(new_n4877));
  nand_5 g04501(.A(new_n4877), .B(new_n4873), .Y(new_n4878));
  xor_4  g04502(.A(new_n4878), .B(new_n4858), .Y(new_n4879));
  nand_5 g04503(.A(pi182), .B(pi033), .Y(new_n4880));
  nand_5 g04504(.A(pi179), .B(pi138), .Y(new_n4881));
  xor_4  g04505(.A(new_n4881), .B(new_n4880), .Y(new_n4882));
  nand_5 g04506(.A(pi162), .B(pi041), .Y(new_n4883));
  xor_4  g04507(.A(new_n4883), .B(new_n4882), .Y(new_n4884));
  nand_5 g04508(.A(pi138), .B(pi033), .Y(new_n4885));
  nand_5 g04509(.A(pi182), .B(pi162), .Y(new_n4886));
  nor_5  g04510(.A(new_n4886), .B(new_n4885), .Y(new_n4887));
  not_8  g04511(.A(new_n4887), .Y(new_n4888));
  nor_5  g04512(.A(new_n4888), .B(new_n4884), .Y(new_n4889));
  nand_5 g04513(.A(pi182), .B(pi179), .Y(new_n4890));
  nand_5 g04514(.A(pi041), .B(pi033), .Y(new_n4891));
  nand_5 g04515(.A(pi216), .B(pi162), .Y(new_n4892));
  xor_4  g04516(.A(new_n4892), .B(new_n4891), .Y(new_n4893));
  xor_4  g04517(.A(new_n4893), .B(new_n4890), .Y(new_n4894));
  nand_5 g04518(.A(pi138), .B(pi048), .Y(new_n4895));
  nand_5 g04519(.A(new_n4881), .B(new_n4880), .Y(new_n4896));
  nand_5 g04520(.A(new_n4883), .B(new_n4882), .Y(new_n4897));
  nand_5 g04521(.A(new_n4897), .B(new_n4896), .Y(new_n4898));
  xor_4  g04522(.A(new_n4898), .B(new_n4895), .Y(new_n4899));
  xor_4  g04523(.A(new_n4899), .B(new_n4894), .Y(new_n4900));
  xor_4  g04524(.A(new_n4900), .B(new_n4889), .Y(new_n4901));
  xnor_4 g04525(.A(new_n4876), .B(new_n4874), .Y(new_n4902));
  xor_4  g04526(.A(new_n4887), .B(new_n4884), .Y(new_n4903));
  nor_5  g04527(.A(new_n4903), .B(new_n4902), .Y(new_n4904));
  xnor_4 g04528(.A(new_n4903), .B(new_n4902), .Y(new_n4905));
  nand_5 g04529(.A(pi162), .B(pi138), .Y(new_n4906));
  xor_4  g04530(.A(new_n4852), .B(new_n4829), .Y(new_n4907));
  not_8  g04531(.A(new_n4907), .Y(new_n4908));
  nor_5  g04532(.A(new_n4908), .B(new_n4906), .Y(new_n4909));
  xor_4  g04533(.A(new_n4886), .B(new_n4885), .Y(new_n4910));
  or_6   g04534(.A(new_n4910), .B(new_n4909), .Y(new_n4911));
  xor_4  g04535(.A(new_n4868), .B(new_n4867), .Y(new_n4912));
  xor_4  g04536(.A(new_n4910), .B(new_n4909), .Y(new_n4913));
  nand_5 g04537(.A(new_n4913), .B(new_n4912), .Y(new_n4914));
  nand_5 g04538(.A(new_n4914), .B(new_n4911), .Y(new_n4915));
  nor_5  g04539(.A(new_n4915), .B(new_n4905), .Y(new_n4916));
  nor_5  g04540(.A(new_n4916), .B(new_n4904), .Y(new_n4917));
  xor_4  g04541(.A(new_n4917), .B(new_n4901), .Y(new_n4918));
  xor_4  g04542(.A(new_n4918), .B(new_n4879), .Y(new_n4919));
  nand_5 g04543(.A(pi057), .B(pi020), .Y(new_n4920));
  nand_5 g04544(.A(pi194), .B(pi160), .Y(new_n4921));
  xor_4  g04545(.A(new_n4921), .B(new_n4920), .Y(new_n4922));
  nand_5 g04546(.A(pi143), .B(pi060), .Y(new_n4923));
  xor_4  g04547(.A(new_n4923), .B(new_n4922), .Y(new_n4924));
  nand_5 g04548(.A(pi160), .B(pi143), .Y(new_n4925));
  or_6   g04549(.A(new_n4925), .B(new_n4920), .Y(new_n4926));
  nor_5  g04550(.A(new_n4926), .B(new_n4924), .Y(new_n4927));
  nand_5 g04551(.A(pi194), .B(pi020), .Y(new_n4928));
  nand_5 g04552(.A(pi223), .B(pi143), .Y(new_n4929));
  nand_5 g04553(.A(pi060), .B(pi057), .Y(new_n4930));
  xor_4  g04554(.A(new_n4930), .B(new_n4929), .Y(new_n4931));
  xor_4  g04555(.A(new_n4931), .B(new_n4928), .Y(new_n4932));
  nand_5 g04556(.A(pi160), .B(pi085), .Y(new_n4933));
  nand_5 g04557(.A(new_n4921), .B(new_n4920), .Y(new_n4934));
  nand_5 g04558(.A(new_n4923), .B(new_n4922), .Y(new_n4935));
  nand_5 g04559(.A(new_n4935), .B(new_n4934), .Y(new_n4936));
  xor_4  g04560(.A(new_n4936), .B(new_n4933), .Y(new_n4937));
  xor_4  g04561(.A(new_n4937), .B(new_n4932), .Y(new_n4938));
  xor_4  g04562(.A(new_n4938), .B(new_n4927), .Y(new_n4939));
  xor_4  g04563(.A(new_n4926), .B(new_n4924), .Y(new_n4940));
  xor_4  g04564(.A(new_n4907), .B(new_n4906), .Y(new_n4941));
  or_6   g04565(.A(new_n4941), .B(new_n4925), .Y(new_n4942));
  nand_5 g04566(.A(pi160), .B(pi057), .Y(new_n4943));
  nand_5 g04567(.A(pi143), .B(pi020), .Y(new_n4944));
  nand_5 g04568(.A(new_n4944), .B(new_n4943), .Y(new_n4945));
  nand_5 g04569(.A(new_n4945), .B(new_n4926), .Y(new_n4946));
  or_6   g04570(.A(new_n4946), .B(new_n4942), .Y(new_n4947));
  xnor_4 g04571(.A(new_n4913), .B(new_n4912), .Y(new_n4948));
  xor_4  g04572(.A(new_n4946), .B(new_n4942), .Y(new_n4949));
  nand_5 g04573(.A(new_n4949), .B(new_n4948), .Y(new_n4950));
  nand_5 g04574(.A(new_n4950), .B(new_n4947), .Y(new_n4951));
  or_6   g04575(.A(new_n4951), .B(new_n4940), .Y(new_n4952));
  xor_4  g04576(.A(new_n4915), .B(new_n4905), .Y(new_n4953));
  not_8  g04577(.A(new_n4953), .Y(new_n4954));
  xor_4  g04578(.A(new_n4951), .B(new_n4940), .Y(new_n4955));
  nand_5 g04579(.A(new_n4955), .B(new_n4954), .Y(new_n4956));
  nand_5 g04580(.A(new_n4956), .B(new_n4952), .Y(new_n4957));
  xor_4  g04581(.A(new_n4957), .B(new_n4939), .Y(new_n4958));
  xor_4  g04582(.A(new_n4958), .B(new_n4919), .Y(po016));
  nand_5 g04583(.A(pi226), .B(pi163), .Y(new_n4960));
  nand_5 g04584(.A(pi109), .B(pi107), .Y(new_n4961));
  nor_5  g04585(.A(new_n4961), .B(new_n4960), .Y(new_n4962));
  nand_5 g04586(.A(pi226), .B(pi148), .Y(new_n4963));
  nand_5 g04587(.A(pi207), .B(pi163), .Y(new_n4964));
  nand_5 g04588(.A(new_n4964), .B(new_n4963), .Y(new_n4965));
  nand_5 g04589(.A(pi207), .B(pi148), .Y(new_n4966));
  nor_5  g04590(.A(new_n4966), .B(new_n4960), .Y(new_n4967));
  not_8  g04591(.A(new_n4967), .Y(new_n4968));
  nand_5 g04592(.A(new_n4968), .B(new_n4965), .Y(new_n4969));
  xor_4  g04593(.A(new_n4969), .B(new_n4962), .Y(new_n4970));
  nand_5 g04594(.A(pi107), .B(pi014), .Y(new_n4971));
  nand_5 g04595(.A(pi171), .B(pi109), .Y(new_n4972));
  nand_5 g04596(.A(new_n4972), .B(new_n4971), .Y(new_n4973));
  nand_5 g04597(.A(pi171), .B(pi014), .Y(new_n4974));
  nor_5  g04598(.A(new_n4974), .B(new_n4961), .Y(new_n4975));
  not_8  g04599(.A(new_n4975), .Y(new_n4976));
  nand_5 g04600(.A(new_n4976), .B(new_n4973), .Y(new_n4977));
  xor_4  g04601(.A(new_n4977), .B(new_n4970), .Y(new_n4978));
  xor_4  g04602(.A(new_n4961), .B(new_n4960), .Y(new_n4979));
  not_8  g04603(.A(new_n4979), .Y(new_n4980));
  nand_5 g04604(.A(pi175), .B(pi132), .Y(new_n4981));
  or_6   g04605(.A(new_n4981), .B(new_n4980), .Y(new_n4982));
  nand_5 g04606(.A(pi186), .B(pi175), .Y(new_n4983));
  nand_5 g04607(.A(pi134), .B(pi132), .Y(new_n4984));
  and_6  g04608(.A(new_n4984), .B(new_n4983), .Y(new_n4985));
  nand_5 g04609(.A(pi186), .B(pi134), .Y(new_n4986));
  nor_5  g04610(.A(new_n4986), .B(new_n4981), .Y(new_n4987));
  or_6   g04611(.A(new_n4987), .B(new_n4985), .Y(new_n4988));
  xor_4  g04612(.A(new_n4988), .B(new_n4982), .Y(new_n4989));
  xor_4  g04613(.A(new_n4989), .B(new_n4978), .Y(new_n4990));
  xor_4  g04614(.A(new_n4981), .B(new_n4979), .Y(new_n4991));
  nand_5 g04615(.A(pi103), .B(pi029), .Y(new_n4992));
  nor_5  g04616(.A(new_n4992), .B(new_n4991), .Y(new_n4993));
  nand_5 g04617(.A(pi117), .B(pi029), .Y(new_n4994));
  nand_5 g04618(.A(pi103), .B(pi069), .Y(new_n4995));
  xor_4  g04619(.A(new_n4995), .B(new_n4994), .Y(new_n4996));
  xor_4  g04620(.A(new_n4996), .B(new_n4993), .Y(new_n4997));
  xor_4  g04621(.A(new_n4997), .B(new_n4990), .Y(po017));
  xor_4  g04622(.A(new_n3113), .B(new_n3112), .Y(po018));
  nand_5 g04623(.A(pi173), .B(pi141), .Y(new_n5000));
  nand_5 g04624(.A(pi090), .B(pi014), .Y(new_n5001));
  nand_5 g04625(.A(pi109), .B(pi047), .Y(new_n5002));
  nand_5 g04626(.A(new_n5002), .B(new_n5001), .Y(new_n5003));
  nand_5 g04627(.A(pi109), .B(pi090), .Y(new_n5004));
  nand_5 g04628(.A(pi047), .B(pi014), .Y(new_n5005));
  or_6   g04629(.A(new_n5005), .B(new_n5004), .Y(new_n5006));
  nand_5 g04630(.A(new_n5006), .B(new_n5003), .Y(new_n5007));
  xor_4  g04631(.A(new_n5007), .B(new_n5000), .Y(new_n5008));
  nand_5 g04632(.A(pi141), .B(pi014), .Y(new_n5009));
  nand_5 g04633(.A(new_n5009), .B(new_n5004), .Y(new_n5010));
  nand_5 g04634(.A(pi173), .B(pi161), .Y(new_n5011));
  xor_4  g04635(.A(new_n5009), .B(new_n5004), .Y(new_n5012));
  nand_5 g04636(.A(new_n5012), .B(new_n5011), .Y(new_n5013));
  nand_5 g04637(.A(new_n5013), .B(new_n5010), .Y(new_n5014));
  xor_4  g04638(.A(new_n5014), .B(new_n5008), .Y(new_n5015));
  nand_5 g04639(.A(pi230), .B(pi161), .Y(new_n5016));
  nand_5 g04640(.A(pi241), .B(pi050), .Y(new_n5017));
  and_6  g04641(.A(new_n5017), .B(new_n5016), .Y(new_n5018));
  nand_5 g04642(.A(pi241), .B(pi230), .Y(new_n5019));
  nand_5 g04643(.A(pi161), .B(pi050), .Y(new_n5020));
  nor_5  g04644(.A(new_n5020), .B(new_n5019), .Y(new_n5021));
  or_6   g04645(.A(new_n5021), .B(new_n5018), .Y(new_n5022));
  xnor_4 g04646(.A(new_n5022), .B(new_n5015), .Y(new_n5023));
  nand_5 g04647(.A(new_n3131), .B(new_n3130), .Y(new_n5024));
  nand_5 g04648(.A(new_n3132), .B(new_n3129), .Y(new_n5025));
  nand_5 g04649(.A(new_n5025), .B(new_n5024), .Y(new_n5026));
  nand_5 g04650(.A(new_n5026), .B(new_n5019), .Y(new_n5027));
  xor_4  g04651(.A(new_n5012), .B(new_n5011), .Y(new_n5028));
  xor_4  g04652(.A(new_n5026), .B(new_n5019), .Y(new_n5029));
  nand_5 g04653(.A(new_n5029), .B(new_n5028), .Y(new_n5030));
  nand_5 g04654(.A(new_n5030), .B(new_n5027), .Y(new_n5031));
  xor_4  g04655(.A(new_n5031), .B(new_n5023), .Y(new_n5032));
  xor_4  g04656(.A(new_n5029), .B(new_n5028), .Y(new_n5033));
  nand_5 g04657(.A(pi236), .B(pi050), .Y(new_n5034));
  or_6   g04658(.A(new_n5034), .B(new_n5033), .Y(new_n5035));
  xor_4  g04659(.A(new_n5034), .B(new_n5033), .Y(new_n5036));
  or_6   g04660(.A(new_n3127), .B(new_n3120), .Y(new_n5037));
  nand_5 g04661(.A(new_n3133), .B(new_n3128), .Y(new_n5038));
  nand_5 g04662(.A(new_n5038), .B(new_n5037), .Y(new_n5039));
  nand_5 g04663(.A(new_n5039), .B(new_n5036), .Y(new_n5040));
  nand_5 g04664(.A(new_n5040), .B(new_n5035), .Y(new_n5041));
  nand_5 g04665(.A(new_n5041), .B(new_n5032), .Y(new_n5042));
  nand_5 g04666(.A(pi173), .B(pi090), .Y(new_n5043));
  nand_5 g04667(.A(pi109), .B(pi018), .Y(new_n5044));
  xor_4  g04668(.A(new_n5044), .B(new_n5043), .Y(new_n5045));
  xor_4  g04669(.A(new_n5045), .B(new_n5005), .Y(new_n5046));
  nand_5 g04670(.A(pi230), .B(pi141), .Y(new_n5047));
  xor_4  g04671(.A(new_n5047), .B(new_n5006), .Y(new_n5048));
  xor_4  g04672(.A(new_n5048), .B(new_n5046), .Y(new_n5049));
  nand_5 g04673(.A(pi253), .B(pi241), .Y(new_n5050));
  nand_5 g04674(.A(pi236), .B(pi074), .Y(new_n5051));
  xor_4  g04675(.A(new_n5051), .B(new_n5050), .Y(new_n5052));
  xor_4  g04676(.A(new_n5052), .B(new_n5020), .Y(new_n5053));
  nand_5 g04677(.A(new_n5007), .B(new_n5000), .Y(new_n5054));
  nand_5 g04678(.A(new_n5014), .B(new_n5008), .Y(new_n5055));
  nand_5 g04679(.A(new_n5055), .B(new_n5054), .Y(new_n5056));
  xor_4  g04680(.A(new_n5056), .B(new_n5053), .Y(new_n5057));
  xnor_4 g04681(.A(new_n5057), .B(new_n5049), .Y(new_n5058));
  nor_5  g04682(.A(new_n5022), .B(new_n5015), .Y(new_n5059));
  nor_5  g04683(.A(new_n5031), .B(new_n5023), .Y(new_n5060));
  xor_4  g04684(.A(new_n5060), .B(new_n5021), .Y(new_n5061));
  nor_5  g04685(.A(new_n5061), .B(new_n5059), .Y(new_n5062));
  xor_4  g04686(.A(new_n5062), .B(new_n5058), .Y(new_n5063));
  xnor_4 g04687(.A(new_n5063), .B(new_n5042), .Y(new_n5064));
  nand_5 g04688(.A(pi253), .B(pi236), .Y(new_n5065));
  nor_5  g04689(.A(new_n3181), .B(new_n3134), .Y(new_n5066));
  xor_4  g04690(.A(new_n5039), .B(new_n5036), .Y(new_n5067));
  nand_5 g04691(.A(new_n5067), .B(new_n5066), .Y(new_n5068));
  nand_5 g04692(.A(new_n5068), .B(new_n5065), .Y(new_n5069));
  xnor_4 g04693(.A(new_n5041), .B(new_n5032), .Y(new_n5070));
  xor_4  g04694(.A(new_n5068), .B(new_n5065), .Y(new_n5071));
  nand_5 g04695(.A(new_n5071), .B(new_n5070), .Y(new_n5072));
  nand_5 g04696(.A(new_n5072), .B(new_n5069), .Y(new_n5073));
  xnor_4 g04697(.A(new_n5073), .B(new_n5064), .Y(new_n5074));
  nand_5 g04698(.A(pi066), .B(pi013), .Y(new_n5075));
  nand_5 g04699(.A(pi207), .B(pi013), .Y(new_n5076));
  nand_5 g04700(.A(pi104), .B(pi066), .Y(new_n5077));
  nand_5 g04701(.A(new_n5077), .B(new_n5076), .Y(new_n5078));
  nand_5 g04702(.A(pi226), .B(pi112), .Y(new_n5079));
  xor_4  g04703(.A(new_n5077), .B(new_n5076), .Y(new_n5080));
  nand_5 g04704(.A(new_n5080), .B(new_n5079), .Y(new_n5081));
  nand_5 g04705(.A(new_n5081), .B(new_n5078), .Y(new_n5082));
  nand_5 g04706(.A(pi226), .B(pi105), .Y(new_n5083));
  nand_5 g04707(.A(pi207), .B(pi112), .Y(new_n5084));
  nand_5 g04708(.A(new_n5084), .B(new_n5083), .Y(new_n5085));
  nand_5 g04709(.A(pi207), .B(pi105), .Y(new_n5086));
  or_6   g04710(.A(new_n5086), .B(new_n5079), .Y(new_n5087));
  nand_5 g04711(.A(new_n5087), .B(new_n5085), .Y(new_n5088));
  xor_4  g04712(.A(new_n5088), .B(new_n5082), .Y(new_n5089));
  xor_4  g04713(.A(new_n5089), .B(new_n5075), .Y(new_n5090));
  nand_5 g04714(.A(pi104), .B(pi055), .Y(new_n5091));
  nand_5 g04715(.A(pi212), .B(pi002), .Y(new_n5092));
  nand_5 g04716(.A(new_n5092), .B(new_n5091), .Y(new_n5093));
  nand_5 g04717(.A(pi212), .B(pi055), .Y(new_n5094));
  nand_5 g04718(.A(pi104), .B(pi002), .Y(new_n5095));
  nor_5  g04719(.A(new_n5095), .B(new_n5094), .Y(new_n5096));
  not_8  g04720(.A(new_n5096), .Y(new_n5097));
  nand_5 g04721(.A(new_n5097), .B(new_n5093), .Y(new_n5098));
  xnor_4 g04722(.A(new_n5098), .B(new_n5090), .Y(new_n5099));
  nand_5 g04723(.A(new_n3151), .B(new_n3150), .Y(new_n5100));
  nand_5 g04724(.A(new_n3152), .B(new_n3149), .Y(new_n5101));
  nand_5 g04725(.A(new_n5101), .B(new_n5100), .Y(new_n5102));
  nand_5 g04726(.A(new_n5102), .B(new_n5094), .Y(new_n5103));
  xor_4  g04727(.A(new_n5080), .B(new_n5079), .Y(new_n5104));
  xor_4  g04728(.A(new_n5102), .B(new_n5094), .Y(new_n5105));
  nand_5 g04729(.A(new_n5105), .B(new_n5104), .Y(new_n5106));
  nand_5 g04730(.A(new_n5106), .B(new_n5103), .Y(new_n5107));
  xor_4  g04731(.A(new_n5107), .B(new_n5099), .Y(new_n5108));
  nand_5 g04732(.A(pi213), .B(pi002), .Y(new_n5109));
  nand_5 g04733(.A(new_n3157), .B(new_n3154), .Y(new_n5110));
  nand_5 g04734(.A(new_n3158), .B(new_n3153), .Y(new_n5111));
  nand_5 g04735(.A(new_n5111), .B(new_n5110), .Y(new_n5112));
  or_6   g04736(.A(new_n5112), .B(new_n5109), .Y(new_n5113));
  xor_4  g04737(.A(new_n5105), .B(new_n5104), .Y(new_n5114));
  not_8  g04738(.A(new_n5114), .Y(new_n5115));
  xor_4  g04739(.A(new_n5112), .B(new_n5109), .Y(new_n5116));
  nand_5 g04740(.A(new_n5116), .B(new_n5115), .Y(new_n5117));
  nand_5 g04741(.A(new_n5117), .B(new_n5113), .Y(new_n5118));
  nand_5 g04742(.A(new_n5118), .B(new_n5108), .Y(new_n5119));
  nand_5 g04743(.A(pi226), .B(pi183), .Y(new_n5120));
  nand_5 g04744(.A(pi112), .B(pi066), .Y(new_n5121));
  xor_4  g04745(.A(new_n5121), .B(new_n5120), .Y(new_n5122));
  xor_4  g04746(.A(new_n5122), .B(new_n5086), .Y(new_n5123));
  nand_5 g04747(.A(pi055), .B(pi013), .Y(new_n5124));
  xor_4  g04748(.A(new_n5124), .B(new_n5087), .Y(new_n5125));
  xor_4  g04749(.A(new_n5125), .B(new_n5123), .Y(new_n5126));
  nand_5 g04750(.A(pi212), .B(pi025), .Y(new_n5127));
  nand_5 g04751(.A(pi239), .B(pi213), .Y(new_n5128));
  xor_4  g04752(.A(new_n5128), .B(new_n5127), .Y(new_n5129));
  xor_4  g04753(.A(new_n5129), .B(new_n5095), .Y(new_n5130));
  nand_5 g04754(.A(new_n5088), .B(new_n5082), .Y(new_n5131));
  nand_5 g04755(.A(new_n5089), .B(new_n5075), .Y(new_n5132));
  nand_5 g04756(.A(new_n5132), .B(new_n5131), .Y(new_n5133));
  xor_4  g04757(.A(new_n5133), .B(new_n5130), .Y(new_n5134));
  xnor_4 g04758(.A(new_n5134), .B(new_n5126), .Y(new_n5135));
  nor_5  g04759(.A(new_n5107), .B(new_n5099), .Y(new_n5136));
  and_6  g04760(.A(new_n5136), .B(new_n5096), .Y(new_n5137));
  or_6   g04761(.A(new_n5098), .B(new_n5090), .Y(new_n5138));
  nand_5 g04762(.A(new_n5138), .B(new_n5097), .Y(new_n5139));
  nor_5  g04763(.A(new_n5139), .B(new_n5136), .Y(new_n5140));
  or_6   g04764(.A(new_n5140), .B(new_n5137), .Y(new_n5141));
  xor_4  g04765(.A(new_n5141), .B(new_n5135), .Y(new_n5142));
  xor_4  g04766(.A(new_n5142), .B(new_n5119), .Y(new_n5143));
  nand_5 g04767(.A(pi213), .B(pi025), .Y(new_n5144));
  xnor_4 g04768(.A(new_n5118), .B(new_n5108), .Y(new_n5145));
  or_6   g04769(.A(new_n5145), .B(new_n5144), .Y(new_n5146));
  nand_5 g04770(.A(new_n3160), .B(new_n3148), .Y(new_n5147));
  xor_4  g04771(.A(new_n5116), .B(new_n5114), .Y(new_n5148));
  nor_5  g04772(.A(new_n5148), .B(new_n5147), .Y(new_n5149));
  xor_4  g04773(.A(new_n5145), .B(new_n5144), .Y(new_n5150));
  nand_5 g04774(.A(new_n5150), .B(new_n5149), .Y(new_n5151));
  nand_5 g04775(.A(new_n5151), .B(new_n5146), .Y(new_n5152));
  xor_4  g04776(.A(new_n5152), .B(new_n5143), .Y(new_n5153));
  xor_4  g04777(.A(new_n5153), .B(new_n5074), .Y(new_n5154));
  xnor_4 g04778(.A(new_n5071), .B(new_n5070), .Y(new_n5155));
  xor_4  g04779(.A(new_n5150), .B(new_n5149), .Y(new_n5156));
  nand_5 g04780(.A(new_n5156), .B(new_n5155), .Y(new_n5157));
  xor_4  g04781(.A(new_n5156), .B(new_n5155), .Y(new_n5158));
  xor_4  g04782(.A(new_n5067), .B(new_n5066), .Y(new_n5159));
  xor_4  g04783(.A(new_n5148), .B(new_n5147), .Y(new_n5160));
  nand_5 g04784(.A(new_n5160), .B(new_n5159), .Y(new_n5161));
  xor_4  g04785(.A(new_n5160), .B(new_n5159), .Y(new_n5162));
  not_8  g04786(.A(new_n3161), .Y(new_n5163));
  nor_5  g04787(.A(new_n5163), .B(new_n3139), .Y(new_n5164));
  nor_5  g04788(.A(new_n3186), .B(new_n3162), .Y(new_n5165));
  nor_5  g04789(.A(new_n5165), .B(new_n5164), .Y(new_n5166));
  not_8  g04790(.A(new_n5166), .Y(new_n5167));
  nand_5 g04791(.A(new_n5167), .B(new_n5162), .Y(new_n5168));
  nand_5 g04792(.A(new_n5168), .B(new_n5161), .Y(new_n5169));
  nand_5 g04793(.A(new_n5169), .B(new_n5158), .Y(new_n5170));
  nand_5 g04794(.A(new_n5170), .B(new_n5157), .Y(new_n5171));
  xnor_4 g04795(.A(new_n5171), .B(new_n5154), .Y(new_n5172));
  nand_5 g04796(.A(pi058), .B(pi035), .Y(new_n5173));
  nand_5 g04797(.A(pi204), .B(pi132), .Y(new_n5174));
  nand_5 g04798(.A(pi186), .B(pi015), .Y(new_n5175));
  nand_5 g04799(.A(new_n5175), .B(new_n5174), .Y(new_n5176));
  nand_5 g04800(.A(pi132), .B(pi015), .Y(new_n5177));
  nand_5 g04801(.A(pi204), .B(pi186), .Y(new_n5178));
  or_6   g04802(.A(new_n5178), .B(new_n5177), .Y(new_n5179));
  nand_5 g04803(.A(new_n5179), .B(new_n5176), .Y(new_n5180));
  xor_4  g04804(.A(new_n5180), .B(new_n5173), .Y(new_n5181));
  nand_5 g04805(.A(pi186), .B(pi035), .Y(new_n5182));
  nand_5 g04806(.A(new_n5182), .B(new_n5177), .Y(new_n5183));
  nand_5 g04807(.A(pi139), .B(pi058), .Y(new_n5184));
  xor_4  g04808(.A(new_n5182), .B(new_n5177), .Y(new_n5185));
  nand_5 g04809(.A(new_n5185), .B(new_n5184), .Y(new_n5186));
  nand_5 g04810(.A(new_n5186), .B(new_n5183), .Y(new_n5187));
  xor_4  g04811(.A(new_n5187), .B(new_n5181), .Y(new_n5188));
  nand_5 g04812(.A(pi211), .B(pi139), .Y(new_n5189));
  nand_5 g04813(.A(pi208), .B(pi199), .Y(new_n5190));
  and_6  g04814(.A(new_n5190), .B(new_n5189), .Y(new_n5191));
  nand_5 g04815(.A(pi211), .B(pi208), .Y(new_n5192));
  nand_5 g04816(.A(pi199), .B(pi139), .Y(new_n5193));
  nor_5  g04817(.A(new_n5193), .B(new_n5192), .Y(new_n5194));
  or_6   g04818(.A(new_n5194), .B(new_n5191), .Y(new_n5195));
  xnor_4 g04819(.A(new_n5195), .B(new_n5188), .Y(new_n5196));
  nand_5 g04820(.A(new_n3203), .B(new_n3202), .Y(new_n5197));
  nand_5 g04821(.A(new_n3204), .B(new_n3201), .Y(new_n5198));
  nand_5 g04822(.A(new_n5198), .B(new_n5197), .Y(new_n5199));
  nand_5 g04823(.A(new_n5199), .B(new_n5192), .Y(new_n5200));
  xor_4  g04824(.A(new_n5185), .B(new_n5184), .Y(new_n5201));
  xor_4  g04825(.A(new_n5199), .B(new_n5192), .Y(new_n5202));
  nand_5 g04826(.A(new_n5202), .B(new_n5201), .Y(new_n5203));
  nand_5 g04827(.A(new_n5203), .B(new_n5200), .Y(new_n5204));
  xor_4  g04828(.A(new_n5204), .B(new_n5196), .Y(new_n5205));
  xor_4  g04829(.A(new_n5202), .B(new_n5201), .Y(new_n5206));
  nand_5 g04830(.A(pi199), .B(pi168), .Y(new_n5207));
  or_6   g04831(.A(new_n5207), .B(new_n5206), .Y(new_n5208));
  xor_4  g04832(.A(new_n5207), .B(new_n5206), .Y(new_n5209));
  or_6   g04833(.A(new_n3199), .B(new_n3196), .Y(new_n5210));
  nand_5 g04834(.A(new_n3205), .B(new_n3200), .Y(new_n5211));
  nand_5 g04835(.A(new_n5211), .B(new_n5210), .Y(new_n5212));
  nand_5 g04836(.A(new_n5212), .B(new_n5209), .Y(new_n5213));
  nand_5 g04837(.A(new_n5213), .B(new_n5208), .Y(new_n5214));
  nand_5 g04838(.A(new_n5214), .B(new_n5205), .Y(new_n5215));
  nand_5 g04839(.A(pi146), .B(pi132), .Y(new_n5216));
  nand_5 g04840(.A(pi058), .B(pi015), .Y(new_n5217));
  xor_4  g04841(.A(new_n5217), .B(new_n5216), .Y(new_n5218));
  xor_4  g04842(.A(new_n5218), .B(new_n5178), .Y(new_n5219));
  nand_5 g04843(.A(pi211), .B(pi035), .Y(new_n5220));
  xor_4  g04844(.A(new_n5220), .B(new_n5179), .Y(new_n5221));
  xor_4  g04845(.A(new_n5221), .B(new_n5219), .Y(new_n5222));
  nand_5 g04846(.A(pi208), .B(pi195), .Y(new_n5223));
  nand_5 g04847(.A(pi218), .B(pi168), .Y(new_n5224));
  xor_4  g04848(.A(new_n5224), .B(new_n5223), .Y(new_n5225));
  xor_4  g04849(.A(new_n5225), .B(new_n5193), .Y(new_n5226));
  nand_5 g04850(.A(new_n5180), .B(new_n5173), .Y(new_n5227));
  nand_5 g04851(.A(new_n5187), .B(new_n5181), .Y(new_n5228));
  nand_5 g04852(.A(new_n5228), .B(new_n5227), .Y(new_n5229));
  xor_4  g04853(.A(new_n5229), .B(new_n5226), .Y(new_n5230));
  xnor_4 g04854(.A(new_n5230), .B(new_n5222), .Y(new_n5231));
  nor_5  g04855(.A(new_n5195), .B(new_n5188), .Y(new_n5232));
  nor_5  g04856(.A(new_n5204), .B(new_n5196), .Y(new_n5233));
  xor_4  g04857(.A(new_n5233), .B(new_n5194), .Y(new_n5234));
  nor_5  g04858(.A(new_n5234), .B(new_n5232), .Y(new_n5235));
  xor_4  g04859(.A(new_n5235), .B(new_n5231), .Y(new_n5236));
  nand_5 g04860(.A(pi195), .B(pi168), .Y(new_n5237));
  nor_5  g04861(.A(new_n3206), .B(new_n3195), .Y(new_n5238));
  xor_4  g04862(.A(new_n5212), .B(new_n5209), .Y(new_n5239));
  nand_5 g04863(.A(new_n5239), .B(new_n5238), .Y(new_n5240));
  nand_5 g04864(.A(new_n5240), .B(new_n5237), .Y(new_n5241));
  xnor_4 g04865(.A(new_n5214), .B(new_n5205), .Y(new_n5242));
  xor_4  g04866(.A(new_n5240), .B(new_n5237), .Y(new_n5243));
  nand_5 g04867(.A(new_n5243), .B(new_n5242), .Y(new_n5244));
  nand_5 g04868(.A(new_n5244), .B(new_n5241), .Y(new_n5245));
  xor_4  g04869(.A(new_n5245), .B(new_n5236), .Y(new_n5246));
  xor_4  g04870(.A(new_n5246), .B(new_n5215), .Y(new_n5247));
  xor_4  g04871(.A(new_n5247), .B(new_n5172), .Y(new_n5248));
  xor_4  g04872(.A(new_n5169), .B(new_n5158), .Y(new_n5249));
  not_8  g04873(.A(new_n5249), .Y(new_n5250));
  xor_4  g04874(.A(new_n5243), .B(new_n5242), .Y(new_n5251));
  or_6   g04875(.A(new_n5251), .B(new_n5250), .Y(new_n5252));
  xor_4  g04876(.A(new_n5251), .B(new_n5250), .Y(new_n5253));
  xor_4  g04877(.A(new_n5167), .B(new_n5162), .Y(new_n5254));
  xor_4  g04878(.A(new_n5239), .B(new_n5238), .Y(new_n5255));
  nand_5 g04879(.A(new_n5255), .B(new_n5254), .Y(new_n5256));
  not_8  g04880(.A(new_n5256), .Y(new_n5257));
  xnor_4 g04881(.A(new_n5255), .B(new_n5254), .Y(new_n5258));
  or_6   g04882(.A(new_n3226), .B(new_n3207), .Y(new_n5259));
  not_8  g04883(.A(new_n3187), .Y(new_n5260));
  nand_5 g04884(.A(new_n3227), .B(new_n5260), .Y(new_n5261));
  nand_5 g04885(.A(new_n5261), .B(new_n5259), .Y(new_n5262));
  nor_5  g04886(.A(new_n5262), .B(new_n5258), .Y(new_n5263));
  nor_5  g04887(.A(new_n5263), .B(new_n5257), .Y(new_n5264));
  not_8  g04888(.A(new_n5264), .Y(new_n5265));
  nand_5 g04889(.A(new_n5265), .B(new_n5253), .Y(new_n5266));
  nand_5 g04890(.A(new_n5266), .B(new_n5252), .Y(new_n5267));
  xnor_4 g04891(.A(new_n5267), .B(new_n5248), .Y(new_n5268));
  nand_5 g04892(.A(pi244), .B(pi133), .Y(new_n5269));
  nand_5 g04893(.A(pi189), .B(pi069), .Y(new_n5270));
  nand_5 g04894(.A(pi064), .B(pi029), .Y(new_n5271));
  nand_5 g04895(.A(new_n5271), .B(new_n5270), .Y(new_n5272));
  nand_5 g04896(.A(pi189), .B(pi029), .Y(new_n5273));
  nand_5 g04897(.A(pi069), .B(pi064), .Y(new_n5274));
  or_6   g04898(.A(new_n5274), .B(new_n5273), .Y(new_n5275));
  nand_5 g04899(.A(new_n5275), .B(new_n5272), .Y(new_n5276));
  xor_4  g04900(.A(new_n5276), .B(new_n5269), .Y(new_n5277));
  nand_5 g04901(.A(pi244), .B(pi077), .Y(new_n5278));
  nand_5 g04902(.A(pi133), .B(pi069), .Y(new_n5279));
  nand_5 g04903(.A(new_n5279), .B(new_n5278), .Y(new_n5280));
  xor_4  g04904(.A(new_n5279), .B(new_n5278), .Y(new_n5281));
  nand_5 g04905(.A(new_n5281), .B(new_n5273), .Y(new_n5282));
  nand_5 g04906(.A(new_n5282), .B(new_n5280), .Y(new_n5283));
  xor_4  g04907(.A(new_n5283), .B(new_n5277), .Y(new_n5284));
  nand_5 g04908(.A(pi150), .B(pi077), .Y(new_n5285));
  nand_5 g04909(.A(pi221), .B(pi052), .Y(new_n5286));
  and_6  g04910(.A(new_n5286), .B(new_n5285), .Y(new_n5287));
  nand_5 g04911(.A(pi150), .B(pi052), .Y(new_n5288));
  nand_5 g04912(.A(pi221), .B(pi077), .Y(new_n5289));
  nor_5  g04913(.A(new_n5289), .B(new_n5288), .Y(new_n5290));
  or_6   g04914(.A(new_n5290), .B(new_n5287), .Y(new_n5291));
  xnor_4 g04915(.A(new_n5291), .B(new_n5284), .Y(new_n5292));
  nand_5 g04916(.A(new_n3240), .B(new_n3239), .Y(new_n5293));
  nand_5 g04917(.A(new_n3241), .B(new_n3238), .Y(new_n5294));
  nand_5 g04918(.A(new_n5294), .B(new_n5293), .Y(new_n5295));
  nand_5 g04919(.A(new_n5295), .B(new_n5288), .Y(new_n5296));
  xor_4  g04920(.A(new_n5281), .B(new_n5273), .Y(new_n5297));
  xor_4  g04921(.A(new_n5295), .B(new_n5288), .Y(new_n5298));
  nand_5 g04922(.A(new_n5298), .B(new_n5297), .Y(new_n5299));
  nand_5 g04923(.A(new_n5299), .B(new_n5296), .Y(new_n5300));
  xor_4  g04924(.A(new_n5300), .B(new_n5292), .Y(new_n5301));
  nand_5 g04925(.A(pi221), .B(pi131), .Y(new_n5302));
  nand_5 g04926(.A(new_n3246), .B(new_n3243), .Y(new_n5303));
  nand_5 g04927(.A(new_n3247), .B(new_n3242), .Y(new_n5304));
  nand_5 g04928(.A(new_n5304), .B(new_n5303), .Y(new_n5305));
  or_6   g04929(.A(new_n5305), .B(new_n5302), .Y(new_n5306));
  xnor_4 g04930(.A(new_n5298), .B(new_n5297), .Y(new_n5307));
  xor_4  g04931(.A(new_n5305), .B(new_n5302), .Y(new_n5308));
  nand_5 g04932(.A(new_n5308), .B(new_n5307), .Y(new_n5309));
  nand_5 g04933(.A(new_n5309), .B(new_n5306), .Y(new_n5310));
  nand_5 g04934(.A(new_n5310), .B(new_n5301), .Y(new_n5311));
  nand_5 g04935(.A(pi084), .B(pi029), .Y(new_n5312));
  nand_5 g04936(.A(pi244), .B(pi189), .Y(new_n5313));
  xor_4  g04937(.A(new_n5313), .B(new_n5312), .Y(new_n5314));
  xor_4  g04938(.A(new_n5314), .B(new_n5274), .Y(new_n5315));
  nand_5 g04939(.A(pi150), .B(pi133), .Y(new_n5316));
  xor_4  g04940(.A(new_n5316), .B(new_n5275), .Y(new_n5317));
  xor_4  g04941(.A(new_n5317), .B(new_n5315), .Y(new_n5318));
  nand_5 g04942(.A(pi196), .B(pi052), .Y(new_n5319));
  nand_5 g04943(.A(pi184), .B(pi131), .Y(new_n5320));
  xor_4  g04944(.A(new_n5320), .B(new_n5319), .Y(new_n5321));
  xor_4  g04945(.A(new_n5321), .B(new_n5289), .Y(new_n5322));
  nand_5 g04946(.A(new_n5276), .B(new_n5269), .Y(new_n5323));
  nand_5 g04947(.A(new_n5283), .B(new_n5277), .Y(new_n5324));
  nand_5 g04948(.A(new_n5324), .B(new_n5323), .Y(new_n5325));
  xor_4  g04949(.A(new_n5325), .B(new_n5322), .Y(new_n5326));
  xnor_4 g04950(.A(new_n5326), .B(new_n5318), .Y(new_n5327));
  nor_5  g04951(.A(new_n5291), .B(new_n5284), .Y(new_n5328));
  nor_5  g04952(.A(new_n5300), .B(new_n5292), .Y(new_n5329));
  xor_4  g04953(.A(new_n5329), .B(new_n5290), .Y(new_n5330));
  nor_5  g04954(.A(new_n5330), .B(new_n5328), .Y(new_n5331));
  not_8  g04955(.A(new_n5331), .Y(new_n5332));
  xor_4  g04956(.A(new_n5332), .B(new_n5327), .Y(new_n5333));
  xor_4  g04957(.A(new_n5333), .B(new_n5311), .Y(new_n5334));
  nand_5 g04958(.A(pi196), .B(pi131), .Y(new_n5335));
  not_8  g04959(.A(new_n3237), .Y(new_n5336));
  nor_5  g04960(.A(new_n3248), .B(new_n5336), .Y(new_n5337));
  xor_4  g04961(.A(new_n5308), .B(new_n5307), .Y(new_n5338));
  nand_5 g04962(.A(new_n5338), .B(new_n5337), .Y(new_n5339));
  nand_5 g04963(.A(new_n5339), .B(new_n5335), .Y(new_n5340));
  xor_4  g04964(.A(new_n5310), .B(new_n5301), .Y(new_n5341));
  not_8  g04965(.A(new_n5341), .Y(new_n5342));
  xor_4  g04966(.A(new_n5339), .B(new_n5335), .Y(new_n5343));
  nand_5 g04967(.A(new_n5343), .B(new_n5342), .Y(new_n5344));
  nand_5 g04968(.A(new_n5344), .B(new_n5340), .Y(new_n5345));
  xor_4  g04969(.A(new_n5345), .B(new_n5334), .Y(new_n5346));
  xor_4  g04970(.A(new_n5346), .B(new_n5268), .Y(new_n5347));
  xor_4  g04971(.A(new_n5264), .B(new_n5253), .Y(new_n5348));
  xor_4  g04972(.A(new_n5338), .B(new_n5337), .Y(new_n5349));
  or_6   g04973(.A(new_n3268), .B(new_n3249), .Y(new_n5350));
  nand_5 g04974(.A(new_n3269), .B(new_n3228), .Y(new_n5351));
  nand_5 g04975(.A(new_n5351), .B(new_n5350), .Y(new_n5352));
  or_6   g04976(.A(new_n5352), .B(new_n5349), .Y(new_n5353));
  xor_4  g04977(.A(new_n5262), .B(new_n5258), .Y(new_n5354));
  not_8  g04978(.A(new_n5354), .Y(new_n5355));
  xor_4  g04979(.A(new_n5352), .B(new_n5349), .Y(new_n5356));
  nand_5 g04980(.A(new_n5356), .B(new_n5355), .Y(new_n5357));
  nand_5 g04981(.A(new_n5357), .B(new_n5353), .Y(new_n5358));
  or_6   g04982(.A(new_n5358), .B(new_n5348), .Y(new_n5359));
  xor_4  g04983(.A(new_n5343), .B(new_n5341), .Y(new_n5360));
  xor_4  g04984(.A(new_n5358), .B(new_n5348), .Y(new_n5361));
  nand_5 g04985(.A(new_n5361), .B(new_n5360), .Y(new_n5362));
  nand_5 g04986(.A(new_n5362), .B(new_n5359), .Y(new_n5363));
  xor_4  g04987(.A(new_n5363), .B(new_n5347), .Y(po019));
  xor_4  g04988(.A(new_n3266), .B(new_n3264), .Y(po020));
  nand_5 g04989(.A(pi087), .B(pi028), .Y(new_n5366));
  nand_5 g04990(.A(pi113), .B(pi102), .Y(new_n5367));
  nand_5 g04991(.A(pi007), .B(pi001), .Y(new_n5368));
  nand_5 g04992(.A(pi122), .B(pi051), .Y(new_n5369));
  nand_5 g04993(.A(pi135), .B(pi042), .Y(new_n5370));
  or_6   g04994(.A(new_n5370), .B(new_n5369), .Y(new_n5371));
  or_6   g04995(.A(new_n5371), .B(new_n5368), .Y(new_n5372));
  nand_5 g04996(.A(pi059), .B(pi051), .Y(new_n5373));
  nand_5 g04997(.A(pi122), .B(pi108), .Y(new_n5374));
  xor_4  g04998(.A(new_n5374), .B(new_n5373), .Y(new_n5375));
  xor_4  g04999(.A(new_n5375), .B(new_n5370), .Y(new_n5376));
  not_8  g05000(.A(new_n5376), .Y(new_n5377));
  xor_4  g05001(.A(new_n5371), .B(new_n5368), .Y(new_n5378));
  nand_5 g05002(.A(new_n5378), .B(new_n5377), .Y(new_n5379));
  nand_5 g05003(.A(new_n5379), .B(new_n5372), .Y(new_n5380));
  xor_4  g05004(.A(new_n5380), .B(new_n5367), .Y(new_n5381));
  nand_5 g05005(.A(pi180), .B(pi060), .Y(new_n5382));
  nand_5 g05006(.A(pi085), .B(pi020), .Y(new_n5383));
  nor_5  g05007(.A(new_n5383), .B(new_n5382), .Y(new_n5384));
  nand_5 g05008(.A(pi223), .B(pi194), .Y(new_n5385));
  nand_5 g05009(.A(pi225), .B(pi143), .Y(new_n5386));
  nand_5 g05010(.A(pi101), .B(pi057), .Y(new_n5387));
  nand_5 g05011(.A(new_n5387), .B(new_n5386), .Y(new_n5388));
  nand_5 g05012(.A(pi143), .B(pi101), .Y(new_n5389));
  nand_5 g05013(.A(pi225), .B(pi057), .Y(new_n5390));
  or_6   g05014(.A(new_n5390), .B(new_n5389), .Y(new_n5391));
  nand_5 g05015(.A(new_n5391), .B(new_n5388), .Y(new_n5392));
  xor_4  g05016(.A(new_n5392), .B(new_n5385), .Y(new_n5393));
  nand_5 g05017(.A(pi223), .B(pi057), .Y(new_n5394));
  nand_5 g05018(.A(new_n5394), .B(new_n5389), .Y(new_n5395));
  nand_5 g05019(.A(pi194), .B(pi060), .Y(new_n5396));
  xor_4  g05020(.A(new_n5394), .B(new_n5389), .Y(new_n5397));
  nand_5 g05021(.A(new_n5397), .B(new_n5396), .Y(new_n5398));
  nand_5 g05022(.A(new_n5398), .B(new_n5395), .Y(new_n5399));
  xor_4  g05023(.A(new_n5399), .B(new_n5393), .Y(new_n5400));
  nand_5 g05024(.A(pi180), .B(pi020), .Y(new_n5401));
  nand_5 g05025(.A(pi085), .B(pi060), .Y(new_n5402));
  and_6  g05026(.A(new_n5402), .B(new_n5401), .Y(new_n5403));
  or_6   g05027(.A(new_n5403), .B(new_n5384), .Y(new_n5404));
  xnor_4 g05028(.A(new_n5404), .B(new_n5400), .Y(new_n5405));
  nand_5 g05029(.A(new_n4930), .B(new_n4929), .Y(new_n5406));
  nand_5 g05030(.A(new_n4931), .B(new_n4928), .Y(new_n5407));
  nand_5 g05031(.A(new_n5407), .B(new_n5406), .Y(new_n5408));
  nand_5 g05032(.A(new_n5408), .B(new_n5383), .Y(new_n5409));
  xor_4  g05033(.A(new_n5397), .B(new_n5396), .Y(new_n5410));
  xor_4  g05034(.A(new_n5408), .B(new_n5383), .Y(new_n5411));
  nand_5 g05035(.A(new_n5411), .B(new_n5410), .Y(new_n5412));
  nand_5 g05036(.A(new_n5412), .B(new_n5409), .Y(new_n5413));
  nor_5  g05037(.A(new_n5413), .B(new_n5405), .Y(new_n5414));
  nand_5 g05038(.A(new_n5414), .B(new_n5384), .Y(new_n5415));
  nand_5 g05039(.A(pi177), .B(pi143), .Y(new_n5416));
  nand_5 g05040(.A(pi194), .B(pi101), .Y(new_n5417));
  xor_4  g05041(.A(new_n5417), .B(new_n5416), .Y(new_n5418));
  xor_4  g05042(.A(new_n5418), .B(new_n5390), .Y(new_n5419));
  nand_5 g05043(.A(pi223), .B(pi085), .Y(new_n5420));
  xor_4  g05044(.A(new_n5420), .B(new_n5391), .Y(new_n5421));
  not_8  g05045(.A(new_n5421), .Y(new_n5422));
  xor_4  g05046(.A(new_n5422), .B(new_n5419), .Y(new_n5423));
  nand_5 g05047(.A(pi160), .B(pi068), .Y(new_n5424));
  nand_5 g05048(.A(pi036), .B(pi020), .Y(new_n5425));
  xor_4  g05049(.A(new_n5425), .B(new_n5424), .Y(new_n5426));
  xor_4  g05050(.A(new_n5426), .B(new_n5382), .Y(new_n5427));
  nand_5 g05051(.A(new_n5392), .B(new_n5385), .Y(new_n5428));
  nand_5 g05052(.A(new_n5399), .B(new_n5393), .Y(new_n5429));
  nand_5 g05053(.A(new_n5429), .B(new_n5428), .Y(new_n5430));
  xor_4  g05054(.A(new_n5430), .B(new_n5427), .Y(new_n5431));
  xor_4  g05055(.A(new_n5431), .B(new_n5423), .Y(new_n5432));
  nor_5  g05056(.A(new_n5404), .B(new_n5400), .Y(new_n5433));
  xor_4  g05057(.A(new_n5414), .B(new_n5384), .Y(new_n5434));
  nor_5  g05058(.A(new_n5434), .B(new_n5433), .Y(new_n5435));
  not_8  g05059(.A(new_n5435), .Y(new_n5436));
  nand_5 g05060(.A(new_n5436), .B(new_n5432), .Y(new_n5437));
  nand_5 g05061(.A(new_n5437), .B(new_n5415), .Y(new_n5438));
  nand_5 g05062(.A(pi143), .B(pi137), .Y(new_n5439));
  nand_5 g05063(.A(pi160), .B(pi046), .Y(new_n5440));
  xnor_4 g05064(.A(new_n5440), .B(new_n5439), .Y(new_n5441));
  xor_4  g05065(.A(new_n5441), .B(new_n5438), .Y(new_n5442));
  nand_5 g05066(.A(new_n5374), .B(new_n5373), .Y(new_n5443));
  nand_5 g05067(.A(new_n5375), .B(new_n5370), .Y(new_n5444));
  nand_5 g05068(.A(new_n5444), .B(new_n5443), .Y(new_n5445));
  xor_4  g05069(.A(new_n5435), .B(new_n5432), .Y(new_n5446));
  nand_5 g05070(.A(pi160), .B(pi036), .Y(new_n5447));
  not_8  g05071(.A(new_n4927), .Y(new_n5448));
  nor_5  g05072(.A(new_n4938), .B(new_n5448), .Y(new_n5449));
  xor_4  g05073(.A(new_n5411), .B(new_n5410), .Y(new_n5450));
  nand_5 g05074(.A(pi180), .B(pi160), .Y(new_n5451));
  xnor_4 g05075(.A(new_n5451), .B(new_n5450), .Y(new_n5452));
  nand_5 g05076(.A(new_n4936), .B(new_n4933), .Y(new_n5453));
  nand_5 g05077(.A(new_n4937), .B(new_n4932), .Y(new_n5454));
  nand_5 g05078(.A(new_n5454), .B(new_n5453), .Y(new_n5455));
  xor_4  g05079(.A(new_n5455), .B(new_n5452), .Y(new_n5456));
  nand_5 g05080(.A(new_n5456), .B(new_n5449), .Y(new_n5457));
  nand_5 g05081(.A(new_n5457), .B(new_n5447), .Y(new_n5458));
  xor_4  g05082(.A(new_n5413), .B(new_n5405), .Y(new_n5459));
  nor_5  g05083(.A(new_n5451), .B(new_n5450), .Y(new_n5460));
  nor_5  g05084(.A(new_n5455), .B(new_n5452), .Y(new_n5461));
  nor_5  g05085(.A(new_n5461), .B(new_n5460), .Y(new_n5462));
  xor_4  g05086(.A(new_n5462), .B(new_n5459), .Y(new_n5463));
  xor_4  g05087(.A(new_n5457), .B(new_n5447), .Y(new_n5464));
  nand_5 g05088(.A(new_n5464), .B(new_n5463), .Y(new_n5465));
  nand_5 g05089(.A(new_n5465), .B(new_n5458), .Y(new_n5466));
  nand_5 g05090(.A(new_n5466), .B(new_n5446), .Y(new_n5467));
  not_8  g05091(.A(new_n5462), .Y(new_n5468));
  nand_5 g05092(.A(new_n5468), .B(new_n5459), .Y(new_n5469));
  xor_4  g05093(.A(new_n5466), .B(new_n5446), .Y(new_n5470));
  nand_5 g05094(.A(new_n5470), .B(new_n5469), .Y(new_n5471));
  nand_5 g05095(.A(new_n5471), .B(new_n5467), .Y(new_n5472));
  xor_4  g05096(.A(new_n5472), .B(new_n5445), .Y(new_n5473));
  xor_4  g05097(.A(new_n5473), .B(new_n5442), .Y(new_n5474));
  nand_5 g05098(.A(pi219), .B(pi038), .Y(new_n5475));
  nand_5 g05099(.A(pi087), .B(pi038), .Y(new_n5476));
  nand_5 g05100(.A(pi219), .B(pi113), .Y(new_n5477));
  nand_5 g05101(.A(new_n5477), .B(new_n5476), .Y(new_n5478));
  nand_5 g05102(.A(pi118), .B(pi102), .Y(new_n5479));
  xor_4  g05103(.A(new_n5477), .B(new_n5476), .Y(new_n5480));
  nand_5 g05104(.A(new_n5480), .B(new_n5479), .Y(new_n5481));
  nand_5 g05105(.A(new_n5481), .B(new_n5478), .Y(new_n5482));
  xor_4  g05106(.A(new_n5480), .B(new_n5479), .Y(new_n5483));
  nand_5 g05107(.A(pi108), .B(pi001), .Y(new_n5484));
  nand_5 g05108(.A(pi122), .B(pi042), .Y(new_n5485));
  nand_5 g05109(.A(pi135), .B(pi051), .Y(new_n5486));
  nand_5 g05110(.A(new_n5486), .B(new_n5485), .Y(new_n5487));
  nand_5 g05111(.A(new_n5487), .B(new_n5371), .Y(new_n5488));
  nand_5 g05112(.A(new_n5488), .B(new_n5484), .Y(new_n5489));
  xor_4  g05113(.A(new_n5488), .B(new_n5484), .Y(new_n5490));
  nand_5 g05114(.A(pi108), .B(pi102), .Y(new_n5491));
  nand_5 g05115(.A(pi042), .B(pi001), .Y(new_n5492));
  nand_5 g05116(.A(new_n5492), .B(new_n5491), .Y(new_n5493));
  xor_4  g05117(.A(new_n5492), .B(new_n5491), .Y(new_n5494));
  nand_5 g05118(.A(new_n5494), .B(new_n5369), .Y(new_n5495));
  nand_5 g05119(.A(new_n5495), .B(new_n5493), .Y(new_n5496));
  nand_5 g05120(.A(new_n5496), .B(new_n5490), .Y(new_n5497));
  nand_5 g05121(.A(new_n5497), .B(new_n5489), .Y(new_n5498));
  or_6   g05122(.A(new_n5498), .B(new_n5483), .Y(new_n5499));
  xor_4  g05123(.A(new_n5378), .B(new_n5377), .Y(new_n5500));
  xor_4  g05124(.A(new_n5498), .B(new_n5483), .Y(new_n5501));
  nand_5 g05125(.A(new_n5501), .B(new_n5500), .Y(new_n5502));
  nand_5 g05126(.A(new_n5502), .B(new_n5499), .Y(new_n5503));
  xor_4  g05127(.A(new_n5503), .B(new_n5482), .Y(new_n5504));
  xor_4  g05128(.A(new_n5470), .B(new_n5469), .Y(new_n5505));
  xor_4  g05129(.A(new_n5464), .B(new_n5463), .Y(new_n5506));
  nand_5 g05130(.A(pi182), .B(pi048), .Y(new_n5507));
  nand_5 g05131(.A(new_n4892), .B(new_n4891), .Y(new_n5508));
  nand_5 g05132(.A(new_n4893), .B(new_n4890), .Y(new_n5509));
  nand_5 g05133(.A(new_n5509), .B(new_n5508), .Y(new_n5510));
  nand_5 g05134(.A(new_n5510), .B(new_n5507), .Y(new_n5511));
  nand_5 g05135(.A(pi162), .B(pi076), .Y(new_n5512));
  nand_5 g05136(.A(pi216), .B(pi033), .Y(new_n5513));
  nand_5 g05137(.A(pi179), .B(pi041), .Y(new_n5514));
  xor_4  g05138(.A(new_n5514), .B(new_n5513), .Y(new_n5515));
  xor_4  g05139(.A(new_n5515), .B(new_n5512), .Y(new_n5516));
  xor_4  g05140(.A(new_n5510), .B(new_n5507), .Y(new_n5517));
  nand_5 g05141(.A(new_n5517), .B(new_n5516), .Y(new_n5518));
  nand_5 g05142(.A(new_n5518), .B(new_n5511), .Y(new_n5519));
  nand_5 g05143(.A(pi216), .B(pi179), .Y(new_n5520));
  nand_5 g05144(.A(pi076), .B(pi033), .Y(new_n5521));
  nand_5 g05145(.A(pi162), .B(pi079), .Y(new_n5522));
  nand_5 g05146(.A(new_n5522), .B(new_n5521), .Y(new_n5523));
  nand_5 g05147(.A(pi079), .B(pi033), .Y(new_n5524));
  or_6   g05148(.A(new_n5524), .B(new_n5512), .Y(new_n5525));
  nand_5 g05149(.A(new_n5525), .B(new_n5523), .Y(new_n5526));
  xor_4  g05150(.A(new_n5526), .B(new_n5520), .Y(new_n5527));
  nand_5 g05151(.A(new_n5514), .B(new_n5513), .Y(new_n5528));
  nand_5 g05152(.A(new_n5515), .B(new_n5512), .Y(new_n5529));
  nand_5 g05153(.A(new_n5529), .B(new_n5528), .Y(new_n5530));
  xor_4  g05154(.A(new_n5530), .B(new_n5527), .Y(new_n5531));
  nand_5 g05155(.A(pi048), .B(pi041), .Y(new_n5532));
  nand_5 g05156(.A(pi237), .B(pi182), .Y(new_n5533));
  nand_5 g05157(.A(new_n5533), .B(new_n5532), .Y(new_n5534));
  nand_5 g05158(.A(pi237), .B(pi041), .Y(new_n5535));
  or_6   g05159(.A(new_n5535), .B(new_n5507), .Y(new_n5536));
  nand_5 g05160(.A(new_n5536), .B(new_n5534), .Y(new_n5537));
  xor_4  g05161(.A(new_n5537), .B(new_n5531), .Y(new_n5538));
  xnor_4 g05162(.A(new_n5538), .B(new_n5519), .Y(new_n5539));
  xor_4  g05163(.A(new_n5517), .B(new_n5516), .Y(new_n5540));
  nand_5 g05164(.A(pi237), .B(pi138), .Y(new_n5541));
  nor_5  g05165(.A(new_n5541), .B(new_n5540), .Y(new_n5542));
  xnor_4 g05166(.A(new_n5541), .B(new_n5540), .Y(new_n5543));
  nand_5 g05167(.A(new_n4898), .B(new_n4895), .Y(new_n5544));
  nand_5 g05168(.A(new_n4899), .B(new_n4894), .Y(new_n5545));
  nand_5 g05169(.A(new_n5545), .B(new_n5544), .Y(new_n5546));
  nor_5  g05170(.A(new_n5546), .B(new_n5543), .Y(new_n5547));
  nor_5  g05171(.A(new_n5547), .B(new_n5542), .Y(new_n5548));
  xor_4  g05172(.A(new_n5548), .B(new_n5539), .Y(new_n5549));
  nand_5 g05173(.A(pi238), .B(pi138), .Y(new_n5550));
  not_8  g05174(.A(new_n4889), .Y(new_n5551));
  nor_5  g05175(.A(new_n4900), .B(new_n5551), .Y(new_n5552));
  xor_4  g05176(.A(new_n5546), .B(new_n5543), .Y(new_n5553));
  nand_5 g05177(.A(new_n5553), .B(new_n5552), .Y(new_n5554));
  xor_4  g05178(.A(new_n5554), .B(new_n5550), .Y(new_n5555));
  xor_4  g05179(.A(new_n5555), .B(new_n5549), .Y(new_n5556));
  nand_5 g05180(.A(pi123), .B(pi061), .Y(new_n5557));
  nand_5 g05181(.A(pi178), .B(pi099), .Y(new_n5558));
  nand_5 g05182(.A(pi188), .B(pi023), .Y(new_n5559));
  nand_5 g05183(.A(new_n5559), .B(new_n5558), .Y(new_n5560));
  nand_5 g05184(.A(pi188), .B(pi099), .Y(new_n5561));
  nand_5 g05185(.A(pi178), .B(pi023), .Y(new_n5562));
  or_6   g05186(.A(new_n5562), .B(new_n5561), .Y(new_n5563));
  nand_5 g05187(.A(new_n5563), .B(new_n5560), .Y(new_n5564));
  xor_4  g05188(.A(new_n5564), .B(new_n5557), .Y(new_n5565));
  nand_5 g05189(.A(pi169), .B(pi061), .Y(new_n5566));
  nand_5 g05190(.A(new_n5566), .B(new_n5561), .Y(new_n5567));
  nand_5 g05191(.A(pi178), .B(pi123), .Y(new_n5568));
  xor_4  g05192(.A(new_n5566), .B(new_n5561), .Y(new_n5569));
  nand_5 g05193(.A(new_n5569), .B(new_n5568), .Y(new_n5570));
  nand_5 g05194(.A(new_n5570), .B(new_n5567), .Y(new_n5571));
  xor_4  g05195(.A(new_n5571), .B(new_n5565), .Y(new_n5572));
  nand_5 g05196(.A(pi169), .B(pi012), .Y(new_n5573));
  nand_5 g05197(.A(pi144), .B(pi071), .Y(new_n5574));
  and_6  g05198(.A(new_n5574), .B(new_n5573), .Y(new_n5575));
  nand_5 g05199(.A(pi071), .B(pi012), .Y(new_n5576));
  nand_5 g05200(.A(pi169), .B(pi144), .Y(new_n5577));
  nor_5  g05201(.A(new_n5577), .B(new_n5576), .Y(new_n5578));
  or_6   g05202(.A(new_n5578), .B(new_n5575), .Y(new_n5579));
  xnor_4 g05203(.A(new_n5579), .B(new_n5572), .Y(new_n5580));
  nand_5 g05204(.A(new_n4846), .B(new_n4845), .Y(new_n5581));
  nand_5 g05205(.A(new_n4847), .B(new_n4844), .Y(new_n5582));
  nand_5 g05206(.A(new_n5582), .B(new_n5581), .Y(new_n5583));
  nand_5 g05207(.A(new_n5583), .B(new_n5576), .Y(new_n5584));
  xor_4  g05208(.A(new_n5569), .B(new_n5568), .Y(new_n5585));
  xor_4  g05209(.A(new_n5583), .B(new_n5576), .Y(new_n5586));
  nand_5 g05210(.A(new_n5586), .B(new_n5585), .Y(new_n5587));
  nand_5 g05211(.A(new_n5587), .B(new_n5584), .Y(new_n5588));
  xor_4  g05212(.A(new_n5588), .B(new_n5580), .Y(new_n5589));
  nand_5 g05213(.A(pi144), .B(pi142), .Y(new_n5590));
  not_8  g05214(.A(new_n5590), .Y(new_n5591));
  or_6   g05215(.A(new_n4842), .B(new_n4841), .Y(new_n5592));
  not_8  g05216(.A(new_n4848), .Y(new_n5593));
  nand_5 g05217(.A(new_n5593), .B(new_n4843), .Y(new_n5594));
  nand_5 g05218(.A(new_n5594), .B(new_n5592), .Y(new_n5595));
  nand_5 g05219(.A(new_n5595), .B(new_n5591), .Y(new_n5596));
  xor_4  g05220(.A(new_n5595), .B(new_n5590), .Y(new_n5597));
  xor_4  g05221(.A(new_n5586), .B(new_n5585), .Y(new_n5598));
  or_6   g05222(.A(new_n5598), .B(new_n5597), .Y(new_n5599));
  nand_5 g05223(.A(new_n5599), .B(new_n5596), .Y(new_n5600));
  xor_4  g05224(.A(new_n5600), .B(new_n5589), .Y(new_n5601));
  nor_5  g05225(.A(new_n4856), .B(new_n4849), .Y(new_n5602));
  xor_4  g05226(.A(new_n5598), .B(new_n5597), .Y(new_n5603));
  nand_5 g05227(.A(new_n5603), .B(new_n5602), .Y(new_n5604));
  nand_5 g05228(.A(pi142), .B(pi098), .Y(new_n5605));
  xor_4  g05229(.A(new_n5605), .B(new_n5604), .Y(new_n5606));
  xor_4  g05230(.A(new_n5606), .B(new_n5601), .Y(new_n5607));
  nor_5  g05231(.A(new_n4833), .B(new_n4826), .Y(new_n5608));
  xor_4  g05232(.A(new_n5494), .B(new_n5369), .Y(new_n5609));
  nand_5 g05233(.A(pi219), .B(pi007), .Y(new_n5610));
  nand_5 g05234(.A(new_n4823), .B(new_n4822), .Y(new_n5611));
  nand_5 g05235(.A(new_n4824), .B(new_n4821), .Y(new_n5612));
  nand_5 g05236(.A(new_n5612), .B(new_n5611), .Y(new_n5613));
  xor_4  g05237(.A(new_n5613), .B(new_n5610), .Y(new_n5614));
  xnor_4 g05238(.A(new_n5614), .B(new_n5609), .Y(new_n5615));
  nand_5 g05239(.A(pi118), .B(pi087), .Y(new_n5616));
  or_6   g05240(.A(new_n4819), .B(new_n4812), .Y(new_n5617));
  nand_5 g05241(.A(new_n4825), .B(new_n4820), .Y(new_n5618));
  nand_5 g05242(.A(new_n5618), .B(new_n5617), .Y(new_n5619));
  xor_4  g05243(.A(new_n5619), .B(new_n5616), .Y(new_n5620));
  xnor_4 g05244(.A(new_n5620), .B(new_n5615), .Y(new_n5621));
  nand_5 g05245(.A(new_n5621), .B(new_n5608), .Y(new_n5622));
  nand_5 g05246(.A(pi113), .B(pi087), .Y(new_n5623));
  xor_4  g05247(.A(new_n5496), .B(new_n5490), .Y(new_n5624));
  nand_5 g05248(.A(pi219), .B(pi118), .Y(new_n5625));
  nand_5 g05249(.A(pi102), .B(pi007), .Y(new_n5626));
  and_6  g05250(.A(new_n5626), .B(new_n5625), .Y(new_n5627));
  nor_5  g05251(.A(new_n5610), .B(new_n5479), .Y(new_n5628));
  or_6   g05252(.A(new_n5628), .B(new_n5627), .Y(new_n5629));
  xnor_4 g05253(.A(new_n5629), .B(new_n5624), .Y(new_n5630));
  nand_5 g05254(.A(new_n5613), .B(new_n5610), .Y(new_n5631));
  nand_5 g05255(.A(new_n5614), .B(new_n5609), .Y(new_n5632));
  nand_5 g05256(.A(new_n5632), .B(new_n5631), .Y(new_n5633));
  xnor_4 g05257(.A(new_n5633), .B(new_n5630), .Y(new_n5634));
  not_8  g05258(.A(new_n5616), .Y(new_n5635));
  nor_5  g05259(.A(new_n5619), .B(new_n5635), .Y(new_n5636));
  nor_5  g05260(.A(new_n5620), .B(new_n5615), .Y(new_n5637));
  nor_5  g05261(.A(new_n5637), .B(new_n5636), .Y(new_n5638));
  xor_4  g05262(.A(new_n5638), .B(new_n5634), .Y(new_n5639));
  xor_4  g05263(.A(new_n5639), .B(new_n5623), .Y(new_n5640));
  not_8  g05264(.A(new_n5640), .Y(new_n5641));
  xor_4  g05265(.A(new_n5641), .B(new_n5622), .Y(new_n5642));
  xor_4  g05266(.A(new_n5642), .B(new_n5607), .Y(new_n5643));
  xor_4  g05267(.A(new_n5621), .B(new_n5608), .Y(new_n5644));
  xor_4  g05268(.A(new_n5603), .B(new_n5602), .Y(new_n5645));
  nor_5  g05269(.A(new_n5645), .B(new_n5644), .Y(new_n5646));
  xnor_4 g05270(.A(new_n5645), .B(new_n5644), .Y(new_n5647));
  nand_5 g05271(.A(new_n4857), .B(new_n4834), .Y(new_n5648));
  nand_5 g05272(.A(new_n4878), .B(new_n4858), .Y(new_n5649));
  nand_5 g05273(.A(new_n5649), .B(new_n5648), .Y(new_n5650));
  nor_5  g05274(.A(new_n5650), .B(new_n5647), .Y(new_n5651));
  nor_5  g05275(.A(new_n5651), .B(new_n5646), .Y(new_n5652));
  xor_4  g05276(.A(new_n5652), .B(new_n5643), .Y(new_n5653));
  xnor_4 g05277(.A(new_n5553), .B(new_n5552), .Y(new_n5654));
  nand_5 g05278(.A(new_n4917), .B(new_n4901), .Y(new_n5655));
  not_8  g05279(.A(new_n4879), .Y(new_n5656));
  nand_5 g05280(.A(new_n4918), .B(new_n5656), .Y(new_n5657));
  nand_5 g05281(.A(new_n5657), .B(new_n5655), .Y(new_n5658));
  or_6   g05282(.A(new_n5658), .B(new_n5654), .Y(new_n5659));
  xnor_4 g05283(.A(new_n5650), .B(new_n5647), .Y(new_n5660));
  xor_4  g05284(.A(new_n5658), .B(new_n5654), .Y(new_n5661));
  nand_5 g05285(.A(new_n5661), .B(new_n5660), .Y(new_n5662));
  nand_5 g05286(.A(new_n5662), .B(new_n5659), .Y(new_n5663));
  xor_4  g05287(.A(new_n5663), .B(new_n5653), .Y(new_n5664));
  xor_4  g05288(.A(new_n5664), .B(new_n5556), .Y(new_n5665));
  nand_5 g05289(.A(new_n5665), .B(new_n5506), .Y(new_n5666));
  xor_4  g05290(.A(new_n5665), .B(new_n5506), .Y(new_n5667));
  xor_4  g05291(.A(new_n5456), .B(new_n5449), .Y(new_n5668));
  or_6   g05292(.A(new_n4957), .B(new_n4939), .Y(new_n5669));
  nand_5 g05293(.A(new_n4958), .B(new_n4919), .Y(new_n5670));
  nand_5 g05294(.A(new_n5670), .B(new_n5669), .Y(new_n5671));
  or_6   g05295(.A(new_n5671), .B(new_n5668), .Y(new_n5672));
  xor_4  g05296(.A(new_n5661), .B(new_n5660), .Y(new_n5673));
  not_8  g05297(.A(new_n5673), .Y(new_n5674));
  xor_4  g05298(.A(new_n5671), .B(new_n5668), .Y(new_n5675));
  nand_5 g05299(.A(new_n5675), .B(new_n5674), .Y(new_n5676));
  nand_5 g05300(.A(new_n5676), .B(new_n5672), .Y(new_n5677));
  nand_5 g05301(.A(new_n5677), .B(new_n5667), .Y(new_n5678));
  nand_5 g05302(.A(new_n5678), .B(new_n5666), .Y(new_n5679));
  nand_5 g05303(.A(new_n5679), .B(new_n5505), .Y(new_n5680));
  not_8  g05304(.A(new_n5638), .Y(new_n5681));
  nor_5  g05305(.A(new_n5681), .B(new_n5634), .Y(new_n5682));
  xor_4  g05306(.A(new_n5501), .B(new_n5500), .Y(new_n5683));
  not_8  g05307(.A(new_n5683), .Y(new_n5684));
  nor_5  g05308(.A(new_n5629), .B(new_n5624), .Y(new_n5685));
  nor_5  g05309(.A(new_n5633), .B(new_n5630), .Y(new_n5686));
  xor_4  g05310(.A(new_n5686), .B(new_n5628), .Y(new_n5687));
  nor_5  g05311(.A(new_n5687), .B(new_n5685), .Y(new_n5688));
  xor_4  g05312(.A(new_n5688), .B(new_n5684), .Y(new_n5689));
  xor_4  g05313(.A(new_n5689), .B(new_n5682), .Y(new_n5690));
  nor_5  g05314(.A(new_n5639), .B(new_n5623), .Y(new_n5691));
  nor_5  g05315(.A(new_n5641), .B(new_n5622), .Y(new_n5692));
  or_6   g05316(.A(new_n5692), .B(new_n5691), .Y(new_n5693));
  xnor_4 g05317(.A(new_n5693), .B(new_n5690), .Y(new_n5694));
  nand_5 g05318(.A(new_n5605), .B(new_n5604), .Y(new_n5695));
  not_8  g05319(.A(new_n5601), .Y(new_n5696));
  nand_5 g05320(.A(new_n5606), .B(new_n5696), .Y(new_n5697));
  nand_5 g05321(.A(new_n5697), .B(new_n5695), .Y(new_n5698));
  nand_5 g05322(.A(new_n5600), .B(new_n5589), .Y(new_n5699));
  nand_5 g05323(.A(pi099), .B(pi061), .Y(new_n5700));
  nand_5 g05324(.A(pi188), .B(pi155), .Y(new_n5701));
  xor_4  g05325(.A(new_n5701), .B(new_n5700), .Y(new_n5702));
  xor_4  g05326(.A(new_n5702), .B(new_n5562), .Y(new_n5703));
  not_8  g05327(.A(new_n5703), .Y(new_n5704));
  nand_5 g05328(.A(pi123), .B(pi012), .Y(new_n5705));
  xor_4  g05329(.A(new_n5705), .B(new_n5563), .Y(new_n5706));
  xor_4  g05330(.A(new_n5706), .B(new_n5704), .Y(new_n5707));
  nand_5 g05331(.A(pi098), .B(pi071), .Y(new_n5708));
  nand_5 g05332(.A(pi142), .B(pi043), .Y(new_n5709));
  xor_4  g05333(.A(new_n5709), .B(new_n5708), .Y(new_n5710));
  xor_4  g05334(.A(new_n5710), .B(new_n5577), .Y(new_n5711));
  nand_5 g05335(.A(new_n5564), .B(new_n5557), .Y(new_n5712));
  nand_5 g05336(.A(new_n5571), .B(new_n5565), .Y(new_n5713));
  nand_5 g05337(.A(new_n5713), .B(new_n5712), .Y(new_n5714));
  xor_4  g05338(.A(new_n5714), .B(new_n5711), .Y(new_n5715));
  xor_4  g05339(.A(new_n5715), .B(new_n5707), .Y(new_n5716));
  nor_5  g05340(.A(new_n5579), .B(new_n5572), .Y(new_n5717));
  nor_5  g05341(.A(new_n5588), .B(new_n5580), .Y(new_n5718));
  xor_4  g05342(.A(new_n5718), .B(new_n5578), .Y(new_n5719));
  nor_5  g05343(.A(new_n5719), .B(new_n5717), .Y(new_n5720));
  xor_4  g05344(.A(new_n5720), .B(new_n5716), .Y(new_n5721));
  xor_4  g05345(.A(new_n5721), .B(new_n5699), .Y(new_n5722));
  xor_4  g05346(.A(new_n5722), .B(new_n5698), .Y(new_n5723));
  xnor_4 g05347(.A(new_n5723), .B(new_n5694), .Y(new_n5724));
  nand_5 g05348(.A(new_n5642), .B(new_n5607), .Y(new_n5725));
  nand_5 g05349(.A(new_n5652), .B(new_n5643), .Y(new_n5726));
  nand_5 g05350(.A(new_n5726), .B(new_n5725), .Y(new_n5727));
  xor_4  g05351(.A(new_n5727), .B(new_n5724), .Y(new_n5728));
  not_8  g05352(.A(new_n5548), .Y(new_n5729));
  nand_5 g05353(.A(new_n5729), .B(new_n5539), .Y(new_n5730));
  nand_5 g05354(.A(pi251), .B(pi162), .Y(new_n5731));
  nand_5 g05355(.A(pi179), .B(pi076), .Y(new_n5732));
  xor_4  g05356(.A(new_n5732), .B(new_n5731), .Y(new_n5733));
  xor_4  g05357(.A(new_n5733), .B(new_n5524), .Y(new_n5734));
  not_8  g05358(.A(new_n5734), .Y(new_n5735));
  nand_5 g05359(.A(pi216), .B(pi048), .Y(new_n5736));
  xor_4  g05360(.A(new_n5736), .B(new_n5525), .Y(new_n5737));
  xor_4  g05361(.A(new_n5737), .B(new_n5735), .Y(new_n5738));
  nand_5 g05362(.A(pi238), .B(pi182), .Y(new_n5739));
  nand_5 g05363(.A(pi193), .B(pi138), .Y(new_n5740));
  xor_4  g05364(.A(new_n5740), .B(new_n5739), .Y(new_n5741));
  xor_4  g05365(.A(new_n5741), .B(new_n5535), .Y(new_n5742));
  nand_5 g05366(.A(new_n5526), .B(new_n5520), .Y(new_n5743));
  nand_5 g05367(.A(new_n5530), .B(new_n5527), .Y(new_n5744));
  nand_5 g05368(.A(new_n5744), .B(new_n5743), .Y(new_n5745));
  xor_4  g05369(.A(new_n5745), .B(new_n5742), .Y(new_n5746));
  xor_4  g05370(.A(new_n5746), .B(new_n5738), .Y(new_n5747));
  nand_5 g05371(.A(new_n5537), .B(new_n5531), .Y(new_n5748));
  nand_5 g05372(.A(new_n5538), .B(new_n5519), .Y(new_n5749));
  nand_5 g05373(.A(new_n5749), .B(new_n5748), .Y(new_n5750));
  xor_4  g05374(.A(new_n5750), .B(new_n5536), .Y(new_n5751));
  xnor_4 g05375(.A(new_n5751), .B(new_n5747), .Y(new_n5752));
  xnor_4 g05376(.A(new_n5752), .B(new_n5730), .Y(new_n5753));
  nand_5 g05377(.A(new_n5554), .B(new_n5550), .Y(new_n5754));
  nand_5 g05378(.A(new_n5555), .B(new_n5549), .Y(new_n5755));
  nand_5 g05379(.A(new_n5755), .B(new_n5754), .Y(new_n5756));
  xor_4  g05380(.A(new_n5756), .B(new_n5753), .Y(new_n5757));
  xor_4  g05381(.A(new_n5757), .B(new_n5728), .Y(new_n5758));
  or_6   g05382(.A(new_n5663), .B(new_n5653), .Y(new_n5759));
  nand_5 g05383(.A(new_n5664), .B(new_n5556), .Y(new_n5760));
  nand_5 g05384(.A(new_n5760), .B(new_n5759), .Y(new_n5761));
  xor_4  g05385(.A(new_n5761), .B(new_n5758), .Y(new_n5762));
  not_8  g05386(.A(new_n5762), .Y(new_n5763));
  xor_4  g05387(.A(new_n5679), .B(new_n5505), .Y(new_n5764));
  nand_5 g05388(.A(new_n5764), .B(new_n5763), .Y(new_n5765));
  nand_5 g05389(.A(new_n5765), .B(new_n5680), .Y(new_n5766));
  xor_4  g05390(.A(new_n5766), .B(new_n5504), .Y(new_n5767));
  xor_4  g05391(.A(new_n5767), .B(new_n5475), .Y(new_n5768));
  xor_4  g05392(.A(new_n5768), .B(new_n5474), .Y(new_n5769));
  xor_4  g05393(.A(new_n5769), .B(new_n5381), .Y(new_n5770));
  xor_4  g05394(.A(new_n5770), .B(new_n5366), .Y(new_n5771));
  nand_5 g05395(.A(new_n5686), .B(new_n5628), .Y(new_n5772));
  or_6   g05396(.A(new_n5688), .B(new_n5684), .Y(new_n5773));
  nand_5 g05397(.A(new_n5773), .B(new_n5772), .Y(new_n5774));
  nand_5 g05398(.A(pi059), .B(pi042), .Y(new_n5775));
  nand_5 g05399(.A(pi135), .B(pi108), .Y(new_n5776));
  xor_4  g05400(.A(new_n5776), .B(new_n5775), .Y(new_n5777));
  xor_4  g05401(.A(new_n5777), .B(new_n5774), .Y(new_n5778));
  nand_5 g05402(.A(new_n5689), .B(new_n5682), .Y(new_n5779));
  nand_5 g05403(.A(new_n5693), .B(new_n5690), .Y(new_n5780));
  nand_5 g05404(.A(new_n5780), .B(new_n5779), .Y(new_n5781));
  nand_5 g05405(.A(pi094), .B(pi051), .Y(new_n5782));
  xor_4  g05406(.A(new_n5782), .B(new_n5781), .Y(new_n5783));
  xor_4  g05407(.A(new_n5783), .B(new_n5778), .Y(new_n5784));
  nand_5 g05408(.A(pi122), .B(pi007), .Y(new_n5785));
  nand_5 g05409(.A(pi118), .B(pi001), .Y(new_n5786));
  xor_4  g05410(.A(new_n5786), .B(new_n5785), .Y(new_n5787));
  nand_5 g05411(.A(new_n5714), .B(new_n5711), .Y(new_n5788));
  not_8  g05412(.A(new_n5707), .Y(new_n5789));
  nand_5 g05413(.A(new_n5715), .B(new_n5789), .Y(new_n5790));
  nand_5 g05414(.A(new_n5790), .B(new_n5788), .Y(new_n5791));
  nand_5 g05415(.A(pi144), .B(pi123), .Y(new_n5792));
  nand_5 g05416(.A(pi071), .B(pi043), .Y(new_n5793));
  nand_5 g05417(.A(pi169), .B(pi098), .Y(new_n5794));
  xnor_4 g05418(.A(new_n5794), .B(new_n5793), .Y(new_n5795));
  xor_4  g05419(.A(new_n5795), .B(new_n5792), .Y(new_n5796));
  xor_4  g05420(.A(new_n5796), .B(new_n5791), .Y(new_n5797));
  nand_5 g05421(.A(new_n5709), .B(new_n5708), .Y(new_n5798));
  nand_5 g05422(.A(new_n5710), .B(new_n5577), .Y(new_n5799));
  nand_5 g05423(.A(new_n5799), .B(new_n5798), .Y(new_n5800));
  or_6   g05424(.A(new_n5705), .B(new_n5563), .Y(new_n5801));
  nand_5 g05425(.A(new_n5706), .B(new_n5704), .Y(new_n5802));
  nand_5 g05426(.A(new_n5802), .B(new_n5801), .Y(new_n5803));
  xor_4  g05427(.A(new_n5803), .B(new_n5800), .Y(new_n5804));
  nand_5 g05428(.A(new_n5701), .B(new_n5700), .Y(new_n5805));
  nand_5 g05429(.A(new_n5702), .B(new_n5562), .Y(new_n5806));
  nand_5 g05430(.A(new_n5806), .B(new_n5805), .Y(new_n5807));
  nand_5 g05431(.A(pi099), .B(pi012), .Y(new_n5808));
  xor_4  g05432(.A(new_n5808), .B(new_n5807), .Y(new_n5809));
  xor_4  g05433(.A(new_n5809), .B(new_n5804), .Y(new_n5810));
  xor_4  g05434(.A(new_n5810), .B(new_n5797), .Y(new_n5811));
  xor_4  g05435(.A(new_n5811), .B(new_n5787), .Y(new_n5812));
  xor_4  g05436(.A(new_n5812), .B(new_n5784), .Y(new_n5813));
  xor_4  g05437(.A(new_n5813), .B(new_n5771), .Y(new_n5814));
  nand_5 g05438(.A(new_n5740), .B(new_n5739), .Y(new_n5815));
  nand_5 g05439(.A(new_n5741), .B(new_n5535), .Y(new_n5816));
  nand_5 g05440(.A(new_n5816), .B(new_n5815), .Y(new_n5817));
  nand_5 g05441(.A(pi237), .B(pi216), .Y(new_n5818));
  nand_5 g05442(.A(pi238), .B(pi041), .Y(new_n5819));
  xor_4  g05443(.A(new_n5819), .B(new_n5818), .Y(new_n5820));
  xor_4  g05444(.A(new_n5820), .B(new_n5817), .Y(new_n5821));
  xor_4  g05445(.A(new_n5821), .B(new_n5814), .Y(new_n5822));
  nand_5 g05446(.A(new_n5721), .B(new_n5699), .Y(new_n5823));
  nand_5 g05447(.A(new_n5722), .B(new_n5698), .Y(new_n5824));
  nand_5 g05448(.A(new_n5824), .B(new_n5823), .Y(new_n5825));
  nand_5 g05449(.A(new_n5718), .B(new_n5578), .Y(new_n5826));
  not_8  g05450(.A(new_n5720), .Y(new_n5827));
  nand_5 g05451(.A(new_n5827), .B(new_n5716), .Y(new_n5828));
  nand_5 g05452(.A(new_n5828), .B(new_n5826), .Y(new_n5829));
  xor_4  g05453(.A(new_n5829), .B(new_n5825), .Y(new_n5830));
  or_6   g05454(.A(new_n5736), .B(new_n5525), .Y(new_n5831));
  nand_5 g05455(.A(new_n5737), .B(new_n5735), .Y(new_n5832));
  nand_5 g05456(.A(new_n5832), .B(new_n5831), .Y(new_n5833));
  nand_5 g05457(.A(new_n5745), .B(new_n5742), .Y(new_n5834));
  not_8  g05458(.A(new_n5738), .Y(new_n5835));
  nand_5 g05459(.A(new_n5746), .B(new_n5835), .Y(new_n5836));
  nand_5 g05460(.A(new_n5836), .B(new_n5834), .Y(new_n5837));
  xor_4  g05461(.A(new_n5837), .B(new_n5833), .Y(new_n5838));
  xor_4  g05462(.A(new_n5838), .B(new_n5830), .Y(new_n5839));
  not_8  g05463(.A(new_n5757), .Y(new_n5840));
  nor_5  g05464(.A(new_n5840), .B(new_n5728), .Y(new_n5841));
  nor_5  g05465(.A(new_n5761), .B(new_n5758), .Y(new_n5842));
  nor_5  g05466(.A(new_n5842), .B(new_n5841), .Y(new_n5843));
  nor_5  g05467(.A(new_n5420), .B(new_n5391), .Y(new_n5844));
  nor_5  g05468(.A(new_n5422), .B(new_n5419), .Y(new_n5845));
  or_6   g05469(.A(new_n5845), .B(new_n5844), .Y(new_n5846));
  nand_5 g05470(.A(pi177), .B(pi057), .Y(new_n5847));
  nand_5 g05471(.A(pi225), .B(pi194), .Y(new_n5848));
  xor_4  g05472(.A(new_n5848), .B(new_n5847), .Y(new_n5849));
  xor_4  g05473(.A(new_n5849), .B(new_n5846), .Y(new_n5850));
  xor_4  g05474(.A(new_n5850), .B(new_n5843), .Y(new_n5851));
  nand_5 g05475(.A(new_n5425), .B(new_n5424), .Y(new_n5852));
  nand_5 g05476(.A(new_n5426), .B(new_n5382), .Y(new_n5853));
  nand_5 g05477(.A(new_n5853), .B(new_n5852), .Y(new_n5854));
  or_6   g05478(.A(new_n5430), .B(new_n5427), .Y(new_n5855));
  nand_5 g05479(.A(new_n5431), .B(new_n5423), .Y(new_n5856));
  nand_5 g05480(.A(new_n5856), .B(new_n5855), .Y(new_n5857));
  xor_4  g05481(.A(new_n5857), .B(new_n5854), .Y(new_n5858));
  nand_5 g05482(.A(pi068), .B(pi020), .Y(new_n5859));
  nand_5 g05483(.A(pi101), .B(pi085), .Y(new_n5860));
  xor_4  g05484(.A(new_n5860), .B(new_n5859), .Y(new_n5861));
  xor_4  g05485(.A(new_n5861), .B(new_n5858), .Y(new_n5862));
  nor_5  g05486(.A(new_n5752), .B(new_n5730), .Y(new_n5863));
  nor_5  g05487(.A(new_n5756), .B(new_n5753), .Y(new_n5864));
  nor_5  g05488(.A(new_n5864), .B(new_n5863), .Y(new_n5865));
  nand_5 g05489(.A(new_n5417), .B(new_n5416), .Y(new_n5866));
  nand_5 g05490(.A(new_n5418), .B(new_n5390), .Y(new_n5867));
  nand_5 g05491(.A(new_n5867), .B(new_n5866), .Y(new_n5868));
  nand_5 g05492(.A(pi223), .B(pi180), .Y(new_n5869));
  xor_4  g05493(.A(new_n5869), .B(new_n5868), .Y(new_n5870));
  xor_4  g05494(.A(new_n5870), .B(new_n5865), .Y(new_n5871));
  xor_4  g05495(.A(new_n5871), .B(new_n5862), .Y(new_n5872));
  nand_5 g05496(.A(pi060), .B(pi036), .Y(new_n5873));
  nand_5 g05497(.A(pi159), .B(pi138), .Y(new_n5874));
  nand_5 g05498(.A(pi251), .B(pi033), .Y(new_n5875));
  nand_5 g05499(.A(pi192), .B(pi162), .Y(new_n5876));
  or_6   g05500(.A(new_n5750), .B(new_n5536), .Y(new_n5877));
  nand_5 g05501(.A(new_n5751), .B(new_n5747), .Y(new_n5878));
  nand_5 g05502(.A(new_n5878), .B(new_n5877), .Y(new_n5879));
  xor_4  g05503(.A(new_n5879), .B(new_n5876), .Y(new_n5880));
  xor_4  g05504(.A(new_n5880), .B(new_n5875), .Y(new_n5881));
  xor_4  g05505(.A(new_n5881), .B(new_n5874), .Y(new_n5882));
  xor_4  g05506(.A(new_n5882), .B(new_n5873), .Y(new_n5883));
  xor_4  g05507(.A(new_n5883), .B(new_n5872), .Y(new_n5884));
  xor_4  g05508(.A(new_n5884), .B(new_n5851), .Y(new_n5885));
  nand_5 g05509(.A(pi076), .B(pi048), .Y(new_n5886));
  nand_5 g05510(.A(pi193), .B(pi182), .Y(new_n5887));
  nand_5 g05511(.A(new_n5732), .B(new_n5731), .Y(new_n5888));
  nand_5 g05512(.A(new_n5733), .B(new_n5524), .Y(new_n5889));
  nand_5 g05513(.A(new_n5889), .B(new_n5888), .Y(new_n5890));
  xor_4  g05514(.A(new_n5890), .B(new_n5887), .Y(new_n5891));
  xor_4  g05515(.A(new_n5891), .B(new_n5886), .Y(new_n5892));
  xor_4  g05516(.A(new_n5892), .B(new_n5885), .Y(new_n5893));
  xor_4  g05517(.A(new_n5893), .B(new_n5839), .Y(new_n5894));
  nand_5 g05518(.A(pi179), .B(pi079), .Y(new_n5895));
  nand_5 g05519(.A(pi188), .B(pi086), .Y(new_n5896));
  nand_5 g05520(.A(pi061), .B(pi023), .Y(new_n5897));
  nand_5 g05521(.A(pi178), .B(pi155), .Y(new_n5898));
  xor_4  g05522(.A(new_n5898), .B(new_n5897), .Y(new_n5899));
  nand_5 g05523(.A(pi142), .B(pi126), .Y(new_n5900));
  nand_5 g05524(.A(new_n5723), .B(new_n5694), .Y(new_n5901));
  or_6   g05525(.A(new_n5727), .B(new_n5724), .Y(new_n5902));
  nand_5 g05526(.A(new_n5902), .B(new_n5901), .Y(new_n5903));
  xor_4  g05527(.A(new_n5903), .B(new_n5900), .Y(new_n5904));
  xor_4  g05528(.A(new_n5904), .B(new_n5899), .Y(new_n5905));
  xor_4  g05529(.A(new_n5905), .B(new_n5896), .Y(new_n5906));
  xor_4  g05530(.A(new_n5906), .B(new_n5895), .Y(new_n5907));
  xor_4  g05531(.A(new_n5907), .B(new_n5894), .Y(new_n5908));
  xor_4  g05532(.A(new_n5908), .B(new_n5822), .Y(po021));
  xor_4  g05533(.A(new_n4806), .B(new_n4799), .Y(po022));
  xor_4  g05534(.A(new_n2575), .B(new_n2539), .Y(po023));
  xor_4  g05535(.A(new_n1815), .B(new_n1813), .Y(po024));
  xnor_4 g05536(.A(new_n3692), .B(new_n3691), .Y(po025));
  xor_4  g05537(.A(new_n5361), .B(new_n5360), .Y(po026));
  nand_5 g05538(.A(pi141), .B(pi089), .Y(new_n5915));
  nand_5 g05539(.A(new_n3335), .B(new_n3334), .Y(new_n5916));
  nand_5 g05540(.A(new_n3336), .B(new_n3333), .Y(new_n5917));
  nand_5 g05541(.A(new_n5917), .B(new_n5916), .Y(new_n5918));
  xor_4  g05542(.A(new_n5918), .B(new_n5915), .Y(new_n5919));
  nand_5 g05543(.A(pi254), .B(pi047), .Y(new_n5920));
  nand_5 g05544(.A(pi158), .B(pi090), .Y(new_n5921));
  nand_5 g05545(.A(new_n5921), .B(new_n5920), .Y(new_n5922));
  nand_5 g05546(.A(pi158), .B(pi047), .Y(new_n5923));
  nor_5  g05547(.A(new_n5923), .B(new_n3335), .Y(new_n5924));
  not_8  g05548(.A(new_n5924), .Y(new_n5925));
  nand_5 g05549(.A(new_n5925), .B(new_n5922), .Y(new_n5926));
  xor_4  g05550(.A(new_n5926), .B(new_n5919), .Y(new_n5927));
  nand_5 g05551(.A(new_n3341), .B(new_n3338), .Y(new_n5928));
  nand_5 g05552(.A(new_n3342), .B(new_n3337), .Y(new_n5929));
  nand_5 g05553(.A(new_n5929), .B(new_n5928), .Y(new_n5930));
  nand_5 g05554(.A(pi161), .B(pi154), .Y(new_n5931));
  nand_5 g05555(.A(pi241), .B(pi095), .Y(new_n5932));
  nand_5 g05556(.A(new_n5932), .B(new_n5931), .Y(new_n5933));
  nand_5 g05557(.A(pi161), .B(pi095), .Y(new_n5934));
  or_6   g05558(.A(new_n5934), .B(new_n3338), .Y(new_n5935));
  nand_5 g05559(.A(new_n5935), .B(new_n5933), .Y(new_n5936));
  xor_4  g05560(.A(new_n5936), .B(new_n5930), .Y(new_n5937));
  xor_4  g05561(.A(new_n5937), .B(new_n5927), .Y(new_n5938));
  not_8  g05562(.A(new_n5938), .Y(new_n5939));
  not_8  g05563(.A(new_n3344), .Y(new_n5940));
  nand_5 g05564(.A(new_n3347), .B(new_n5940), .Y(new_n5941));
  or_6   g05565(.A(new_n3348), .B(new_n3343), .Y(new_n5942));
  nand_5 g05566(.A(new_n5942), .B(new_n5941), .Y(new_n5943));
  nand_5 g05567(.A(new_n5943), .B(new_n5939), .Y(new_n5944));
  nand_5 g05568(.A(pi090), .B(pi089), .Y(new_n5945));
  nand_5 g05569(.A(pi254), .B(pi018), .Y(new_n5946));
  xor_4  g05570(.A(new_n5946), .B(new_n5945), .Y(new_n5947));
  xor_4  g05571(.A(new_n5947), .B(new_n5923), .Y(new_n5948));
  nand_5 g05572(.A(pi154), .B(pi141), .Y(new_n5949));
  xor_4  g05573(.A(new_n5949), .B(new_n5925), .Y(new_n5950));
  not_8  g05574(.A(new_n5950), .Y(new_n5951));
  xor_4  g05575(.A(new_n5951), .B(new_n5948), .Y(new_n5952));
  nand_5 g05576(.A(pi241), .B(pi006), .Y(new_n5953));
  nand_5 g05577(.A(pi236), .B(pi209), .Y(new_n5954));
  xor_4  g05578(.A(new_n5954), .B(new_n5953), .Y(new_n5955));
  xor_4  g05579(.A(new_n5955), .B(new_n5934), .Y(new_n5956));
  nand_5 g05580(.A(new_n5918), .B(new_n5915), .Y(new_n5957));
  nand_5 g05581(.A(new_n5926), .B(new_n5919), .Y(new_n5958));
  nand_5 g05582(.A(new_n5958), .B(new_n5957), .Y(new_n5959));
  xor_4  g05583(.A(new_n5959), .B(new_n5956), .Y(new_n5960));
  xor_4  g05584(.A(new_n5960), .B(new_n5952), .Y(new_n5961));
  nand_5 g05585(.A(new_n5936), .B(new_n5930), .Y(new_n5962));
  nand_5 g05586(.A(new_n5937), .B(new_n5927), .Y(new_n5963));
  nand_5 g05587(.A(new_n5963), .B(new_n5962), .Y(new_n5964));
  xor_4  g05588(.A(new_n5964), .B(new_n5935), .Y(new_n5965));
  xnor_4 g05589(.A(new_n5965), .B(new_n5961), .Y(new_n5966));
  or_6   g05590(.A(new_n5966), .B(new_n5944), .Y(new_n5967));
  xor_4  g05591(.A(new_n5966), .B(new_n5944), .Y(new_n5968));
  nand_5 g05592(.A(pi236), .B(pi006), .Y(new_n5969));
  xor_4  g05593(.A(new_n5943), .B(new_n5938), .Y(new_n5970));
  nor_5  g05594(.A(new_n5970), .B(new_n5969), .Y(new_n5971));
  nand_5 g05595(.A(new_n3349), .B(new_n3332), .Y(new_n5972));
  xor_4  g05596(.A(new_n5970), .B(new_n5969), .Y(new_n5973));
  not_8  g05597(.A(new_n5973), .Y(new_n5974));
  nor_5  g05598(.A(new_n5974), .B(new_n5972), .Y(new_n5975));
  or_6   g05599(.A(new_n5975), .B(new_n5971), .Y(new_n5976));
  nand_5 g05600(.A(new_n5976), .B(new_n5968), .Y(new_n5977));
  nand_5 g05601(.A(new_n5977), .B(new_n5967), .Y(new_n5978));
  nand_5 g05602(.A(pi229), .B(pi133), .Y(new_n5979));
  nand_5 g05603(.A(new_n3470), .B(new_n3469), .Y(new_n5980));
  nand_5 g05604(.A(new_n3471), .B(new_n3468), .Y(new_n5981));
  nand_5 g05605(.A(new_n5981), .B(new_n5980), .Y(new_n5982));
  xor_4  g05606(.A(new_n5982), .B(new_n5979), .Y(new_n5983));
  nand_5 g05607(.A(pi189), .B(pi092), .Y(new_n5984));
  nand_5 g05608(.A(pi190), .B(pi064), .Y(new_n5985));
  nand_5 g05609(.A(new_n5985), .B(new_n5984), .Y(new_n5986));
  nand_5 g05610(.A(pi092), .B(pi064), .Y(new_n5987));
  or_6   g05611(.A(new_n5987), .B(new_n3470), .Y(new_n5988));
  nand_5 g05612(.A(new_n5988), .B(new_n5986), .Y(new_n5989));
  xor_4  g05613(.A(new_n5989), .B(new_n5983), .Y(new_n5990));
  nand_5 g05614(.A(pi077), .B(pi067), .Y(new_n5991));
  nand_5 g05615(.A(pi053), .B(pi052), .Y(new_n5992));
  and_6  g05616(.A(new_n5992), .B(new_n5991), .Y(new_n5993));
  nand_5 g05617(.A(pi077), .B(pi053), .Y(new_n5994));
  nor_5  g05618(.A(new_n5994), .B(new_n3473), .Y(new_n5995));
  or_6   g05619(.A(new_n5995), .B(new_n5993), .Y(new_n5996));
  xnor_4 g05620(.A(new_n5996), .B(new_n5990), .Y(new_n5997));
  nand_5 g05621(.A(new_n3476), .B(new_n3473), .Y(new_n5998));
  nand_5 g05622(.A(new_n3477), .B(new_n3472), .Y(new_n5999));
  nand_5 g05623(.A(new_n5999), .B(new_n5998), .Y(new_n6000));
  xor_4  g05624(.A(new_n6000), .B(new_n5997), .Y(new_n6001));
  not_8  g05625(.A(new_n3479), .Y(new_n6002));
  nand_5 g05626(.A(new_n3482), .B(new_n6002), .Y(new_n6003));
  or_6   g05627(.A(new_n3483), .B(new_n3478), .Y(new_n6004));
  nand_5 g05628(.A(new_n6004), .B(new_n6003), .Y(new_n6005));
  nand_5 g05629(.A(new_n6005), .B(new_n6001), .Y(new_n6006));
  nand_5 g05630(.A(pi229), .B(pi189), .Y(new_n6007));
  nand_5 g05631(.A(pi190), .B(pi084), .Y(new_n6008));
  xor_4  g05632(.A(new_n6008), .B(new_n6007), .Y(new_n6009));
  xor_4  g05633(.A(new_n6009), .B(new_n5987), .Y(new_n6010));
  nand_5 g05634(.A(pi133), .B(pi067), .Y(new_n6011));
  xor_4  g05635(.A(new_n6011), .B(new_n5988), .Y(new_n6012));
  xor_4  g05636(.A(new_n6012), .B(new_n6010), .Y(new_n6013));
  nand_5 g05637(.A(pi185), .B(pi052), .Y(new_n6014));
  nand_5 g05638(.A(pi131), .B(pi030), .Y(new_n6015));
  xor_4  g05639(.A(new_n6015), .B(new_n5994), .Y(new_n6016));
  xor_4  g05640(.A(new_n6016), .B(new_n6014), .Y(new_n6017));
  nand_5 g05641(.A(new_n5982), .B(new_n5979), .Y(new_n6018));
  nand_5 g05642(.A(new_n5989), .B(new_n5983), .Y(new_n6019));
  nand_5 g05643(.A(new_n6019), .B(new_n6018), .Y(new_n6020));
  xor_4  g05644(.A(new_n6020), .B(new_n6017), .Y(new_n6021));
  xnor_4 g05645(.A(new_n6021), .B(new_n6013), .Y(new_n6022));
  nor_5  g05646(.A(new_n5996), .B(new_n5990), .Y(new_n6023));
  nor_5  g05647(.A(new_n6000), .B(new_n5997), .Y(new_n6024));
  xor_4  g05648(.A(new_n6024), .B(new_n5995), .Y(new_n6025));
  nor_5  g05649(.A(new_n6025), .B(new_n6023), .Y(new_n6026));
  xor_4  g05650(.A(new_n6026), .B(new_n6022), .Y(new_n6027));
  xnor_4 g05651(.A(new_n6027), .B(new_n6006), .Y(new_n6028));
  nand_5 g05652(.A(new_n3484), .B(new_n3467), .Y(new_n6029));
  nand_5 g05653(.A(pi185), .B(pi131), .Y(new_n6030));
  nand_5 g05654(.A(new_n6030), .B(new_n6029), .Y(new_n6031));
  xnor_4 g05655(.A(new_n6005), .B(new_n6001), .Y(new_n6032));
  xor_4  g05656(.A(new_n6030), .B(new_n6029), .Y(new_n6033));
  nand_5 g05657(.A(new_n6033), .B(new_n6032), .Y(new_n6034));
  nand_5 g05658(.A(new_n6034), .B(new_n6031), .Y(new_n6035));
  xor_4  g05659(.A(new_n6035), .B(new_n6028), .Y(new_n6036));
  nand_5 g05660(.A(pi073), .B(pi013), .Y(new_n6037));
  nand_5 g05661(.A(pi112), .B(pi004), .Y(new_n6038));
  nand_5 g05662(.A(pi170), .B(pi105), .Y(new_n6039));
  nand_5 g05663(.A(new_n6039), .B(new_n6038), .Y(new_n6040));
  nand_5 g05664(.A(pi105), .B(pi004), .Y(new_n6041));
  or_6   g05665(.A(new_n6041), .B(new_n3295), .Y(new_n6042));
  nand_5 g05666(.A(new_n6042), .B(new_n6040), .Y(new_n6043));
  xor_4  g05667(.A(new_n6043), .B(new_n6037), .Y(new_n6044));
  nand_5 g05668(.A(new_n3296), .B(new_n3295), .Y(new_n6045));
  nand_5 g05669(.A(new_n3297), .B(new_n3294), .Y(new_n6046));
  nand_5 g05670(.A(new_n6046), .B(new_n6045), .Y(new_n6047));
  xor_4  g05671(.A(new_n6047), .B(new_n6044), .Y(new_n6048));
  nand_5 g05672(.A(pi212), .B(pi130), .Y(new_n6049));
  nand_5 g05673(.A(pi104), .B(pi003), .Y(new_n6050));
  nand_5 g05674(.A(new_n6050), .B(new_n6049), .Y(new_n6051));
  nand_5 g05675(.A(pi130), .B(pi104), .Y(new_n6052));
  nor_5  g05676(.A(new_n6052), .B(new_n3299), .Y(new_n6053));
  not_8  g05677(.A(new_n6053), .Y(new_n6054));
  nand_5 g05678(.A(new_n6054), .B(new_n6051), .Y(new_n6055));
  xnor_4 g05679(.A(new_n6055), .B(new_n6048), .Y(new_n6056));
  nand_5 g05680(.A(new_n3302), .B(new_n3299), .Y(new_n6057));
  nand_5 g05681(.A(new_n3303), .B(new_n3298), .Y(new_n6058));
  nand_5 g05682(.A(new_n6058), .B(new_n6057), .Y(new_n6059));
  xnor_4 g05683(.A(new_n6059), .B(new_n6056), .Y(new_n6060));
  not_8  g05684(.A(new_n3305), .Y(new_n6061));
  nor_5  g05685(.A(new_n3309), .B(new_n6061), .Y(new_n6062));
  nor_5  g05686(.A(new_n3310), .B(new_n3304), .Y(new_n6063));
  nor_5  g05687(.A(new_n6063), .B(new_n6062), .Y(new_n6064));
  not_8  g05688(.A(new_n6064), .Y(new_n6065));
  nor_5  g05689(.A(new_n6065), .B(new_n6060), .Y(new_n6066));
  not_8  g05690(.A(new_n6066), .Y(new_n6067));
  nand_5 g05691(.A(pi183), .B(pi170), .Y(new_n6068));
  nand_5 g05692(.A(pi112), .B(pi073), .Y(new_n6069));
  xor_4  g05693(.A(new_n6069), .B(new_n6068), .Y(new_n6070));
  xor_4  g05694(.A(new_n6070), .B(new_n6041), .Y(new_n6071));
  nand_5 g05695(.A(pi013), .B(pi003), .Y(new_n6072));
  xor_4  g05696(.A(new_n6072), .B(new_n6042), .Y(new_n6073));
  xor_4  g05697(.A(new_n6073), .B(new_n6071), .Y(new_n6074));
  nand_5 g05698(.A(pi215), .B(pi213), .Y(new_n6075));
  nand_5 g05699(.A(pi212), .B(pi124), .Y(new_n6076));
  xor_4  g05700(.A(new_n6076), .B(new_n6052), .Y(new_n6077));
  xor_4  g05701(.A(new_n6077), .B(new_n6075), .Y(new_n6078));
  nand_5 g05702(.A(new_n6043), .B(new_n6037), .Y(new_n6079));
  nand_5 g05703(.A(new_n6047), .B(new_n6044), .Y(new_n6080));
  nand_5 g05704(.A(new_n6080), .B(new_n6079), .Y(new_n6081));
  xor_4  g05705(.A(new_n6081), .B(new_n6078), .Y(new_n6082));
  xnor_4 g05706(.A(new_n6082), .B(new_n6074), .Y(new_n6083));
  nor_5  g05707(.A(new_n6059), .B(new_n6056), .Y(new_n6084));
  and_6  g05708(.A(new_n6084), .B(new_n6053), .Y(new_n6085));
  or_6   g05709(.A(new_n6055), .B(new_n6048), .Y(new_n6086));
  nand_5 g05710(.A(new_n6086), .B(new_n6054), .Y(new_n6087));
  nor_5  g05711(.A(new_n6087), .B(new_n6084), .Y(new_n6088));
  or_6   g05712(.A(new_n6088), .B(new_n6085), .Y(new_n6089));
  xor_4  g05713(.A(new_n6089), .B(new_n6083), .Y(new_n6090));
  xor_4  g05714(.A(new_n6090), .B(new_n6067), .Y(new_n6091));
  nand_5 g05715(.A(pi213), .B(pi124), .Y(new_n6092));
  xor_4  g05716(.A(new_n6064), .B(new_n6060), .Y(new_n6093));
  or_6   g05717(.A(new_n6093), .B(new_n6092), .Y(new_n6094));
  not_8  g05718(.A(new_n3311), .Y(new_n6095));
  nand_5 g05719(.A(new_n6095), .B(new_n3293), .Y(new_n6096));
  not_8  g05720(.A(new_n6096), .Y(new_n6097));
  xor_4  g05721(.A(new_n6093), .B(new_n6092), .Y(new_n6098));
  nand_5 g05722(.A(new_n6098), .B(new_n6097), .Y(new_n6099));
  nand_5 g05723(.A(new_n6099), .B(new_n6094), .Y(new_n6100));
  xor_4  g05724(.A(new_n6100), .B(new_n6091), .Y(new_n6101));
  xor_4  g05725(.A(new_n5974), .B(new_n5972), .Y(new_n6102));
  xor_4  g05726(.A(new_n6098), .B(new_n6097), .Y(new_n6103));
  nand_5 g05727(.A(new_n6103), .B(new_n6102), .Y(new_n6104));
  not_8  g05728(.A(new_n6104), .Y(new_n6105));
  xnor_4 g05729(.A(new_n6103), .B(new_n6102), .Y(new_n6106));
  or_6   g05730(.A(new_n3377), .B(new_n3350), .Y(new_n6107));
  nand_5 g05731(.A(new_n3378), .B(new_n3312), .Y(new_n6108));
  nand_5 g05732(.A(new_n6108), .B(new_n6107), .Y(new_n6109));
  nor_5  g05733(.A(new_n6109), .B(new_n6106), .Y(new_n6110));
  nor_5  g05734(.A(new_n6110), .B(new_n6105), .Y(new_n6111));
  not_8  g05735(.A(new_n6111), .Y(new_n6112));
  xor_4  g05736(.A(new_n6112), .B(new_n6101), .Y(new_n6113));
  xor_4  g05737(.A(new_n5976), .B(new_n5968), .Y(new_n6114));
  xnor_4 g05738(.A(new_n6114), .B(new_n6113), .Y(new_n6115));
  nand_5 g05739(.A(new_n3410), .B(new_n3407), .Y(new_n6116));
  nand_5 g05740(.A(new_n3411), .B(new_n3406), .Y(new_n6117));
  nand_5 g05741(.A(new_n6117), .B(new_n6116), .Y(new_n6118));
  nand_5 g05742(.A(pi120), .B(pi035), .Y(new_n6119));
  nand_5 g05743(.A(new_n3404), .B(new_n3403), .Y(new_n6120));
  nand_5 g05744(.A(new_n3405), .B(new_n3402), .Y(new_n6121));
  nand_5 g05745(.A(new_n6121), .B(new_n6120), .Y(new_n6122));
  xor_4  g05746(.A(new_n6122), .B(new_n6119), .Y(new_n6123));
  nand_5 g05747(.A(pi062), .B(pi015), .Y(new_n6124));
  nand_5 g05748(.A(pi204), .B(pi065), .Y(new_n6125));
  nand_5 g05749(.A(new_n6125), .B(new_n6124), .Y(new_n6126));
  nand_5 g05750(.A(pi204), .B(pi062), .Y(new_n6127));
  nor_5  g05751(.A(new_n6127), .B(new_n3404), .Y(new_n6128));
  not_8  g05752(.A(new_n6128), .Y(new_n6129));
  nand_5 g05753(.A(new_n6129), .B(new_n6126), .Y(new_n6130));
  xor_4  g05754(.A(new_n6130), .B(new_n6123), .Y(new_n6131));
  nand_5 g05755(.A(pi172), .B(pi139), .Y(new_n6132));
  nand_5 g05756(.A(pi208), .B(pi198), .Y(new_n6133));
  nand_5 g05757(.A(new_n6133), .B(new_n6132), .Y(new_n6134));
  nand_5 g05758(.A(pi198), .B(pi139), .Y(new_n6135));
  or_6   g05759(.A(new_n6135), .B(new_n3407), .Y(new_n6136));
  nand_5 g05760(.A(new_n6136), .B(new_n6134), .Y(new_n6137));
  xor_4  g05761(.A(new_n6137), .B(new_n6131), .Y(new_n6138));
  xor_4  g05762(.A(new_n6138), .B(new_n6118), .Y(new_n6139));
  not_8  g05763(.A(new_n6139), .Y(new_n6140));
  not_8  g05764(.A(new_n3413), .Y(new_n6141));
  nand_5 g05765(.A(new_n3416), .B(new_n6141), .Y(new_n6142));
  or_6   g05766(.A(new_n3417), .B(new_n3412), .Y(new_n6143));
  nand_5 g05767(.A(new_n6143), .B(new_n6142), .Y(new_n6144));
  nand_5 g05768(.A(new_n6144), .B(new_n6140), .Y(new_n6145));
  nand_5 g05769(.A(pi120), .B(pi015), .Y(new_n6146));
  nand_5 g05770(.A(pi146), .B(pi065), .Y(new_n6147));
  xor_4  g05771(.A(new_n6147), .B(new_n6146), .Y(new_n6148));
  xor_4  g05772(.A(new_n6148), .B(new_n6127), .Y(new_n6149));
  nand_5 g05773(.A(pi172), .B(pi035), .Y(new_n6150));
  xor_4  g05774(.A(new_n6150), .B(new_n6129), .Y(new_n6151));
  not_8  g05775(.A(new_n6151), .Y(new_n6152));
  xor_4  g05776(.A(new_n6152), .B(new_n6149), .Y(new_n6153));
  nand_5 g05777(.A(pi197), .B(pi168), .Y(new_n6154));
  nand_5 g05778(.A(pi208), .B(pi165), .Y(new_n6155));
  xor_4  g05779(.A(new_n6155), .B(new_n6154), .Y(new_n6156));
  xor_4  g05780(.A(new_n6156), .B(new_n6135), .Y(new_n6157));
  nand_5 g05781(.A(new_n6122), .B(new_n6119), .Y(new_n6158));
  nand_5 g05782(.A(new_n6130), .B(new_n6123), .Y(new_n6159));
  nand_5 g05783(.A(new_n6159), .B(new_n6158), .Y(new_n6160));
  xor_4  g05784(.A(new_n6160), .B(new_n6157), .Y(new_n6161));
  xor_4  g05785(.A(new_n6161), .B(new_n6153), .Y(new_n6162));
  nand_5 g05786(.A(new_n6137), .B(new_n6131), .Y(new_n6163));
  nand_5 g05787(.A(new_n6138), .B(new_n6118), .Y(new_n6164));
  nand_5 g05788(.A(new_n6164), .B(new_n6163), .Y(new_n6165));
  xor_4  g05789(.A(new_n6165), .B(new_n6136), .Y(new_n6166));
  xnor_4 g05790(.A(new_n6166), .B(new_n6162), .Y(new_n6167));
  xor_4  g05791(.A(new_n6167), .B(new_n6145), .Y(new_n6168));
  nand_5 g05792(.A(pi168), .B(pi165), .Y(new_n6169));
  xor_4  g05793(.A(new_n6144), .B(new_n6139), .Y(new_n6170));
  nor_5  g05794(.A(new_n6170), .B(new_n6169), .Y(new_n6171));
  nand_5 g05795(.A(new_n3418), .B(new_n3401), .Y(new_n6172));
  xor_4  g05796(.A(new_n6170), .B(new_n6169), .Y(new_n6173));
  not_8  g05797(.A(new_n6173), .Y(new_n6174));
  nor_5  g05798(.A(new_n6174), .B(new_n6172), .Y(new_n6175));
  or_6   g05799(.A(new_n6175), .B(new_n6171), .Y(new_n6176));
  xor_4  g05800(.A(new_n6176), .B(new_n6168), .Y(new_n6177));
  xor_4  g05801(.A(new_n6177), .B(new_n6115), .Y(new_n6178));
  xor_4  g05802(.A(new_n6109), .B(new_n6106), .Y(new_n6179));
  xor_4  g05803(.A(new_n6174), .B(new_n6172), .Y(new_n6180));
  nand_5 g05804(.A(new_n6180), .B(new_n6179), .Y(new_n6181));
  or_6   g05805(.A(new_n3444), .B(new_n3419), .Y(new_n6182));
  nand_5 g05806(.A(new_n3445), .B(new_n3379), .Y(new_n6183));
  nand_5 g05807(.A(new_n6183), .B(new_n6182), .Y(new_n6184));
  xor_4  g05808(.A(new_n6180), .B(new_n6179), .Y(new_n6185));
  nand_5 g05809(.A(new_n6185), .B(new_n6184), .Y(new_n6186));
  nand_5 g05810(.A(new_n6186), .B(new_n6181), .Y(new_n6187));
  xor_4  g05811(.A(new_n6187), .B(new_n6178), .Y(new_n6188));
  not_8  g05812(.A(new_n6188), .Y(new_n6189));
  nand_5 g05813(.A(new_n6189), .B(new_n6036), .Y(new_n6190));
  xor_4  g05814(.A(new_n6189), .B(new_n6036), .Y(new_n6191));
  not_8  g05815(.A(new_n6191), .Y(new_n6192));
  xor_4  g05816(.A(new_n6185), .B(new_n6184), .Y(new_n6193));
  xor_4  g05817(.A(new_n6033), .B(new_n6032), .Y(new_n6194));
  not_8  g05818(.A(new_n6194), .Y(new_n6195));
  nand_5 g05819(.A(new_n6195), .B(new_n6193), .Y(new_n6196));
  not_8  g05820(.A(new_n6196), .Y(new_n6197));
  xor_4  g05821(.A(new_n6194), .B(new_n6193), .Y(new_n6198));
  or_6   g05822(.A(new_n3510), .B(new_n3485), .Y(new_n6199));
  not_8  g05823(.A(new_n3446), .Y(new_n6200));
  nand_5 g05824(.A(new_n3511), .B(new_n6200), .Y(new_n6201));
  nand_5 g05825(.A(new_n6201), .B(new_n6199), .Y(new_n6202));
  nor_5  g05826(.A(new_n6202), .B(new_n6198), .Y(new_n6203));
  nor_5  g05827(.A(new_n6203), .B(new_n6197), .Y(new_n6204));
  or_6   g05828(.A(new_n6204), .B(new_n6192), .Y(new_n6205));
  nand_5 g05829(.A(new_n6205), .B(new_n6190), .Y(new_n6206));
  nand_5 g05830(.A(pi172), .B(pi015), .Y(new_n6207));
  nand_5 g05831(.A(new_n6160), .B(new_n6157), .Y(new_n6208));
  not_8  g05832(.A(new_n6153), .Y(new_n6209));
  nand_5 g05833(.A(new_n6161), .B(new_n6209), .Y(new_n6210));
  nand_5 g05834(.A(new_n6210), .B(new_n6208), .Y(new_n6211));
  xor_4  g05835(.A(new_n6211), .B(new_n6207), .Y(new_n6212));
  xor_4  g05836(.A(new_n6212), .B(new_n6206), .Y(new_n6213));
  xor_4  g05837(.A(new_n6213), .B(new_n5978), .Y(new_n6214));
  nand_5 g05838(.A(pi154), .B(pi090), .Y(new_n6215));
  nand_5 g05839(.A(pi141), .B(pi095), .Y(new_n6216));
  xor_4  g05840(.A(new_n6216), .B(new_n6215), .Y(new_n6217));
  or_6   g05841(.A(new_n6072), .B(new_n6042), .Y(new_n6218));
  not_8  g05842(.A(new_n6071), .Y(new_n6219));
  nand_5 g05843(.A(new_n6073), .B(new_n6219), .Y(new_n6220));
  nand_5 g05844(.A(new_n6220), .B(new_n6218), .Y(new_n6221));
  nand_5 g05845(.A(new_n6069), .B(new_n6068), .Y(new_n6222));
  nand_5 g05846(.A(new_n6070), .B(new_n6041), .Y(new_n6223));
  nand_5 g05847(.A(new_n6223), .B(new_n6222), .Y(new_n6224));
  xor_4  g05848(.A(new_n6224), .B(new_n6221), .Y(new_n6225));
  nand_5 g05849(.A(pi124), .B(pi104), .Y(new_n6226));
  nand_5 g05850(.A(pi215), .B(pi212), .Y(new_n6227));
  xor_4  g05851(.A(new_n6227), .B(new_n6226), .Y(new_n6228));
  xor_4  g05852(.A(new_n6228), .B(new_n6225), .Y(new_n6229));
  nand_5 g05853(.A(pi130), .B(pi013), .Y(new_n6230));
  nand_5 g05854(.A(new_n6076), .B(new_n6052), .Y(new_n6231));
  nand_5 g05855(.A(new_n6077), .B(new_n6075), .Y(new_n6232));
  nand_5 g05856(.A(new_n6232), .B(new_n6231), .Y(new_n6233));
  xor_4  g05857(.A(new_n6233), .B(new_n6230), .Y(new_n6234));
  nand_5 g05858(.A(pi112), .B(pi003), .Y(new_n6235));
  xor_4  g05859(.A(new_n6235), .B(new_n6234), .Y(new_n6236));
  xor_4  g05860(.A(new_n6236), .B(new_n6229), .Y(new_n6237));
  xor_4  g05861(.A(new_n6237), .B(new_n6217), .Y(new_n6238));
  nand_5 g05862(.A(new_n6081), .B(new_n6078), .Y(new_n6239));
  nand_5 g05863(.A(new_n6082), .B(new_n6074), .Y(new_n6240));
  nand_5 g05864(.A(new_n6240), .B(new_n6239), .Y(new_n6241));
  nand_5 g05865(.A(pi158), .B(pi018), .Y(new_n6242));
  xor_4  g05866(.A(new_n6242), .B(new_n6241), .Y(new_n6243));
  xor_4  g05867(.A(new_n6243), .B(new_n6238), .Y(new_n6244));
  or_6   g05868(.A(new_n5964), .B(new_n5935), .Y(new_n6245));
  nand_5 g05869(.A(new_n5965), .B(new_n5961), .Y(new_n6246));
  nand_5 g05870(.A(new_n6246), .B(new_n6245), .Y(new_n6247));
  nand_5 g05871(.A(pi236), .B(pi153), .Y(new_n6248));
  xor_4  g05872(.A(new_n6248), .B(new_n6247), .Y(new_n6249));
  xor_4  g05873(.A(new_n6249), .B(new_n6244), .Y(new_n6250));
  nor_5  g05874(.A(new_n6027), .B(new_n6006), .Y(new_n6251));
  nor_5  g05875(.A(new_n6035), .B(new_n6028), .Y(new_n6252));
  nor_5  g05876(.A(new_n6252), .B(new_n6251), .Y(new_n6253));
  nand_5 g05877(.A(pi161), .B(pi006), .Y(new_n6254));
  nor_5  g05878(.A(new_n5949), .B(new_n5925), .Y(new_n6255));
  nor_5  g05879(.A(new_n5951), .B(new_n5948), .Y(new_n6256));
  or_6   g05880(.A(new_n6256), .B(new_n6255), .Y(new_n6257));
  xor_4  g05881(.A(new_n6257), .B(new_n6254), .Y(new_n6258));
  nand_5 g05882(.A(new_n5959), .B(new_n5956), .Y(new_n6259));
  not_8  g05883(.A(new_n5952), .Y(new_n6260));
  nand_5 g05884(.A(new_n5960), .B(new_n6260), .Y(new_n6261));
  nand_5 g05885(.A(new_n6261), .B(new_n6259), .Y(new_n6262));
  nand_5 g05886(.A(new_n5954), .B(new_n5953), .Y(new_n6263));
  nand_5 g05887(.A(new_n5955), .B(new_n5934), .Y(new_n6264));
  nand_5 g05888(.A(new_n6264), .B(new_n6263), .Y(new_n6265));
  xor_4  g05889(.A(new_n6265), .B(new_n6262), .Y(new_n6266));
  nand_5 g05890(.A(new_n5946), .B(new_n5945), .Y(new_n6267));
  nand_5 g05891(.A(new_n5947), .B(new_n5923), .Y(new_n6268));
  nand_5 g05892(.A(new_n6268), .B(new_n6267), .Y(new_n6269));
  xor_4  g05893(.A(new_n6269), .B(new_n6266), .Y(new_n6270));
  nand_5 g05894(.A(pi241), .B(pi209), .Y(new_n6271));
  nand_5 g05895(.A(pi190), .B(pi034), .Y(new_n6272));
  nand_5 g05896(.A(pi220), .B(pi131), .Y(new_n6273));
  xor_4  g05897(.A(new_n6273), .B(new_n6272), .Y(new_n6274));
  nand_5 g05898(.A(new_n6024), .B(new_n5995), .Y(new_n6275));
  not_8  g05899(.A(new_n6026), .Y(new_n6276));
  nand_5 g05900(.A(new_n6276), .B(new_n6022), .Y(new_n6277));
  nand_5 g05901(.A(new_n6277), .B(new_n6275), .Y(new_n6278));
  xor_4  g05902(.A(new_n6278), .B(new_n6274), .Y(new_n6279));
  xor_4  g05903(.A(new_n6279), .B(new_n6271), .Y(new_n6280));
  xor_4  g05904(.A(new_n6280), .B(new_n6270), .Y(new_n6281));
  xor_4  g05905(.A(new_n6281), .B(new_n6258), .Y(new_n6282));
  nand_5 g05906(.A(pi089), .B(pi047), .Y(new_n6283));
  nand_5 g05907(.A(pi254), .B(pi128), .Y(new_n6284));
  xor_4  g05908(.A(new_n6284), .B(new_n6283), .Y(new_n6285));
  xor_4  g05909(.A(new_n6285), .B(new_n6282), .Y(new_n6286));
  xor_4  g05910(.A(new_n6286), .B(new_n6253), .Y(new_n6287));
  xor_4  g05911(.A(new_n6287), .B(new_n6250), .Y(new_n6288));
  nand_5 g05912(.A(new_n6112), .B(new_n6101), .Y(new_n6289));
  nand_5 g05913(.A(new_n6114), .B(new_n6113), .Y(new_n6290));
  nand_5 g05914(.A(new_n6290), .B(new_n6289), .Y(new_n6291));
  nand_5 g05915(.A(pi198), .B(pi035), .Y(new_n6292));
  nand_5 g05916(.A(pi165), .B(pi139), .Y(new_n6293));
  xor_4  g05917(.A(new_n6293), .B(new_n6292), .Y(new_n6294));
  xor_4  g05918(.A(new_n6294), .B(new_n6291), .Y(new_n6295));
  nand_5 g05919(.A(pi204), .B(pi120), .Y(new_n6296));
  not_8  g05920(.A(new_n6177), .Y(new_n6297));
  nand_5 g05921(.A(new_n6297), .B(new_n6115), .Y(new_n6298));
  or_6   g05922(.A(new_n6187), .B(new_n6178), .Y(new_n6299));
  nand_5 g05923(.A(new_n6299), .B(new_n6298), .Y(new_n6300));
  nand_5 g05924(.A(pi229), .B(pi064), .Y(new_n6301));
  nand_5 g05925(.A(pi185), .B(pi077), .Y(new_n6302));
  nand_5 g05926(.A(pi052), .B(pi030), .Y(new_n6303));
  xor_4  g05927(.A(new_n6303), .B(new_n6302), .Y(new_n6304));
  xor_4  g05928(.A(new_n6304), .B(new_n6301), .Y(new_n6305));
  xor_4  g05929(.A(new_n6305), .B(new_n6300), .Y(new_n6306));
  nand_5 g05930(.A(new_n6020), .B(new_n6017), .Y(new_n6307));
  nand_5 g05931(.A(new_n6021), .B(new_n6013), .Y(new_n6308));
  nand_5 g05932(.A(new_n6308), .B(new_n6307), .Y(new_n6309));
  nand_5 g05933(.A(new_n6015), .B(new_n5994), .Y(new_n6310));
  nand_5 g05934(.A(new_n6016), .B(new_n6014), .Y(new_n6311));
  nand_5 g05935(.A(new_n6311), .B(new_n6310), .Y(new_n6312));
  xor_4  g05936(.A(new_n6312), .B(new_n6309), .Y(new_n6313));
  nand_5 g05937(.A(pi189), .B(pi067), .Y(new_n6314));
  nand_5 g05938(.A(pi133), .B(pi053), .Y(new_n6315));
  xor_4  g05939(.A(new_n6315), .B(new_n6314), .Y(new_n6316));
  xor_4  g05940(.A(new_n6316), .B(new_n6313), .Y(new_n6317));
  or_6   g05941(.A(new_n6167), .B(new_n6145), .Y(new_n6318));
  nand_5 g05942(.A(new_n6176), .B(new_n6168), .Y(new_n6319));
  nand_5 g05943(.A(new_n6319), .B(new_n6318), .Y(new_n6320));
  nand_5 g05944(.A(pi092), .B(pi084), .Y(new_n6321));
  xor_4  g05945(.A(new_n6321), .B(new_n6320), .Y(new_n6322));
  xor_4  g05946(.A(new_n6322), .B(new_n6317), .Y(new_n6323));
  nand_5 g05947(.A(pi146), .B(pi062), .Y(new_n6324));
  nand_5 g05948(.A(pi168), .B(pi078), .Y(new_n6325));
  xor_4  g05949(.A(new_n6325), .B(new_n6324), .Y(new_n6326));
  nand_5 g05950(.A(pi152), .B(pi065), .Y(new_n6327));
  or_6   g05951(.A(new_n6165), .B(new_n6136), .Y(new_n6328));
  nand_5 g05952(.A(new_n6166), .B(new_n6162), .Y(new_n6329));
  nand_5 g05953(.A(new_n6329), .B(new_n6328), .Y(new_n6330));
  xor_4  g05954(.A(new_n6330), .B(new_n6327), .Y(new_n6331));
  xor_4  g05955(.A(new_n6331), .B(new_n6326), .Y(new_n6332));
  nand_5 g05956(.A(new_n6008), .B(new_n6007), .Y(new_n6333));
  nand_5 g05957(.A(new_n6009), .B(new_n5987), .Y(new_n6334));
  nand_5 g05958(.A(new_n6334), .B(new_n6333), .Y(new_n6335));
  or_6   g05959(.A(new_n6011), .B(new_n5988), .Y(new_n6336));
  not_8  g05960(.A(new_n6010), .Y(new_n6337));
  nand_5 g05961(.A(new_n6012), .B(new_n6337), .Y(new_n6338));
  nand_5 g05962(.A(new_n6338), .B(new_n6336), .Y(new_n6339));
  xor_4  g05963(.A(new_n6339), .B(new_n6335), .Y(new_n6340));
  xor_4  g05964(.A(new_n6340), .B(new_n6332), .Y(new_n6341));
  xor_4  g05965(.A(new_n6341), .B(new_n6323), .Y(new_n6342));
  xor_4  g05966(.A(new_n6342), .B(new_n6306), .Y(new_n6343));
  xor_4  g05967(.A(new_n6343), .B(new_n6296), .Y(new_n6344));
  xor_4  g05968(.A(new_n6344), .B(new_n6295), .Y(new_n6345));
  nand_5 g05969(.A(pi213), .B(pi022), .Y(new_n6346));
  or_6   g05970(.A(new_n6090), .B(new_n6067), .Y(new_n6347));
  nand_5 g05971(.A(new_n6100), .B(new_n6091), .Y(new_n6348));
  nand_5 g05972(.A(new_n6348), .B(new_n6347), .Y(new_n6349));
  xor_4  g05973(.A(new_n6349), .B(new_n6346), .Y(new_n6350));
  nand_5 g05974(.A(new_n6155), .B(new_n6154), .Y(new_n6351));
  nand_5 g05975(.A(new_n6156), .B(new_n6135), .Y(new_n6352));
  nand_5 g05976(.A(new_n6352), .B(new_n6351), .Y(new_n6353));
  nor_5  g05977(.A(new_n6089), .B(new_n6083), .Y(new_n6354));
  nor_5  g05978(.A(new_n6354), .B(new_n6088), .Y(new_n6355));
  xor_4  g05979(.A(new_n6355), .B(new_n6353), .Y(new_n6356));
  nand_5 g05980(.A(pi183), .B(pi004), .Y(new_n6357));
  nand_5 g05981(.A(pi105), .B(pi073), .Y(new_n6358));
  xor_4  g05982(.A(new_n6358), .B(new_n6357), .Y(new_n6359));
  nand_5 g05983(.A(pi170), .B(pi088), .Y(new_n6360));
  xor_4  g05984(.A(new_n6360), .B(new_n6359), .Y(new_n6361));
  xor_4  g05985(.A(new_n6361), .B(new_n6356), .Y(new_n6362));
  xor_4  g05986(.A(new_n6362), .B(new_n6350), .Y(new_n6363));
  nand_5 g05987(.A(pi208), .B(pi197), .Y(new_n6364));
  nand_5 g05988(.A(new_n6147), .B(new_n6146), .Y(new_n6365));
  nand_5 g05989(.A(new_n6148), .B(new_n6127), .Y(new_n6366));
  nand_5 g05990(.A(new_n6366), .B(new_n6365), .Y(new_n6367));
  nor_5  g05991(.A(new_n6150), .B(new_n6129), .Y(new_n6368));
  nor_5  g05992(.A(new_n6152), .B(new_n6149), .Y(new_n6369));
  or_6   g05993(.A(new_n6369), .B(new_n6368), .Y(new_n6370));
  xor_4  g05994(.A(new_n6370), .B(new_n6367), .Y(new_n6371));
  xor_4  g05995(.A(new_n6371), .B(new_n6364), .Y(new_n6372));
  xor_4  g05996(.A(new_n6372), .B(new_n6363), .Y(new_n6373));
  xor_4  g05997(.A(new_n6373), .B(new_n6345), .Y(new_n6374));
  xor_4  g05998(.A(new_n6374), .B(new_n6288), .Y(new_n6375));
  xor_4  g05999(.A(new_n6375), .B(new_n6214), .Y(po027));
  nand_5 g06000(.A(pi141), .B(pi108), .Y(new_n6377));
  nand_5 g06001(.A(new_n4599), .B(new_n4598), .Y(new_n6378));
  nand_5 g06002(.A(new_n4600), .B(new_n4597), .Y(new_n6379));
  nand_5 g06003(.A(new_n6379), .B(new_n6378), .Y(new_n6380));
  xnor_4 g06004(.A(new_n6380), .B(new_n6377), .Y(new_n6381));
  nand_5 g06005(.A(pi090), .B(pi042), .Y(new_n6382));
  nand_5 g06006(.A(pi051), .B(pi047), .Y(new_n6383));
  nand_5 g06007(.A(new_n6383), .B(new_n6382), .Y(new_n6384));
  nand_5 g06008(.A(pi047), .B(pi042), .Y(new_n6385));
  or_6   g06009(.A(new_n6385), .B(new_n4598), .Y(new_n6386));
  nand_5 g06010(.A(new_n6386), .B(new_n6384), .Y(new_n6387));
  xnor_4 g06011(.A(new_n6387), .B(new_n6381), .Y(new_n6388));
  nand_5 g06012(.A(pi161), .B(pi007), .Y(new_n6389));
  nand_5 g06013(.A(pi241), .B(pi118), .Y(new_n6390));
  and_6  g06014(.A(new_n6390), .B(new_n6389), .Y(new_n6391));
  nand_5 g06015(.A(pi161), .B(pi118), .Y(new_n6392));
  nor_5  g06016(.A(new_n6392), .B(new_n4602), .Y(new_n6393));
  or_6   g06017(.A(new_n6393), .B(new_n6391), .Y(new_n6394));
  xnor_4 g06018(.A(new_n6394), .B(new_n6388), .Y(new_n6395));
  nand_5 g06019(.A(new_n4605), .B(new_n4602), .Y(new_n6396));
  nand_5 g06020(.A(new_n4606), .B(new_n4601), .Y(new_n6397));
  nand_5 g06021(.A(new_n6397), .B(new_n6396), .Y(new_n6398));
  xor_4  g06022(.A(new_n6398), .B(new_n6395), .Y(new_n6399));
  not_8  g06023(.A(new_n4608), .Y(new_n6400));
  nand_5 g06024(.A(new_n4612), .B(new_n6400), .Y(new_n6401));
  or_6   g06025(.A(new_n4613), .B(new_n4607), .Y(new_n6402));
  nand_5 g06026(.A(new_n6402), .B(new_n6401), .Y(new_n6403));
  xnor_4 g06027(.A(new_n6403), .B(new_n6399), .Y(new_n6404));
  nand_5 g06028(.A(new_n4614), .B(new_n4596), .Y(new_n6405));
  nand_5 g06029(.A(pi236), .B(pi113), .Y(new_n6406));
  xor_4  g06030(.A(new_n6406), .B(new_n6405), .Y(new_n6407));
  xnor_4 g06031(.A(new_n6407), .B(new_n6404), .Y(new_n6408));
  or_6   g06032(.A(new_n4652), .B(new_n4635), .Y(new_n6409));
  nand_5 g06033(.A(pi061), .B(pi013), .Y(new_n6410));
  nand_5 g06034(.A(pi188), .B(pi105), .Y(new_n6411));
  nand_5 g06035(.A(pi178), .B(pi112), .Y(new_n6412));
  nand_5 g06036(.A(new_n6412), .B(new_n6411), .Y(new_n6413));
  nand_5 g06037(.A(pi178), .B(pi105), .Y(new_n6414));
  or_6   g06038(.A(new_n6414), .B(new_n4636), .Y(new_n6415));
  nand_5 g06039(.A(new_n6415), .B(new_n6413), .Y(new_n6416));
  xor_4  g06040(.A(new_n6416), .B(new_n6410), .Y(new_n6417));
  nand_5 g06041(.A(new_n4638), .B(new_n4637), .Y(new_n6418));
  nand_5 g06042(.A(new_n4639), .B(new_n4636), .Y(new_n6419));
  nand_5 g06043(.A(new_n6419), .B(new_n6418), .Y(new_n6420));
  xor_4  g06044(.A(new_n6420), .B(new_n6417), .Y(new_n6421));
  nand_5 g06045(.A(pi104), .B(pi012), .Y(new_n6422));
  nand_5 g06046(.A(pi212), .B(pi144), .Y(new_n6423));
  and_6  g06047(.A(new_n6423), .B(new_n6422), .Y(new_n6424));
  nand_5 g06048(.A(pi144), .B(pi104), .Y(new_n6425));
  nor_5  g06049(.A(new_n6425), .B(new_n4641), .Y(new_n6426));
  or_6   g06050(.A(new_n6426), .B(new_n6424), .Y(new_n6427));
  xnor_4 g06051(.A(new_n6427), .B(new_n6421), .Y(new_n6428));
  nand_5 g06052(.A(new_n4644), .B(new_n4641), .Y(new_n6429));
  nand_5 g06053(.A(new_n4645), .B(new_n4640), .Y(new_n6430));
  nand_5 g06054(.A(new_n6430), .B(new_n6429), .Y(new_n6431));
  xor_4  g06055(.A(new_n6431), .B(new_n6428), .Y(new_n6432));
  or_6   g06056(.A(new_n4650), .B(new_n4647), .Y(new_n6433));
  nand_5 g06057(.A(new_n4651), .B(new_n4646), .Y(new_n6434));
  nand_5 g06058(.A(new_n6434), .B(new_n6433), .Y(new_n6435));
  xnor_4 g06059(.A(new_n6435), .B(new_n6432), .Y(new_n6436));
  nand_5 g06060(.A(pi213), .B(pi098), .Y(new_n6437));
  xor_4  g06061(.A(new_n6437), .B(new_n6436), .Y(new_n6438));
  xor_4  g06062(.A(new_n6438), .B(new_n6409), .Y(new_n6439));
  xor_4  g06063(.A(new_n6439), .B(new_n6408), .Y(new_n6440));
  nand_5 g06064(.A(new_n4653), .B(new_n4615), .Y(new_n6441));
  not_8  g06065(.A(new_n4681), .Y(new_n6442));
  nand_5 g06066(.A(new_n6442), .B(new_n4654), .Y(new_n6443));
  nand_5 g06067(.A(new_n6443), .B(new_n6441), .Y(new_n6444));
  xnor_4 g06068(.A(new_n6444), .B(new_n6440), .Y(new_n6445));
  nand_5 g06069(.A(pi179), .B(pi035), .Y(new_n6446));
  nand_5 g06070(.A(pi033), .B(pi015), .Y(new_n6447));
  nand_5 g06071(.A(pi204), .B(pi162), .Y(new_n6448));
  nand_5 g06072(.A(new_n6448), .B(new_n6447), .Y(new_n6449));
  nand_5 g06073(.A(pi204), .B(pi033), .Y(new_n6450));
  or_6   g06074(.A(new_n6450), .B(new_n4705), .Y(new_n6451));
  nand_5 g06075(.A(new_n6451), .B(new_n6449), .Y(new_n6452));
  xor_4  g06076(.A(new_n6452), .B(new_n6446), .Y(new_n6453));
  nand_5 g06077(.A(new_n4705), .B(new_n4704), .Y(new_n6454));
  nand_5 g06078(.A(new_n4706), .B(new_n4703), .Y(new_n6455));
  nand_5 g06079(.A(new_n6455), .B(new_n6454), .Y(new_n6456));
  xor_4  g06080(.A(new_n6456), .B(new_n6453), .Y(new_n6457));
  nand_5 g06081(.A(pi139), .B(pi048), .Y(new_n6458));
  nand_5 g06082(.A(pi237), .B(pi208), .Y(new_n6459));
  and_6  g06083(.A(new_n6459), .B(new_n6458), .Y(new_n6460));
  nand_5 g06084(.A(pi237), .B(pi139), .Y(new_n6461));
  nor_5  g06085(.A(new_n6461), .B(new_n4708), .Y(new_n6462));
  or_6   g06086(.A(new_n6462), .B(new_n6460), .Y(new_n6463));
  xnor_4 g06087(.A(new_n6463), .B(new_n6457), .Y(new_n6464));
  nand_5 g06088(.A(new_n4711), .B(new_n4708), .Y(new_n6465));
  nand_5 g06089(.A(new_n4712), .B(new_n4707), .Y(new_n6466));
  nand_5 g06090(.A(new_n6466), .B(new_n6465), .Y(new_n6467));
  xor_4  g06091(.A(new_n6467), .B(new_n6464), .Y(new_n6468));
  not_8  g06092(.A(new_n4714), .Y(new_n6469));
  nand_5 g06093(.A(new_n4717), .B(new_n6469), .Y(new_n6470));
  or_6   g06094(.A(new_n4718), .B(new_n4713), .Y(new_n6471));
  nand_5 g06095(.A(new_n6471), .B(new_n6470), .Y(new_n6472));
  xnor_4 g06096(.A(new_n6472), .B(new_n6468), .Y(new_n6473));
  nand_5 g06097(.A(new_n4719), .B(new_n4702), .Y(new_n6474));
  nand_5 g06098(.A(pi238), .B(pi168), .Y(new_n6475));
  xor_4  g06099(.A(new_n6475), .B(new_n6474), .Y(new_n6476));
  xor_4  g06100(.A(new_n6476), .B(new_n6473), .Y(new_n6477));
  or_6   g06101(.A(new_n4745), .B(new_n4720), .Y(new_n6478));
  nand_5 g06102(.A(new_n4746), .B(new_n4682), .Y(new_n6479));
  nand_5 g06103(.A(new_n6479), .B(new_n6478), .Y(new_n6480));
  xor_4  g06104(.A(new_n6480), .B(new_n6477), .Y(new_n6481));
  xor_4  g06105(.A(new_n6481), .B(new_n6445), .Y(new_n6482));
  nand_5 g06106(.A(pi194), .B(pi133), .Y(new_n6483));
  nand_5 g06107(.A(pi143), .B(pi064), .Y(new_n6484));
  nand_5 g06108(.A(pi189), .B(pi057), .Y(new_n6485));
  nand_5 g06109(.A(new_n6485), .B(new_n6484), .Y(new_n6486));
  nand_5 g06110(.A(pi064), .B(pi057), .Y(new_n6487));
  or_6   g06111(.A(new_n6487), .B(new_n4772), .Y(new_n6488));
  nand_5 g06112(.A(new_n6488), .B(new_n6486), .Y(new_n6489));
  xor_4  g06113(.A(new_n6489), .B(new_n6483), .Y(new_n6490));
  nand_5 g06114(.A(new_n4773), .B(new_n4772), .Y(new_n6491));
  nand_5 g06115(.A(new_n4774), .B(new_n4771), .Y(new_n6492));
  nand_5 g06116(.A(new_n6492), .B(new_n6491), .Y(new_n6493));
  xor_4  g06117(.A(new_n6493), .B(new_n6490), .Y(new_n6494));
  nand_5 g06118(.A(pi085), .B(pi077), .Y(new_n6495));
  nand_5 g06119(.A(pi180), .B(pi052), .Y(new_n6496));
  nand_5 g06120(.A(new_n6496), .B(new_n6495), .Y(new_n6497));
  nand_5 g06121(.A(pi180), .B(pi077), .Y(new_n6498));
  nor_5  g06122(.A(new_n6498), .B(new_n4776), .Y(new_n6499));
  not_8  g06123(.A(new_n6499), .Y(new_n6500));
  nand_5 g06124(.A(new_n6500), .B(new_n6497), .Y(new_n6501));
  xnor_4 g06125(.A(new_n6501), .B(new_n6494), .Y(new_n6502));
  nand_5 g06126(.A(new_n4779), .B(new_n4776), .Y(new_n6503));
  nand_5 g06127(.A(new_n4780), .B(new_n4775), .Y(new_n6504));
  nand_5 g06128(.A(new_n6504), .B(new_n6503), .Y(new_n6505));
  xor_4  g06129(.A(new_n6505), .B(new_n6502), .Y(new_n6506));
  or_6   g06130(.A(new_n4782), .B(new_n4781), .Y(new_n6507));
  nand_5 g06131(.A(new_n4786), .B(new_n4783), .Y(new_n6508));
  nand_5 g06132(.A(new_n6508), .B(new_n6507), .Y(new_n6509));
  xnor_4 g06133(.A(new_n6509), .B(new_n6506), .Y(new_n6510));
  nand_5 g06134(.A(new_n4787), .B(new_n4770), .Y(new_n6511));
  nand_5 g06135(.A(pi131), .B(pi036), .Y(new_n6512));
  xor_4  g06136(.A(new_n6512), .B(new_n6511), .Y(new_n6513));
  xor_4  g06137(.A(new_n6513), .B(new_n6510), .Y(new_n6514));
  not_8  g06138(.A(new_n4788), .Y(new_n6515));
  nor_5  g06139(.A(new_n6515), .B(new_n4747), .Y(new_n6516));
  nor_5  g06140(.A(new_n4810), .B(new_n4789), .Y(new_n6517));
  nor_5  g06141(.A(new_n6517), .B(new_n6516), .Y(new_n6518));
  xor_4  g06142(.A(new_n6518), .B(new_n6514), .Y(new_n6519));
  xor_4  g06143(.A(new_n6519), .B(new_n6482), .Y(po028));
  xnor_4 g06144(.A(new_n881), .B(new_n880), .Y(po029));
  xor_4  g06145(.A(new_n1820), .B(new_n1819), .Y(po030));
  nand_5 g06146(.A(pi210), .B(pi163), .Y(new_n6523));
  nand_5 g06147(.A(pi242), .B(pi107), .Y(new_n6524));
  xor_4  g06148(.A(new_n6524), .B(new_n6523), .Y(new_n6525));
  nand_5 g06149(.A(pi249), .B(pi175), .Y(new_n6526));
  xor_4  g06150(.A(new_n6526), .B(new_n6525), .Y(new_n6527));
  nand_5 g06151(.A(pi217), .B(pi103), .Y(new_n6528));
  xor_4  g06152(.A(new_n6528), .B(new_n6527), .Y(po031));
  xor_4  g06153(.A(new_n2569), .B(new_n2551), .Y(po032));
  nand_5 g06154(.A(pi171), .B(pi140), .Y(new_n6531));
  nand_5 g06155(.A(pi252), .B(pi107), .Y(new_n6532));
  xor_4  g06156(.A(new_n6532), .B(new_n6531), .Y(new_n6533));
  nand_5 g06157(.A(pi242), .B(pi049), .Y(new_n6534));
  xor_4  g06158(.A(new_n6534), .B(new_n6533), .Y(new_n6535));
  nor_5  g06159(.A(new_n6531), .B(new_n6524), .Y(new_n6536));
  xor_4  g06160(.A(new_n6536), .B(new_n6535), .Y(new_n6537));
  not_8  g06161(.A(new_n6523), .Y(new_n6538));
  nand_5 g06162(.A(pi148), .B(pi111), .Y(new_n6539));
  nor_5  g06163(.A(new_n6539), .B(new_n6538), .Y(new_n6540));
  nand_5 g06164(.A(pi228), .B(pi210), .Y(new_n6541));
  nand_5 g06165(.A(pi163), .B(pi024), .Y(new_n6542));
  nand_5 g06166(.A(new_n6542), .B(new_n6541), .Y(new_n6543));
  or_6   g06167(.A(new_n6542), .B(new_n6541), .Y(new_n6544));
  and_6  g06168(.A(new_n6544), .B(new_n6543), .Y(new_n6545));
  or_6   g06169(.A(new_n6545), .B(new_n6540), .Y(new_n6546));
  nand_5 g06170(.A(new_n6543), .B(new_n6540), .Y(new_n6547));
  nand_5 g06171(.A(new_n6547), .B(new_n6546), .Y(new_n6548));
  xor_4  g06172(.A(new_n6548), .B(new_n6537), .Y(new_n6549));
  or_6   g06173(.A(new_n6524), .B(new_n6523), .Y(new_n6550));
  nand_5 g06174(.A(pi210), .B(pi148), .Y(new_n6551));
  nand_5 g06175(.A(pi163), .B(pi111), .Y(new_n6552));
  nand_5 g06176(.A(new_n6552), .B(new_n6551), .Y(new_n6553));
  or_6   g06177(.A(new_n6539), .B(new_n6523), .Y(new_n6554));
  nand_5 g06178(.A(new_n6554), .B(new_n6553), .Y(new_n6555));
  nor_5  g06179(.A(new_n6555), .B(new_n6550), .Y(new_n6556));
  xnor_4 g06180(.A(new_n6555), .B(new_n6550), .Y(new_n6557));
  not_8  g06181(.A(new_n6536), .Y(new_n6558));
  nand_5 g06182(.A(pi140), .B(pi107), .Y(new_n6559));
  nand_5 g06183(.A(pi242), .B(pi171), .Y(new_n6560));
  nand_5 g06184(.A(new_n6560), .B(new_n6559), .Y(new_n6561));
  nand_5 g06185(.A(new_n6561), .B(new_n6558), .Y(new_n6562));
  nor_5  g06186(.A(new_n6562), .B(new_n6557), .Y(new_n6563));
  nor_5  g06187(.A(new_n6563), .B(new_n6556), .Y(new_n6564));
  not_8  g06188(.A(new_n6564), .Y(new_n6565));
  xor_4  g06189(.A(new_n6565), .B(new_n6549), .Y(new_n6566));
  not_8  g06190(.A(new_n6525), .Y(new_n6567));
  nor_5  g06191(.A(new_n6526), .B(new_n6567), .Y(new_n6568));
  nand_5 g06192(.A(pi249), .B(pi134), .Y(new_n6569));
  nand_5 g06193(.A(pi222), .B(pi175), .Y(new_n6570));
  xor_4  g06194(.A(new_n6570), .B(new_n6569), .Y(new_n6571));
  or_6   g06195(.A(new_n6571), .B(new_n6568), .Y(new_n6572));
  xor_4  g06196(.A(new_n6562), .B(new_n6557), .Y(new_n6573));
  not_8  g06197(.A(new_n6573), .Y(new_n6574));
  xor_4  g06198(.A(new_n6571), .B(new_n6568), .Y(new_n6575));
  nand_5 g06199(.A(new_n6575), .B(new_n6574), .Y(new_n6576));
  nand_5 g06200(.A(new_n6576), .B(new_n6572), .Y(new_n6577));
  nand_5 g06201(.A(pi249), .B(pi240), .Y(new_n6578));
  nand_5 g06202(.A(pi175), .B(pi125), .Y(new_n6579));
  nand_5 g06203(.A(new_n6579), .B(new_n6578), .Y(new_n6580));
  not_8  g06204(.A(new_n6580), .Y(new_n6581));
  nand_5 g06205(.A(pi222), .B(pi134), .Y(new_n6582));
  not_8  g06206(.A(new_n6582), .Y(new_n6583));
  nand_5 g06207(.A(new_n6583), .B(new_n6526), .Y(new_n6584));
  nor_5  g06208(.A(new_n6584), .B(new_n6581), .Y(new_n6585));
  nand_5 g06209(.A(new_n6584), .B(new_n6581), .Y(new_n6586));
  or_6   g06210(.A(new_n6579), .B(new_n6578), .Y(new_n6587));
  nand_5 g06211(.A(new_n6587), .B(new_n6586), .Y(new_n6588));
  or_6   g06212(.A(new_n6588), .B(new_n6585), .Y(new_n6589));
  xor_4  g06213(.A(new_n6589), .B(new_n6577), .Y(new_n6590));
  not_8  g06214(.A(new_n6590), .Y(new_n6591));
  xor_4  g06215(.A(new_n6591), .B(new_n6566), .Y(new_n6592));
  or_6   g06216(.A(new_n6528), .B(new_n6527), .Y(new_n6593));
  nand_5 g06217(.A(pi103), .B(pi100), .Y(new_n6594));
  nand_5 g06218(.A(pi217), .B(pi117), .Y(new_n6595));
  nand_5 g06219(.A(new_n6595), .B(new_n6594), .Y(new_n6596));
  nand_5 g06220(.A(pi117), .B(pi100), .Y(new_n6597));
  or_6   g06221(.A(new_n6597), .B(new_n6528), .Y(new_n6598));
  nand_5 g06222(.A(new_n6598), .B(new_n6596), .Y(new_n6599));
  or_6   g06223(.A(new_n6599), .B(new_n6593), .Y(new_n6600));
  xor_4  g06224(.A(new_n6575), .B(new_n6573), .Y(new_n6601));
  xor_4  g06225(.A(new_n6599), .B(new_n6593), .Y(new_n6602));
  nand_5 g06226(.A(new_n6602), .B(new_n6601), .Y(new_n6603));
  nand_5 g06227(.A(new_n6603), .B(new_n6600), .Y(new_n6604));
  not_8  g06228(.A(new_n6528), .Y(new_n6605));
  nor_5  g06229(.A(new_n6597), .B(new_n6605), .Y(new_n6606));
  nand_5 g06230(.A(pi227), .B(pi103), .Y(new_n6607));
  nand_5 g06231(.A(pi217), .B(pi016), .Y(new_n6608));
  nand_5 g06232(.A(new_n6608), .B(new_n6607), .Y(new_n6609));
  or_6   g06233(.A(new_n6608), .B(new_n6607), .Y(new_n6610));
  and_6  g06234(.A(new_n6610), .B(new_n6609), .Y(new_n6611));
  nor_5  g06235(.A(new_n6611), .B(new_n6606), .Y(new_n6612));
  not_8  g06236(.A(new_n6612), .Y(new_n6613));
  nand_5 g06237(.A(new_n6609), .B(new_n6606), .Y(new_n6614));
  and_6  g06238(.A(new_n6614), .B(new_n6613), .Y(new_n6615));
  xor_4  g06239(.A(new_n6615), .B(new_n6604), .Y(new_n6616));
  xnor_4 g06240(.A(new_n6616), .B(new_n6592), .Y(po033));
  xor_4  g06241(.A(new_n4566), .B(new_n4564), .Y(po034));
  xor_4  g06242(.A(new_n4041), .B(new_n4040), .Y(po035));
  nand_5 g06243(.A(pi227), .B(pi080), .Y(new_n6620));
  nand_5 g06244(.A(pi234), .B(pi217), .Y(new_n6621));
  nand_5 g06245(.A(pi247), .B(pi100), .Y(new_n6622));
  nand_5 g06246(.A(new_n6622), .B(new_n6621), .Y(new_n6623));
  nand_5 g06247(.A(pi247), .B(pi217), .Y(new_n6624));
  nand_5 g06248(.A(pi234), .B(pi100), .Y(new_n6625));
  or_6   g06249(.A(new_n6625), .B(new_n6624), .Y(new_n6626));
  nand_5 g06250(.A(new_n6626), .B(new_n6623), .Y(new_n6627));
  xor_4  g06251(.A(new_n6627), .B(new_n6620), .Y(new_n6628));
  nand_5 g06252(.A(pi227), .B(pi016), .Y(new_n6629));
  nand_5 g06253(.A(pi100), .B(pi080), .Y(new_n6630));
  nand_5 g06254(.A(new_n6630), .B(new_n6629), .Y(new_n6631));
  xor_4  g06255(.A(new_n6630), .B(new_n6629), .Y(new_n6632));
  nand_5 g06256(.A(new_n6632), .B(new_n6624), .Y(new_n6633));
  nand_5 g06257(.A(new_n6633), .B(new_n6631), .Y(new_n6634));
  xor_4  g06258(.A(new_n6634), .B(new_n6628), .Y(new_n6635));
  nand_5 g06259(.A(pi081), .B(pi016), .Y(new_n6636));
  nand_5 g06260(.A(pi117), .B(pi106), .Y(new_n6637));
  nand_5 g06261(.A(new_n6637), .B(new_n6636), .Y(new_n6638));
  nand_5 g06262(.A(pi106), .B(pi016), .Y(new_n6639));
  nand_5 g06263(.A(pi117), .B(pi081), .Y(new_n6640));
  nor_5  g06264(.A(new_n6640), .B(new_n6639), .Y(new_n6641));
  not_8  g06265(.A(new_n6641), .Y(new_n6642));
  nand_5 g06266(.A(new_n6642), .B(new_n6638), .Y(new_n6643));
  xnor_4 g06267(.A(new_n6643), .B(new_n6635), .Y(new_n6644));
  nand_5 g06268(.A(pi100), .B(pi016), .Y(new_n6645));
  nand_5 g06269(.A(pi217), .B(pi080), .Y(new_n6646));
  nand_5 g06270(.A(new_n6646), .B(new_n6645), .Y(new_n6647));
  nand_5 g06271(.A(pi227), .B(pi117), .Y(new_n6648));
  xor_4  g06272(.A(new_n6646), .B(new_n6645), .Y(new_n6649));
  nand_5 g06273(.A(new_n6649), .B(new_n6648), .Y(new_n6650));
  nand_5 g06274(.A(new_n6650), .B(new_n6647), .Y(new_n6651));
  nand_5 g06275(.A(new_n6651), .B(new_n6640), .Y(new_n6652));
  xor_4  g06276(.A(new_n6632), .B(new_n6624), .Y(new_n6653));
  xor_4  g06277(.A(new_n6651), .B(new_n6640), .Y(new_n6654));
  nand_5 g06278(.A(new_n6654), .B(new_n6653), .Y(new_n6655));
  nand_5 g06279(.A(new_n6655), .B(new_n6652), .Y(new_n6656));
  xor_4  g06280(.A(new_n6656), .B(new_n6644), .Y(new_n6657));
  xor_4  g06281(.A(new_n6654), .B(new_n6653), .Y(new_n6658));
  nand_5 g06282(.A(pi106), .B(pi103), .Y(new_n6659));
  or_6   g06283(.A(new_n6659), .B(new_n6658), .Y(new_n6660));
  xor_4  g06284(.A(new_n6659), .B(new_n6658), .Y(new_n6661));
  nand_5 g06285(.A(pi103), .B(pi081), .Y(new_n6662));
  nand_5 g06286(.A(new_n6610), .B(new_n6597), .Y(new_n6663));
  nand_5 g06287(.A(new_n6663), .B(new_n6609), .Y(new_n6664));
  or_6   g06288(.A(new_n6664), .B(new_n6662), .Y(new_n6665));
  xnor_4 g06289(.A(new_n6649), .B(new_n6648), .Y(new_n6666));
  xor_4  g06290(.A(new_n6664), .B(new_n6662), .Y(new_n6667));
  nand_5 g06291(.A(new_n6667), .B(new_n6666), .Y(new_n6668));
  nand_5 g06292(.A(new_n6668), .B(new_n6665), .Y(new_n6669));
  nand_5 g06293(.A(new_n6669), .B(new_n6661), .Y(new_n6670));
  nand_5 g06294(.A(new_n6670), .B(new_n6660), .Y(new_n6671));
  nand_5 g06295(.A(new_n6671), .B(new_n6657), .Y(new_n6672));
  nand_5 g06296(.A(pi217), .B(pi214), .Y(new_n6673));
  nand_5 g06297(.A(pi247), .B(pi227), .Y(new_n6674));
  xor_4  g06298(.A(new_n6674), .B(new_n6673), .Y(new_n6675));
  xor_4  g06299(.A(new_n6675), .B(new_n6625), .Y(new_n6676));
  nand_5 g06300(.A(pi081), .B(pi080), .Y(new_n6677));
  xor_4  g06301(.A(new_n6677), .B(new_n6626), .Y(new_n6678));
  xor_4  g06302(.A(new_n6678), .B(new_n6676), .Y(new_n6679));
  nand_5 g06303(.A(pi233), .B(pi117), .Y(new_n6680));
  nand_5 g06304(.A(pi187), .B(pi103), .Y(new_n6681));
  xor_4  g06305(.A(new_n6681), .B(new_n6680), .Y(new_n6682));
  xor_4  g06306(.A(new_n6682), .B(new_n6639), .Y(new_n6683));
  nand_5 g06307(.A(new_n6627), .B(new_n6620), .Y(new_n6684));
  nand_5 g06308(.A(new_n6634), .B(new_n6628), .Y(new_n6685));
  nand_5 g06309(.A(new_n6685), .B(new_n6684), .Y(new_n6686));
  xor_4  g06310(.A(new_n6686), .B(new_n6683), .Y(new_n6687));
  xnor_4 g06311(.A(new_n6687), .B(new_n6679), .Y(new_n6688));
  nor_5  g06312(.A(new_n6656), .B(new_n6644), .Y(new_n6689));
  and_6  g06313(.A(new_n6689), .B(new_n6641), .Y(new_n6690));
  or_6   g06314(.A(new_n6643), .B(new_n6635), .Y(new_n6691));
  nand_5 g06315(.A(new_n6691), .B(new_n6642), .Y(new_n6692));
  nor_5  g06316(.A(new_n6692), .B(new_n6689), .Y(new_n6693));
  or_6   g06317(.A(new_n6693), .B(new_n6690), .Y(new_n6694));
  xor_4  g06318(.A(new_n6694), .B(new_n6688), .Y(new_n6695));
  xnor_4 g06319(.A(new_n6695), .B(new_n6672), .Y(new_n6696));
  nand_5 g06320(.A(pi233), .B(pi103), .Y(new_n6697));
  xor_4  g06321(.A(new_n6667), .B(new_n6666), .Y(new_n6698));
  nor_5  g06322(.A(new_n6613), .B(new_n6598), .Y(new_n6699));
  nand_5 g06323(.A(new_n6699), .B(new_n6698), .Y(new_n6700));
  not_8  g06324(.A(new_n6700), .Y(new_n6701));
  xor_4  g06325(.A(new_n6669), .B(new_n6661), .Y(new_n6702));
  nand_5 g06326(.A(new_n6702), .B(new_n6701), .Y(new_n6703));
  nand_5 g06327(.A(new_n6703), .B(new_n6697), .Y(new_n6704));
  xnor_4 g06328(.A(new_n6671), .B(new_n6657), .Y(new_n6705));
  xor_4  g06329(.A(new_n6703), .B(new_n6697), .Y(new_n6706));
  nand_5 g06330(.A(new_n6706), .B(new_n6705), .Y(new_n6707));
  nand_5 g06331(.A(new_n6707), .B(new_n6704), .Y(new_n6708));
  xor_4  g06332(.A(new_n6708), .B(new_n6696), .Y(new_n6709));
  or_6   g06333(.A(new_n6558), .B(new_n6535), .Y(new_n6710));
  nand_5 g06334(.A(pi121), .B(pi107), .Y(new_n6711));
  nand_5 g06335(.A(new_n6532), .B(new_n6531), .Y(new_n6712));
  nand_5 g06336(.A(new_n6534), .B(new_n6533), .Y(new_n6713));
  nand_5 g06337(.A(new_n6713), .B(new_n6712), .Y(new_n6714));
  xor_4  g06338(.A(new_n6714), .B(new_n6711), .Y(new_n6715));
  nand_5 g06339(.A(pi252), .B(pi171), .Y(new_n6716));
  nand_5 g06340(.A(pi245), .B(pi242), .Y(new_n6717));
  nand_5 g06341(.A(pi140), .B(pi049), .Y(new_n6718));
  xor_4  g06342(.A(new_n6718), .B(new_n6717), .Y(new_n6719));
  xnor_4 g06343(.A(new_n6719), .B(new_n6716), .Y(new_n6720));
  xnor_4 g06344(.A(new_n6720), .B(new_n6715), .Y(new_n6721));
  nor_5  g06345(.A(new_n6721), .B(new_n6710), .Y(new_n6722));
  nand_5 g06346(.A(pi252), .B(pi049), .Y(new_n6723));
  nand_5 g06347(.A(pi242), .B(pi201), .Y(new_n6724));
  nand_5 g06348(.A(pi245), .B(pi140), .Y(new_n6725));
  xor_4  g06349(.A(new_n6725), .B(new_n6724), .Y(new_n6726));
  xor_4  g06350(.A(new_n6726), .B(new_n6723), .Y(new_n6727));
  nand_5 g06351(.A(pi171), .B(pi121), .Y(new_n6728));
  nand_5 g06352(.A(new_n6718), .B(new_n6717), .Y(new_n6729));
  nand_5 g06353(.A(new_n6719), .B(new_n6716), .Y(new_n6730));
  nand_5 g06354(.A(new_n6730), .B(new_n6729), .Y(new_n6731));
  xor_4  g06355(.A(new_n6731), .B(new_n6728), .Y(new_n6732));
  xor_4  g06356(.A(new_n6732), .B(new_n6727), .Y(new_n6733));
  nand_5 g06357(.A(pi231), .B(pi107), .Y(new_n6734));
  or_6   g06358(.A(new_n6714), .B(new_n6711), .Y(new_n6735));
  nand_5 g06359(.A(new_n6720), .B(new_n6715), .Y(new_n6736));
  nand_5 g06360(.A(new_n6736), .B(new_n6735), .Y(new_n6737));
  xor_4  g06361(.A(new_n6737), .B(new_n6734), .Y(new_n6738));
  xor_4  g06362(.A(new_n6738), .B(new_n6733), .Y(new_n6739));
  xnor_4 g06363(.A(new_n6739), .B(new_n6722), .Y(new_n6740));
  nand_5 g06364(.A(pi210), .B(pi039), .Y(new_n6741));
  nand_5 g06365(.A(pi228), .B(pi111), .Y(new_n6742));
  nand_5 g06366(.A(pi148), .B(pi024), .Y(new_n6743));
  xor_4  g06367(.A(new_n6743), .B(new_n6742), .Y(new_n6744));
  xor_4  g06368(.A(new_n6744), .B(new_n6741), .Y(new_n6745));
  nand_5 g06369(.A(new_n6544), .B(new_n6539), .Y(new_n6746));
  nand_5 g06370(.A(new_n6746), .B(new_n6543), .Y(new_n6747));
  nand_5 g06371(.A(pi224), .B(pi163), .Y(new_n6748));
  xor_4  g06372(.A(new_n6748), .B(new_n6747), .Y(new_n6749));
  xor_4  g06373(.A(new_n6749), .B(new_n6745), .Y(new_n6750));
  nor_5  g06374(.A(new_n6554), .B(new_n6546), .Y(new_n6751));
  not_8  g06375(.A(new_n6751), .Y(new_n6752));
  nor_5  g06376(.A(new_n6752), .B(new_n6750), .Y(new_n6753));
  nand_5 g06377(.A(pi210), .B(pi116), .Y(new_n6754));
  nand_5 g06378(.A(pi228), .B(pi024), .Y(new_n6755));
  nand_5 g06379(.A(pi111), .B(pi039), .Y(new_n6756));
  xor_4  g06380(.A(new_n6756), .B(new_n6755), .Y(new_n6757));
  xor_4  g06381(.A(new_n6757), .B(new_n6754), .Y(new_n6758));
  nand_5 g06382(.A(pi224), .B(pi148), .Y(new_n6759));
  nand_5 g06383(.A(new_n6743), .B(new_n6742), .Y(new_n6760));
  nand_5 g06384(.A(new_n6744), .B(new_n6741), .Y(new_n6761));
  nand_5 g06385(.A(new_n6761), .B(new_n6760), .Y(new_n6762));
  xor_4  g06386(.A(new_n6762), .B(new_n6759), .Y(new_n6763));
  xnor_4 g06387(.A(new_n6763), .B(new_n6758), .Y(new_n6764));
  nand_5 g06388(.A(pi255), .B(pi163), .Y(new_n6765));
  nand_5 g06389(.A(new_n6748), .B(new_n6747), .Y(new_n6766));
  nand_5 g06390(.A(new_n6749), .B(new_n6745), .Y(new_n6767));
  nand_5 g06391(.A(new_n6767), .B(new_n6766), .Y(new_n6768));
  xor_4  g06392(.A(new_n6768), .B(new_n6765), .Y(new_n6769));
  xnor_4 g06393(.A(new_n6769), .B(new_n6764), .Y(new_n6770));
  xor_4  g06394(.A(new_n6770), .B(new_n6753), .Y(new_n6771));
  xor_4  g06395(.A(new_n6721), .B(new_n6710), .Y(new_n6772));
  or_6   g06396(.A(new_n6548), .B(new_n6537), .Y(new_n6773));
  nand_5 g06397(.A(new_n6565), .B(new_n6549), .Y(new_n6774));
  nand_5 g06398(.A(new_n6774), .B(new_n6773), .Y(new_n6775));
  or_6   g06399(.A(new_n6775), .B(new_n6772), .Y(new_n6776));
  xor_4  g06400(.A(new_n6752), .B(new_n6750), .Y(new_n6777));
  not_8  g06401(.A(new_n6777), .Y(new_n6778));
  xor_4  g06402(.A(new_n6775), .B(new_n6772), .Y(new_n6779));
  nand_5 g06403(.A(new_n6779), .B(new_n6778), .Y(new_n6780));
  nand_5 g06404(.A(new_n6780), .B(new_n6776), .Y(new_n6781));
  xor_4  g06405(.A(new_n6781), .B(new_n6771), .Y(new_n6782));
  xnor_4 g06406(.A(new_n6782), .B(new_n6740), .Y(new_n6783));
  nand_5 g06407(.A(pi249), .B(pi149), .Y(new_n6784));
  nand_5 g06408(.A(pi240), .B(pi222), .Y(new_n6785));
  nand_5 g06409(.A(pi134), .B(pi125), .Y(new_n6786));
  xor_4  g06410(.A(new_n6786), .B(new_n6785), .Y(new_n6787));
  xnor_4 g06411(.A(new_n6787), .B(new_n6784), .Y(new_n6788));
  nand_5 g06412(.A(new_n6587), .B(new_n6582), .Y(new_n6789));
  nand_5 g06413(.A(new_n6789), .B(new_n6580), .Y(new_n6790));
  nand_5 g06414(.A(pi176), .B(pi175), .Y(new_n6791));
  xor_4  g06415(.A(new_n6791), .B(new_n6790), .Y(new_n6792));
  xor_4  g06416(.A(new_n6792), .B(new_n6788), .Y(new_n6793));
  not_8  g06417(.A(new_n6793), .Y(new_n6794));
  nand_5 g06418(.A(new_n6588), .B(new_n6583), .Y(new_n6795));
  nor_5  g06419(.A(new_n6795), .B(new_n6794), .Y(new_n6796));
  nand_5 g06420(.A(pi249), .B(pi167), .Y(new_n6797));
  nand_5 g06421(.A(pi240), .B(pi125), .Y(new_n6798));
  nand_5 g06422(.A(pi222), .B(pi149), .Y(new_n6799));
  xor_4  g06423(.A(new_n6799), .B(new_n6798), .Y(new_n6800));
  xor_4  g06424(.A(new_n6800), .B(new_n6797), .Y(new_n6801));
  nand_5 g06425(.A(pi176), .B(pi134), .Y(new_n6802));
  nand_5 g06426(.A(new_n6786), .B(new_n6785), .Y(new_n6803));
  nand_5 g06427(.A(new_n6787), .B(new_n6784), .Y(new_n6804));
  nand_5 g06428(.A(new_n6804), .B(new_n6803), .Y(new_n6805));
  xor_4  g06429(.A(new_n6805), .B(new_n6802), .Y(new_n6806));
  xor_4  g06430(.A(new_n6806), .B(new_n6801), .Y(new_n6807));
  nand_5 g06431(.A(pi175), .B(pi040), .Y(new_n6808));
  xor_4  g06432(.A(new_n6808), .B(new_n6807), .Y(new_n6809));
  or_6   g06433(.A(new_n6791), .B(new_n6790), .Y(new_n6810));
  nand_5 g06434(.A(new_n6792), .B(new_n6788), .Y(new_n6811));
  nand_5 g06435(.A(new_n6811), .B(new_n6810), .Y(new_n6812));
  xor_4  g06436(.A(new_n6812), .B(new_n6809), .Y(new_n6813));
  xor_4  g06437(.A(new_n6813), .B(new_n6796), .Y(new_n6814));
  nor_5  g06438(.A(new_n6814), .B(new_n6783), .Y(new_n6815));
  xor_4  g06439(.A(new_n6814), .B(new_n6783), .Y(new_n6816));
  not_8  g06440(.A(new_n6816), .Y(new_n6817));
  xor_4  g06441(.A(new_n6795), .B(new_n6793), .Y(new_n6818));
  nand_5 g06442(.A(new_n6589), .B(new_n6577), .Y(new_n6819));
  or_6   g06443(.A(new_n6591), .B(new_n6566), .Y(new_n6820));
  nand_5 g06444(.A(new_n6820), .B(new_n6819), .Y(new_n6821));
  or_6   g06445(.A(new_n6821), .B(new_n6818), .Y(new_n6822));
  xor_4  g06446(.A(new_n6779), .B(new_n6777), .Y(new_n6823));
  xor_4  g06447(.A(new_n6821), .B(new_n6818), .Y(new_n6824));
  nand_5 g06448(.A(new_n6824), .B(new_n6823), .Y(new_n6825));
  nand_5 g06449(.A(new_n6825), .B(new_n6822), .Y(new_n6826));
  nor_5  g06450(.A(new_n6826), .B(new_n6817), .Y(new_n6827));
  nor_5  g06451(.A(new_n6827), .B(new_n6815), .Y(new_n6828));
  nand_5 g06452(.A(pi149), .B(pi125), .Y(new_n6829));
  nand_5 g06453(.A(pi222), .B(pi167), .Y(new_n6830));
  nand_5 g06454(.A(pi249), .B(pi181), .Y(new_n6831));
  nand_5 g06455(.A(new_n6831), .B(new_n6830), .Y(new_n6832));
  nand_5 g06456(.A(pi222), .B(pi181), .Y(new_n6833));
  or_6   g06457(.A(new_n6833), .B(new_n6797), .Y(new_n6834));
  nand_5 g06458(.A(new_n6834), .B(new_n6832), .Y(new_n6835));
  xor_4  g06459(.A(new_n6835), .B(new_n6829), .Y(new_n6836));
  nand_5 g06460(.A(new_n6799), .B(new_n6798), .Y(new_n6837));
  nand_5 g06461(.A(new_n6800), .B(new_n6797), .Y(new_n6838));
  nand_5 g06462(.A(new_n6838), .B(new_n6837), .Y(new_n6839));
  xor_4  g06463(.A(new_n6839), .B(new_n6836), .Y(new_n6840));
  nand_5 g06464(.A(new_n6805), .B(new_n6802), .Y(new_n6841));
  nand_5 g06465(.A(new_n6806), .B(new_n6801), .Y(new_n6842));
  nand_5 g06466(.A(new_n6842), .B(new_n6841), .Y(new_n6843));
  nand_5 g06467(.A(pi240), .B(pi176), .Y(new_n6844));
  nand_5 g06468(.A(pi134), .B(pi040), .Y(new_n6845));
  nand_5 g06469(.A(new_n6845), .B(new_n6844), .Y(new_n6846));
  nand_5 g06470(.A(pi240), .B(pi040), .Y(new_n6847));
  or_6   g06471(.A(new_n6847), .B(new_n6802), .Y(new_n6848));
  nand_5 g06472(.A(new_n6848), .B(new_n6846), .Y(new_n6849));
  xor_4  g06473(.A(new_n6849), .B(new_n6843), .Y(new_n6850));
  xnor_4 g06474(.A(new_n6850), .B(new_n6840), .Y(new_n6851));
  or_6   g06475(.A(new_n6808), .B(new_n6807), .Y(new_n6852));
  nand_5 g06476(.A(new_n6812), .B(new_n6809), .Y(new_n6853));
  nand_5 g06477(.A(new_n6853), .B(new_n6852), .Y(new_n6854));
  xnor_4 g06478(.A(new_n6854), .B(new_n6851), .Y(new_n6855));
  nand_5 g06479(.A(new_n6813), .B(new_n6796), .Y(new_n6856));
  nand_5 g06480(.A(pi175), .B(pi174), .Y(new_n6857));
  xor_4  g06481(.A(new_n6857), .B(new_n6856), .Y(new_n6858));
  xnor_4 g06482(.A(new_n6858), .B(new_n6855), .Y(new_n6859));
  not_8  g06483(.A(new_n6753), .Y(new_n6860));
  nor_5  g06484(.A(new_n6770), .B(new_n6860), .Y(new_n6861));
  nand_5 g06485(.A(pi163), .B(pi127), .Y(new_n6862));
  nand_5 g06486(.A(pi039), .B(pi024), .Y(new_n6863));
  nand_5 g06487(.A(pi116), .B(pi111), .Y(new_n6864));
  nand_5 g06488(.A(pi210), .B(pi070), .Y(new_n6865));
  nand_5 g06489(.A(new_n6865), .B(new_n6864), .Y(new_n6866));
  nand_5 g06490(.A(pi111), .B(pi070), .Y(new_n6867));
  or_6   g06491(.A(new_n6867), .B(new_n6754), .Y(new_n6868));
  nand_5 g06492(.A(new_n6868), .B(new_n6866), .Y(new_n6869));
  xor_4  g06493(.A(new_n6869), .B(new_n6863), .Y(new_n6870));
  nand_5 g06494(.A(new_n6756), .B(new_n6755), .Y(new_n6871));
  nand_5 g06495(.A(new_n6757), .B(new_n6754), .Y(new_n6872));
  nand_5 g06496(.A(new_n6872), .B(new_n6871), .Y(new_n6873));
  xor_4  g06497(.A(new_n6873), .B(new_n6870), .Y(new_n6874));
  nand_5 g06498(.A(pi228), .B(pi224), .Y(new_n6875));
  nand_5 g06499(.A(pi255), .B(pi148), .Y(new_n6876));
  and_6  g06500(.A(new_n6876), .B(new_n6875), .Y(new_n6877));
  nand_5 g06501(.A(pi255), .B(pi228), .Y(new_n6878));
  nor_5  g06502(.A(new_n6878), .B(new_n6759), .Y(new_n6879));
  or_6   g06503(.A(new_n6879), .B(new_n6877), .Y(new_n6880));
  xnor_4 g06504(.A(new_n6880), .B(new_n6874), .Y(new_n6881));
  nand_5 g06505(.A(new_n6762), .B(new_n6759), .Y(new_n6882));
  nand_5 g06506(.A(new_n6763), .B(new_n6758), .Y(new_n6883));
  nand_5 g06507(.A(new_n6883), .B(new_n6882), .Y(new_n6884));
  xor_4  g06508(.A(new_n6884), .B(new_n6881), .Y(new_n6885));
  or_6   g06509(.A(new_n6768), .B(new_n6765), .Y(new_n6886));
  nand_5 g06510(.A(new_n6769), .B(new_n6764), .Y(new_n6887));
  nand_5 g06511(.A(new_n6887), .B(new_n6886), .Y(new_n6888));
  xnor_4 g06512(.A(new_n6888), .B(new_n6885), .Y(new_n6889));
  xor_4  g06513(.A(new_n6889), .B(new_n6862), .Y(new_n6890));
  xnor_4 g06514(.A(new_n6890), .B(new_n6861), .Y(new_n6891));
  nand_5 g06515(.A(new_n6739), .B(new_n6722), .Y(new_n6892));
  not_8  g06516(.A(new_n6892), .Y(new_n6893));
  nand_5 g06517(.A(pi107), .B(pi005), .Y(new_n6894));
  nand_5 g06518(.A(pi252), .B(pi245), .Y(new_n6895));
  nand_5 g06519(.A(new_n6725), .B(new_n6724), .Y(new_n6896));
  nand_5 g06520(.A(new_n6726), .B(new_n6723), .Y(new_n6897));
  nand_5 g06521(.A(new_n6897), .B(new_n6896), .Y(new_n6898));
  xor_4  g06522(.A(new_n6898), .B(new_n6895), .Y(new_n6899));
  nand_5 g06523(.A(pi201), .B(pi140), .Y(new_n6900));
  nand_5 g06524(.A(pi242), .B(pi156), .Y(new_n6901));
  nand_5 g06525(.A(new_n6901), .B(new_n6900), .Y(new_n6902));
  nand_5 g06526(.A(pi156), .B(pi140), .Y(new_n6903));
  nor_5  g06527(.A(new_n6903), .B(new_n6724), .Y(new_n6904));
  not_8  g06528(.A(new_n6904), .Y(new_n6905));
  nand_5 g06529(.A(new_n6905), .B(new_n6902), .Y(new_n6906));
  xor_4  g06530(.A(new_n6906), .B(new_n6899), .Y(new_n6907));
  nand_5 g06531(.A(pi231), .B(pi171), .Y(new_n6908));
  nand_5 g06532(.A(pi121), .B(pi049), .Y(new_n6909));
  and_6  g06533(.A(new_n6909), .B(new_n6908), .Y(new_n6910));
  nand_5 g06534(.A(pi231), .B(pi049), .Y(new_n6911));
  nor_5  g06535(.A(new_n6911), .B(new_n6728), .Y(new_n6912));
  or_6   g06536(.A(new_n6912), .B(new_n6910), .Y(new_n6913));
  xnor_4 g06537(.A(new_n6913), .B(new_n6907), .Y(new_n6914));
  nand_5 g06538(.A(new_n6731), .B(new_n6728), .Y(new_n6915));
  nand_5 g06539(.A(new_n6732), .B(new_n6727), .Y(new_n6916));
  nand_5 g06540(.A(new_n6916), .B(new_n6915), .Y(new_n6917));
  xor_4  g06541(.A(new_n6917), .B(new_n6914), .Y(new_n6918));
  not_8  g06542(.A(new_n6734), .Y(new_n6919));
  nand_5 g06543(.A(new_n6737), .B(new_n6919), .Y(new_n6920));
  or_6   g06544(.A(new_n6738), .B(new_n6733), .Y(new_n6921));
  nand_5 g06545(.A(new_n6921), .B(new_n6920), .Y(new_n6922));
  xnor_4 g06546(.A(new_n6922), .B(new_n6918), .Y(new_n6923));
  xor_4  g06547(.A(new_n6923), .B(new_n6894), .Y(new_n6924));
  xor_4  g06548(.A(new_n6924), .B(new_n6893), .Y(new_n6925));
  xor_4  g06549(.A(new_n6925), .B(new_n6891), .Y(new_n6926));
  nand_5 g06550(.A(new_n6781), .B(new_n6771), .Y(new_n6927));
  nand_5 g06551(.A(new_n6782), .B(new_n6740), .Y(new_n6928));
  nand_5 g06552(.A(new_n6928), .B(new_n6927), .Y(new_n6929));
  xor_4  g06553(.A(new_n6929), .B(new_n6926), .Y(new_n6930));
  xor_4  g06554(.A(new_n6930), .B(new_n6859), .Y(new_n6931));
  xor_4  g06555(.A(new_n6931), .B(new_n6828), .Y(new_n6932));
  not_8  g06556(.A(new_n6932), .Y(new_n6933));
  xor_4  g06557(.A(new_n6706), .B(new_n6705), .Y(new_n6934));
  or_6   g06558(.A(new_n6934), .B(new_n6933), .Y(new_n6935));
  xor_4  g06559(.A(new_n6934), .B(new_n6933), .Y(new_n6936));
  xor_4  g06560(.A(new_n6702), .B(new_n6700), .Y(new_n6937));
  xnor_4 g06561(.A(new_n6699), .B(new_n6698), .Y(new_n6938));
  or_6   g06562(.A(new_n6615), .B(new_n6604), .Y(new_n6939));
  nand_5 g06563(.A(new_n6616), .B(new_n6592), .Y(new_n6940));
  nand_5 g06564(.A(new_n6940), .B(new_n6939), .Y(new_n6941));
  nand_5 g06565(.A(new_n6941), .B(new_n6938), .Y(new_n6942));
  xor_4  g06566(.A(new_n6824), .B(new_n6823), .Y(new_n6943));
  not_8  g06567(.A(new_n6943), .Y(new_n6944));
  xor_4  g06568(.A(new_n6941), .B(new_n6938), .Y(new_n6945));
  nand_5 g06569(.A(new_n6945), .B(new_n6944), .Y(new_n6946));
  nand_5 g06570(.A(new_n6946), .B(new_n6942), .Y(new_n6947));
  or_6   g06571(.A(new_n6947), .B(new_n6937), .Y(new_n6948));
  xor_4  g06572(.A(new_n6826), .B(new_n6816), .Y(new_n6949));
  xor_4  g06573(.A(new_n6947), .B(new_n6937), .Y(new_n6950));
  nand_5 g06574(.A(new_n6950), .B(new_n6949), .Y(new_n6951));
  nand_5 g06575(.A(new_n6951), .B(new_n6948), .Y(new_n6952));
  nand_5 g06576(.A(new_n6952), .B(new_n6936), .Y(new_n6953));
  nand_5 g06577(.A(new_n6953), .B(new_n6935), .Y(new_n6954));
  or_6   g06578(.A(new_n6954), .B(new_n6709), .Y(new_n6955));
  not_8  g06579(.A(new_n6925), .Y(new_n6956));
  nor_5  g06580(.A(new_n6956), .B(new_n6891), .Y(new_n6957));
  nor_5  g06581(.A(new_n6929), .B(new_n6926), .Y(new_n6958));
  nor_5  g06582(.A(new_n6958), .B(new_n6957), .Y(new_n6959));
  nand_5 g06583(.A(new_n6888), .B(new_n6885), .Y(new_n6960));
  nand_5 g06584(.A(pi210), .B(pi115), .Y(new_n6961));
  nand_5 g06585(.A(pi116), .B(pi024), .Y(new_n6962));
  xor_4  g06586(.A(new_n6962), .B(new_n6961), .Y(new_n6963));
  xor_4  g06587(.A(new_n6963), .B(new_n6867), .Y(new_n6964));
  not_8  g06588(.A(new_n6964), .Y(new_n6965));
  nand_5 g06589(.A(pi224), .B(pi039), .Y(new_n6966));
  xor_4  g06590(.A(new_n6966), .B(new_n6868), .Y(new_n6967));
  xor_4  g06591(.A(new_n6967), .B(new_n6965), .Y(new_n6968));
  nand_5 g06592(.A(pi232), .B(pi163), .Y(new_n6969));
  nand_5 g06593(.A(pi148), .B(pi127), .Y(new_n6970));
  xor_4  g06594(.A(new_n6970), .B(new_n6969), .Y(new_n6971));
  xor_4  g06595(.A(new_n6971), .B(new_n6878), .Y(new_n6972));
  nand_5 g06596(.A(new_n6869), .B(new_n6863), .Y(new_n6973));
  nand_5 g06597(.A(new_n6873), .B(new_n6870), .Y(new_n6974));
  nand_5 g06598(.A(new_n6974), .B(new_n6973), .Y(new_n6975));
  xor_4  g06599(.A(new_n6975), .B(new_n6972), .Y(new_n6976));
  xor_4  g06600(.A(new_n6976), .B(new_n6968), .Y(new_n6977));
  nor_5  g06601(.A(new_n6884), .B(new_n6881), .Y(new_n6978));
  nand_5 g06602(.A(new_n6978), .B(new_n6879), .Y(new_n6979));
  nor_5  g06603(.A(new_n6880), .B(new_n6874), .Y(new_n6980));
  or_6   g06604(.A(new_n6980), .B(new_n6879), .Y(new_n6981));
  or_6   g06605(.A(new_n6981), .B(new_n6978), .Y(new_n6982));
  nand_5 g06606(.A(new_n6982), .B(new_n6979), .Y(new_n6983));
  xor_4  g06607(.A(new_n6983), .B(new_n6977), .Y(new_n6984));
  xor_4  g06608(.A(new_n6984), .B(new_n6960), .Y(new_n6985));
  or_6   g06609(.A(new_n6889), .B(new_n6862), .Y(new_n6986));
  nand_5 g06610(.A(new_n6890), .B(new_n6861), .Y(new_n6987));
  nand_5 g06611(.A(new_n6987), .B(new_n6986), .Y(new_n6988));
  xor_4  g06612(.A(new_n6988), .B(new_n6985), .Y(new_n6989));
  nand_5 g06613(.A(new_n6922), .B(new_n6918), .Y(new_n6990));
  nand_5 g06614(.A(pi242), .B(pi063), .Y(new_n6991));
  nand_5 g06615(.A(pi252), .B(pi201), .Y(new_n6992));
  xor_4  g06616(.A(new_n6992), .B(new_n6991), .Y(new_n6993));
  xor_4  g06617(.A(new_n6993), .B(new_n6903), .Y(new_n6994));
  nand_5 g06618(.A(pi245), .B(pi121), .Y(new_n6995));
  xor_4  g06619(.A(new_n6995), .B(new_n6905), .Y(new_n6996));
  not_8  g06620(.A(new_n6996), .Y(new_n6997));
  xor_4  g06621(.A(new_n6997), .B(new_n6994), .Y(new_n6998));
  nand_5 g06622(.A(pi107), .B(pi021), .Y(new_n6999));
  nand_5 g06623(.A(pi171), .B(pi005), .Y(new_n7000));
  xor_4  g06624(.A(new_n7000), .B(new_n6999), .Y(new_n7001));
  xor_4  g06625(.A(new_n7001), .B(new_n6911), .Y(new_n7002));
  nand_5 g06626(.A(new_n6898), .B(new_n6895), .Y(new_n7003));
  nand_5 g06627(.A(new_n6906), .B(new_n6899), .Y(new_n7004));
  nand_5 g06628(.A(new_n7004), .B(new_n7003), .Y(new_n7005));
  xor_4  g06629(.A(new_n7005), .B(new_n7002), .Y(new_n7006));
  xor_4  g06630(.A(new_n7006), .B(new_n6998), .Y(new_n7007));
  nor_5  g06631(.A(new_n6917), .B(new_n6914), .Y(new_n7008));
  nand_5 g06632(.A(new_n7008), .B(new_n6912), .Y(new_n7009));
  nor_5  g06633(.A(new_n6913), .B(new_n6907), .Y(new_n7010));
  or_6   g06634(.A(new_n7010), .B(new_n6912), .Y(new_n7011));
  or_6   g06635(.A(new_n7011), .B(new_n7008), .Y(new_n7012));
  nand_5 g06636(.A(new_n7012), .B(new_n7009), .Y(new_n7013));
  xor_4  g06637(.A(new_n7013), .B(new_n7007), .Y(new_n7014));
  xor_4  g06638(.A(new_n7014), .B(new_n6990), .Y(new_n7015));
  or_6   g06639(.A(new_n6923), .B(new_n6894), .Y(new_n7016));
  nand_5 g06640(.A(new_n6924), .B(new_n6893), .Y(new_n7017));
  nand_5 g06641(.A(new_n7017), .B(new_n7016), .Y(new_n7018));
  xor_4  g06642(.A(new_n7018), .B(new_n7015), .Y(new_n7019));
  xor_4  g06643(.A(new_n7019), .B(new_n6989), .Y(new_n7020));
  xnor_4 g06644(.A(new_n7020), .B(new_n6959), .Y(new_n7021));
  nand_5 g06645(.A(new_n6854), .B(new_n6851), .Y(new_n7022));
  nand_5 g06646(.A(pi249), .B(pi200), .Y(new_n7023));
  nand_5 g06647(.A(pi167), .B(pi125), .Y(new_n7024));
  xor_4  g06648(.A(new_n7024), .B(new_n7023), .Y(new_n7025));
  xor_4  g06649(.A(new_n7025), .B(new_n6833), .Y(new_n7026));
  not_8  g06650(.A(new_n7026), .Y(new_n7027));
  nand_5 g06651(.A(pi176), .B(pi149), .Y(new_n7028));
  xor_4  g06652(.A(new_n7028), .B(new_n6834), .Y(new_n7029));
  xor_4  g06653(.A(new_n7029), .B(new_n7027), .Y(new_n7030));
  nand_5 g06654(.A(pi175), .B(pi157), .Y(new_n7031));
  nand_5 g06655(.A(pi174), .B(pi134), .Y(new_n7032));
  xor_4  g06656(.A(new_n7032), .B(new_n7031), .Y(new_n7033));
  xor_4  g06657(.A(new_n7033), .B(new_n6847), .Y(new_n7034));
  nand_5 g06658(.A(new_n6835), .B(new_n6829), .Y(new_n7035));
  nand_5 g06659(.A(new_n6839), .B(new_n6836), .Y(new_n7036));
  nand_5 g06660(.A(new_n7036), .B(new_n7035), .Y(new_n7037));
  xor_4  g06661(.A(new_n7037), .B(new_n7034), .Y(new_n7038));
  xor_4  g06662(.A(new_n7038), .B(new_n7030), .Y(new_n7039));
  not_8  g06663(.A(new_n7039), .Y(new_n7040));
  nand_5 g06664(.A(new_n6849), .B(new_n6843), .Y(new_n7041));
  nand_5 g06665(.A(new_n6850), .B(new_n6840), .Y(new_n7042));
  nand_5 g06666(.A(new_n7042), .B(new_n7041), .Y(new_n7043));
  xor_4  g06667(.A(new_n7043), .B(new_n6848), .Y(new_n7044));
  xor_4  g06668(.A(new_n7044), .B(new_n7040), .Y(new_n7045));
  xnor_4 g06669(.A(new_n7045), .B(new_n7022), .Y(new_n7046));
  nand_5 g06670(.A(new_n6857), .B(new_n6856), .Y(new_n7047));
  nand_5 g06671(.A(new_n6858), .B(new_n6855), .Y(new_n7048));
  nand_5 g06672(.A(new_n7048), .B(new_n7047), .Y(new_n7049));
  xor_4  g06673(.A(new_n7049), .B(new_n7046), .Y(new_n7050));
  xor_4  g06674(.A(new_n7050), .B(new_n7021), .Y(new_n7051));
  nand_5 g06675(.A(new_n6930), .B(new_n6859), .Y(new_n7052));
  nand_5 g06676(.A(new_n6931), .B(new_n6828), .Y(new_n7053));
  nand_5 g06677(.A(new_n7053), .B(new_n7052), .Y(new_n7054));
  xor_4  g06678(.A(new_n7054), .B(new_n7051), .Y(new_n7055));
  not_8  g06679(.A(new_n7055), .Y(new_n7056));
  xor_4  g06680(.A(new_n6954), .B(new_n6709), .Y(new_n7057));
  nand_5 g06681(.A(new_n7057), .B(new_n7056), .Y(new_n7058));
  nand_5 g06682(.A(new_n7058), .B(new_n6955), .Y(new_n7059));
  nand_5 g06683(.A(pi171), .B(pi021), .Y(new_n7060));
  nand_5 g06684(.A(new_n6992), .B(new_n6991), .Y(new_n7061));
  nand_5 g06685(.A(new_n6993), .B(new_n6903), .Y(new_n7062));
  nand_5 g06686(.A(new_n7062), .B(new_n7061), .Y(new_n7063));
  xor_4  g06687(.A(new_n7063), .B(new_n7060), .Y(new_n7064));
  nor_5  g06688(.A(new_n6694), .B(new_n6688), .Y(new_n7065));
  nor_5  g06689(.A(new_n7065), .B(new_n6693), .Y(new_n7066));
  nand_5 g06690(.A(pi255), .B(pi039), .Y(new_n7067));
  nand_5 g06691(.A(new_n6970), .B(new_n6969), .Y(new_n7068));
  nand_5 g06692(.A(new_n6971), .B(new_n6878), .Y(new_n7069));
  nand_5 g06693(.A(new_n7069), .B(new_n7068), .Y(new_n7070));
  xor_4  g06694(.A(new_n7070), .B(new_n7067), .Y(new_n7071));
  or_6   g06695(.A(new_n7013), .B(new_n7007), .Y(new_n7072));
  nand_5 g06696(.A(new_n7072), .B(new_n7012), .Y(new_n7073));
  nand_5 g06697(.A(pi201), .B(pi121), .Y(new_n7074));
  nand_5 g06698(.A(pi245), .B(pi231), .Y(new_n7075));
  xor_4  g06699(.A(new_n7075), .B(new_n7074), .Y(new_n7076));
  xor_4  g06700(.A(new_n7076), .B(new_n7073), .Y(new_n7077));
  xor_4  g06701(.A(new_n7077), .B(new_n7071), .Y(new_n7078));
  xor_4  g06702(.A(new_n7078), .B(new_n7066), .Y(new_n7079));
  xor_4  g06703(.A(new_n7079), .B(new_n7064), .Y(new_n7080));
  xor_4  g06704(.A(new_n7080), .B(new_n7059), .Y(new_n7081));
  or_6   g06705(.A(new_n7014), .B(new_n6990), .Y(new_n7082));
  nand_5 g06706(.A(new_n7018), .B(new_n7015), .Y(new_n7083));
  nand_5 g06707(.A(new_n7083), .B(new_n7082), .Y(new_n7084));
  nor_5  g06708(.A(new_n6695), .B(new_n6672), .Y(new_n7085));
  nor_5  g06709(.A(new_n6708), .B(new_n6696), .Y(new_n7086));
  or_6   g06710(.A(new_n7086), .B(new_n7085), .Y(new_n7087));
  xor_4  g06711(.A(new_n7087), .B(new_n7084), .Y(new_n7088));
  nor_5  g06712(.A(new_n6995), .B(new_n6905), .Y(new_n7089));
  nor_5  g06713(.A(new_n6997), .B(new_n6994), .Y(new_n7090));
  or_6   g06714(.A(new_n7090), .B(new_n7089), .Y(new_n7091));
  xor_4  g06715(.A(new_n7091), .B(new_n7088), .Y(new_n7092));
  nand_5 g06716(.A(pi181), .B(pi125), .Y(new_n7093));
  nand_5 g06717(.A(pi210), .B(pi000), .Y(new_n7094));
  nand_5 g06718(.A(pi070), .B(pi024), .Y(new_n7095));
  nand_5 g06719(.A(pi115), .B(pi111), .Y(new_n7096));
  xor_4  g06720(.A(new_n7096), .B(new_n7095), .Y(new_n7097));
  nand_5 g06721(.A(pi191), .B(pi163), .Y(new_n7098));
  or_6   g06722(.A(new_n7019), .B(new_n6989), .Y(new_n7099));
  nand_5 g06723(.A(new_n7020), .B(new_n6959), .Y(new_n7100));
  nand_5 g06724(.A(new_n7100), .B(new_n7099), .Y(new_n7101));
  xor_4  g06725(.A(new_n7101), .B(new_n7098), .Y(new_n7102));
  xor_4  g06726(.A(new_n7102), .B(new_n7097), .Y(new_n7103));
  xor_4  g06727(.A(new_n7103), .B(new_n7094), .Y(new_n7104));
  xor_4  g06728(.A(new_n7104), .B(new_n7093), .Y(new_n7105));
  nand_5 g06729(.A(pi176), .B(pi167), .Y(new_n7106));
  or_6   g06730(.A(new_n7028), .B(new_n6834), .Y(new_n7107));
  nand_5 g06731(.A(new_n7029), .B(new_n7027), .Y(new_n7108));
  nand_5 g06732(.A(new_n7108), .B(new_n7107), .Y(new_n7109));
  xor_4  g06733(.A(new_n7109), .B(new_n7106), .Y(new_n7110));
  or_6   g06734(.A(new_n6984), .B(new_n6960), .Y(new_n7111));
  nand_5 g06735(.A(new_n6988), .B(new_n6985), .Y(new_n7112));
  nand_5 g06736(.A(new_n7112), .B(new_n7111), .Y(new_n7113));
  nand_5 g06737(.A(pi157), .B(pi134), .Y(new_n7114));
  nand_5 g06738(.A(new_n7024), .B(new_n7023), .Y(new_n7115));
  nand_5 g06739(.A(new_n7025), .B(new_n6833), .Y(new_n7116));
  nand_5 g06740(.A(new_n7116), .B(new_n7115), .Y(new_n7117));
  or_6   g06741(.A(new_n7037), .B(new_n7034), .Y(new_n7118));
  nand_5 g06742(.A(new_n7038), .B(new_n7030), .Y(new_n7119));
  nand_5 g06743(.A(new_n7119), .B(new_n7118), .Y(new_n7120));
  xor_4  g06744(.A(new_n7120), .B(new_n7117), .Y(new_n7121));
  xor_4  g06745(.A(new_n7121), .B(new_n7114), .Y(new_n7122));
  xor_4  g06746(.A(new_n7122), .B(new_n7113), .Y(new_n7123));
  xor_4  g06747(.A(new_n7123), .B(new_n7110), .Y(new_n7124));
  or_6   g06748(.A(new_n6983), .B(new_n6977), .Y(new_n7125));
  nand_5 g06749(.A(new_n7125), .B(new_n6982), .Y(new_n7126));
  nand_5 g06750(.A(new_n7032), .B(new_n7031), .Y(new_n7127));
  nand_5 g06751(.A(new_n7033), .B(new_n6847), .Y(new_n7128));
  nand_5 g06752(.A(new_n7128), .B(new_n7127), .Y(new_n7129));
  xor_4  g06753(.A(new_n7129), .B(new_n7126), .Y(new_n7130));
  nand_5 g06754(.A(pi149), .B(pi040), .Y(new_n7131));
  nand_5 g06755(.A(pi240), .B(pi174), .Y(new_n7132));
  xor_4  g06756(.A(new_n7132), .B(new_n7131), .Y(new_n7133));
  xor_4  g06757(.A(new_n7133), .B(new_n7130), .Y(new_n7134));
  xor_4  g06758(.A(new_n7134), .B(new_n7124), .Y(new_n7135));
  xor_4  g06759(.A(new_n7135), .B(new_n7105), .Y(new_n7136));
  nand_5 g06760(.A(pi187), .B(pi117), .Y(new_n7137));
  nand_5 g06761(.A(pi214), .B(pi100), .Y(new_n7138));
  xor_4  g06762(.A(new_n7138), .B(new_n7137), .Y(new_n7139));
  xor_4  g06763(.A(new_n7139), .B(new_n7136), .Y(new_n7140));
  nand_5 g06764(.A(new_n6674), .B(new_n6673), .Y(new_n7141));
  nand_5 g06765(.A(new_n6675), .B(new_n6625), .Y(new_n7142));
  nand_5 g06766(.A(new_n7142), .B(new_n7141), .Y(new_n7143));
  nand_5 g06767(.A(pi247), .B(pi081), .Y(new_n7144));
  nand_5 g06768(.A(pi106), .B(pi080), .Y(new_n7145));
  xor_4  g06769(.A(new_n7145), .B(new_n7144), .Y(new_n7146));
  xor_4  g06770(.A(new_n7146), .B(new_n7143), .Y(new_n7147));
  nand_5 g06771(.A(pi233), .B(pi016), .Y(new_n7148));
  nor_5  g06772(.A(new_n7045), .B(new_n7022), .Y(new_n7149));
  nor_5  g06773(.A(new_n7049), .B(new_n7046), .Y(new_n7150));
  or_6   g06774(.A(new_n7150), .B(new_n7149), .Y(new_n7151));
  nand_5 g06775(.A(pi249), .B(pi203), .Y(new_n7152));
  xor_4  g06776(.A(new_n7152), .B(new_n7151), .Y(new_n7153));
  nand_5 g06777(.A(new_n7043), .B(new_n6848), .Y(new_n7154));
  nand_5 g06778(.A(new_n7044), .B(new_n7040), .Y(new_n7155));
  nand_5 g06779(.A(new_n7155), .B(new_n7154), .Y(new_n7156));
  nand_5 g06780(.A(new_n6686), .B(new_n6683), .Y(new_n7157));
  nand_5 g06781(.A(new_n6687), .B(new_n6679), .Y(new_n7158));
  nand_5 g06782(.A(new_n7158), .B(new_n7157), .Y(new_n7159));
  nand_5 g06783(.A(new_n6681), .B(new_n6680), .Y(new_n7160));
  nand_5 g06784(.A(new_n6682), .B(new_n6639), .Y(new_n7161));
  nand_5 g06785(.A(new_n7161), .B(new_n7160), .Y(new_n7162));
  nand_5 g06786(.A(pi222), .B(pi200), .Y(new_n7163));
  nand_5 g06787(.A(pi175), .B(pi017), .Y(new_n7164));
  xor_4  g06788(.A(new_n7164), .B(new_n7163), .Y(new_n7165));
  xor_4  g06789(.A(new_n7165), .B(new_n7162), .Y(new_n7166));
  xor_4  g06790(.A(new_n7166), .B(new_n7159), .Y(new_n7167));
  xor_4  g06791(.A(new_n7167), .B(new_n7156), .Y(new_n7168));
  xor_4  g06792(.A(new_n7168), .B(new_n7153), .Y(new_n7169));
  xor_4  g06793(.A(new_n7169), .B(new_n7148), .Y(new_n7170));
  xor_4  g06794(.A(new_n7170), .B(new_n7147), .Y(new_n7171));
  or_6   g06795(.A(new_n6677), .B(new_n6626), .Y(new_n7172));
  not_8  g06796(.A(new_n6676), .Y(new_n7173));
  nand_5 g06797(.A(new_n6678), .B(new_n7173), .Y(new_n7174));
  nand_5 g06798(.A(new_n7174), .B(new_n7172), .Y(new_n7175));
  nand_5 g06799(.A(pi234), .B(pi227), .Y(new_n7176));
  xor_4  g06800(.A(new_n7176), .B(new_n7175), .Y(new_n7177));
  xor_4  g06801(.A(new_n7177), .B(new_n7171), .Y(new_n7178));
  xor_4  g06802(.A(new_n7178), .B(new_n7140), .Y(new_n7179));
  nand_5 g06803(.A(new_n7000), .B(new_n6999), .Y(new_n7180));
  nand_5 g06804(.A(new_n7001), .B(new_n6911), .Y(new_n7181));
  nand_5 g06805(.A(new_n7181), .B(new_n7180), .Y(new_n7182));
  or_6   g06806(.A(new_n7005), .B(new_n7002), .Y(new_n7183));
  nand_5 g06807(.A(new_n7006), .B(new_n6998), .Y(new_n7184));
  nand_5 g06808(.A(new_n7184), .B(new_n7183), .Y(new_n7185));
  xor_4  g06809(.A(new_n7185), .B(new_n7182), .Y(new_n7186));
  nand_5 g06810(.A(pi049), .B(pi005), .Y(new_n7187));
  xor_4  g06811(.A(new_n7187), .B(new_n7186), .Y(new_n7188));
  xor_4  g06812(.A(new_n7188), .B(new_n7179), .Y(new_n7189));
  xor_4  g06813(.A(new_n7189), .B(new_n7092), .Y(new_n7190));
  nand_5 g06814(.A(new_n7050), .B(new_n7021), .Y(new_n7191));
  nand_5 g06815(.A(new_n7054), .B(new_n7051), .Y(new_n7192));
  nand_5 g06816(.A(new_n7192), .B(new_n7191), .Y(new_n7193));
  nand_5 g06817(.A(pi217), .B(pi202), .Y(new_n7194));
  nand_5 g06818(.A(pi129), .B(pi103), .Y(new_n7195));
  xor_4  g06819(.A(new_n7195), .B(new_n7194), .Y(new_n7196));
  or_6   g06820(.A(new_n6975), .B(new_n6972), .Y(new_n7197));
  nand_5 g06821(.A(new_n6976), .B(new_n6968), .Y(new_n7198));
  nand_5 g06822(.A(new_n7198), .B(new_n7197), .Y(new_n7199));
  xor_4  g06823(.A(new_n7199), .B(new_n7196), .Y(new_n7200));
  nand_5 g06824(.A(pi224), .B(pi116), .Y(new_n7201));
  or_6   g06825(.A(new_n6966), .B(new_n6868), .Y(new_n7202));
  nand_5 g06826(.A(new_n6967), .B(new_n6965), .Y(new_n7203));
  nand_5 g06827(.A(new_n7203), .B(new_n7202), .Y(new_n7204));
  nand_5 g06828(.A(new_n6962), .B(new_n6961), .Y(new_n7205));
  nand_5 g06829(.A(new_n6963), .B(new_n6867), .Y(new_n7206));
  nand_5 g06830(.A(new_n7206), .B(new_n7205), .Y(new_n7207));
  xor_4  g06831(.A(new_n7207), .B(new_n7204), .Y(new_n7208));
  nand_5 g06832(.A(pi232), .B(pi148), .Y(new_n7209));
  nand_5 g06833(.A(pi228), .B(pi127), .Y(new_n7210));
  xor_4  g06834(.A(new_n7210), .B(new_n7209), .Y(new_n7211));
  xor_4  g06835(.A(new_n7211), .B(new_n7208), .Y(new_n7212));
  xor_4  g06836(.A(new_n7212), .B(new_n7201), .Y(new_n7213));
  nand_5 g06837(.A(pi140), .B(pi063), .Y(new_n7214));
  nand_5 g06838(.A(pi107), .B(pi082), .Y(new_n7215));
  nand_5 g06839(.A(pi252), .B(pi156), .Y(new_n7216));
  nand_5 g06840(.A(pi242), .B(pi083), .Y(new_n7217));
  xor_4  g06841(.A(new_n7217), .B(new_n7216), .Y(new_n7218));
  xor_4  g06842(.A(new_n7218), .B(new_n7215), .Y(new_n7219));
  xor_4  g06843(.A(new_n7219), .B(new_n7214), .Y(new_n7220));
  xor_4  g06844(.A(new_n7220), .B(new_n7213), .Y(new_n7221));
  xor_4  g06845(.A(new_n7221), .B(new_n7200), .Y(new_n7222));
  xor_4  g06846(.A(new_n7222), .B(new_n7193), .Y(new_n7223));
  xor_4  g06847(.A(new_n7223), .B(new_n7190), .Y(new_n7224));
  xor_4  g06848(.A(new_n7224), .B(new_n7081), .Y(po036));
  xor_4  g06849(.A(new_n6952), .B(new_n6936), .Y(po037));
  xnor_4 g06850(.A(new_n3260), .B(new_n3259), .Y(po038));
  nand_5 g06851(.A(pi145), .B(pi013), .Y(new_n7228));
  nand_5 g06852(.A(pi164), .B(pi112), .Y(new_n7229));
  nand_5 g06853(.A(pi206), .B(pi105), .Y(new_n7230));
  or_6   g06854(.A(new_n7230), .B(new_n7229), .Y(new_n7231));
  or_6   g06855(.A(new_n7231), .B(new_n7228), .Y(new_n7232));
  nand_5 g06856(.A(pi183), .B(pi164), .Y(new_n7233));
  nand_5 g06857(.A(pi112), .B(pi032), .Y(new_n7234));
  xor_4  g06858(.A(new_n7234), .B(new_n7233), .Y(new_n7235));
  xor_4  g06859(.A(new_n7235), .B(new_n7230), .Y(new_n7236));
  not_8  g06860(.A(new_n7236), .Y(new_n7237));
  xor_4  g06861(.A(new_n7231), .B(new_n7228), .Y(new_n7238));
  nand_5 g06862(.A(new_n7238), .B(new_n7237), .Y(new_n7239));
  nand_5 g06863(.A(new_n7239), .B(new_n7232), .Y(new_n7240));
  nand_5 g06864(.A(pi077), .B(pi054), .Y(new_n7241));
  nand_5 g06865(.A(pi052), .B(pi044), .Y(new_n7242));
  nor_5  g06866(.A(new_n7242), .B(new_n7241), .Y(new_n7243));
  nand_5 g06867(.A(pi250), .B(pi133), .Y(new_n7244));
  nand_5 g06868(.A(pi189), .B(pi045), .Y(new_n7245));
  nand_5 g06869(.A(pi119), .B(pi064), .Y(new_n7246));
  nand_5 g06870(.A(new_n7246), .B(new_n7245), .Y(new_n7247));
  nand_5 g06871(.A(pi189), .B(pi119), .Y(new_n7248));
  nand_5 g06872(.A(pi064), .B(pi045), .Y(new_n7249));
  or_6   g06873(.A(new_n7249), .B(new_n7248), .Y(new_n7250));
  nand_5 g06874(.A(new_n7250), .B(new_n7247), .Y(new_n7251));
  xor_4  g06875(.A(new_n7251), .B(new_n7244), .Y(new_n7252));
  nand_5 g06876(.A(pi250), .B(pi077), .Y(new_n7253));
  nand_5 g06877(.A(new_n7253), .B(new_n7248), .Y(new_n7254));
  nand_5 g06878(.A(pi133), .B(pi045), .Y(new_n7255));
  xor_4  g06879(.A(new_n7253), .B(new_n7248), .Y(new_n7256));
  nand_5 g06880(.A(new_n7256), .B(new_n7255), .Y(new_n7257));
  nand_5 g06881(.A(new_n7257), .B(new_n7254), .Y(new_n7258));
  xor_4  g06882(.A(new_n7258), .B(new_n7252), .Y(new_n7259));
  nand_5 g06883(.A(pi077), .B(pi044), .Y(new_n7260));
  nand_5 g06884(.A(pi054), .B(pi052), .Y(new_n7261));
  and_6  g06885(.A(new_n7261), .B(new_n7260), .Y(new_n7262));
  or_6   g06886(.A(new_n7262), .B(new_n7243), .Y(new_n7263));
  xnor_4 g06887(.A(new_n7263), .B(new_n7259), .Y(new_n7264));
  nand_5 g06888(.A(pi133), .B(pi119), .Y(new_n7265));
  nand_5 g06889(.A(pi077), .B(pi045), .Y(new_n7266));
  nand_5 g06890(.A(new_n7266), .B(new_n7265), .Y(new_n7267));
  nand_5 g06891(.A(pi250), .B(pi052), .Y(new_n7268));
  xor_4  g06892(.A(new_n7266), .B(new_n7265), .Y(new_n7269));
  nand_5 g06893(.A(new_n7269), .B(new_n7268), .Y(new_n7270));
  nand_5 g06894(.A(new_n7270), .B(new_n7267), .Y(new_n7271));
  nand_5 g06895(.A(new_n7271), .B(new_n7242), .Y(new_n7272));
  xor_4  g06896(.A(new_n7256), .B(new_n7255), .Y(new_n7273));
  xor_4  g06897(.A(new_n7271), .B(new_n7242), .Y(new_n7274));
  nand_5 g06898(.A(new_n7274), .B(new_n7273), .Y(new_n7275));
  nand_5 g06899(.A(new_n7275), .B(new_n7272), .Y(new_n7276));
  nor_5  g06900(.A(new_n7276), .B(new_n7264), .Y(new_n7277));
  nand_5 g06901(.A(new_n7277), .B(new_n7243), .Y(new_n7278));
  nand_5 g06902(.A(pi250), .B(pi189), .Y(new_n7279));
  nand_5 g06903(.A(pi119), .B(pi084), .Y(new_n7280));
  xor_4  g06904(.A(new_n7280), .B(new_n7279), .Y(new_n7281));
  xor_4  g06905(.A(new_n7281), .B(new_n7249), .Y(new_n7282));
  nand_5 g06906(.A(pi133), .B(pi044), .Y(new_n7283));
  xor_4  g06907(.A(new_n7283), .B(new_n7250), .Y(new_n7284));
  xor_4  g06908(.A(new_n7284), .B(new_n7282), .Y(new_n7285));
  nand_5 g06909(.A(pi072), .B(pi052), .Y(new_n7286));
  nand_5 g06910(.A(pi248), .B(pi131), .Y(new_n7287));
  xor_4  g06911(.A(new_n7287), .B(new_n7286), .Y(new_n7288));
  xor_4  g06912(.A(new_n7288), .B(new_n7241), .Y(new_n7289));
  nand_5 g06913(.A(new_n7251), .B(new_n7244), .Y(new_n7290));
  nand_5 g06914(.A(new_n7258), .B(new_n7252), .Y(new_n7291));
  nand_5 g06915(.A(new_n7291), .B(new_n7290), .Y(new_n7292));
  xor_4  g06916(.A(new_n7292), .B(new_n7289), .Y(new_n7293));
  xnor_4 g06917(.A(new_n7293), .B(new_n7285), .Y(new_n7294));
  nor_5  g06918(.A(new_n7263), .B(new_n7259), .Y(new_n7295));
  xor_4  g06919(.A(new_n7277), .B(new_n7243), .Y(new_n7296));
  nor_5  g06920(.A(new_n7296), .B(new_n7295), .Y(new_n7297));
  not_8  g06921(.A(new_n7297), .Y(new_n7298));
  nand_5 g06922(.A(new_n7298), .B(new_n7294), .Y(new_n7299));
  nand_5 g06923(.A(new_n7299), .B(new_n7278), .Y(new_n7300));
  nand_5 g06924(.A(pi241), .B(pi235), .Y(new_n7301));
  xor_4  g06925(.A(new_n7276), .B(new_n7264), .Y(new_n7302));
  nand_5 g06926(.A(pi131), .B(pi054), .Y(new_n7303));
  nand_5 g06927(.A(pi131), .B(pi044), .Y(new_n7304));
  nand_5 g06928(.A(pi250), .B(pi131), .Y(new_n7305));
  nand_5 g06929(.A(pi052), .B(pi045), .Y(new_n7306));
  nand_5 g06930(.A(new_n7306), .B(new_n7305), .Y(new_n7307));
  nand_5 g06931(.A(pi119), .B(pi077), .Y(new_n7308));
  xor_4  g06932(.A(new_n7306), .B(new_n7305), .Y(new_n7309));
  nand_5 g06933(.A(new_n7309), .B(new_n7308), .Y(new_n7310));
  nand_5 g06934(.A(new_n7310), .B(new_n7307), .Y(new_n7311));
  nand_5 g06935(.A(new_n7311), .B(new_n7304), .Y(new_n7312));
  xor_4  g06936(.A(new_n7269), .B(new_n7268), .Y(new_n7313));
  xor_4  g06937(.A(new_n7311), .B(new_n7304), .Y(new_n7314));
  nand_5 g06938(.A(new_n7314), .B(new_n7313), .Y(new_n7315));
  nand_5 g06939(.A(new_n7315), .B(new_n7312), .Y(new_n7316));
  or_6   g06940(.A(new_n7316), .B(new_n7303), .Y(new_n7317));
  xor_4  g06941(.A(new_n7316), .B(new_n7303), .Y(new_n7318));
  xnor_4 g06942(.A(new_n7274), .B(new_n7273), .Y(new_n7319));
  nand_5 g06943(.A(new_n7319), .B(new_n7318), .Y(new_n7320));
  nand_5 g06944(.A(new_n7320), .B(new_n7317), .Y(new_n7321));
  xor_4  g06945(.A(new_n7321), .B(new_n7302), .Y(new_n7322));
  nand_5 g06946(.A(pi131), .B(pi072), .Y(new_n7323));
  xor_4  g06947(.A(new_n7309), .B(new_n7308), .Y(new_n7324));
  nand_5 g06948(.A(pi131), .B(pi045), .Y(new_n7325));
  nand_5 g06949(.A(pi119), .B(pi052), .Y(new_n7326));
  nor_5  g06950(.A(new_n7326), .B(new_n7325), .Y(new_n7327));
  not_8  g06951(.A(new_n7327), .Y(new_n7328));
  or_6   g06952(.A(new_n7328), .B(new_n7324), .Y(new_n7329));
  xor_4  g06953(.A(new_n7314), .B(new_n7313), .Y(new_n7330));
  nor_5  g06954(.A(new_n7330), .B(new_n7329), .Y(new_n7331));
  xor_4  g06955(.A(new_n7319), .B(new_n7318), .Y(new_n7332));
  nand_5 g06956(.A(new_n7332), .B(new_n7331), .Y(new_n7333));
  xor_4  g06957(.A(new_n7333), .B(new_n7323), .Y(new_n7334));
  xor_4  g06958(.A(new_n7334), .B(new_n7322), .Y(new_n7335));
  xor_4  g06959(.A(new_n7332), .B(new_n7331), .Y(new_n7336));
  not_8  g06960(.A(new_n7336), .Y(new_n7337));
  nand_5 g06961(.A(pi164), .B(pi104), .Y(new_n7338));
  nand_5 g06962(.A(pi212), .B(pi206), .Y(new_n7339));
  nand_5 g06963(.A(pi213), .B(pi032), .Y(new_n7340));
  xor_4  g06964(.A(new_n7340), .B(new_n7339), .Y(new_n7341));
  xor_4  g06965(.A(new_n7341), .B(new_n7338), .Y(new_n7342));
  or_6   g06966(.A(new_n7339), .B(new_n378), .Y(new_n7343));
  or_6   g06967(.A(new_n7343), .B(new_n7342), .Y(new_n7344));
  nand_5 g06968(.A(pi212), .B(pi032), .Y(new_n7345));
  nand_5 g06969(.A(pi206), .B(pi104), .Y(new_n7346));
  nand_5 g06970(.A(pi164), .B(pi013), .Y(new_n7347));
  xor_4  g06971(.A(new_n7347), .B(new_n7346), .Y(new_n7348));
  xor_4  g06972(.A(new_n7348), .B(new_n7345), .Y(new_n7349));
  nand_5 g06973(.A(pi213), .B(pi145), .Y(new_n7350));
  nand_5 g06974(.A(new_n7340), .B(new_n7339), .Y(new_n7351));
  nand_5 g06975(.A(new_n7341), .B(new_n7338), .Y(new_n7352));
  nand_5 g06976(.A(new_n7352), .B(new_n7351), .Y(new_n7353));
  xor_4  g06977(.A(new_n7353), .B(new_n7350), .Y(new_n7354));
  xor_4  g06978(.A(new_n7354), .B(new_n7349), .Y(new_n7355));
  nor_5  g06979(.A(new_n7355), .B(new_n7344), .Y(new_n7356));
  nand_5 g06980(.A(pi104), .B(pi032), .Y(new_n7357));
  nand_5 g06981(.A(pi206), .B(pi013), .Y(new_n7358));
  xor_4  g06982(.A(new_n7358), .B(new_n7357), .Y(new_n7359));
  xor_4  g06983(.A(new_n7359), .B(new_n7229), .Y(new_n7360));
  nand_5 g06984(.A(pi212), .B(pi145), .Y(new_n7361));
  nand_5 g06985(.A(new_n7347), .B(new_n7346), .Y(new_n7362));
  nand_5 g06986(.A(new_n7348), .B(new_n7345), .Y(new_n7363));
  nand_5 g06987(.A(new_n7363), .B(new_n7362), .Y(new_n7364));
  xor_4  g06988(.A(new_n7364), .B(new_n7361), .Y(new_n7365));
  xor_4  g06989(.A(new_n7365), .B(new_n7360), .Y(new_n7366));
  nand_5 g06990(.A(pi246), .B(pi213), .Y(new_n7367));
  xnor_4 g06991(.A(new_n7367), .B(new_n7366), .Y(new_n7368));
  nand_5 g06992(.A(new_n7353), .B(new_n7350), .Y(new_n7369));
  nand_5 g06993(.A(new_n7354), .B(new_n7349), .Y(new_n7370));
  nand_5 g06994(.A(new_n7370), .B(new_n7369), .Y(new_n7371));
  xor_4  g06995(.A(new_n7371), .B(new_n7368), .Y(new_n7372));
  xnor_4 g06996(.A(new_n7372), .B(new_n7356), .Y(new_n7373));
  nand_5 g06997(.A(pi161), .B(pi027), .Y(new_n7374));
  nand_5 g06998(.A(pi236), .B(pi008), .Y(new_n7375));
  nand_5 g06999(.A(new_n7375), .B(new_n7374), .Y(new_n7376));
  nand_5 g07000(.A(pi241), .B(pi026), .Y(new_n7377));
  or_6   g07001(.A(new_n7375), .B(new_n7374), .Y(new_n7378));
  nand_5 g07002(.A(new_n7378), .B(new_n7377), .Y(new_n7379));
  nand_5 g07003(.A(new_n7379), .B(new_n7376), .Y(new_n7380));
  nand_5 g07004(.A(pi236), .B(pi056), .Y(new_n7381));
  xor_4  g07005(.A(new_n7381), .B(new_n7380), .Y(new_n7382));
  nand_5 g07006(.A(pi161), .B(pi026), .Y(new_n7383));
  nand_5 g07007(.A(pi141), .B(pi027), .Y(new_n7384));
  nand_5 g07008(.A(pi241), .B(pi008), .Y(new_n7385));
  xor_4  g07009(.A(new_n7385), .B(new_n7384), .Y(new_n7386));
  xor_4  g07010(.A(new_n7386), .B(new_n7383), .Y(new_n7387));
  xor_4  g07011(.A(new_n7387), .B(new_n7382), .Y(new_n7388));
  not_8  g07012(.A(new_n7377), .Y(new_n7389));
  not_8  g07013(.A(new_n7376), .Y(new_n7390));
  nand_5 g07014(.A(new_n7389), .B(new_n377), .Y(new_n7391));
  nand_5 g07015(.A(new_n7391), .B(new_n7390), .Y(new_n7392));
  nand_5 g07016(.A(new_n7392), .B(new_n7378), .Y(new_n7393));
  nand_5 g07017(.A(new_n7393), .B(new_n7389), .Y(new_n7394));
  nor_5  g07018(.A(new_n7394), .B(new_n7388), .Y(new_n7395));
  nand_5 g07019(.A(pi161), .B(pi008), .Y(new_n7396));
  nand_5 g07020(.A(pi090), .B(pi027), .Y(new_n7397));
  nand_5 g07021(.A(pi141), .B(pi026), .Y(new_n7398));
  xor_4  g07022(.A(new_n7398), .B(new_n7397), .Y(new_n7399));
  xor_4  g07023(.A(new_n7399), .B(new_n7396), .Y(new_n7400));
  nand_5 g07024(.A(pi241), .B(pi056), .Y(new_n7401));
  nand_5 g07025(.A(new_n7385), .B(new_n7384), .Y(new_n7402));
  nand_5 g07026(.A(new_n7386), .B(new_n7383), .Y(new_n7403));
  nand_5 g07027(.A(new_n7403), .B(new_n7402), .Y(new_n7404));
  xor_4  g07028(.A(new_n7404), .B(new_n7401), .Y(new_n7405));
  xor_4  g07029(.A(new_n7405), .B(new_n7400), .Y(new_n7406));
  nand_5 g07030(.A(pi236), .B(pi136), .Y(new_n7407));
  xor_4  g07031(.A(new_n7407), .B(new_n7406), .Y(new_n7408));
  or_6   g07032(.A(new_n7381), .B(new_n7380), .Y(new_n7409));
  not_8  g07033(.A(new_n7387), .Y(new_n7410));
  nand_5 g07034(.A(new_n7410), .B(new_n7382), .Y(new_n7411));
  nand_5 g07035(.A(new_n7411), .B(new_n7409), .Y(new_n7412));
  xor_4  g07036(.A(new_n7412), .B(new_n7408), .Y(new_n7413));
  xnor_4 g07037(.A(new_n7413), .B(new_n7395), .Y(new_n7414));
  xor_4  g07038(.A(new_n7394), .B(new_n7388), .Y(new_n7415));
  xor_4  g07039(.A(new_n7343), .B(new_n7342), .Y(new_n7416));
  nor_5  g07040(.A(new_n7391), .B(new_n7390), .Y(new_n7417));
  nor_5  g07041(.A(new_n7417), .B(new_n7393), .Y(new_n7418));
  nand_5 g07042(.A(new_n7418), .B(new_n7416), .Y(new_n7419));
  xor_4  g07043(.A(new_n7418), .B(new_n7416), .Y(new_n7420));
  nor_5  g07044(.A(new_n378), .B(new_n377), .Y(new_n7421));
  nand_5 g07045(.A(pi241), .B(pi027), .Y(new_n7422));
  nand_5 g07046(.A(pi236), .B(pi026), .Y(new_n7423));
  xor_4  g07047(.A(new_n7423), .B(new_n7422), .Y(new_n7424));
  nand_5 g07048(.A(new_n7424), .B(new_n7421), .Y(new_n7425));
  xnor_4 g07049(.A(new_n7424), .B(new_n7421), .Y(new_n7426));
  nand_5 g07050(.A(pi213), .B(pi206), .Y(new_n7427));
  nand_5 g07051(.A(pi212), .B(pi164), .Y(new_n7428));
  nand_5 g07052(.A(new_n7428), .B(new_n7427), .Y(new_n7429));
  nand_5 g07053(.A(new_n7429), .B(new_n7343), .Y(new_n7430));
  or_6   g07054(.A(new_n7430), .B(new_n7426), .Y(new_n7431));
  nand_5 g07055(.A(new_n7431), .B(new_n7425), .Y(new_n7432));
  nand_5 g07056(.A(new_n7432), .B(new_n7420), .Y(new_n7433));
  nand_5 g07057(.A(new_n7433), .B(new_n7419), .Y(new_n7434));
  or_6   g07058(.A(new_n7434), .B(new_n7415), .Y(new_n7435));
  xnor_4 g07059(.A(new_n7355), .B(new_n7344), .Y(new_n7436));
  xor_4  g07060(.A(new_n7434), .B(new_n7415), .Y(new_n7437));
  nand_5 g07061(.A(new_n7437), .B(new_n7436), .Y(new_n7438));
  nand_5 g07062(.A(new_n7438), .B(new_n7435), .Y(new_n7439));
  xor_4  g07063(.A(new_n7439), .B(new_n7414), .Y(new_n7440));
  xor_4  g07064(.A(new_n7440), .B(new_n7373), .Y(new_n7441));
  nand_5 g07065(.A(pi147), .B(pi035), .Y(new_n7442));
  nand_5 g07066(.A(pi208), .B(pi019), .Y(new_n7443));
  nand_5 g07067(.A(pi151), .B(pi139), .Y(new_n7444));
  xor_4  g07068(.A(new_n7444), .B(new_n7443), .Y(new_n7445));
  xnor_4 g07069(.A(new_n7445), .B(new_n7442), .Y(new_n7446));
  nand_5 g07070(.A(pi168), .B(pi019), .Y(new_n7447));
  nand_5 g07071(.A(pi147), .B(pi139), .Y(new_n7448));
  nand_5 g07072(.A(new_n7448), .B(new_n7447), .Y(new_n7449));
  nand_5 g07073(.A(pi208), .B(pi151), .Y(new_n7450));
  or_6   g07074(.A(new_n7448), .B(new_n7447), .Y(new_n7451));
  nand_5 g07075(.A(new_n7451), .B(new_n7450), .Y(new_n7452));
  nand_5 g07076(.A(new_n7452), .B(new_n7449), .Y(new_n7453));
  nand_5 g07077(.A(pi168), .B(pi097), .Y(new_n7454));
  xor_4  g07078(.A(new_n7454), .B(new_n7453), .Y(new_n7455));
  xnor_4 g07079(.A(new_n7455), .B(new_n7446), .Y(new_n7456));
  not_8  g07080(.A(new_n7450), .Y(new_n7457));
  not_8  g07081(.A(new_n7449), .Y(new_n7458));
  nand_5 g07082(.A(new_n7457), .B(new_n380), .Y(new_n7459));
  nand_5 g07083(.A(new_n7459), .B(new_n7458), .Y(new_n7460));
  nand_5 g07084(.A(new_n7460), .B(new_n7451), .Y(new_n7461));
  nand_5 g07085(.A(new_n7461), .B(new_n7457), .Y(new_n7462));
  nor_5  g07086(.A(new_n7462), .B(new_n7456), .Y(new_n7463));
  nand_5 g07087(.A(pi139), .B(pi019), .Y(new_n7464));
  nand_5 g07088(.A(pi151), .B(pi035), .Y(new_n7465));
  nand_5 g07089(.A(pi147), .B(pi015), .Y(new_n7466));
  xor_4  g07090(.A(new_n7466), .B(new_n7465), .Y(new_n7467));
  xor_4  g07091(.A(new_n7467), .B(new_n7464), .Y(new_n7468));
  nand_5 g07092(.A(pi208), .B(pi097), .Y(new_n7469));
  nand_5 g07093(.A(new_n7444), .B(new_n7443), .Y(new_n7470));
  nand_5 g07094(.A(new_n7445), .B(new_n7442), .Y(new_n7471));
  nand_5 g07095(.A(new_n7471), .B(new_n7470), .Y(new_n7472));
  xor_4  g07096(.A(new_n7472), .B(new_n7469), .Y(new_n7473));
  xor_4  g07097(.A(new_n7473), .B(new_n7468), .Y(new_n7474));
  nand_5 g07098(.A(pi168), .B(pi075), .Y(new_n7475));
  or_6   g07099(.A(new_n7454), .B(new_n7453), .Y(new_n7476));
  nand_5 g07100(.A(new_n7455), .B(new_n7446), .Y(new_n7477));
  nand_5 g07101(.A(new_n7477), .B(new_n7476), .Y(new_n7478));
  xor_4  g07102(.A(new_n7478), .B(new_n7475), .Y(new_n7479));
  xor_4  g07103(.A(new_n7479), .B(new_n7474), .Y(new_n7480));
  xor_4  g07104(.A(new_n7480), .B(new_n7463), .Y(new_n7481));
  not_8  g07105(.A(new_n7481), .Y(new_n7482));
  xor_4  g07106(.A(new_n7482), .B(new_n7441), .Y(new_n7483));
  xor_4  g07107(.A(new_n7437), .B(new_n7436), .Y(new_n7484));
  xor_4  g07108(.A(new_n7462), .B(new_n7456), .Y(new_n7485));
  not_8  g07109(.A(new_n7485), .Y(new_n7486));
  nand_5 g07110(.A(new_n7486), .B(new_n7484), .Y(new_n7487));
  xor_4  g07111(.A(new_n7486), .B(new_n7484), .Y(new_n7488));
  xor_4  g07112(.A(new_n7432), .B(new_n7420), .Y(new_n7489));
  nor_5  g07113(.A(new_n7459), .B(new_n7458), .Y(new_n7490));
  nor_5  g07114(.A(new_n7490), .B(new_n7461), .Y(new_n7491));
  or_6   g07115(.A(new_n7491), .B(new_n7489), .Y(new_n7492));
  xor_4  g07116(.A(new_n7491), .B(new_n7489), .Y(new_n7493));
  not_8  g07117(.A(new_n379), .Y(new_n7494));
  nor_5  g07118(.A(new_n380), .B(new_n7494), .Y(new_n7495));
  nand_5 g07119(.A(pi168), .B(pi151), .Y(new_n7496));
  nand_5 g07120(.A(pi208), .B(pi147), .Y(new_n7497));
  xor_4  g07121(.A(new_n7497), .B(new_n7496), .Y(new_n7498));
  or_6   g07122(.A(new_n7498), .B(new_n7495), .Y(new_n7499));
  xnor_4 g07123(.A(new_n7430), .B(new_n7426), .Y(new_n7500));
  xor_4  g07124(.A(new_n7498), .B(new_n7495), .Y(new_n7501));
  nand_5 g07125(.A(new_n7501), .B(new_n7500), .Y(new_n7502));
  nand_5 g07126(.A(new_n7502), .B(new_n7499), .Y(new_n7503));
  nand_5 g07127(.A(new_n7503), .B(new_n7493), .Y(new_n7504));
  nand_5 g07128(.A(new_n7504), .B(new_n7492), .Y(new_n7505));
  nand_5 g07129(.A(new_n7505), .B(new_n7488), .Y(new_n7506));
  nand_5 g07130(.A(new_n7506), .B(new_n7487), .Y(new_n7507));
  xor_4  g07131(.A(new_n7507), .B(new_n7483), .Y(new_n7508));
  nor_5  g07132(.A(new_n7508), .B(new_n7337), .Y(new_n7509));
  xor_4  g07133(.A(new_n7508), .B(new_n7337), .Y(new_n7510));
  not_8  g07134(.A(new_n7510), .Y(new_n7511));
  xor_4  g07135(.A(new_n7330), .B(new_n7329), .Y(new_n7512));
  not_8  g07136(.A(new_n7512), .Y(new_n7513));
  xor_4  g07137(.A(new_n7505), .B(new_n7488), .Y(new_n7514));
  nor_5  g07138(.A(new_n7514), .B(new_n7513), .Y(new_n7515));
  xor_4  g07139(.A(new_n7514), .B(new_n7512), .Y(new_n7516));
  xor_4  g07140(.A(new_n7503), .B(new_n7493), .Y(new_n7517));
  nor_5  g07141(.A(new_n382), .B(new_n381), .Y(new_n7518));
  xor_4  g07142(.A(new_n7326), .B(new_n7325), .Y(new_n7519));
  or_6   g07143(.A(new_n7519), .B(new_n7518), .Y(new_n7520));
  xor_4  g07144(.A(new_n7501), .B(new_n7500), .Y(new_n7521));
  xor_4  g07145(.A(new_n7519), .B(new_n7518), .Y(new_n7522));
  nand_5 g07146(.A(new_n7522), .B(new_n7521), .Y(new_n7523));
  nand_5 g07147(.A(new_n7523), .B(new_n7520), .Y(new_n7524));
  nand_5 g07148(.A(new_n7524), .B(new_n7517), .Y(new_n7525));
  xor_4  g07149(.A(new_n7328), .B(new_n7324), .Y(new_n7526));
  not_8  g07150(.A(new_n7526), .Y(new_n7527));
  xor_4  g07151(.A(new_n7524), .B(new_n7517), .Y(new_n7528));
  nand_5 g07152(.A(new_n7528), .B(new_n7527), .Y(new_n7529));
  nand_5 g07153(.A(new_n7529), .B(new_n7525), .Y(new_n7530));
  nor_5  g07154(.A(new_n7530), .B(new_n7516), .Y(new_n7531));
  nor_5  g07155(.A(new_n7531), .B(new_n7515), .Y(new_n7532));
  nor_5  g07156(.A(new_n7532), .B(new_n7511), .Y(new_n7533));
  or_6   g07157(.A(new_n7533), .B(new_n7509), .Y(new_n7534));
  nand_5 g07158(.A(new_n7534), .B(new_n7335), .Y(new_n7535));
  nand_5 g07159(.A(pi032), .B(pi013), .Y(new_n7536));
  nand_5 g07160(.A(pi206), .B(pi112), .Y(new_n7537));
  nand_5 g07161(.A(pi164), .B(pi105), .Y(new_n7538));
  nand_5 g07162(.A(new_n7538), .B(new_n7537), .Y(new_n7539));
  nand_5 g07163(.A(new_n7539), .B(new_n7231), .Y(new_n7540));
  xor_4  g07164(.A(new_n7540), .B(new_n7536), .Y(new_n7541));
  nand_5 g07165(.A(new_n7358), .B(new_n7357), .Y(new_n7542));
  nand_5 g07166(.A(new_n7359), .B(new_n7229), .Y(new_n7543));
  nand_5 g07167(.A(new_n7543), .B(new_n7542), .Y(new_n7544));
  xor_4  g07168(.A(new_n7544), .B(new_n7541), .Y(new_n7545));
  nand_5 g07169(.A(pi145), .B(pi104), .Y(new_n7546));
  nand_5 g07170(.A(pi246), .B(pi212), .Y(new_n7547));
  and_6  g07171(.A(new_n7547), .B(new_n7546), .Y(new_n7548));
  nand_5 g07172(.A(pi246), .B(pi104), .Y(new_n7549));
  nor_5  g07173(.A(new_n7549), .B(new_n7361), .Y(new_n7550));
  or_6   g07174(.A(new_n7550), .B(new_n7548), .Y(new_n7551));
  xnor_4 g07175(.A(new_n7551), .B(new_n7545), .Y(new_n7552));
  nand_5 g07176(.A(new_n7364), .B(new_n7361), .Y(new_n7553));
  nand_5 g07177(.A(new_n7365), .B(new_n7360), .Y(new_n7554));
  nand_5 g07178(.A(new_n7554), .B(new_n7553), .Y(new_n7555));
  xor_4  g07179(.A(new_n7555), .B(new_n7552), .Y(new_n7556));
  nor_5  g07180(.A(new_n7367), .B(new_n7366), .Y(new_n7557));
  nor_5  g07181(.A(new_n7371), .B(new_n7368), .Y(new_n7558));
  nor_5  g07182(.A(new_n7558), .B(new_n7557), .Y(new_n7559));
  xor_4  g07183(.A(new_n7559), .B(new_n7556), .Y(new_n7560));
  nand_5 g07184(.A(new_n7372), .B(new_n7356), .Y(new_n7561));
  nand_5 g07185(.A(pi213), .B(pi114), .Y(new_n7562));
  xor_4  g07186(.A(new_n7562), .B(new_n7561), .Y(new_n7563));
  xor_4  g07187(.A(new_n7563), .B(new_n7560), .Y(new_n7564));
  nand_5 g07188(.A(pi141), .B(pi008), .Y(new_n7565));
  nand_5 g07189(.A(pi090), .B(pi026), .Y(new_n7566));
  nand_5 g07190(.A(pi047), .B(pi027), .Y(new_n7567));
  nand_5 g07191(.A(new_n7567), .B(new_n7566), .Y(new_n7568));
  nand_5 g07192(.A(pi047), .B(pi026), .Y(new_n7569));
  or_6   g07193(.A(new_n7569), .B(new_n7397), .Y(new_n7570));
  nand_5 g07194(.A(new_n7570), .B(new_n7568), .Y(new_n7571));
  xor_4  g07195(.A(new_n7571), .B(new_n7565), .Y(new_n7572));
  nand_5 g07196(.A(new_n7398), .B(new_n7397), .Y(new_n7573));
  nand_5 g07197(.A(new_n7399), .B(new_n7396), .Y(new_n7574));
  nand_5 g07198(.A(new_n7574), .B(new_n7573), .Y(new_n7575));
  xor_4  g07199(.A(new_n7575), .B(new_n7572), .Y(new_n7576));
  nand_5 g07200(.A(pi241), .B(pi136), .Y(new_n7577));
  nand_5 g07201(.A(pi161), .B(pi056), .Y(new_n7578));
  and_6  g07202(.A(new_n7578), .B(new_n7577), .Y(new_n7579));
  nand_5 g07203(.A(pi161), .B(pi136), .Y(new_n7580));
  nor_5  g07204(.A(new_n7580), .B(new_n7401), .Y(new_n7581));
  or_6   g07205(.A(new_n7581), .B(new_n7579), .Y(new_n7582));
  xnor_4 g07206(.A(new_n7582), .B(new_n7576), .Y(new_n7583));
  nand_5 g07207(.A(new_n7404), .B(new_n7401), .Y(new_n7584));
  nand_5 g07208(.A(new_n7405), .B(new_n7400), .Y(new_n7585));
  nand_5 g07209(.A(new_n7585), .B(new_n7584), .Y(new_n7586));
  xor_4  g07210(.A(new_n7586), .B(new_n7583), .Y(new_n7587));
  or_6   g07211(.A(new_n7407), .B(new_n7406), .Y(new_n7588));
  nand_5 g07212(.A(new_n7412), .B(new_n7408), .Y(new_n7589));
  nand_5 g07213(.A(new_n7589), .B(new_n7588), .Y(new_n7590));
  xnor_4 g07214(.A(new_n7590), .B(new_n7587), .Y(new_n7591));
  nand_5 g07215(.A(new_n7413), .B(new_n7395), .Y(new_n7592));
  nand_5 g07216(.A(pi236), .B(pi096), .Y(new_n7593));
  xor_4  g07217(.A(new_n7593), .B(new_n7592), .Y(new_n7594));
  xor_4  g07218(.A(new_n7594), .B(new_n7591), .Y(new_n7595));
  xnor_4 g07219(.A(new_n7595), .B(new_n7564), .Y(new_n7596));
  nand_5 g07220(.A(new_n7439), .B(new_n7414), .Y(new_n7597));
  nand_5 g07221(.A(new_n7440), .B(new_n7373), .Y(new_n7598));
  nand_5 g07222(.A(new_n7598), .B(new_n7597), .Y(new_n7599));
  xnor_4 g07223(.A(new_n7599), .B(new_n7596), .Y(new_n7600));
  nand_5 g07224(.A(new_n7472), .B(new_n7469), .Y(new_n7601));
  nand_5 g07225(.A(new_n7473), .B(new_n7468), .Y(new_n7602));
  nand_5 g07226(.A(new_n7602), .B(new_n7601), .Y(new_n7603));
  nand_5 g07227(.A(pi035), .B(pi019), .Y(new_n7604));
  nand_5 g07228(.A(new_n7466), .B(new_n7465), .Y(new_n7605));
  nand_5 g07229(.A(new_n7467), .B(new_n7464), .Y(new_n7606));
  nand_5 g07230(.A(new_n7606), .B(new_n7605), .Y(new_n7607));
  xor_4  g07231(.A(new_n7607), .B(new_n7604), .Y(new_n7608));
  nand_5 g07232(.A(pi151), .B(pi015), .Y(new_n7609));
  nand_5 g07233(.A(pi204), .B(pi147), .Y(new_n7610));
  nand_5 g07234(.A(new_n7610), .B(new_n7609), .Y(new_n7611));
  nand_5 g07235(.A(pi204), .B(pi151), .Y(new_n7612));
  nor_5  g07236(.A(new_n7612), .B(new_n7466), .Y(new_n7613));
  not_8  g07237(.A(new_n7613), .Y(new_n7614));
  nand_5 g07238(.A(new_n7614), .B(new_n7611), .Y(new_n7615));
  xor_4  g07239(.A(new_n7615), .B(new_n7608), .Y(new_n7616));
  nand_5 g07240(.A(pi139), .B(pi097), .Y(new_n7617));
  nand_5 g07241(.A(pi208), .B(pi075), .Y(new_n7618));
  nand_5 g07242(.A(new_n7618), .B(new_n7617), .Y(new_n7619));
  nand_5 g07243(.A(pi139), .B(pi075), .Y(new_n7620));
  or_6   g07244(.A(new_n7620), .B(new_n7469), .Y(new_n7621));
  nand_5 g07245(.A(new_n7621), .B(new_n7619), .Y(new_n7622));
  xor_4  g07246(.A(new_n7622), .B(new_n7616), .Y(new_n7623));
  xor_4  g07247(.A(new_n7623), .B(new_n7603), .Y(new_n7624));
  not_8  g07248(.A(new_n7475), .Y(new_n7625));
  nand_5 g07249(.A(new_n7478), .B(new_n7625), .Y(new_n7626));
  or_6   g07250(.A(new_n7479), .B(new_n7474), .Y(new_n7627));
  nand_5 g07251(.A(new_n7627), .B(new_n7626), .Y(new_n7628));
  xor_4  g07252(.A(new_n7628), .B(new_n7624), .Y(new_n7629));
  nand_5 g07253(.A(new_n7480), .B(new_n7463), .Y(new_n7630));
  nand_5 g07254(.A(pi168), .B(pi093), .Y(new_n7631));
  xor_4  g07255(.A(new_n7631), .B(new_n7630), .Y(new_n7632));
  xor_4  g07256(.A(new_n7632), .B(new_n7629), .Y(new_n7633));
  xor_4  g07257(.A(new_n7633), .B(new_n7600), .Y(new_n7634));
  nand_5 g07258(.A(new_n7482), .B(new_n7441), .Y(new_n7635));
  nand_5 g07259(.A(new_n7507), .B(new_n7483), .Y(new_n7636));
  nand_5 g07260(.A(new_n7636), .B(new_n7635), .Y(new_n7637));
  xnor_4 g07261(.A(new_n7637), .B(new_n7634), .Y(new_n7638));
  xor_4  g07262(.A(new_n7534), .B(new_n7335), .Y(new_n7639));
  nand_5 g07263(.A(new_n7639), .B(new_n7638), .Y(new_n7640));
  nand_5 g07264(.A(new_n7640), .B(new_n7535), .Y(new_n7641));
  nand_5 g07265(.A(new_n7333), .B(new_n7323), .Y(new_n7642));
  not_8  g07266(.A(new_n7322), .Y(new_n7643));
  nand_5 g07267(.A(new_n7334), .B(new_n7643), .Y(new_n7644));
  nand_5 g07268(.A(new_n7644), .B(new_n7642), .Y(new_n7645));
  nand_5 g07269(.A(new_n7321), .B(new_n7302), .Y(new_n7646));
  xor_4  g07270(.A(new_n7297), .B(new_n7294), .Y(new_n7647));
  xor_4  g07271(.A(new_n7647), .B(new_n7646), .Y(new_n7648));
  xnor_4 g07272(.A(new_n7648), .B(new_n7645), .Y(new_n7649));
  or_6   g07273(.A(new_n7649), .B(new_n7641), .Y(new_n7650));
  not_8  g07274(.A(new_n7559), .Y(new_n7651));
  nand_5 g07275(.A(new_n7651), .B(new_n7556), .Y(new_n7652));
  xor_4  g07276(.A(new_n7238), .B(new_n7236), .Y(new_n7653));
  nand_5 g07277(.A(pi212), .B(pi114), .Y(new_n7654));
  nand_5 g07278(.A(pi213), .B(pi091), .Y(new_n7655));
  xor_4  g07279(.A(new_n7655), .B(new_n7654), .Y(new_n7656));
  xor_4  g07280(.A(new_n7656), .B(new_n7549), .Y(new_n7657));
  nand_5 g07281(.A(new_n7540), .B(new_n7536), .Y(new_n7658));
  nand_5 g07282(.A(new_n7544), .B(new_n7541), .Y(new_n7659));
  nand_5 g07283(.A(new_n7659), .B(new_n7658), .Y(new_n7660));
  xor_4  g07284(.A(new_n7660), .B(new_n7657), .Y(new_n7661));
  xnor_4 g07285(.A(new_n7661), .B(new_n7653), .Y(new_n7662));
  nor_5  g07286(.A(new_n7551), .B(new_n7545), .Y(new_n7663));
  nor_5  g07287(.A(new_n7555), .B(new_n7552), .Y(new_n7664));
  xor_4  g07288(.A(new_n7664), .B(new_n7550), .Y(new_n7665));
  nor_5  g07289(.A(new_n7665), .B(new_n7663), .Y(new_n7666));
  xor_4  g07290(.A(new_n7666), .B(new_n7662), .Y(new_n7667));
  xnor_4 g07291(.A(new_n7667), .B(new_n7652), .Y(new_n7668));
  nand_5 g07292(.A(new_n7562), .B(new_n7561), .Y(new_n7669));
  nand_5 g07293(.A(new_n7563), .B(new_n7560), .Y(new_n7670));
  nand_5 g07294(.A(new_n7670), .B(new_n7669), .Y(new_n7671));
  xnor_4 g07295(.A(new_n7671), .B(new_n7668), .Y(new_n7672));
  nand_5 g07296(.A(new_n7590), .B(new_n7587), .Y(new_n7673));
  nand_5 g07297(.A(pi027), .B(pi018), .Y(new_n7674));
  nand_5 g07298(.A(pi090), .B(pi008), .Y(new_n7675));
  xor_4  g07299(.A(new_n7675), .B(new_n7674), .Y(new_n7676));
  xor_4  g07300(.A(new_n7676), .B(new_n7569), .Y(new_n7677));
  nand_5 g07301(.A(pi141), .B(pi056), .Y(new_n7678));
  xor_4  g07302(.A(new_n7678), .B(new_n7570), .Y(new_n7679));
  xor_4  g07303(.A(new_n7679), .B(new_n7677), .Y(new_n7680));
  nand_5 g07304(.A(pi241), .B(pi096), .Y(new_n7681));
  nand_5 g07305(.A(pi236), .B(pi235), .Y(new_n7682));
  xor_4  g07306(.A(new_n7682), .B(new_n7681), .Y(new_n7683));
  xor_4  g07307(.A(new_n7683), .B(new_n7580), .Y(new_n7684));
  nand_5 g07308(.A(new_n7571), .B(new_n7565), .Y(new_n7685));
  nand_5 g07309(.A(new_n7575), .B(new_n7572), .Y(new_n7686));
  nand_5 g07310(.A(new_n7686), .B(new_n7685), .Y(new_n7687));
  xor_4  g07311(.A(new_n7687), .B(new_n7684), .Y(new_n7688));
  xnor_4 g07312(.A(new_n7688), .B(new_n7680), .Y(new_n7689));
  nor_5  g07313(.A(new_n7582), .B(new_n7576), .Y(new_n7690));
  nor_5  g07314(.A(new_n7586), .B(new_n7583), .Y(new_n7691));
  xor_4  g07315(.A(new_n7691), .B(new_n7581), .Y(new_n7692));
  nor_5  g07316(.A(new_n7692), .B(new_n7690), .Y(new_n7693));
  xor_4  g07317(.A(new_n7693), .B(new_n7689), .Y(new_n7694));
  xnor_4 g07318(.A(new_n7694), .B(new_n7673), .Y(new_n7695));
  nand_5 g07319(.A(new_n7593), .B(new_n7592), .Y(new_n7696));
  nand_5 g07320(.A(new_n7594), .B(new_n7591), .Y(new_n7697));
  nand_5 g07321(.A(new_n7697), .B(new_n7696), .Y(new_n7698));
  xor_4  g07322(.A(new_n7698), .B(new_n7695), .Y(new_n7699));
  not_8  g07323(.A(new_n7699), .Y(new_n7700));
  xor_4  g07324(.A(new_n7700), .B(new_n7672), .Y(new_n7701));
  nor_5  g07325(.A(new_n7595), .B(new_n7564), .Y(new_n7702));
  nor_5  g07326(.A(new_n7599), .B(new_n7596), .Y(new_n7703));
  nor_5  g07327(.A(new_n7703), .B(new_n7702), .Y(new_n7704));
  xor_4  g07328(.A(new_n7704), .B(new_n7701), .Y(new_n7705));
  not_8  g07329(.A(new_n7624), .Y(new_n7706));
  nand_5 g07330(.A(new_n7628), .B(new_n7706), .Y(new_n7707));
  nand_5 g07331(.A(pi147), .B(pi146), .Y(new_n7708));
  nand_5 g07332(.A(pi019), .B(pi015), .Y(new_n7709));
  xor_4  g07333(.A(new_n7709), .B(new_n7708), .Y(new_n7710));
  xor_4  g07334(.A(new_n7710), .B(new_n7612), .Y(new_n7711));
  nand_5 g07335(.A(pi097), .B(pi035), .Y(new_n7712));
  xor_4  g07336(.A(new_n7712), .B(new_n7614), .Y(new_n7713));
  not_8  g07337(.A(new_n7713), .Y(new_n7714));
  xor_4  g07338(.A(new_n7714), .B(new_n7711), .Y(new_n7715));
  nand_5 g07339(.A(pi208), .B(pi093), .Y(new_n7716));
  nand_5 g07340(.A(pi168), .B(pi166), .Y(new_n7717));
  xor_4  g07341(.A(new_n7717), .B(new_n7716), .Y(new_n7718));
  xor_4  g07342(.A(new_n7718), .B(new_n7620), .Y(new_n7719));
  nand_5 g07343(.A(new_n7607), .B(new_n7604), .Y(new_n7720));
  nand_5 g07344(.A(new_n7615), .B(new_n7608), .Y(new_n7721));
  nand_5 g07345(.A(new_n7721), .B(new_n7720), .Y(new_n7722));
  xor_4  g07346(.A(new_n7722), .B(new_n7719), .Y(new_n7723));
  xor_4  g07347(.A(new_n7723), .B(new_n7715), .Y(new_n7724));
  nand_5 g07348(.A(new_n7622), .B(new_n7616), .Y(new_n7725));
  nand_5 g07349(.A(new_n7623), .B(new_n7603), .Y(new_n7726));
  nand_5 g07350(.A(new_n7726), .B(new_n7725), .Y(new_n7727));
  xor_4  g07351(.A(new_n7727), .B(new_n7621), .Y(new_n7728));
  xnor_4 g07352(.A(new_n7728), .B(new_n7724), .Y(new_n7729));
  xnor_4 g07353(.A(new_n7729), .B(new_n7707), .Y(new_n7730));
  nand_5 g07354(.A(new_n7631), .B(new_n7630), .Y(new_n7731));
  nand_5 g07355(.A(new_n7632), .B(new_n7629), .Y(new_n7732));
  nand_5 g07356(.A(new_n7732), .B(new_n7731), .Y(new_n7733));
  xor_4  g07357(.A(new_n7733), .B(new_n7730), .Y(new_n7734));
  not_8  g07358(.A(new_n7734), .Y(new_n7735));
  xor_4  g07359(.A(new_n7735), .B(new_n7705), .Y(new_n7736));
  nand_5 g07360(.A(new_n7633), .B(new_n7600), .Y(new_n7737));
  nand_5 g07361(.A(new_n7637), .B(new_n7634), .Y(new_n7738));
  nand_5 g07362(.A(new_n7738), .B(new_n7737), .Y(new_n7739));
  xor_4  g07363(.A(new_n7739), .B(new_n7736), .Y(new_n7740));
  xor_4  g07364(.A(new_n7649), .B(new_n7641), .Y(new_n7741));
  nand_5 g07365(.A(new_n7741), .B(new_n7740), .Y(new_n7742));
  nand_5 g07366(.A(new_n7742), .B(new_n7650), .Y(new_n7743));
  xor_4  g07367(.A(new_n7743), .B(new_n7301), .Y(new_n7744));
  xor_4  g07368(.A(new_n7744), .B(new_n7300), .Y(new_n7745));
  nand_5 g07369(.A(pi131), .B(pi009), .Y(new_n7746));
  nand_5 g07370(.A(new_n7647), .B(new_n7646), .Y(new_n7747));
  nand_5 g07371(.A(new_n7648), .B(new_n7645), .Y(new_n7748));
  nand_5 g07372(.A(new_n7748), .B(new_n7747), .Y(new_n7749));
  nand_5 g07373(.A(pi119), .B(pi034), .Y(new_n7750));
  xor_4  g07374(.A(new_n7750), .B(new_n7749), .Y(new_n7751));
  xor_4  g07375(.A(new_n7751), .B(new_n7746), .Y(new_n7752));
  nand_5 g07376(.A(new_n7675), .B(new_n7674), .Y(new_n7753));
  nand_5 g07377(.A(new_n7676), .B(new_n7569), .Y(new_n7754));
  nand_5 g07378(.A(new_n7754), .B(new_n7753), .Y(new_n7755));
  or_6   g07379(.A(new_n7678), .B(new_n7570), .Y(new_n7756));
  not_8  g07380(.A(new_n7677), .Y(new_n7757));
  nand_5 g07381(.A(new_n7679), .B(new_n7757), .Y(new_n7758));
  nand_5 g07382(.A(new_n7758), .B(new_n7756), .Y(new_n7759));
  nand_5 g07383(.A(new_n7687), .B(new_n7684), .Y(new_n7760));
  nand_5 g07384(.A(new_n7688), .B(new_n7680), .Y(new_n7761));
  nand_5 g07385(.A(new_n7761), .B(new_n7760), .Y(new_n7762));
  nand_5 g07386(.A(new_n7682), .B(new_n7681), .Y(new_n7763));
  nand_5 g07387(.A(new_n7683), .B(new_n7580), .Y(new_n7764));
  nand_5 g07388(.A(new_n7764), .B(new_n7763), .Y(new_n7765));
  xor_4  g07389(.A(new_n7765), .B(new_n7762), .Y(new_n7766));
  nand_5 g07390(.A(pi161), .B(pi096), .Y(new_n7767));
  xor_4  g07391(.A(new_n7767), .B(new_n7766), .Y(new_n7768));
  xor_4  g07392(.A(new_n7768), .B(new_n7759), .Y(new_n7769));
  xor_4  g07393(.A(new_n7769), .B(new_n7755), .Y(new_n7770));
  xor_4  g07394(.A(new_n7770), .B(new_n7752), .Y(new_n7771));
  xor_4  g07395(.A(new_n7771), .B(new_n7745), .Y(new_n7772));
  xor_4  g07396(.A(new_n7772), .B(new_n7240), .Y(new_n7773));
  nand_5 g07397(.A(new_n7655), .B(new_n7654), .Y(new_n7774));
  nand_5 g07398(.A(new_n7656), .B(new_n7549), .Y(new_n7775));
  nand_5 g07399(.A(new_n7775), .B(new_n7774), .Y(new_n7776));
  nor_5  g07400(.A(new_n7694), .B(new_n7673), .Y(new_n7777));
  nor_5  g07401(.A(new_n7698), .B(new_n7695), .Y(new_n7778));
  nor_5  g07402(.A(new_n7778), .B(new_n7777), .Y(new_n7779));
  xor_4  g07403(.A(new_n7779), .B(new_n7776), .Y(new_n7780));
  nand_5 g07404(.A(pi212), .B(pi091), .Y(new_n7781));
  nand_5 g07405(.A(pi114), .B(pi104), .Y(new_n7782));
  xor_4  g07406(.A(new_n7782), .B(new_n7781), .Y(new_n7783));
  nand_5 g07407(.A(new_n7691), .B(new_n7581), .Y(new_n7784));
  not_8  g07408(.A(new_n7693), .Y(new_n7785));
  nand_5 g07409(.A(new_n7785), .B(new_n7689), .Y(new_n7786));
  nand_5 g07410(.A(new_n7786), .B(new_n7784), .Y(new_n7787));
  nand_5 g07411(.A(pi090), .B(pi056), .Y(new_n7788));
  nand_5 g07412(.A(pi141), .B(pi136), .Y(new_n7789));
  xor_4  g07413(.A(new_n7789), .B(new_n7788), .Y(new_n7790));
  xor_4  g07414(.A(new_n7790), .B(new_n7787), .Y(new_n7791));
  nand_5 g07415(.A(pi047), .B(pi008), .Y(new_n7792));
  nand_5 g07416(.A(pi236), .B(pi110), .Y(new_n7793));
  nand_5 g07417(.A(pi026), .B(pi018), .Y(new_n7794));
  nand_5 g07418(.A(pi128), .B(pi027), .Y(new_n7795));
  xor_4  g07419(.A(new_n7795), .B(new_n7794), .Y(new_n7796));
  xor_4  g07420(.A(new_n7796), .B(new_n7793), .Y(new_n7797));
  xor_4  g07421(.A(new_n7797), .B(new_n7792), .Y(new_n7798));
  xor_4  g07422(.A(new_n7798), .B(new_n7791), .Y(new_n7799));
  xor_4  g07423(.A(new_n7799), .B(new_n7783), .Y(new_n7800));
  xor_4  g07424(.A(new_n7800), .B(new_n7780), .Y(new_n7801));
  nand_5 g07425(.A(pi164), .B(pi088), .Y(new_n7802));
  nand_5 g07426(.A(pi206), .B(pi183), .Y(new_n7803));
  nand_5 g07427(.A(pi105), .B(pi032), .Y(new_n7804));
  xor_4  g07428(.A(new_n7804), .B(new_n7803), .Y(new_n7805));
  nand_5 g07429(.A(pi213), .B(pi031), .Y(new_n7806));
  nand_5 g07430(.A(new_n7700), .B(new_n7672), .Y(new_n7807));
  nand_5 g07431(.A(new_n7704), .B(new_n7701), .Y(new_n7808));
  nand_5 g07432(.A(new_n7808), .B(new_n7807), .Y(new_n7809));
  xor_4  g07433(.A(new_n7809), .B(new_n7806), .Y(new_n7810));
  xor_4  g07434(.A(new_n7810), .B(new_n7805), .Y(new_n7811));
  xor_4  g07435(.A(new_n7811), .B(new_n7802), .Y(new_n7812));
  nand_5 g07436(.A(pi075), .B(pi035), .Y(new_n7813));
  nand_5 g07437(.A(pi139), .B(pi093), .Y(new_n7814));
  xor_4  g07438(.A(new_n7814), .B(new_n7813), .Y(new_n7815));
  nand_5 g07439(.A(pi204), .B(pi019), .Y(new_n7816));
  xor_4  g07440(.A(new_n7816), .B(new_n7815), .Y(new_n7817));
  nand_5 g07441(.A(pi208), .B(pi166), .Y(new_n7818));
  nand_5 g07442(.A(new_n7709), .B(new_n7708), .Y(new_n7819));
  nand_5 g07443(.A(new_n7710), .B(new_n7612), .Y(new_n7820));
  nand_5 g07444(.A(new_n7820), .B(new_n7819), .Y(new_n7821));
  nor_5  g07445(.A(new_n7712), .B(new_n7614), .Y(new_n7822));
  nor_5  g07446(.A(new_n7714), .B(new_n7711), .Y(new_n7823));
  or_6   g07447(.A(new_n7823), .B(new_n7822), .Y(new_n7824));
  xor_4  g07448(.A(new_n7824), .B(new_n7821), .Y(new_n7825));
  xor_4  g07449(.A(new_n7825), .B(new_n7818), .Y(new_n7826));
  xor_4  g07450(.A(new_n7826), .B(new_n7817), .Y(new_n7827));
  xor_4  g07451(.A(new_n7827), .B(new_n7812), .Y(new_n7828));
  nand_5 g07452(.A(new_n7664), .B(new_n7550), .Y(new_n7829));
  not_8  g07453(.A(new_n7666), .Y(new_n7830));
  nand_5 g07454(.A(new_n7830), .B(new_n7662), .Y(new_n7831));
  nand_5 g07455(.A(new_n7831), .B(new_n7829), .Y(new_n7832));
  nor_5  g07456(.A(new_n7667), .B(new_n7652), .Y(new_n7833));
  nor_5  g07457(.A(new_n7671), .B(new_n7668), .Y(new_n7834));
  or_6   g07458(.A(new_n7834), .B(new_n7833), .Y(new_n7835));
  xor_4  g07459(.A(new_n7835), .B(new_n7832), .Y(new_n7836));
  nand_5 g07460(.A(new_n7717), .B(new_n7716), .Y(new_n7837));
  nand_5 g07461(.A(new_n7718), .B(new_n7620), .Y(new_n7838));
  nand_5 g07462(.A(new_n7838), .B(new_n7837), .Y(new_n7839));
  nand_5 g07463(.A(pi097), .B(pi015), .Y(new_n7840));
  nand_5 g07464(.A(new_n7722), .B(new_n7719), .Y(new_n7841));
  not_8  g07465(.A(new_n7715), .Y(new_n7842));
  nand_5 g07466(.A(new_n7723), .B(new_n7842), .Y(new_n7843));
  nand_5 g07467(.A(new_n7843), .B(new_n7841), .Y(new_n7844));
  xor_4  g07468(.A(new_n7844), .B(new_n7840), .Y(new_n7845));
  xor_4  g07469(.A(new_n7845), .B(new_n7839), .Y(new_n7846));
  xor_4  g07470(.A(new_n7846), .B(new_n7836), .Y(new_n7847));
  xor_4  g07471(.A(new_n7847), .B(new_n7828), .Y(new_n7848));
  nand_5 g07472(.A(pi084), .B(pi045), .Y(new_n7849));
  nand_5 g07473(.A(pi248), .B(pi052), .Y(new_n7850));
  nand_5 g07474(.A(pi077), .B(pi072), .Y(new_n7851));
  xor_4  g07475(.A(new_n7851), .B(new_n7850), .Y(new_n7852));
  xor_4  g07476(.A(new_n7852), .B(new_n7849), .Y(new_n7853));
  xor_4  g07477(.A(new_n7853), .B(new_n7848), .Y(new_n7854));
  nand_5 g07478(.A(new_n7292), .B(new_n7289), .Y(new_n7855));
  nand_5 g07479(.A(new_n7293), .B(new_n7285), .Y(new_n7856));
  nand_5 g07480(.A(new_n7856), .B(new_n7855), .Y(new_n7857));
  nand_5 g07481(.A(new_n7287), .B(new_n7286), .Y(new_n7858));
  nand_5 g07482(.A(new_n7288), .B(new_n7241), .Y(new_n7859));
  nand_5 g07483(.A(new_n7859), .B(new_n7858), .Y(new_n7860));
  xor_4  g07484(.A(new_n7860), .B(new_n7857), .Y(new_n7861));
  nand_5 g07485(.A(pi189), .B(pi044), .Y(new_n7862));
  nand_5 g07486(.A(pi133), .B(pi054), .Y(new_n7863));
  xor_4  g07487(.A(new_n7863), .B(new_n7862), .Y(new_n7864));
  xor_4  g07488(.A(new_n7864), .B(new_n7861), .Y(new_n7865));
  nor_5  g07489(.A(new_n7729), .B(new_n7707), .Y(new_n7866));
  nor_5  g07490(.A(new_n7733), .B(new_n7730), .Y(new_n7867));
  nor_5  g07491(.A(new_n7867), .B(new_n7866), .Y(new_n7868));
  nand_5 g07492(.A(pi250), .B(pi064), .Y(new_n7869));
  xor_4  g07493(.A(new_n7869), .B(new_n7868), .Y(new_n7870));
  xor_4  g07494(.A(new_n7870), .B(new_n7865), .Y(new_n7871));
  or_6   g07495(.A(new_n7727), .B(new_n7621), .Y(new_n7872));
  nand_5 g07496(.A(new_n7728), .B(new_n7724), .Y(new_n7873));
  nand_5 g07497(.A(new_n7873), .B(new_n7872), .Y(new_n7874));
  nand_5 g07498(.A(pi168), .B(pi011), .Y(new_n7875));
  xor_4  g07499(.A(new_n7875), .B(new_n7874), .Y(new_n7876));
  nand_5 g07500(.A(pi152), .B(pi147), .Y(new_n7877));
  nand_5 g07501(.A(pi151), .B(pi146), .Y(new_n7878));
  xor_4  g07502(.A(new_n7878), .B(new_n7877), .Y(new_n7879));
  xor_4  g07503(.A(new_n7879), .B(new_n7876), .Y(new_n7880));
  nand_5 g07504(.A(new_n7280), .B(new_n7279), .Y(new_n7881));
  nand_5 g07505(.A(new_n7281), .B(new_n7249), .Y(new_n7882));
  nand_5 g07506(.A(new_n7882), .B(new_n7881), .Y(new_n7883));
  or_6   g07507(.A(new_n7283), .B(new_n7250), .Y(new_n7884));
  not_8  g07508(.A(new_n7282), .Y(new_n7885));
  nand_5 g07509(.A(new_n7284), .B(new_n7885), .Y(new_n7886));
  nand_5 g07510(.A(new_n7886), .B(new_n7884), .Y(new_n7887));
  xor_4  g07511(.A(new_n7887), .B(new_n7883), .Y(new_n7888));
  xor_4  g07512(.A(new_n7888), .B(new_n7880), .Y(new_n7889));
  xor_4  g07513(.A(new_n7889), .B(new_n7871), .Y(new_n7890));
  xor_4  g07514(.A(new_n7890), .B(new_n7854), .Y(new_n7891));
  nand_5 g07515(.A(pi246), .B(pi013), .Y(new_n7892));
  nand_5 g07516(.A(new_n7660), .B(new_n7657), .Y(new_n7893));
  nand_5 g07517(.A(new_n7661), .B(new_n7653), .Y(new_n7894));
  nand_5 g07518(.A(new_n7894), .B(new_n7893), .Y(new_n7895));
  xor_4  g07519(.A(new_n7895), .B(new_n7892), .Y(new_n7896));
  nand_5 g07520(.A(pi145), .B(pi112), .Y(new_n7897));
  xor_4  g07521(.A(new_n7897), .B(new_n7896), .Y(new_n7898));
  xor_4  g07522(.A(new_n7898), .B(new_n7891), .Y(new_n7899));
  xor_4  g07523(.A(new_n7899), .B(new_n7801), .Y(new_n7900));
  nand_5 g07524(.A(new_n7735), .B(new_n7705), .Y(new_n7901));
  nand_5 g07525(.A(new_n7739), .B(new_n7736), .Y(new_n7902));
  nand_5 g07526(.A(new_n7902), .B(new_n7901), .Y(new_n7903));
  nand_5 g07527(.A(new_n7234), .B(new_n7233), .Y(new_n7904));
  nand_5 g07528(.A(new_n7235), .B(new_n7230), .Y(new_n7905));
  nand_5 g07529(.A(new_n7905), .B(new_n7904), .Y(new_n7906));
  xor_4  g07530(.A(new_n7906), .B(new_n7903), .Y(new_n7907));
  xor_4  g07531(.A(new_n7907), .B(new_n7900), .Y(new_n7908));
  xor_4  g07532(.A(new_n7908), .B(new_n7773), .Y(po039));
  xor_4  g07533(.A(new_n7639), .B(new_n7638), .Y(po040));
  nand_5 g07534(.A(pi163), .B(pi066), .Y(new_n7911));
  xor_4  g07535(.A(new_n7911), .B(new_n4966), .Y(new_n7912));
  nand_5 g07536(.A(pi228), .B(pi226), .Y(new_n7913));
  xor_4  g07537(.A(new_n7913), .B(new_n7912), .Y(new_n7914));
  or_6   g07538(.A(new_n7914), .B(new_n4968), .Y(new_n7915));
  nand_5 g07539(.A(pi228), .B(pi207), .Y(new_n7916));
  nand_5 g07540(.A(pi148), .B(pi066), .Y(new_n7917));
  nand_5 g07541(.A(pi226), .B(pi039), .Y(new_n7918));
  xor_4  g07542(.A(new_n7918), .B(new_n7917), .Y(new_n7919));
  xor_4  g07543(.A(new_n7919), .B(new_n7916), .Y(new_n7920));
  nand_5 g07544(.A(pi163), .B(pi055), .Y(new_n7921));
  nand_5 g07545(.A(new_n7911), .B(new_n4966), .Y(new_n7922));
  nand_5 g07546(.A(new_n7913), .B(new_n7912), .Y(new_n7923));
  nand_5 g07547(.A(new_n7923), .B(new_n7922), .Y(new_n7924));
  xor_4  g07548(.A(new_n7924), .B(new_n7921), .Y(new_n7925));
  xor_4  g07549(.A(new_n7925), .B(new_n7920), .Y(new_n7926));
  or_6   g07550(.A(new_n7926), .B(new_n7915), .Y(new_n7927));
  nand_5 g07551(.A(pi163), .B(pi002), .Y(new_n7928));
  nand_5 g07552(.A(new_n7924), .B(new_n7921), .Y(new_n7929));
  nand_5 g07553(.A(new_n7925), .B(new_n7920), .Y(new_n7930));
  nand_5 g07554(.A(new_n7930), .B(new_n7929), .Y(new_n7931));
  xor_4  g07555(.A(new_n7931), .B(new_n7928), .Y(new_n7932));
  nand_5 g07556(.A(pi226), .B(pi116), .Y(new_n7933));
  nand_5 g07557(.A(pi228), .B(pi066), .Y(new_n7934));
  nand_5 g07558(.A(pi207), .B(pi039), .Y(new_n7935));
  xor_4  g07559(.A(new_n7935), .B(new_n7934), .Y(new_n7936));
  xor_4  g07560(.A(new_n7936), .B(new_n7933), .Y(new_n7937));
  nand_5 g07561(.A(pi148), .B(pi055), .Y(new_n7938));
  nand_5 g07562(.A(new_n7918), .B(new_n7917), .Y(new_n7939));
  nand_5 g07563(.A(new_n7919), .B(new_n7916), .Y(new_n7940));
  nand_5 g07564(.A(new_n7940), .B(new_n7939), .Y(new_n7941));
  xor_4  g07565(.A(new_n7941), .B(new_n7938), .Y(new_n7942));
  xnor_4 g07566(.A(new_n7942), .B(new_n7937), .Y(new_n7943));
  xnor_4 g07567(.A(new_n7943), .B(new_n7932), .Y(new_n7944));
  xor_4  g07568(.A(new_n7944), .B(new_n7927), .Y(new_n7945));
  nand_5 g07569(.A(pi173), .B(pi107), .Y(new_n7946));
  xor_4  g07570(.A(new_n7946), .B(new_n4974), .Y(new_n7947));
  nand_5 g07571(.A(pi109), .B(pi049), .Y(new_n7948));
  xor_4  g07572(.A(new_n7948), .B(new_n7947), .Y(new_n7949));
  or_6   g07573(.A(new_n7949), .B(new_n4976), .Y(new_n7950));
  nand_5 g07574(.A(pi173), .B(pi171), .Y(new_n7951));
  nand_5 g07575(.A(pi245), .B(pi109), .Y(new_n7952));
  nand_5 g07576(.A(pi049), .B(pi014), .Y(new_n7953));
  xor_4  g07577(.A(new_n7953), .B(new_n7952), .Y(new_n7954));
  xor_4  g07578(.A(new_n7954), .B(new_n7951), .Y(new_n7955));
  nand_5 g07579(.A(pi230), .B(pi107), .Y(new_n7956));
  nand_5 g07580(.A(new_n7946), .B(new_n4974), .Y(new_n7957));
  nand_5 g07581(.A(new_n7948), .B(new_n7947), .Y(new_n7958));
  nand_5 g07582(.A(new_n7958), .B(new_n7957), .Y(new_n7959));
  xor_4  g07583(.A(new_n7959), .B(new_n7956), .Y(new_n7960));
  xor_4  g07584(.A(new_n7960), .B(new_n7955), .Y(new_n7961));
  nor_5  g07585(.A(new_n7961), .B(new_n7950), .Y(new_n7962));
  nand_5 g07586(.A(pi173), .B(pi049), .Y(new_n7963));
  nand_5 g07587(.A(pi245), .B(pi014), .Y(new_n7964));
  nand_5 g07588(.A(pi201), .B(pi109), .Y(new_n7965));
  xor_4  g07589(.A(new_n7965), .B(new_n7964), .Y(new_n7966));
  xor_4  g07590(.A(new_n7966), .B(new_n7963), .Y(new_n7967));
  nand_5 g07591(.A(pi230), .B(pi171), .Y(new_n7968));
  nand_5 g07592(.A(new_n7953), .B(new_n7952), .Y(new_n7969));
  nand_5 g07593(.A(new_n7954), .B(new_n7951), .Y(new_n7970));
  nand_5 g07594(.A(new_n7970), .B(new_n7969), .Y(new_n7971));
  xor_4  g07595(.A(new_n7971), .B(new_n7968), .Y(new_n7972));
  xnor_4 g07596(.A(new_n7972), .B(new_n7967), .Y(new_n7973));
  nand_5 g07597(.A(pi107), .B(pi050), .Y(new_n7974));
  nand_5 g07598(.A(new_n7959), .B(new_n7956), .Y(new_n7975));
  nand_5 g07599(.A(new_n7960), .B(new_n7955), .Y(new_n7976));
  nand_5 g07600(.A(new_n7976), .B(new_n7975), .Y(new_n7977));
  xor_4  g07601(.A(new_n7977), .B(new_n7974), .Y(new_n7978));
  xor_4  g07602(.A(new_n7978), .B(new_n7973), .Y(new_n7979));
  xor_4  g07603(.A(new_n7979), .B(new_n7962), .Y(new_n7980));
  xor_4  g07604(.A(new_n7980), .B(new_n7945), .Y(new_n7981));
  xor_4  g07605(.A(new_n7961), .B(new_n7950), .Y(new_n7982));
  xor_4  g07606(.A(new_n7926), .B(new_n7915), .Y(new_n7983));
  nand_5 g07607(.A(new_n7983), .B(new_n7982), .Y(new_n7984));
  not_8  g07608(.A(new_n7984), .Y(new_n7985));
  xnor_4 g07609(.A(new_n7983), .B(new_n7982), .Y(new_n7986));
  xor_4  g07610(.A(new_n7949), .B(new_n4975), .Y(new_n7987));
  not_8  g07611(.A(new_n4962), .Y(new_n7988));
  nor_5  g07612(.A(new_n4969), .B(new_n7988), .Y(new_n7989));
  nor_5  g07613(.A(new_n4977), .B(new_n4970), .Y(new_n7990));
  nor_5  g07614(.A(new_n7990), .B(new_n7989), .Y(new_n7991));
  nand_5 g07615(.A(new_n7991), .B(new_n7987), .Y(new_n7992));
  xor_4  g07616(.A(new_n7914), .B(new_n4968), .Y(new_n7993));
  not_8  g07617(.A(new_n7993), .Y(new_n7994));
  xor_4  g07618(.A(new_n7991), .B(new_n7987), .Y(new_n7995));
  nand_5 g07619(.A(new_n7995), .B(new_n7994), .Y(new_n7996));
  nand_5 g07620(.A(new_n7996), .B(new_n7992), .Y(new_n7997));
  nor_5  g07621(.A(new_n7997), .B(new_n7986), .Y(new_n7998));
  nor_5  g07622(.A(new_n7998), .B(new_n7985), .Y(new_n7999));
  not_8  g07623(.A(new_n7999), .Y(new_n8000));
  xor_4  g07624(.A(new_n8000), .B(new_n7981), .Y(new_n8001));
  nand_5 g07625(.A(pi175), .B(pi058), .Y(new_n8002));
  xor_4  g07626(.A(new_n8002), .B(new_n4986), .Y(new_n8003));
  nand_5 g07627(.A(pi240), .B(pi132), .Y(new_n8004));
  xor_4  g07628(.A(new_n8004), .B(new_n8003), .Y(new_n8005));
  not_8  g07629(.A(new_n8005), .Y(new_n8006));
  nand_5 g07630(.A(new_n8006), .B(new_n4987), .Y(new_n8007));
  nand_5 g07631(.A(pi211), .B(pi175), .Y(new_n8008));
  nand_5 g07632(.A(new_n8002), .B(new_n4986), .Y(new_n8009));
  nand_5 g07633(.A(new_n8004), .B(new_n8003), .Y(new_n8010));
  nand_5 g07634(.A(new_n8010), .B(new_n8009), .Y(new_n8011));
  xor_4  g07635(.A(new_n8011), .B(new_n8008), .Y(new_n8012));
  nand_5 g07636(.A(pi134), .B(pi058), .Y(new_n8013));
  nand_5 g07637(.A(pi149), .B(pi132), .Y(new_n8014));
  nand_5 g07638(.A(pi240), .B(pi186), .Y(new_n8015));
  xor_4  g07639(.A(new_n8015), .B(new_n8014), .Y(new_n8016));
  xor_4  g07640(.A(new_n8016), .B(new_n8013), .Y(new_n8017));
  xor_4  g07641(.A(new_n8017), .B(new_n8012), .Y(new_n8018));
  nor_5  g07642(.A(new_n8018), .B(new_n8007), .Y(new_n8019));
  nand_5 g07643(.A(pi240), .B(pi058), .Y(new_n8020));
  nand_5 g07644(.A(pi186), .B(pi149), .Y(new_n8021));
  nand_5 g07645(.A(pi167), .B(pi132), .Y(new_n8022));
  xor_4  g07646(.A(new_n8022), .B(new_n8021), .Y(new_n8023));
  xor_4  g07647(.A(new_n8023), .B(new_n8020), .Y(new_n8024));
  nand_5 g07648(.A(pi211), .B(pi134), .Y(new_n8025));
  nand_5 g07649(.A(new_n8015), .B(new_n8014), .Y(new_n8026));
  nand_5 g07650(.A(new_n8016), .B(new_n8013), .Y(new_n8027));
  nand_5 g07651(.A(new_n8027), .B(new_n8026), .Y(new_n8028));
  xor_4  g07652(.A(new_n8028), .B(new_n8025), .Y(new_n8029));
  xor_4  g07653(.A(new_n8029), .B(new_n8024), .Y(new_n8030));
  nand_5 g07654(.A(pi199), .B(pi175), .Y(new_n8031));
  or_6   g07655(.A(new_n8011), .B(new_n8008), .Y(new_n8032));
  not_8  g07656(.A(new_n8017), .Y(new_n8033));
  nand_5 g07657(.A(new_n8033), .B(new_n8012), .Y(new_n8034));
  nand_5 g07658(.A(new_n8034), .B(new_n8032), .Y(new_n8035));
  xor_4  g07659(.A(new_n8035), .B(new_n8031), .Y(new_n8036));
  xor_4  g07660(.A(new_n8036), .B(new_n8030), .Y(new_n8037));
  xor_4  g07661(.A(new_n8037), .B(new_n8019), .Y(new_n8038));
  xor_4  g07662(.A(new_n8038), .B(new_n8001), .Y(new_n8039));
  xor_4  g07663(.A(new_n7997), .B(new_n7986), .Y(new_n8040));
  xor_4  g07664(.A(new_n8018), .B(new_n8007), .Y(new_n8041));
  nand_5 g07665(.A(new_n8041), .B(new_n8040), .Y(new_n8042));
  xor_4  g07666(.A(new_n8041), .B(new_n8040), .Y(new_n8043));
  xor_4  g07667(.A(new_n8005), .B(new_n4987), .Y(new_n8044));
  nand_5 g07668(.A(new_n4988), .B(new_n4982), .Y(new_n8045));
  not_8  g07669(.A(new_n4978), .Y(new_n8046));
  nand_5 g07670(.A(new_n4989), .B(new_n8046), .Y(new_n8047));
  nand_5 g07671(.A(new_n8047), .B(new_n8045), .Y(new_n8048));
  or_6   g07672(.A(new_n8048), .B(new_n8044), .Y(new_n8049));
  xor_4  g07673(.A(new_n7995), .B(new_n7993), .Y(new_n8050));
  xor_4  g07674(.A(new_n8048), .B(new_n8044), .Y(new_n8051));
  nand_5 g07675(.A(new_n8051), .B(new_n8050), .Y(new_n8052));
  nand_5 g07676(.A(new_n8052), .B(new_n8049), .Y(new_n8053));
  nand_5 g07677(.A(new_n8053), .B(new_n8043), .Y(new_n8054));
  nand_5 g07678(.A(new_n8054), .B(new_n8042), .Y(new_n8055));
  xor_4  g07679(.A(new_n8055), .B(new_n8039), .Y(new_n8056));
  nand_5 g07680(.A(pi150), .B(pi103), .Y(new_n8057));
  nand_5 g07681(.A(pi244), .B(pi103), .Y(new_n8058));
  nand_5 g07682(.A(pi029), .B(pi016), .Y(new_n8059));
  nand_5 g07683(.A(new_n8059), .B(new_n8058), .Y(new_n8060));
  nand_5 g07684(.A(pi117), .B(pi069), .Y(new_n8061));
  or_6   g07685(.A(new_n8059), .B(new_n8058), .Y(new_n8062));
  nand_5 g07686(.A(new_n8062), .B(new_n8061), .Y(new_n8063));
  nand_5 g07687(.A(new_n8063), .B(new_n8060), .Y(new_n8064));
  xor_4  g07688(.A(new_n8064), .B(new_n8057), .Y(new_n8065));
  nand_5 g07689(.A(pi069), .B(pi016), .Y(new_n8066));
  nand_5 g07690(.A(pi080), .B(pi029), .Y(new_n8067));
  nand_5 g07691(.A(pi244), .B(pi117), .Y(new_n8068));
  xor_4  g07692(.A(new_n8068), .B(new_n8067), .Y(new_n8069));
  xor_4  g07693(.A(new_n8069), .B(new_n8066), .Y(new_n8070));
  xor_4  g07694(.A(new_n8070), .B(new_n8065), .Y(new_n8071));
  not_8  g07695(.A(new_n8061), .Y(new_n8072));
  not_8  g07696(.A(new_n8060), .Y(new_n8073));
  nand_5 g07697(.A(new_n8072), .B(new_n4992), .Y(new_n8074));
  nand_5 g07698(.A(new_n8074), .B(new_n8073), .Y(new_n8075));
  nand_5 g07699(.A(new_n8075), .B(new_n8062), .Y(new_n8076));
  nand_5 g07700(.A(new_n8076), .B(new_n8072), .Y(new_n8077));
  nor_5  g07701(.A(new_n8077), .B(new_n8071), .Y(new_n8078));
  nand_5 g07702(.A(pi244), .B(pi016), .Y(new_n8079));
  nand_5 g07703(.A(pi080), .B(pi069), .Y(new_n8080));
  nand_5 g07704(.A(pi247), .B(pi029), .Y(new_n8081));
  xor_4  g07705(.A(new_n8081), .B(new_n8080), .Y(new_n8082));
  xor_4  g07706(.A(new_n8082), .B(new_n8079), .Y(new_n8083));
  nand_5 g07707(.A(pi150), .B(pi117), .Y(new_n8084));
  nand_5 g07708(.A(new_n8068), .B(new_n8067), .Y(new_n8085));
  nand_5 g07709(.A(new_n8069), .B(new_n8066), .Y(new_n8086));
  nand_5 g07710(.A(new_n8086), .B(new_n8085), .Y(new_n8087));
  xor_4  g07711(.A(new_n8087), .B(new_n8084), .Y(new_n8088));
  xnor_4 g07712(.A(new_n8088), .B(new_n8083), .Y(new_n8089));
  nand_5 g07713(.A(pi221), .B(pi103), .Y(new_n8090));
  or_6   g07714(.A(new_n8064), .B(new_n8057), .Y(new_n8091));
  not_8  g07715(.A(new_n8070), .Y(new_n8092));
  nand_5 g07716(.A(new_n8092), .B(new_n8065), .Y(new_n8093));
  nand_5 g07717(.A(new_n8093), .B(new_n8091), .Y(new_n8094));
  xor_4  g07718(.A(new_n8094), .B(new_n8090), .Y(new_n8095));
  xor_4  g07719(.A(new_n8095), .B(new_n8089), .Y(new_n8096));
  xor_4  g07720(.A(new_n8096), .B(new_n8078), .Y(new_n8097));
  xor_4  g07721(.A(new_n8077), .B(new_n8071), .Y(new_n8098));
  nor_5  g07722(.A(new_n8074), .B(new_n8073), .Y(new_n8099));
  nor_5  g07723(.A(new_n8099), .B(new_n8076), .Y(new_n8100));
  nand_5 g07724(.A(new_n4996), .B(new_n4993), .Y(new_n8101));
  nand_5 g07725(.A(new_n4997), .B(new_n4990), .Y(new_n8102));
  nand_5 g07726(.A(new_n8102), .B(new_n8101), .Y(new_n8103));
  nand_5 g07727(.A(new_n8103), .B(new_n8100), .Y(new_n8104));
  xor_4  g07728(.A(new_n8051), .B(new_n8050), .Y(new_n8105));
  xor_4  g07729(.A(new_n8103), .B(new_n8100), .Y(new_n8106));
  nand_5 g07730(.A(new_n8106), .B(new_n8105), .Y(new_n8107));
  nand_5 g07731(.A(new_n8107), .B(new_n8104), .Y(new_n8108));
  or_6   g07732(.A(new_n8108), .B(new_n8098), .Y(new_n8109));
  xor_4  g07733(.A(new_n8053), .B(new_n8043), .Y(new_n8110));
  not_8  g07734(.A(new_n8110), .Y(new_n8111));
  xor_4  g07735(.A(new_n8108), .B(new_n8098), .Y(new_n8112));
  nand_5 g07736(.A(new_n8112), .B(new_n8111), .Y(new_n8113));
  nand_5 g07737(.A(new_n8113), .B(new_n8109), .Y(new_n8114));
  xor_4  g07738(.A(new_n8114), .B(new_n8097), .Y(new_n8115));
  xor_4  g07739(.A(new_n8115), .B(new_n8056), .Y(po041));
  xor_4  g07740(.A(new_n6945), .B(new_n6943), .Y(po042));
  xor_4  g07741(.A(new_n4955), .B(new_n4953), .Y(po043));
  xor_4  g07742(.A(new_n1036), .B(new_n1019), .Y(po044));
  xor_4  g07743(.A(new_n2573), .B(new_n2543), .Y(po045));
  xor_4  g07744(.A(new_n4941), .B(new_n4925), .Y(po046));
  nand_5 g07745(.A(pi205), .B(pi107), .Y(new_n8122));
  nand_5 g07746(.A(pi253), .B(pi171), .Y(new_n8123));
  nand_5 g07747(.A(pi107), .B(pi074), .Y(new_n8124));
  nand_5 g07748(.A(new_n8124), .B(new_n8123), .Y(new_n8125));
  nand_5 g07749(.A(pi050), .B(pi049), .Y(new_n8126));
  xor_4  g07750(.A(new_n8124), .B(new_n8123), .Y(new_n8127));
  nand_5 g07751(.A(new_n8127), .B(new_n8126), .Y(new_n8128));
  nand_5 g07752(.A(new_n8128), .B(new_n8125), .Y(new_n8129));
  nand_5 g07753(.A(pi171), .B(pi074), .Y(new_n8130));
  nand_5 g07754(.A(pi109), .B(pi063), .Y(new_n8131));
  nand_5 g07755(.A(pi201), .B(pi173), .Y(new_n8132));
  nand_5 g07756(.A(new_n8132), .B(new_n8131), .Y(new_n8133));
  nand_5 g07757(.A(pi156), .B(pi014), .Y(new_n8134));
  xor_4  g07758(.A(new_n8132), .B(new_n8131), .Y(new_n8135));
  nand_5 g07759(.A(new_n8135), .B(new_n8134), .Y(new_n8136));
  nand_5 g07760(.A(new_n8136), .B(new_n8133), .Y(new_n8137));
  xor_4  g07761(.A(new_n8137), .B(new_n8130), .Y(new_n8138));
  xor_4  g07762(.A(new_n8138), .B(new_n8129), .Y(new_n8139));
  nand_5 g07763(.A(pi202), .B(pi029), .Y(new_n8140));
  nand_5 g07764(.A(pi244), .B(pi080), .Y(new_n8141));
  nand_5 g07765(.A(new_n8081), .B(new_n8080), .Y(new_n8142));
  nand_5 g07766(.A(new_n8082), .B(new_n8079), .Y(new_n8143));
  nand_5 g07767(.A(new_n8143), .B(new_n8142), .Y(new_n8144));
  xor_4  g07768(.A(new_n8144), .B(new_n8141), .Y(new_n8145));
  nand_5 g07769(.A(pi247), .B(pi069), .Y(new_n8146));
  nand_5 g07770(.A(pi234), .B(pi029), .Y(new_n8147));
  nand_5 g07771(.A(new_n8147), .B(new_n8146), .Y(new_n8148));
  nand_5 g07772(.A(pi234), .B(pi069), .Y(new_n8149));
  nor_5  g07773(.A(new_n8149), .B(new_n8081), .Y(new_n8150));
  not_8  g07774(.A(new_n8150), .Y(new_n8151));
  nand_5 g07775(.A(new_n8151), .B(new_n8148), .Y(new_n8152));
  xor_4  g07776(.A(new_n8152), .B(new_n8145), .Y(new_n8153));
  nand_5 g07777(.A(pi150), .B(pi016), .Y(new_n8154));
  nand_5 g07778(.A(pi221), .B(pi117), .Y(new_n8155));
  nand_5 g07779(.A(new_n8155), .B(new_n8154), .Y(new_n8156));
  nand_5 g07780(.A(pi221), .B(pi016), .Y(new_n8157));
  or_6   g07781(.A(new_n8157), .B(new_n8084), .Y(new_n8158));
  nand_5 g07782(.A(new_n8158), .B(new_n8156), .Y(new_n8159));
  xor_4  g07783(.A(new_n8159), .B(new_n8153), .Y(new_n8160));
  nand_5 g07784(.A(new_n8087), .B(new_n8084), .Y(new_n8161));
  nand_5 g07785(.A(new_n8088), .B(new_n8083), .Y(new_n8162));
  nand_5 g07786(.A(new_n8162), .B(new_n8161), .Y(new_n8163));
  xor_4  g07787(.A(new_n8163), .B(new_n8160), .Y(new_n8164));
  not_8  g07788(.A(new_n8090), .Y(new_n8165));
  nor_5  g07789(.A(new_n8094), .B(new_n8165), .Y(new_n8166));
  nor_5  g07790(.A(new_n8095), .B(new_n8089), .Y(new_n8167));
  nor_5  g07791(.A(new_n8167), .B(new_n8166), .Y(new_n8168));
  not_8  g07792(.A(new_n8168), .Y(new_n8169));
  nor_5  g07793(.A(new_n8169), .B(new_n8164), .Y(new_n8170));
  nand_5 g07794(.A(pi247), .B(pi244), .Y(new_n8171));
  nand_5 g07795(.A(pi214), .B(pi029), .Y(new_n8172));
  xor_4  g07796(.A(new_n8172), .B(new_n8149), .Y(new_n8173));
  xor_4  g07797(.A(new_n8173), .B(new_n8171), .Y(new_n8174));
  nand_5 g07798(.A(pi150), .B(pi080), .Y(new_n8175));
  xor_4  g07799(.A(new_n8175), .B(new_n8151), .Y(new_n8176));
  not_8  g07800(.A(new_n8176), .Y(new_n8177));
  xor_4  g07801(.A(new_n8177), .B(new_n8174), .Y(new_n8178));
  nand_5 g07802(.A(pi196), .B(pi117), .Y(new_n8179));
  nand_5 g07803(.A(pi184), .B(pi103), .Y(new_n8180));
  xor_4  g07804(.A(new_n8180), .B(new_n8179), .Y(new_n8181));
  xor_4  g07805(.A(new_n8181), .B(new_n8157), .Y(new_n8182));
  nand_5 g07806(.A(new_n8144), .B(new_n8141), .Y(new_n8183));
  nand_5 g07807(.A(new_n8152), .B(new_n8145), .Y(new_n8184));
  nand_5 g07808(.A(new_n8184), .B(new_n8183), .Y(new_n8185));
  xor_4  g07809(.A(new_n8185), .B(new_n8182), .Y(new_n8186));
  xor_4  g07810(.A(new_n8186), .B(new_n8178), .Y(new_n8187));
  nand_5 g07811(.A(new_n8159), .B(new_n8153), .Y(new_n8188));
  nand_5 g07812(.A(new_n8163), .B(new_n8160), .Y(new_n8189));
  nand_5 g07813(.A(new_n8189), .B(new_n8188), .Y(new_n8190));
  xor_4  g07814(.A(new_n8190), .B(new_n8158), .Y(new_n8191));
  xor_4  g07815(.A(new_n8191), .B(new_n8187), .Y(new_n8192));
  nand_5 g07816(.A(new_n8192), .B(new_n8170), .Y(new_n8193));
  xor_4  g07817(.A(new_n8192), .B(new_n8170), .Y(new_n8194));
  nand_5 g07818(.A(pi196), .B(pi103), .Y(new_n8195));
  xor_4  g07819(.A(new_n8168), .B(new_n8164), .Y(new_n8196));
  or_6   g07820(.A(new_n8196), .B(new_n8195), .Y(new_n8197));
  not_8  g07821(.A(new_n8078), .Y(new_n8198));
  nor_5  g07822(.A(new_n8096), .B(new_n8198), .Y(new_n8199));
  xor_4  g07823(.A(new_n8196), .B(new_n8195), .Y(new_n8200));
  nand_5 g07824(.A(new_n8200), .B(new_n8199), .Y(new_n8201));
  nand_5 g07825(.A(new_n8201), .B(new_n8197), .Y(new_n8202));
  nand_5 g07826(.A(new_n8202), .B(new_n8194), .Y(new_n8203));
  nand_5 g07827(.A(new_n8203), .B(new_n8193), .Y(new_n8204));
  xor_4  g07828(.A(new_n8204), .B(new_n8140), .Y(new_n8205));
  nand_5 g07829(.A(pi103), .B(pi010), .Y(new_n8206));
  xor_4  g07830(.A(new_n8206), .B(new_n8205), .Y(new_n8207));
  or_6   g07831(.A(new_n8190), .B(new_n8158), .Y(new_n8208));
  nand_5 g07832(.A(new_n8191), .B(new_n8187), .Y(new_n8209));
  nand_5 g07833(.A(new_n8209), .B(new_n8208), .Y(new_n8210));
  nand_5 g07834(.A(pi253), .B(pi049), .Y(new_n8211));
  nand_5 g07835(.A(pi245), .B(pi230), .Y(new_n8212));
  or_6   g07836(.A(new_n8134), .B(new_n7965), .Y(new_n8213));
  or_6   g07837(.A(new_n8213), .B(new_n8212), .Y(new_n8214));
  xor_4  g07838(.A(new_n8135), .B(new_n8134), .Y(new_n8215));
  not_8  g07839(.A(new_n8215), .Y(new_n8216));
  xor_4  g07840(.A(new_n8213), .B(new_n8212), .Y(new_n8217));
  nand_5 g07841(.A(new_n8217), .B(new_n8216), .Y(new_n8218));
  nand_5 g07842(.A(new_n8218), .B(new_n8214), .Y(new_n8219));
  xor_4  g07843(.A(new_n8219), .B(new_n8211), .Y(new_n8220));
  xor_4  g07844(.A(new_n8220), .B(new_n8210), .Y(new_n8221));
  xor_4  g07845(.A(new_n8221), .B(new_n8207), .Y(new_n8222));
  xor_4  g07846(.A(new_n8202), .B(new_n8194), .Y(new_n8223));
  not_8  g07847(.A(new_n8223), .Y(new_n8224));
  nand_5 g07848(.A(new_n8037), .B(new_n8019), .Y(new_n8225));
  nand_5 g07849(.A(pi195), .B(pi175), .Y(new_n8226));
  nand_5 g07850(.A(new_n8226), .B(new_n8225), .Y(new_n8227));
  nand_5 g07851(.A(pi149), .B(pi058), .Y(new_n8228));
  nand_5 g07852(.A(new_n8022), .B(new_n8021), .Y(new_n8229));
  nand_5 g07853(.A(new_n8023), .B(new_n8020), .Y(new_n8230));
  nand_5 g07854(.A(new_n8230), .B(new_n8229), .Y(new_n8231));
  xor_4  g07855(.A(new_n8231), .B(new_n8228), .Y(new_n8232));
  nand_5 g07856(.A(pi186), .B(pi167), .Y(new_n8233));
  nand_5 g07857(.A(pi181), .B(pi132), .Y(new_n8234));
  nand_5 g07858(.A(new_n8234), .B(new_n8233), .Y(new_n8235));
  nand_5 g07859(.A(pi186), .B(pi181), .Y(new_n8236));
  nor_5  g07860(.A(new_n8236), .B(new_n8022), .Y(new_n8237));
  not_8  g07861(.A(new_n8237), .Y(new_n8238));
  nand_5 g07862(.A(new_n8238), .B(new_n8235), .Y(new_n8239));
  xor_4  g07863(.A(new_n8239), .B(new_n8232), .Y(new_n8240));
  nand_5 g07864(.A(pi240), .B(pi211), .Y(new_n8241));
  nand_5 g07865(.A(pi199), .B(pi134), .Y(new_n8242));
  and_6  g07866(.A(new_n8242), .B(new_n8241), .Y(new_n8243));
  nand_5 g07867(.A(pi240), .B(pi199), .Y(new_n8244));
  nor_5  g07868(.A(new_n8244), .B(new_n8025), .Y(new_n8245));
  or_6   g07869(.A(new_n8245), .B(new_n8243), .Y(new_n8246));
  xnor_4 g07870(.A(new_n8246), .B(new_n8240), .Y(new_n8247));
  nand_5 g07871(.A(new_n8028), .B(new_n8025), .Y(new_n8248));
  nand_5 g07872(.A(new_n8029), .B(new_n8024), .Y(new_n8249));
  nand_5 g07873(.A(new_n8249), .B(new_n8248), .Y(new_n8250));
  xor_4  g07874(.A(new_n8250), .B(new_n8247), .Y(new_n8251));
  not_8  g07875(.A(new_n8031), .Y(new_n8252));
  nand_5 g07876(.A(new_n8035), .B(new_n8252), .Y(new_n8253));
  or_6   g07877(.A(new_n8036), .B(new_n8030), .Y(new_n8254));
  nand_5 g07878(.A(new_n8254), .B(new_n8253), .Y(new_n8255));
  xor_4  g07879(.A(new_n8255), .B(new_n8251), .Y(new_n8256));
  not_8  g07880(.A(new_n8256), .Y(new_n8257));
  xor_4  g07881(.A(new_n8226), .B(new_n8225), .Y(new_n8258));
  nand_5 g07882(.A(new_n8258), .B(new_n8257), .Y(new_n8259));
  nand_5 g07883(.A(new_n8259), .B(new_n8227), .Y(new_n8260));
  nand_5 g07884(.A(new_n8255), .B(new_n8251), .Y(new_n8261));
  nand_5 g07885(.A(pi200), .B(pi132), .Y(new_n8262));
  nand_5 g07886(.A(pi167), .B(pi058), .Y(new_n8263));
  xor_4  g07887(.A(new_n8263), .B(new_n8262), .Y(new_n8264));
  xor_4  g07888(.A(new_n8264), .B(new_n8236), .Y(new_n8265));
  nand_5 g07889(.A(pi211), .B(pi149), .Y(new_n8266));
  xor_4  g07890(.A(new_n8266), .B(new_n8238), .Y(new_n8267));
  not_8  g07891(.A(new_n8267), .Y(new_n8268));
  xor_4  g07892(.A(new_n8268), .B(new_n8265), .Y(new_n8269));
  nand_5 g07893(.A(pi195), .B(pi134), .Y(new_n8270));
  nand_5 g07894(.A(pi218), .B(pi175), .Y(new_n8271));
  xor_4  g07895(.A(new_n8271), .B(new_n8270), .Y(new_n8272));
  xor_4  g07896(.A(new_n8272), .B(new_n8244), .Y(new_n8273));
  nand_5 g07897(.A(new_n8231), .B(new_n8228), .Y(new_n8274));
  nand_5 g07898(.A(new_n8239), .B(new_n8232), .Y(new_n8275));
  nand_5 g07899(.A(new_n8275), .B(new_n8274), .Y(new_n8276));
  xor_4  g07900(.A(new_n8276), .B(new_n8273), .Y(new_n8277));
  xor_4  g07901(.A(new_n8277), .B(new_n8269), .Y(new_n8278));
  nor_5  g07902(.A(new_n8246), .B(new_n8240), .Y(new_n8279));
  nor_5  g07903(.A(new_n8250), .B(new_n8247), .Y(new_n8280));
  xor_4  g07904(.A(new_n8280), .B(new_n8245), .Y(new_n8281));
  nor_5  g07905(.A(new_n8281), .B(new_n8279), .Y(new_n8282));
  xor_4  g07906(.A(new_n8282), .B(new_n8278), .Y(new_n8283));
  xor_4  g07907(.A(new_n8283), .B(new_n8261), .Y(new_n8284));
  xor_4  g07908(.A(new_n8284), .B(new_n8260), .Y(new_n8285));
  nand_5 g07909(.A(pi245), .B(pi173), .Y(new_n8286));
  nand_5 g07910(.A(pi201), .B(pi014), .Y(new_n8287));
  nand_5 g07911(.A(pi156), .B(pi109), .Y(new_n8288));
  nand_5 g07912(.A(new_n8288), .B(new_n8287), .Y(new_n8289));
  nand_5 g07913(.A(new_n8289), .B(new_n8213), .Y(new_n8290));
  xor_4  g07914(.A(new_n8290), .B(new_n8286), .Y(new_n8291));
  nand_5 g07915(.A(new_n7965), .B(new_n7964), .Y(new_n8292));
  nand_5 g07916(.A(new_n7966), .B(new_n7963), .Y(new_n8293));
  nand_5 g07917(.A(new_n8293), .B(new_n8292), .Y(new_n8294));
  xor_4  g07918(.A(new_n8294), .B(new_n8291), .Y(new_n8295));
  nand_5 g07919(.A(pi230), .B(pi049), .Y(new_n8296));
  nand_5 g07920(.A(pi171), .B(pi050), .Y(new_n8297));
  and_6  g07921(.A(new_n8297), .B(new_n8296), .Y(new_n8298));
  nor_5  g07922(.A(new_n8126), .B(new_n7968), .Y(new_n8299));
  or_6   g07923(.A(new_n8299), .B(new_n8298), .Y(new_n8300));
  xnor_4 g07924(.A(new_n8300), .B(new_n8295), .Y(new_n8301));
  nand_5 g07925(.A(new_n7971), .B(new_n7968), .Y(new_n8302));
  nand_5 g07926(.A(new_n7972), .B(new_n7967), .Y(new_n8303));
  nand_5 g07927(.A(new_n8303), .B(new_n8302), .Y(new_n8304));
  xor_4  g07928(.A(new_n8304), .B(new_n8301), .Y(new_n8305));
  or_6   g07929(.A(new_n7977), .B(new_n7974), .Y(new_n8306));
  nand_5 g07930(.A(new_n7978), .B(new_n7973), .Y(new_n8307));
  nand_5 g07931(.A(new_n8307), .B(new_n8306), .Y(new_n8308));
  nand_5 g07932(.A(new_n8308), .B(new_n8305), .Y(new_n8309));
  xor_4  g07933(.A(new_n8217), .B(new_n8215), .Y(new_n8310));
  xor_4  g07934(.A(new_n8127), .B(new_n8126), .Y(new_n8311));
  nand_5 g07935(.A(new_n8290), .B(new_n8286), .Y(new_n8312));
  nand_5 g07936(.A(new_n8294), .B(new_n8291), .Y(new_n8313));
  nand_5 g07937(.A(new_n8313), .B(new_n8312), .Y(new_n8314));
  xor_4  g07938(.A(new_n8314), .B(new_n8311), .Y(new_n8315));
  xnor_4 g07939(.A(new_n8315), .B(new_n8310), .Y(new_n8316));
  nor_5  g07940(.A(new_n8300), .B(new_n8295), .Y(new_n8317));
  nor_5  g07941(.A(new_n8304), .B(new_n8301), .Y(new_n8318));
  xor_4  g07942(.A(new_n8318), .B(new_n8299), .Y(new_n8319));
  nor_5  g07943(.A(new_n8319), .B(new_n8317), .Y(new_n8320));
  xor_4  g07944(.A(new_n8320), .B(new_n8316), .Y(new_n8321));
  xnor_4 g07945(.A(new_n8321), .B(new_n8309), .Y(new_n8322));
  nand_5 g07946(.A(new_n7979), .B(new_n7962), .Y(new_n8323));
  nand_5 g07947(.A(pi253), .B(pi107), .Y(new_n8324));
  nand_5 g07948(.A(new_n8324), .B(new_n8323), .Y(new_n8325));
  xnor_4 g07949(.A(new_n8308), .B(new_n8305), .Y(new_n8326));
  xor_4  g07950(.A(new_n8324), .B(new_n8323), .Y(new_n8327));
  nand_5 g07951(.A(new_n8327), .B(new_n8326), .Y(new_n8328));
  nand_5 g07952(.A(new_n8328), .B(new_n8325), .Y(new_n8329));
  xnor_4 g07953(.A(new_n8329), .B(new_n8322), .Y(new_n8330));
  nor_5  g07954(.A(new_n7944), .B(new_n7927), .Y(new_n8331));
  not_8  g07955(.A(new_n8331), .Y(new_n8332));
  nand_5 g07956(.A(pi163), .B(pi025), .Y(new_n8333));
  nand_5 g07957(.A(new_n8333), .B(new_n8332), .Y(new_n8334));
  nand_5 g07958(.A(pi066), .B(pi039), .Y(new_n8335));
  nand_5 g07959(.A(pi207), .B(pi116), .Y(new_n8336));
  nand_5 g07960(.A(pi226), .B(pi070), .Y(new_n8337));
  nand_5 g07961(.A(new_n8337), .B(new_n8336), .Y(new_n8338));
  nand_5 g07962(.A(pi207), .B(pi070), .Y(new_n8339));
  or_6   g07963(.A(new_n8339), .B(new_n7933), .Y(new_n8340));
  nand_5 g07964(.A(new_n8340), .B(new_n8338), .Y(new_n8341));
  xor_4  g07965(.A(new_n8341), .B(new_n8335), .Y(new_n8342));
  nand_5 g07966(.A(new_n7935), .B(new_n7934), .Y(new_n8343));
  nand_5 g07967(.A(new_n7936), .B(new_n7933), .Y(new_n8344));
  nand_5 g07968(.A(new_n8344), .B(new_n8343), .Y(new_n8345));
  xor_4  g07969(.A(new_n8345), .B(new_n8342), .Y(new_n8346));
  nand_5 g07970(.A(new_n7941), .B(new_n7938), .Y(new_n8347));
  nand_5 g07971(.A(new_n7942), .B(new_n7937), .Y(new_n8348));
  nand_5 g07972(.A(new_n8348), .B(new_n8347), .Y(new_n8349));
  nand_5 g07973(.A(pi228), .B(pi055), .Y(new_n8350));
  nand_5 g07974(.A(pi148), .B(pi002), .Y(new_n8351));
  nand_5 g07975(.A(new_n8351), .B(new_n8350), .Y(new_n8352));
  nand_5 g07976(.A(pi228), .B(pi002), .Y(new_n8353));
  or_6   g07977(.A(new_n8353), .B(new_n7938), .Y(new_n8354));
  nand_5 g07978(.A(new_n8354), .B(new_n8352), .Y(new_n8355));
  xor_4  g07979(.A(new_n8355), .B(new_n8349), .Y(new_n8356));
  xor_4  g07980(.A(new_n8356), .B(new_n8346), .Y(new_n8357));
  or_6   g07981(.A(new_n7931), .B(new_n7928), .Y(new_n8358));
  nand_5 g07982(.A(new_n7943), .B(new_n7932), .Y(new_n8359));
  nand_5 g07983(.A(new_n8359), .B(new_n8358), .Y(new_n8360));
  xor_4  g07984(.A(new_n8360), .B(new_n8357), .Y(new_n8361));
  xor_4  g07985(.A(new_n8333), .B(new_n8332), .Y(new_n8362));
  nand_5 g07986(.A(new_n8362), .B(new_n8361), .Y(new_n8363));
  nand_5 g07987(.A(new_n8363), .B(new_n8334), .Y(new_n8364));
  not_8  g07988(.A(new_n8357), .Y(new_n8365));
  nand_5 g07989(.A(new_n8360), .B(new_n8365), .Y(new_n8366));
  nand_5 g07990(.A(pi226), .B(pi115), .Y(new_n8367));
  nand_5 g07991(.A(pi116), .B(pi066), .Y(new_n8368));
  xor_4  g07992(.A(new_n8368), .B(new_n8367), .Y(new_n8369));
  xor_4  g07993(.A(new_n8369), .B(new_n8339), .Y(new_n8370));
  not_8  g07994(.A(new_n8370), .Y(new_n8371));
  nand_5 g07995(.A(pi055), .B(pi039), .Y(new_n8372));
  xor_4  g07996(.A(new_n8372), .B(new_n8340), .Y(new_n8373));
  xor_4  g07997(.A(new_n8373), .B(new_n8371), .Y(new_n8374));
  nand_5 g07998(.A(pi239), .B(pi163), .Y(new_n8375));
  nand_5 g07999(.A(pi148), .B(pi025), .Y(new_n8376));
  xor_4  g08000(.A(new_n8376), .B(new_n8375), .Y(new_n8377));
  xor_4  g08001(.A(new_n8377), .B(new_n8353), .Y(new_n8378));
  nand_5 g08002(.A(new_n8341), .B(new_n8335), .Y(new_n8379));
  nand_5 g08003(.A(new_n8345), .B(new_n8342), .Y(new_n8380));
  nand_5 g08004(.A(new_n8380), .B(new_n8379), .Y(new_n8381));
  xor_4  g08005(.A(new_n8381), .B(new_n8378), .Y(new_n8382));
  xor_4  g08006(.A(new_n8382), .B(new_n8374), .Y(new_n8383));
  nand_5 g08007(.A(new_n8355), .B(new_n8349), .Y(new_n8384));
  nand_5 g08008(.A(new_n8356), .B(new_n8346), .Y(new_n8385));
  nand_5 g08009(.A(new_n8385), .B(new_n8384), .Y(new_n8386));
  xor_4  g08010(.A(new_n8386), .B(new_n8354), .Y(new_n8387));
  xnor_4 g08011(.A(new_n8387), .B(new_n8383), .Y(new_n8388));
  xor_4  g08012(.A(new_n8388), .B(new_n8366), .Y(new_n8389));
  xor_4  g08013(.A(new_n8389), .B(new_n8364), .Y(new_n8390));
  xor_4  g08014(.A(new_n8390), .B(new_n8330), .Y(new_n8391));
  xnor_4 g08015(.A(new_n8362), .B(new_n8361), .Y(new_n8392));
  nand_5 g08016(.A(new_n7980), .B(new_n7945), .Y(new_n8393));
  nand_5 g08017(.A(new_n8000), .B(new_n7981), .Y(new_n8394));
  nand_5 g08018(.A(new_n8394), .B(new_n8393), .Y(new_n8395));
  nand_5 g08019(.A(new_n8395), .B(new_n8392), .Y(new_n8396));
  xnor_4 g08020(.A(new_n8327), .B(new_n8326), .Y(new_n8397));
  xor_4  g08021(.A(new_n8395), .B(new_n8392), .Y(new_n8398));
  nand_5 g08022(.A(new_n8398), .B(new_n8397), .Y(new_n8399));
  nand_5 g08023(.A(new_n8399), .B(new_n8396), .Y(new_n8400));
  xor_4  g08024(.A(new_n8400), .B(new_n8391), .Y(new_n8401));
  xor_4  g08025(.A(new_n8258), .B(new_n8256), .Y(new_n8402));
  nand_5 g08026(.A(new_n8038), .B(new_n8001), .Y(new_n8403));
  nand_5 g08027(.A(new_n8055), .B(new_n8039), .Y(new_n8404));
  nand_5 g08028(.A(new_n8404), .B(new_n8403), .Y(new_n8405));
  nand_5 g08029(.A(new_n8405), .B(new_n8402), .Y(new_n8406));
  xor_4  g08030(.A(new_n8398), .B(new_n8397), .Y(new_n8407));
  xor_4  g08031(.A(new_n8405), .B(new_n8402), .Y(new_n8408));
  nand_5 g08032(.A(new_n8408), .B(new_n8407), .Y(new_n8409));
  nand_5 g08033(.A(new_n8409), .B(new_n8406), .Y(new_n8410));
  xor_4  g08034(.A(new_n8410), .B(new_n8401), .Y(new_n8411));
  xor_4  g08035(.A(new_n8411), .B(new_n8285), .Y(new_n8412));
  nor_5  g08036(.A(new_n8412), .B(new_n8224), .Y(new_n8413));
  xor_4  g08037(.A(new_n8412), .B(new_n8223), .Y(new_n8414));
  xnor_4 g08038(.A(new_n8200), .B(new_n8199), .Y(new_n8415));
  nand_5 g08039(.A(new_n8114), .B(new_n8097), .Y(new_n8416));
  not_8  g08040(.A(new_n8056), .Y(new_n8417));
  nand_5 g08041(.A(new_n8115), .B(new_n8417), .Y(new_n8418));
  nand_5 g08042(.A(new_n8418), .B(new_n8416), .Y(new_n8419));
  nand_5 g08043(.A(new_n8419), .B(new_n8415), .Y(new_n8420));
  xor_4  g08044(.A(new_n8408), .B(new_n8407), .Y(new_n8421));
  not_8  g08045(.A(new_n8421), .Y(new_n8422));
  xor_4  g08046(.A(new_n8419), .B(new_n8415), .Y(new_n8423));
  nand_5 g08047(.A(new_n8423), .B(new_n8422), .Y(new_n8424));
  nand_5 g08048(.A(new_n8424), .B(new_n8420), .Y(new_n8425));
  nor_5  g08049(.A(new_n8425), .B(new_n8414), .Y(new_n8426));
  nor_5  g08050(.A(new_n8426), .B(new_n8413), .Y(new_n8427));
  nand_5 g08051(.A(new_n8314), .B(new_n8311), .Y(new_n8428));
  nand_5 g08052(.A(new_n8315), .B(new_n8310), .Y(new_n8429));
  nand_5 g08053(.A(new_n8429), .B(new_n8428), .Y(new_n8430));
  xor_4  g08054(.A(new_n8430), .B(new_n8427), .Y(new_n8431));
  xor_4  g08055(.A(new_n8431), .B(new_n8222), .Y(new_n8432));
  xor_4  g08056(.A(new_n8432), .B(new_n8139), .Y(new_n8433));
  xor_4  g08057(.A(new_n8433), .B(new_n8122), .Y(new_n8434));
  nand_5 g08058(.A(pi063), .B(pi014), .Y(new_n8435));
  nand_5 g08059(.A(pi173), .B(pi156), .Y(new_n8436));
  xor_4  g08060(.A(new_n8436), .B(new_n8435), .Y(new_n8437));
  nand_5 g08061(.A(new_n8381), .B(new_n8378), .Y(new_n8438));
  not_8  g08062(.A(new_n8374), .Y(new_n8439));
  nand_5 g08063(.A(new_n8382), .B(new_n8439), .Y(new_n8440));
  nand_5 g08064(.A(new_n8440), .B(new_n8438), .Y(new_n8441));
  nand_5 g08065(.A(pi116), .B(pi055), .Y(new_n8442));
  xor_4  g08066(.A(new_n8442), .B(new_n8441), .Y(new_n8443));
  nand_5 g08067(.A(new_n8368), .B(new_n8367), .Y(new_n8444));
  nand_5 g08068(.A(new_n8369), .B(new_n8339), .Y(new_n8445));
  nand_5 g08069(.A(new_n8445), .B(new_n8444), .Y(new_n8446));
  nand_5 g08070(.A(new_n8376), .B(new_n8375), .Y(new_n8447));
  nand_5 g08071(.A(new_n8377), .B(new_n8353), .Y(new_n8448));
  nand_5 g08072(.A(new_n8448), .B(new_n8447), .Y(new_n8449));
  nand_5 g08073(.A(pi039), .B(pi002), .Y(new_n8450));
  xor_4  g08074(.A(new_n8450), .B(new_n8449), .Y(new_n8451));
  xor_4  g08075(.A(new_n8451), .B(new_n8446), .Y(new_n8452));
  or_6   g08076(.A(new_n8372), .B(new_n8340), .Y(new_n8453));
  nand_5 g08077(.A(new_n8373), .B(new_n8371), .Y(new_n8454));
  nand_5 g08078(.A(new_n8454), .B(new_n8453), .Y(new_n8455));
  nand_5 g08079(.A(pi239), .B(pi148), .Y(new_n8456));
  nand_5 g08080(.A(pi228), .B(pi025), .Y(new_n8457));
  xnor_4 g08081(.A(new_n8457), .B(new_n8456), .Y(new_n8458));
  xor_4  g08082(.A(new_n8458), .B(new_n8455), .Y(new_n8459));
  xor_4  g08083(.A(new_n8459), .B(new_n8452), .Y(new_n8460));
  xor_4  g08084(.A(new_n8460), .B(new_n8443), .Y(new_n8461));
  xor_4  g08085(.A(new_n8461), .B(new_n8437), .Y(new_n8462));
  nor_5  g08086(.A(new_n8321), .B(new_n8309), .Y(new_n8463));
  nor_5  g08087(.A(new_n8329), .B(new_n8322), .Y(new_n8464));
  nor_5  g08088(.A(new_n8464), .B(new_n8463), .Y(new_n8465));
  nand_5 g08089(.A(pi109), .B(pi083), .Y(new_n8466));
  xor_4  g08090(.A(new_n8466), .B(new_n8465), .Y(new_n8467));
  xor_4  g08091(.A(new_n8467), .B(new_n8462), .Y(new_n8468));
  nand_5 g08092(.A(new_n8318), .B(new_n8299), .Y(new_n8469));
  not_8  g08093(.A(new_n8320), .Y(new_n8470));
  nand_5 g08094(.A(new_n8470), .B(new_n8316), .Y(new_n8471));
  nand_5 g08095(.A(new_n8471), .B(new_n8469), .Y(new_n8472));
  nand_5 g08096(.A(pi230), .B(pi201), .Y(new_n8473));
  nand_5 g08097(.A(pi245), .B(pi050), .Y(new_n8474));
  xor_4  g08098(.A(new_n8474), .B(new_n8473), .Y(new_n8475));
  xor_4  g08099(.A(new_n8475), .B(new_n8472), .Y(new_n8476));
  xor_4  g08100(.A(new_n8476), .B(new_n8468), .Y(new_n8477));
  xor_4  g08101(.A(new_n8477), .B(new_n8434), .Y(new_n8478));
  nand_5 g08102(.A(pi200), .B(pi186), .Y(new_n8479));
  nand_5 g08103(.A(pi203), .B(pi132), .Y(new_n8480));
  nand_5 g08104(.A(new_n8280), .B(new_n8245), .Y(new_n8481));
  not_8  g08105(.A(new_n8282), .Y(new_n8482));
  nand_5 g08106(.A(new_n8482), .B(new_n8278), .Y(new_n8483));
  nand_5 g08107(.A(new_n8483), .B(new_n8481), .Y(new_n8484));
  xor_4  g08108(.A(new_n8484), .B(new_n8480), .Y(new_n8485));
  nand_5 g08109(.A(pi175), .B(pi037), .Y(new_n8486));
  nand_5 g08110(.A(new_n8283), .B(new_n8261), .Y(new_n8487));
  nand_5 g08111(.A(new_n8284), .B(new_n8260), .Y(new_n8488));
  nand_5 g08112(.A(new_n8488), .B(new_n8487), .Y(new_n8489));
  xor_4  g08113(.A(new_n8489), .B(new_n8486), .Y(new_n8490));
  xor_4  g08114(.A(new_n8490), .B(new_n8485), .Y(new_n8491));
  xor_4  g08115(.A(new_n8491), .B(new_n8479), .Y(new_n8492));
  nand_5 g08116(.A(new_n8172), .B(new_n8149), .Y(new_n8493));
  nand_5 g08117(.A(new_n8173), .B(new_n8171), .Y(new_n8494));
  nand_5 g08118(.A(new_n8494), .B(new_n8493), .Y(new_n8495));
  nor_5  g08119(.A(new_n8175), .B(new_n8151), .Y(new_n8496));
  nor_5  g08120(.A(new_n8177), .B(new_n8174), .Y(new_n8497));
  or_6   g08121(.A(new_n8497), .B(new_n8496), .Y(new_n8498));
  xor_4  g08122(.A(new_n8498), .B(new_n8495), .Y(new_n8499));
  xor_4  g08123(.A(new_n8499), .B(new_n8492), .Y(new_n8500));
  xor_4  g08124(.A(new_n8500), .B(new_n8478), .Y(new_n8501));
  or_6   g08125(.A(new_n8386), .B(new_n8354), .Y(new_n8502));
  nand_5 g08126(.A(new_n8387), .B(new_n8383), .Y(new_n8503));
  nand_5 g08127(.A(new_n8503), .B(new_n8502), .Y(new_n8504));
  nand_5 g08128(.A(new_n8388), .B(new_n8366), .Y(new_n8505));
  nand_5 g08129(.A(new_n8389), .B(new_n8364), .Y(new_n8506));
  nand_5 g08130(.A(new_n8506), .B(new_n8505), .Y(new_n8507));
  xor_4  g08131(.A(new_n8507), .B(new_n8504), .Y(new_n8508));
  nand_5 g08132(.A(pi199), .B(pi149), .Y(new_n8509));
  nand_5 g08133(.A(pi240), .B(pi195), .Y(new_n8510));
  xor_4  g08134(.A(new_n8510), .B(new_n8509), .Y(new_n8511));
  nand_5 g08135(.A(pi211), .B(pi167), .Y(new_n8512));
  nand_5 g08136(.A(new_n8276), .B(new_n8273), .Y(new_n8513));
  not_8  g08137(.A(new_n8269), .Y(new_n8514));
  nand_5 g08138(.A(new_n8277), .B(new_n8514), .Y(new_n8515));
  nand_5 g08139(.A(new_n8515), .B(new_n8513), .Y(new_n8516));
  xnor_4 g08140(.A(new_n8516), .B(new_n8512), .Y(new_n8517));
  xor_4  g08141(.A(new_n8517), .B(new_n8511), .Y(new_n8518));
  xor_4  g08142(.A(new_n8518), .B(new_n8508), .Y(new_n8519));
  nand_5 g08143(.A(new_n8263), .B(new_n8262), .Y(new_n8520));
  nand_5 g08144(.A(new_n8264), .B(new_n8236), .Y(new_n8521));
  nand_5 g08145(.A(new_n8521), .B(new_n8520), .Y(new_n8522));
  nand_5 g08146(.A(pi218), .B(pi134), .Y(new_n8523));
  nand_5 g08147(.A(new_n8271), .B(new_n8270), .Y(new_n8524));
  nand_5 g08148(.A(new_n8272), .B(new_n8244), .Y(new_n8525));
  nand_5 g08149(.A(new_n8525), .B(new_n8524), .Y(new_n8526));
  xor_4  g08150(.A(new_n8526), .B(new_n8523), .Y(new_n8527));
  xor_4  g08151(.A(new_n8527), .B(new_n8522), .Y(new_n8528));
  nor_5  g08152(.A(new_n8266), .B(new_n8238), .Y(new_n8529));
  nor_5  g08153(.A(new_n8268), .B(new_n8265), .Y(new_n8530));
  or_6   g08154(.A(new_n8530), .B(new_n8529), .Y(new_n8531));
  nand_5 g08155(.A(pi181), .B(pi058), .Y(new_n8532));
  xor_4  g08156(.A(new_n8532), .B(new_n8531), .Y(new_n8533));
  xor_4  g08157(.A(new_n8533), .B(new_n8528), .Y(new_n8534));
  xor_4  g08158(.A(new_n8534), .B(new_n8519), .Y(new_n8535));
  nand_5 g08159(.A(pi214), .B(pi069), .Y(new_n8536));
  nand_5 g08160(.A(pi247), .B(pi150), .Y(new_n8537));
  xor_4  g08161(.A(new_n8537), .B(new_n8536), .Y(new_n8538));
  xor_4  g08162(.A(new_n8538), .B(new_n8535), .Y(new_n8539));
  or_6   g08163(.A(new_n8410), .B(new_n8401), .Y(new_n8540));
  nand_5 g08164(.A(new_n8411), .B(new_n8285), .Y(new_n8541));
  nand_5 g08165(.A(new_n8541), .B(new_n8540), .Y(new_n8542));
  nand_5 g08166(.A(new_n8185), .B(new_n8182), .Y(new_n8543));
  not_8  g08167(.A(new_n8178), .Y(new_n8544));
  nand_5 g08168(.A(new_n8186), .B(new_n8544), .Y(new_n8545));
  nand_5 g08169(.A(new_n8545), .B(new_n8543), .Y(new_n8546));
  nand_5 g08170(.A(new_n8180), .B(new_n8179), .Y(new_n8547));
  nand_5 g08171(.A(new_n8181), .B(new_n8157), .Y(new_n8548));
  nand_5 g08172(.A(new_n8548), .B(new_n8547), .Y(new_n8549));
  xor_4  g08173(.A(new_n8549), .B(new_n8546), .Y(new_n8550));
  nand_5 g08174(.A(pi221), .B(pi080), .Y(new_n8551));
  xor_4  g08175(.A(new_n8551), .B(new_n8550), .Y(new_n8552));
  xor_4  g08176(.A(new_n8552), .B(new_n8542), .Y(new_n8553));
  xor_4  g08177(.A(new_n8553), .B(new_n8539), .Y(new_n8554));
  nand_5 g08178(.A(pi226), .B(pi000), .Y(new_n8555));
  nand_5 g08179(.A(pi207), .B(pi115), .Y(new_n8556));
  nand_5 g08180(.A(pi070), .B(pi066), .Y(new_n8557));
  xor_4  g08181(.A(new_n8557), .B(new_n8556), .Y(new_n8558));
  nand_5 g08182(.A(pi243), .B(pi163), .Y(new_n8559));
  nand_5 g08183(.A(new_n8390), .B(new_n8330), .Y(new_n8560));
  not_8  g08184(.A(new_n8391), .Y(new_n8561));
  or_6   g08185(.A(new_n8400), .B(new_n8561), .Y(new_n8562));
  nand_5 g08186(.A(new_n8562), .B(new_n8560), .Y(new_n8563));
  xor_4  g08187(.A(new_n8563), .B(new_n8559), .Y(new_n8564));
  xor_4  g08188(.A(new_n8564), .B(new_n8558), .Y(new_n8565));
  xor_4  g08189(.A(new_n8565), .B(new_n8555), .Y(new_n8566));
  nand_5 g08190(.A(pi244), .B(pi234), .Y(new_n8567));
  nand_5 g08191(.A(pi184), .B(pi117), .Y(new_n8568));
  nand_5 g08192(.A(pi196), .B(pi016), .Y(new_n8569));
  xor_4  g08193(.A(new_n8569), .B(new_n8568), .Y(new_n8570));
  xor_4  g08194(.A(new_n8570), .B(new_n8567), .Y(new_n8571));
  xor_4  g08195(.A(new_n8571), .B(new_n8566), .Y(new_n8572));
  xor_4  g08196(.A(new_n8572), .B(new_n8554), .Y(new_n8573));
  xor_4  g08197(.A(new_n8573), .B(new_n8501), .Y(po047));
  xnor_4 g08198(.A(new_n4808), .B(new_n4794), .Y(po048));
  xor_4  g08199(.A(new_n3095), .B(new_n3094), .Y(po049));
  nor_5  g08200(.A(new_n1104), .B(new_n1097), .Y(new_n8577));
  nand_5 g08201(.A(pi252), .B(pi161), .Y(new_n8578));
  nand_5 g08202(.A(pi242), .B(pi090), .Y(new_n8579));
  nand_5 g08203(.A(pi141), .B(pi140), .Y(new_n8580));
  xor_4  g08204(.A(new_n8580), .B(new_n8579), .Y(new_n8581));
  xor_4  g08205(.A(new_n8581), .B(new_n8578), .Y(new_n8582));
  nand_5 g08206(.A(pi241), .B(pi121), .Y(new_n8583));
  nand_5 g08207(.A(new_n1094), .B(new_n1093), .Y(new_n8584));
  nand_5 g08208(.A(new_n1095), .B(new_n1092), .Y(new_n8585));
  nand_5 g08209(.A(new_n8585), .B(new_n8584), .Y(new_n8586));
  xor_4  g08210(.A(new_n8586), .B(new_n8583), .Y(new_n8587));
  xor_4  g08211(.A(new_n8587), .B(new_n8582), .Y(new_n8588));
  nand_5 g08212(.A(pi236), .B(pi231), .Y(new_n8589));
  or_6   g08213(.A(new_n1090), .B(new_n1089), .Y(new_n8590));
  nand_5 g08214(.A(new_n1096), .B(new_n1091), .Y(new_n8591));
  nand_5 g08215(.A(new_n8591), .B(new_n8590), .Y(new_n8592));
  xor_4  g08216(.A(new_n8592), .B(new_n8589), .Y(new_n8593));
  xor_4  g08217(.A(new_n8593), .B(new_n8588), .Y(new_n8594));
  xor_4  g08218(.A(new_n8594), .B(new_n8577), .Y(new_n8595));
  nor_5  g08219(.A(new_n1127), .B(new_n1120), .Y(new_n8596));
  nand_5 g08220(.A(pi104), .B(pi024), .Y(new_n8597));
  nand_5 g08221(.A(pi210), .B(pi112), .Y(new_n8598));
  nand_5 g08222(.A(pi111), .B(pi013), .Y(new_n8599));
  xor_4  g08223(.A(new_n8599), .B(new_n8598), .Y(new_n8600));
  xor_4  g08224(.A(new_n8600), .B(new_n8597), .Y(new_n8601));
  nand_5 g08225(.A(pi224), .B(pi212), .Y(new_n8602));
  nand_5 g08226(.A(new_n1108), .B(new_n1107), .Y(new_n8603));
  nand_5 g08227(.A(new_n1109), .B(new_n1106), .Y(new_n8604));
  nand_5 g08228(.A(new_n8604), .B(new_n8603), .Y(new_n8605));
  xor_4  g08229(.A(new_n8605), .B(new_n8602), .Y(new_n8606));
  xnor_4 g08230(.A(new_n8606), .B(new_n8601), .Y(new_n8607));
  nand_5 g08231(.A(pi255), .B(pi213), .Y(new_n8608));
  nand_5 g08232(.A(new_n1118), .B(new_n1117), .Y(new_n8609));
  nand_5 g08233(.A(new_n1119), .B(new_n1110), .Y(new_n8610));
  nand_5 g08234(.A(new_n8610), .B(new_n8609), .Y(new_n8611));
  xor_4  g08235(.A(new_n8611), .B(new_n8608), .Y(new_n8612));
  xor_4  g08236(.A(new_n8612), .B(new_n8607), .Y(new_n8613));
  xnor_4 g08237(.A(new_n8613), .B(new_n8596), .Y(new_n8614));
  not_8  g08238(.A(new_n1128), .Y(new_n8615));
  nor_5  g08239(.A(new_n8615), .B(new_n1105), .Y(new_n8616));
  nor_5  g08240(.A(new_n1150), .B(new_n1129), .Y(new_n8617));
  nor_5  g08241(.A(new_n8617), .B(new_n8616), .Y(new_n8618));
  xor_4  g08242(.A(new_n8618), .B(new_n8614), .Y(new_n8619));
  xor_4  g08243(.A(new_n8619), .B(new_n8595), .Y(new_n8620));
  or_6   g08244(.A(new_n1081), .B(new_n1070), .Y(new_n8621));
  nand_5 g08245(.A(pi249), .B(pi015), .Y(new_n8622));
  nand_5 g08246(.A(pi222), .B(pi035), .Y(new_n8623));
  nand_5 g08247(.A(pi139), .B(pi125), .Y(new_n8624));
  xor_4  g08248(.A(new_n8624), .B(new_n8623), .Y(new_n8625));
  xor_4  g08249(.A(new_n8625), .B(new_n8622), .Y(new_n8626));
  nand_5 g08250(.A(pi208), .B(pi176), .Y(new_n8627));
  nand_5 g08251(.A(new_n1073), .B(new_n1072), .Y(new_n8628));
  nand_5 g08252(.A(new_n1074), .B(new_n1071), .Y(new_n8629));
  nand_5 g08253(.A(new_n8629), .B(new_n8628), .Y(new_n8630));
  xor_4  g08254(.A(new_n8630), .B(new_n8627), .Y(new_n8631));
  xnor_4 g08255(.A(new_n8631), .B(new_n8626), .Y(new_n8632));
  nand_5 g08256(.A(pi168), .B(pi040), .Y(new_n8633));
  nand_5 g08257(.A(new_n1079), .B(new_n1076), .Y(new_n8634));
  nand_5 g08258(.A(new_n1080), .B(new_n1075), .Y(new_n8635));
  nand_5 g08259(.A(new_n8635), .B(new_n8634), .Y(new_n8636));
  xor_4  g08260(.A(new_n8636), .B(new_n8633), .Y(new_n8637));
  xnor_4 g08261(.A(new_n8637), .B(new_n8632), .Y(new_n8638));
  xor_4  g08262(.A(new_n8638), .B(new_n8621), .Y(new_n8639));
  nand_5 g08263(.A(new_n1151), .B(new_n1082), .Y(new_n8640));
  nand_5 g08264(.A(new_n1171), .B(new_n1152), .Y(new_n8641));
  nand_5 g08265(.A(new_n8641), .B(new_n8640), .Y(new_n8642));
  xor_4  g08266(.A(new_n8642), .B(new_n8639), .Y(new_n8643));
  xnor_4 g08267(.A(new_n8643), .B(new_n8620), .Y(new_n8644));
  nor_5  g08268(.A(new_n1194), .B(new_n1187), .Y(new_n8645));
  nand_5 g08269(.A(pi131), .B(pi106), .Y(new_n8646));
  nand_5 g08270(.A(new_n1185), .B(new_n1184), .Y(new_n8647));
  nand_5 g08271(.A(new_n1186), .B(new_n1177), .Y(new_n8648));
  nand_5 g08272(.A(new_n8648), .B(new_n8647), .Y(new_n8649));
  xor_4  g08273(.A(new_n8649), .B(new_n8646), .Y(new_n8650));
  nand_5 g08274(.A(pi133), .B(pi100), .Y(new_n8651));
  nand_5 g08275(.A(pi227), .B(pi077), .Y(new_n8652));
  nand_5 g08276(.A(pi217), .B(pi189), .Y(new_n8653));
  xor_4  g08277(.A(new_n8653), .B(new_n8652), .Y(new_n8654));
  xor_4  g08278(.A(new_n8654), .B(new_n8651), .Y(new_n8655));
  nand_5 g08279(.A(pi081), .B(pi052), .Y(new_n8656));
  nand_5 g08280(.A(new_n1175), .B(new_n1174), .Y(new_n8657));
  nand_5 g08281(.A(new_n1176), .B(new_n1173), .Y(new_n8658));
  nand_5 g08282(.A(new_n8658), .B(new_n8657), .Y(new_n8659));
  xor_4  g08283(.A(new_n8659), .B(new_n8656), .Y(new_n8660));
  xnor_4 g08284(.A(new_n8660), .B(new_n8655), .Y(new_n8661));
  xor_4  g08285(.A(new_n8661), .B(new_n8650), .Y(new_n8662));
  xor_4  g08286(.A(new_n8662), .B(new_n8645), .Y(new_n8663));
  not_8  g08287(.A(new_n8663), .Y(new_n8664));
  xor_4  g08288(.A(new_n8664), .B(new_n8644), .Y(new_n8665));
  nand_5 g08289(.A(new_n1213), .B(new_n1195), .Y(new_n8666));
  not_8  g08290(.A(new_n1172), .Y(new_n8667));
  nand_5 g08291(.A(new_n1214), .B(new_n8667), .Y(new_n8668));
  nand_5 g08292(.A(new_n8668), .B(new_n8666), .Y(new_n8669));
  xnor_4 g08293(.A(new_n8669), .B(new_n8665), .Y(po050));
  nand_5 g08294(.A(pi216), .B(pi125), .Y(new_n8671));
  nand_5 g08295(.A(pi222), .B(pi076), .Y(new_n8672));
  nand_5 g08296(.A(pi249), .B(pi079), .Y(new_n8673));
  nand_5 g08297(.A(new_n8673), .B(new_n8672), .Y(new_n8674));
  nand_5 g08298(.A(pi249), .B(pi076), .Y(new_n8675));
  nand_5 g08299(.A(pi222), .B(pi079), .Y(new_n8676));
  or_6   g08300(.A(new_n8676), .B(new_n8675), .Y(new_n8677));
  nand_5 g08301(.A(new_n8677), .B(new_n8674), .Y(new_n8678));
  xor_4  g08302(.A(new_n8678), .B(new_n8671), .Y(new_n8679));
  nand_5 g08303(.A(pi125), .B(pi041), .Y(new_n8680));
  nand_5 g08304(.A(new_n8680), .B(new_n8675), .Y(new_n8681));
  nand_5 g08305(.A(pi222), .B(pi216), .Y(new_n8682));
  xor_4  g08306(.A(new_n8680), .B(new_n8675), .Y(new_n8683));
  nand_5 g08307(.A(new_n8683), .B(new_n8682), .Y(new_n8684));
  nand_5 g08308(.A(new_n8684), .B(new_n8681), .Y(new_n8685));
  xor_4  g08309(.A(new_n8685), .B(new_n8679), .Y(new_n8686));
  nand_5 g08310(.A(pi182), .B(pi176), .Y(new_n8687));
  nand_5 g08311(.A(pi222), .B(pi041), .Y(new_n8688));
  nand_5 g08312(.A(pi249), .B(pi216), .Y(new_n8689));
  nand_5 g08313(.A(new_n8689), .B(new_n8688), .Y(new_n8690));
  nand_5 g08314(.A(pi182), .B(pi125), .Y(new_n8691));
  xor_4  g08315(.A(new_n8689), .B(new_n8688), .Y(new_n8692));
  nand_5 g08316(.A(new_n8692), .B(new_n8691), .Y(new_n8693));
  nand_5 g08317(.A(new_n8693), .B(new_n8690), .Y(new_n8694));
  nand_5 g08318(.A(new_n8694), .B(new_n8687), .Y(new_n8695));
  xor_4  g08319(.A(new_n8683), .B(new_n8682), .Y(new_n8696));
  xor_4  g08320(.A(new_n8694), .B(new_n8687), .Y(new_n8697));
  nand_5 g08321(.A(new_n8697), .B(new_n8696), .Y(new_n8698));
  nand_5 g08322(.A(new_n8698), .B(new_n8695), .Y(new_n8699));
  nand_5 g08323(.A(pi176), .B(pi041), .Y(new_n8700));
  nand_5 g08324(.A(pi182), .B(pi040), .Y(new_n8701));
  nand_5 g08325(.A(new_n8701), .B(new_n8700), .Y(new_n8702));
  nand_5 g08326(.A(pi041), .B(pi040), .Y(new_n8703));
  or_6   g08327(.A(new_n8703), .B(new_n8687), .Y(new_n8704));
  nand_5 g08328(.A(new_n8704), .B(new_n8702), .Y(new_n8705));
  xor_4  g08329(.A(new_n8705), .B(new_n8699), .Y(new_n8706));
  xor_4  g08330(.A(new_n8706), .B(new_n8686), .Y(new_n8707));
  not_8  g08331(.A(new_n8707), .Y(new_n8708));
  xor_4  g08332(.A(new_n8697), .B(new_n8696), .Y(new_n8709));
  nand_5 g08333(.A(pi138), .B(pi040), .Y(new_n8710));
  or_6   g08334(.A(new_n8710), .B(new_n8709), .Y(new_n8711));
  xor_4  g08335(.A(new_n8710), .B(new_n8709), .Y(new_n8712));
  nand_5 g08336(.A(pi249), .B(pi041), .Y(new_n8713));
  nand_5 g08337(.A(pi138), .B(pi125), .Y(new_n8714));
  nand_5 g08338(.A(new_n8714), .B(new_n8713), .Y(new_n8715));
  nand_5 g08339(.A(pi222), .B(pi182), .Y(new_n8716));
  or_6   g08340(.A(new_n8714), .B(new_n8713), .Y(new_n8717));
  nand_5 g08341(.A(new_n8717), .B(new_n8716), .Y(new_n8718));
  nand_5 g08342(.A(new_n8718), .B(new_n8715), .Y(new_n8719));
  nand_5 g08343(.A(pi176), .B(pi138), .Y(new_n8720));
  or_6   g08344(.A(new_n8720), .B(new_n8719), .Y(new_n8721));
  xnor_4 g08345(.A(new_n8692), .B(new_n8691), .Y(new_n8722));
  xor_4  g08346(.A(new_n8720), .B(new_n8719), .Y(new_n8723));
  nand_5 g08347(.A(new_n8723), .B(new_n8722), .Y(new_n8724));
  nand_5 g08348(.A(new_n8724), .B(new_n8721), .Y(new_n8725));
  nand_5 g08349(.A(new_n8725), .B(new_n8712), .Y(new_n8726));
  nand_5 g08350(.A(new_n8726), .B(new_n8711), .Y(new_n8727));
  nand_5 g08351(.A(new_n8727), .B(new_n8708), .Y(new_n8728));
  nand_5 g08352(.A(pi125), .B(pi076), .Y(new_n8729));
  nand_5 g08353(.A(pi251), .B(pi249), .Y(new_n8730));
  xor_4  g08354(.A(new_n8730), .B(new_n8729), .Y(new_n8731));
  xor_4  g08355(.A(new_n8731), .B(new_n8676), .Y(new_n8732));
  not_8  g08356(.A(new_n8732), .Y(new_n8733));
  nand_5 g08357(.A(pi216), .B(pi176), .Y(new_n8734));
  xor_4  g08358(.A(new_n8734), .B(new_n8677), .Y(new_n8735));
  xor_4  g08359(.A(new_n8735), .B(new_n8733), .Y(new_n8736));
  nand_5 g08360(.A(pi182), .B(pi174), .Y(new_n8737));
  nand_5 g08361(.A(pi157), .B(pi138), .Y(new_n8738));
  xor_4  g08362(.A(new_n8738), .B(new_n8737), .Y(new_n8739));
  xor_4  g08363(.A(new_n8739), .B(new_n8703), .Y(new_n8740));
  nand_5 g08364(.A(new_n8678), .B(new_n8671), .Y(new_n8741));
  nand_5 g08365(.A(new_n8685), .B(new_n8679), .Y(new_n8742));
  nand_5 g08366(.A(new_n8742), .B(new_n8741), .Y(new_n8743));
  xor_4  g08367(.A(new_n8743), .B(new_n8740), .Y(new_n8744));
  xor_4  g08368(.A(new_n8744), .B(new_n8736), .Y(new_n8745));
  nand_5 g08369(.A(new_n8705), .B(new_n8699), .Y(new_n8746));
  nand_5 g08370(.A(new_n8706), .B(new_n8686), .Y(new_n8747));
  nand_5 g08371(.A(new_n8747), .B(new_n8746), .Y(new_n8748));
  xor_4  g08372(.A(new_n8748), .B(new_n8704), .Y(new_n8749));
  xnor_4 g08373(.A(new_n8749), .B(new_n8745), .Y(new_n8750));
  xnor_4 g08374(.A(new_n8750), .B(new_n8728), .Y(new_n8751));
  nand_5 g08375(.A(pi174), .B(pi138), .Y(new_n8752));
  xor_4  g08376(.A(new_n8725), .B(new_n8712), .Y(new_n8753));
  xnor_4 g08377(.A(new_n8723), .B(new_n8722), .Y(new_n8754));
  not_8  g08378(.A(new_n8716), .Y(new_n8755));
  not_8  g08379(.A(new_n8715), .Y(new_n8756));
  nand_5 g08380(.A(pi249), .B(pi138), .Y(new_n8757));
  nand_5 g08381(.A(new_n8757), .B(new_n8755), .Y(new_n8758));
  nand_5 g08382(.A(new_n8758), .B(new_n8756), .Y(new_n8759));
  nand_5 g08383(.A(new_n8759), .B(new_n8717), .Y(new_n8760));
  nand_5 g08384(.A(new_n8760), .B(new_n8755), .Y(new_n8761));
  nor_5  g08385(.A(new_n8761), .B(new_n8754), .Y(new_n8762));
  nand_5 g08386(.A(new_n8762), .B(new_n8753), .Y(new_n8763));
  nand_5 g08387(.A(new_n8763), .B(new_n8752), .Y(new_n8764));
  xor_4  g08388(.A(new_n8727), .B(new_n8707), .Y(new_n8765));
  xor_4  g08389(.A(new_n8763), .B(new_n8752), .Y(new_n8766));
  nand_5 g08390(.A(new_n8766), .B(new_n8765), .Y(new_n8767));
  nand_5 g08391(.A(new_n8767), .B(new_n8764), .Y(new_n8768));
  xor_4  g08392(.A(new_n8768), .B(new_n8751), .Y(new_n8769));
  nand_5 g08393(.A(pi123), .B(pi024), .Y(new_n8770));
  nand_5 g08394(.A(pi210), .B(pi023), .Y(new_n8771));
  nand_5 g08395(.A(pi111), .B(pi099), .Y(new_n8772));
  nand_5 g08396(.A(new_n8772), .B(new_n8771), .Y(new_n8773));
  nand_5 g08397(.A(pi210), .B(pi099), .Y(new_n8774));
  nand_5 g08398(.A(pi111), .B(pi023), .Y(new_n8775));
  or_6   g08399(.A(new_n8775), .B(new_n8774), .Y(new_n8776));
  nand_5 g08400(.A(new_n8776), .B(new_n8773), .Y(new_n8777));
  xor_4  g08401(.A(new_n8777), .B(new_n8770), .Y(new_n8778));
  nand_5 g08402(.A(pi169), .B(pi024), .Y(new_n8779));
  nand_5 g08403(.A(pi123), .B(pi111), .Y(new_n8780));
  nand_5 g08404(.A(new_n8780), .B(new_n8779), .Y(new_n8781));
  xor_4  g08405(.A(new_n8780), .B(new_n8779), .Y(new_n8782));
  nand_5 g08406(.A(new_n8782), .B(new_n8774), .Y(new_n8783));
  nand_5 g08407(.A(new_n8783), .B(new_n8781), .Y(new_n8784));
  xor_4  g08408(.A(new_n8784), .B(new_n8778), .Y(new_n8785));
  nand_5 g08409(.A(pi224), .B(pi169), .Y(new_n8786));
  nand_5 g08410(.A(pi255), .B(pi071), .Y(new_n8787));
  and_6  g08411(.A(new_n8787), .B(new_n8786), .Y(new_n8788));
  nand_5 g08412(.A(pi224), .B(pi071), .Y(new_n8789));
  nand_5 g08413(.A(pi255), .B(pi169), .Y(new_n8790));
  nor_5  g08414(.A(new_n8790), .B(new_n8789), .Y(new_n8791));
  or_6   g08415(.A(new_n8791), .B(new_n8788), .Y(new_n8792));
  xnor_4 g08416(.A(new_n8792), .B(new_n8785), .Y(new_n8793));
  nand_5 g08417(.A(pi169), .B(pi111), .Y(new_n8794));
  nand_5 g08418(.A(pi071), .B(pi024), .Y(new_n8795));
  nand_5 g08419(.A(new_n8795), .B(new_n8794), .Y(new_n8796));
  nand_5 g08420(.A(pi210), .B(pi123), .Y(new_n8797));
  xor_4  g08421(.A(new_n8795), .B(new_n8794), .Y(new_n8798));
  nand_5 g08422(.A(new_n8798), .B(new_n8797), .Y(new_n8799));
  nand_5 g08423(.A(new_n8799), .B(new_n8796), .Y(new_n8800));
  nand_5 g08424(.A(new_n8800), .B(new_n8789), .Y(new_n8801));
  xor_4  g08425(.A(new_n8782), .B(new_n8774), .Y(new_n8802));
  xor_4  g08426(.A(new_n8800), .B(new_n8789), .Y(new_n8803));
  nand_5 g08427(.A(new_n8803), .B(new_n8802), .Y(new_n8804));
  nand_5 g08428(.A(new_n8804), .B(new_n8801), .Y(new_n8805));
  xor_4  g08429(.A(new_n8805), .B(new_n8793), .Y(new_n8806));
  nand_5 g08430(.A(pi255), .B(pi142), .Y(new_n8807));
  not_8  g08431(.A(new_n8807), .Y(new_n8808));
  nand_5 g08432(.A(pi210), .B(pi169), .Y(new_n8809));
  nand_5 g08433(.A(pi142), .B(pi024), .Y(new_n8810));
  nand_5 g08434(.A(new_n8810), .B(new_n8809), .Y(new_n8811));
  nand_5 g08435(.A(pi111), .B(pi071), .Y(new_n8812));
  or_6   g08436(.A(new_n8810), .B(new_n8809), .Y(new_n8813));
  nand_5 g08437(.A(new_n8813), .B(new_n8812), .Y(new_n8814));
  nand_5 g08438(.A(new_n8814), .B(new_n8811), .Y(new_n8815));
  nand_5 g08439(.A(pi224), .B(pi142), .Y(new_n8816));
  or_6   g08440(.A(new_n8816), .B(new_n8815), .Y(new_n8817));
  xor_4  g08441(.A(new_n8816), .B(new_n8815), .Y(new_n8818));
  xnor_4 g08442(.A(new_n8798), .B(new_n8797), .Y(new_n8819));
  nand_5 g08443(.A(new_n8819), .B(new_n8818), .Y(new_n8820));
  nand_5 g08444(.A(new_n8820), .B(new_n8817), .Y(new_n8821));
  nand_5 g08445(.A(new_n8821), .B(new_n8808), .Y(new_n8822));
  xor_4  g08446(.A(new_n8821), .B(new_n8807), .Y(new_n8823));
  xor_4  g08447(.A(new_n8803), .B(new_n8802), .Y(new_n8824));
  or_6   g08448(.A(new_n8824), .B(new_n8823), .Y(new_n8825));
  nand_5 g08449(.A(new_n8825), .B(new_n8822), .Y(new_n8826));
  nand_5 g08450(.A(new_n8826), .B(new_n8806), .Y(new_n8827));
  nand_5 g08451(.A(pi099), .B(pi024), .Y(new_n8828));
  nand_5 g08452(.A(pi210), .B(pi155), .Y(new_n8829));
  xor_4  g08453(.A(new_n8829), .B(new_n8775), .Y(new_n8830));
  xor_4  g08454(.A(new_n8830), .B(new_n8828), .Y(new_n8831));
  nand_5 g08455(.A(pi224), .B(pi123), .Y(new_n8832));
  xor_4  g08456(.A(new_n8832), .B(new_n8776), .Y(new_n8833));
  xor_4  g08457(.A(new_n8833), .B(new_n8831), .Y(new_n8834));
  nand_5 g08458(.A(pi127), .B(pi071), .Y(new_n8835));
  nand_5 g08459(.A(pi232), .B(pi142), .Y(new_n8836));
  xor_4  g08460(.A(new_n8836), .B(new_n8835), .Y(new_n8837));
  xor_4  g08461(.A(new_n8837), .B(new_n8790), .Y(new_n8838));
  nand_5 g08462(.A(new_n8777), .B(new_n8770), .Y(new_n8839));
  nand_5 g08463(.A(new_n8784), .B(new_n8778), .Y(new_n8840));
  nand_5 g08464(.A(new_n8840), .B(new_n8839), .Y(new_n8841));
  xor_4  g08465(.A(new_n8841), .B(new_n8838), .Y(new_n8842));
  xnor_4 g08466(.A(new_n8842), .B(new_n8834), .Y(new_n8843));
  nor_5  g08467(.A(new_n8805), .B(new_n8793), .Y(new_n8844));
  nand_5 g08468(.A(new_n8844), .B(new_n8791), .Y(new_n8845));
  nor_5  g08469(.A(new_n8792), .B(new_n8785), .Y(new_n8846));
  or_6   g08470(.A(new_n8846), .B(new_n8791), .Y(new_n8847));
  or_6   g08471(.A(new_n8847), .B(new_n8844), .Y(new_n8848));
  nand_5 g08472(.A(new_n8848), .B(new_n8845), .Y(new_n8849));
  xor_4  g08473(.A(new_n8849), .B(new_n8843), .Y(new_n8850));
  xnor_4 g08474(.A(new_n8850), .B(new_n8827), .Y(new_n8851));
  nand_5 g08475(.A(pi142), .B(pi127), .Y(new_n8852));
  xnor_4 g08476(.A(new_n8819), .B(new_n8818), .Y(new_n8853));
  not_8  g08477(.A(new_n8812), .Y(new_n8854));
  not_8  g08478(.A(new_n8811), .Y(new_n8855));
  nand_5 g08479(.A(pi210), .B(pi142), .Y(new_n8856));
  nand_5 g08480(.A(new_n8856), .B(new_n8854), .Y(new_n8857));
  nand_5 g08481(.A(new_n8857), .B(new_n8855), .Y(new_n8858));
  nand_5 g08482(.A(new_n8858), .B(new_n8813), .Y(new_n8859));
  nand_5 g08483(.A(new_n8859), .B(new_n8854), .Y(new_n8860));
  nor_5  g08484(.A(new_n8860), .B(new_n8853), .Y(new_n8861));
  xor_4  g08485(.A(new_n8824), .B(new_n8823), .Y(new_n8862));
  nand_5 g08486(.A(new_n8862), .B(new_n8861), .Y(new_n8863));
  nand_5 g08487(.A(new_n8863), .B(new_n8852), .Y(new_n8864));
  xnor_4 g08488(.A(new_n8826), .B(new_n8806), .Y(new_n8865));
  xor_4  g08489(.A(new_n8863), .B(new_n8852), .Y(new_n8866));
  nand_5 g08490(.A(new_n8866), .B(new_n8865), .Y(new_n8867));
  nand_5 g08491(.A(new_n8867), .B(new_n8864), .Y(new_n8868));
  xor_4  g08492(.A(new_n8868), .B(new_n8851), .Y(new_n8869));
  nand_5 g08493(.A(pi140), .B(pi135), .Y(new_n8870));
  nand_5 g08494(.A(pi252), .B(pi122), .Y(new_n8871));
  nand_5 g08495(.A(pi242), .B(pi059), .Y(new_n8872));
  xor_4  g08496(.A(new_n8872), .B(new_n8871), .Y(new_n8873));
  xor_4  g08497(.A(new_n8873), .B(new_n8870), .Y(new_n8874));
  not_8  g08498(.A(new_n8874), .Y(new_n8875));
  nand_5 g08499(.A(pi121), .B(pi001), .Y(new_n8876));
  nand_5 g08500(.A(pi242), .B(pi122), .Y(new_n8877));
  or_6   g08501(.A(new_n8877), .B(new_n8870), .Y(new_n8878));
  xor_4  g08502(.A(new_n8878), .B(new_n8876), .Y(new_n8879));
  xor_4  g08503(.A(new_n8879), .B(new_n8875), .Y(new_n8880));
  nand_5 g08504(.A(pi231), .B(pi102), .Y(new_n8881));
  nand_5 g08505(.A(pi087), .B(pi021), .Y(new_n8882));
  nand_5 g08506(.A(pi219), .B(pi005), .Y(new_n8883));
  xor_4  g08507(.A(new_n8883), .B(new_n8882), .Y(new_n8884));
  xor_4  g08508(.A(new_n8884), .B(new_n8881), .Y(new_n8885));
  nand_5 g08509(.A(pi252), .B(pi001), .Y(new_n8886));
  nand_5 g08510(.A(pi140), .B(pi122), .Y(new_n8887));
  nand_5 g08511(.A(pi242), .B(pi135), .Y(new_n8888));
  nand_5 g08512(.A(new_n8888), .B(new_n8887), .Y(new_n8889));
  nand_5 g08513(.A(new_n8889), .B(new_n8878), .Y(new_n8890));
  nand_5 g08514(.A(new_n8890), .B(new_n8886), .Y(new_n8891));
  xor_4  g08515(.A(new_n8890), .B(new_n8886), .Y(new_n8892));
  nand_5 g08516(.A(pi140), .B(pi001), .Y(new_n8893));
  nand_5 g08517(.A(new_n8893), .B(new_n8877), .Y(new_n8894));
  nand_5 g08518(.A(pi252), .B(pi102), .Y(new_n8895));
  xor_4  g08519(.A(new_n8893), .B(new_n8877), .Y(new_n8896));
  nand_5 g08520(.A(new_n8896), .B(new_n8895), .Y(new_n8897));
  nand_5 g08521(.A(new_n8897), .B(new_n8894), .Y(new_n8898));
  nand_5 g08522(.A(new_n8898), .B(new_n8892), .Y(new_n8899));
  nand_5 g08523(.A(new_n8899), .B(new_n8891), .Y(new_n8900));
  xor_4  g08524(.A(new_n8900), .B(new_n8885), .Y(new_n8901));
  xor_4  g08525(.A(new_n8901), .B(new_n8880), .Y(new_n8902));
  not_8  g08526(.A(new_n8902), .Y(new_n8903));
  nand_5 g08527(.A(pi219), .B(pi121), .Y(new_n8904));
  or_6   g08528(.A(new_n8904), .B(new_n8881), .Y(new_n8905));
  nand_5 g08529(.A(pi242), .B(pi001), .Y(new_n8906));
  nand_5 g08530(.A(pi252), .B(pi219), .Y(new_n8907));
  nand_5 g08531(.A(new_n8907), .B(new_n8906), .Y(new_n8908));
  nand_5 g08532(.A(pi140), .B(pi102), .Y(new_n8909));
  xor_4  g08533(.A(new_n8907), .B(new_n8906), .Y(new_n8910));
  nand_5 g08534(.A(new_n8910), .B(new_n8909), .Y(new_n8911));
  nand_5 g08535(.A(new_n8911), .B(new_n8908), .Y(new_n8912));
  nand_5 g08536(.A(new_n8912), .B(new_n8904), .Y(new_n8913));
  xor_4  g08537(.A(new_n8896), .B(new_n8895), .Y(new_n8914));
  xor_4  g08538(.A(new_n8912), .B(new_n8904), .Y(new_n8915));
  nand_5 g08539(.A(new_n8915), .B(new_n8914), .Y(new_n8916));
  nand_5 g08540(.A(new_n8916), .B(new_n8913), .Y(new_n8917));
  nand_5 g08541(.A(pi121), .B(pi102), .Y(new_n8918));
  nand_5 g08542(.A(pi231), .B(pi219), .Y(new_n8919));
  nand_5 g08543(.A(new_n8919), .B(new_n8918), .Y(new_n8920));
  nand_5 g08544(.A(new_n8920), .B(new_n8905), .Y(new_n8921));
  nand_5 g08545(.A(new_n8921), .B(new_n8917), .Y(new_n8922));
  xor_4  g08546(.A(new_n8898), .B(new_n8892), .Y(new_n8923));
  xor_4  g08547(.A(new_n8921), .B(new_n8917), .Y(new_n8924));
  nand_5 g08548(.A(new_n8924), .B(new_n8923), .Y(new_n8925));
  nand_5 g08549(.A(new_n8925), .B(new_n8922), .Y(new_n8926));
  xor_4  g08550(.A(new_n8926), .B(new_n8905), .Y(new_n8927));
  xor_4  g08551(.A(new_n8927), .B(new_n8903), .Y(new_n8928));
  xor_4  g08552(.A(new_n8924), .B(new_n8923), .Y(new_n8929));
  not_8  g08553(.A(new_n8929), .Y(new_n8930));
  nand_5 g08554(.A(pi231), .B(pi087), .Y(new_n8931));
  not_8  g08555(.A(new_n8931), .Y(new_n8932));
  nand_5 g08556(.A(pi242), .B(pi102), .Y(new_n8933));
  nand_5 g08557(.A(pi252), .B(pi087), .Y(new_n8934));
  nand_5 g08558(.A(new_n8934), .B(new_n8933), .Y(new_n8935));
  nand_5 g08559(.A(pi219), .B(pi140), .Y(new_n8936));
  or_6   g08560(.A(new_n8934), .B(new_n8933), .Y(new_n8937));
  nand_5 g08561(.A(new_n8937), .B(new_n8936), .Y(new_n8938));
  nand_5 g08562(.A(new_n8938), .B(new_n8935), .Y(new_n8939));
  nand_5 g08563(.A(pi121), .B(pi087), .Y(new_n8940));
  or_6   g08564(.A(new_n8940), .B(new_n8939), .Y(new_n8941));
  xor_4  g08565(.A(new_n8940), .B(new_n8939), .Y(new_n8942));
  xnor_4 g08566(.A(new_n8910), .B(new_n8909), .Y(new_n8943));
  nand_5 g08567(.A(new_n8943), .B(new_n8942), .Y(new_n8944));
  nand_5 g08568(.A(new_n8944), .B(new_n8941), .Y(new_n8945));
  nand_5 g08569(.A(new_n8945), .B(new_n8932), .Y(new_n8946));
  xor_4  g08570(.A(new_n8915), .B(new_n8914), .Y(new_n8947));
  xor_4  g08571(.A(new_n8945), .B(new_n8931), .Y(new_n8948));
  or_6   g08572(.A(new_n8948), .B(new_n8947), .Y(new_n8949));
  nand_5 g08573(.A(new_n8949), .B(new_n8946), .Y(new_n8950));
  nand_5 g08574(.A(new_n8950), .B(new_n8930), .Y(new_n8951));
  xnor_4 g08575(.A(new_n8943), .B(new_n8942), .Y(new_n8952));
  not_8  g08576(.A(new_n8936), .Y(new_n8953));
  not_8  g08577(.A(new_n8935), .Y(new_n8954));
  nand_5 g08578(.A(pi242), .B(pi087), .Y(new_n8955));
  nand_5 g08579(.A(new_n8955), .B(new_n8953), .Y(new_n8956));
  nand_5 g08580(.A(new_n8956), .B(new_n8954), .Y(new_n8957));
  nand_5 g08581(.A(new_n8957), .B(new_n8937), .Y(new_n8958));
  nand_5 g08582(.A(new_n8958), .B(new_n8953), .Y(new_n8959));
  nor_5  g08583(.A(new_n8959), .B(new_n8952), .Y(new_n8960));
  xor_4  g08584(.A(new_n8948), .B(new_n8947), .Y(new_n8961));
  nand_5 g08585(.A(new_n8961), .B(new_n8960), .Y(new_n8962));
  nand_5 g08586(.A(pi087), .B(pi005), .Y(new_n8963));
  xor_4  g08587(.A(new_n8950), .B(new_n8929), .Y(new_n8964));
  xnor_4 g08588(.A(new_n8964), .B(new_n8963), .Y(new_n8965));
  nor_5  g08589(.A(new_n8965), .B(new_n8962), .Y(new_n8966));
  not_8  g08590(.A(new_n8966), .Y(new_n8967));
  nor_5  g08591(.A(new_n8967), .B(new_n8951), .Y(new_n8968));
  or_6   g08592(.A(new_n8964), .B(new_n8963), .Y(new_n8969));
  nand_5 g08593(.A(new_n8969), .B(new_n8951), .Y(new_n8970));
  nor_5  g08594(.A(new_n8970), .B(new_n8966), .Y(new_n8971));
  nor_5  g08595(.A(new_n8971), .B(new_n8968), .Y(new_n8972));
  xor_4  g08596(.A(new_n8972), .B(new_n8928), .Y(new_n8973));
  not_8  g08597(.A(new_n8973), .Y(new_n8974));
  xor_4  g08598(.A(new_n8974), .B(new_n8869), .Y(new_n8975));
  xnor_4 g08599(.A(new_n8866), .B(new_n8865), .Y(new_n8976));
  xor_4  g08600(.A(new_n8965), .B(new_n8962), .Y(new_n8977));
  nand_5 g08601(.A(new_n8977), .B(new_n8976), .Y(new_n8978));
  xor_4  g08602(.A(new_n8977), .B(new_n8976), .Y(new_n8979));
  xor_4  g08603(.A(new_n8961), .B(new_n8960), .Y(new_n8980));
  xor_4  g08604(.A(new_n8862), .B(new_n8861), .Y(new_n8981));
  nand_5 g08605(.A(new_n8981), .B(new_n8980), .Y(new_n8982));
  not_8  g08606(.A(new_n8982), .Y(new_n8983));
  xnor_4 g08607(.A(new_n8981), .B(new_n8980), .Y(new_n8984));
  xnor_4 g08608(.A(new_n8959), .B(new_n8952), .Y(new_n8985));
  nor_5  g08609(.A(new_n8857), .B(new_n8855), .Y(new_n8986));
  or_6   g08610(.A(new_n8986), .B(new_n8859), .Y(new_n8987));
  nor_5  g08611(.A(new_n8956), .B(new_n8954), .Y(new_n8988));
  nor_5  g08612(.A(new_n8988), .B(new_n8958), .Y(new_n8989));
  not_8  g08613(.A(new_n8989), .Y(new_n8990));
  nand_5 g08614(.A(new_n8990), .B(new_n8987), .Y(new_n8991));
  xor_4  g08615(.A(new_n8989), .B(new_n8987), .Y(new_n8992));
  nand_5 g08616(.A(pi142), .B(pi111), .Y(new_n8993));
  nand_5 g08617(.A(pi210), .B(pi071), .Y(new_n8994));
  xor_4  g08618(.A(new_n8994), .B(new_n8993), .Y(new_n8995));
  nor_5  g08619(.A(new_n8955), .B(new_n8856), .Y(new_n8996));
  nand_5 g08620(.A(new_n8996), .B(new_n8995), .Y(new_n8997));
  nand_5 g08621(.A(pi242), .B(pi219), .Y(new_n8998));
  nand_5 g08622(.A(pi140), .B(pi087), .Y(new_n8999));
  xor_4  g08623(.A(new_n8999), .B(new_n8998), .Y(new_n9000));
  xor_4  g08624(.A(new_n8996), .B(new_n8995), .Y(new_n9001));
  nand_5 g08625(.A(new_n9001), .B(new_n9000), .Y(new_n9002));
  nand_5 g08626(.A(new_n9002), .B(new_n8997), .Y(new_n9003));
  or_6   g08627(.A(new_n9003), .B(new_n8992), .Y(new_n9004));
  nand_5 g08628(.A(new_n9004), .B(new_n8991), .Y(new_n9005));
  nand_5 g08629(.A(new_n9005), .B(new_n8985), .Y(new_n9006));
  xor_4  g08630(.A(new_n8860), .B(new_n8853), .Y(new_n9007));
  not_8  g08631(.A(new_n9007), .Y(new_n9008));
  xor_4  g08632(.A(new_n9005), .B(new_n8985), .Y(new_n9009));
  nand_5 g08633(.A(new_n9009), .B(new_n9008), .Y(new_n9010));
  nand_5 g08634(.A(new_n9010), .B(new_n9006), .Y(new_n9011));
  nor_5  g08635(.A(new_n9011), .B(new_n8984), .Y(new_n9012));
  nor_5  g08636(.A(new_n9012), .B(new_n8983), .Y(new_n9013));
  not_8  g08637(.A(new_n9013), .Y(new_n9014));
  nand_5 g08638(.A(new_n9014), .B(new_n8979), .Y(new_n9015));
  nand_5 g08639(.A(new_n9015), .B(new_n8978), .Y(new_n9016));
  xor_4  g08640(.A(new_n9016), .B(new_n8975), .Y(new_n9017));
  xor_4  g08641(.A(new_n9017), .B(new_n8769), .Y(new_n9018));
  xor_4  g08642(.A(new_n9013), .B(new_n8979), .Y(new_n9019));
  xor_4  g08643(.A(new_n8766), .B(new_n8765), .Y(new_n9020));
  nor_5  g08644(.A(new_n9020), .B(new_n9019), .Y(new_n9021));
  xnor_4 g08645(.A(new_n9020), .B(new_n9019), .Y(new_n9022));
  xor_4  g08646(.A(new_n8762), .B(new_n8753), .Y(new_n9023));
  xor_4  g08647(.A(new_n8761), .B(new_n8754), .Y(new_n9024));
  xor_4  g08648(.A(new_n9009), .B(new_n9008), .Y(new_n9025));
  not_8  g08649(.A(new_n9025), .Y(new_n9026));
  nor_5  g08650(.A(new_n9026), .B(new_n9024), .Y(new_n9027));
  xor_4  g08651(.A(new_n9025), .B(new_n9024), .Y(new_n9028));
  xor_4  g08652(.A(new_n9003), .B(new_n8992), .Y(new_n9029));
  xor_4  g08653(.A(new_n8955), .B(new_n8856), .Y(new_n9030));
  not_8  g08654(.A(new_n9030), .Y(new_n9031));
  nor_5  g08655(.A(new_n9031), .B(new_n8757), .Y(new_n9032));
  nand_5 g08656(.A(pi222), .B(pi138), .Y(new_n9033));
  nand_5 g08657(.A(pi249), .B(pi182), .Y(new_n9034));
  xor_4  g08658(.A(new_n9034), .B(new_n9033), .Y(new_n9035));
  or_6   g08659(.A(new_n9035), .B(new_n9032), .Y(new_n9036));
  xnor_4 g08660(.A(new_n9001), .B(new_n9000), .Y(new_n9037));
  xor_4  g08661(.A(new_n9035), .B(new_n9032), .Y(new_n9038));
  nand_5 g08662(.A(new_n9038), .B(new_n9037), .Y(new_n9039));
  nand_5 g08663(.A(new_n9039), .B(new_n9036), .Y(new_n9040));
  or_6   g08664(.A(new_n9040), .B(new_n9029), .Y(new_n9041));
  xor_4  g08665(.A(new_n9040), .B(new_n9029), .Y(new_n9042));
  nor_5  g08666(.A(new_n8758), .B(new_n8756), .Y(new_n9043));
  nor_5  g08667(.A(new_n9043), .B(new_n8760), .Y(new_n9044));
  nand_5 g08668(.A(new_n9044), .B(new_n9042), .Y(new_n9045));
  nand_5 g08669(.A(new_n9045), .B(new_n9041), .Y(new_n9046));
  nor_5  g08670(.A(new_n9046), .B(new_n9028), .Y(new_n9047));
  nor_5  g08671(.A(new_n9047), .B(new_n9027), .Y(new_n9048));
  or_6   g08672(.A(new_n9048), .B(new_n9023), .Y(new_n9049));
  xor_4  g08673(.A(new_n9011), .B(new_n8984), .Y(new_n9050));
  not_8  g08674(.A(new_n9050), .Y(new_n9051));
  xor_4  g08675(.A(new_n9048), .B(new_n9023), .Y(new_n9052));
  nand_5 g08676(.A(new_n9052), .B(new_n9051), .Y(new_n9053));
  nand_5 g08677(.A(new_n9053), .B(new_n9049), .Y(new_n9054));
  nor_5  g08678(.A(new_n9054), .B(new_n9022), .Y(new_n9055));
  nor_5  g08679(.A(new_n9055), .B(new_n9021), .Y(new_n9056));
  xor_4  g08680(.A(new_n9056), .B(new_n9018), .Y(new_n9057));
  nand_5 g08681(.A(pi233), .B(pi160), .Y(new_n9058));
  nand_5 g08682(.A(pi217), .B(pi060), .Y(new_n9059));
  nand_5 g08683(.A(pi227), .B(pi160), .Y(new_n9060));
  nand_5 g08684(.A(pi100), .B(pi020), .Y(new_n9061));
  xor_4  g08685(.A(new_n9061), .B(new_n9060), .Y(new_n9062));
  xor_4  g08686(.A(new_n9062), .B(new_n9059), .Y(new_n9063));
  nand_5 g08687(.A(pi160), .B(pi100), .Y(new_n9064));
  nand_5 g08688(.A(pi217), .B(pi020), .Y(new_n9065));
  nor_5  g08689(.A(new_n9065), .B(new_n9064), .Y(new_n9066));
  not_8  g08690(.A(new_n9066), .Y(new_n9067));
  nor_5  g08691(.A(new_n9067), .B(new_n9063), .Y(new_n9068));
  not_8  g08692(.A(new_n9068), .Y(new_n9069));
  nand_5 g08693(.A(pi227), .B(pi020), .Y(new_n9070));
  nand_5 g08694(.A(pi223), .B(pi217), .Y(new_n9071));
  nand_5 g08695(.A(pi100), .B(pi060), .Y(new_n9072));
  xor_4  g08696(.A(new_n9072), .B(new_n9071), .Y(new_n9073));
  xnor_4 g08697(.A(new_n9073), .B(new_n9070), .Y(new_n9074));
  nand_5 g08698(.A(pi160), .B(pi081), .Y(new_n9075));
  nand_5 g08699(.A(new_n9061), .B(new_n9060), .Y(new_n9076));
  nand_5 g08700(.A(new_n9062), .B(new_n9059), .Y(new_n9077));
  nand_5 g08701(.A(new_n9077), .B(new_n9076), .Y(new_n9078));
  xor_4  g08702(.A(new_n9078), .B(new_n9075), .Y(new_n9079));
  xnor_4 g08703(.A(new_n9079), .B(new_n9074), .Y(new_n9080));
  nor_5  g08704(.A(new_n9080), .B(new_n9069), .Y(new_n9081));
  nand_5 g08705(.A(pi227), .B(pi060), .Y(new_n9082));
  nand_5 g08706(.A(pi223), .B(pi100), .Y(new_n9083));
  nand_5 g08707(.A(pi217), .B(pi101), .Y(new_n9084));
  xor_4  g08708(.A(new_n9084), .B(new_n9083), .Y(new_n9085));
  xor_4  g08709(.A(new_n9085), .B(new_n9082), .Y(new_n9086));
  nand_5 g08710(.A(pi081), .B(pi020), .Y(new_n9087));
  nand_5 g08711(.A(new_n9072), .B(new_n9071), .Y(new_n9088));
  nand_5 g08712(.A(new_n9073), .B(new_n9070), .Y(new_n9089));
  nand_5 g08713(.A(new_n9089), .B(new_n9088), .Y(new_n9090));
  xor_4  g08714(.A(new_n9090), .B(new_n9087), .Y(new_n9091));
  xor_4  g08715(.A(new_n9091), .B(new_n9086), .Y(new_n9092));
  nand_5 g08716(.A(pi160), .B(pi106), .Y(new_n9093));
  xor_4  g08717(.A(new_n9093), .B(new_n9092), .Y(new_n9094));
  or_6   g08718(.A(new_n9078), .B(new_n9075), .Y(new_n9095));
  nand_5 g08719(.A(new_n9079), .B(new_n9074), .Y(new_n9096));
  nand_5 g08720(.A(new_n9096), .B(new_n9095), .Y(new_n9097));
  xor_4  g08721(.A(new_n9097), .B(new_n9094), .Y(new_n9098));
  nand_5 g08722(.A(new_n9098), .B(new_n9081), .Y(new_n9099));
  nand_5 g08723(.A(new_n9099), .B(new_n9058), .Y(new_n9100));
  nand_5 g08724(.A(pi227), .B(pi223), .Y(new_n9101));
  nand_5 g08725(.A(pi225), .B(pi217), .Y(new_n9102));
  nand_5 g08726(.A(pi101), .B(pi100), .Y(new_n9103));
  nand_5 g08727(.A(new_n9103), .B(new_n9102), .Y(new_n9104));
  nand_5 g08728(.A(pi225), .B(pi100), .Y(new_n9105));
  or_6   g08729(.A(new_n9105), .B(new_n9084), .Y(new_n9106));
  nand_5 g08730(.A(new_n9106), .B(new_n9104), .Y(new_n9107));
  xor_4  g08731(.A(new_n9107), .B(new_n9101), .Y(new_n9108));
  nand_5 g08732(.A(new_n9084), .B(new_n9083), .Y(new_n9109));
  nand_5 g08733(.A(new_n9085), .B(new_n9082), .Y(new_n9110));
  nand_5 g08734(.A(new_n9110), .B(new_n9109), .Y(new_n9111));
  xor_4  g08735(.A(new_n9111), .B(new_n9108), .Y(new_n9112));
  nand_5 g08736(.A(pi081), .B(pi060), .Y(new_n9113));
  nand_5 g08737(.A(pi106), .B(pi020), .Y(new_n9114));
  and_6  g08738(.A(new_n9114), .B(new_n9113), .Y(new_n9115));
  nand_5 g08739(.A(pi106), .B(pi060), .Y(new_n9116));
  nor_5  g08740(.A(new_n9116), .B(new_n9087), .Y(new_n9117));
  or_6   g08741(.A(new_n9117), .B(new_n9115), .Y(new_n9118));
  xnor_4 g08742(.A(new_n9118), .B(new_n9112), .Y(new_n9119));
  nand_5 g08743(.A(new_n9090), .B(new_n9087), .Y(new_n9120));
  nand_5 g08744(.A(new_n9091), .B(new_n9086), .Y(new_n9121));
  nand_5 g08745(.A(new_n9121), .B(new_n9120), .Y(new_n9122));
  xor_4  g08746(.A(new_n9122), .B(new_n9119), .Y(new_n9123));
  or_6   g08747(.A(new_n9093), .B(new_n9092), .Y(new_n9124));
  nand_5 g08748(.A(new_n9097), .B(new_n9094), .Y(new_n9125));
  nand_5 g08749(.A(new_n9125), .B(new_n9124), .Y(new_n9126));
  xnor_4 g08750(.A(new_n9126), .B(new_n9123), .Y(new_n9127));
  xor_4  g08751(.A(new_n9099), .B(new_n9058), .Y(new_n9128));
  nand_5 g08752(.A(new_n9128), .B(new_n9127), .Y(new_n9129));
  nand_5 g08753(.A(new_n9129), .B(new_n9100), .Y(new_n9130));
  nand_5 g08754(.A(new_n9126), .B(new_n9123), .Y(new_n9131));
  nand_5 g08755(.A(pi227), .B(pi101), .Y(new_n9132));
  nand_5 g08756(.A(pi217), .B(pi177), .Y(new_n9133));
  xor_4  g08757(.A(new_n9133), .B(new_n9132), .Y(new_n9134));
  xor_4  g08758(.A(new_n9134), .B(new_n9105), .Y(new_n9135));
  nand_5 g08759(.A(pi223), .B(pi081), .Y(new_n9136));
  xor_4  g08760(.A(new_n9136), .B(new_n9106), .Y(new_n9137));
  xor_4  g08761(.A(new_n9137), .B(new_n9135), .Y(new_n9138));
  nand_5 g08762(.A(pi233), .B(pi020), .Y(new_n9139));
  nand_5 g08763(.A(pi187), .B(pi160), .Y(new_n9140));
  xor_4  g08764(.A(new_n9140), .B(new_n9139), .Y(new_n9141));
  xor_4  g08765(.A(new_n9141), .B(new_n9116), .Y(new_n9142));
  nand_5 g08766(.A(new_n9107), .B(new_n9101), .Y(new_n9143));
  nand_5 g08767(.A(new_n9111), .B(new_n9108), .Y(new_n9144));
  nand_5 g08768(.A(new_n9144), .B(new_n9143), .Y(new_n9145));
  xor_4  g08769(.A(new_n9145), .B(new_n9142), .Y(new_n9146));
  xnor_4 g08770(.A(new_n9146), .B(new_n9138), .Y(new_n9147));
  nor_5  g08771(.A(new_n9118), .B(new_n9112), .Y(new_n9148));
  nor_5  g08772(.A(new_n9122), .B(new_n9119), .Y(new_n9149));
  xor_4  g08773(.A(new_n9149), .B(new_n9117), .Y(new_n9150));
  nor_5  g08774(.A(new_n9150), .B(new_n9148), .Y(new_n9151));
  xor_4  g08775(.A(new_n9151), .B(new_n9147), .Y(new_n9152));
  xor_4  g08776(.A(new_n9152), .B(new_n9131), .Y(new_n9153));
  xor_4  g08777(.A(new_n9153), .B(new_n9130), .Y(new_n9154));
  or_6   g08778(.A(new_n9154), .B(new_n9057), .Y(new_n9155));
  xor_4  g08779(.A(new_n9054), .B(new_n9022), .Y(new_n9156));
  not_8  g08780(.A(new_n9156), .Y(new_n9157));
  xor_4  g08781(.A(new_n9128), .B(new_n9127), .Y(new_n9158));
  or_6   g08782(.A(new_n9158), .B(new_n9157), .Y(new_n9159));
  xor_4  g08783(.A(new_n9158), .B(new_n9157), .Y(new_n9160));
  xnor_4 g08784(.A(new_n9098), .B(new_n9081), .Y(new_n9161));
  xor_4  g08785(.A(new_n9046), .B(new_n9028), .Y(new_n9162));
  xor_4  g08786(.A(new_n9066), .B(new_n9063), .Y(new_n9163));
  nand_5 g08787(.A(pi217), .B(pi160), .Y(new_n9164));
  xor_4  g08788(.A(new_n9030), .B(new_n8757), .Y(new_n9165));
  nor_5  g08789(.A(new_n9165), .B(new_n9164), .Y(new_n9166));
  xor_4  g08790(.A(new_n9065), .B(new_n9064), .Y(new_n9167));
  or_6   g08791(.A(new_n9167), .B(new_n9166), .Y(new_n9168));
  xor_4  g08792(.A(new_n9038), .B(new_n9037), .Y(new_n9169));
  xor_4  g08793(.A(new_n9167), .B(new_n9166), .Y(new_n9170));
  nand_5 g08794(.A(new_n9170), .B(new_n9169), .Y(new_n9171));
  nand_5 g08795(.A(new_n9171), .B(new_n9168), .Y(new_n9172));
  nand_5 g08796(.A(new_n9172), .B(new_n9163), .Y(new_n9173));
  xor_4  g08797(.A(new_n9044), .B(new_n9042), .Y(new_n9174));
  not_8  g08798(.A(new_n9174), .Y(new_n9175));
  xor_4  g08799(.A(new_n9172), .B(new_n9163), .Y(new_n9176));
  nand_5 g08800(.A(new_n9176), .B(new_n9175), .Y(new_n9177));
  nand_5 g08801(.A(new_n9177), .B(new_n9173), .Y(new_n9178));
  nand_5 g08802(.A(new_n9178), .B(new_n9162), .Y(new_n9179));
  xor_4  g08803(.A(new_n9080), .B(new_n9069), .Y(new_n9180));
  not_8  g08804(.A(new_n9180), .Y(new_n9181));
  xor_4  g08805(.A(new_n9178), .B(new_n9162), .Y(new_n9182));
  nand_5 g08806(.A(new_n9182), .B(new_n9181), .Y(new_n9183));
  nand_5 g08807(.A(new_n9183), .B(new_n9179), .Y(new_n9184));
  or_6   g08808(.A(new_n9184), .B(new_n9161), .Y(new_n9185));
  xor_4  g08809(.A(new_n9052), .B(new_n9050), .Y(new_n9186));
  xor_4  g08810(.A(new_n9184), .B(new_n9161), .Y(new_n9187));
  nand_5 g08811(.A(new_n9187), .B(new_n9186), .Y(new_n9188));
  nand_5 g08812(.A(new_n9188), .B(new_n9185), .Y(new_n9189));
  nand_5 g08813(.A(new_n9189), .B(new_n9160), .Y(new_n9190));
  nand_5 g08814(.A(new_n9190), .B(new_n9159), .Y(new_n9191));
  xor_4  g08815(.A(new_n9154), .B(new_n9057), .Y(new_n9192));
  nand_5 g08816(.A(new_n9192), .B(new_n9191), .Y(new_n9193));
  nand_5 g08817(.A(new_n9193), .B(new_n9155), .Y(new_n9194));
  nand_5 g08818(.A(new_n9152), .B(new_n9131), .Y(new_n9195));
  nand_5 g08819(.A(new_n9153), .B(new_n9130), .Y(new_n9196));
  nand_5 g08820(.A(new_n9196), .B(new_n9195), .Y(new_n9197));
  xor_4  g08821(.A(new_n9197), .B(new_n9194), .Y(new_n9198));
  nand_5 g08822(.A(pi155), .B(pi111), .Y(new_n9199));
  nand_5 g08823(.A(pi024), .B(pi023), .Y(new_n9200));
  xor_4  g08824(.A(new_n9200), .B(new_n9199), .Y(new_n9201));
  nand_5 g08825(.A(pi176), .B(pi076), .Y(new_n9202));
  or_6   g08826(.A(new_n8734), .B(new_n8677), .Y(new_n9203));
  nand_5 g08827(.A(new_n8735), .B(new_n8733), .Y(new_n9204));
  nand_5 g08828(.A(new_n9204), .B(new_n9203), .Y(new_n9205));
  xor_4  g08829(.A(new_n9205), .B(new_n9202), .Y(new_n9206));
  nand_5 g08830(.A(pi216), .B(pi040), .Y(new_n9207));
  nand_5 g08831(.A(pi174), .B(pi041), .Y(new_n9208));
  xor_4  g08832(.A(new_n9208), .B(new_n9207), .Y(new_n9209));
  nand_5 g08833(.A(pi125), .B(pi079), .Y(new_n9210));
  xor_4  g08834(.A(new_n9210), .B(new_n9209), .Y(new_n9211));
  nand_5 g08835(.A(pi182), .B(pi157), .Y(new_n9212));
  nand_5 g08836(.A(new_n8730), .B(new_n8729), .Y(new_n9213));
  nand_5 g08837(.A(new_n8731), .B(new_n8676), .Y(new_n9214));
  nand_5 g08838(.A(new_n9214), .B(new_n9213), .Y(new_n9215));
  nand_5 g08839(.A(new_n8743), .B(new_n8740), .Y(new_n9216));
  not_8  g08840(.A(new_n8736), .Y(new_n9217));
  nand_5 g08841(.A(new_n8744), .B(new_n9217), .Y(new_n9218));
  nand_5 g08842(.A(new_n9218), .B(new_n9216), .Y(new_n9219));
  xor_4  g08843(.A(new_n9219), .B(new_n9215), .Y(new_n9220));
  xor_4  g08844(.A(new_n9220), .B(new_n9212), .Y(new_n9221));
  xor_4  g08845(.A(new_n9221), .B(new_n9211), .Y(new_n9222));
  xor_4  g08846(.A(new_n9222), .B(new_n9206), .Y(new_n9223));
  xor_4  g08847(.A(new_n9223), .B(new_n9201), .Y(new_n9224));
  xor_4  g08848(.A(new_n9224), .B(new_n9198), .Y(new_n9225));
  nand_5 g08849(.A(pi191), .B(pi142), .Y(new_n9226));
  nand_5 g08850(.A(new_n8738), .B(new_n8737), .Y(new_n9227));
  nand_5 g08851(.A(new_n8739), .B(new_n8703), .Y(new_n9228));
  nand_5 g08852(.A(new_n9228), .B(new_n9227), .Y(new_n9229));
  xor_4  g08853(.A(new_n9229), .B(new_n9226), .Y(new_n9230));
  nand_5 g08854(.A(pi138), .B(pi017), .Y(new_n9231));
  nand_5 g08855(.A(new_n9145), .B(new_n9142), .Y(new_n9232));
  nand_5 g08856(.A(new_n9146), .B(new_n9138), .Y(new_n9233));
  nand_5 g08857(.A(new_n9233), .B(new_n9232), .Y(new_n9234));
  xor_4  g08858(.A(new_n9234), .B(new_n9231), .Y(new_n9235));
  nand_5 g08859(.A(new_n9140), .B(new_n9139), .Y(new_n9236));
  nand_5 g08860(.A(new_n9141), .B(new_n9116), .Y(new_n9237));
  nand_5 g08861(.A(new_n9237), .B(new_n9236), .Y(new_n9238));
  nand_5 g08862(.A(pi249), .B(pi192), .Y(new_n9239));
  or_6   g08863(.A(new_n8748), .B(new_n8704), .Y(new_n9240));
  nand_5 g08864(.A(new_n8749), .B(new_n8745), .Y(new_n9241));
  nand_5 g08865(.A(new_n9241), .B(new_n9240), .Y(new_n9242));
  xor_4  g08866(.A(new_n9242), .B(new_n9239), .Y(new_n9243));
  nand_5 g08867(.A(pi251), .B(pi222), .Y(new_n9244));
  xor_4  g08868(.A(new_n9244), .B(new_n9243), .Y(new_n9245));
  xor_4  g08869(.A(new_n9245), .B(new_n9238), .Y(new_n9246));
  xor_4  g08870(.A(new_n9246), .B(new_n9235), .Y(new_n9247));
  nand_5 g08871(.A(new_n9133), .B(new_n9132), .Y(new_n9248));
  nand_5 g08872(.A(new_n9134), .B(new_n9105), .Y(new_n9249));
  nand_5 g08873(.A(new_n9249), .B(new_n9248), .Y(new_n9250));
  or_6   g08874(.A(new_n9136), .B(new_n9106), .Y(new_n9251));
  not_8  g08875(.A(new_n9135), .Y(new_n9252));
  nand_5 g08876(.A(new_n9137), .B(new_n9252), .Y(new_n9253));
  nand_5 g08877(.A(new_n9253), .B(new_n9251), .Y(new_n9254));
  xor_4  g08878(.A(new_n9254), .B(new_n9250), .Y(new_n9255));
  xor_4  g08879(.A(new_n9255), .B(new_n9247), .Y(new_n9256));
  xor_4  g08880(.A(new_n9256), .B(new_n9230), .Y(new_n9257));
  or_6   g08881(.A(new_n9017), .B(new_n8769), .Y(new_n9258));
  nand_5 g08882(.A(new_n9056), .B(new_n9018), .Y(new_n9259));
  nand_5 g08883(.A(new_n9259), .B(new_n9258), .Y(new_n9260));
  nand_5 g08884(.A(pi122), .B(pi121), .Y(new_n9261));
  nand_5 g08885(.A(pi231), .B(pi001), .Y(new_n9262));
  xor_4  g08886(.A(new_n9262), .B(new_n9261), .Y(new_n9263));
  nand_5 g08887(.A(new_n8841), .B(new_n8838), .Y(new_n9264));
  nand_5 g08888(.A(new_n8842), .B(new_n8834), .Y(new_n9265));
  nand_5 g08889(.A(new_n9265), .B(new_n9264), .Y(new_n9266));
  nand_5 g08890(.A(pi224), .B(pi099), .Y(new_n9267));
  xor_4  g08891(.A(new_n9267), .B(new_n9266), .Y(new_n9268));
  nand_5 g08892(.A(new_n8829), .B(new_n8775), .Y(new_n9269));
  nand_5 g08893(.A(new_n8830), .B(new_n8828), .Y(new_n9270));
  nand_5 g08894(.A(new_n9270), .B(new_n9269), .Y(new_n9271));
  nand_5 g08895(.A(new_n8836), .B(new_n8835), .Y(new_n9272));
  nand_5 g08896(.A(new_n8837), .B(new_n8790), .Y(new_n9273));
  nand_5 g08897(.A(new_n9273), .B(new_n9272), .Y(new_n9274));
  nand_5 g08898(.A(pi255), .B(pi123), .Y(new_n9275));
  xor_4  g08899(.A(new_n9275), .B(new_n9274), .Y(new_n9276));
  xor_4  g08900(.A(new_n9276), .B(new_n9271), .Y(new_n9277));
  or_6   g08901(.A(new_n8832), .B(new_n8776), .Y(new_n9278));
  not_8  g08902(.A(new_n8831), .Y(new_n9279));
  nand_5 g08903(.A(new_n8833), .B(new_n9279), .Y(new_n9280));
  nand_5 g08904(.A(new_n9280), .B(new_n9278), .Y(new_n9281));
  nand_5 g08905(.A(pi232), .B(pi071), .Y(new_n9282));
  nand_5 g08906(.A(pi169), .B(pi127), .Y(new_n9283));
  xor_4  g08907(.A(new_n9283), .B(new_n9282), .Y(new_n9284));
  xor_4  g08908(.A(new_n9284), .B(new_n9281), .Y(new_n9285));
  xor_4  g08909(.A(new_n9285), .B(new_n9277), .Y(new_n9286));
  xor_4  g08910(.A(new_n9286), .B(new_n9268), .Y(new_n9287));
  xor_4  g08911(.A(new_n9287), .B(new_n9263), .Y(new_n9288));
  xor_4  g08912(.A(new_n9288), .B(new_n9260), .Y(new_n9289));
  nand_5 g08913(.A(new_n8926), .B(new_n8905), .Y(new_n9290));
  nand_5 g08914(.A(new_n8927), .B(new_n8903), .Y(new_n9291));
  nand_5 g08915(.A(new_n9291), .B(new_n9290), .Y(new_n9292));
  nand_5 g08916(.A(pi087), .B(pi082), .Y(new_n9293));
  xor_4  g08917(.A(new_n9293), .B(new_n9292), .Y(new_n9294));
  and_6  g08918(.A(new_n8972), .B(new_n8928), .Y(new_n9295));
  or_6   g08919(.A(new_n9295), .B(new_n8971), .Y(new_n9296));
  nand_5 g08920(.A(pi140), .B(pi059), .Y(new_n9297));
  nand_5 g08921(.A(pi242), .B(pi094), .Y(new_n9298));
  xor_4  g08922(.A(new_n9298), .B(new_n9297), .Y(new_n9299));
  xor_4  g08923(.A(new_n9299), .B(new_n9296), .Y(new_n9300));
  xor_4  g08924(.A(new_n9300), .B(new_n9294), .Y(new_n9301));
  nand_5 g08925(.A(pi252), .B(pi135), .Y(new_n9302));
  nand_5 g08926(.A(pi217), .B(pi137), .Y(new_n9303));
  nand_5 g08927(.A(pi160), .B(pi129), .Y(new_n9304));
  xor_4  g08928(.A(new_n9304), .B(new_n9303), .Y(new_n9305));
  or_6   g08929(.A(new_n8900), .B(new_n8885), .Y(new_n9306));
  nand_5 g08930(.A(new_n8901), .B(new_n8880), .Y(new_n9307));
  nand_5 g08931(.A(new_n9307), .B(new_n9306), .Y(new_n9308));
  nand_5 g08932(.A(pi219), .B(pi021), .Y(new_n9309));
  nand_5 g08933(.A(pi102), .B(pi005), .Y(new_n9310));
  xor_4  g08934(.A(new_n9310), .B(new_n9309), .Y(new_n9311));
  xor_4  g08935(.A(new_n9311), .B(new_n9308), .Y(new_n9312));
  xor_4  g08936(.A(new_n9312), .B(new_n9305), .Y(new_n9313));
  nand_5 g08937(.A(new_n9149), .B(new_n9117), .Y(new_n9314));
  not_8  g08938(.A(new_n9151), .Y(new_n9315));
  nand_5 g08939(.A(new_n9315), .B(new_n9147), .Y(new_n9316));
  nand_5 g08940(.A(new_n9316), .B(new_n9314), .Y(new_n9317));
  nand_5 g08941(.A(new_n8872), .B(new_n8871), .Y(new_n9318));
  nand_5 g08942(.A(new_n8873), .B(new_n8870), .Y(new_n9319));
  nand_5 g08943(.A(new_n9319), .B(new_n9318), .Y(new_n9320));
  nand_5 g08944(.A(new_n8883), .B(new_n8882), .Y(new_n9321));
  nand_5 g08945(.A(new_n8884), .B(new_n8881), .Y(new_n9322));
  nand_5 g08946(.A(new_n9322), .B(new_n9321), .Y(new_n9323));
  xnor_4 g08947(.A(new_n9323), .B(new_n9320), .Y(new_n9324));
  or_6   g08948(.A(new_n8878), .B(new_n8876), .Y(new_n9325));
  nand_5 g08949(.A(new_n8879), .B(new_n8875), .Y(new_n9326));
  nand_5 g08950(.A(new_n9326), .B(new_n9325), .Y(new_n9327));
  xor_4  g08951(.A(new_n9327), .B(new_n9324), .Y(new_n9328));
  xor_4  g08952(.A(new_n9328), .B(new_n9317), .Y(new_n9329));
  xor_4  g08953(.A(new_n9329), .B(new_n9313), .Y(new_n9330));
  xor_4  g08954(.A(new_n9330), .B(new_n9302), .Y(new_n9331));
  xor_4  g08955(.A(new_n9331), .B(new_n9301), .Y(new_n9332));
  xor_4  g08956(.A(new_n9332), .B(new_n9289), .Y(new_n9333));
  nand_5 g08957(.A(pi177), .B(pi100), .Y(new_n9334));
  nor_5  g08958(.A(new_n8750), .B(new_n8728), .Y(new_n9335));
  nor_5  g08959(.A(new_n8768), .B(new_n8751), .Y(new_n9336));
  or_6   g08960(.A(new_n9336), .B(new_n9335), .Y(new_n9337));
  nand_5 g08961(.A(pi101), .B(pi081), .Y(new_n9338));
  nand_5 g08962(.A(pi223), .B(pi106), .Y(new_n9339));
  xor_4  g08963(.A(new_n9339), .B(new_n9338), .Y(new_n9340));
  xor_4  g08964(.A(new_n9340), .B(new_n9337), .Y(new_n9341));
  xor_4  g08965(.A(new_n9341), .B(new_n9334), .Y(new_n9342));
  nand_5 g08966(.A(pi227), .B(pi225), .Y(new_n9343));
  nand_5 g08967(.A(pi187), .B(pi020), .Y(new_n9344));
  nand_5 g08968(.A(pi233), .B(pi060), .Y(new_n9345));
  xor_4  g08969(.A(new_n9345), .B(new_n9344), .Y(new_n9346));
  xor_4  g08970(.A(new_n9346), .B(new_n9343), .Y(new_n9347));
  xor_4  g08971(.A(new_n9347), .B(new_n9342), .Y(new_n9348));
  xor_4  g08972(.A(new_n9348), .B(new_n9333), .Y(new_n9349));
  xor_4  g08973(.A(new_n9349), .B(new_n9257), .Y(new_n9350));
  nand_5 g08974(.A(pi210), .B(pi086), .Y(new_n9351));
  or_6   g08975(.A(new_n8849), .B(new_n8843), .Y(new_n9352));
  nand_5 g08976(.A(new_n9352), .B(new_n8848), .Y(new_n9353));
  nor_5  g08977(.A(new_n8850), .B(new_n8827), .Y(new_n9354));
  nor_5  g08978(.A(new_n8868), .B(new_n8851), .Y(new_n9355));
  nor_5  g08979(.A(new_n9355), .B(new_n9354), .Y(new_n9356));
  nand_5 g08980(.A(new_n8974), .B(new_n8869), .Y(new_n9357));
  nand_5 g08981(.A(new_n9016), .B(new_n8975), .Y(new_n9358));
  nand_5 g08982(.A(new_n9358), .B(new_n9357), .Y(new_n9359));
  xor_4  g08983(.A(new_n9359), .B(new_n9356), .Y(new_n9360));
  xor_4  g08984(.A(new_n9360), .B(new_n9353), .Y(new_n9361));
  xor_4  g08985(.A(new_n9361), .B(new_n9351), .Y(new_n9362));
  xor_4  g08986(.A(new_n9362), .B(new_n9350), .Y(new_n9363));
  xor_4  g08987(.A(new_n9363), .B(new_n9225), .Y(po051));
  xor_4  g08988(.A(new_n3251), .B(new_n3234), .Y(po052));
  xor_4  g08989(.A(new_n3492), .B(new_n3452), .Y(po053));
  xor_4  g08990(.A(new_n872), .B(new_n846), .Y(po054));
  xor_4  g08991(.A(new_n7530), .B(new_n7516), .Y(po055));
  xor_4  g08992(.A(new_n3938), .B(new_n3937), .Y(po056));
  xor_4  g08993(.A(new_n1809), .B(new_n1807), .Y(po057));
  xor_4  g08994(.A(new_n3750), .B(new_n3749), .Y(po058));
  xor_4  g08995(.A(new_n5356), .B(new_n5354), .Y(po059));
  xor_4  g08996(.A(new_n2571), .B(new_n2547), .Y(po060));
  xor_4  g08997(.A(new_n2567), .B(new_n2566), .Y(po061));
  nand_5 g08998(.A(new_n8659), .B(new_n8656), .Y(new_n9375));
  nand_5 g08999(.A(new_n8660), .B(new_n8655), .Y(new_n9376));
  nand_5 g09000(.A(new_n9376), .B(new_n9375), .Y(new_n9377));
  nand_5 g09001(.A(pi227), .B(pi133), .Y(new_n9378));
  nand_5 g09002(.A(new_n8653), .B(new_n8652), .Y(new_n9379));
  nand_5 g09003(.A(new_n8654), .B(new_n8651), .Y(new_n9380));
  nand_5 g09004(.A(new_n9380), .B(new_n9379), .Y(new_n9381));
  nand_5 g09005(.A(pi189), .B(pi100), .Y(new_n9382));
  nand_5 g09006(.A(pi217), .B(pi064), .Y(new_n9383));
  nand_5 g09007(.A(new_n9383), .B(new_n9382), .Y(new_n9384));
  nand_5 g09008(.A(pi100), .B(pi064), .Y(new_n9385));
  or_6   g09009(.A(new_n9385), .B(new_n8653), .Y(new_n9386));
  nand_5 g09010(.A(new_n9386), .B(new_n9384), .Y(new_n9387));
  xor_4  g09011(.A(new_n9387), .B(new_n9381), .Y(new_n9388));
  xor_4  g09012(.A(new_n9388), .B(new_n9378), .Y(new_n9389));
  nand_5 g09013(.A(pi081), .B(pi077), .Y(new_n9390));
  nand_5 g09014(.A(pi106), .B(pi052), .Y(new_n9391));
  nand_5 g09015(.A(new_n9391), .B(new_n9390), .Y(new_n9392));
  nand_5 g09016(.A(pi106), .B(pi077), .Y(new_n9393));
  or_6   g09017(.A(new_n9393), .B(new_n8656), .Y(new_n9394));
  nand_5 g09018(.A(new_n9394), .B(new_n9392), .Y(new_n9395));
  xor_4  g09019(.A(new_n9395), .B(new_n9389), .Y(new_n9396));
  xor_4  g09020(.A(new_n9396), .B(new_n9377), .Y(new_n9397));
  not_8  g09021(.A(new_n9397), .Y(new_n9398));
  or_6   g09022(.A(new_n8649), .B(new_n8646), .Y(new_n9399));
  nand_5 g09023(.A(new_n8661), .B(new_n8650), .Y(new_n9400));
  nand_5 g09024(.A(new_n9400), .B(new_n9399), .Y(new_n9401));
  nand_5 g09025(.A(new_n9401), .B(new_n9398), .Y(new_n9402));
  nand_5 g09026(.A(new_n9395), .B(new_n9389), .Y(new_n9403));
  nand_5 g09027(.A(new_n9396), .B(new_n9377), .Y(new_n9404));
  nand_5 g09028(.A(new_n9404), .B(new_n9403), .Y(new_n9405));
  xor_4  g09029(.A(new_n9405), .B(new_n9394), .Y(new_n9406));
  nand_5 g09030(.A(pi227), .B(pi189), .Y(new_n9407));
  nand_5 g09031(.A(pi217), .B(pi084), .Y(new_n9408));
  xor_4  g09032(.A(new_n9408), .B(new_n9407), .Y(new_n9409));
  xor_4  g09033(.A(new_n9409), .B(new_n9385), .Y(new_n9410));
  nand_5 g09034(.A(pi133), .B(pi081), .Y(new_n9411));
  xor_4  g09035(.A(new_n9411), .B(new_n9386), .Y(new_n9412));
  xor_4  g09036(.A(new_n9412), .B(new_n9410), .Y(new_n9413));
  nand_5 g09037(.A(pi187), .B(pi131), .Y(new_n9414));
  nand_5 g09038(.A(pi233), .B(pi052), .Y(new_n9415));
  xor_4  g09039(.A(new_n9415), .B(new_n9414), .Y(new_n9416));
  xor_4  g09040(.A(new_n9416), .B(new_n9393), .Y(new_n9417));
  nand_5 g09041(.A(new_n9387), .B(new_n9381), .Y(new_n9418));
  nand_5 g09042(.A(new_n9388), .B(new_n9378), .Y(new_n9419));
  nand_5 g09043(.A(new_n9419), .B(new_n9418), .Y(new_n9420));
  xor_4  g09044(.A(new_n9420), .B(new_n9417), .Y(new_n9421));
  xor_4  g09045(.A(new_n9421), .B(new_n9413), .Y(new_n9422));
  xor_4  g09046(.A(new_n9422), .B(new_n9406), .Y(new_n9423));
  nand_5 g09047(.A(new_n8662), .B(new_n8645), .Y(new_n9424));
  nand_5 g09048(.A(pi233), .B(pi131), .Y(new_n9425));
  nand_5 g09049(.A(new_n9425), .B(new_n9424), .Y(new_n9426));
  xor_4  g09050(.A(new_n9401), .B(new_n9397), .Y(new_n9427));
  xor_4  g09051(.A(new_n9425), .B(new_n9424), .Y(new_n9428));
  nand_5 g09052(.A(new_n9428), .B(new_n9427), .Y(new_n9429));
  nand_5 g09053(.A(new_n9429), .B(new_n9426), .Y(new_n9430));
  xnor_4 g09054(.A(new_n9430), .B(new_n9423), .Y(new_n9431));
  xor_4  g09055(.A(new_n9431), .B(new_n9402), .Y(new_n9432));
  nand_5 g09056(.A(pi125), .B(pi035), .Y(new_n9433));
  nand_5 g09057(.A(new_n8624), .B(new_n8623), .Y(new_n9434));
  nand_5 g09058(.A(new_n8625), .B(new_n8622), .Y(new_n9435));
  nand_5 g09059(.A(new_n9435), .B(new_n9434), .Y(new_n9436));
  nand_5 g09060(.A(pi249), .B(pi204), .Y(new_n9437));
  nand_5 g09061(.A(pi222), .B(pi015), .Y(new_n9438));
  nand_5 g09062(.A(new_n9438), .B(new_n9437), .Y(new_n9439));
  nand_5 g09063(.A(pi222), .B(pi204), .Y(new_n9440));
  or_6   g09064(.A(new_n9440), .B(new_n8622), .Y(new_n9441));
  nand_5 g09065(.A(new_n9441), .B(new_n9439), .Y(new_n9442));
  xor_4  g09066(.A(new_n9442), .B(new_n9436), .Y(new_n9443));
  xor_4  g09067(.A(new_n9443), .B(new_n9433), .Y(new_n9444));
  nand_5 g09068(.A(new_n8630), .B(new_n8627), .Y(new_n9445));
  nand_5 g09069(.A(new_n8631), .B(new_n8626), .Y(new_n9446));
  nand_5 g09070(.A(new_n9446), .B(new_n9445), .Y(new_n9447));
  nand_5 g09071(.A(new_n9447), .B(new_n9444), .Y(new_n9448));
  or_6   g09072(.A(new_n9447), .B(new_n9444), .Y(new_n9449));
  and_6  g09073(.A(new_n9449), .B(new_n9448), .Y(new_n9450));
  nand_5 g09074(.A(pi176), .B(pi139), .Y(new_n9451));
  nand_5 g09075(.A(pi208), .B(pi040), .Y(new_n9452));
  nand_5 g09076(.A(new_n9452), .B(new_n9451), .Y(new_n9453));
  nand_5 g09077(.A(pi139), .B(pi040), .Y(new_n9454));
  or_6   g09078(.A(new_n9454), .B(new_n8627), .Y(new_n9455));
  nand_5 g09079(.A(new_n9455), .B(new_n9453), .Y(new_n9456));
  xor_4  g09080(.A(new_n9456), .B(new_n9450), .Y(new_n9457));
  not_8  g09081(.A(new_n9457), .Y(new_n9458));
  or_6   g09082(.A(new_n8636), .B(new_n8633), .Y(new_n9459));
  nand_5 g09083(.A(new_n8637), .B(new_n8632), .Y(new_n9460));
  nand_5 g09084(.A(new_n9460), .B(new_n9459), .Y(new_n9461));
  nand_5 g09085(.A(new_n9461), .B(new_n9458), .Y(new_n9462));
  nand_5 g09086(.A(pi249), .B(pi146), .Y(new_n9463));
  nand_5 g09087(.A(pi125), .B(pi015), .Y(new_n9464));
  xor_4  g09088(.A(new_n9464), .B(new_n9463), .Y(new_n9465));
  xor_4  g09089(.A(new_n9465), .B(new_n9440), .Y(new_n9466));
  nand_5 g09090(.A(pi176), .B(pi035), .Y(new_n9467));
  xor_4  g09091(.A(new_n9467), .B(new_n9441), .Y(new_n9468));
  xor_4  g09092(.A(new_n9468), .B(new_n9466), .Y(new_n9469));
  nand_5 g09093(.A(pi208), .B(pi174), .Y(new_n9470));
  nand_5 g09094(.A(pi168), .B(pi157), .Y(new_n9471));
  xor_4  g09095(.A(new_n9471), .B(new_n9470), .Y(new_n9472));
  xor_4  g09096(.A(new_n9472), .B(new_n9454), .Y(new_n9473));
  nand_5 g09097(.A(new_n9442), .B(new_n9436), .Y(new_n9474));
  nand_5 g09098(.A(new_n9443), .B(new_n9433), .Y(new_n9475));
  nand_5 g09099(.A(new_n9475), .B(new_n9474), .Y(new_n9476));
  xor_4  g09100(.A(new_n9476), .B(new_n9473), .Y(new_n9477));
  xor_4  g09101(.A(new_n9477), .B(new_n9469), .Y(new_n9478));
  nand_5 g09102(.A(new_n9456), .B(new_n9450), .Y(new_n9479));
  nand_5 g09103(.A(new_n9479), .B(new_n9448), .Y(new_n9480));
  and_6  g09104(.A(new_n9480), .B(new_n9455), .Y(new_n9481));
  nor_5  g09105(.A(new_n9455), .B(new_n9449), .Y(new_n9482));
  or_6   g09106(.A(new_n9482), .B(new_n9481), .Y(new_n9483));
  xnor_4 g09107(.A(new_n9483), .B(new_n9478), .Y(new_n9484));
  xor_4  g09108(.A(new_n9484), .B(new_n9462), .Y(new_n9485));
  nand_5 g09109(.A(pi174), .B(pi168), .Y(new_n9486));
  xor_4  g09110(.A(new_n9461), .B(new_n9457), .Y(new_n9487));
  or_6   g09111(.A(new_n9487), .B(new_n9486), .Y(new_n9488));
  nor_5  g09112(.A(new_n8638), .B(new_n8621), .Y(new_n9489));
  xor_4  g09113(.A(new_n9487), .B(new_n9486), .Y(new_n9490));
  nand_5 g09114(.A(new_n9490), .B(new_n9489), .Y(new_n9491));
  nand_5 g09115(.A(new_n9491), .B(new_n9488), .Y(new_n9492));
  xnor_4 g09116(.A(new_n9492), .B(new_n9485), .Y(new_n9493));
  xor_4  g09117(.A(new_n9490), .B(new_n9489), .Y(new_n9494));
  nand_5 g09118(.A(new_n8642), .B(new_n8639), .Y(new_n9495));
  nand_5 g09119(.A(new_n8643), .B(new_n8620), .Y(new_n9496));
  nand_5 g09120(.A(new_n9496), .B(new_n9495), .Y(new_n9497));
  or_6   g09121(.A(new_n9497), .B(new_n9494), .Y(new_n9498));
  xor_4  g09122(.A(new_n9497), .B(new_n9494), .Y(new_n9499));
  nand_5 g09123(.A(new_n8594), .B(new_n8577), .Y(new_n9500));
  nand_5 g09124(.A(pi252), .B(pi141), .Y(new_n9501));
  nand_5 g09125(.A(pi140), .B(pi090), .Y(new_n9502));
  nand_5 g09126(.A(pi242), .B(pi047), .Y(new_n9503));
  nand_5 g09127(.A(new_n9503), .B(new_n9502), .Y(new_n9504));
  nand_5 g09128(.A(pi140), .B(pi047), .Y(new_n9505));
  or_6   g09129(.A(new_n9505), .B(new_n8579), .Y(new_n9506));
  nand_5 g09130(.A(new_n9506), .B(new_n9504), .Y(new_n9507));
  xor_4  g09131(.A(new_n9507), .B(new_n9501), .Y(new_n9508));
  nand_5 g09132(.A(new_n8580), .B(new_n8579), .Y(new_n9509));
  nand_5 g09133(.A(new_n8581), .B(new_n8578), .Y(new_n9510));
  nand_5 g09134(.A(new_n9510), .B(new_n9509), .Y(new_n9511));
  xor_4  g09135(.A(new_n9511), .B(new_n9508), .Y(new_n9512));
  nand_5 g09136(.A(pi161), .B(pi121), .Y(new_n9513));
  nand_5 g09137(.A(pi241), .B(pi231), .Y(new_n9514));
  and_6  g09138(.A(new_n9514), .B(new_n9513), .Y(new_n9515));
  nand_5 g09139(.A(pi231), .B(pi161), .Y(new_n9516));
  nor_5  g09140(.A(new_n9516), .B(new_n8583), .Y(new_n9517));
  or_6   g09141(.A(new_n9517), .B(new_n9515), .Y(new_n9518));
  xnor_4 g09142(.A(new_n9518), .B(new_n9512), .Y(new_n9519));
  nand_5 g09143(.A(new_n8586), .B(new_n8583), .Y(new_n9520));
  nand_5 g09144(.A(new_n8587), .B(new_n8582), .Y(new_n9521));
  nand_5 g09145(.A(new_n9521), .B(new_n9520), .Y(new_n9522));
  xor_4  g09146(.A(new_n9522), .B(new_n9519), .Y(new_n9523));
  not_8  g09147(.A(new_n8589), .Y(new_n9524));
  nand_5 g09148(.A(new_n8592), .B(new_n9524), .Y(new_n9525));
  or_6   g09149(.A(new_n8593), .B(new_n8588), .Y(new_n9526));
  nand_5 g09150(.A(new_n9526), .B(new_n9525), .Y(new_n9527));
  xnor_4 g09151(.A(new_n9527), .B(new_n9523), .Y(new_n9528));
  nand_5 g09152(.A(pi236), .B(pi005), .Y(new_n9529));
  xor_4  g09153(.A(new_n9529), .B(new_n9528), .Y(new_n9530));
  xor_4  g09154(.A(new_n9530), .B(new_n9500), .Y(new_n9531));
  nand_5 g09155(.A(new_n8605), .B(new_n8602), .Y(new_n9532));
  nand_5 g09156(.A(new_n8606), .B(new_n8601), .Y(new_n9533));
  nand_5 g09157(.A(new_n9533), .B(new_n9532), .Y(new_n9534));
  nand_5 g09158(.A(pi024), .B(pi013), .Y(new_n9535));
  nand_5 g09159(.A(new_n8599), .B(new_n8598), .Y(new_n9536));
  nand_5 g09160(.A(new_n8600), .B(new_n8597), .Y(new_n9537));
  nand_5 g09161(.A(new_n9537), .B(new_n9536), .Y(new_n9538));
  nand_5 g09162(.A(pi112), .B(pi111), .Y(new_n9539));
  nand_5 g09163(.A(pi210), .B(pi105), .Y(new_n9540));
  nand_5 g09164(.A(new_n9540), .B(new_n9539), .Y(new_n9541));
  nand_5 g09165(.A(pi111), .B(pi105), .Y(new_n9542));
  or_6   g09166(.A(new_n9542), .B(new_n8598), .Y(new_n9543));
  nand_5 g09167(.A(new_n9543), .B(new_n9541), .Y(new_n9544));
  xor_4  g09168(.A(new_n9544), .B(new_n9538), .Y(new_n9545));
  xor_4  g09169(.A(new_n9545), .B(new_n9535), .Y(new_n9546));
  nand_5 g09170(.A(pi224), .B(pi104), .Y(new_n9547));
  nand_5 g09171(.A(pi255), .B(pi212), .Y(new_n9548));
  nand_5 g09172(.A(new_n9548), .B(new_n9547), .Y(new_n9549));
  nand_5 g09173(.A(pi255), .B(pi104), .Y(new_n9550));
  or_6   g09174(.A(new_n9550), .B(new_n8602), .Y(new_n9551));
  nand_5 g09175(.A(new_n9551), .B(new_n9549), .Y(new_n9552));
  xor_4  g09176(.A(new_n9552), .B(new_n9546), .Y(new_n9553));
  xor_4  g09177(.A(new_n9553), .B(new_n9534), .Y(new_n9554));
  or_6   g09178(.A(new_n8611), .B(new_n8608), .Y(new_n9555));
  nand_5 g09179(.A(new_n8612), .B(new_n8607), .Y(new_n9556));
  nand_5 g09180(.A(new_n9556), .B(new_n9555), .Y(new_n9557));
  xor_4  g09181(.A(new_n9557), .B(new_n9554), .Y(new_n9558));
  nand_5 g09182(.A(new_n8613), .B(new_n8596), .Y(new_n9559));
  nand_5 g09183(.A(pi213), .B(pi127), .Y(new_n9560));
  xor_4  g09184(.A(new_n9560), .B(new_n9559), .Y(new_n9561));
  xor_4  g09185(.A(new_n9561), .B(new_n9558), .Y(new_n9562));
  xor_4  g09186(.A(new_n9562), .B(new_n9531), .Y(new_n9563));
  nand_5 g09187(.A(new_n8618), .B(new_n8614), .Y(new_n9564));
  not_8  g09188(.A(new_n8595), .Y(new_n9565));
  nand_5 g09189(.A(new_n8619), .B(new_n9565), .Y(new_n9566));
  nand_5 g09190(.A(new_n9566), .B(new_n9564), .Y(new_n9567));
  xor_4  g09191(.A(new_n9567), .B(new_n9563), .Y(new_n9568));
  nand_5 g09192(.A(new_n9568), .B(new_n9499), .Y(new_n9569));
  nand_5 g09193(.A(new_n9569), .B(new_n9498), .Y(new_n9570));
  xor_4  g09194(.A(new_n9570), .B(new_n9493), .Y(new_n9571));
  not_8  g09195(.A(new_n9571), .Y(new_n9572));
  not_8  g09196(.A(new_n9554), .Y(new_n9573));
  nand_5 g09197(.A(new_n9557), .B(new_n9573), .Y(new_n9574));
  nand_5 g09198(.A(pi210), .B(pi183), .Y(new_n9575));
  nand_5 g09199(.A(pi112), .B(pi024), .Y(new_n9576));
  xor_4  g09200(.A(new_n9576), .B(new_n9575), .Y(new_n9577));
  xor_4  g09201(.A(new_n9577), .B(new_n9542), .Y(new_n9578));
  not_8  g09202(.A(new_n9578), .Y(new_n9579));
  nand_5 g09203(.A(pi224), .B(pi013), .Y(new_n9580));
  xor_4  g09204(.A(new_n9580), .B(new_n9543), .Y(new_n9581));
  xor_4  g09205(.A(new_n9581), .B(new_n9579), .Y(new_n9582));
  nand_5 g09206(.A(pi212), .B(pi127), .Y(new_n9583));
  nand_5 g09207(.A(pi232), .B(pi213), .Y(new_n9584));
  xor_4  g09208(.A(new_n9584), .B(new_n9583), .Y(new_n9585));
  xor_4  g09209(.A(new_n9585), .B(new_n9550), .Y(new_n9586));
  nand_5 g09210(.A(new_n9544), .B(new_n9538), .Y(new_n9587));
  nand_5 g09211(.A(new_n9545), .B(new_n9535), .Y(new_n9588));
  nand_5 g09212(.A(new_n9588), .B(new_n9587), .Y(new_n9589));
  xor_4  g09213(.A(new_n9589), .B(new_n9586), .Y(new_n9590));
  xor_4  g09214(.A(new_n9590), .B(new_n9582), .Y(new_n9591));
  nand_5 g09215(.A(new_n9552), .B(new_n9546), .Y(new_n9592));
  nand_5 g09216(.A(new_n9553), .B(new_n9534), .Y(new_n9593));
  nand_5 g09217(.A(new_n9593), .B(new_n9592), .Y(new_n9594));
  xor_4  g09218(.A(new_n9594), .B(new_n9551), .Y(new_n9595));
  xnor_4 g09219(.A(new_n9595), .B(new_n9591), .Y(new_n9596));
  xnor_4 g09220(.A(new_n9596), .B(new_n9574), .Y(new_n9597));
  nand_5 g09221(.A(new_n9560), .B(new_n9559), .Y(new_n9598));
  nand_5 g09222(.A(new_n9561), .B(new_n9558), .Y(new_n9599));
  nand_5 g09223(.A(new_n9599), .B(new_n9598), .Y(new_n9600));
  xnor_4 g09224(.A(new_n9600), .B(new_n9597), .Y(new_n9601));
  nand_5 g09225(.A(new_n9527), .B(new_n9523), .Y(new_n9602));
  nand_5 g09226(.A(pi242), .B(pi018), .Y(new_n9603));
  nand_5 g09227(.A(pi252), .B(pi090), .Y(new_n9604));
  xor_4  g09228(.A(new_n9604), .B(new_n9603), .Y(new_n9605));
  xor_4  g09229(.A(new_n9605), .B(new_n9505), .Y(new_n9606));
  not_8  g09230(.A(new_n9606), .Y(new_n9607));
  nand_5 g09231(.A(pi141), .B(pi121), .Y(new_n9608));
  xor_4  g09232(.A(new_n9608), .B(new_n9506), .Y(new_n9609));
  xor_4  g09233(.A(new_n9609), .B(new_n9607), .Y(new_n9610));
  nand_5 g09234(.A(pi236), .B(pi021), .Y(new_n9611));
  nand_5 g09235(.A(pi241), .B(pi005), .Y(new_n9612));
  xor_4  g09236(.A(new_n9612), .B(new_n9611), .Y(new_n9613));
  xor_4  g09237(.A(new_n9613), .B(new_n9516), .Y(new_n9614));
  nand_5 g09238(.A(new_n9507), .B(new_n9501), .Y(new_n9615));
  nand_5 g09239(.A(new_n9511), .B(new_n9508), .Y(new_n9616));
  nand_5 g09240(.A(new_n9616), .B(new_n9615), .Y(new_n9617));
  xor_4  g09241(.A(new_n9617), .B(new_n9614), .Y(new_n9618));
  xor_4  g09242(.A(new_n9618), .B(new_n9610), .Y(new_n9619));
  nor_5  g09243(.A(new_n9522), .B(new_n9519), .Y(new_n9620));
  nand_5 g09244(.A(new_n9620), .B(new_n9517), .Y(new_n9621));
  nor_5  g09245(.A(new_n9518), .B(new_n9512), .Y(new_n9622));
  or_6   g09246(.A(new_n9622), .B(new_n9517), .Y(new_n9623));
  or_6   g09247(.A(new_n9623), .B(new_n9620), .Y(new_n9624));
  nand_5 g09248(.A(new_n9624), .B(new_n9621), .Y(new_n9625));
  xor_4  g09249(.A(new_n9625), .B(new_n9619), .Y(new_n9626));
  xor_4  g09250(.A(new_n9626), .B(new_n9602), .Y(new_n9627));
  or_6   g09251(.A(new_n9529), .B(new_n9528), .Y(new_n9628));
  not_8  g09252(.A(new_n9500), .Y(new_n9629));
  nand_5 g09253(.A(new_n9530), .B(new_n9629), .Y(new_n9630));
  nand_5 g09254(.A(new_n9630), .B(new_n9628), .Y(new_n9631));
  xor_4  g09255(.A(new_n9631), .B(new_n9627), .Y(new_n9632));
  not_8  g09256(.A(new_n9632), .Y(new_n9633));
  xor_4  g09257(.A(new_n9633), .B(new_n9601), .Y(new_n9634));
  nand_5 g09258(.A(new_n9562), .B(new_n9531), .Y(new_n9635));
  nand_5 g09259(.A(new_n9567), .B(new_n9563), .Y(new_n9636));
  nand_5 g09260(.A(new_n9636), .B(new_n9635), .Y(new_n9637));
  xor_4  g09261(.A(new_n9637), .B(new_n9634), .Y(new_n9638));
  xor_4  g09262(.A(new_n9638), .B(new_n9572), .Y(new_n9639));
  xor_4  g09263(.A(new_n9639), .B(new_n9432), .Y(new_n9640));
  xor_4  g09264(.A(new_n9428), .B(new_n9427), .Y(new_n9641));
  nand_5 g09265(.A(new_n8664), .B(new_n8644), .Y(new_n9642));
  nand_5 g09266(.A(new_n8669), .B(new_n8665), .Y(new_n9643));
  nand_5 g09267(.A(new_n9643), .B(new_n9642), .Y(new_n9644));
  or_6   g09268(.A(new_n9644), .B(new_n9641), .Y(new_n9645));
  xnor_4 g09269(.A(new_n9568), .B(new_n9499), .Y(new_n9646));
  xor_4  g09270(.A(new_n9644), .B(new_n9641), .Y(new_n9647));
  nand_5 g09271(.A(new_n9647), .B(new_n9646), .Y(new_n9648));
  nand_5 g09272(.A(new_n9648), .B(new_n9645), .Y(new_n9649));
  xor_4  g09273(.A(new_n9649), .B(new_n9640), .Y(po062));
  xor_4  g09274(.A(new_n9165), .B(new_n9164), .Y(po063));
  nor_5  g09275(.A(new_n3080), .B(new_n2978), .Y(new_n9652));
  not_8  g09276(.A(new_n3081), .Y(new_n9653));
  nor_5  g09277(.A(new_n3118), .B(new_n9653), .Y(new_n9654));
  nor_5  g09278(.A(new_n9654), .B(new_n9652), .Y(new_n9655));
  nor_5  g09279(.A(new_n2875), .B(new_n2852), .Y(new_n9656));
  nor_5  g09280(.A(new_n2893), .B(new_n2876), .Y(new_n9657));
  nor_5  g09281(.A(new_n9657), .B(new_n9656), .Y(new_n9658));
  nand_5 g09282(.A(pi197), .B(pi182), .Y(new_n9659));
  nand_5 g09283(.A(new_n2654), .B(new_n2653), .Y(new_n9660));
  nand_5 g09284(.A(new_n2655), .B(new_n2601), .Y(new_n9661));
  nand_5 g09285(.A(new_n9661), .B(new_n9660), .Y(new_n9662));
  or_6   g09286(.A(new_n2667), .B(new_n2664), .Y(new_n9663));
  nand_5 g09287(.A(new_n2668), .B(new_n2660), .Y(new_n9664));
  nand_5 g09288(.A(new_n9664), .B(new_n9663), .Y(new_n9665));
  xor_4  g09289(.A(new_n9665), .B(new_n9662), .Y(new_n9666));
  xor_4  g09290(.A(new_n9666), .B(new_n9659), .Y(new_n9667));
  xor_4  g09291(.A(new_n9667), .B(new_n9658), .Y(new_n9668));
  xor_4  g09292(.A(new_n9668), .B(new_n9655), .Y(new_n9669));
  nand_5 g09293(.A(pi216), .B(pi198), .Y(new_n9670));
  nand_5 g09294(.A(new_n2894), .B(new_n2794), .Y(new_n9671));
  nand_5 g09295(.A(new_n2936), .B(new_n2895), .Y(new_n9672));
  nand_5 g09296(.A(new_n9672), .B(new_n9671), .Y(new_n9673));
  nand_5 g09297(.A(pi229), .B(pi225), .Y(new_n9674));
  nand_5 g09298(.A(pi030), .B(pi020), .Y(new_n9675));
  nand_5 g09299(.A(pi185), .B(pi060), .Y(new_n9676));
  xor_4  g09300(.A(new_n9676), .B(new_n9675), .Y(new_n9677));
  xor_4  g09301(.A(new_n9677), .B(new_n9674), .Y(new_n9678));
  xor_4  g09302(.A(new_n9678), .B(new_n9673), .Y(new_n9679));
  nand_5 g09303(.A(new_n3052), .B(new_n3051), .Y(new_n9680));
  nand_5 g09304(.A(new_n3053), .B(new_n3031), .Y(new_n9681));
  nand_5 g09305(.A(new_n9681), .B(new_n9680), .Y(new_n9682));
  nand_5 g09306(.A(pi101), .B(pi067), .Y(new_n9683));
  nand_5 g09307(.A(pi223), .B(pi053), .Y(new_n9684));
  xor_4  g09308(.A(new_n9684), .B(new_n9683), .Y(new_n9685));
  xor_4  g09309(.A(new_n9685), .B(new_n9682), .Y(new_n9686));
  nor_5  g09310(.A(new_n2676), .B(new_n2652), .Y(new_n9687));
  nor_5  g09311(.A(new_n2692), .B(new_n2677), .Y(new_n9688));
  or_6   g09312(.A(new_n9688), .B(new_n9687), .Y(new_n9689));
  nand_5 g09313(.A(pi177), .B(pi092), .Y(new_n9690));
  xor_4  g09314(.A(new_n9690), .B(new_n9689), .Y(new_n9691));
  xor_4  g09315(.A(new_n9691), .B(new_n9686), .Y(new_n9692));
  nand_5 g09316(.A(new_n3057), .B(new_n3054), .Y(new_n9693));
  nand_5 g09317(.A(new_n3058), .B(new_n3050), .Y(new_n9694));
  nand_5 g09318(.A(new_n9694), .B(new_n9693), .Y(new_n9695));
  nand_5 g09319(.A(pi251), .B(pi062), .Y(new_n9696));
  nand_5 g09320(.A(pi138), .B(pi078), .Y(new_n9697));
  xor_4  g09321(.A(new_n9697), .B(new_n9696), .Y(new_n9698));
  nand_5 g09322(.A(pi192), .B(pi065), .Y(new_n9699));
  or_6   g09323(.A(new_n2675), .B(new_n2669), .Y(new_n9700));
  nand_5 g09324(.A(new_n9700), .B(new_n2674), .Y(new_n9701));
  xor_4  g09325(.A(new_n9701), .B(new_n9699), .Y(new_n9702));
  xor_4  g09326(.A(new_n9702), .B(new_n9698), .Y(new_n9703));
  xor_4  g09327(.A(new_n9703), .B(new_n9695), .Y(new_n9704));
  nand_5 g09328(.A(new_n3045), .B(new_n3044), .Y(new_n9705));
  nand_5 g09329(.A(new_n3046), .B(new_n3019), .Y(new_n9706));
  nand_5 g09330(.A(new_n9706), .B(new_n9705), .Y(new_n9707));
  or_6   g09331(.A(new_n3048), .B(new_n3020), .Y(new_n9708));
  not_8  g09332(.A(new_n3047), .Y(new_n9709));
  nand_5 g09333(.A(new_n3049), .B(new_n9709), .Y(new_n9710));
  nand_5 g09334(.A(new_n9710), .B(new_n9708), .Y(new_n9711));
  xor_4  g09335(.A(new_n9711), .B(new_n9707), .Y(new_n9712));
  xor_4  g09336(.A(new_n9712), .B(new_n9704), .Y(new_n9713));
  xor_4  g09337(.A(new_n9713), .B(new_n9692), .Y(new_n9714));
  xor_4  g09338(.A(new_n9714), .B(new_n9679), .Y(new_n9715));
  xor_4  g09339(.A(new_n9715), .B(new_n9670), .Y(new_n9716));
  nor_5  g09340(.A(new_n2775), .B(new_n2751), .Y(new_n9717));
  nor_5  g09341(.A(new_n2793), .B(new_n2776), .Y(new_n9718));
  nor_5  g09342(.A(new_n9718), .B(new_n9717), .Y(new_n9719));
  nor_5  g09343(.A(new_n3060), .B(new_n3036), .Y(new_n9720));
  nor_5  g09344(.A(new_n3079), .B(new_n3061), .Y(new_n9721));
  nor_5  g09345(.A(new_n9721), .B(new_n9720), .Y(new_n9722));
  xor_4  g09346(.A(new_n9722), .B(new_n9719), .Y(new_n9723));
  nand_5 g09347(.A(new_n2753), .B(new_n2752), .Y(new_n9724));
  nand_5 g09348(.A(new_n2754), .B(new_n2706), .Y(new_n9725));
  nand_5 g09349(.A(new_n9725), .B(new_n9724), .Y(new_n9726));
  xor_4  g09350(.A(new_n9726), .B(new_n9723), .Y(new_n9727));
  nand_5 g09351(.A(pi219), .B(pi209), .Y(new_n9728));
  nor_5  g09352(.A(new_n2756), .B(new_n2708), .Y(new_n9729));
  nor_5  g09353(.A(new_n2758), .B(new_n2755), .Y(new_n9730));
  or_6   g09354(.A(new_n9730), .B(new_n9729), .Y(new_n9731));
  xor_4  g09355(.A(new_n9731), .B(new_n9728), .Y(new_n9732));
  nand_5 g09356(.A(pi130), .B(pi123), .Y(new_n9733));
  or_6   g09357(.A(new_n2774), .B(new_n2768), .Y(new_n9734));
  nand_5 g09358(.A(new_n9734), .B(new_n2773), .Y(new_n9735));
  nand_5 g09359(.A(pi154), .B(pi122), .Y(new_n9736));
  nand_5 g09360(.A(pi095), .B(pi001), .Y(new_n9737));
  xor_4  g09361(.A(new_n9737), .B(new_n9736), .Y(new_n9738));
  xor_4  g09362(.A(new_n9738), .B(new_n9735), .Y(new_n9739));
  nand_5 g09363(.A(pi135), .B(pi089), .Y(new_n9740));
  nand_5 g09364(.A(pi153), .B(pi087), .Y(new_n9741));
  nand_5 g09365(.A(pi158), .B(pi059), .Y(new_n9742));
  nand_5 g09366(.A(pi254), .B(pi094), .Y(new_n9743));
  xnor_4 g09367(.A(new_n9743), .B(new_n9742), .Y(new_n9744));
  xor_4  g09368(.A(new_n9744), .B(new_n9741), .Y(new_n9745));
  xor_4  g09369(.A(new_n9745), .B(new_n9740), .Y(new_n9746));
  xor_4  g09370(.A(new_n9746), .B(new_n9739), .Y(new_n9747));
  xor_4  g09371(.A(new_n9747), .B(new_n9733), .Y(new_n9748));
  nand_5 g09372(.A(new_n2854), .B(new_n2853), .Y(new_n9749));
  nand_5 g09373(.A(new_n2855), .B(new_n2820), .Y(new_n9750));
  nand_5 g09374(.A(new_n9750), .B(new_n9749), .Y(new_n9751));
  nand_5 g09375(.A(new_n2862), .B(new_n2861), .Y(new_n9752));
  nand_5 g09376(.A(new_n2863), .B(new_n2828), .Y(new_n9753));
  nand_5 g09377(.A(new_n9753), .B(new_n9752), .Y(new_n9754));
  nor_5  g09378(.A(new_n2857), .B(new_n2822), .Y(new_n9755));
  nor_5  g09379(.A(new_n2859), .B(new_n2856), .Y(new_n9756));
  or_6   g09380(.A(new_n9756), .B(new_n9755), .Y(new_n9757));
  xor_4  g09381(.A(new_n9757), .B(new_n9754), .Y(new_n9758));
  xor_4  g09382(.A(new_n9758), .B(new_n9751), .Y(new_n9759));
  nand_5 g09383(.A(pi215), .B(pi071), .Y(new_n9760));
  nand_5 g09384(.A(pi169), .B(pi124), .Y(new_n9761));
  xor_4  g09385(.A(new_n9761), .B(new_n9760), .Y(new_n9762));
  nand_5 g09386(.A(pi099), .B(pi003), .Y(new_n9763));
  xor_4  g09387(.A(new_n9763), .B(new_n9762), .Y(new_n9764));
  xor_4  g09388(.A(new_n9764), .B(new_n9759), .Y(new_n9765));
  xor_4  g09389(.A(new_n9765), .B(new_n9748), .Y(new_n9766));
  nand_5 g09390(.A(pi102), .B(pi006), .Y(new_n9767));
  nand_5 g09391(.A(pi190), .B(pi137), .Y(new_n9768));
  nand_5 g09392(.A(pi220), .B(pi160), .Y(new_n9769));
  xor_4  g09393(.A(new_n9769), .B(new_n9768), .Y(new_n9770));
  or_6   g09394(.A(new_n3059), .B(new_n3043), .Y(new_n9771));
  nand_5 g09395(.A(new_n9771), .B(new_n3040), .Y(new_n9772));
  xor_4  g09396(.A(new_n9772), .B(new_n9770), .Y(new_n9773));
  xor_4  g09397(.A(new_n9773), .B(new_n9767), .Y(new_n9774));
  xor_4  g09398(.A(new_n9774), .B(new_n9766), .Y(new_n9775));
  xor_4  g09399(.A(new_n9775), .B(new_n9732), .Y(new_n9776));
  or_6   g09400(.A(new_n2867), .B(new_n2864), .Y(new_n9777));
  nand_5 g09401(.A(new_n2868), .B(new_n2860), .Y(new_n9778));
  nand_5 g09402(.A(new_n9778), .B(new_n9777), .Y(new_n9779));
  nand_5 g09403(.A(new_n2761), .B(new_n2715), .Y(new_n9780));
  nand_5 g09404(.A(new_n2762), .B(new_n2760), .Y(new_n9781));
  nand_5 g09405(.A(new_n9781), .B(new_n9780), .Y(new_n9782));
  or_6   g09406(.A(new_n2766), .B(new_n2763), .Y(new_n9783));
  nand_5 g09407(.A(new_n2767), .B(new_n2759), .Y(new_n9784));
  nand_5 g09408(.A(new_n9784), .B(new_n9783), .Y(new_n9785));
  xor_4  g09409(.A(new_n9785), .B(new_n9782), .Y(new_n9786));
  xor_4  g09410(.A(new_n9786), .B(new_n9779), .Y(new_n9787));
  xor_4  g09411(.A(new_n9787), .B(new_n9776), .Y(new_n9788));
  xor_4  g09412(.A(new_n9788), .B(new_n9727), .Y(new_n9789));
  nand_5 g09413(.A(pi120), .B(pi079), .Y(new_n9790));
  nand_5 g09414(.A(pi172), .B(pi076), .Y(new_n9791));
  xor_4  g09415(.A(new_n9791), .B(new_n9790), .Y(new_n9792));
  nand_5 g09416(.A(new_n2873), .B(new_n2829), .Y(new_n9793));
  nand_5 g09417(.A(new_n2874), .B(new_n2870), .Y(new_n9794));
  nand_5 g09418(.A(new_n9794), .B(new_n9793), .Y(new_n9795));
  nand_5 g09419(.A(pi073), .B(pi023), .Y(new_n9796));
  nand_5 g09420(.A(pi155), .B(pi004), .Y(new_n9797));
  xor_4  g09421(.A(new_n9797), .B(new_n9796), .Y(new_n9798));
  xor_4  g09422(.A(new_n9798), .B(new_n9795), .Y(new_n9799));
  nand_5 g09423(.A(pi142), .B(pi022), .Y(new_n9800));
  nand_5 g09424(.A(new_n2662), .B(new_n2661), .Y(new_n9801));
  nand_5 g09425(.A(new_n2663), .B(new_n2616), .Y(new_n9802));
  nand_5 g09426(.A(new_n9802), .B(new_n9801), .Y(new_n9803));
  xor_4  g09427(.A(new_n9803), .B(new_n9800), .Y(new_n9804));
  nand_5 g09428(.A(pi170), .B(pi086), .Y(new_n9805));
  xor_4  g09429(.A(new_n9805), .B(new_n9804), .Y(new_n9806));
  xor_4  g09430(.A(new_n9806), .B(new_n9799), .Y(new_n9807));
  xor_4  g09431(.A(new_n9807), .B(new_n9792), .Y(new_n9808));
  xor_4  g09432(.A(new_n9808), .B(new_n9789), .Y(new_n9809));
  xor_4  g09433(.A(new_n9809), .B(new_n9716), .Y(new_n9810));
  or_6   g09434(.A(new_n2937), .B(new_n2693), .Y(new_n9811));
  nand_5 g09435(.A(new_n2977), .B(new_n2938), .Y(new_n9812));
  nand_5 g09436(.A(new_n9812), .B(new_n9811), .Y(new_n9813));
  nand_5 g09437(.A(pi165), .B(pi041), .Y(new_n9814));
  or_6   g09438(.A(new_n2658), .B(new_n2602), .Y(new_n9815));
  nand_5 g09439(.A(new_n2659), .B(new_n2657), .Y(new_n9816));
  nand_5 g09440(.A(new_n9816), .B(new_n9815), .Y(new_n9817));
  xor_4  g09441(.A(new_n9817), .B(new_n9814), .Y(new_n9818));
  xor_4  g09442(.A(new_n9818), .B(new_n9813), .Y(new_n9819));
  xor_4  g09443(.A(new_n9819), .B(new_n9810), .Y(new_n9820));
  xor_4  g09444(.A(new_n9820), .B(new_n9669), .Y(po064));
  xor_4  g09445(.A(new_n9176), .B(new_n9174), .Y(po065));
  xor_4  g09446(.A(new_n3103), .B(new_n3101), .Y(po066));
  xor_4  g09447(.A(new_n4992), .B(new_n4991), .Y(po067));
  xor_4  g09448(.A(new_n6950), .B(new_n6949), .Y(po068));
  xor_4  g09449(.A(new_n3824), .B(new_n3822), .Y(po069));
  xnor_4 g09450(.A(new_n1211), .B(new_n1210), .Y(po070));
  xor_4  g09451(.A(new_n9182), .B(new_n9180), .Y(po071));
  nand_5 g09452(.A(pi141), .B(pi007), .Y(new_n9829));
  or_6   g09453(.A(new_n9829), .B(new_n6386), .Y(new_n9830));
  nand_5 g09454(.A(pi051), .B(pi018), .Y(new_n9831));
  nand_5 g09455(.A(pi108), .B(pi090), .Y(new_n9832));
  xor_4  g09456(.A(new_n9832), .B(new_n9831), .Y(new_n9833));
  xor_4  g09457(.A(new_n9833), .B(new_n6385), .Y(new_n9834));
  not_8  g09458(.A(new_n9834), .Y(new_n9835));
  xor_4  g09459(.A(new_n9829), .B(new_n6386), .Y(new_n9836));
  nand_5 g09460(.A(new_n9836), .B(new_n9835), .Y(new_n9837));
  nand_5 g09461(.A(new_n9837), .B(new_n9830), .Y(new_n9838));
  nand_5 g09462(.A(new_n6406), .B(new_n6405), .Y(new_n9839));
  nand_5 g09463(.A(new_n6407), .B(new_n6404), .Y(new_n9840));
  nand_5 g09464(.A(new_n9840), .B(new_n9839), .Y(new_n9841));
  nand_5 g09465(.A(new_n6403), .B(new_n6399), .Y(new_n9842));
  xor_4  g09466(.A(new_n9836), .B(new_n9834), .Y(new_n9843));
  nand_5 g09467(.A(pi241), .B(pi113), .Y(new_n9844));
  nand_5 g09468(.A(pi236), .B(pi038), .Y(new_n9845));
  xor_4  g09469(.A(new_n9845), .B(new_n9844), .Y(new_n9846));
  xor_4  g09470(.A(new_n9846), .B(new_n6392), .Y(new_n9847));
  nor_5  g09471(.A(new_n6380), .B(new_n6377), .Y(new_n9848));
  nor_5  g09472(.A(new_n6387), .B(new_n6381), .Y(new_n9849));
  nor_5  g09473(.A(new_n9849), .B(new_n9848), .Y(new_n9850));
  xor_4  g09474(.A(new_n9850), .B(new_n9847), .Y(new_n9851));
  xnor_4 g09475(.A(new_n9851), .B(new_n9843), .Y(new_n9852));
  nor_5  g09476(.A(new_n6394), .B(new_n6388), .Y(new_n9853));
  nor_5  g09477(.A(new_n6398), .B(new_n6395), .Y(new_n9854));
  xor_4  g09478(.A(new_n9854), .B(new_n6393), .Y(new_n9855));
  nor_5  g09479(.A(new_n9855), .B(new_n9853), .Y(new_n9856));
  xor_4  g09480(.A(new_n9856), .B(new_n9852), .Y(new_n9857));
  xor_4  g09481(.A(new_n9857), .B(new_n9842), .Y(new_n9858));
  xnor_4 g09482(.A(new_n9858), .B(new_n9841), .Y(new_n9859));
  nand_5 g09483(.A(new_n6435), .B(new_n6432), .Y(new_n9860));
  nand_5 g09484(.A(pi188), .B(pi183), .Y(new_n9861));
  nand_5 g09485(.A(pi112), .B(pi061), .Y(new_n9862));
  xor_4  g09486(.A(new_n9862), .B(new_n9861), .Y(new_n9863));
  xor_4  g09487(.A(new_n9863), .B(new_n6414), .Y(new_n9864));
  nand_5 g09488(.A(pi013), .B(pi012), .Y(new_n9865));
  xor_4  g09489(.A(new_n9865), .B(new_n6415), .Y(new_n9866));
  xor_4  g09490(.A(new_n9866), .B(new_n9864), .Y(new_n9867));
  nand_5 g09491(.A(pi212), .B(pi098), .Y(new_n9868));
  nand_5 g09492(.A(pi213), .B(pi043), .Y(new_n9869));
  xor_4  g09493(.A(new_n9869), .B(new_n9868), .Y(new_n9870));
  xor_4  g09494(.A(new_n9870), .B(new_n6425), .Y(new_n9871));
  nand_5 g09495(.A(new_n6416), .B(new_n6410), .Y(new_n9872));
  nand_5 g09496(.A(new_n6420), .B(new_n6417), .Y(new_n9873));
  nand_5 g09497(.A(new_n9873), .B(new_n9872), .Y(new_n9874));
  xor_4  g09498(.A(new_n9874), .B(new_n9871), .Y(new_n9875));
  xnor_4 g09499(.A(new_n9875), .B(new_n9867), .Y(new_n9876));
  nor_5  g09500(.A(new_n6427), .B(new_n6421), .Y(new_n9877));
  nor_5  g09501(.A(new_n6431), .B(new_n6428), .Y(new_n9878));
  xor_4  g09502(.A(new_n9878), .B(new_n6426), .Y(new_n9879));
  nor_5  g09503(.A(new_n9879), .B(new_n9877), .Y(new_n9880));
  not_8  g09504(.A(new_n9880), .Y(new_n9881));
  xor_4  g09505(.A(new_n9881), .B(new_n9876), .Y(new_n9882));
  xor_4  g09506(.A(new_n9882), .B(new_n9860), .Y(new_n9883));
  nand_5 g09507(.A(new_n6437), .B(new_n6436), .Y(new_n9884));
  nand_5 g09508(.A(new_n6438), .B(new_n6409), .Y(new_n9885));
  nand_5 g09509(.A(new_n9885), .B(new_n9884), .Y(new_n9886));
  xor_4  g09510(.A(new_n9886), .B(new_n9883), .Y(new_n9887));
  xor_4  g09511(.A(new_n9887), .B(new_n9859), .Y(new_n9888));
  not_8  g09512(.A(new_n6439), .Y(new_n9889));
  nor_5  g09513(.A(new_n9889), .B(new_n6408), .Y(new_n9890));
  nor_5  g09514(.A(new_n6444), .B(new_n6440), .Y(new_n9891));
  nor_5  g09515(.A(new_n9891), .B(new_n9890), .Y(new_n9892));
  xor_4  g09516(.A(new_n9892), .B(new_n9888), .Y(new_n9893));
  nand_5 g09517(.A(new_n6472), .B(new_n6468), .Y(new_n9894));
  nand_5 g09518(.A(pi179), .B(pi015), .Y(new_n9895));
  nand_5 g09519(.A(pi162), .B(pi146), .Y(new_n9896));
  xor_4  g09520(.A(new_n9896), .B(new_n9895), .Y(new_n9897));
  xor_4  g09521(.A(new_n9897), .B(new_n6450), .Y(new_n9898));
  not_8  g09522(.A(new_n9898), .Y(new_n9899));
  nand_5 g09523(.A(pi048), .B(pi035), .Y(new_n9900));
  xor_4  g09524(.A(new_n9900), .B(new_n6451), .Y(new_n9901));
  xor_4  g09525(.A(new_n9901), .B(new_n9899), .Y(new_n9902));
  nand_5 g09526(.A(pi193), .B(pi168), .Y(new_n9903));
  nand_5 g09527(.A(pi238), .B(pi208), .Y(new_n9904));
  xor_4  g09528(.A(new_n9904), .B(new_n9903), .Y(new_n9905));
  xor_4  g09529(.A(new_n9905), .B(new_n6461), .Y(new_n9906));
  nand_5 g09530(.A(new_n6452), .B(new_n6446), .Y(new_n9907));
  nand_5 g09531(.A(new_n6456), .B(new_n6453), .Y(new_n9908));
  nand_5 g09532(.A(new_n9908), .B(new_n9907), .Y(new_n9909));
  xor_4  g09533(.A(new_n9909), .B(new_n9906), .Y(new_n9910));
  xor_4  g09534(.A(new_n9910), .B(new_n9902), .Y(new_n9911));
  nor_5  g09535(.A(new_n6467), .B(new_n6464), .Y(new_n9912));
  nand_5 g09536(.A(new_n9912), .B(new_n6462), .Y(new_n9913));
  nor_5  g09537(.A(new_n6463), .B(new_n6457), .Y(new_n9914));
  or_6   g09538(.A(new_n9914), .B(new_n6462), .Y(new_n9915));
  or_6   g09539(.A(new_n9915), .B(new_n9912), .Y(new_n9916));
  nand_5 g09540(.A(new_n9916), .B(new_n9913), .Y(new_n9917));
  xor_4  g09541(.A(new_n9917), .B(new_n9911), .Y(new_n9918));
  xnor_4 g09542(.A(new_n9918), .B(new_n9894), .Y(new_n9919));
  nand_5 g09543(.A(new_n6475), .B(new_n6474), .Y(new_n9920));
  nand_5 g09544(.A(new_n6476), .B(new_n6473), .Y(new_n9921));
  nand_5 g09545(.A(new_n9921), .B(new_n9920), .Y(new_n9922));
  xor_4  g09546(.A(new_n9922), .B(new_n9919), .Y(new_n9923));
  nor_5  g09547(.A(new_n9923), .B(new_n9893), .Y(new_n9924));
  or_6   g09548(.A(new_n6480), .B(new_n6477), .Y(new_n9925));
  nand_5 g09549(.A(new_n6481), .B(new_n6445), .Y(new_n9926));
  nand_5 g09550(.A(new_n9926), .B(new_n9925), .Y(new_n9927));
  xnor_4 g09551(.A(new_n9923), .B(new_n9893), .Y(new_n9928));
  nor_5  g09552(.A(new_n9928), .B(new_n9927), .Y(new_n9929));
  nor_5  g09553(.A(new_n9929), .B(new_n9924), .Y(new_n9930));
  nand_5 g09554(.A(pi194), .B(pi064), .Y(new_n9931));
  nand_5 g09555(.A(pi068), .B(pi052), .Y(new_n9932));
  nand_5 g09556(.A(pi077), .B(pi036), .Y(new_n9933));
  xor_4  g09557(.A(new_n9933), .B(new_n9932), .Y(new_n9934));
  xor_4  g09558(.A(new_n9934), .B(new_n9931), .Y(new_n9935));
  xor_4  g09559(.A(new_n9935), .B(new_n9930), .Y(new_n9936));
  nand_5 g09560(.A(pi131), .B(pi068), .Y(new_n9937));
  nand_5 g09561(.A(pi052), .B(pi036), .Y(new_n9938));
  nand_5 g09562(.A(new_n9938), .B(new_n9937), .Y(new_n9939));
  xor_4  g09563(.A(new_n9938), .B(new_n9937), .Y(new_n9940));
  nand_5 g09564(.A(new_n9940), .B(new_n6498), .Y(new_n9941));
  nand_5 g09565(.A(new_n9941), .B(new_n9939), .Y(new_n9942));
  xor_4  g09566(.A(new_n9940), .B(new_n6498), .Y(new_n9943));
  nand_5 g09567(.A(new_n6489), .B(new_n6483), .Y(new_n9944));
  nand_5 g09568(.A(new_n6493), .B(new_n6490), .Y(new_n9945));
  nand_5 g09569(.A(new_n9945), .B(new_n9944), .Y(new_n9946));
  or_6   g09570(.A(new_n9946), .B(new_n9943), .Y(new_n9947));
  nand_5 g09571(.A(pi194), .B(pi189), .Y(new_n9948));
  nand_5 g09572(.A(pi143), .B(pi084), .Y(new_n9949));
  xor_4  g09573(.A(new_n9949), .B(new_n9948), .Y(new_n9950));
  xor_4  g09574(.A(new_n9950), .B(new_n6487), .Y(new_n9951));
  not_8  g09575(.A(new_n9951), .Y(new_n9952));
  nand_5 g09576(.A(pi133), .B(pi085), .Y(new_n9953));
  xor_4  g09577(.A(new_n9953), .B(new_n6488), .Y(new_n9954));
  xor_4  g09578(.A(new_n9954), .B(new_n9952), .Y(new_n9955));
  xor_4  g09579(.A(new_n9946), .B(new_n9943), .Y(new_n9956));
  nand_5 g09580(.A(new_n9956), .B(new_n9955), .Y(new_n9957));
  nand_5 g09581(.A(new_n9957), .B(new_n9947), .Y(new_n9958));
  xor_4  g09582(.A(new_n9958), .B(new_n9942), .Y(new_n9959));
  nand_5 g09583(.A(pi189), .B(pi085), .Y(new_n9960));
  nand_5 g09584(.A(pi180), .B(pi133), .Y(new_n9961));
  xor_4  g09585(.A(new_n9961), .B(new_n9960), .Y(new_n9962));
  xor_4  g09586(.A(new_n9962), .B(new_n9959), .Y(new_n9963));
  nor_5  g09587(.A(new_n9918), .B(new_n9894), .Y(new_n9964));
  nor_5  g09588(.A(new_n9922), .B(new_n9919), .Y(new_n9965));
  nor_5  g09589(.A(new_n9965), .B(new_n9964), .Y(new_n9966));
  nand_5 g09590(.A(pi084), .B(pi057), .Y(new_n9967));
  xor_4  g09591(.A(new_n9967), .B(new_n9966), .Y(new_n9968));
  xor_4  g09592(.A(new_n9968), .B(new_n9963), .Y(new_n9969));
  nand_5 g09593(.A(pi168), .B(pi159), .Y(new_n9970));
  nand_5 g09594(.A(pi146), .B(pi033), .Y(new_n9971));
  nand_5 g09595(.A(pi162), .B(pi152), .Y(new_n9972));
  or_6   g09596(.A(new_n9917), .B(new_n9911), .Y(new_n9973));
  nand_5 g09597(.A(new_n9973), .B(new_n9916), .Y(new_n9974));
  xor_4  g09598(.A(new_n9974), .B(new_n9972), .Y(new_n9975));
  xor_4  g09599(.A(new_n9975), .B(new_n9971), .Y(new_n9976));
  xor_4  g09600(.A(new_n9976), .B(new_n9970), .Y(new_n9977));
  nand_5 g09601(.A(new_n9949), .B(new_n9948), .Y(new_n9978));
  nand_5 g09602(.A(new_n9950), .B(new_n6487), .Y(new_n9979));
  nand_5 g09603(.A(new_n9979), .B(new_n9978), .Y(new_n9980));
  or_6   g09604(.A(new_n9953), .B(new_n6488), .Y(new_n9981));
  nand_5 g09605(.A(new_n9954), .B(new_n9952), .Y(new_n9982));
  nand_5 g09606(.A(new_n9982), .B(new_n9981), .Y(new_n9983));
  xor_4  g09607(.A(new_n9983), .B(new_n9980), .Y(new_n9984));
  xor_4  g09608(.A(new_n9984), .B(new_n9977), .Y(new_n9985));
  xor_4  g09609(.A(new_n9985), .B(new_n9969), .Y(new_n9986));
  xor_4  g09610(.A(new_n9986), .B(new_n9936), .Y(new_n9987));
  nand_5 g09611(.A(pi144), .B(pi013), .Y(new_n9988));
  nand_5 g09612(.A(new_n9874), .B(new_n9871), .Y(new_n9989));
  nand_5 g09613(.A(new_n9875), .B(new_n9867), .Y(new_n9990));
  nand_5 g09614(.A(new_n9990), .B(new_n9989), .Y(new_n9991));
  xor_4  g09615(.A(new_n9991), .B(new_n9988), .Y(new_n9992));
  nand_5 g09616(.A(pi112), .B(pi012), .Y(new_n9993));
  xor_4  g09617(.A(new_n9993), .B(new_n9992), .Y(new_n9994));
  xor_4  g09618(.A(new_n9994), .B(new_n9987), .Y(new_n9995));
  or_6   g09619(.A(new_n9900), .B(new_n6451), .Y(new_n9996));
  nand_5 g09620(.A(new_n9901), .B(new_n9899), .Y(new_n9997));
  nand_5 g09621(.A(new_n9997), .B(new_n9996), .Y(new_n9998));
  nand_5 g09622(.A(pi237), .B(pi035), .Y(new_n9999));
  nand_5 g09623(.A(pi238), .B(pi139), .Y(new_n10000));
  xor_4  g09624(.A(new_n10000), .B(new_n9999), .Y(new_n10001));
  xor_4  g09625(.A(new_n10001), .B(new_n9998), .Y(new_n10002));
  nand_5 g09626(.A(new_n9878), .B(new_n6426), .Y(new_n10003));
  nand_5 g09627(.A(new_n9881), .B(new_n9876), .Y(new_n10004));
  nand_5 g09628(.A(new_n10004), .B(new_n10003), .Y(new_n10005));
  nand_5 g09629(.A(pi204), .B(pi179), .Y(new_n10006));
  xor_4  g09630(.A(new_n10006), .B(new_n10005), .Y(new_n10007));
  xor_4  g09631(.A(new_n10007), .B(new_n10002), .Y(new_n10008));
  or_6   g09632(.A(new_n9909), .B(new_n9906), .Y(new_n10009));
  nand_5 g09633(.A(new_n9910), .B(new_n9902), .Y(new_n10010));
  nand_5 g09634(.A(new_n10010), .B(new_n10009), .Y(new_n10011));
  nand_5 g09635(.A(new_n9896), .B(new_n9895), .Y(new_n10012));
  nand_5 g09636(.A(new_n9897), .B(new_n6450), .Y(new_n10013));
  nand_5 g09637(.A(new_n10013), .B(new_n10012), .Y(new_n10014));
  xor_4  g09638(.A(new_n10014), .B(new_n10011), .Y(new_n10015));
  xor_4  g09639(.A(new_n10015), .B(new_n10008), .Y(new_n10016));
  nand_5 g09640(.A(new_n9862), .B(new_n9861), .Y(new_n10017));
  nand_5 g09641(.A(new_n9863), .B(new_n6414), .Y(new_n10018));
  nand_5 g09642(.A(new_n10018), .B(new_n10017), .Y(new_n10019));
  or_6   g09643(.A(new_n9865), .B(new_n6415), .Y(new_n10020));
  not_8  g09644(.A(new_n9864), .Y(new_n10021));
  nand_5 g09645(.A(new_n9866), .B(new_n10021), .Y(new_n10022));
  nand_5 g09646(.A(new_n10022), .B(new_n10020), .Y(new_n10023));
  xor_4  g09647(.A(new_n10023), .B(new_n10019), .Y(new_n10024));
  nand_5 g09648(.A(new_n9887), .B(new_n9859), .Y(new_n10025));
  nand_5 g09649(.A(new_n9892), .B(new_n9888), .Y(new_n10026));
  nand_5 g09650(.A(new_n10026), .B(new_n10025), .Y(new_n10027));
  nand_5 g09651(.A(pi213), .B(pi126), .Y(new_n10028));
  xor_4  g09652(.A(new_n10028), .B(new_n10027), .Y(new_n10029));
  nand_5 g09653(.A(new_n9904), .B(new_n9903), .Y(new_n10030));
  nand_5 g09654(.A(new_n9905), .B(new_n6461), .Y(new_n10031));
  nand_5 g09655(.A(new_n10031), .B(new_n10030), .Y(new_n10032));
  nand_5 g09656(.A(pi188), .B(pi088), .Y(new_n10033));
  not_8  g09657(.A(new_n9882), .Y(new_n10034));
  nor_5  g09658(.A(new_n10034), .B(new_n9860), .Y(new_n10035));
  nor_5  g09659(.A(new_n9886), .B(new_n9883), .Y(new_n10036));
  or_6   g09660(.A(new_n10036), .B(new_n10035), .Y(new_n10037));
  nand_5 g09661(.A(pi183), .B(pi178), .Y(new_n10038));
  nand_5 g09662(.A(pi105), .B(pi061), .Y(new_n10039));
  xor_4  g09663(.A(new_n10039), .B(new_n10038), .Y(new_n10040));
  xor_4  g09664(.A(new_n10040), .B(new_n10037), .Y(new_n10041));
  xor_4  g09665(.A(new_n10041), .B(new_n10033), .Y(new_n10042));
  xor_4  g09666(.A(new_n10042), .B(new_n10032), .Y(new_n10043));
  xor_4  g09667(.A(new_n10043), .B(new_n10029), .Y(new_n10044));
  nand_5 g09668(.A(pi208), .B(pi193), .Y(new_n10045));
  nand_5 g09669(.A(pi048), .B(pi015), .Y(new_n10046));
  xor_4  g09670(.A(new_n10046), .B(new_n10045), .Y(new_n10047));
  xor_4  g09671(.A(new_n10047), .B(new_n10044), .Y(new_n10048));
  xor_4  g09672(.A(new_n10048), .B(new_n10024), .Y(new_n10049));
  xor_4  g09673(.A(new_n10049), .B(new_n10016), .Y(new_n10050));
  nand_5 g09674(.A(new_n9869), .B(new_n9868), .Y(new_n10051));
  nand_5 g09675(.A(new_n9870), .B(new_n6425), .Y(new_n10052));
  nand_5 g09676(.A(new_n10052), .B(new_n10051), .Y(new_n10053));
  nand_5 g09677(.A(new_n9857), .B(new_n9842), .Y(new_n10054));
  nand_5 g09678(.A(new_n9858), .B(new_n9841), .Y(new_n10055));
  nand_5 g09679(.A(new_n10055), .B(new_n10054), .Y(new_n10056));
  xor_4  g09680(.A(new_n10056), .B(new_n10053), .Y(new_n10057));
  nand_5 g09681(.A(pi212), .B(pi043), .Y(new_n10058));
  nand_5 g09682(.A(pi104), .B(pi098), .Y(new_n10059));
  xor_4  g09683(.A(new_n10059), .B(new_n10058), .Y(new_n10060));
  nand_5 g09684(.A(new_n9854), .B(new_n6393), .Y(new_n10061));
  not_8  g09685(.A(new_n9856), .Y(new_n10062));
  nand_5 g09686(.A(new_n10062), .B(new_n9852), .Y(new_n10063));
  nand_5 g09687(.A(new_n10063), .B(new_n10061), .Y(new_n10064));
  nand_5 g09688(.A(pi090), .B(pi007), .Y(new_n10065));
  nand_5 g09689(.A(pi141), .B(pi118), .Y(new_n10066));
  xor_4  g09690(.A(new_n10066), .B(new_n10065), .Y(new_n10067));
  xor_4  g09691(.A(new_n10067), .B(new_n10064), .Y(new_n10068));
  nand_5 g09692(.A(pi108), .B(pi047), .Y(new_n10069));
  nand_5 g09693(.A(pi236), .B(pi028), .Y(new_n10070));
  nand_5 g09694(.A(pi042), .B(pi018), .Y(new_n10071));
  nand_5 g09695(.A(pi128), .B(pi051), .Y(new_n10072));
  xnor_4 g09696(.A(new_n10072), .B(new_n10071), .Y(new_n10073));
  xor_4  g09697(.A(new_n10073), .B(new_n10070), .Y(new_n10074));
  xor_4  g09698(.A(new_n10074), .B(new_n10069), .Y(new_n10075));
  xor_4  g09699(.A(new_n10075), .B(new_n10068), .Y(new_n10076));
  xor_4  g09700(.A(new_n10076), .B(new_n10060), .Y(new_n10077));
  xor_4  g09701(.A(new_n10077), .B(new_n10057), .Y(new_n10078));
  xor_4  g09702(.A(new_n10078), .B(new_n10050), .Y(new_n10079));
  xor_4  g09703(.A(new_n10079), .B(new_n9995), .Y(new_n10080));
  xor_4  g09704(.A(new_n10080), .B(new_n9838), .Y(new_n10081));
  nand_5 g09705(.A(new_n9832), .B(new_n9831), .Y(new_n10082));
  nand_5 g09706(.A(new_n9833), .B(new_n6385), .Y(new_n10083));
  nand_5 g09707(.A(new_n10083), .B(new_n10082), .Y(new_n10084));
  xor_4  g09708(.A(new_n9928), .B(new_n9927), .Y(new_n10085));
  nand_5 g09709(.A(new_n6509), .B(new_n6506), .Y(new_n10086));
  xor_4  g09710(.A(new_n9956), .B(new_n9955), .Y(new_n10087));
  nor_5  g09711(.A(new_n6505), .B(new_n6502), .Y(new_n10088));
  and_6  g09712(.A(new_n10088), .B(new_n6499), .Y(new_n10089));
  or_6   g09713(.A(new_n6501), .B(new_n6494), .Y(new_n10090));
  nand_5 g09714(.A(new_n10090), .B(new_n6500), .Y(new_n10091));
  nor_5  g09715(.A(new_n10091), .B(new_n10088), .Y(new_n10092));
  or_6   g09716(.A(new_n10092), .B(new_n10089), .Y(new_n10093));
  xor_4  g09717(.A(new_n10093), .B(new_n10087), .Y(new_n10094));
  xnor_4 g09718(.A(new_n10094), .B(new_n10086), .Y(new_n10095));
  nand_5 g09719(.A(new_n6512), .B(new_n6511), .Y(new_n10096));
  nand_5 g09720(.A(new_n6513), .B(new_n6510), .Y(new_n10097));
  nand_5 g09721(.A(new_n10097), .B(new_n10096), .Y(new_n10098));
  xor_4  g09722(.A(new_n10098), .B(new_n10095), .Y(new_n10099));
  not_8  g09723(.A(new_n10099), .Y(new_n10100));
  nor_5  g09724(.A(new_n10100), .B(new_n10085), .Y(new_n10101));
  xor_4  g09725(.A(new_n10099), .B(new_n10085), .Y(new_n10102));
  nand_5 g09726(.A(new_n6518), .B(new_n6514), .Y(new_n10103));
  not_8  g09727(.A(new_n6482), .Y(new_n10104));
  nand_5 g09728(.A(new_n6519), .B(new_n10104), .Y(new_n10105));
  nand_5 g09729(.A(new_n10105), .B(new_n10103), .Y(new_n10106));
  nor_5  g09730(.A(new_n10106), .B(new_n10102), .Y(new_n10107));
  nor_5  g09731(.A(new_n10107), .B(new_n10101), .Y(new_n10108));
  nand_5 g09732(.A(new_n9850), .B(new_n9847), .Y(new_n10109));
  nand_5 g09733(.A(new_n9851), .B(new_n9843), .Y(new_n10110));
  nand_5 g09734(.A(new_n10110), .B(new_n10109), .Y(new_n10111));
  nand_5 g09735(.A(new_n9845), .B(new_n9844), .Y(new_n10112));
  nand_5 g09736(.A(new_n9846), .B(new_n6392), .Y(new_n10113));
  nand_5 g09737(.A(new_n10113), .B(new_n10112), .Y(new_n10114));
  xor_4  g09738(.A(new_n10114), .B(new_n10111), .Y(new_n10115));
  xor_4  g09739(.A(new_n10115), .B(new_n10108), .Y(new_n10116));
  xor_4  g09740(.A(new_n10116), .B(new_n10084), .Y(new_n10117));
  nand_5 g09741(.A(pi241), .B(pi038), .Y(new_n10118));
  nand_5 g09742(.A(pi161), .B(pi113), .Y(new_n10119));
  xor_4  g09743(.A(new_n10119), .B(new_n10118), .Y(new_n10120));
  nand_5 g09744(.A(pi143), .B(pi034), .Y(new_n10121));
  nand_5 g09745(.A(pi131), .B(pi046), .Y(new_n10122));
  xor_4  g09746(.A(new_n10122), .B(new_n10121), .Y(new_n10123));
  nor_5  g09747(.A(new_n10093), .B(new_n10087), .Y(new_n10124));
  nor_5  g09748(.A(new_n10124), .B(new_n10092), .Y(new_n10125));
  nor_5  g09749(.A(new_n10094), .B(new_n10086), .Y(new_n10126));
  nor_5  g09750(.A(new_n10098), .B(new_n10095), .Y(new_n10127));
  nor_5  g09751(.A(new_n10127), .B(new_n10126), .Y(new_n10128));
  xor_4  g09752(.A(new_n10128), .B(new_n10125), .Y(new_n10129));
  xor_4  g09753(.A(new_n10129), .B(new_n10123), .Y(new_n10130));
  xor_4  g09754(.A(new_n10130), .B(new_n10120), .Y(new_n10131));
  xor_4  g09755(.A(new_n10131), .B(new_n10117), .Y(new_n10132));
  xor_4  g09756(.A(new_n10132), .B(new_n10081), .Y(po072));
  xor_4  g09757(.A(new_n895), .B(new_n894), .Y(po073));
  xor_4  g09758(.A(new_n6202), .B(new_n6198), .Y(po074));
  xor_4  g09759(.A(new_n7532), .B(new_n7511), .Y(po075));
  xor_4  g09760(.A(new_n6602), .B(new_n6601), .Y(po076));
  xor_4  g09761(.A(new_n1196), .B(new_n1190), .Y(po077));
  xor_4  g09762(.A(new_n1832), .B(new_n1831), .Y(po078));
  xor_4  g09763(.A(new_n5675), .B(new_n5673), .Y(po079));
  xnor_4 g09764(.A(new_n9170), .B(new_n9169), .Y(po080));
  xor_4  g09765(.A(new_n7528), .B(new_n7526), .Y(po081));
  xor_4  g09766(.A(new_n6204), .B(new_n6192), .Y(po082));
  xor_4  g09767(.A(new_n1204), .B(new_n1202), .Y(po083));
  not_8  g09768(.A(new_n722), .Y(new_n10145));
  nand_5 g09769(.A(new_n10145), .B(new_n622), .Y(new_n10146));
  or_6   g09770(.A(new_n760), .B(new_n723), .Y(new_n10147));
  nand_5 g09771(.A(new_n10147), .B(new_n10146), .Y(new_n10148));
  nand_5 g09772(.A(pi167), .B(pi097), .Y(new_n10149));
  nand_5 g09773(.A(pi166), .B(pi134), .Y(new_n10150));
  nand_5 g09774(.A(new_n683), .B(new_n682), .Y(new_n10151));
  nand_5 g09775(.A(new_n684), .B(new_n628), .Y(new_n10152));
  nand_5 g09776(.A(new_n10152), .B(new_n10151), .Y(new_n10153));
  xor_4  g09777(.A(new_n10153), .B(new_n10150), .Y(new_n10154));
  xor_4  g09778(.A(new_n10154), .B(new_n10149), .Y(new_n10155));
  xor_4  g09779(.A(new_n10155), .B(new_n10148), .Y(new_n10156));
  nand_5 g09780(.A(new_n690), .B(new_n689), .Y(new_n10157));
  nand_5 g09781(.A(new_n691), .B(new_n643), .Y(new_n10158));
  nand_5 g09782(.A(new_n10158), .B(new_n10157), .Y(new_n10159));
  nand_5 g09783(.A(pi149), .B(pi075), .Y(new_n10160));
  nand_5 g09784(.A(pi240), .B(pi093), .Y(new_n10161));
  xor_4  g09785(.A(new_n10161), .B(new_n10160), .Y(new_n10162));
  xor_4  g09786(.A(new_n10162), .B(new_n10159), .Y(new_n10163));
  nand_5 g09787(.A(pi181), .B(pi019), .Y(new_n10164));
  nand_5 g09788(.A(pi164), .B(pi000), .Y(new_n10165));
  nand_5 g09789(.A(pi206), .B(pi115), .Y(new_n10166));
  nand_5 g09790(.A(pi070), .B(pi032), .Y(new_n10167));
  xor_4  g09791(.A(new_n10167), .B(new_n10166), .Y(new_n10168));
  nand_5 g09792(.A(pi163), .B(pi031), .Y(new_n10169));
  nand_5 g09793(.A(new_n580), .B(new_n483), .Y(new_n10170));
  not_8  g09794(.A(new_n621), .Y(new_n10171));
  nand_5 g09795(.A(new_n10171), .B(new_n581), .Y(new_n10172));
  nand_5 g09796(.A(new_n10172), .B(new_n10170), .Y(new_n10173));
  xor_4  g09797(.A(new_n10173), .B(new_n10169), .Y(new_n10174));
  xor_4  g09798(.A(new_n10174), .B(new_n10168), .Y(new_n10175));
  xor_4  g09799(.A(new_n10175), .B(new_n10165), .Y(new_n10176));
  xor_4  g09800(.A(new_n10176), .B(new_n10164), .Y(new_n10177));
  xor_4  g09801(.A(new_n10177), .B(new_n10163), .Y(new_n10178));
  nand_5 g09802(.A(new_n558), .B(new_n505), .Y(new_n10179));
  nand_5 g09803(.A(new_n561), .B(new_n556), .Y(new_n10180));
  nand_5 g09804(.A(new_n10180), .B(new_n10179), .Y(new_n10181));
  not_8  g09805(.A(new_n562), .Y(new_n10182));
  nor_5  g09806(.A(new_n10182), .B(new_n540), .Y(new_n10183));
  nor_5  g09807(.A(new_n579), .B(new_n563), .Y(new_n10184));
  nor_5  g09808(.A(new_n10184), .B(new_n10183), .Y(new_n10185));
  xor_4  g09809(.A(new_n10185), .B(new_n10181), .Y(new_n10186));
  or_6   g09810(.A(new_n686), .B(new_n629), .Y(new_n10187));
  not_8  g09811(.A(new_n685), .Y(new_n10188));
  nand_5 g09812(.A(new_n687), .B(new_n10188), .Y(new_n10189));
  nand_5 g09813(.A(new_n10189), .B(new_n10187), .Y(new_n10190));
  nand_5 g09814(.A(new_n695), .B(new_n692), .Y(new_n10191));
  nand_5 g09815(.A(new_n696), .B(new_n688), .Y(new_n10192));
  nand_5 g09816(.A(new_n10192), .B(new_n10191), .Y(new_n10193));
  xor_4  g09817(.A(new_n10193), .B(new_n10190), .Y(new_n10194));
  xor_4  g09818(.A(new_n10194), .B(new_n10186), .Y(new_n10195));
  xor_4  g09819(.A(new_n10195), .B(new_n10178), .Y(new_n10196));
  xor_4  g09820(.A(new_n10196), .B(new_n10156), .Y(new_n10197));
  nand_5 g09821(.A(pi250), .B(pi234), .Y(new_n10198));
  nand_5 g09822(.A(new_n821), .B(new_n820), .Y(new_n10199));
  nand_5 g09823(.A(new_n822), .B(new_n774), .Y(new_n10200));
  nand_5 g09824(.A(new_n10200), .B(new_n10199), .Y(new_n10201));
  xor_4  g09825(.A(new_n10201), .B(new_n10198), .Y(new_n10202));
  xor_4  g09826(.A(new_n10202), .B(new_n10197), .Y(new_n10203));
  nand_5 g09827(.A(new_n829), .B(new_n783), .Y(new_n10204));
  nand_5 g09828(.A(new_n830), .B(new_n828), .Y(new_n10205));
  nand_5 g09829(.A(new_n10205), .B(new_n10204), .Y(new_n10206));
  nand_5 g09830(.A(pi247), .B(pi044), .Y(new_n10207));
  nand_5 g09831(.A(pi080), .B(pi054), .Y(new_n10208));
  xor_4  g09832(.A(new_n10208), .B(new_n10207), .Y(new_n10209));
  xor_4  g09833(.A(new_n10209), .B(new_n10206), .Y(new_n10210));
  or_6   g09834(.A(new_n702), .B(new_n681), .Y(new_n10211));
  nand_5 g09835(.A(new_n721), .B(new_n703), .Y(new_n10212));
  nand_5 g09836(.A(new_n10212), .B(new_n10211), .Y(new_n10213));
  nand_5 g09837(.A(pi214), .B(pi045), .Y(new_n10214));
  xor_4  g09838(.A(new_n10214), .B(new_n10213), .Y(new_n10215));
  xor_4  g09839(.A(new_n10215), .B(new_n10210), .Y(new_n10216));
  nand_5 g09840(.A(pi200), .B(pi151), .Y(new_n10217));
  nand_5 g09841(.A(pi203), .B(pi147), .Y(new_n10218));
  nand_5 g09842(.A(new_n699), .B(new_n644), .Y(new_n10219));
  not_8  g09843(.A(new_n701), .Y(new_n10220));
  nand_5 g09844(.A(new_n10220), .B(new_n697), .Y(new_n10221));
  nand_5 g09845(.A(new_n10221), .B(new_n10219), .Y(new_n10222));
  xor_4  g09846(.A(new_n10222), .B(new_n10218), .Y(new_n10223));
  xor_4  g09847(.A(new_n10223), .B(new_n10217), .Y(new_n10224));
  nand_5 g09848(.A(pi175), .B(pi011), .Y(new_n10225));
  or_6   g09849(.A(new_n834), .B(new_n831), .Y(new_n10226));
  nand_5 g09850(.A(new_n835), .B(new_n827), .Y(new_n10227));
  nand_5 g09851(.A(new_n10227), .B(new_n10226), .Y(new_n10228));
  xor_4  g09852(.A(new_n10228), .B(new_n10225), .Y(new_n10229));
  xor_4  g09853(.A(new_n10229), .B(new_n10224), .Y(new_n10230));
  nand_5 g09854(.A(pi072), .B(pi016), .Y(new_n10231));
  nand_5 g09855(.A(pi248), .B(pi117), .Y(new_n10232));
  nor_5  g09856(.A(new_n824), .B(new_n776), .Y(new_n10233));
  nor_5  g09857(.A(new_n826), .B(new_n823), .Y(new_n10234));
  or_6   g09858(.A(new_n10234), .B(new_n10233), .Y(new_n10235));
  xor_4  g09859(.A(new_n10235), .B(new_n10232), .Y(new_n10236));
  xor_4  g09860(.A(new_n10236), .B(new_n10231), .Y(new_n10237));
  xor_4  g09861(.A(new_n10237), .B(new_n10230), .Y(new_n10238));
  xor_4  g09862(.A(new_n10238), .B(new_n10216), .Y(new_n10239));
  xor_4  g09863(.A(new_n10239), .B(new_n10203), .Y(new_n10240));
  or_6   g09864(.A(new_n842), .B(new_n836), .Y(new_n10241));
  nand_5 g09865(.A(new_n10241), .B(new_n841), .Y(new_n10242));
  nand_5 g09866(.A(new_n444), .B(new_n443), .Y(new_n10243));
  nand_5 g09867(.A(new_n445), .B(new_n389), .Y(new_n10244));
  nand_5 g09868(.A(new_n10244), .B(new_n10243), .Y(new_n10245));
  xor_4  g09869(.A(new_n10245), .B(new_n10242), .Y(new_n10246));
  xor_4  g09870(.A(new_n10246), .B(new_n10240), .Y(new_n10247));
  nor_5  g09871(.A(new_n843), .B(new_n819), .Y(new_n10248));
  nor_5  g09872(.A(new_n861), .B(new_n844), .Y(new_n10249));
  nor_5  g09873(.A(new_n10249), .B(new_n10248), .Y(new_n10250));
  nand_5 g09874(.A(new_n452), .B(new_n451), .Y(new_n10251));
  nand_5 g09875(.A(new_n453), .B(new_n416), .Y(new_n10252));
  nand_5 g09876(.A(new_n10252), .B(new_n10251), .Y(new_n10253));
  nand_5 g09877(.A(pi096), .B(pi049), .Y(new_n10254));
  xor_4  g09878(.A(new_n10254), .B(new_n10253), .Y(new_n10255));
  xor_4  g09879(.A(new_n10255), .B(new_n10250), .Y(new_n10256));
  nand_5 g09880(.A(new_n863), .B(new_n761), .Y(new_n10257));
  nand_5 g09881(.A(new_n903), .B(new_n864), .Y(new_n10258));
  nand_5 g09882(.A(new_n10258), .B(new_n10257), .Y(new_n10259));
  nand_5 g09883(.A(pi202), .B(pi119), .Y(new_n10260));
  nand_5 g09884(.A(pi103), .B(pi009), .Y(new_n10261));
  xor_4  g09885(.A(new_n10261), .B(new_n10260), .Y(new_n10262));
  or_6   g09886(.A(new_n448), .B(new_n390), .Y(new_n10263));
  nand_5 g09887(.A(new_n449), .B(new_n447), .Y(new_n10264));
  nand_5 g09888(.A(new_n10264), .B(new_n10263), .Y(new_n10265));
  xor_4  g09889(.A(new_n10265), .B(new_n10262), .Y(new_n10266));
  xor_4  g09890(.A(new_n10266), .B(new_n10259), .Y(new_n10267));
  xor_4  g09891(.A(new_n10267), .B(new_n10256), .Y(new_n10268));
  nor_5  g09892(.A(new_n464), .B(new_n442), .Y(new_n10269));
  nor_5  g09893(.A(new_n482), .B(new_n465), .Y(new_n10270));
  nor_5  g09894(.A(new_n10270), .B(new_n10269), .Y(new_n10271));
  nand_5 g09895(.A(pi201), .B(pi056), .Y(new_n10272));
  nand_5 g09896(.A(pi245), .B(pi136), .Y(new_n10273));
  xor_4  g09897(.A(new_n10273), .B(new_n10272), .Y(new_n10274));
  xor_4  g09898(.A(new_n10274), .B(new_n10271), .Y(new_n10275));
  nand_5 g09899(.A(pi110), .B(pi107), .Y(new_n10276));
  nand_5 g09900(.A(pi083), .B(pi027), .Y(new_n10277));
  nand_5 g09901(.A(pi063), .B(pi026), .Y(new_n10278));
  nand_5 g09902(.A(pi156), .B(pi008), .Y(new_n10279));
  xor_4  g09903(.A(new_n10279), .B(new_n10278), .Y(new_n10280));
  nand_5 g09904(.A(new_n542), .B(new_n541), .Y(new_n10281));
  nand_5 g09905(.A(new_n543), .B(new_n489), .Y(new_n10282));
  nand_5 g09906(.A(new_n10282), .B(new_n10281), .Y(new_n10283));
  nand_5 g09907(.A(new_n549), .B(new_n548), .Y(new_n10284));
  nand_5 g09908(.A(new_n550), .B(new_n504), .Y(new_n10285));
  nand_5 g09909(.A(new_n10285), .B(new_n10284), .Y(new_n10286));
  xor_4  g09910(.A(new_n10286), .B(new_n10283), .Y(new_n10287));
  nand_5 g09911(.A(pi145), .B(pi116), .Y(new_n10288));
  xor_4  g09912(.A(new_n10288), .B(new_n10287), .Y(new_n10289));
  or_6   g09913(.A(new_n545), .B(new_n490), .Y(new_n10290));
  not_8  g09914(.A(new_n544), .Y(new_n10291));
  nand_5 g09915(.A(new_n546), .B(new_n10291), .Y(new_n10292));
  nand_5 g09916(.A(new_n10292), .B(new_n10290), .Y(new_n10293));
  or_6   g09917(.A(new_n462), .B(new_n417), .Y(new_n10294));
  nand_5 g09918(.A(new_n463), .B(new_n459), .Y(new_n10295));
  nand_5 g09919(.A(new_n10295), .B(new_n10294), .Y(new_n10296));
  xor_4  g09920(.A(new_n10296), .B(new_n10293), .Y(new_n10297));
  nand_5 g09921(.A(pi148), .B(pi091), .Y(new_n10298));
  nand_5 g09922(.A(pi228), .B(pi114), .Y(new_n10299));
  xor_4  g09923(.A(new_n10299), .B(new_n10298), .Y(new_n10300));
  nand_5 g09924(.A(pi246), .B(pi039), .Y(new_n10301));
  nand_5 g09925(.A(new_n554), .B(new_n551), .Y(new_n10302));
  nand_5 g09926(.A(new_n555), .B(new_n547), .Y(new_n10303));
  nand_5 g09927(.A(new_n10303), .B(new_n10302), .Y(new_n10304));
  xnor_4 g09928(.A(new_n10304), .B(new_n10301), .Y(new_n10305));
  xor_4  g09929(.A(new_n10305), .B(new_n10300), .Y(new_n10306));
  xor_4  g09930(.A(new_n10306), .B(new_n10297), .Y(new_n10307));
  xor_4  g09931(.A(new_n10307), .B(new_n10289), .Y(new_n10308));
  xor_4  g09932(.A(new_n10308), .B(new_n10280), .Y(new_n10309));
  xor_4  g09933(.A(new_n10309), .B(new_n10277), .Y(new_n10310));
  xor_4  g09934(.A(new_n10310), .B(new_n10276), .Y(new_n10311));
  xor_4  g09935(.A(new_n10311), .B(new_n10275), .Y(new_n10312));
  nand_5 g09936(.A(pi235), .B(pi171), .Y(new_n10313));
  nand_5 g09937(.A(new_n457), .B(new_n454), .Y(new_n10314));
  not_8  g09938(.A(new_n450), .Y(new_n10315));
  nand_5 g09939(.A(new_n458), .B(new_n10315), .Y(new_n10316));
  nand_5 g09940(.A(new_n10316), .B(new_n10314), .Y(new_n10317));
  xor_4  g09941(.A(new_n10317), .B(new_n10313), .Y(new_n10318));
  xor_4  g09942(.A(new_n10318), .B(new_n10312), .Y(new_n10319));
  xor_4  g09943(.A(new_n10319), .B(new_n10268), .Y(new_n10320));
  xor_4  g09944(.A(new_n10320), .B(new_n10247), .Y(po084));
  xor_4  g09945(.A(new_n10106), .B(new_n10102), .Y(po085));
  nand_5 g09946(.A(new_n9612), .B(new_n9611), .Y(new_n10323));
  nand_5 g09947(.A(new_n9613), .B(new_n9516), .Y(new_n10324));
  nand_5 g09948(.A(new_n10324), .B(new_n10323), .Y(new_n10325));
  or_6   g09949(.A(new_n9608), .B(new_n9506), .Y(new_n10326));
  nand_5 g09950(.A(new_n9609), .B(new_n9607), .Y(new_n10327));
  nand_5 g09951(.A(new_n10327), .B(new_n10326), .Y(new_n10328));
  xor_4  g09952(.A(new_n10328), .B(new_n10325), .Y(new_n10329));
  nor_5  g09953(.A(new_n9430), .B(new_n9423), .Y(new_n10330));
  nor_5  g09954(.A(new_n9431), .B(new_n9402), .Y(new_n10331));
  nor_5  g09955(.A(new_n10331), .B(new_n10330), .Y(new_n10332));
  nand_5 g09956(.A(pi210), .B(pi088), .Y(new_n10333));
  nand_5 g09957(.A(pi183), .B(pi111), .Y(new_n10334));
  nand_5 g09958(.A(pi105), .B(pi024), .Y(new_n10335));
  xor_4  g09959(.A(new_n10335), .B(new_n10334), .Y(new_n10336));
  nand_5 g09960(.A(pi213), .B(pi191), .Y(new_n10337));
  nand_5 g09961(.A(new_n9633), .B(new_n9601), .Y(new_n10338));
  nand_5 g09962(.A(new_n9637), .B(new_n9634), .Y(new_n10339));
  nand_5 g09963(.A(new_n10339), .B(new_n10338), .Y(new_n10340));
  xor_4  g09964(.A(new_n10340), .B(new_n10337), .Y(new_n10341));
  xor_4  g09965(.A(new_n10341), .B(new_n10336), .Y(new_n10342));
  xor_4  g09966(.A(new_n10342), .B(new_n10333), .Y(new_n10343));
  nand_5 g09967(.A(new_n9415), .B(new_n9414), .Y(new_n10344));
  nand_5 g09968(.A(new_n9416), .B(new_n9393), .Y(new_n10345));
  nand_5 g09969(.A(new_n10345), .B(new_n10344), .Y(new_n10346));
  nand_5 g09970(.A(pi133), .B(pi106), .Y(new_n10347));
  nand_5 g09971(.A(new_n9408), .B(new_n9407), .Y(new_n10348));
  nand_5 g09972(.A(new_n9409), .B(new_n9385), .Y(new_n10349));
  nand_5 g09973(.A(new_n10349), .B(new_n10348), .Y(new_n10350));
  xor_4  g09974(.A(new_n10350), .B(new_n10347), .Y(new_n10351));
  xor_4  g09975(.A(new_n10351), .B(new_n10346), .Y(new_n10352));
  xor_4  g09976(.A(new_n10352), .B(new_n10343), .Y(new_n10353));
  nand_5 g09977(.A(pi168), .B(pi017), .Y(new_n10354));
  nand_5 g09978(.A(new_n9420), .B(new_n9417), .Y(new_n10355));
  nand_5 g09979(.A(new_n9421), .B(new_n9413), .Y(new_n10356));
  nand_5 g09980(.A(new_n10356), .B(new_n10355), .Y(new_n10357));
  xor_4  g09981(.A(new_n10357), .B(new_n10354), .Y(new_n10358));
  or_6   g09982(.A(new_n9594), .B(new_n9551), .Y(new_n10359));
  nand_5 g09983(.A(new_n9595), .B(new_n9591), .Y(new_n10360));
  nand_5 g09984(.A(new_n10360), .B(new_n10359), .Y(new_n10361));
  nor_5  g09985(.A(new_n9596), .B(new_n9574), .Y(new_n10362));
  nor_5  g09986(.A(new_n9600), .B(new_n9597), .Y(new_n10363));
  nor_5  g09987(.A(new_n10363), .B(new_n10362), .Y(new_n10364));
  xor_4  g09988(.A(new_n10364), .B(new_n10361), .Y(new_n10365));
  nand_5 g09989(.A(pi208), .B(pi157), .Y(new_n10366));
  nand_5 g09990(.A(new_n9464), .B(new_n9463), .Y(new_n10367));
  nand_5 g09991(.A(new_n9465), .B(new_n9440), .Y(new_n10368));
  nand_5 g09992(.A(new_n10368), .B(new_n10367), .Y(new_n10369));
  or_6   g09993(.A(new_n9467), .B(new_n9441), .Y(new_n10370));
  not_8  g09994(.A(new_n9466), .Y(new_n10371));
  nand_5 g09995(.A(new_n9468), .B(new_n10371), .Y(new_n10372));
  nand_5 g09996(.A(new_n10372), .B(new_n10370), .Y(new_n10373));
  xor_4  g09997(.A(new_n10373), .B(new_n10369), .Y(new_n10374));
  xor_4  g09998(.A(new_n10374), .B(new_n10366), .Y(new_n10375));
  xor_4  g09999(.A(new_n10375), .B(new_n10365), .Y(new_n10376));
  nand_5 g10000(.A(pi204), .B(pi125), .Y(new_n10377));
  nand_5 g10001(.A(new_n9471), .B(new_n9470), .Y(new_n10378));
  nand_5 g10002(.A(new_n9472), .B(new_n9454), .Y(new_n10379));
  nand_5 g10003(.A(new_n10379), .B(new_n10378), .Y(new_n10380));
  nand_5 g10004(.A(pi040), .B(pi035), .Y(new_n10381));
  nand_5 g10005(.A(pi174), .B(pi139), .Y(new_n10382));
  xor_4  g10006(.A(new_n10382), .B(new_n10381), .Y(new_n10383));
  xor_4  g10007(.A(new_n10383), .B(new_n10380), .Y(new_n10384));
  xor_4  g10008(.A(new_n10384), .B(new_n10377), .Y(new_n10385));
  nand_5 g10009(.A(pi176), .B(pi015), .Y(new_n10386));
  nand_5 g10010(.A(new_n9476), .B(new_n9473), .Y(new_n10387));
  nand_5 g10011(.A(new_n9477), .B(new_n9469), .Y(new_n10388));
  nand_5 g10012(.A(new_n10388), .B(new_n10387), .Y(new_n10389));
  xor_4  g10013(.A(new_n10389), .B(new_n10386), .Y(new_n10390));
  xor_4  g10014(.A(new_n10390), .B(new_n10385), .Y(new_n10391));
  xor_4  g10015(.A(new_n10391), .B(new_n10376), .Y(new_n10392));
  nand_5 g10016(.A(pi222), .B(pi146), .Y(new_n10393));
  nand_5 g10017(.A(pi249), .B(pi152), .Y(new_n10394));
  nor_5  g10018(.A(new_n9483), .B(new_n9478), .Y(new_n10395));
  nor_5  g10019(.A(new_n10395), .B(new_n9482), .Y(new_n10396));
  xor_4  g10020(.A(new_n10396), .B(new_n10394), .Y(new_n10397));
  xor_4  g10021(.A(new_n10397), .B(new_n10393), .Y(new_n10398));
  xor_4  g10022(.A(new_n10398), .B(new_n10392), .Y(new_n10399));
  xor_4  g10023(.A(new_n10399), .B(new_n10358), .Y(new_n10400));
  or_6   g10024(.A(new_n9484), .B(new_n9462), .Y(new_n10401));
  nand_5 g10025(.A(new_n9492), .B(new_n9485), .Y(new_n10402));
  nand_5 g10026(.A(new_n10402), .B(new_n10401), .Y(new_n10403));
  nand_5 g10027(.A(pi227), .B(pi064), .Y(new_n10404));
  nand_5 g10028(.A(pi100), .B(pi084), .Y(new_n10405));
  xor_4  g10029(.A(new_n10405), .B(new_n10404), .Y(new_n10406));
  nand_5 g10030(.A(pi189), .B(pi081), .Y(new_n10407));
  xor_4  g10031(.A(new_n10407), .B(new_n10406), .Y(new_n10408));
  nand_5 g10032(.A(pi187), .B(pi052), .Y(new_n10409));
  or_6   g10033(.A(new_n9411), .B(new_n9386), .Y(new_n10410));
  not_8  g10034(.A(new_n9410), .Y(new_n10411));
  nand_5 g10035(.A(new_n9412), .B(new_n10411), .Y(new_n10412));
  nand_5 g10036(.A(new_n10412), .B(new_n10410), .Y(new_n10413));
  xor_4  g10037(.A(new_n10413), .B(new_n10409), .Y(new_n10414));
  nand_5 g10038(.A(pi233), .B(pi077), .Y(new_n10415));
  xor_4  g10039(.A(new_n10415), .B(new_n10414), .Y(new_n10416));
  xor_4  g10040(.A(new_n10416), .B(new_n10408), .Y(new_n10417));
  xor_4  g10041(.A(new_n10417), .B(new_n10403), .Y(new_n10418));
  xor_4  g10042(.A(new_n10418), .B(new_n10400), .Y(new_n10419));
  xor_4  g10043(.A(new_n10419), .B(new_n10353), .Y(new_n10420));
  xor_4  g10044(.A(new_n10420), .B(new_n10332), .Y(new_n10421));
  xor_4  g10045(.A(new_n10421), .B(new_n10329), .Y(new_n10422));
  nand_5 g10046(.A(new_n9604), .B(new_n9603), .Y(new_n10423));
  nand_5 g10047(.A(new_n9605), .B(new_n9505), .Y(new_n10424));
  nand_5 g10048(.A(new_n10424), .B(new_n10423), .Y(new_n10425));
  or_6   g10049(.A(new_n9617), .B(new_n9614), .Y(new_n10426));
  nand_5 g10050(.A(new_n9618), .B(new_n9610), .Y(new_n10427));
  nand_5 g10051(.A(new_n10427), .B(new_n10426), .Y(new_n10428));
  nand_5 g10052(.A(pi241), .B(pi021), .Y(new_n10429));
  nand_5 g10053(.A(pi161), .B(pi005), .Y(new_n10430));
  xor_4  g10054(.A(new_n10430), .B(new_n10429), .Y(new_n10431));
  xor_4  g10055(.A(new_n10431), .B(new_n10428), .Y(new_n10432));
  xor_4  g10056(.A(new_n10432), .B(new_n10425), .Y(new_n10433));
  nand_5 g10057(.A(new_n9405), .B(new_n9394), .Y(new_n10434));
  nand_5 g10058(.A(new_n9422), .B(new_n9406), .Y(new_n10435));
  nand_5 g10059(.A(new_n10435), .B(new_n10434), .Y(new_n10436));
  nand_5 g10060(.A(pi252), .B(pi047), .Y(new_n10437));
  nand_5 g10061(.A(new_n9576), .B(new_n9575), .Y(new_n10438));
  nand_5 g10062(.A(new_n9577), .B(new_n9542), .Y(new_n10439));
  nand_5 g10063(.A(new_n10439), .B(new_n10438), .Y(new_n10440));
  nand_5 g10064(.A(new_n9584), .B(new_n9583), .Y(new_n10441));
  nand_5 g10065(.A(new_n9585), .B(new_n9550), .Y(new_n10442));
  nand_5 g10066(.A(new_n10442), .B(new_n10441), .Y(new_n10443));
  xor_4  g10067(.A(new_n10443), .B(new_n10440), .Y(new_n10444));
  nand_5 g10068(.A(pi224), .B(pi112), .Y(new_n10445));
  xor_4  g10069(.A(new_n10445), .B(new_n10444), .Y(new_n10446));
  or_6   g10070(.A(new_n9580), .B(new_n9543), .Y(new_n10447));
  nand_5 g10071(.A(new_n9581), .B(new_n9579), .Y(new_n10448));
  nand_5 g10072(.A(new_n10448), .B(new_n10447), .Y(new_n10449));
  nand_5 g10073(.A(pi232), .B(pi212), .Y(new_n10450));
  nand_5 g10074(.A(pi127), .B(pi104), .Y(new_n10451));
  xor_4  g10075(.A(new_n10451), .B(new_n10450), .Y(new_n10452));
  nand_5 g10076(.A(pi255), .B(pi013), .Y(new_n10453));
  nand_5 g10077(.A(new_n9589), .B(new_n9586), .Y(new_n10454));
  not_8  g10078(.A(new_n9582), .Y(new_n10455));
  nand_5 g10079(.A(new_n9590), .B(new_n10455), .Y(new_n10456));
  nand_5 g10080(.A(new_n10456), .B(new_n10454), .Y(new_n10457));
  xnor_4 g10081(.A(new_n10457), .B(new_n10453), .Y(new_n10458));
  xor_4  g10082(.A(new_n10458), .B(new_n10452), .Y(new_n10459));
  xor_4  g10083(.A(new_n10459), .B(new_n10449), .Y(new_n10460));
  xor_4  g10084(.A(new_n10460), .B(new_n10446), .Y(new_n10461));
  xor_4  g10085(.A(new_n10461), .B(new_n10437), .Y(new_n10462));
  xor_4  g10086(.A(new_n10462), .B(new_n10436), .Y(new_n10463));
  nand_5 g10087(.A(new_n9639), .B(new_n9432), .Y(new_n10464));
  nand_5 g10088(.A(new_n9649), .B(new_n9640), .Y(new_n10465));
  nand_5 g10089(.A(new_n10465), .B(new_n10464), .Y(new_n10466));
  nand_5 g10090(.A(pi140), .B(pi018), .Y(new_n10467));
  nand_5 g10091(.A(pi242), .B(pi128), .Y(new_n10468));
  xor_4  g10092(.A(new_n10468), .B(new_n10467), .Y(new_n10469));
  or_6   g10093(.A(new_n9626), .B(new_n9602), .Y(new_n10470));
  nand_5 g10094(.A(new_n9631), .B(new_n9627), .Y(new_n10471));
  nand_5 g10095(.A(new_n10471), .B(new_n10470), .Y(new_n10472));
  nand_5 g10096(.A(pi236), .B(pi082), .Y(new_n10473));
  xor_4  g10097(.A(new_n10473), .B(new_n10472), .Y(new_n10474));
  xor_4  g10098(.A(new_n10474), .B(new_n10469), .Y(new_n10475));
  or_6   g10099(.A(new_n9625), .B(new_n9619), .Y(new_n10476));
  nand_5 g10100(.A(new_n10476), .B(new_n9624), .Y(new_n10477));
  nand_5 g10101(.A(pi121), .B(pi090), .Y(new_n10478));
  nand_5 g10102(.A(pi231), .B(pi141), .Y(new_n10479));
  xor_4  g10103(.A(new_n10479), .B(new_n10478), .Y(new_n10480));
  xor_4  g10104(.A(new_n10480), .B(new_n10477), .Y(new_n10481));
  xor_4  g10105(.A(new_n10481), .B(new_n10475), .Y(new_n10482));
  xor_4  g10106(.A(new_n10482), .B(new_n10466), .Y(new_n10483));
  xor_4  g10107(.A(new_n10483), .B(new_n10463), .Y(new_n10484));
  nor_5  g10108(.A(new_n9570), .B(new_n9493), .Y(new_n10485));
  nor_5  g10109(.A(new_n9638), .B(new_n9572), .Y(new_n10486));
  or_6   g10110(.A(new_n10486), .B(new_n10485), .Y(new_n10487));
  nand_5 g10111(.A(pi217), .B(pi034), .Y(new_n10488));
  nand_5 g10112(.A(pi131), .B(pi129), .Y(new_n10489));
  xor_4  g10113(.A(new_n10489), .B(new_n10488), .Y(new_n10490));
  xor_4  g10114(.A(new_n10490), .B(new_n10487), .Y(new_n10491));
  xor_4  g10115(.A(new_n10491), .B(new_n10484), .Y(new_n10492));
  xor_4  g10116(.A(new_n10492), .B(new_n10433), .Y(new_n10493));
  xor_4  g10117(.A(new_n10493), .B(new_n10422), .Y(po086));
  xnor_4 g10118(.A(new_n7522), .B(new_n7521), .Y(po087));
  xnor_4 g10119(.A(new_n4804), .B(new_n4803), .Y(po088));
  xor_4  g10120(.A(new_n3088), .B(new_n3067), .Y(po089));
  xor_4  g10121(.A(new_n2562), .B(new_n2561), .Y(po090));
  xor_4  g10122(.A(new_n3501), .B(new_n3499), .Y(po091));
  xnor_4 g10123(.A(new_n5677), .B(new_n5667), .Y(po092));
  xor_4  g10124(.A(new_n9189), .B(new_n9160), .Y(po093));
  xor_4  g10125(.A(new_n901), .B(new_n899), .Y(po094));
  xor_4  g10126(.A(new_n1050), .B(new_n1049), .Y(po095));
  xor_4  g10127(.A(new_n3506), .B(new_n3505), .Y(po096));
  nand_5 g10128(.A(pi243), .B(pi213), .Y(new_n10505));
  or_6   g10129(.A(new_n5142), .B(new_n5119), .Y(new_n10506));
  nand_5 g10130(.A(new_n5152), .B(new_n5143), .Y(new_n10507));
  nand_5 g10131(.A(new_n10507), .B(new_n10506), .Y(new_n10508));
  nor_5  g10132(.A(new_n5141), .B(new_n5135), .Y(new_n10509));
  nor_5  g10133(.A(new_n10509), .B(new_n5140), .Y(new_n10510));
  xor_4  g10134(.A(new_n10510), .B(new_n10508), .Y(new_n10511));
  xor_4  g10135(.A(new_n10511), .B(new_n10505), .Y(new_n10512));
  nand_5 g10136(.A(pi207), .B(pi183), .Y(new_n10513));
  nand_5 g10137(.A(pi105), .B(pi066), .Y(new_n10514));
  xor_4  g10138(.A(new_n10514), .B(new_n10513), .Y(new_n10515));
  nand_5 g10139(.A(pi226), .B(pi088), .Y(new_n10516));
  xor_4  g10140(.A(new_n10516), .B(new_n10515), .Y(new_n10517));
  nand_5 g10141(.A(new_n5224), .B(new_n5223), .Y(new_n10518));
  nand_5 g10142(.A(new_n5225), .B(new_n5193), .Y(new_n10519));
  nand_5 g10143(.A(new_n10519), .B(new_n10518), .Y(new_n10520));
  not_8  g10144(.A(new_n5153), .Y(new_n10521));
  nand_5 g10145(.A(new_n10521), .B(new_n5074), .Y(new_n10522));
  or_6   g10146(.A(new_n5171), .B(new_n5154), .Y(new_n10523));
  nand_5 g10147(.A(new_n10523), .B(new_n10522), .Y(new_n10524));
  xor_4  g10148(.A(new_n10524), .B(new_n10520), .Y(new_n10525));
  xor_4  g10149(.A(new_n10525), .B(new_n10517), .Y(new_n10526));
  xor_4  g10150(.A(new_n10526), .B(new_n10512), .Y(new_n10527));
  nand_5 g10151(.A(pi218), .B(pi208), .Y(new_n10528));
  nand_5 g10152(.A(new_n5217), .B(new_n5216), .Y(new_n10529));
  nand_5 g10153(.A(new_n5218), .B(new_n5178), .Y(new_n10530));
  nand_5 g10154(.A(new_n10530), .B(new_n10529), .Y(new_n10531));
  or_6   g10155(.A(new_n5220), .B(new_n5179), .Y(new_n10532));
  not_8  g10156(.A(new_n5219), .Y(new_n10533));
  nand_5 g10157(.A(new_n5221), .B(new_n10533), .Y(new_n10534));
  nand_5 g10158(.A(new_n10534), .B(new_n10532), .Y(new_n10535));
  xor_4  g10159(.A(new_n10535), .B(new_n10531), .Y(new_n10536));
  xor_4  g10160(.A(new_n10536), .B(new_n10528), .Y(new_n10537));
  xor_4  g10161(.A(new_n10537), .B(new_n10527), .Y(new_n10538));
  nand_5 g10162(.A(pi204), .B(pi058), .Y(new_n10539));
  or_6   g10163(.A(new_n5316), .B(new_n5275), .Y(new_n10540));
  not_8  g10164(.A(new_n5315), .Y(new_n10541));
  nand_5 g10165(.A(new_n5317), .B(new_n10541), .Y(new_n10542));
  nand_5 g10166(.A(new_n10542), .B(new_n10540), .Y(new_n10543));
  nand_5 g10167(.A(pi199), .B(pi035), .Y(new_n10544));
  nand_5 g10168(.A(pi195), .B(pi139), .Y(new_n10545));
  xor_4  g10169(.A(new_n10545), .B(new_n10544), .Y(new_n10546));
  xor_4  g10170(.A(new_n10546), .B(new_n10543), .Y(new_n10547));
  xor_4  g10171(.A(new_n10547), .B(new_n10539), .Y(new_n10548));
  nand_5 g10172(.A(pi211), .B(pi015), .Y(new_n10549));
  nand_5 g10173(.A(new_n5229), .B(new_n5226), .Y(new_n10550));
  nand_5 g10174(.A(new_n5230), .B(new_n5222), .Y(new_n10551));
  nand_5 g10175(.A(new_n10551), .B(new_n10550), .Y(new_n10552));
  xor_4  g10176(.A(new_n10552), .B(new_n10549), .Y(new_n10553));
  xor_4  g10177(.A(new_n10553), .B(new_n10548), .Y(new_n10554));
  xor_4  g10178(.A(new_n10554), .B(new_n10538), .Y(new_n10555));
  nand_5 g10179(.A(new_n5044), .B(new_n5043), .Y(new_n10556));
  nand_5 g10180(.A(new_n5045), .B(new_n5005), .Y(new_n10557));
  nand_5 g10181(.A(new_n10557), .B(new_n10556), .Y(new_n10558));
  nand_5 g10182(.A(new_n5051), .B(new_n5050), .Y(new_n10559));
  nand_5 g10183(.A(new_n5052), .B(new_n5020), .Y(new_n10560));
  nand_5 g10184(.A(new_n10560), .B(new_n10559), .Y(new_n10561));
  xor_4  g10185(.A(new_n10561), .B(new_n10558), .Y(new_n10562));
  or_6   g10186(.A(new_n5047), .B(new_n5006), .Y(new_n10563));
  not_8  g10187(.A(new_n5046), .Y(new_n10564));
  nand_5 g10188(.A(new_n5048), .B(new_n10564), .Y(new_n10565));
  nand_5 g10189(.A(new_n10565), .B(new_n10563), .Y(new_n10566));
  xor_4  g10190(.A(new_n10566), .B(new_n10562), .Y(new_n10567));
  xor_4  g10191(.A(new_n10567), .B(new_n10555), .Y(new_n10568));
  nand_5 g10192(.A(new_n5329), .B(new_n5290), .Y(new_n10569));
  nand_5 g10193(.A(new_n5332), .B(new_n5327), .Y(new_n10570));
  nand_5 g10194(.A(new_n10570), .B(new_n10569), .Y(new_n10571));
  not_8  g10195(.A(new_n5333), .Y(new_n10572));
  nor_5  g10196(.A(new_n10572), .B(new_n5311), .Y(new_n10573));
  nor_5  g10197(.A(new_n5345), .B(new_n5334), .Y(new_n10574));
  nor_5  g10198(.A(new_n10574), .B(new_n10573), .Y(new_n10575));
  xor_4  g10199(.A(new_n10575), .B(new_n10571), .Y(new_n10576));
  nand_5 g10200(.A(pi034), .B(pi029), .Y(new_n10577));
  nand_5 g10201(.A(pi131), .B(pi010), .Y(new_n10578));
  xor_4  g10202(.A(new_n10578), .B(new_n10577), .Y(new_n10579));
  nand_5 g10203(.A(new_n5056), .B(new_n5053), .Y(new_n10580));
  nand_5 g10204(.A(new_n5057), .B(new_n5049), .Y(new_n10581));
  nand_5 g10205(.A(new_n10581), .B(new_n10580), .Y(new_n10582));
  nand_5 g10206(.A(pi241), .B(pi074), .Y(new_n10583));
  nand_5 g10207(.A(pi253), .B(pi161), .Y(new_n10584));
  xor_4  g10208(.A(new_n10584), .B(new_n10583), .Y(new_n10585));
  xor_4  g10209(.A(new_n10585), .B(new_n10582), .Y(new_n10586));
  xor_4  g10210(.A(new_n10586), .B(new_n10579), .Y(new_n10587));
  xor_4  g10211(.A(new_n10587), .B(new_n10576), .Y(new_n10588));
  xor_4  g10212(.A(new_n10588), .B(new_n10568), .Y(new_n10589));
  nand_5 g10213(.A(pi084), .B(pi069), .Y(new_n10590));
  nand_5 g10214(.A(new_n5313), .B(new_n5312), .Y(new_n10591));
  nand_5 g10215(.A(new_n5314), .B(new_n5274), .Y(new_n10592));
  nand_5 g10216(.A(new_n10592), .B(new_n10591), .Y(new_n10593));
  xor_4  g10217(.A(new_n10593), .B(new_n10590), .Y(new_n10594));
  xor_4  g10218(.A(new_n10594), .B(new_n10589), .Y(new_n10595));
  nand_5 g10219(.A(new_n5245), .B(new_n5236), .Y(new_n10596));
  nand_5 g10220(.A(new_n5246), .B(new_n5215), .Y(new_n10597));
  nand_5 g10221(.A(new_n10597), .B(new_n10596), .Y(new_n10598));
  nand_5 g10222(.A(pi189), .B(pi150), .Y(new_n10599));
  nand_5 g10223(.A(pi221), .B(pi133), .Y(new_n10600));
  xor_4  g10224(.A(new_n10600), .B(new_n10599), .Y(new_n10601));
  xor_4  g10225(.A(new_n10601), .B(new_n10598), .Y(new_n10602));
  not_8  g10226(.A(new_n5247), .Y(new_n10603));
  nor_5  g10227(.A(new_n10603), .B(new_n5172), .Y(new_n10604));
  nor_5  g10228(.A(new_n5267), .B(new_n5248), .Y(new_n10605));
  nor_5  g10229(.A(new_n10605), .B(new_n10604), .Y(new_n10606));
  nand_5 g10230(.A(pi244), .B(pi064), .Y(new_n10607));
  xor_4  g10231(.A(new_n10607), .B(new_n10606), .Y(new_n10608));
  xor_4  g10232(.A(new_n10608), .B(new_n10602), .Y(new_n10609));
  nand_5 g10233(.A(pi184), .B(pi052), .Y(new_n10610));
  nand_5 g10234(.A(pi196), .B(pi077), .Y(new_n10611));
  xor_4  g10235(.A(new_n10611), .B(new_n10610), .Y(new_n10612));
  nand_5 g10236(.A(new_n5325), .B(new_n5322), .Y(new_n10613));
  nand_5 g10237(.A(new_n5326), .B(new_n5318), .Y(new_n10614));
  nand_5 g10238(.A(new_n10614), .B(new_n10613), .Y(new_n10615));
  nand_5 g10239(.A(pi186), .B(pi146), .Y(new_n10616));
  nand_5 g10240(.A(pi168), .B(pi037), .Y(new_n10617));
  xor_4  g10241(.A(new_n10617), .B(new_n10616), .Y(new_n10618));
  xor_4  g10242(.A(new_n10618), .B(new_n10615), .Y(new_n10619));
  nand_5 g10243(.A(pi152), .B(pi132), .Y(new_n10620));
  nand_5 g10244(.A(new_n5233), .B(new_n5194), .Y(new_n10621));
  not_8  g10245(.A(new_n5235), .Y(new_n10622));
  nand_5 g10246(.A(new_n10622), .B(new_n5231), .Y(new_n10623));
  nand_5 g10247(.A(new_n10623), .B(new_n10621), .Y(new_n10624));
  xor_4  g10248(.A(new_n10624), .B(new_n10620), .Y(new_n10625));
  nand_5 g10249(.A(new_n5320), .B(new_n5319), .Y(new_n10626));
  nand_5 g10250(.A(new_n5321), .B(new_n5289), .Y(new_n10627));
  nand_5 g10251(.A(new_n10627), .B(new_n10626), .Y(new_n10628));
  xor_4  g10252(.A(new_n10628), .B(new_n10625), .Y(new_n10629));
  xor_4  g10253(.A(new_n10629), .B(new_n10619), .Y(new_n10630));
  xor_4  g10254(.A(new_n10630), .B(new_n10612), .Y(new_n10631));
  xor_4  g10255(.A(new_n10631), .B(new_n10609), .Y(new_n10632));
  xor_4  g10256(.A(new_n10632), .B(new_n10595), .Y(new_n10633));
  nand_5 g10257(.A(new_n5060), .B(new_n5021), .Y(new_n10634));
  not_8  g10258(.A(new_n5062), .Y(new_n10635));
  nand_5 g10259(.A(new_n10635), .B(new_n5058), .Y(new_n10636));
  nand_5 g10260(.A(new_n10636), .B(new_n10634), .Y(new_n10637));
  nand_5 g10261(.A(pi173), .B(pi047), .Y(new_n10638));
  nand_5 g10262(.A(pi018), .B(pi014), .Y(new_n10639));
  xor_4  g10263(.A(new_n10639), .B(new_n10638), .Y(new_n10640));
  xor_4  g10264(.A(new_n10640), .B(new_n10637), .Y(new_n10641));
  xor_4  g10265(.A(new_n10641), .B(new_n10633), .Y(new_n10642));
  nand_5 g10266(.A(pi230), .B(pi090), .Y(new_n10643));
  nand_5 g10267(.A(pi141), .B(pi050), .Y(new_n10644));
  xor_4  g10268(.A(new_n10644), .B(new_n10643), .Y(new_n10645));
  nand_5 g10269(.A(new_n5133), .B(new_n5130), .Y(new_n10646));
  nand_5 g10270(.A(new_n5134), .B(new_n5126), .Y(new_n10647));
  nand_5 g10271(.A(new_n10647), .B(new_n10646), .Y(new_n10648));
  nand_5 g10272(.A(new_n5128), .B(new_n5127), .Y(new_n10649));
  nand_5 g10273(.A(new_n5129), .B(new_n5095), .Y(new_n10650));
  nand_5 g10274(.A(new_n10650), .B(new_n10649), .Y(new_n10651));
  xor_4  g10275(.A(new_n10651), .B(new_n10648), .Y(new_n10652));
  nand_5 g10276(.A(pi112), .B(pi055), .Y(new_n10653));
  or_6   g10277(.A(new_n5124), .B(new_n5087), .Y(new_n10654));
  not_8  g10278(.A(new_n5123), .Y(new_n10655));
  nand_5 g10279(.A(new_n5125), .B(new_n10655), .Y(new_n10656));
  nand_5 g10280(.A(new_n10656), .B(new_n10654), .Y(new_n10657));
  nand_5 g10281(.A(pi239), .B(pi212), .Y(new_n10658));
  nand_5 g10282(.A(pi104), .B(pi025), .Y(new_n10659));
  xor_4  g10283(.A(new_n10659), .B(new_n10658), .Y(new_n10660));
  xor_4  g10284(.A(new_n10660), .B(new_n10657), .Y(new_n10661));
  xor_4  g10285(.A(new_n10661), .B(new_n10653), .Y(new_n10662));
  nand_5 g10286(.A(pi013), .B(pi002), .Y(new_n10663));
  nand_5 g10287(.A(new_n5121), .B(new_n5120), .Y(new_n10664));
  nand_5 g10288(.A(new_n5122), .B(new_n5086), .Y(new_n10665));
  nand_5 g10289(.A(new_n10665), .B(new_n10664), .Y(new_n10666));
  xor_4  g10290(.A(new_n10666), .B(new_n10663), .Y(new_n10667));
  xor_4  g10291(.A(new_n10667), .B(new_n10662), .Y(new_n10668));
  xor_4  g10292(.A(new_n10668), .B(new_n10652), .Y(new_n10669));
  xor_4  g10293(.A(new_n10669), .B(new_n10645), .Y(new_n10670));
  nor_5  g10294(.A(new_n5346), .B(new_n5268), .Y(new_n10671));
  not_8  g10295(.A(new_n5347), .Y(new_n10672));
  nor_5  g10296(.A(new_n5363), .B(new_n10672), .Y(new_n10673));
  nor_5  g10297(.A(new_n10673), .B(new_n10671), .Y(new_n10674));
  nand_5 g10298(.A(pi236), .B(pi205), .Y(new_n10675));
  xor_4  g10299(.A(new_n10675), .B(new_n10674), .Y(new_n10676));
  xor_4  g10300(.A(new_n10676), .B(new_n10670), .Y(new_n10677));
  nor_5  g10301(.A(new_n5063), .B(new_n5042), .Y(new_n10678));
  nor_5  g10302(.A(new_n5073), .B(new_n5064), .Y(new_n10679));
  nor_5  g10303(.A(new_n10679), .B(new_n10678), .Y(new_n10680));
  nand_5 g10304(.A(pi128), .B(pi109), .Y(new_n10681));
  xor_4  g10305(.A(new_n10681), .B(new_n10680), .Y(new_n10682));
  xor_4  g10306(.A(new_n10682), .B(new_n10677), .Y(new_n10683));
  xor_4  g10307(.A(new_n10683), .B(new_n10642), .Y(po097));
  xor_4  g10308(.A(new_n1803), .B(new_n1801), .Y(po098));
  xnor_4 g10309(.A(new_n7741), .B(new_n7740), .Y(po099));
  xnor_4 g10310(.A(new_n890), .B(new_n889), .Y(po100));
  xor_4  g10311(.A(new_n887), .B(new_n885), .Y(po101));
  xor_4  g10312(.A(new_n1045), .B(new_n1043), .Y(po102));
  xor_4  g10313(.A(new_n3116), .B(new_n3115), .Y(po103));
  xor_4  g10314(.A(new_n2554), .B(new_n1986), .Y(po104));
  xnor_4 g10315(.A(new_n3695), .B(new_n3694), .Y(po105));
  xor_4  g10316(.A(new_n5764), .B(new_n5762), .Y(po106));
  xor_4  g10317(.A(new_n9192), .B(new_n9191), .Y(po107));
  xor_4  g10318(.A(new_n3683), .B(new_n3607), .Y(po108));
  or_6   g10319(.A(new_n4530), .B(new_n4496), .Y(new_n10696));
  not_8  g10320(.A(new_n4529), .Y(new_n10697));
  nand_5 g10321(.A(new_n4531), .B(new_n10697), .Y(new_n10698));
  nand_5 g10322(.A(new_n10698), .B(new_n10696), .Y(new_n10699));
  nand_5 g10323(.A(pi103), .B(pi046), .Y(new_n10700));
  nor_5  g10324(.A(new_n4546), .B(new_n4525), .Y(new_n10701));
  not_8  g10325(.A(new_n4547), .Y(new_n10702));
  nor_5  g10326(.A(new_n4556), .B(new_n10702), .Y(new_n10703));
  nor_5  g10327(.A(new_n10703), .B(new_n10701), .Y(new_n10704));
  xor_4  g10328(.A(new_n10704), .B(new_n10700), .Y(new_n10705));
  xor_4  g10329(.A(new_n10705), .B(new_n10699), .Y(new_n10706));
  nand_5 g10330(.A(pi188), .B(pi000), .Y(new_n10707));
  nand_5 g10331(.A(pi178), .B(pi115), .Y(new_n10708));
  nand_5 g10332(.A(pi070), .B(pi061), .Y(new_n10709));
  xor_4  g10333(.A(new_n10709), .B(new_n10708), .Y(new_n10710));
  nand_5 g10334(.A(new_n4439), .B(new_n4438), .Y(new_n10711));
  nand_5 g10335(.A(new_n4440), .B(new_n4407), .Y(new_n10712));
  nand_5 g10336(.A(new_n10712), .B(new_n10711), .Y(new_n10713));
  nand_5 g10337(.A(pi167), .B(pi048), .Y(new_n10714));
  or_6   g10338(.A(new_n4435), .B(new_n4400), .Y(new_n10715));
  not_8  g10339(.A(new_n4434), .Y(new_n10716));
  nand_5 g10340(.A(new_n4436), .B(new_n10716), .Y(new_n10717));
  nand_5 g10341(.A(new_n10717), .B(new_n10715), .Y(new_n10718));
  xor_4  g10342(.A(new_n10718), .B(new_n10714), .Y(new_n10719));
  xor_4  g10343(.A(new_n10719), .B(new_n10713), .Y(new_n10720));
  nand_5 g10344(.A(new_n4353), .B(new_n4313), .Y(new_n10721));
  nand_5 g10345(.A(new_n4356), .B(new_n4351), .Y(new_n10722));
  nand_5 g10346(.A(new_n10722), .B(new_n10721), .Y(new_n10723));
  nand_5 g10347(.A(pi237), .B(pi149), .Y(new_n10724));
  nand_5 g10348(.A(pi240), .B(pi238), .Y(new_n10725));
  xor_4  g10349(.A(new_n10725), .B(new_n10724), .Y(new_n10726));
  nand_5 g10350(.A(pi181), .B(pi179), .Y(new_n10727));
  xor_4  g10351(.A(new_n10727), .B(new_n10726), .Y(new_n10728));
  nand_5 g10352(.A(pi193), .B(pi134), .Y(new_n10729));
  nand_5 g10353(.A(new_n4444), .B(new_n4441), .Y(new_n10730));
  nand_5 g10354(.A(new_n4445), .B(new_n4437), .Y(new_n10731));
  nand_5 g10355(.A(new_n10731), .B(new_n10730), .Y(new_n10732));
  xor_4  g10356(.A(new_n10732), .B(new_n10729), .Y(new_n10733));
  nand_5 g10357(.A(new_n4432), .B(new_n4431), .Y(new_n10734));
  nand_5 g10358(.A(new_n4433), .B(new_n4399), .Y(new_n10735));
  nand_5 g10359(.A(new_n10735), .B(new_n10734), .Y(new_n10736));
  xor_4  g10360(.A(new_n10736), .B(new_n10733), .Y(new_n10737));
  xor_4  g10361(.A(new_n10737), .B(new_n10728), .Y(new_n10738));
  xor_4  g10362(.A(new_n10738), .B(new_n10723), .Y(new_n10739));
  xor_4  g10363(.A(new_n10739), .B(new_n10720), .Y(new_n10740));
  xor_4  g10364(.A(new_n10740), .B(new_n10710), .Y(new_n10741));
  xor_4  g10365(.A(new_n10741), .B(new_n10707), .Y(new_n10742));
  not_8  g10366(.A(new_n4452), .Y(new_n10743));
  nor_5  g10367(.A(new_n10743), .B(new_n4430), .Y(new_n10744));
  nor_5  g10368(.A(new_n4463), .B(new_n4453), .Y(new_n10745));
  nor_5  g10369(.A(new_n10745), .B(new_n10744), .Y(new_n10746));
  nand_5 g10370(.A(new_n4527), .B(new_n4526), .Y(new_n10747));
  nand_5 g10371(.A(new_n4528), .B(new_n4495), .Y(new_n10748));
  nand_5 g10372(.A(new_n10748), .B(new_n10747), .Y(new_n10749));
  nand_5 g10373(.A(new_n4539), .B(new_n4536), .Y(new_n10750));
  nand_5 g10374(.A(new_n4540), .B(new_n4532), .Y(new_n10751));
  nand_5 g10375(.A(new_n10751), .B(new_n10750), .Y(new_n10752));
  xor_4  g10376(.A(new_n10752), .B(new_n10749), .Y(new_n10753));
  nand_5 g10377(.A(pi117), .B(pi068), .Y(new_n10754));
  nand_5 g10378(.A(pi036), .B(pi016), .Y(new_n10755));
  xor_4  g10379(.A(new_n10755), .B(new_n10754), .Y(new_n10756));
  nand_5 g10380(.A(pi214), .B(pi057), .Y(new_n10757));
  xor_4  g10381(.A(new_n10757), .B(new_n10756), .Y(new_n10758));
  xor_4  g10382(.A(new_n10758), .B(new_n10753), .Y(new_n10759));
  xor_4  g10383(.A(new_n10759), .B(new_n10746), .Y(new_n10760));
  xor_4  g10384(.A(new_n10760), .B(new_n10742), .Y(new_n10761));
  nand_5 g10385(.A(new_n4464), .B(new_n4386), .Y(new_n10762));
  nand_5 g10386(.A(new_n4481), .B(new_n4465), .Y(new_n10763));
  nand_5 g10387(.A(new_n10763), .B(new_n10762), .Y(new_n10764));
  nand_5 g10388(.A(pi163), .B(pi126), .Y(new_n10765));
  not_8  g10389(.A(new_n4357), .Y(new_n10766));
  nor_5  g10390(.A(new_n10766), .B(new_n4335), .Y(new_n10767));
  nor_5  g10391(.A(new_n4367), .B(new_n4358), .Y(new_n10768));
  or_6   g10392(.A(new_n10768), .B(new_n10767), .Y(new_n10769));
  xor_4  g10393(.A(new_n10769), .B(new_n10765), .Y(new_n10770));
  nand_5 g10394(.A(new_n4369), .B(new_n4291), .Y(new_n10771));
  nand_5 g10395(.A(new_n4385), .B(new_n4370), .Y(new_n10772));
  nand_5 g10396(.A(new_n10772), .B(new_n10771), .Y(new_n10773));
  nand_5 g10397(.A(pi203), .B(pi162), .Y(new_n10774));
  nand_5 g10398(.A(new_n4448), .B(new_n4408), .Y(new_n10775));
  nand_5 g10399(.A(new_n4451), .B(new_n4446), .Y(new_n10776));
  nand_5 g10400(.A(new_n10776), .B(new_n10775), .Y(new_n10777));
  xor_4  g10401(.A(new_n10777), .B(new_n10774), .Y(new_n10778));
  nand_5 g10402(.A(pi200), .B(pi033), .Y(new_n10779));
  nand_5 g10403(.A(pi175), .B(pi159), .Y(new_n10780));
  xor_4  g10404(.A(new_n10780), .B(new_n10779), .Y(new_n10781));
  nand_5 g10405(.A(new_n4534), .B(new_n4533), .Y(new_n10782));
  nand_5 g10406(.A(new_n4535), .B(new_n4503), .Y(new_n10783));
  nand_5 g10407(.A(new_n10783), .B(new_n10782), .Y(new_n10784));
  xor_4  g10408(.A(new_n10784), .B(new_n10781), .Y(new_n10785));
  xor_4  g10409(.A(new_n10785), .B(new_n10778), .Y(new_n10786));
  nand_5 g10410(.A(pi234), .B(pi194), .Y(new_n10787));
  nand_5 g10411(.A(pi247), .B(pi085), .Y(new_n10788));
  nand_5 g10412(.A(pi180), .B(pi080), .Y(new_n10789));
  xor_4  g10413(.A(new_n10789), .B(new_n10788), .Y(new_n10790));
  xor_4  g10414(.A(new_n10790), .B(new_n10787), .Y(new_n10791));
  xor_4  g10415(.A(new_n10791), .B(new_n10786), .Y(new_n10792));
  xor_4  g10416(.A(new_n10792), .B(new_n10773), .Y(new_n10793));
  xor_4  g10417(.A(new_n10793), .B(new_n10770), .Y(new_n10794));
  xor_4  g10418(.A(new_n10794), .B(new_n10764), .Y(new_n10795));
  xor_4  g10419(.A(new_n10795), .B(new_n10761), .Y(new_n10796));
  nand_5 g10420(.A(new_n4344), .B(new_n4343), .Y(new_n10797));
  nand_5 g10421(.A(new_n4345), .B(new_n4312), .Y(new_n10798));
  nand_5 g10422(.A(new_n10798), .B(new_n10797), .Y(new_n10799));
  or_6   g10423(.A(new_n4340), .B(new_n4298), .Y(new_n10800));
  not_8  g10424(.A(new_n4339), .Y(new_n10801));
  nand_5 g10425(.A(new_n4341), .B(new_n10801), .Y(new_n10802));
  nand_5 g10426(.A(new_n10802), .B(new_n10800), .Y(new_n10803));
  xor_4  g10427(.A(new_n10803), .B(new_n10799), .Y(new_n10804));
  nand_5 g10428(.A(new_n4337), .B(new_n4336), .Y(new_n10805));
  nand_5 g10429(.A(new_n4338), .B(new_n4297), .Y(new_n10806));
  nand_5 g10430(.A(new_n10806), .B(new_n10805), .Y(new_n10807));
  nand_5 g10431(.A(pi116), .B(pi012), .Y(new_n10808));
  xor_4  g10432(.A(new_n10808), .B(new_n10807), .Y(new_n10809));
  xor_4  g10433(.A(new_n10809), .B(new_n10804), .Y(new_n10810));
  nand_5 g10434(.A(new_n4543), .B(new_n4504), .Y(new_n10811));
  not_8  g10435(.A(new_n4545), .Y(new_n10812));
  nand_5 g10436(.A(new_n10812), .B(new_n4541), .Y(new_n10813));
  nand_5 g10437(.A(new_n10813), .B(new_n10811), .Y(new_n10814));
  nand_5 g10438(.A(pi156), .B(pi108), .Y(new_n10815));
  nand_5 g10439(.A(pi083), .B(pi051), .Y(new_n10816));
  nand_5 g10440(.A(pi107), .B(pi028), .Y(new_n10817));
  xor_4  g10441(.A(new_n10817), .B(new_n10816), .Y(new_n10818));
  xor_4  g10442(.A(new_n10818), .B(new_n10815), .Y(new_n10819));
  nand_5 g10443(.A(pi201), .B(pi007), .Y(new_n10820));
  nand_5 g10444(.A(pi245), .B(pi118), .Y(new_n10821));
  xor_4  g10445(.A(new_n10821), .B(new_n10820), .Y(new_n10822));
  nand_5 g10446(.A(pi063), .B(pi042), .Y(new_n10823));
  xor_4  g10447(.A(new_n10823), .B(new_n10822), .Y(new_n10824));
  nand_5 g10448(.A(new_n4286), .B(new_n4252), .Y(new_n10825));
  not_8  g10449(.A(new_n4288), .Y(new_n10826));
  nand_5 g10450(.A(new_n10826), .B(new_n4284), .Y(new_n10827));
  nand_5 g10451(.A(new_n10827), .B(new_n10825), .Y(new_n10828));
  nand_5 g10452(.A(new_n4289), .B(new_n4267), .Y(new_n10829));
  nand_5 g10453(.A(new_n4290), .B(new_n4266), .Y(new_n10830));
  nand_5 g10454(.A(new_n10830), .B(new_n10829), .Y(new_n10831));
  xor_4  g10455(.A(new_n10831), .B(new_n10828), .Y(new_n10832));
  xor_4  g10456(.A(new_n10832), .B(new_n10824), .Y(new_n10833));
  xor_4  g10457(.A(new_n10833), .B(new_n10819), .Y(new_n10834));
  nand_5 g10458(.A(pi148), .B(pi043), .Y(new_n10835));
  nand_5 g10459(.A(pi228), .B(pi098), .Y(new_n10836));
  xor_4  g10460(.A(new_n10836), .B(new_n10835), .Y(new_n10837));
  nand_5 g10461(.A(pi144), .B(pi039), .Y(new_n10838));
  nand_5 g10462(.A(new_n4349), .B(new_n4346), .Y(new_n10839));
  nand_5 g10463(.A(new_n4350), .B(new_n4342), .Y(new_n10840));
  nand_5 g10464(.A(new_n10840), .B(new_n10839), .Y(new_n10841));
  xor_4  g10465(.A(new_n10841), .B(new_n10838), .Y(new_n10842));
  xor_4  g10466(.A(new_n10842), .B(new_n10837), .Y(new_n10843));
  xor_4  g10467(.A(new_n10843), .B(new_n10834), .Y(new_n10844));
  xor_4  g10468(.A(new_n10844), .B(new_n10814), .Y(new_n10845));
  xor_4  g10469(.A(new_n10845), .B(new_n10810), .Y(new_n10846));
  nand_5 g10470(.A(pi202), .B(pi143), .Y(new_n10847));
  nand_5 g10471(.A(new_n4574), .B(new_n4557), .Y(new_n10848));
  not_8  g10472(.A(new_n4482), .Y(new_n10849));
  nand_5 g10473(.A(new_n4575), .B(new_n10849), .Y(new_n10850));
  nand_5 g10474(.A(new_n10850), .B(new_n10848), .Y(new_n10851));
  nand_5 g10475(.A(pi171), .B(pi038), .Y(new_n10852));
  nand_5 g10476(.A(pi113), .B(pi049), .Y(new_n10853));
  xor_4  g10477(.A(new_n10853), .B(new_n10852), .Y(new_n10854));
  xor_4  g10478(.A(new_n10854), .B(new_n10851), .Y(new_n10855));
  or_6   g10479(.A(new_n4273), .B(new_n4241), .Y(new_n10856));
  nand_5 g10480(.A(new_n4274), .B(new_n4272), .Y(new_n10857));
  nand_5 g10481(.A(new_n10857), .B(new_n10856), .Y(new_n10858));
  or_6   g10482(.A(new_n4282), .B(new_n4279), .Y(new_n10859));
  nand_5 g10483(.A(new_n4283), .B(new_n4275), .Y(new_n10860));
  nand_5 g10484(.A(new_n10860), .B(new_n10859), .Y(new_n10861));
  nand_5 g10485(.A(new_n4269), .B(new_n4268), .Y(new_n10862));
  nand_5 g10486(.A(new_n4270), .B(new_n4240), .Y(new_n10863));
  nand_5 g10487(.A(new_n10863), .B(new_n10862), .Y(new_n10864));
  nand_5 g10488(.A(new_n4277), .B(new_n4276), .Y(new_n10865));
  nand_5 g10489(.A(new_n4278), .B(new_n4251), .Y(new_n10866));
  nand_5 g10490(.A(new_n10866), .B(new_n10865), .Y(new_n10867));
  xor_4  g10491(.A(new_n10867), .B(new_n10864), .Y(new_n10868));
  xor_4  g10492(.A(new_n10868), .B(new_n10861), .Y(new_n10869));
  xor_4  g10493(.A(new_n10869), .B(new_n10858), .Y(new_n10870));
  xor_4  g10494(.A(new_n10870), .B(new_n10855), .Y(new_n10871));
  xor_4  g10495(.A(new_n10871), .B(new_n10847), .Y(new_n10872));
  xor_4  g10496(.A(new_n10872), .B(new_n10846), .Y(new_n10873));
  xor_4  g10497(.A(new_n10873), .B(new_n10796), .Y(new_n10874));
  xor_4  g10498(.A(new_n10874), .B(new_n10706), .Y(po109));
  xor_4  g10499(.A(new_n4949), .B(new_n4948), .Y(po110));
  xor_4  g10500(.A(new_n3108), .B(new_n3107), .Y(po111));
  xor_4  g10501(.A(new_n8106), .B(new_n8105), .Y(po112));
  xor_4  g10502(.A(new_n8112), .B(new_n8110), .Y(po113));
  xor_4  g10503(.A(new_n8423), .B(new_n8421), .Y(po114));
  xor_4  g10504(.A(new_n7057), .B(new_n7055), .Y(po115));
  xor_4  g10505(.A(new_n9187), .B(new_n9186), .Y(po116));
  xor_4  g10506(.A(new_n9647), .B(new_n9646), .Y(po117));
  xor_4  g10507(.A(new_n8425), .B(new_n8414), .Y(po118));
  xor_4  g10508(.A(new_n4572), .B(new_n4570), .Y(po119));
endmodule


