module top_809698493_843330999_809698999_896665269_4392119
//module top_809698492_843330999_809698999_896665269_4392119
// module top_809698491_826291639_762447541_4392120
( n45 , n112 , n137 , n159 , n217 , n226 , n381 , n397 , n405 , 
n447 , n503 , n521 , n533 , n615 , n658 , n671 , n753 , n783 , n806 , 
n837 , n844 , n911 , n992 , n996 , n1020 , n1067 , n1094 , n1097 , n1136 , 
n1138 , n1198 , n1199 , n1209 , n1269 , n1333 , n1353 , n1357 , n1471 , n1478 , 
n1510 , n1512 , n1523 , n1564 , n1576 , n1658 , n1798 , n1835 , n1847 , n1906 , 
n1980 , n2024 , n2087 , n2096 , n2131 , n2226 , n2253 , n2278 , n2301 , n2316 , 
n2347 , n2383 , n2393 , n2425 , n2431 , n2433 , n2434 , n2464 , n2498 , n2507 , 
n2508 , n2509 , n2512 , n2515 , n2522 , n2530 , n2551 , n2558 , n2564 , n2577 , 
n2581 , n2585 , n2624 , n2679 , n2708 , n2749 , n2802 , n2818 , n2879 , n2902 , 
n3022 , n3071 , n3124 , n3146 , n3172 , n3214 , n3230 , n3272 , n3287 , n3339 , 
n3342 , n3456 , n3602 , n3616 , n3627 , n3654 , n3661 , n3677 , n3719 , n3754 , 
n3842 , n3849 , n3865 , n3932 , n3986 , n3992 , n4005 , n4086 , n4088 , n4094 , 
n4141 , n4155 , n4159 , n4187 , n4189 , n4190 , n4203 , n4226 , n4230 , n4300 , 
n4312 , n4326 , n4333 , n4370 , n4378 , n4397 , n4436 , n4499 , n4516 , n4553 , 
n4634 , n4686 , n4689 , n4722 , n4733 , n4757 , n4805 , n4817 , n4826 , n4828 , 
n4903 , n4921 , n4928 , n4938 , n4970 , n4971 , n5030 , n5034 , n5069 , n5094 , 
n5105 , n5132 , n5153 , n5191 , n5198 , n5212 , n5240 , n5257 , n5283 , n5305 , 
n5314 , n5319 , n5320 , n5331 , n5411 , n5435 , n5579 , n5641 , n5645 , n5670 , 
n5693 , n5694 , n5760 , n5767 , n5798 , n5814 , n5857 , n5860 , n5934 , n5964 , 
n6016 , n6038 , n6089 , n6126 , n6192 , n6254 , n6273 , n6294 , n6358 , n6359 , 
n6429 , n6431 , n6441 , n6445 , n6578 , n6604 , n6611 , n6645 , n6687 , n6689 , 
n6703 , n6742 , n6770 , n6776 , n6797 , n6806 , n6809 , n6822 , n6826 , n6860 , 
n6877 , n6986 , n7159 , n7160 , n7193 , n7236 , n7265 , n7270 , n7294 , n7320 , 
n7354 , n7388 , n7436 , n7456 , n7500 , n7523 , n7546 , n7568 , n7610 , n7646 , 
n7676 , n7690 , n7730 , n7733 , n7823 , n7862 , n7891 , n7946 , n7965 , n7966 , 
n7981 , n8028 , n8065 , n8100 , n8138 , n8202 , n8236 , n8276 , n8303 , n8336 , 
n8384 , n8398 , n8433 , n8476 , n8595 , n8665 , n8717 , n8759 , n8819 , n9080 , 
n9111 , n9137 , n9189 , n9195 , n9241 , n9387 , n9400 , n9457 , n9571 , n9578 , 
n9583 , n9637 , n9640 , n9706 , n9725 , n9756 , n9763 , n9767 , n9820 , n9920 , 
n9938 , n9956 , n10022 , n10174 , n10217 , n10223 , n10278 , n10327 , n10391 , n10439 , 
n10451 , n10476 , n10510 , n10545 , n10547 , n10589 , n10644 , n10678 , n10685 , n10695 , 
n10789 , n10848 , n10851 , n10898 , n10913 , n10928 , n10949 , n10965 , n10990 , n11023 , 
n11153 , n11216 , n11222 , n11257 , n11296 , n11311 , n11326 , n11407 , n11423 , n11478 , 
n11536 , n11662 , n11707 , n11728 , n11755 , n11757 , n11780 , n11791 , n11821 , n11876 , 
n11877 , n11892 , n11917 , n11919 , n11922 , n11967 , n11999 , n12000 , n12005 , n12014 , 
n12020 , n12025 , n12044 , n12069 , n12076 , n12111 , n12145 , n12221 , n12247 , n12299 , 
n12391 , n12444 , n12489 , n12511 , n12591 , n12648 , n12704 , n12705 , n12706 , n12709 , 
n12720 , n12753 , n12777 , n12807 , n12826 , n12925 , n12947 );
    input n45 , n137 , n159 , n217 , n405 , n447 , n503 , n521 , n533 , 
n615 , n753 , n783 , n806 , n996 , n1067 , n1094 , n1097 , n1198 , n1199 , 
n1209 , n1333 , n1353 , n1357 , n1471 , n1478 , n1510 , n1512 , n1564 , n1576 , 
n1798 , n1835 , n1906 , n1980 , n2024 , n2087 , n2226 , n2253 , n2278 , n2347 , 
n2393 , n2433 , n2464 , n2498 , n2507 , n2508 , n2509 , n2512 , n2515 , n2522 , 
n2530 , n2551 , n2558 , n2564 , n2577 , n2585 , n2749 , n2802 , n2879 , n3022 , 
n3146 , n3172 , n3342 , n3602 , n3616 , n3627 , n3719 , n3754 , n3842 , n3865 , 
n3932 , n3986 , n3992 , n4005 , n4086 , n4094 , n4141 , n4187 , n4189 , n4190 , 
n4203 , n4312 , n4370 , n4436 , n4499 , n4516 , n4634 , n4722 , n4805 , n4817 , 
n4826 , n4828 , n4903 , n4921 , n4928 , n4938 , n4970 , n5069 , n5105 , n5153 , 
n5198 , n5212 , n5240 , n5283 , n5305 , n5314 , n5319 , n5320 , n5331 , n5579 , 
n5645 , n5694 , n5760 , n5767 , n5798 , n5814 , n5857 , n5860 , n5964 , n6016 , 
n6038 , n6126 , n6254 , n6294 , n6358 , n6359 , n6429 , n6431 , n6441 , n6578 , 
n6604 , n6611 , n6687 , n6703 , n6770 , n6776 , n6797 , n6806 , n6826 , n6877 , 
n6986 , n7159 , n7160 , n7236 , n7265 , n7270 , n7294 , n7320 , n7354 , n7388 , 
n7436 , n7456 , n7500 , n7523 , n7546 , n7610 , n7646 , n7690 , n7730 , n7733 , 
n7823 , n7862 , n7891 , n7946 , n7965 , n8028 , n8065 , n8236 , n8276 , n8336 , 
n8384 , n8433 , n8476 , n8595 , n8665 , n8717 , n8759 , n8819 , n9080 , n9111 , 
n9189 , n9195 , n9241 , n9400 , n9457 , n9583 , n9637 , n9640 , n9725 , n9763 , 
n9920 , n9956 , n10022 , n10174 , n10217 , n10223 , n10278 , n10327 , n10391 , n10439 , 
n10451 , n10510 , n10545 , n10547 , n10644 , n10678 , n10685 , n10848 , n10898 , n10928 , 
n10965 , n10990 , n11023 , n11153 , n11222 , n11257 , n11296 , n11311 , n11407 , n11423 , 
n11478 , n11536 , n11662 , n11728 , n11757 , n11791 , n11821 , n11876 , n11877 , n11892 , 
n11917 , n11922 , n11967 , n11999 , n12000 , n12025 , n12044 , n12069 , n12145 , n12221 , 
n12247 , n12299 , n12391 , n12489 , n12511 , n12591 , n12648 , n12704 , n12705 , n12706 , 
n12709 , n12720 , n12753 , n12777 , n12826 , n12925 , n12947 ;
    output n112 , n226 , n381 , n397 , n658 , n671 , n837 , n844 , n911 , 
n992 , n1020 , n1136 , n1138 , n1269 , n1523 , n1658 , n1847 , n2096 , n2131 , 
n2301 , n2316 , n2383 , n2425 , n2431 , n2434 , n2581 , n2624 , n2679 , n2708 , 
n2818 , n2902 , n3071 , n3124 , n3214 , n3230 , n3272 , n3287 , n3339 , n3456 , 
n3654 , n3661 , n3677 , n3849 , n4088 , n4155 , n4159 , n4226 , n4230 , n4300 , 
n4326 , n4333 , n4378 , n4397 , n4553 , n4686 , n4689 , n4733 , n4757 , n4971 , 
n5030 , n5034 , n5094 , n5132 , n5191 , n5257 , n5411 , n5435 , n5641 , n5670 , 
n5693 , n5934 , n6089 , n6192 , n6273 , n6445 , n6645 , n6689 , n6742 , n6809 , 
n6822 , n6860 , n7193 , n7568 , n7676 , n7966 , n7981 , n8100 , n8138 , n8202 , 
n8303 , n8398 , n9137 , n9387 , n9571 , n9578 , n9706 , n9756 , n9767 , n9820 , 
n9938 , n10476 , n10589 , n10695 , n10789 , n10851 , n10913 , n10949 , n11216 , n11326 , 
n11707 , n11755 , n11780 , n11919 , n12005 , n12014 , n12020 , n12076 , n12111 , n12444 , 
n12807 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , 
n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , 
n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , 
n39 , n40 , n41 , n42 , n43 , n44 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
n131 , n132 , n133 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , 
n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , 
n152 , n153 , n154 , n155 , n156 , n157 , n158 , n160 , n161 , n162 , 
n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , 
n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , 
n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , 
n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , 
n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , 
n213 , n214 , n215 , n216 , n218 , n219 , n220 , n221 , n222 , n223 , 
n224 , n225 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , 
n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , 
n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , 
n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , 
n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , 
n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , 
n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , 
n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , 
n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , 
n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , 
n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , 
n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , 
n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , 
n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , 
n375 , n376 , n377 , n378 , n379 , n380 , n382 , n383 , n384 , n385 , 
n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , 
n396 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n406 , n407 , 
n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , 
n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , 
n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , 
n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n448 , 
n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , 
n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , 
n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , 
n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , 
n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , 
n499 , n500 , n501 , n502 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
n531 , n532 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , 
n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , 
n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , 
n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , 
n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , 
n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , 
n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , 
n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , 
n612 , n613 , n614 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , 
n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , 
n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , 
n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , 
n653 , n654 , n655 , n656 , n657 , n659 , n660 , n661 , n662 , n663 , 
n664 , n665 , n666 , n667 , n668 , n669 , n670 , n672 , n673 , n674 , 
n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n754 , n755 , 
n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , 
n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , 
n776 , n777 , n778 , n779 , n780 , n781 , n782 , n784 , n785 , n786 , 
n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n807 , 
n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , 
n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , 
n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n838 , 
n839 , n840 , n841 , n842 , n843 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
n991 , n993 , n994 , n995 , n997 , n998 , n999 , n1000 , n1001 , n1002 , 
n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , 
n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1021 , n1022 , n1023 , 
n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , 
n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , 
n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , 
n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , 
n1064 , n1065 , n1066 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1095 , 
n1096 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , 
n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , 
n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1137 , 
n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , 
n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , 
n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , 
n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , 
n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , 
n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1200 , 
n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1210 , n1211 , 
n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , 
n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , 
n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , 
n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , 
n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , 
n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1270 , n1271 , n1272 , 
n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , 
n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , 
n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , 
n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , 
n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , 
n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , 
n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , 
n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1354 , 
n1355 , n1356 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , 
n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , 
n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , 
n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , 
n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , 
n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , 
n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , 
n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , 
n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , 
n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , 
n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , 
n1466 , n1467 , n1468 , n1469 , n1470 , n1472 , n1473 , n1474 , n1475 , n1476 , 
n1477 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , 
n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , 
n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , 
n1508 , n1509 , n1511 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
n1561 , n1562 , n1563 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , 
n1572 , n1573 , n1574 , n1575 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , 
n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , 
n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , 
n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , 
n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , 
n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , 
n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , 
n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , 
n1653 , n1654 , n1655 , n1656 , n1657 , n1659 , n1660 , n1661 , n1662 , n1663 , 
n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , 
n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , 
n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , 
n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , 
n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , 
n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , 
n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , 
n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , 
n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , 
n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , 
n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , 
n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , 
n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , 
n1794 , n1795 , n1796 , n1797 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , 
n1846 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , 
n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , 
n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , 
n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , 
n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , 
n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1907 , 
n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , 
n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , 
n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , 
n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , 
n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , 
n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , 
n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , 
n1978 , n1979 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , 
n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , 
n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , 
n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , 
n2019 , n2020 , n2021 , n2022 , n2023 , n2025 , n2026 , n2027 , n2028 , n2029 , 
n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2088 , n2089 , n2090 , 
n2091 , n2092 , n2093 , n2094 , n2095 , n2097 , n2098 , n2099 , n2100 , n2101 , 
n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , 
n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , 
n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2132 , 
n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , 
n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , 
n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , 
n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , 
n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , 
n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , 
n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , 
n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
n2223 , n2224 , n2225 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , 
n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , 
n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2254 , 
n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , 
n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , 
n2275 , n2276 , n2277 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , 
n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , 
n2296 , n2297 , n2298 , n2299 , n2300 , n2302 , n2303 , n2304 , n2305 , n2306 , 
n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2317 , 
n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , 
n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , 
n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2348 , 
n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , 
n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , 
n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
n2379 , n2380 , n2381 , n2382 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
n2390 , n2391 , n2392 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
n2421 , n2422 , n2423 , n2424 , n2426 , n2427 , n2428 , n2429 , n2430 , n2432 , 
n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , 
n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2465 , 
n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , 
n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , 
n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , 
n2496 , n2497 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , 
n2510 , n2511 , n2513 , n2514 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , 
n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2531 , n2532 , n2533 , 
n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , 
n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2552 , n2553 , n2554 , 
n2555 , n2556 , n2557 , n2559 , n2560 , n2561 , n2562 , n2563 , n2565 , n2566 , 
n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , 
n2578 , n2579 , n2580 , n2582 , n2583 , n2584 , n2586 , n2587 , n2588 , n2589 , 
n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
n2620 , n2621 , n2622 , n2623 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2680 , n2681 , 
n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , 
n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , 
n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2709 , n2710 , n2711 , n2712 , 
n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2750 , n2751 , n2752 , n2753 , 
n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , 
n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , 
n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , 
n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , 
n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2803 , n2804 , 
n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , 
n2815 , n2816 , n2817 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , 
n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , 
n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , 
n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , 
n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , 
n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , 
n2876 , n2877 , n2878 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , 
n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , 
n2897 , n2898 , n2899 , n2900 , n2901 , n2903 , n2904 , n2905 , n2906 , n2907 , 
n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , 
n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , 
n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , 
n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , 
n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , 
n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , 
n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , 
n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , 
n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , 
n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , 
n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , 
n3018 , n3019 , n3020 , n3021 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , 
n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , 
n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , 
n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , 
n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , 
n3069 , n3070 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
n3120 , n3121 , n3122 , n3123 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
n3141 , n3142 , n3143 , n3144 , n3145 , n3147 , n3148 , n3149 , n3150 , n3151 , 
n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , 
n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , 
n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
n3213 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , 
n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3231 , n3232 , n3233 , n3234 , 
n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , 
n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3273 , n3274 , n3275 , 
n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , 
n3286 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , 
n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , 
n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , 
n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , 
n3337 , n3338 , n3340 , n3341 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , 
n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , 
n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , 
n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , 
n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , 
n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , 
n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , 
n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , 
n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , 
n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , 
n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , 
n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3457 , n3458 , n3459 , 
n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
n3600 , n3601 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
n3611 , n3612 , n3613 , n3614 , n3615 , n3617 , n3618 , n3619 , n3620 , n3621 , 
n3622 , n3623 , n3624 , n3625 , n3626 , n3628 , n3629 , n3630 , n3631 , n3632 , 
n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , 
n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , 
n3653 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3662 , n3663 , n3664 , 
n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , 
n3675 , n3676 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , 
n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , 
n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , 
n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , 
n3716 , n3717 , n3718 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3755 , n3756 , n3757 , 
n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , 
n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , 
n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , 
n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , 
n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , 
n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , 
n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , 
n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , 
n3838 , n3839 , n3840 , n3841 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , 
n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
n3860 , n3861 , n3862 , n3863 , n3864 , n3866 , n3867 , n3868 , n3869 , n3870 , 
n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
n3931 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , 
n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , 
n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , 
n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , 
n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , 
n3982 , n3983 , n3984 , n3985 , n3987 , n3988 , n3989 , n3990 , n3991 , n3993 , 
n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , 
n4004 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , 
n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , 
n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , 
n4085 , n4087 , n4089 , n4090 , n4091 , n4092 , n4093 , n4095 , n4096 , n4097 , 
n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , 
n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , 
n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , 
n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , 
n4138 , n4139 , n4140 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , 
n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4156 , n4157 , n4158 , n4160 , 
n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4188 , n4191 , n4192 , n4193 , 
n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4204 , 
n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , 
n4225 , n4227 , n4228 , n4229 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , 
n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , 
n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , 
n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , 
n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , 
n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
n4297 , n4298 , n4299 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , 
n4308 , n4309 , n4310 , n4311 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , 
n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4327 , n4328 , n4329 , 
n4330 , n4331 , n4332 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4371 , 
n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4379 , n4380 , n4381 , n4382 , 
n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , 
n4393 , n4394 , n4395 , n4396 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , 
n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , 
n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , 
n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , 
n4434 , n4435 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , 
n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , 
n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , 
n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , 
n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , 
n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , 
n4495 , n4496 , n4497 , n4498 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , 
n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , 
n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , 
n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , 
n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , 
n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4554 , n4555 , n4556 , n4557 , 
n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , 
n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , 
n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , 
n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , 
n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , 
n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , 
n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , 
n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4635 , n4636 , n4637 , n4638 , 
n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4687 , n4688 , n4690 , 
n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
n4721 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , 
n4732 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , 
n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , 
n4753 , n4754 , n4755 , n4756 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , 
n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , 
n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , 
n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , 
n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , 
n4804 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , 
n4815 , n4816 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , 
n4827 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , 
n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , 
n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , 
n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , 
n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , 
n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , 
n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , 
n4898 , n4899 , n4900 , n4901 , n4902 , n4904 , n4905 , n4906 , n4907 , n4908 , 
n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
n4919 , n4920 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4929 , n4930 , 
n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4939 , n4940 , n4941 , 
n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , 
n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , 
n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4972 , n4973 , 
n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , 
n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , 
n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , 
n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , 
n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , 
n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5031 , n5032 , n5033 , n5035 , 
n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , 
n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , 
n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , 
n5066 , n5067 , n5068 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , 
n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5095 , n5096 , n5097 , 
n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5106 , n5107 , n5108 , 
n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , 
n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , 
n5129 , n5130 , n5131 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
n5150 , n5151 , n5152 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5199 , n5200 , n5201 , n5202 , 
n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5213 , 
n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , 
n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , 
n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5241 , n5242 , n5243 , n5244 , 
n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , 
n5255 , n5256 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , 
n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , 
n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5284 , n5285 , n5286 , 
n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , 
n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5306 , n5307 , 
n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5315 , n5316 , n5317 , n5318 , 
n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , 
n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , 
n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , 
n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , 
n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , 
n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , 
n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , 
n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5412 , 
n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , 
n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , 
n5433 , n5434 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , 
n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , 
n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , 
n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , 
n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , 
n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , 
n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , 
n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , 
n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , 
n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , 
n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , 
n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , 
n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , 
n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , 
n5574 , n5575 , n5576 , n5577 , n5578 , n5580 , n5581 , n5582 , n5583 , n5584 , 
n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , 
n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , 
n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , 
n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , 
n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , 
n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5642 , n5643 , n5644 , n5646 , 
n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , 
n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , 
n5667 , n5668 , n5669 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , 
n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , 
n5688 , n5689 , n5690 , n5691 , n5692 , n5695 , n5696 , n5697 , n5698 , n5699 , 
n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5768 , n5769 , n5770 , n5771 , 
n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , 
n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , 
n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5799 , n5800 , n5801 , n5802 , 
n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , 
n5813 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , 
n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , 
n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , 
n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , 
n5854 , n5855 , n5856 , n5858 , n5859 , n5861 , n5862 , n5863 , n5864 , n5865 , 
n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , 
n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , 
n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , 
n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , 
n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , 
n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , 
n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5935 , n5936 , 
n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , 
n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , 
n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5965 , n5966 , n5967 , 
n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , 
n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , 
n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , 
n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , 
n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6017 , n6018 , 
n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6039 , 
n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6090 , 
n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
n6121 , n6122 , n6123 , n6124 , n6125 , n6127 , n6128 , n6129 , n6130 , n6131 , 
n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , 
n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , 
n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , 
n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , 
n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , 
n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , 
n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , 
n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , 
n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , 
n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , 
n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , 
n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , 
n6253 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , 
n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6274 , 
n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , 
n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6295 , 
n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , 
n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , 
n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , 
n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , 
n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , 
n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , 
n6356 , n6357 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , 
n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , 
n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , 
n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , 
n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , 
n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , 
n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , 
n6428 , n6430 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
n6440 , n6442 , n6443 , n6444 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , 
n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , 
n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , 
n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , 
n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , 
n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , 
n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , 
n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , 
n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , 
n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , 
n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , 
n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , 
n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , 
n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6579 , n6580 , n6581 , n6582 , 
n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , 
n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , 
n6603 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6612 , n6613 , n6614 , 
n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , 
n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , 
n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , 
n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , 
n6686 , n6688 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , 
n6698 , n6699 , n6700 , n6701 , n6702 , n6704 , n6705 , n6706 , n6707 , n6708 , 
n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , 
n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , 
n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , 
n6739 , n6740 , n6741 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
n6771 , n6772 , n6773 , n6774 , n6775 , n6777 , n6778 , n6779 , n6780 , n6781 , 
n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , 
n6792 , n6793 , n6794 , n6795 , n6796 , n6798 , n6799 , n6800 , n6801 , n6802 , 
n6803 , n6804 , n6805 , n6807 , n6808 , n6810 , n6811 , n6812 , n6813 , n6814 , 
n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6823 , n6824 , n6825 , 
n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , 
n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , 
n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , 
n6857 , n6858 , n6859 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , 
n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6878 , 
n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6987 , n6988 , n6989 , 
n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7161 , 
n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , 
n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , 
n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , 
n7192 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , 
n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , 
n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , 
n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , 
n7233 , n7234 , n7235 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , 
n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , 
n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , 
n7264 , n7266 , n7267 , n7268 , n7269 , n7271 , n7272 , n7273 , n7274 , n7275 , 
n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , 
n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7295 , n7296 , 
n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , 
n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , 
n7317 , n7318 , n7319 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , 
n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , 
n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , 
n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7355 , n7356 , n7357 , n7358 , 
n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7389 , 
n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7437 , n7438 , n7439 , n7440 , 
n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
n7451 , n7452 , n7453 , n7454 , n7455 , n7457 , n7458 , n7459 , n7460 , n7461 , 
n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , 
n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , 
n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , 
n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7501 , n7502 , 
n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , 
n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , 
n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , 
n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , 
n7544 , n7545 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
n7565 , n7566 , n7567 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , 
n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , 
n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , 
n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , 
n7606 , n7607 , n7608 , n7609 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , 
n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , 
n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , 
n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7647 , 
n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , 
n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , 
n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7677 , n7678 , 
n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , 
n7689 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
n7731 , n7732 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , 
n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , 
n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , 
n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , 
n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , 
n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , 
n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , 
n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , 
n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , 
n7822 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , 
n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , 
n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , 
n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7863 , 
n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , 
n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , 
n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7892 , n7893 , n7894 , 
n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , 
n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , 
n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , 
n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , 
n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , 
n7945 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , 
n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7967 , 
n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , 
n7978 , n7979 , n7980 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , 
n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , 
n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , 
n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8029 , 
n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
n8060 , n8061 , n8062 , n8063 , n8064 , n8066 , n8067 , n8068 , n8069 , n8070 , 
n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8101 , 
n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , 
n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , 
n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , 
n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8139 , n8140 , n8141 , n8142 , 
n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , 
n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , 
n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , 
n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , 
n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , 
n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8203 , 
n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , 
n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , 
n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , 
n8234 , n8235 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , 
n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , 
n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , 
n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , 
n8275 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , 
n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , 
n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8304 , n8305 , n8306 , 
n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , 
n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , 
n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8337 , 
n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , 
n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , 
n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , 
n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , 
n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8385 , n8386 , n8387 , n8388 , 
n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8399 , 
n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
n8430 , n8431 , n8432 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
n8471 , n8472 , n8473 , n8474 , n8475 , n8477 , n8478 , n8479 , n8480 , n8481 , 
n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , 
n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , 
n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , 
n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , 
n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , 
n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , 
n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , 
n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , 
n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , 
n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , 
n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , 
n8592 , n8593 , n8594 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , 
n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , 
n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , 
n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , 
n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , 
n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , 
n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , 
n8663 , n8664 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , 
n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , 
n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , 
n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , 
n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , 
n8714 , n8715 , n8716 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , 
n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , 
n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , 
n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , 
n8755 , n8756 , n8757 , n8758 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , 
n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , 
n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , 
n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , 
n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , 
n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , 
n8816 , n8817 , n8818 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , 
n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , 
n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , 
n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , 
n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , 
n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , 
n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , 
n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , 
n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , 
n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , 
n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , 
n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , 
n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , 
n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , 
n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , 
n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , 
n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , 
n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , 
n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , 
n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , 
n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , 
n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , 
n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , 
n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , 
n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , 
n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , 
n9077 , n9078 , n9079 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , 
n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , 
n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , 
n9108 , n9109 , n9110 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , 
n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9138 , n9139 , 
n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9190 , 
n9191 , n9192 , n9193 , n9194 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , 
n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , 
n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , 
n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , 
n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9242 , 
n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , 
n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , 
n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , 
n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , 
n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , 
n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , 
n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , 
n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , 
n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , 
n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , 
n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , 
n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , 
n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , 
n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , 
n9383 , n9384 , n9385 , n9386 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , 
n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9401 , n9402 , n9403 , n9404 , 
n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , 
n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , 
n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , 
n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , 
n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , 
n9455 , n9456 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , 
n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , 
n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , 
n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , 
n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , 
n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , 
n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , 
n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , 
n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , 
n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , 
n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , 
n9566 , n9567 , n9568 , n9569 , n9570 , n9572 , n9573 , n9574 , n9575 , n9576 , 
n9577 , n9579 , n9580 , n9581 , n9582 , n9584 , n9585 , n9586 , n9587 , n9588 , 
n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , 
n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , 
n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , 
n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , 
n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9638 , n9639 , 
n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
n9701 , n9702 , n9703 , n9704 , n9705 , n9707 , n9708 , n9709 , n9710 , n9711 , 
n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , 
n9722 , n9723 , n9724 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , 
n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , 
n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , 
n9753 , n9754 , n9755 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9764 , 
n9765 , n9766 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , 
n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , 
n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , 
n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , 
n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , 
n9816 , n9817 , n9818 , n9819 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
n9917 , n9918 , n9919 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , 
n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , 
n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , 
n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9957 , n9958 , n9959 , 
n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
n10020 , n10021 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
n10171 , n10172 , n10173 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , 
n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , 
n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , 
n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , 
n10212 , n10213 , n10214 , n10215 , n10216 , n10218 , n10219 , n10220 , n10221 , n10222 , 
n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , 
n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , 
n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , 
n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , 
n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , 
n10274 , n10275 , n10276 , n10277 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , 
n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , 
n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , 
n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , 
n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , 
n10325 , n10326 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , 
n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , 
n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , 
n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , 
n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , 
n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , 
n10386 , n10387 , n10388 , n10389 , n10390 , n10392 , n10393 , n10394 , n10395 , n10396 , 
n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
n10437 , n10438 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , 
n10448 , n10449 , n10450 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , 
n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , 
n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10477 , n10478 , n10479 , 
n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , 
n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , 
n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , 
n10541 , n10542 , n10543 , n10544 , n10546 , n10548 , n10549 , n10550 , n10551 , n10552 , 
n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , 
n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , 
n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , 
n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10590 , n10591 , n10592 , n10593 , 
n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , 
n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , 
n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , 
n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , 
n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , 
n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , 
n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , 
n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , 
n10675 , n10676 , n10677 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10686 , 
n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10696 , n10697 , 
n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , 
n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , 
n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , 
n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , 
n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , 
n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , 
n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , 
n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , 
n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , 
n10788 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10849 , 
n10850 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , 
n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , 
n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , 
n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10899 , n10900 , n10901 , 
n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , 
n10912 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , 
n10923 , n10924 , n10925 , n10926 , n10927 , n10929 , n10930 , n10931 , n10932 , n10933 , 
n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , 
n10944 , n10945 , n10946 , n10947 , n10948 , n10950 , n10951 , n10952 , n10953 , n10954 , 
n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , 
n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , 
n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , 
n10986 , n10987 , n10988 , n10989 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , 
n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , 
n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , 
n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11024 , n11025 , n11026 , n11027 , 
n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , 
n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , 
n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , 
n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , 
n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , 
n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , 
n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , 
n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , 
n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , 
n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , 
n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , 
n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , 
n11148 , n11149 , n11150 , n11151 , n11152 , n11154 , n11155 , n11156 , n11157 , n11158 , 
n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , 
n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , 
n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11217 , n11218 , n11219 , 
n11220 , n11221 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , 
n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11258 , n11259 , n11260 , n11261 , 
n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , 
n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , 
n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , 
n11292 , n11293 , n11294 , n11295 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , 
n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11312 , n11313 , 
n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , 
n11324 , n11325 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , 
n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , 
n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , 
n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , 
n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , 
n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , 
n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , 
n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , 
n11405 , n11406 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , 
n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11424 , n11425 , n11426 , 
n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , 
n11477 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , 
n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , 
n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , 
n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , 
n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , 
n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11537 , n11538 , 
n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
n11659 , n11660 , n11661 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11708 , n11709 , n11710 , 
n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , 
n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11729 , n11730 , n11731 , 
n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , 
n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , 
n11752 , n11753 , n11754 , n11756 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , 
n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , 
n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11781 , n11782 , n11783 , n11784 , 
n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11792 , n11793 , n11794 , n11795 , 
n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , 
n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , 
n11816 , n11817 , n11818 , n11819 , n11820 , n11822 , n11823 , n11824 , n11825 , n11826 , 
n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , 
n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , 
n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , 
n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , 
n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11878 , 
n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , 
n11889 , n11890 , n11891 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11918 , n11920 , n11921 , 
n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , 
n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , 
n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , 
n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , 
n11963 , n11964 , n11965 , n11966 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , 
n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , 
n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , 
n11994 , n11995 , n11996 , n11997 , n11998 , n12001 , n12002 , n12003 , n12004 , n12006 , 
n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12015 , n12016 , n12017 , 
n12018 , n12019 , n12021 , n12022 , n12023 , n12024 , n12026 , n12027 , n12028 , n12029 , 
n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
n12040 , n12041 , n12042 , n12043 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12070 , n12071 , 
n12072 , n12073 , n12074 , n12075 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , 
n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , 
n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , 
n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12112 , n12113 , 
n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , 
n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , 
n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , 
n12144 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , 
n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , 
n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , 
n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , 
n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , 
n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , 
n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , 
n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12222 , n12223 , n12224 , n12225 , 
n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , 
n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , 
n12246 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
n12297 , n12298 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , 
n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , 
n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , 
n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , 
n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , 
n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , 
n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , 
n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , 
n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , 
n12388 , n12389 , n12390 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , 
n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , 
n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , 
n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , 
n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , 
n12439 , n12440 , n12441 , n12442 , n12443 , n12445 , n12446 , n12447 , n12448 , n12449 , 
n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , 
n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12490 , 
n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , 
n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , 
n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , 
n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , 
n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , 
n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , 
n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , 
n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , 
n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12592 , 
n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , 
n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , 
n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , 
n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , 
n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , 
n12643 , n12644 , n12645 , n12646 , n12647 , n12649 , n12650 , n12651 , n12652 , n12653 , 
n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , 
n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , 
n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , 
n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , 
n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , 
n12707 , n12708 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , 
n12718 , n12719 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , 
n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , 
n12749 , n12750 , n12751 , n12752 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12778 , n12779 , n12780 , 
n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , 
n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , 
n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12808 , n12809 , n12810 , n12811 , 
n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , 
n12822 , n12823 , n12824 , n12825 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , 
n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , 
n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , 
n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , 
n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , 
n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , 
n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , 
n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , 
n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , 
n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , 
n12923 , n12924 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , 
n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , 
n12944 , n12945 , n12946 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , 
n12955 , n12956 , n12957 , n12958 , n12959 , n12960 ;
    and g0 ( n2141 , n2530 , n521 );
    xnor g1 ( n206 , n491 , n5906 );
    and g2 ( n3102 , n4112 , n2282 );
    or g3 ( n2523 , n12144 , n5251 );
    or g4 ( n2468 , n491 , n9006 );
    nor g5 ( n5935 , n5205 , n1662 );
    and g6 ( n12452 , n3831 , n6309 );
    or g7 ( n3584 , n9389 , n6402 );
    xnor g8 ( n12769 , n12488 , n2077 );
    xnor g9 ( n9132 , n8037 , n4937 );
    xnor g10 ( n8628 , n8093 , n65 );
    xnor g11 ( n7698 , n8387 , n966 );
    not g12 ( n490 , n5531 );
    or g13 ( n999 , n9750 , n4371 );
    nor g14 ( n5811 , n7893 , n291 );
    nor g15 ( n4271 , n3168 , n10348 );
    or g16 ( n12068 , n636 , n12735 );
    not g17 ( n2076 , n12706 );
    xnor g18 ( n10627 , n9510 , n851 );
    xnor g19 ( n8741 , n5885 , n10164 );
    or g20 ( n6963 , n9723 , n12736 );
    or g21 ( n5770 , n10925 , n11911 );
    xnor g22 ( n2237 , n6664 , n8627 );
    not g23 ( n7708 , n10979 );
    and g24 ( n8228 , n6073 , n8947 );
    xnor g25 ( n8420 , n6208 , n6269 );
    not g26 ( n1335 , n12713 );
    nor g27 ( n6572 , n1342 , n7497 );
    xnor g28 ( n12308 , n5629 , n8716 );
    and g29 ( n3369 , n12792 , n2220 );
    xnor g30 ( n3113 , n9048 , n5993 );
    xnor g31 ( n5819 , n10889 , n7455 );
    xnor g32 ( n5150 , n7321 , n2104 );
    and g33 ( n6886 , n9202 , n7379 );
    xnor g34 ( n6118 , n10013 , n9298 );
    not g35 ( n171 , n8009 );
    and g36 ( n10492 , n638 , n7227 );
    xnor g37 ( n9668 , n2213 , n1443 );
    and g38 ( n10042 , n7236 , n11876 );
    and g39 ( n12212 , n1392 , n2337 );
    or g40 ( n3581 , n11073 , n5965 );
    and g41 ( n6875 , n246 , n5633 );
    nor g42 ( n12285 , n1762 , n5238 );
    or g43 ( n2936 , n8903 , n5834 );
    xnor g44 ( n8724 , n11543 , n924 );
    or g45 ( n11838 , n989 , n1546 );
    xnor g46 ( n4629 , n11708 , n11243 );
    or g47 ( n4319 , n7130 , n2371 );
    or g48 ( n8111 , n12237 , n12535 );
    xnor g49 ( n6562 , n11596 , n5864 );
    and g50 ( n2487 , n1989 , n3600 );
    xnor g51 ( n6692 , n10970 , n11448 );
    xnor g52 ( n3458 , n2834 , n2017 );
    xnor g53 ( n10494 , n638 , n1446 );
    xnor g54 ( n2545 , n9828 , n952 );
    xnor g55 ( n9965 , n5371 , n1780 );
    nor g56 ( n8178 , n5532 , n2604 );
    or g57 ( n11147 , n11923 , n4527 );
    xnor g58 ( n1622 , n4430 , n2054 );
    or g59 ( n1082 , n11026 , n10916 );
    or g60 ( n8348 , n2099 , n1163 );
    and g61 ( n8486 , n3207 , n10957 );
    or g62 ( n1757 , n7749 , n8602 );
    or g63 ( n10124 , n4250 , n7101 );
    nor g64 ( n2478 , n3943 , n7708 );
    xnor g65 ( n1228 , n9428 , n9981 );
    xnor g66 ( n4157 , n8423 , n7315 );
    xnor g67 ( n8463 , n3767 , n8601 );
    xnor g68 ( n9317 , n2340 , n6152 );
    xor g69 ( n8303 , n5732 , n5336 );
    and g70 ( n10085 , n9122 , n4460 );
    or g71 ( n8631 , n242 , n12250 );
    nor g72 ( n10958 , n3380 , n4252 );
    or g73 ( n1579 , n1699 , n6071 );
    and g74 ( n5316 , n4358 , n10165 );
    xnor g75 ( n10473 , n9382 , n3001 );
    or g76 ( n2321 , n8428 , n2815 );
    and g77 ( n4965 , n9271 , n1866 );
    and g78 ( n3103 , n7916 , n2642 );
    not g79 ( n8152 , n5213 );
    xnor g80 ( n3034 , n8018 , n744 );
    or g81 ( n10839 , n9370 , n12328 );
    xnor g82 ( n10454 , n1661 , n6545 );
    or g83 ( n10310 , n4175 , n457 );
    or g84 ( n6142 , n1653 , n10896 );
    xnor g85 ( n4910 , n6400 , n2360 );
    not g86 ( n8690 , n7121 );
    or g87 ( n10461 , n6718 , n12120 );
    not g88 ( n11803 , n6866 );
    and g89 ( n372 , n5350 , n3540 );
    not g90 ( n9377 , n6787 );
    or g91 ( n4958 , n9561 , n11702 );
    or g92 ( n6911 , n1937 , n12816 );
    or g93 ( n8730 , n6510 , n49 );
    xnor g94 ( n2061 , n5956 , n2369 );
    xnor g95 ( n11117 , n1930 , n9047 );
    and g96 ( n2307 , n3655 , n4653 );
    nor g97 ( n12594 , n7659 , n9923 );
    xnor g98 ( n8651 , n6335 , n5728 );
    and g99 ( n7187 , n8623 , n7113 );
    not g100 ( n2050 , n8938 );
    or g101 ( n3442 , n3127 , n10419 );
    xnor g102 ( n5257 , n10357 , n5568 );
    and g103 ( n5834 , n5489 , n10173 );
    xnor g104 ( n2462 , n4717 , n12433 );
    xnor g105 ( n7483 , n3418 , n2490 );
    or g106 ( n7076 , n3218 , n3846 );
    xnor g107 ( n4520 , n1033 , n617 );
    not g108 ( n5455 , n11016 );
    or g109 ( n9277 , n12138 , n7132 );
    nor g110 ( n12377 , n11098 , n2315 );
    nor g111 ( n11028 , n1179 , n7664 );
    xnor g112 ( n1103 , n12125 , n1204 );
    and g113 ( n12342 , n11892 , n217 );
    xnor g114 ( n6480 , n2246 , n9569 );
    not g115 ( n9422 , n8937 );
    nor g116 ( n4639 , n3509 , n727 );
    nor g117 ( n221 , n5107 , n258 );
    or g118 ( n9126 , n2956 , n6653 );
    xnor g119 ( n11397 , n842 , n10764 );
    or g120 ( n1049 , n12442 , n10382 );
    not g121 ( n3740 , n6165 );
    and g122 ( n1169 , n4760 , n10105 );
    and g123 ( n12150 , n8181 , n8485 );
    not g124 ( n4048 , n11265 );
    or g125 ( n2984 , n10904 , n126 );
    or g126 ( n8290 , n1183 , n10854 );
    not g127 ( n8158 , n5745 );
    not g128 ( n6389 , n2879 );
    or g129 ( n7837 , n295 , n8415 );
    xnor g130 ( n9153 , n9388 , n6619 );
    not g131 ( n5683 , n4809 );
    or g132 ( n3724 , n12398 , n4655 );
    and g133 ( n1355 , n9512 , n5173 );
    or g134 ( n8260 , n3127 , n8524 );
    or g135 ( n12831 , n2099 , n12441 );
    xnor g136 ( n8029 , n6075 , n12581 );
    or g137 ( n7347 , n2671 , n9678 );
    nor g138 ( n8443 , n4210 , n5871 );
    or g139 ( n8006 , n1146 , n8593 );
    xnor g140 ( n12126 , n7468 , n271 );
    xnor g141 ( n7882 , n8058 , n6323 );
    xnor g142 ( n4258 , n8581 , n4231 );
    xnor g143 ( n8100 , n750 , n863 );
    or g144 ( n2201 , n6577 , n8414 );
    not g145 ( n1179 , n7009 );
    or g146 ( n9690 , n8042 , n1905 );
    and g147 ( n9775 , n7843 , n3005 );
    not g148 ( n8929 , n2945 );
    nor g149 ( n8182 , n2474 , n6830 );
    or g150 ( n1955 , n4456 , n10442 );
    or g151 ( n11129 , n5659 , n366 );
    and g152 ( n7119 , n12862 , n5595 );
    or g153 ( n661 , n6349 , n8350 );
    and g154 ( n3565 , n4744 , n171 );
    not g155 ( n3098 , n9572 );
    or g156 ( n7791 , n11923 , n9078 );
    and g157 ( n8763 , n11892 , n2749 );
    xnor g158 ( n9184 , n9621 , n1490 );
    nor g159 ( n1142 , n2600 , n12332 );
    or g160 ( n10231 , n9878 , n10854 );
    and g161 ( n6119 , n7046 , n11778 );
    and g162 ( n3993 , n1998 , n6081 );
    xnor g163 ( n9684 , n10144 , n10484 );
    or g164 ( n7261 , n10546 , n1307 );
    or g165 ( n5800 , n3757 , n10363 );
    and g166 ( n12481 , n5559 , n496 );
    xnor g167 ( n2007 , n2086 , n7547 );
    xnor g168 ( n6659 , n7359 , n8616 );
    or g169 ( n11289 , n4498 , n5497 );
    nor g170 ( n10195 , n2608 , n4615 );
    not g171 ( n1467 , n670 );
    xnor g172 ( n12265 , n11377 , n4052 );
    or g173 ( n9114 , n3096 , n6197 );
    xnor g174 ( n12106 , n887 , n8942 );
    xnor g175 ( n12785 , n9065 , n141 );
    xnor g176 ( n11886 , n4999 , n4897 );
    xnor g177 ( n2345 , n3978 , n3515 );
    or g178 ( n11694 , n7391 , n1851 );
    and g179 ( n1064 , n118 , n5957 );
    not g180 ( n11474 , n7519 );
    and g181 ( n6846 , n2125 , n9796 );
    xnor g182 ( n12160 , n5177 , n4626 );
    or g183 ( n9081 , n11026 , n9568 );
    not g184 ( n9402 , n5697 );
    not g185 ( n5261 , n9539 );
    or g186 ( n4451 , n1941 , n11820 );
    xnor g187 ( n12075 , n747 , n4069 );
    and g188 ( n1443 , n5436 , n6471 );
    not g189 ( n676 , n9677 );
    and g190 ( n7897 , n12406 , n5121 );
    and g191 ( n9592 , n6030 , n3866 );
    xnor g192 ( n6858 , n5377 , n10765 );
    nor g193 ( n1968 , n1557 , n7030 );
    xnor g194 ( n10924 , n176 , n6873 );
    xnor g195 ( n10008 , n1689 , n9950 );
    or g196 ( n1682 , n7449 , n6922 );
    or g197 ( n4784 , n9978 , n2489 );
    and g198 ( n2632 , n3992 , n8433 );
    or g199 ( n5703 , n8535 , n2410 );
    nor g200 ( n9494 , n4980 , n8875 );
    or g201 ( n9082 , n7391 , n7881 );
    or g202 ( n4696 , n7116 , n12816 );
    not g203 ( n7725 , n716 );
    and g204 ( n11913 , n1161 , n134 );
    or g205 ( n12192 , n11434 , n10153 );
    nor g206 ( n3185 , n12347 , n9480 );
    and g207 ( n1397 , n10545 , n7159 );
    xnor g208 ( n3564 , n10959 , n3879 );
    or g209 ( n8596 , n10142 , n2076 );
    or g210 ( n500 , n10657 , n11861 );
    and g211 ( n9942 , n7363 , n10684 );
    or g212 ( n3555 , n9004 , n3164 );
    xnor g213 ( n8213 , n10527 , n4227 );
    or g214 ( n2670 , n994 , n1162 );
    xnor g215 ( n1528 , n1139 , n5098 );
    and g216 ( n5190 , n11969 , n5585 );
    and g217 ( n5526 , n12391 , n2558 );
    not g218 ( n6193 , n1185 );
    and g219 ( n12583 , n5395 , n1952 );
    xnor g220 ( n10722 , n8066 , n9294 );
    xnor g221 ( n8639 , n4777 , n7475 );
    xnor g222 ( n10497 , n6177 , n10713 );
    xnor g223 ( n141 , n9073 , n4641 );
    not g224 ( n7553 , n270 );
    or g225 ( n3900 , n3562 , n10796 );
    and g226 ( n7127 , n6601 , n7223 );
    and g227 ( n5167 , n11736 , n569 );
    and g228 ( n7230 , n12675 , n11381 );
    and g229 ( n10258 , n11204 , n243 );
    xnor g230 ( n6464 , n12351 , n5804 );
    or g231 ( n4032 , n3967 , n8057 );
    or g232 ( n6740 , n3746 , n11820 );
    and g233 ( n9773 , n4966 , n5161 );
    nor g234 ( n442 , n690 , n11084 );
    xnor g235 ( n1693 , n12004 , n5033 );
    xnor g236 ( n9719 , n4012 , n1971 );
    and g237 ( n5673 , n9199 , n2302 );
    xnor g238 ( n2623 , n8863 , n7766 );
    or g239 ( n839 , n6590 , n11930 );
    not g240 ( n11893 , n9547 );
    and g241 ( n7577 , n4787 , n1889 );
    or g242 ( n3734 , n7810 , n4538 );
    or g243 ( n9652 , n6718 , n9144 );
    and g244 ( n9954 , n2995 , n10800 );
    not g245 ( n1130 , n1584 );
    or g246 ( n6681 , n5530 , n5326 );
    and g247 ( n7139 , n12803 , n11117 );
    xnor g248 ( n12032 , n11324 , n12756 );
    xnor g249 ( n639 , n2381 , n8506 );
    or g250 ( n1461 , n2456 , n6071 );
    and g251 ( n3623 , n10435 , n4895 );
    xnor g252 ( n11001 , n8123 , n6774 );
    xnor g253 ( n10036 , n9152 , n9509 );
    or g254 ( n5449 , n7906 , n9794 );
    or g255 ( n2236 , n12930 , n6947 );
    nor g256 ( n886 , n2837 , n5360 );
    or g257 ( n8020 , n4960 , n4945 );
    or g258 ( n5473 , n9373 , n12771 );
    not g259 ( n1311 , n1594 );
    and g260 ( n186 , n12705 , n3932 );
    not g261 ( n10142 , n6687 );
    or g262 ( n9203 , n11923 , n2020 );
    or g263 ( n9070 , n2056 , n10008 );
    xnor g264 ( n10747 , n5294 , n4748 );
    or g265 ( n2654 , n4579 , n1167 );
    or g266 ( n11602 , n8216 , n10480 );
    or g267 ( n9159 , n5160 , n9283 );
    xnor g268 ( n1496 , n6993 , n8633 );
    or g269 ( n5652 , n4628 , n530 );
    nor g270 ( n1005 , n11813 , n8922 );
    and g271 ( n64 , n2842 , n6424 );
    or g272 ( n10675 , n6032 , n3801 );
    not g273 ( n8405 , n6578 );
    xnor g274 ( n11788 , n11610 , n2547 );
    and g275 ( n4774 , n4972 , n2542 );
    or g276 ( n11068 , n5945 , n2232 );
    or g277 ( n8169 , n2382 , n948 );
    nor g278 ( n4396 , n5092 , n3074 );
    or g279 ( n1714 , n12610 , n7794 );
    or g280 ( n11266 , n11923 , n4875 );
    or g281 ( n11608 , n3127 , n11827 );
    not g282 ( n8210 , n8772 );
    and g283 ( n9482 , n12273 , n9256 );
    or g284 ( n6458 , n5788 , n7673 );
    xnor g285 ( n7728 , n2009 , n12921 );
    and g286 ( n5978 , n4481 , n10634 );
    not g287 ( n4176 , n6751 );
    or g288 ( n6028 , n11941 , n4793 );
    nor g289 ( n12190 , n9490 , n767 );
    nor g290 ( n1730 , n5559 , n496 );
    nor g291 ( n11371 , n6067 , n8182 );
    and g292 ( n1151 , n4275 , n9813 );
    not g293 ( n7449 , n7388 );
    xnor g294 ( n3704 , n6984 , n2543 );
    xnor g295 ( n1366 , n4714 , n1118 );
    not g296 ( n5735 , n10425 );
    xnor g297 ( n8668 , n10743 , n8721 );
    or g298 ( n8135 , n288 , n11386 );
    or g299 ( n10134 , n3829 , n10384 );
    xnor g300 ( n12158 , n1091 , n10497 );
    xnor g301 ( n7652 , n4794 , n7799 );
    or g302 ( n3389 , n4247 , n554 );
    or g303 ( n4228 , n10196 , n8643 );
    or g304 ( n1547 , n10824 , n6501 );
    not g305 ( n2262 , n10831 );
    xnor g306 ( n2825 , n5454 , n9125 );
    and g307 ( n1686 , n1261 , n2366 );
    and g308 ( n12867 , n7683 , n12954 );
    or g309 ( n10831 , n2093 , n6102 );
    and g310 ( n3359 , n9829 , n5541 );
    not g311 ( n4421 , n5207 );
    xnor g312 ( n11610 , n5784 , n10591 );
    xnor g313 ( n9902 , n8484 , n4363 );
    xnor g314 ( n5983 , n11624 , n3484 );
    or g315 ( n2045 , n8428 , n6197 );
    and g316 ( n5276 , n3627 , n6038 );
    xnor g317 ( n8357 , n6135 , n12459 );
    nor g318 ( n4122 , n12931 , n9495 );
    or g319 ( n8649 , n27 , n1050 );
    xnor g320 ( n8783 , n6467 , n11860 );
    or g321 ( n3278 , n11923 , n4864 );
    nor g322 ( n7199 , n4512 , n11170 );
    or g323 ( n10118 , n5765 , n9144 );
    nor g324 ( n2353 , n2549 , n1680 );
    nor g325 ( n2093 , n7115 , n310 );
    not g326 ( n5045 , n7464 );
    nor g327 ( n8328 , n5647 , n10263 );
    not g328 ( n2589 , n2278 );
    or g329 ( n4046 , n6072 , n891 );
    and g330 ( n12401 , n3251 , n1274 );
    xnor g331 ( n3705 , n2906 , n6699 );
    or g332 ( n1292 , n12722 , n1763 );
    and g333 ( n12759 , n3491 , n8543 );
    or g334 ( n12122 , n2099 , n9188 );
    xnor g335 ( n10981 , n5109 , n12295 );
    or g336 ( n2187 , n8229 , n1276 );
    xnor g337 ( n416 , n7504 , n224 );
    not g338 ( n12307 , n12664 );
    xnor g339 ( n2949 , n1760 , n12766 );
    not g340 ( n7022 , n4386 );
    or g341 ( n8096 , n11552 , n8830 );
    and g342 ( n2795 , n9379 , n1356 );
    or g343 ( n2663 , n7116 , n8768 );
    xnor g344 ( n9745 , n2314 , n268 );
    xnor g345 ( n2765 , n2644 , n12810 );
    or g346 ( n6843 , n7283 , n9589 );
    or g347 ( n1239 , n7243 , n2460 );
    xnor g348 ( n6803 , n8118 , n11933 );
    or g349 ( n10530 , n8583 , n9144 );
    and g350 ( n1494 , n4347 , n6375 );
    and g351 ( n1602 , n4369 , n467 );
    nor g352 ( n8141 , n4717 , n12302 );
    and g353 ( n2705 , n11328 , n6043 );
    xnor g354 ( n11482 , n7551 , n9867 );
    nor g355 ( n5091 , n8163 , n3914 );
    xnor g356 ( n12323 , n11550 , n5176 );
    xnor g357 ( n6479 , n1654 , n8571 );
    or g358 ( n2455 , n6574 , n8331 );
    or g359 ( n7550 , n10843 , n11295 );
    xnor g360 ( n2352 , n11617 , n8400 );
    not g361 ( n8505 , n2500 );
    xnor g362 ( n2119 , n10456 , n32 );
    not g363 ( n3216 , n9437 );
    or g364 ( n2113 , n4059 , n561 );
    or g365 ( n307 , n4492 , n11901 );
    and g366 ( n11355 , n9905 , n10792 );
    and g367 ( n10096 , n2687 , n7153 );
    and g368 ( n10752 , n2159 , n12822 );
    nor g369 ( n12184 , n1637 , n11325 );
    nor g370 ( n163 , n10497 , n1091 );
    xnor g371 ( n1819 , n7763 , n185 );
    or g372 ( n2988 , n12727 , n8005 );
    or g373 ( n6836 , n2217 , n1476 );
    or g374 ( n12416 , n12853 , n8109 );
    xnor g375 ( n7622 , n4137 , n4640 );
    and g376 ( n11950 , n12699 , n4113 );
    or g377 ( n10182 , n7116 , n11122 );
    or g378 ( n4842 , n9136 , n7642 );
    xnor g379 ( n3749 , n2674 , n11847 );
    xnor g380 ( n4558 , n3769 , n3070 );
    xnor g381 ( n7215 , n5887 , n11904 );
    not g382 ( n11812 , n255 );
    or g383 ( n3757 , n5765 , n1047 );
    xnor g384 ( n11320 , n9000 , n11598 );
    or g385 ( n12746 , n5355 , n4400 );
    xnor g386 ( n9672 , n11646 , n1203 );
    not g387 ( n826 , n5645 );
    nor g388 ( n2185 , n10639 , n6479 );
    not g389 ( n9950 , n4967 );
    xnor g390 ( n42 , n12508 , n2994 );
    xnor g391 ( n409 , n715 , n4000 );
    and g392 ( n6489 , n1985 , n4186 );
    xnor g393 ( n7796 , n2307 , n12902 );
    xnor g394 ( n12480 , n3541 , n11067 );
    xnor g395 ( n11720 , n817 , n9361 );
    and g396 ( n6409 , n6642 , n1893 );
    not g397 ( n7063 , n10556 );
    xnor g398 ( n10319 , n6580 , n5304 );
    xnor g399 ( n11105 , n11280 , n8825 );
    xnor g400 ( n2679 , n68 , n1876 );
    xnor g401 ( n8406 , n11983 , n1036 );
    xnor g402 ( n4978 , n4669 , n9650 );
    xnor g403 ( n2004 , n3148 , n6821 );
    xnor g404 ( n7775 , n5983 , n9347 );
    or g405 ( n260 , n10208 , n11932 );
    xnor g406 ( n1400 , n7686 , n10079 );
    and g407 ( n10621 , n41 , n1255 );
    and g408 ( n10953 , n9529 , n7950 );
    xnor g409 ( n8567 , n2432 , n213 );
    and g410 ( n9812 , n5108 , n9198 );
    or g411 ( n878 , n756 , n12428 );
    not g412 ( n3433 , n4270 );
    or g413 ( n12098 , n6373 , n4875 );
    or g414 ( n12419 , n6001 , n1152 );
    or g415 ( n584 , n4994 , n2980 );
    xnor g416 ( n534 , n6889 , n6179 );
    and g417 ( n8356 , n3627 , n11407 );
    nor g418 ( n4467 , n7684 , n12162 );
    xnor g419 ( n7743 , n2717 , n5282 );
    xnor g420 ( n8151 , n8055 , n8344 );
    not g421 ( n727 , n7528 );
    or g422 ( n724 , n3275 , n9293 );
    and g423 ( n9475 , n8753 , n5752 );
    xnor g424 ( n3448 , n3068 , n12058 );
    and g425 ( n7346 , n4716 , n7 );
    xnor g426 ( n1120 , n633 , n1221 );
    and g427 ( n1220 , n5960 , n10664 );
    or g428 ( n12316 , n994 , n9589 );
    xnor g429 ( n5113 , n9903 , n7362 );
    xnor g430 ( n5603 , n6964 , n2143 );
    and g431 ( n11455 , n5589 , n11291 );
    or g432 ( n906 , n4453 , n4706 );
    and g433 ( n9658 , n11535 , n11767 );
    or g434 ( n4061 , n10750 , n6071 );
    xnor g435 ( n8378 , n9863 , n12860 );
    or g436 ( n7033 , n921 , n8298 );
    and g437 ( n6069 , n2838 , n6164 );
    or g438 ( n1019 , n9389 , n11746 );
    and g439 ( n3815 , n10640 , n5223 );
    and g440 ( n7778 , n6358 , n217 );
    or g441 ( n545 , n333 , n487 );
    and g442 ( n8987 , n8490 , n5321 );
    and g443 ( n7813 , n8945 , n1859 );
    and g444 ( n3337 , n8158 , n5616 );
    xnor g445 ( n11399 , n6515 , n11471 );
    or g446 ( n4013 , n2045 , n11274 );
    and g447 ( n3333 , n0 , n9322 );
    or g448 ( n7378 , n4911 , n1455 );
    xnor g449 ( n425 , n75 , n1823 );
    and g450 ( n8933 , n8363 , n5806 );
    not g451 ( n8407 , n2695 );
    or g452 ( n8451 , n12924 , n1124 );
    and g453 ( n4891 , n10843 , n11295 );
    xnor g454 ( n11833 , n408 , n11082 );
    and g455 ( n813 , n7306 , n10584 );
    xnor g456 ( n10366 , n2457 , n2517 );
    or g457 ( n2667 , n2266 , n11618 );
    xnor g458 ( n5722 , n11021 , n9660 );
    or g459 ( n6945 , n8583 , n8830 );
    and g460 ( n2085 , n12299 , n8819 );
    nor g461 ( n3413 , n9709 , n2015 );
    or g462 ( n10485 , n11108 , n11637 );
    or g463 ( n779 , n10642 , n9973 );
    nor g464 ( n12774 , n11137 , n470 );
    and g465 ( n10176 , n8758 , n12630 );
    or g466 ( n523 , n2367 , n4474 );
    not g467 ( n2252 , n8447 );
    xnor g468 ( n3269 , n12210 , n12536 );
    xnor g469 ( n9535 , n1062 , n12811 );
    or g470 ( n11902 , n5466 , n4578 );
    or g471 ( n5663 , n1808 , n2210 );
    xnor g472 ( n11496 , n4742 , n8621 );
    nor g473 ( n6113 , n9298 , n10013 );
    xnor g474 ( n9436 , n6161 , n12599 );
    or g475 ( n938 , n10354 , n1502 );
    not g476 ( n6696 , n9391 );
    xnor g477 ( n4526 , n9493 , n10069 );
    or g478 ( n428 , n4121 , n11975 );
    or g479 ( n6093 , n2013 , n8542 );
    xnor g480 ( n4749 , n9079 , n6695 );
    xnor g481 ( n7024 , n1242 , n6378 );
    xnor g482 ( n12728 , n3225 , n7099 );
    or g483 ( n2814 , n11358 , n6201 );
    or g484 ( n7169 , n11416 , n2535 );
    and g485 ( n9803 , n11832 , n9681 );
    xnor g486 ( n12148 , n4703 , n11570 );
    or g487 ( n9925 , n9802 , n9220 );
    xnor g488 ( n12850 , n9368 , n809 );
    or g489 ( n2695 , n12503 , n2020 );
    nor g490 ( n10909 , n7441 , n3009 );
    xnor g491 ( n8765 , n11563 , n5192 );
    nor g492 ( n8034 , n7579 , n10073 );
    not g493 ( n3538 , n733 );
    xnor g494 ( n3101 , n5016 , n12202 );
    not g495 ( n3434 , n3443 );
    xnor g496 ( n4231 , n771 , n1829 );
    or g497 ( n12242 , n10835 , n9160 );
    or g498 ( n3793 , n3837 , n9096 );
    or g499 ( n9797 , n10835 , n10916 );
    not g500 ( n4610 , n4784 );
    or g501 ( n8264 , n5847 , n136 );
    nor g502 ( n6933 , n645 , n4043 );
    not g503 ( n1184 , n6474 );
    or g504 ( n6893 , n10874 , n1300 );
    xnor g505 ( n2764 , n11538 , n8798 );
    xnor g506 ( n12610 , n12118 , n3721 );
    xnor g507 ( n2369 , n522 , n8401 );
    or g508 ( n3050 , n10835 , n1047 );
    and g509 ( n9670 , n5384 , n12652 );
    or g510 ( n5592 , n8115 , n1106 );
    or g511 ( n2351 , n8467 , n8231 );
    or g512 ( n7266 , n11271 , n8239 );
    and g513 ( n9060 , n9119 , n1182 );
    and g514 ( n1542 , n10326 , n9618 );
    or g515 ( n10619 , n11719 , n10066 );
    not g516 ( n5902 , n6826 );
    and g517 ( n9345 , n9236 , n1559 );
    xnor g518 ( n1538 , n11605 , n3278 );
    not g519 ( n9235 , n3460 );
    nor g520 ( n1976 , n10746 , n10577 );
    and g521 ( n11124 , n3381 , n10811 );
    nor g522 ( n5218 , n11548 , n4523 );
    xnor g523 ( n11467 , n6907 , n3610 );
    xnor g524 ( n8434 , n3840 , n4151 );
    xnor g525 ( n4333 , n8792 , n6372 );
    or g526 ( n9794 , n9878 , n12535 );
    not g527 ( n8962 , n8732 );
    not g528 ( n2012 , n8790 );
    not g529 ( n3522 , n1027 );
    xnor g530 ( n1661 , n2063 , n7466 );
    or g531 ( n1445 , n8959 , n6197 );
    or g532 ( n10573 , n12237 , n3224 );
    xnor g533 ( n5617 , n12195 , n4622 );
    and g534 ( n10225 , n10336 , n11677 );
    xnor g535 ( n11469 , n1248 , n8440 );
    not g536 ( n11350 , n10914 );
    not g537 ( n10641 , n9738 );
    xnor g538 ( n6556 , n3085 , n2554 );
    or g539 ( n947 , n8152 , n11942 );
    or g540 ( n9432 , n5355 , n7703 );
    xnor g541 ( n1168 , n6413 , n12778 );
    xnor g542 ( n8107 , n9358 , n547 );
    xnor g543 ( n8956 , n7092 , n4030 );
    not g544 ( n1871 , n3978 );
    or g545 ( n10673 , n5384 , n12652 );
    not g546 ( n2221 , n1611 );
    xnor g547 ( n837 , n5483 , n5072 );
    or g548 ( n1043 , n6577 , n9741 );
    or g549 ( n7768 , n2097 , n3792 );
    nor g550 ( n1406 , n6889 , n9422 );
    and g551 ( n12290 , n9368 , n809 );
    xnor g552 ( n12928 , n11234 , n2359 );
    xnor g553 ( n4284 , n2069 , n10458 );
    not g554 ( n5851 , n3865 );
    xnor g555 ( n5772 , n8287 , n10188 );
    or g556 ( n2600 , n12119 , n12446 );
    nor g557 ( n9689 , n7070 , n10571 );
    and g558 ( n3765 , n9933 , n8729 );
    and g559 ( n8705 , n3771 , n3302 );
    or g560 ( n11299 , n2497 , n9001 );
    and g561 ( n566 , n6934 , n1377 );
    xnor g562 ( n6799 , n4926 , n2745 );
    xnor g563 ( n1038 , n7285 , n6498 );
    and g564 ( n11093 , n3766 , n11974 );
    or g565 ( n1917 , n849 , n4575 );
    and g566 ( n3814 , n3581 , n6230 );
    and g567 ( n2441 , n3236 , n3067 );
    xnor g568 ( n7696 , n3517 , n823 );
    nor g569 ( n3751 , n1252 , n9565 );
    and g570 ( n8854 , n196 , n11477 );
    nor g571 ( n5829 , n6794 , n3545 );
    or g572 ( n3652 , n6550 , n5792 );
    or g573 ( n10418 , n8071 , n7595 );
    or g574 ( n8137 , n5850 , n1347 );
    or g575 ( n4264 , n6977 , n5012 );
    not g576 ( n11031 , n11501 );
    or g577 ( n3405 , n1051 , n12816 );
    not g578 ( n11775 , n3602 );
    not g579 ( n5594 , n6087 );
    xnor g580 ( n1520 , n11112 , n5123 );
    not g581 ( n12843 , n4921 );
    xnor g582 ( n7279 , n9194 , n2480 );
    and g583 ( n1911 , n7735 , n1324 );
    nor g584 ( n4801 , n7817 , n9118 );
    and g585 ( n7096 , n10742 , n12001 );
    not g586 ( n10101 , n1515 );
    or g587 ( n3739 , n6766 , n395 );
    xnor g588 ( n3214 , n4583 , n4276 );
    not g589 ( n7326 , n12710 );
    xnor g590 ( n3301 , n7746 , n4743 );
    or g591 ( n1317 , n2217 , n9160 );
    or g592 ( n270 , n12531 , n5565 );
    or g593 ( n2395 , n5915 , n3224 );
    or g594 ( n3166 , n10142 , n4400 );
    or g595 ( n5192 , n7449 , n9521 );
    and g596 ( n6287 , n9570 , n12050 );
    or g597 ( n4849 , n4059 , n1455 );
    not g598 ( n11369 , n12632 );
    xnor g599 ( n6942 , n3985 , n5112 );
    or g600 ( n4369 , n10551 , n7988 );
    or g601 ( n8282 , n6977 , n8414 );
    and g602 ( n8459 , n9896 , n9815 );
    xnor g603 ( n3151 , n11343 , n6106 );
    or g604 ( n10632 , n9262 , n4474 );
    nor g605 ( n6602 , n10525 , n9466 );
    not g606 ( n8684 , n7143 );
    xnor g607 ( n9783 , n12142 , n12061 );
    or g608 ( n11232 , n3746 , n7395 );
    not g609 ( n6985 , n4079 );
    and g610 ( n10472 , n4202 , n9496 );
    or g611 ( n11794 , n3324 , n1509 );
    nor g612 ( n1348 , n9063 , n9580 );
    xnor g613 ( n1201 , n3584 , n4037 );
    and g614 ( n5606 , n11950 , n5127 );
    and g615 ( n3465 , n4187 , n3602 );
    nor g616 ( n2277 , n221 , n3529 );
    not g617 ( n1448 , n10904 );
    xnor g618 ( n12409 , n2912 , n4192 );
    and g619 ( n9882 , n11152 , n10482 );
    xnor g620 ( n469 , n6220 , n59 );
    xnor g621 ( n12589 , n10983 , n91 );
    or g622 ( n11505 , n10108 , n11827 );
    nor g623 ( n12407 , n5424 , n9337 );
    or g624 ( n9433 , n7221 , n6453 );
    or g625 ( n10312 , n2593 , n8497 );
    xnor g626 ( n12268 , n7386 , n8651 );
    xnor g627 ( n8606 , n3077 , n2627 );
    xnor g628 ( n3272 , n5354 , n6014 );
    xnor g629 ( n10562 , n1785 , n12143 );
    xnor g630 ( n2387 , n2637 , n8950 );
    xnor g631 ( n4771 , n6090 , n1698 );
    or g632 ( n2982 , n5089 , n10823 );
    or g633 ( n3589 , n7905 , n12431 );
    nor g634 ( n10384 , n721 , n9327 );
    xnor g635 ( n12094 , n7483 , n5297 );
    nor g636 ( n10980 , n4541 , n7995 );
    or g637 ( n10128 , n3324 , n4474 );
    or g638 ( n3541 , n10508 , n10930 );
    or g639 ( n10636 , n10199 , n7637 );
    nor g640 ( n6597 , n9446 , n9051 );
    or g641 ( n11384 , n1705 , n12251 );
    and g642 ( n11501 , n12815 , n10109 );
    xnor g643 ( n6127 , n10744 , n5913 );
    xnor g644 ( n9874 , n9145 , n12649 );
    xnor g645 ( n4887 , n9499 , n11096 );
    and g646 ( n4414 , n12069 , n1564 );
    and g647 ( n4668 , n3265 , n1454 );
    and g648 ( n323 , n12879 , n7792 );
    not g649 ( n7512 , n2640 );
    nor g650 ( n9278 , n2011 , n4899 );
    xor g651 ( n10087 , n6087 , n3134 );
    xnor g652 ( n5106 , n6168 , n4418 );
    and g653 ( n10741 , n5289 , n6166 );
    not g654 ( n12363 , n11842 );
    and g655 ( n9112 , n4013 , n9800 );
    xnor g656 ( n382 , n8140 , n10253 );
    and g657 ( n11508 , n6776 , n6703 );
    or g658 ( n3426 , n3693 , n12795 );
    nor g659 ( n9989 , n4930 , n12448 );
    not g660 ( n5098 , n6683 );
    nor g661 ( n10704 , n9278 , n12352 );
    xnor g662 ( n10681 , n10815 , n9254 );
    xnor g663 ( n5217 , n7244 , n2890 );
    not g664 ( n5541 , n11256 );
    or g665 ( n7287 , n11425 , n6025 );
    xnor g666 ( n11768 , n5846 , n12628 );
    or g667 ( n9796 , n12283 , n8333 );
    xnor g668 ( n691 , n7496 , n3436 );
    xnor g669 ( n10843 , n11533 , n12068 );
    xnor g670 ( n3367 , n2488 , n6203 );
    or g671 ( n9806 , n5809 , n12080 );
    or g672 ( n8191 , n7283 , n2076 );
    and g673 ( n4803 , n5231 , n5217 );
    xnor g674 ( n12449 , n8313 , n879 );
    or g675 ( n4238 , n10735 , n4091 );
    xnor g676 ( n3285 , n3884 , n734 );
    xnor g677 ( n8084 , n12203 , n10593 );
    and g678 ( n4034 , n3274 , n3755 );
    nor g679 ( n350 , n1065 , n4039 );
    and g680 ( n8900 , n7236 , n5760 );
    or g681 ( n8782 , n7271 , n11263 );
    nor g682 ( n2639 , n10918 , n12900 );
    and g683 ( n1561 , n5020 , n3916 );
    xnor g684 ( n5721 , n12873 , n10513 );
    and g685 ( n6384 , n8176 , n2388 );
    or g686 ( n8789 , n5575 , n11896 );
    or g687 ( n7437 , n4428 , n8797 );
    or g688 ( n1745 , n1507 , n9168 );
    or g689 ( n134 , n10521 , n1828 );
    and g690 ( n699 , n8903 , n5834 );
    or g691 ( n10822 , n3666 , n7068 );
    xnor g692 ( n12100 , n10091 , n3560 );
    xnor g693 ( n12091 , n6195 , n7571 );
    xnor g694 ( n1551 , n5284 , n12676 );
    or g695 ( n12443 , n994 , n1079 );
    not g696 ( n4052 , n10042 );
    or g697 ( n2188 , n9797 , n2900 );
    not g698 ( n8293 , n10741 );
    xnor g699 ( n1361 , n8027 , n228 );
    xnor g700 ( n5325 , n1408 , n11875 );
    not g701 ( n7395 , n10278 );
    or g702 ( n10075 , n11462 , n11148 );
    or g703 ( n976 , n2651 , n4394 );
    not g704 ( n9636 , n10080 );
    xnor g705 ( n3536 , n11568 , n8846 );
    or g706 ( n3729 , n3746 , n10919 );
    nor g707 ( n4453 , n6485 , n1187 );
    xnor g708 ( n368 , n1571 , n9891 );
    or g709 ( n10633 , n4522 , n4656 );
    or g710 ( n10774 , n5204 , n283 );
    not g711 ( n7705 , n5432 );
    xnor g712 ( n7653 , n5795 , n6118 );
    or g713 ( n7846 , n7283 , n1738 );
    xnor g714 ( n5846 , n10393 , n2540 );
    nor g715 ( n5932 , n1989 , n3600 );
    xnor g716 ( n10024 , n10457 , n7820 );
    and g717 ( n893 , n5026 , n9139 );
    or g718 ( n4466 , n8941 , n1418 );
    and g719 ( n7776 , n12658 , n6327 );
    not g720 ( n1931 , n7312 );
    not g721 ( n4811 , n10517 );
    xnor g722 ( n3546 , n11267 , n4751 );
    not g723 ( n4952 , n6203 );
    or g724 ( n11358 , n7168 , n3047 );
    and g725 ( n10742 , n9920 , n4921 );
    and g726 ( n2145 , n991 , n354 );
    and g727 ( n5376 , n1215 , n5055 );
    xnor g728 ( n8744 , n7146 , n9552 );
    not g729 ( n11377 , n2824 );
    not g730 ( n4841 , n8773 );
    nor g731 ( n9471 , n2739 , n1033 );
    xnor g732 ( n5651 , n6857 , n4544 );
    and g733 ( n3017 , n11892 , n11791 );
    not g734 ( n9534 , n11468 );
    or g735 ( n11200 , n10332 , n12934 );
    or g736 ( n6539 , n3746 , n11122 );
    or g737 ( n11394 , n5493 , n5019 );
    not g738 ( n2849 , n4 );
    or g739 ( n7674 , n9075 , n4840 );
    xnor g740 ( n512 , n4233 , n11553 );
    and g741 ( n7820 , n7453 , n2059 );
    nor g742 ( n7040 , n3651 , n3183 );
    xnor g743 ( n8535 , n4655 , n4825 );
    and g744 ( n8528 , n2427 , n1157 );
    xnor g745 ( n7636 , n1050 , n2544 );
    xnor g746 ( n10907 , n10297 , n2983 );
    or g747 ( n3618 , n12474 , n881 );
    xnor g748 ( n5317 , n7844 , n12378 );
    xnor g749 ( n6499 , n5501 , n4792 );
    xnor g750 ( n6588 , n5848 , n3913 );
    not g751 ( n4864 , n1510 );
    xnor g752 ( n454 , n10904 , n5789 );
    or g753 ( n8255 , n817 , n9817 );
    xnor g754 ( n6110 , n12867 , n3443 );
    xnor g755 ( n4128 , n8189 , n5797 );
    xnor g756 ( n1750 , n11564 , n5015 );
    xnor g757 ( n2388 , n5009 , n821 );
    and g758 ( n4105 , n3992 , n8028 );
    xnor g759 ( n8172 , n2272 , n10258 );
    nor g760 ( n6332 , n2625 , n4874 );
    or g761 ( n5522 , n11887 , n9188 );
    or g762 ( n5625 , n4780 , n10436 );
    and g763 ( n2227 , n12680 , n3783 );
    xnor g764 ( n3758 , n775 , n11071 );
    xnor g765 ( n516 , n11417 , n1314 );
    xnor g766 ( n195 , n9999 , n7478 );
    xnor g767 ( n4998 , n5942 , n11064 );
    and g768 ( n6444 , n3964 , n1334 );
    and g769 ( n80 , n6801 , n6011 );
    or g770 ( n11212 , n4628 , n5781 );
    or g771 ( n3944 , n1699 , n1932 );
    or g772 ( n9192 , n213 , n2432 );
    and g773 ( n8540 , n11422 , n10028 );
    xnor g774 ( n3019 , n10441 , n12904 );
    and g775 ( n10424 , n2901 , n2938 );
    xnor g776 ( n4689 , n595 , n10785 );
    and g777 ( n2590 , n12723 , n1130 );
    xnor g778 ( n4678 , n669 , n10559 );
    and g779 ( n5457 , n7284 , n10144 );
    not g780 ( n7803 , n12162 );
    xnor g781 ( n11708 , n3592 , n12383 );
    xnor g782 ( n1001 , n2979 , n9476 );
    xnor g783 ( n8296 , n7608 , n10632 );
    xnor g784 ( n6633 , n3600 , n8107 );
    nor g785 ( n10263 , n610 , n469 );
    xnor g786 ( n6176 , n6098 , n1845 );
    not g787 ( n5840 , n6824 );
    not g788 ( n7358 , n10947 );
    xnor g789 ( n9595 , n4886 , n5135 );
    nor g790 ( n7150 , n12875 , n6875 );
    xnor g791 ( n8060 , n11036 , n5252 );
    nor g792 ( n12612 , n9244 , n4025 );
    or g793 ( n11850 , n6738 , n11179 );
    and g794 ( n2738 , n11259 , n6119 );
    and g795 ( n5561 , n4184 , n3169 );
    not g796 ( n5704 , n5236 );
    xnor g797 ( n11412 , n6945 , n7023 );
    or g798 ( n5016 , n8026 , n10903 );
    or g799 ( n10730 , n7839 , n2815 );
    xnor g800 ( n4524 , n1366 , n8351 );
    or g801 ( n3303 , n7161 , n8765 );
    nor g802 ( n10888 , n901 , n11252 );
    or g803 ( n4459 , n11593 , n4584 );
    or g804 ( n2659 , n5915 , n826 );
    or g805 ( n9889 , n2832 , n6389 );
    xnor g806 ( n12810 , n4413 , n10803 );
    xnor g807 ( n10254 , n9649 , n12726 );
    xnor g808 ( n8804 , n2611 , n286 );
    xnor g809 ( n5956 , n3523 , n9682 );
    or g810 ( n9228 , n1051 , n2815 );
    and g811 ( n9858 , n4828 , n2498 );
    and g812 ( n3064 , n12299 , n2522 );
    and g813 ( n12737 , n7668 , n9130 );
    or g814 ( n1342 , n5765 , n8285 );
    or g815 ( n367 , n9795 , n9719 );
    xnor g816 ( n3320 , n8092 , n8358 );
    and g817 ( n2409 , n6590 , n11930 );
    nor g818 ( n9914 , n12294 , n6665 );
    or g819 ( n586 , n10838 , n3060 );
    or g820 ( n8757 , n10157 , n3606 );
    not g821 ( n5970 , n5192 );
    xnor g822 ( n10658 , n8790 , n4089 );
    not g823 ( n1857 , n1949 );
    or g824 ( n8108 , n6931 , n4506 );
    or g825 ( n9638 , n11028 , n8 );
    xnor g826 ( n7632 , n2874 , n9587 );
    and g827 ( n5774 , n222 , n9742 );
    not g828 ( n1286 , n12159 );
    or g829 ( n10462 , n6373 , n609 );
    xnor g830 ( n7428 , n7794 , n11888 );
    and g831 ( n2916 , n8011 , n4866 );
    xnor g832 ( n6285 , n2629 , n8062 );
    not g833 ( n2417 , n7043 );
    not g834 ( n4848 , n11878 );
    xnor g835 ( n1672 , n8712 , n10344 );
    or g836 ( n809 , n5765 , n9160 );
    or g837 ( n92 , n7407 , n10662 );
    not g838 ( n12034 , n6520 );
    xnor g839 ( n6760 , n10580 , n9095 );
    or g840 ( n11182 , n8428 , n7425 );
    or g841 ( n9972 , n8428 , n8414 );
    xnor g842 ( n12682 , n11694 , n4377 );
    xnor g843 ( n5165 , n12772 , n9264 );
    and g844 ( n6974 , n7826 , n12034 );
    or g845 ( n10306 , n12797 , n7876 );
    xnor g846 ( n268 , n3006 , n2446 );
    not g847 ( n2620 , n5327 );
    and g848 ( n5346 , n8844 , n302 );
    or g849 ( n3457 , n7449 , n4654 );
    or g850 ( n1360 , n9331 , n1592 );
    not g851 ( n5715 , n7024 );
    xnor g852 ( n4416 , n11995 , n8168 );
    or g853 ( n9497 , n8738 , n12771 );
    or g854 ( n12849 , n12260 , n1501 );
    or g855 ( n5214 , n4059 , n7881 );
    xnor g856 ( n9545 , n9749 , n7513 );
    or g857 ( n6817 , n4498 , n1915 );
    or g858 ( n2945 , n12237 , n8109 );
    and g859 ( n9619 , n12731 , n2110 );
    or g860 ( n8610 , n4815 , n5729 );
    xnor g861 ( n1281 , n12736 , n2764 );
    or g862 ( n3885 , n1051 , n10903 );
    xnor g863 ( n4730 , n3704 , n9396 );
    xnor g864 ( n5513 , n11259 , n6119 );
    xnor g865 ( n2092 , n4469 , n1428 );
    or g866 ( n8119 , n5809 , n5326 );
    xnor g867 ( n5026 , n11750 , n10935 );
    xnor g868 ( n2909 , n12911 , n2198 );
    and g869 ( n11734 , n7082 , n10579 );
    or g870 ( n5215 , n1675 , n344 );
    or g871 ( n6684 , n3241 , n6236 );
    xnor g872 ( n9234 , n5542 , n11232 );
    xnor g873 ( n3 , n1451 , n9676 );
    xnor g874 ( n6668 , n7035 , n11168 );
    xnor g875 ( n7975 , n12490 , n6916 );
    or g876 ( n9573 , n11172 , n6019 );
    or g877 ( n10643 , n3746 , n6169 );
    xnor g878 ( n7623 , n7526 , n4988 );
    or g879 ( n6166 , n7001 , n6401 );
    or g880 ( n3295 , n10565 , n10570 );
    or g881 ( n10926 , n4059 , n1851 );
    and g882 ( n138 , n6589 , n4049 );
    or g883 ( n6601 , n9108 , n3983 );
    xnor g884 ( n2882 , n5931 , n4617 );
    and g885 ( n8319 , n7832 , n11869 );
    and g886 ( n4897 , n4201 , n11762 );
    or g887 ( n4731 , n113 , n10259 );
    xnor g888 ( n9602 , n6368 , n12416 );
    or g889 ( n1270 , n2367 , n2020 );
    or g890 ( n7282 , n5064 , n8974 );
    not g891 ( n9448 , n7779 );
    xnor g892 ( n216 , n8035 , n6322 );
    not g893 ( n5068 , n12319 );
    xnor g894 ( n4170 , n9794 , n4954 );
    and g895 ( n10017 , n4531 , n4885 );
    not g896 ( n1394 , n6904 );
    xnor g897 ( n3738 , n459 , n8609 );
    and g898 ( n3327 , n8555 , n11568 );
    xnor g899 ( n11771 , n4366 , n10752 );
    xnor g900 ( n7677 , n10160 , n12201 );
    and g901 ( n5913 , n2289 , n12192 );
    and g902 ( n5697 , n9472 , n9462 );
    not g903 ( n6307 , n1706 );
    xnor g904 ( n761 , n6244 , n4042 );
    xnor g905 ( n1245 , n11246 , n7814 );
    xnor g906 ( n9154 , n808 , n5849 );
    or g907 ( n6011 , n8026 , n10919 );
    and g908 ( n12241 , n8759 , n3719 );
    not g909 ( n11428 , n11882 );
    and g910 ( n11465 , n3455 , n5392 );
    and g911 ( n6781 , n7626 , n7913 );
    xnor g912 ( n12893 , n745 , n10583 );
    or g913 ( n2215 , n2099 , n12686 );
    xnor g914 ( n9944 , n4860 , n1497 );
    xnor g915 ( n4489 , n5022 , n2864 );
    xnor g916 ( n7772 , n4790 , n3029 );
    nor g917 ( n5548 , n7710 , n3531 );
    xnor g918 ( n4606 , n7874 , n4992 );
    or g919 ( n4478 , n2269 , n6987 );
    and g920 ( n5318 , n3337 , n10736 );
    nor g921 ( n181 , n808 , n9934 );
    or g922 ( n1623 , n2003 , n12762 );
    and g923 ( n6866 , n7891 , n7610 );
    or g924 ( n3984 , n10142 , n10419 );
    and g925 ( n2348 , n11694 , n4377 );
    and g926 ( n5740 , n3570 , n9972 );
    and g927 ( n5194 , n3219 , n1956 );
    not g928 ( n3743 , n7236 );
    or g929 ( n10365 , n8187 , n1851 );
    not g930 ( n5383 , n6367 );
    xnor g931 ( n11512 , n12006 , n5953 );
    xnor g932 ( n3971 , n2791 , n278 );
    xnor g933 ( n10968 , n7154 , n7994 );
    not g934 ( n3622 , n7684 );
    xnor g935 ( n4194 , n4263 , n8131 );
    or g936 ( n9667 , n499 , n819 );
    or g937 ( n12205 , n1417 , n12331 );
    not g938 ( n7136 , n10965 );
    or g939 ( n7032 , n4778 , n8740 );
    or g940 ( n7853 , n5945 , n5012 );
    or g941 ( n10811 , n994 , n6389 );
    or g942 ( n1358 , n7391 , n8524 );
    xnor g943 ( n12827 , n7958 , n9537 );
    and g944 ( n10528 , n4189 , n7456 );
    nor g945 ( n4394 , n7511 , n12711 );
    and g946 ( n6794 , n6425 , n10409 );
    xnor g947 ( n6233 , n103 , n1273 );
    xnor g948 ( n5302 , n706 , n12314 );
    not g949 ( n12441 , n7546 );
    or g950 ( n2973 , n11742 , n11342 );
    and g951 ( n2147 , n11680 , n5625 );
    or g952 ( n4098 , n8687 , n795 );
    or g953 ( n5654 , n2127 , n3333 );
    xnor g954 ( n7411 , n10999 , n1976 );
    xnor g955 ( n9712 , n7925 , n5545 );
    or g956 ( n4403 , n6583 , n10700 );
    xnor g957 ( n2914 , n12053 , n4464 );
    not g958 ( n12809 , n290 );
    xnor g959 ( n10317 , n12189 , n4476 );
    or g960 ( n12837 , n1044 , n6668 );
    or g961 ( n3832 , n7640 , n1489 );
    xnor g962 ( n1652 , n7484 , n10495 );
    and g963 ( n6361 , n3171 , n8421 );
    xnor g964 ( n6223 , n8913 , n4605 );
    and g965 ( n10964 , n10692 , n1210 );
    and g966 ( n10714 , n6044 , n12521 );
    xnor g967 ( n1958 , n10012 , n5837 );
    or g968 ( n12213 , n9878 , n12735 );
    or g969 ( n5696 , n6287 , n10666 );
    nor g970 ( n9040 , n7217 , n11996 );
    and g971 ( n5329 , n1675 , n344 );
    or g972 ( n8617 , n3743 , n9280 );
    or g973 ( n3014 , n3115 , n8324 );
    xnor g974 ( n12216 , n7166 , n7878 );
    not g975 ( n9525 , n2346 );
    xnor g976 ( n1732 , n7024 , n1942 );
    xnor g977 ( n3436 , n703 , n9491 );
    and g978 ( n11554 , n11272 , n9192 );
    not g979 ( n10961 , n6010 );
    nor g980 ( n4043 , n4475 , n7910 );
    xnor g981 ( n6052 , n8122 , n1466 );
    or g982 ( n3304 , n12461 , n8212 );
    not g983 ( n11748 , n3831 );
    and g984 ( n12844 , n6901 , n12638 );
    nor g985 ( n9446 , n7693 , n3330 );
    or g986 ( n2575 , n4001 , n592 );
    nor g987 ( n6225 , n7969 , n3357 );
    and g988 ( n6143 , n11799 , n8502 );
    and g989 ( n2336 , n7236 , n10898 );
    not g990 ( n12274 , n7823 );
    xnor g991 ( n7627 , n10837 , n10968 );
    not g992 ( n6589 , n11554 );
    and g993 ( n6954 , n9875 , n7674 );
    and g994 ( n12611 , n4104 , n8504 );
    or g995 ( n411 , n5925 , n4882 );
    or g996 ( n11543 , n2357 , n12434 );
    or g997 ( n7466 , n10622 , n4876 );
    or g998 ( n4986 , n8187 , n10066 );
    xnor g999 ( n7794 , n10140 , n11763 );
    xnor g1000 ( n2276 , n4358 , n10715 );
    or g1001 ( n224 , n6977 , n2232 );
    nor g1002 ( n12392 , n7929 , n732 );
    not g1003 ( n11631 , n3006 );
    not g1004 ( n3911 , n1798 );
    or g1005 ( n1852 , n686 , n1413 );
    or g1006 ( n11364 , n9319 , n5751 );
    or g1007 ( n4186 , n1057 , n2441 );
    or g1008 ( n5550 , n9584 , n795 );
    xnor g1009 ( n7753 , n9976 , n11224 );
    nor g1010 ( n10985 , n9701 , n2799 );
    not g1011 ( n4055 , n7171 );
    xnor g1012 ( n3111 , n1515 , n6366 );
    and g1013 ( n8653 , n6461 , n3148 );
    and g1014 ( n3774 , n144 , n7137 );
    or g1015 ( n9368 , n2217 , n9144 );
    not g1016 ( n9532 , n492 );
    or g1017 ( n12660 , n5918 , n11409 );
    or g1018 ( n3688 , n2069 , n10458 );
    not g1019 ( n10653 , n4727 );
    or g1020 ( n8373 , n9218 , n10559 );
    or g1021 ( n12545 , n8583 , n7506 );
    or g1022 ( n2631 , n8794 , n2257 );
    and g1023 ( n5748 , n12935 , n9808 );
    xnor g1024 ( n4714 , n11179 , n10232 );
    or g1025 ( n2071 , n12361 , n11820 );
    or g1026 ( n10568 , n8127 , n7881 );
    or g1027 ( n10049 , n7504 , n224 );
    xnor g1028 ( n6904 , n10537 , n9412 );
    and g1029 ( n8906 , n7967 , n7261 );
    nor g1030 ( n12755 , n11029 , n11685 );
    xnor g1031 ( n12064 , n9829 , n11256 );
    xnor g1032 ( n8857 , n7980 , n6183 );
    not g1033 ( n10465 , n7209 );
    and g1034 ( n9054 , n10270 , n6999 );
    or g1035 ( n6283 , n2217 , n12120 );
    xnor g1036 ( n1227 , n10555 , n2162 );
    xnor g1037 ( n11190 , n3375 , n1986 );
    or g1038 ( n4243 , n12071 , n9046 );
    and g1039 ( n7377 , n11047 , n7479 );
    xnor g1040 ( n4363 , n6985 , n11077 );
    or g1041 ( n10860 , n9878 , n12686 );
    and g1042 ( n9862 , n6767 , n6250 );
    or g1043 ( n10646 , n8354 , n12535 );
    or g1044 ( n11589 , n8583 , n12120 );
    nor g1045 ( n11847 , n590 , n9762 );
    not g1046 ( n6144 , n11414 );
    or g1047 ( n9450 , n8583 , n4642 );
    or g1048 ( n4299 , n5690 , n1607 );
    or g1049 ( n281 , n8374 , n7235 );
    or g1050 ( n3379 , n11154 , n9405 );
    and g1051 ( n484 , n7587 , n2343 );
    or g1052 ( n1926 , n9997 , n12576 );
    and g1053 ( n7971 , n9176 , n12409 );
    not g1054 ( n4534 , n7664 );
    or g1055 ( n7243 , n3743 , n12120 );
    or g1056 ( n6538 , n12147 , n85 );
    xnor g1057 ( n12169 , n4676 , n8590 );
    not g1058 ( n9312 , n12404 );
    xnor g1059 ( n9177 , n6564 , n2896 );
    and g1060 ( n11131 , n11674 , n2726 );
    or g1061 ( n4939 , n4674 , n6513 );
    xnor g1062 ( n1059 , n8899 , n8565 );
    nor g1063 ( n1165 , n4461 , n10766 );
    and g1064 ( n9921 , n1423 , n5471 );
    and g1065 ( n10533 , n5423 , n1528 );
    nor g1066 ( n4902 , n9205 , n8089 );
    and g1067 ( n1670 , n7661 , n8724 );
    nor g1068 ( n12017 , n1874 , n8233 );
    or g1069 ( n6642 , n4782 , n4554 );
    and g1070 ( n2621 , n2448 , n3799 );
    and g1071 ( n3797 , n8025 , n3280 );
    not g1072 ( n3267 , n6548 );
    or g1073 ( n5883 , n807 , n11775 );
    or g1074 ( n4770 , n896 , n10155 );
    and g1075 ( n4659 , n12404 , n6493 );
    xnor g1076 ( n5177 , n2752 , n9236 );
    or g1077 ( n9949 , n3569 , n2707 );
    or g1078 ( n5850 , n5915 , n8655 );
    and g1079 ( n11002 , n2406 , n8073 );
    xnor g1080 ( n2644 , n5147 , n8691 );
    xnor g1081 ( n4991 , n789 , n1056 );
    or g1082 ( n9937 , n8127 , n7341 );
    or g1083 ( n9688 , n9373 , n4875 );
    not g1084 ( n5359 , n10608 );
    xnor g1085 ( n8266 , n9683 , n6559 );
    nor g1086 ( n12176 , n2192 , n11761 );
    or g1087 ( n180 , n7209 , n6807 );
    not g1088 ( n6951 , n2385 );
    xnor g1089 ( n10579 , n10416 , n4569 );
    xnor g1090 ( n11303 , n9196 , n4996 );
    xnor g1091 ( n1866 , n12473 , n10784 );
    xnor g1092 ( n12644 , n8526 , n12250 );
    or g1093 ( n12327 , n9370 , n1079 );
    nor g1094 ( n7808 , n1121 , n11510 );
    nor g1095 ( n3708 , n4045 , n1635 );
    xnor g1096 ( n12791 , n5959 , n10748 );
    xnor g1097 ( n3595 , n7939 , n11065 );
    or g1098 ( n12369 , n962 , n12771 );
    or g1099 ( n3706 , n3743 , n5914 );
    or g1100 ( n2300 , n9148 , n4417 );
    not g1101 ( n9138 , n1338 );
    nor g1102 ( n2154 , n11834 , n12355 );
    or g1103 ( n370 , n12119 , n2259 );
    nor g1104 ( n5116 , n11233 , n5078 );
    xnor g1105 ( n8058 , n11928 , n11308 );
    or g1106 ( n19 , n8990 , n1720 );
    nor g1107 ( n4274 , n6944 , n8783 );
    or g1108 ( n4124 , n2217 , n6138 );
    xnor g1109 ( n6623 , n8139 , n1473 );
    or g1110 ( n5060 , n11927 , n8157 );
    or g1111 ( n5429 , n9308 , n9562 );
    or g1112 ( n129 , n636 , n10422 );
    or g1113 ( n2870 , n2541 , n10427 );
    or g1114 ( n11356 , n191 , n8735 );
    xnor g1115 ( n1331 , n9854 , n10430 );
    or g1116 ( n11959 , n7283 , n5851 );
    xnor g1117 ( n7787 , n4304 , n3074 );
    xnor g1118 ( n8292 , n11372 , n6918 );
    and g1119 ( n5379 , n3659 , n4993 );
    xnor g1120 ( n6690 , n6579 , n9997 );
    or g1121 ( n8011 , n10157 , n9144 );
    xnor g1122 ( n6334 , n2600 , n12332 );
    or g1123 ( n9421 , n6174 , n157 );
    or g1124 ( n4693 , n3625 , n9031 );
    xnor g1125 ( n3237 , n6636 , n6991 );
    xnor g1126 ( n6735 , n10779 , n1902 );
    nor g1127 ( n7110 , n9924 , n2185 );
    and g1128 ( n3899 , n11874 , n6793 );
    or g1129 ( n7902 , n3078 , n6895 );
    xnor g1130 ( n7080 , n3171 , n2831 );
    xnor g1131 ( n10638 , n10362 , n1251 );
    and g1132 ( n6092 , n8946 , n1593 );
    not g1133 ( n9844 , n3546 );
    xnor g1134 ( n10977 , n2064 , n2267 );
    and g1135 ( n3082 , n1574 , n7706 );
    xnor g1136 ( n1487 , n6519 , n5549 );
    nor g1137 ( n3357 , n9657 , n1807 );
    or g1138 ( n6881 , n752 , n6197 );
    nor g1139 ( n212 , n1759 , n11817 );
    not g1140 ( n892 , n11166 );
    xnor g1141 ( n6483 , n4010 , n6300 );
    or g1142 ( n8920 , n3127 , n1079 );
    or g1143 ( n4630 , n807 , n7876 );
    or g1144 ( n4615 , n7449 , n4864 );
    or g1145 ( n7893 , n2832 , n3911 );
    and g1146 ( n7030 , n5027 , n10477 );
    xnor g1147 ( n10083 , n11613 , n5928 );
    nor g1148 ( n4044 , n12844 , n9183 );
    xnor g1149 ( n355 , n4492 , n6521 );
    or g1150 ( n5159 , n8631 , n1453 );
    xnor g1151 ( n7452 , n12956 , n11030 );
    xnor g1152 ( n11660 , n11959 , n8659 );
    xnor g1153 ( n11114 , n5216 , n8306 );
    nor g1154 ( n2972 , n9141 , n5149 );
    and g1155 ( n11633 , n6247 , n6973 );
    xnor g1156 ( n7719 , n8897 , n9213 );
    and g1157 ( n5943 , n7037 , n3232 );
    or g1158 ( n599 , n7057 , n3489 );
    nor g1159 ( n2703 , n7267 , n8470 );
    and g1160 ( n8864 , n2047 , n12130 );
    or g1161 ( n244 , n9754 , n4491 );
    nor g1162 ( n8352 , n330 , n2628 );
    or g1163 ( n10435 , n191 , n1915 );
    xnor g1164 ( n8893 , n7133 , n9918 );
    or g1165 ( n41 , n1937 , n995 );
    and g1166 ( n7681 , n9240 , n11264 );
    or g1167 ( n9752 , n962 , n4875 );
    xnor g1168 ( n11136 , n939 , n12824 );
    not g1169 ( n5334 , n9739 );
    or g1170 ( n6168 , n2872 , n6169 );
    nor g1171 ( n8419 , n3619 , n7592 );
    or g1172 ( n1302 , n10668 , n2397 );
    nor g1173 ( n6281 , n10352 , n8815 );
    and g1174 ( n5168 , n8120 , n4248 );
    and g1175 ( n9297 , n9807 , n6295 );
    not g1176 ( n466 , n11800 );
    not g1177 ( n7391 , n4312 );
    and g1178 ( n2784 , n11311 , n8819 );
    xnor g1179 ( n6715 , n2626 , n4041 );
    and g1180 ( n6297 , n301 , n3154 );
    nor g1181 ( n2785 , n12759 , n7915 );
    nor g1182 ( n2656 , n11784 , n9281 );
    not g1183 ( n3415 , n773 );
    and g1184 ( n6823 , n1978 , n5237 );
    xnor g1185 ( n6568 , n4859 , n8618 );
    or g1186 ( n687 , n8793 , n7736 );
    not g1187 ( n6396 , n5174 );
    xnor g1188 ( n5229 , n2337 , n9930 );
    xnor g1189 ( n8464 , n7992 , n8569 );
    and g1190 ( n4074 , n8173 , n3834 );
    and g1191 ( n3118 , n4510 , n6410 );
    xnor g1192 ( n11663 , n12659 , n6846 );
    and g1193 ( n1441 , n12647 , n11313 );
    and g1194 ( n2128 , n12069 , n1067 );
    or g1195 ( n7757 , n11347 , n6405 );
    or g1196 ( n11521 , n11443 , n11237 );
    and g1197 ( n597 , n870 , n1257 );
    xnor g1198 ( n12595 , n3954 , n8955 );
    or g1199 ( n6720 , n5455 , n7785 );
    or g1200 ( n7130 , n5915 , n9188 );
    xnor g1201 ( n445 , n12491 , n6657 );
    not g1202 ( n11282 , n9438 );
    xnor g1203 ( n4914 , n5582 , n1691 );
    and g1204 ( n8952 , n5314 , n806 );
    and g1205 ( n10020 , n1031 , n8378 );
    xnor g1206 ( n1629 , n3216 , n3120 );
    nor g1207 ( n6976 , n4057 , n176 );
    or g1208 ( n1708 , n4628 , n8655 );
    or g1209 ( n6304 , n1298 , n11303 );
    xnor g1210 ( n8412 , n1850 , n12356 );
    and g1211 ( n1469 , n1890 , n3343 );
    not g1212 ( n6595 , n3000 );
    xnor g1213 ( n11340 , n9836 , n249 );
    xnor g1214 ( n9620 , n7867 , n2545 );
    not g1215 ( n8801 , n4337 );
    xnor g1216 ( n7844 , n10884 , n3143 );
    not g1217 ( n7116 , n2226 );
    xnor g1218 ( n11385 , n7871 , n6817 );
    xnor g1219 ( n10253 , n2533 , n3099 );
    not g1220 ( n5362 , n8670 );
    and g1221 ( n5558 , n5236 , n10301 );
    xnor g1222 ( n9938 , n7323 , n7518 );
    or g1223 ( n11525 , n1432 , n4923 );
    and g1224 ( n4798 , n7774 , n7127 );
    nor g1225 ( n4461 , n3196 , n2274 );
    or g1226 ( n7309 , n5355 , n12843 );
    xnor g1227 ( n435 , n2234 , n12414 );
    xnor g1228 ( n7189 , n10980 , n4614 );
    and g1229 ( n12895 , n2476 , n9102 );
    nor g1230 ( n7481 , n9383 , n8195 );
    or g1231 ( n1995 , n686 , n5540 );
    and g1232 ( n2787 , n7550 , n12390 );
    nor g1233 ( n2655 , n8603 , n6969 );
    or g1234 ( n4103 , n11905 , n11186 );
    nor g1235 ( n1293 , n12914 , n10920 );
    or g1236 ( n5374 , n11292 , n9517 );
    and g1237 ( n10291 , n2784 , n12315 );
    nor g1238 ( n10746 , n11613 , n10710 );
    or g1239 ( n8397 , n11966 , n5091 );
    not g1240 ( n6354 , n6318 );
    not g1241 ( n2082 , n7699 );
    and g1242 ( n2533 , n1825 , n3229 );
    not g1243 ( n10331 , n9130 );
    and g1244 ( n11873 , n4057 , n176 );
    not g1245 ( n5994 , n2610 );
    or g1246 ( n4816 , n9487 , n3897 );
    or g1247 ( n12009 , n10993 , n8928 );
    or g1248 ( n12177 , n3746 , n7952 );
    xnor g1249 ( n1939 , n3646 , n1201 );
    or g1250 ( n4993 , n6577 , n11122 );
    and g1251 ( n7951 , n10139 , n3615 );
    xnor g1252 ( n5588 , n4908 , n12345 );
    or g1253 ( n7591 , n10535 , n1457 );
    and g1254 ( n3302 , n4018 , n9159 );
    xnor g1255 ( n4513 , n5241 , n245 );
    or g1256 ( n2712 , n8034 , n5868 );
    xnor g1257 ( n9442 , n9337 , n5587 );
    xnor g1258 ( n1876 , n11760 , n1301 );
    nor g1259 ( n3537 , n2684 , n9962 );
    or g1260 ( n61 , n5765 , n6138 );
    and g1261 ( n6903 , n11843 , n6440 );
    not g1262 ( n9420 , n6899 );
    or g1263 ( n144 , n12119 , n12883 );
    xnor g1264 ( n1329 , n7563 , n6609 );
    or g1265 ( n9948 , n9918 , n7575 );
    nor g1266 ( n9717 , n2885 , n11989 );
    or g1267 ( n6929 , n10835 , n5086 );
    or g1268 ( n7672 , n4911 , n12843 );
    or g1269 ( n5370 , n11887 , n1932 );
    and g1270 ( n10753 , n2606 , n11485 );
    xnor g1271 ( n5454 , n452 , n12646 );
    xnor g1272 ( n2199 , n8180 , n761 );
    xnor g1273 ( n8500 , n9974 , n3392 );
    xnor g1274 ( n479 , n679 , n9045 );
    or g1275 ( n8511 , n7944 , n2594 );
    or g1276 ( n7750 , n10729 , n8018 );
    not g1277 ( n5803 , n12081 );
    xnor g1278 ( n4879 , n9538 , n10503 );
    or g1279 ( n9479 , n8354 , n3224 );
    and g1280 ( n2808 , n3018 , n6810 );
    xnor g1281 ( n8159 , n2043 , n7717 );
    or g1282 ( n3822 , n6560 , n3741 );
    xnor g1283 ( n4491 , n4815 , n10041 );
    not g1284 ( n11926 , n7984 );
    xnor g1285 ( n10550 , n3131 , n10813 );
    or g1286 ( n4250 , n8428 , n3903 );
    nor g1287 ( n5129 , n1123 , n396 );
    not g1288 ( n1144 , n7200 );
    and g1289 ( n3511 , n11613 , n10710 );
    or g1290 ( n6582 , n319 , n1234 );
    or g1291 ( n10590 , n2217 , n9280 );
    or g1292 ( n5560 , n7380 , n1634 );
    nor g1293 ( n10251 , n11280 , n6141 );
    not g1294 ( n8302 , n1213 );
    xnor g1295 ( n4898 , n6248 , n3497 );
    and g1296 ( n4472 , n2424 , n12846 );
    or g1297 ( n9770 , n2217 , n3451 );
    not g1298 ( n4818 , n2802 );
    xor g1299 ( n4682 , n2176 , n4779 );
    xnor g1300 ( n7451 , n1598 , n8724 );
    and g1301 ( n5865 , n1272 , n8761 );
    or g1302 ( n2854 , n12853 , n3924 );
    or g1303 ( n175 , n1659 , n4714 );
    or g1304 ( n6199 , n5365 , n479 );
    xnor g1305 ( n2691 , n11499 , n1216 );
    not g1306 ( n5782 , n4233 );
    or g1307 ( n11984 , n191 , n1546 );
    not g1308 ( n12465 , n6723 );
    or g1309 ( n8194 , n9170 , n1851 );
    or g1310 ( n2616 , n7391 , n5497 );
    not g1311 ( n5185 , n1339 );
    or g1312 ( n3816 , n5828 , n5186 );
    nor g1313 ( n1340 , n8052 , n7989 );
    or g1314 ( n9881 , n4002 , n6061 );
    xnor g1315 ( n9330 , n3386 , n9746 );
    or g1316 ( n6375 , n9459 , n2193 );
    and g1317 ( n4772 , n2931 , n4376 );
    and g1318 ( n5059 , n12541 , n12031 );
    xnor g1319 ( n11479 , n4918 , n1268 );
    not g1320 ( n10935 , n11201 );
    xnor g1321 ( n3085 , n6892 , n12469 );
    xnor g1322 ( n7910 , n12522 , n12928 );
    or g1323 ( n7107 , n9836 , n8081 );
    not g1324 ( n2734 , n8702 );
    or g1325 ( n5281 , n2872 , n6455 );
    or g1326 ( n1057 , n3746 , n11775 );
    and g1327 ( n8555 , n5895 , n11374 );
    or g1328 ( n91 , n3127 , n1162 );
    xnor g1329 ( n3888 , n1590 , n1954 );
    not g1330 ( n1549 , n8562 );
    nor g1331 ( n6557 , n7481 , n9494 );
    not g1332 ( n8570 , n3219 );
    xnor g1333 ( n11982 , n8159 , n2238 );
    or g1334 ( n12512 , n2534 , n4747 );
    xnor g1335 ( n1295 , n9266 , n8711 );
    or g1336 ( n560 , n2140 , n12656 );
    and g1337 ( n4475 , n9450 , n8067 );
    xnor g1338 ( n2758 , n3943 , n4262 );
    or g1339 ( n10202 , n10157 , n4875 );
    xnor g1340 ( n8754 , n5604 , n8837 );
    xnor g1341 ( n5446 , n6697 , n12225 );
    xnor g1342 ( n7349 , n610 , n5647 );
    or g1343 ( n8926 , n9670 , n10048 );
    and g1344 ( n10389 , n8674 , n5642 );
    xnor g1345 ( n11499 , n9153 , n8379 );
    xnor g1346 ( n3209 , n4730 , n12060 );
    xnor g1347 ( n859 , n12355 , n10125 );
    xnor g1348 ( n2372 , n5267 , n9406 );
    nor g1349 ( n1666 , n2359 , n3212 );
    or g1350 ( n12182 , n7116 , n1413 );
    or g1351 ( n6527 , n191 , n11827 );
    and g1352 ( n12558 , n11134 , n401 );
    not g1353 ( n1000 , n8631 );
    xnor g1354 ( n11609 , n4905 , n620 );
    not g1355 ( n5527 , n8816 );
    nor g1356 ( n1768 , n3689 , n9332 );
    xnor g1357 ( n11447 , n4961 , n231 );
    and g1358 ( n10845 , n7862 , n1798 );
    not g1359 ( n7974 , n1241 );
    not g1360 ( n11343 , n6626 );
    or g1361 ( n10288 , n9373 , n12120 );
    or g1362 ( n3193 , n10040 , n7990 );
    xnor g1363 ( n1138 , n12461 , n12672 );
    not g1364 ( n9023 , n1648 );
    xnor g1365 ( n3319 , n10585 , n8728 );
    and g1366 ( n11936 , n7160 , n11922 );
    xnor g1367 ( n12272 , n6929 , n275 );
    xnor g1368 ( n11398 , n6836 , n332 );
    xnor g1369 ( n8571 , n2618 , n4564 );
    xnor g1370 ( n2342 , n2721 , n11628 );
    xnor g1371 ( n3268 , n12306 , n9351 );
    not g1372 ( n8183 , n3689 );
    not g1373 ( n5406 , n7096 );
    or g1374 ( n5682 , n8175 , n11003 );
    not g1375 ( n12021 , n11275 );
    or g1376 ( n3154 , n4603 , n10468 );
    xnor g1377 ( n8437 , n2677 , n9579 );
    or g1378 ( n7982 , n9301 , n2028 );
    or g1379 ( n1660 , n3127 , n6389 );
    or g1380 ( n2056 , n8870 , n3924 );
    not g1381 ( n989 , n2564 );
    and g1382 ( n2709 , n6625 , n12959 );
    and g1383 ( n6390 , n11278 , n441 );
    xnor g1384 ( n1690 , n10202 , n6271 );
    nor g1385 ( n8427 , n3538 , n682 );
    or g1386 ( n2952 , n10879 , n5497 );
    xnor g1387 ( n11918 , n3689 , n206 );
    and g1388 ( n11378 , n4314 , n9089 );
    not g1389 ( n5463 , n8990 );
    and g1390 ( n1187 , n1337 , n4054 );
    or g1391 ( n2014 , n3252 , n12542 );
    and g1392 ( n8148 , n337 , n12329 );
    not g1393 ( n463 , n1872 );
    or g1394 ( n3274 , n8737 , n5874 );
    and g1395 ( n625 , n3648 , n9664 );
    not g1396 ( n8365 , n4771 );
    and g1397 ( n9512 , n6294 , n2498 );
    xnor g1398 ( n5433 , n2599 , n1083 );
    and g1399 ( n3577 , n10463 , n5119 );
    xnor g1400 ( n12582 , n3062 , n2242 );
    xnor g1401 ( n6619 , n3007 , n8561 );
    xnor g1402 ( n322 , n5169 , n42 );
    or g1403 ( n313 , n5765 , n2020 );
    or g1404 ( n4697 , n3127 , n4242 );
    and g1405 ( n6465 , n4085 , n6000 );
    not g1406 ( n7933 , n7716 );
    xnor g1407 ( n2489 , n11530 , n8625 );
    or g1408 ( n7906 , n1699 , n8655 );
    xnor g1409 ( n4296 , n8732 , n1280 );
    not g1410 ( n12029 , n4742 );
    or g1411 ( n10749 , n7370 , n3125 );
    xnor g1412 ( n1674 , n1953 , n10276 );
    and g1413 ( n7307 , n10555 , n7791 );
    and g1414 ( n10706 , n5107 , n258 );
    or g1415 ( n10810 , n994 , n8859 );
    xnor g1416 ( n104 , n1687 , n3785 );
    and g1417 ( n10470 , n1461 , n3374 );
    and g1418 ( n937 , n10847 , n12626 );
    and g1419 ( n11345 , n1102 , n468 );
    and g1420 ( n7390 , n12518 , n10688 );
    or g1421 ( n7432 , n9834 , n7467 );
    xnor g1422 ( n10873 , n3857 , n9008 );
    xnor g1423 ( n2172 , n5144 , n5705 );
    xnor g1424 ( n9910 , n2250 , n1977 );
    or g1425 ( n3937 , n7978 , n9566 );
    xnor g1426 ( n3063 , n969 , n5046 );
    and g1427 ( n3170 , n11290 , n497 );
    and g1428 ( n4550 , n8416 , n2933 );
    or g1429 ( n8308 , n5809 , n7382 );
    or g1430 ( n12786 , n10378 , n2620 );
    and g1431 ( n908 , n279 , n2876 );
    or g1432 ( n7100 , n5575 , n7952 );
    and g1433 ( n1743 , n12881 , n10884 );
    or g1434 ( n10737 , n8354 , n5468 );
    xnor g1435 ( n2880 , n4846 , n11562 );
    xnor g1436 ( n6228 , n1029 , n8639 );
    or g1437 ( n9208 , n1746 , n2404 );
    and g1438 ( n9174 , n6078 , n2672 );
    not g1439 ( n1557 , n6834 );
    or g1440 ( n1101 , n4290 , n10113 );
    xor g1441 ( n4553 , n253 , n11227 );
    and g1442 ( n6628 , n12757 , n5057 );
    xnor g1443 ( n7863 , n7407 , n10662 );
    and g1444 ( n2950 , n5735 , n1058 );
    or g1445 ( n5166 , n2217 , n795 );
    and g1446 ( n5291 , n8276 , n9640 );
    nor g1447 ( n1758 , n908 , n6976 );
    xnor g1448 ( n8769 , n12033 , n6781 );
    xnor g1449 ( n10776 , n5333 , n257 );
    not g1450 ( n9826 , n9662 );
    or g1451 ( n2332 , n5765 , n10916 );
    and g1452 ( n7782 , n10169 , n1411 );
    xnor g1453 ( n10014 , n6486 , n1464 );
    not g1454 ( n198 , n5608 );
    xnor g1455 ( n79 , n8295 , n2862 );
    xnor g1456 ( n8197 , n352 , n8973 );
    and g1457 ( n6714 , n4635 , n12369 );
    not g1458 ( n4149 , n3775 );
    not g1459 ( n2454 , n3710 );
    or g1460 ( n12935 , n2217 , n8830 );
    and g1461 ( n11966 , n2822 , n5265 );
    or g1462 ( n1737 , n7864 , n8099 );
    nor g1463 ( n2048 , n5108 , n9198 );
    and g1464 ( n12642 , n10620 , n11302 );
    and g1465 ( n12571 , n4145 , n11459 );
    or g1466 ( n7318 , n3820 , n2020 );
    and g1467 ( n670 , n3465 , n9147 );
    xnor g1468 ( n10666 , n1899 , n9575 );
    xnor g1469 ( n7514 , n2424 , n8822 );
    or g1470 ( n7643 , n11958 , n6114 );
    xnor g1471 ( n2568 , n2130 , n2037 );
    not g1472 ( n1116 , n10423 );
    not g1473 ( n12479 , n10255 );
    and g1474 ( n9265 , n8384 , n806 );
    or g1475 ( n3131 , n2099 , n530 );
    xnor g1476 ( n5260 , n3030 , n8394 );
    or g1477 ( n8453 , n9674 , n2691 );
    nor g1478 ( n9604 , n5229 , n12653 );
    xnor g1479 ( n2233 , n8591 , n3731 );
    nor g1480 ( n1477 , n8960 , n12466 );
    or g1481 ( n8232 , n8026 , n3468 );
    or g1482 ( n1085 , n4943 , n3189 );
    and g1483 ( n49 , n3674 , n1636 );
    xnor g1484 ( n6655 , n9638 , n3555 );
    xnor g1485 ( n4988 , n4554 , n3935 );
    xnor g1486 ( n1429 , n11641 , n6333 );
    nor g1487 ( n3598 , n11353 , n10000 );
    or g1488 ( n6871 , n11285 , n6537 );
    or g1489 ( n3290 , n78 , n1934 );
    or g1490 ( n12703 , n7495 , n7424 );
    or g1491 ( n6909 , n3591 , n8082 );
    not g1492 ( n6360 , n3330 );
    and g1493 ( n7940 , n12172 , n7096 );
    not g1494 ( n967 , n2717 );
    or g1495 ( n3364 , n5171 , n4317 );
    and g1496 ( n5196 , n10103 , n411 );
    not g1497 ( n1967 , n12087 );
    or g1498 ( n6914 , n3746 , n7425 );
    and g1499 ( n3853 , n11335 , n6518 );
    xnor g1500 ( n6983 , n1206 , n5300 );
    or g1501 ( n9776 , n11433 , n2232 );
    nor g1502 ( n1779 , n2557 , n10923 );
    xnor g1503 ( n9032 , n128 , n5460 );
    not g1504 ( n2120 , n157 );
    and g1505 ( n9246 , n7388 , n12947 );
    xnor g1506 ( n5842 , n11745 , n4969 );
    and g1507 ( n6786 , n12391 , n6806 );
    or g1508 ( n7527 , n8583 , n8643 );
    xnor g1509 ( n5595 , n8568 , n9116 );
    nor g1510 ( n7980 , n12901 , n8105 );
    or g1511 ( n8691 , n11719 , n11746 );
    or g1512 ( n2801 , n4445 , n11105 );
    xnor g1513 ( n1769 , n6500 , n6593 );
    not g1514 ( n9886 , n8284 );
    or g1515 ( n5793 , n12119 , n6071 );
    nor g1516 ( n1785 , n5310 , n5912 );
    xnor g1517 ( n3419 , n6669 , n3568 );
    and g1518 ( n4079 , n11222 , n9111 );
    xnor g1519 ( n983 , n12795 , n9407 );
    not g1520 ( n11103 , n3296 );
    nor g1521 ( n2809 , n6292 , n9824 );
    xnor g1522 ( n3535 , n5273 , n108 );
    and g1523 ( n3351 , n1726 , n3718 );
    or g1524 ( n2791 , n3743 , n7921 );
    not g1525 ( n11389 , n5048 );
    or g1526 ( n290 , n10006 , n10659 );
    xnor g1527 ( n123 , n3509 , n1188 );
    and g1528 ( n2669 , n2447 , n9150 );
    xnor g1529 ( n8827 , n787 , n12944 );
    or g1530 ( n4002 , n10142 , n561 );
    or g1531 ( n9105 , n6777 , n2908 );
    xnor g1532 ( n52 , n11856 , n11998 );
    and g1533 ( n7217 , n9172 , n11949 );
    xnor g1534 ( n7174 , n2285 , n7801 );
    or g1535 ( n3194 , n8127 , n11827 );
    or g1536 ( n8382 , n7123 , n10074 );
    or g1537 ( n1161 , n4956 , n5000 );
    xnor g1538 ( n3662 , n8810 , n318 );
    or g1539 ( n2727 , n1599 , n11816 );
    and g1540 ( n8035 , n3939 , n1368 );
    xnor g1541 ( n2132 , n12457 , n3366 );
    and g1542 ( n5096 , n9000 , n5391 );
    or g1543 ( n4555 , n7760 , n11617 );
    or g1544 ( n10402 , n12237 , n10854 );
    or g1545 ( n6859 , n2808 , n11903 );
    or g1546 ( n905 , n4498 , n1079 );
    xnor g1547 ( n8874 , n99 , n11008 );
    and g1548 ( n8812 , n9900 , n5063 );
    or g1549 ( n306 , n9373 , n1509 );
    or g1550 ( n7143 , n686 , n12816 );
    or g1551 ( n6065 , n4824 , n11273 );
    or g1552 ( n6531 , n3746 , n1413 );
    not g1553 ( n9370 , n3172 );
    xnor g1554 ( n10324 , n12165 , n2720 );
    xnor g1555 ( n10421 , n3189 , n6176 );
    and g1556 ( n8784 , n10572 , n2741 );
    or g1557 ( n4929 , n5739 , n10241 );
    or g1558 ( n3428 , n3096 , n2232 );
    nor g1559 ( n5520 , n6449 , n4626 );
    xnor g1560 ( n3031 , n856 , n7324 );
    or g1561 ( n2379 , n12797 , n6169 );
    xnor g1562 ( n1795 , n9925 , n8658 );
    nor g1563 ( n12798 , n3018 , n6810 );
    or g1564 ( n7234 , n12361 , n11410 );
    not g1565 ( n12958 , n8912 );
    not g1566 ( n4782 , n9967 );
    or g1567 ( n4713 , n6718 , n609 );
    nor g1568 ( n12848 , n4741 , n4384 );
    or g1569 ( n811 , n5224 , n3851 );
    or g1570 ( n4197 , n9801 , n8528 );
    xnor g1571 ( n5480 , n12691 , n306 );
    or g1572 ( n9576 , n11552 , n8643 );
    nor g1573 ( n6649 , n6129 , n4700 );
    or g1574 ( n5687 , n8498 , n7279 );
    not g1575 ( n6000 , n10245 );
    nor g1576 ( n4823 , n1730 , n1772 );
    not g1577 ( n7816 , n3204 );
    and g1578 ( n8329 , n9690 , n5546 );
    and g1579 ( n9263 , n2107 , n5239 );
    xnor g1580 ( n2484 , n9296 , n2712 );
    and g1581 ( n8538 , n12231 , n3958 );
    or g1582 ( n2696 , n7912 , n4136 );
    or g1583 ( n12504 , n4668 , n5572 );
    or g1584 ( n5928 , n962 , n1509 );
    xnor g1585 ( n4868 , n3513 , n10491 );
    xnor g1586 ( n106 , n5947 , n5261 );
    nor g1587 ( n8346 , n6379 , n9484 );
    xnor g1588 ( n8133 , n10613 , n12740 );
    or g1589 ( n8208 , n11958 , n2754 );
    xnor g1590 ( n7873 , n219 , n10523 );
    and g1591 ( n12794 , n10770 , n4048 );
    or g1592 ( n8506 , n11747 , n4058 );
    or g1593 ( n8279 , n37 , n11316 );
    xnor g1594 ( n11016 , n4512 , n9986 );
    xnor g1595 ( n8015 , n847 , n11950 );
    and g1596 ( n8446 , n9758 , n9408 );
    or g1597 ( n8306 , n931 , n1735 );
    and g1598 ( n10635 , n9420 , n5665 );
    or g1599 ( n11882 , n11433 , n6169 );
    not g1600 ( n6212 , n10778 );
    not g1601 ( n11418 , n1776 );
    xnor g1602 ( n10189 , n8677 , n1369 );
    xnor g1603 ( n2389 , n4462 , n11363 );
    or g1604 ( n10286 , n4678 , n10234 );
    or g1605 ( n1583 , n1670 , n8700 );
    xnor g1606 ( n2586 , n9865 , n8654 );
    xnor g1607 ( n7342 , n7566 , n2932 );
    xnor g1608 ( n3182 , n5998 , n9577 );
    xnor g1609 ( n11276 , n9205 , n1069 );
    xnor g1610 ( n4192 , n8310 , n8450 );
    xnor g1611 ( n4847 , n10926 , n5600 );
    or g1612 ( n12740 , n9584 , n4474 );
    and g1613 ( n6371 , n855 , n10699 );
    xnor g1614 ( n8289 , n4484 , n1777 );
    xnor g1615 ( n6445 , n9566 , n336 );
    xnor g1616 ( n3844 , n9937 , n6224 );
    or g1617 ( n2810 , n3746 , n184 );
    nor g1618 ( n9220 , n4649 , n8075 );
    xnor g1619 ( n4963 , n8536 , n1656 );
    and g1620 ( n4584 , n8189 , n5797 );
    and g1621 ( n590 , n4434 , n1584 );
    and g1622 ( n6798 , n8757 , n3021 );
    xnor g1623 ( n4807 , n2948 , n11083 );
    or g1624 ( n683 , n12853 , n12080 );
    and g1625 ( n9171 , n7501 , n1628 );
    or g1626 ( n496 , n5915 , n530 );
    and g1627 ( n802 , n9887 , n9226 );
    and g1628 ( n5206 , n7258 , n2988 );
    xnor g1629 ( n5021 , n1552 , n2091 );
    or g1630 ( n11874 , n12691 , n6543 );
    nor g1631 ( n3040 , n1563 , n7062 );
    xnor g1632 ( n286 , n4070 , n4017 );
    nor g1633 ( n4937 , n7118 , n4093 );
    xnor g1634 ( n146 , n10243 , n9707 );
    not g1635 ( n1399 , n4581 );
    xnor g1636 ( n10218 , n1439 , n4412 );
    xnor g1637 ( n12902 , n4497 , n731 );
    or g1638 ( n3872 , n12180 , n4558 );
    not g1639 ( n5017 , n6328 );
    nor g1640 ( n11871 , n6652 , n6046 );
    or g1641 ( n6939 , n10142 , n4775 );
    or g1642 ( n8964 , n9389 , n1455 );
    or g1643 ( n6059 , n4843 , n11314 );
    xnor g1644 ( n10243 , n7640 , n2396 );
    or g1645 ( n6625 , n5530 , n8648 );
    and g1646 ( n3250 , n6797 , n12489 );
    and g1647 ( n4119 , n8656 , n3144 );
    or g1648 ( n2249 , n2703 , n850 );
    nor g1649 ( n1816 , n7501 , n1628 );
    and g1650 ( n7232 , n11400 , n7590 );
    not g1651 ( n341 , n8754 );
    xnor g1652 ( n408 , n2228 , n5286 );
    nor g1653 ( n968 , n10795 , n12909 );
    or g1654 ( n12557 , n10835 , n8745 );
    xnor g1655 ( n12765 , n11140 , n7163 );
    and g1656 ( n7173 , n11445 , n247 );
    xnor g1657 ( n755 , n9674 , n2691 );
    and g1658 ( n12502 , n9341 , n8154 );
    and g1659 ( n12688 , n2693 , n11525 );
    or g1660 ( n1784 , n6373 , n4474 );
    xnor g1661 ( n5707 , n8372 , n1480 );
    or g1662 ( n5841 , n6977 , n7425 );
    xnor g1663 ( n5807 , n1088 , n1479 );
    xnor g1664 ( n2360 , n1398 , n2338 );
    and g1665 ( n5598 , n4022 , n9318 );
    or g1666 ( n3093 , n9389 , n4400 );
    not g1667 ( n10183 , n8743 );
    and g1668 ( n8272 , n5179 , n8417 );
    xnor g1669 ( n6994 , n3368 , n1326 );
    not g1670 ( n12555 , n10493 );
    or g1671 ( n9821 , n12910 , n5296 );
    and g1672 ( n1285 , n928 , n6381 );
    and g1673 ( n85 , n7895 , n89 );
    not g1674 ( n6764 , n9872 );
    not g1675 ( n5092 , n4304 );
    xnor g1676 ( n3683 , n589 , n12321 );
    or g1677 ( n8711 , n5915 , n5468 );
    nor g1678 ( n5138 , n10070 , n7997 );
    or g1679 ( n10412 , n8894 , n10256 );
    xnor g1680 ( n4023 , n11429 , n9761 );
    and g1681 ( n12770 , n3970 , n1364 );
    xnor g1682 ( n650 , n12601 , n4149 );
    and g1683 ( n7091 , n1305 , n1928 );
    or g1684 ( n885 , n2099 , n12124 );
    not g1685 ( n12451 , n10448 );
    and g1686 ( n6173 , n2711 , n2807 );
    xnor g1687 ( n6192 , n7079 , n9911 );
    nor g1688 ( n8001 , n11741 , n1447 );
    not g1689 ( n12613 , n9419 );
    not g1690 ( n12942 , n2828 );
    and g1691 ( n10941 , n6618 , n12588 );
    nor g1692 ( n2710 , n392 , n9940 );
    and g1693 ( n1216 , n12197 , n8637 );
    and g1694 ( n10397 , n8896 , n4710 );
    and g1695 ( n6349 , n10338 , n6123 );
    xnor g1696 ( n8542 , n4268 , n5586 );
    and g1697 ( n5950 , n9074 , n972 );
    nor g1698 ( n11606 , n3336 , n3752 );
    and g1699 ( n11706 , n12694 , n7386 );
    nor g1700 ( n11865 , n7146 , n7691 );
    xnor g1701 ( n5539 , n9034 , n11359 );
    nor g1702 ( n12016 , n7819 , n7339 );
    or g1703 ( n12814 , n8118 , n9965 );
    or g1704 ( n11438 , n111 , n4618 );
    not g1705 ( n12546 , n6556 );
    xnor g1706 ( n12295 , n6746 , n3119 );
    not g1707 ( n5960 , n11345 );
    or g1708 ( n4763 , n10339 , n8740 );
    not g1709 ( n11376 , n6262 );
    xnor g1710 ( n11086 , n9016 , n10026 );
    xnor g1711 ( n9162 , n8268 , n10669 );
    xnor g1712 ( n7257 , n11415 , n12606 );
    not g1713 ( n5862 , n9380 );
    nor g1714 ( n5877 , n7620 , n1724 );
    xnor g1715 ( n8625 , n2400 , n2705 );
    nor g1716 ( n8007 , n10403 , n6870 );
    or g1717 ( n10374 , n5355 , n11430 );
    nor g1718 ( n4876 , n6406 , n3542 );
    and g1719 ( n312 , n2762 , n5782 );
    xnor g1720 ( n3543 , n6187 , n7403 );
    nor g1721 ( n12833 , n6390 , n8238 );
    and g1722 ( n8507 , n1396 , n10946 );
    or g1723 ( n7223 , n10147 , n12838 );
    and g1724 ( n6006 , n9079 , n6414 );
    xnor g1725 ( n8917 , n2957 , n3671 );
    or g1726 ( n5058 , n11043 , n9721 );
    not g1727 ( n6878 , n11749 );
    and g1728 ( n6998 , n678 , n1703 );
    xnor g1729 ( n3423 , n4346 , n1308 );
    xnor g1730 ( n8681 , n10036 , n3526 );
    xnor g1731 ( n11172 , n7229 , n10749 );
    not g1732 ( n5426 , n1373 );
    or g1733 ( n12400 , n249 , n11480 );
    xnor g1734 ( n12008 , n6081 , n12609 );
    xnor g1735 ( n7463 , n9581 , n10924 );
    xnor g1736 ( n887 , n12258 , n4705 );
    or g1737 ( n5348 , n9373 , n28 );
    and g1738 ( n12623 , n5303 , n3393 );
    or g1739 ( n4075 , n807 , n2815 );
    not g1740 ( n12397 , n3895 );
    xnor g1741 ( n5220 , n229 , n11915 );
    or g1742 ( n1433 , n1941 , n11896 );
    or g1743 ( n10045 , n2459 , n4594 );
    and g1744 ( n7081 , n5677 , n11125 );
    xnor g1745 ( n3863 , n6237 , n12917 );
    xnor g1746 ( n3315 , n12308 , n227 );
    xnor g1747 ( n11515 , n8999 , n11371 );
    xnor g1748 ( n9553 , n11724 , n9919 );
    and g1749 ( n3510 , n2602 , n4014 );
    nor g1750 ( n11979 , n5277 , n7517 );
    xnor g1751 ( n5613 , n4700 , n6129 );
    and g1752 ( n10404 , n3326 , n2364 );
    xnor g1753 ( n11337 , n7401 , n6412 );
    xnor g1754 ( n5135 , n4247 , n554 );
    or g1755 ( n2599 , n5575 , n11410 );
    xnor g1756 ( n3752 , n1859 , n12339 );
    xnor g1757 ( n6748 , n1878 , n10861 );
    or g1758 ( n12873 , n7449 , n6138 );
    xnor g1759 ( n2708 , n7749 , n3281 );
    and g1760 ( n12056 , n4602 , n2676 );
    or g1761 ( n11801 , n11026 , n4875 );
    xnor g1762 ( n2532 , n1722 , n1055 );
    or g1763 ( n773 , n11389 , n1159 );
    not g1764 ( n9302 , n7177 );
    xnor g1765 ( n460 , n1339 , n6299 );
    nor g1766 ( n4025 , n6569 , n12796 );
    or g1767 ( n4 , n270 , n11231 );
    or g1768 ( n8966 , n6031 , n3787 );
    xnor g1769 ( n6438 , n7564 , n8019 );
    or g1770 ( n7544 , n1966 , n7784 );
    xnor g1771 ( n7262 , n1672 , n2553 );
    xnor g1772 ( n3942 , n2345 , n8444 );
    xnor g1773 ( n3173 , n2555 , n12042 );
    or g1774 ( n204 , n4777 , n7475 );
    not g1775 ( n7367 , n3604 );
    or g1776 ( n2597 , n7688 , n11465 );
    not g1777 ( n10582 , n1151 );
    or g1778 ( n1099 , n763 , n5976 );
    not g1779 ( n5057 , n12118 );
    not g1780 ( n4692 , n1687 );
    nor g1781 ( n1891 , n3048 , n5978 );
    xnor g1782 ( n6791 , n2854 , n7701 );
    xnor g1783 ( n7821 , n292 , n2428 );
    or g1784 ( n11381 , n8438 , n12190 );
    not g1785 ( n11011 , n6209 );
    xnor g1786 ( n6497 , n1348 , n10372 );
    not g1787 ( n4599 , n8963 );
    and g1788 ( n784 , n8481 , n1048 );
    and g1789 ( n9579 , n8572 , n11579 );
    or g1790 ( n11534 , n3558 , n1927 );
    or g1791 ( n3260 , n989 , n1162 );
    not g1792 ( n12888 , n39 );
    not g1793 ( n378 , n10155 );
    nor g1794 ( n9168 , n10061 , n10316 );
    not g1795 ( n9417 , n10362 );
    xnor g1796 ( n9994 , n3620 , n5718 );
    xnor g1797 ( n4733 , n12019 , n8661 );
    xnor g1798 ( n10605 , n12464 , n2122 );
    and g1799 ( n1582 , n1871 , n3515 );
    xnor g1800 ( n5504 , n495 , n1189 );
    or g1801 ( n2840 , n5414 , n10759 );
    not g1802 ( n109 , n5517 );
    xnor g1803 ( n4523 , n4514 , n7677 );
    nor g1804 ( n2770 , n2842 , n6424 );
    xnor g1805 ( n9045 , n5328 , n2683 );
    or g1806 ( n695 , n2217 , n4864 );
    not g1807 ( n9389 , n4189 );
    and g1808 ( n12022 , n12960 , n10487 );
    and g1809 ( n542 , n725 , n8146 );
    or g1810 ( n3569 , n5765 , n28 );
    xnor g1811 ( n4341 , n10180 , n4234 );
    and g1812 ( n5046 , n7439 , n5891 );
    xnor g1813 ( n12600 , n10226 , n9680 );
    and g1814 ( n6861 , n607 , n419 );
    xnor g1815 ( n5435 , n1385 , n4009 );
    xnor g1816 ( n4213 , n588 , n156 );
    not g1817 ( n3048 , n37 );
    xnor g1818 ( n314 , n8789 , n1733 );
    or g1819 ( n11468 , n6718 , n4642 );
    not g1820 ( n9147 , n7131 );
    not g1821 ( n11611 , n1865 );
    not g1822 ( n7786 , n1264 );
    xnor g1823 ( n179 , n5023 , n10401 );
    and g1824 ( n7920 , n11220 , n7829 );
    nor g1825 ( n11786 , n3879 , n10499 );
    and g1826 ( n9014 , n2479 , n2317 );
    not g1827 ( n4587 , n7642 );
    or g1828 ( n11884 , n4565 , n1281 );
    not g1829 ( n11191 , n2861 );
    or g1830 ( n5757 , n9370 , n510 );
    and g1831 ( n9817 , n24 , n7334 );
    nor g1832 ( n9769 , n8232 , n7679 );
    xnor g1833 ( n6326 , n6233 , n11513 );
    xnor g1834 ( n2273 , n5423 , n9921 );
    or g1835 ( n11930 , n9370 , n11746 );
    not g1836 ( n10966 , n2311 );
    not g1837 ( n5339 , n7775 );
    xnor g1838 ( n1650 , n7864 , n8099 );
    or g1839 ( n3310 , n7116 , n11775 );
    or g1840 ( n7393 , n5530 , n12883 );
    xnor g1841 ( n8863 , n6694 , n11733 );
    nor g1842 ( n11639 , n10876 , n10982 );
    and g1843 ( n5884 , n5679 , n2963 );
    not g1844 ( n4164 , n4920 );
    xnor g1845 ( n12779 , n2903 , n10734 );
    or g1846 ( n6534 , n8026 , n3903 );
    xnor g1847 ( n6392 , n10341 , n6357 );
    xnor g1848 ( n4422 , n5090 , n1993 );
    xnor g1849 ( n9453 , n12658 , n8392 );
    or g1850 ( n10453 , n2832 , n1455 );
    nor g1851 ( n3645 , n4580 , n7561 );
    and g1852 ( n9348 , n7028 , n898 );
    xnor g1853 ( n9911 , n3811 , n7135 );
    not g1854 ( n6114 , n7730 );
    and g1855 ( n6474 , n9052 , n2716 );
    or g1856 ( n2163 , n4343 , n6513 );
    and g1857 ( n2429 , n4605 , n1678 );
    or g1858 ( n6900 , n8428 , n7395 );
    xnor g1859 ( n2205 , n1341 , n3362 );
    xnor g1860 ( n2778 , n2045 , n11274 );
    or g1861 ( n7284 , n2456 , n8655 );
    not g1862 ( n7767 , n4529 );
    xnor g1863 ( n12783 , n12091 , n12682 );
    xnor g1864 ( n6322 , n5149 , n6035 );
    not g1865 ( n4875 , n4086 );
    and g1866 ( n6430 , n7834 , n8364 );
    xnor g1867 ( n5235 , n7121 , n8944 );
    or g1868 ( n2036 , n5915 , n3924 );
    or g1869 ( n688 , n1051 , n995 );
    not g1870 ( n6485 , n9054 );
    and g1871 ( n4068 , n9027 , n1588 );
    or g1872 ( n1726 , n10142 , n1851 );
    xnor g1873 ( n3238 , n12563 , n9703 );
    xnor g1874 ( n4429 , n1411 , n1925 );
    xnor g1875 ( n12042 , n12035 , n6063 );
    and g1876 ( n6551 , n8690 , n3904 );
    xnor g1877 ( n4942 , n8219 , n6815 );
    or g1878 ( n12513 , n7449 , n609 );
    xnor g1879 ( n909 , n4525 , n11382 );
    and g1880 ( n11353 , n1025 , n4933 );
    or g1881 ( n9216 , n15 , n5218 );
    xnor g1882 ( n11298 , n3665 , n9355 );
    xnor g1883 ( n5870 , n12571 , n619 );
    xnor g1884 ( n9020 , n1583 , n4473 );
    or g1885 ( n2305 , n752 , n5540 );
    xnor g1886 ( n5624 , n940 , n9984 );
    or g1887 ( n11680 , n1043 , n11532 );
    nor g1888 ( n1530 , n1754 , n2291 );
    and g1889 ( n7656 , n11576 , n1712 );
    xnor g1890 ( n9711 , n8331 , n5351 );
    and g1891 ( n5459 , n12497 , n7033 );
    xnor g1892 ( n4984 , n2610 , n9541 );
    or g1893 ( n7303 , n2456 , n4913 );
    or g1894 ( n7964 , n2136 , n10652 );
    nor g1895 ( n11718 , n7448 , n3231 );
    not g1896 ( n8257 , n12571 );
    xnor g1897 ( n5308 , n2447 , n2313 );
    and g1898 ( n9996 , n5680 , n4883 );
    xnor g1899 ( n9868 , n7487 , n8251 );
    and g1900 ( n6298 , n9564 , n706 );
    or g1901 ( n4980 , n10339 , n6513 );
    xnor g1902 ( n10708 , n9245 , n8383 );
    and g1903 ( n12231 , n3989 , n5970 );
    or g1904 ( n10934 , n5765 , n9280 );
    or g1905 ( n7599 , n8738 , n4654 );
    or g1906 ( n7271 , n3743 , n9078 );
    and g1907 ( n10900 , n12142 , n4458 );
    or g1908 ( n6814 , n5355 , n1738 );
    not g1909 ( n1539 , n2087 );
    or g1910 ( n11709 , n6863 , n4427 );
    or g1911 ( n6219 , n2376 , n3679 );
    or g1912 ( n2630 , n12748 , n1336 );
    or g1913 ( n4992 , n9389 , n5497 );
    xnor g1914 ( n267 , n956 , n8680 );
    and g1915 ( n3176 , n5738 , n9642 );
    and g1916 ( n1821 , n7562 , n12889 );
    xnor g1917 ( n8776 , n8975 , n1619 );
    and g1918 ( n12425 , n7713 , n4012 );
    and g1919 ( n6506 , n5689 , n10134 );
    xnor g1920 ( n11380 , n7920 , n8715 );
    not g1921 ( n4411 , n1723 );
    or g1922 ( n266 , n2865 , n1942 );
    nor g1923 ( n3041 , n4446 , n1491 );
    or g1924 ( n5011 , n4559 , n10651 );
    or g1925 ( n493 , n6395 , n2806 );
    nor g1926 ( n643 , n5087 , n5357 );
    and g1927 ( n558 , n11069 , n10056 );
    or g1928 ( n7113 , n7624 , n3139 );
    xnor g1929 ( n8424 , n5673 , n8784 );
    or g1930 ( n4519 , n22 , n5261 );
    and g1931 ( n12303 , n8211 , n12745 );
    or g1932 ( n11278 , n526 , n12480 );
    xnor g1933 ( n2241 , n122 , n11504 );
    and g1934 ( n3276 , n1886 , n4382 );
    xnor g1935 ( n8586 , n3749 , n8995 );
    xnor g1936 ( n3263 , n140 , n7811 );
    xnor g1937 ( n7442 , n3807 , n1967 );
    or g1938 ( n7947 , n9231 , n6051 );
    not g1939 ( n1134 , n634 );
    or g1940 ( n6857 , n6373 , n3606 );
    nor g1941 ( n9597 , n694 , n1527 );
    xnor g1942 ( n11052 , n4122 , n4225 );
    and g1943 ( n634 , n556 , n9483 );
    and g1944 ( n3846 , n5850 , n1347 );
    and g1945 ( n9603 , n11478 , n12489 );
    not g1946 ( n8301 , n1242 );
    or g1947 ( n613 , n10142 , n12843 );
    not g1948 ( n406 , n8914 );
    or g1949 ( n11544 , n10157 , n6922 );
    and g1950 ( n8064 , n5542 , n7234 );
    xnor g1951 ( n11081 , n11276 , n5298 );
    and g1952 ( n9795 , n10199 , n7637 );
    not g1953 ( n12617 , n9519 );
    xnor g1954 ( n10875 , n2781 , n2132 );
    xnor g1955 ( n2544 , n11679 , n1702 );
    nor g1956 ( n12538 , n3065 , n577 );
    or g1957 ( n10105 , n5999 , n7753 );
    xnor g1958 ( n4276 , n12788 , n1120 );
    or g1959 ( n969 , n7391 , n1079 );
    xnor g1960 ( n7103 , n9887 , n9226 );
    or g1961 ( n6377 , n1881 , n3482 );
    or g1962 ( n5488 , n3051 , n2323 );
    or g1963 ( n12227 , n4628 , n3924 );
    not g1964 ( n12186 , n10644 );
    not g1965 ( n5946 , n935 );
    xnor g1966 ( n353 , n8242 , n6266 );
    xnor g1967 ( n8440 , n3138 , n5747 );
    xnor g1968 ( n4087 , n9228 , n776 );
    xnor g1969 ( n3966 , n8534 , n12791 );
    or g1970 ( n1425 , n6571 , n11787 );
    xnor g1971 ( n417 , n7501 , n5037 );
    not g1972 ( n4540 , n8163 );
    and g1973 ( n10917 , n8097 , n3621 );
    xnor g1974 ( n11522 , n331 , n9121 );
    and g1975 ( n10146 , n9431 , n421 );
    and g1976 ( n6351 , n6635 , n9863 );
    or g1977 ( n10995 , n12797 , n2815 );
    and g1978 ( n881 , n12933 , n4152 );
    xnor g1979 ( n1847 , n3521 , n6605 );
    or g1980 ( n11327 , n10251 , n7741 );
    and g1981 ( n9507 , n10551 , n7988 );
    xnor g1982 ( n1262 , n9784 , n945 );
    and g1983 ( n4727 , n8336 , n12709 );
    and g1984 ( n6824 , n12141 , n11811 );
    or g1985 ( n2223 , n5809 , n12735 );
    not g1986 ( n8519 , n4650 );
    and g1987 ( n9485 , n11821 , n1798 );
    xnor g1988 ( n12174 , n1808 , n2210 );
    nor g1989 ( n1846 , n3474 , n5126 );
    nor g1990 ( n6512 , n4017 , n4070 );
    and g1991 ( n338 , n11782 , n5114 );
    xnor g1992 ( n12270 , n5791 , n3300 );
    not g1993 ( n9104 , n6988 );
    or g1994 ( n158 , n4911 , n7881 );
    xor g1995 ( n11858 , n3196 , n10766 );
    or g1996 ( n8903 , n5575 , n10903 );
    not g1997 ( n1717 , n5948 );
    and g1998 ( n11678 , n4961 , n231 );
    not g1999 ( n11627 , n9395 );
    or g2000 ( n10642 , n8921 , n1555 );
    or g2001 ( n1072 , n5355 , n6402 );
    and g2002 ( n6501 , n4243 , n8520 );
    nor g2003 ( n921 , n7936 , n1021 );
    and g2004 ( n5642 , n3756 , n2970 );
    or g2005 ( n9530 , n10196 , n4474 );
    or g2006 ( n5771 , n1462 , n10617 );
    and g2007 ( n9572 , n6376 , n7343 );
    not g2008 ( n12499 , n9896 );
    nor g2009 ( n6448 , n8675 , n9295 );
    and g2010 ( n8392 , n6888 , n11121 );
    and g2011 ( n8794 , n7058 , n6484 );
    xnor g2012 ( n9647 , n11392 , n10994 );
    xnor g2013 ( n6405 , n2303 , n6676 );
    and g2014 ( n7277 , n11126 , n687 );
    not g2015 ( n8969 , n4756 );
    or g2016 ( n9786 , n2595 , n920 );
    or g2017 ( n11109 , n6977 , n3421 );
    or g2018 ( n3218 , n8552 , n10854 );
    xnor g2019 ( n9646 , n11094 , n7005 );
    xnor g2020 ( n11258 , n9176 , n11849 );
    xnor g2021 ( n3575 , n7527 , n5344 );
    or g2022 ( n899 , n10157 , n5759 );
    and g2023 ( n2378 , n1663 , n4964 );
    xnor g2024 ( n1490 , n3403 , n3675 );
    or g2025 ( n4347 , n12841 , n6563 );
    or g2026 ( n7912 , n7283 , n7881 );
    or g2027 ( n8048 , n659 , n2151 );
    xnor g2028 ( n2110 , n5358 , n764 );
    and g2029 ( n9872 , n7177 , n8407 );
    xnor g2030 ( n11561 , n9894 , n5047 );
    xnor g2031 ( n12863 , n10377 , n11 );
    and g2032 ( n4827 , n6931 , n4506 );
    or g2033 ( n2209 , n5355 , n11827 );
    and g2034 ( n4908 , n2538 , n2861 );
    or g2035 ( n8585 , n12119 , n10854 );
    and g2036 ( n12576 , n6579 , n3093 );
    or g2037 ( n5340 , n8371 , n4073 );
    xnor g2038 ( n6178 , n8579 , n1647 );
    and g2039 ( n1439 , n6743 , n4503 );
    or g2040 ( n9875 , n9653 , n3928 );
    xnor g2041 ( n9356 , n4949 , n3083 );
    not g2042 ( n4096 , n5380 );
    xnor g2043 ( n8483 , n9799 , n12802 );
    or g2044 ( n3087 , n10750 , n826 );
    or g2045 ( n3954 , n12237 , n1932 );
    xnor g2046 ( n9139 , n2028 , n3245 );
    xnor g2047 ( n8930 , n7587 , n10511 );
    xnor g2048 ( n12072 , n5523 , n12349 );
    not g2049 ( n11238 , n8660 );
    or g2050 ( n9151 , n9835 , n11151 );
    not g2051 ( n254 , n4135 );
    and g2052 ( n10570 , n7899 , n5485 );
    not g2053 ( n12580 , n3945 );
    not g2054 ( n11887 , n6797 );
    xnor g2055 ( n1194 , n12155 , n10506 );
    or g2056 ( n7916 , n10142 , n9589 );
    and g2057 ( n7797 , n9849 , n8268 );
    xnor g2058 ( n8444 , n4110 , n11565 );
    and g2059 ( n1856 , n6277 , n8368 );
    not g2060 ( n6505 , n5869 );
    xnor g2061 ( n6116 , n4360 , n702 );
    xnor g2062 ( n7247 , n11899 , n477 );
    or g2063 ( n11074 , n4932 , n12548 );
    and g2064 ( n11388 , n9454 , n6302 );
    nor g2065 ( n3794 , n5877 , n653 );
    or g2066 ( n2807 , n11608 , n6029 );
    or g2067 ( n2816 , n8617 , n2375 );
    and g2068 ( n10290 , n11521 , n7438 );
    not g2069 ( n5351 , n6574 );
    and g2070 ( n11711 , n3197 , n6057 );
    and g2071 ( n10639 , n12178 , n5402 );
    or g2072 ( n11653 , n2579 , n4751 );
    not g2073 ( n3275 , n4664 );
    not g2074 ( n3636 , n12068 );
    or g2075 ( n7718 , n11923 , n4474 );
    or g2076 ( n12665 , n854 , n1710 );
    and g2077 ( n9590 , n12299 , n11023 );
    or g2078 ( n6132 , n8738 , n28 );
    xnor g2079 ( n798 , n1853 , n1577 );
    xnor g2080 ( n710 , n2777 , n10319 );
    xnor g2081 ( n8892 , n4998 , n6646 );
    xnor g2082 ( n10214 , n82 , n3917 );
    or g2083 ( n7895 , n1629 , n11103 );
    or g2084 ( n4974 , n3461 , n8923 );
    xnor g2085 ( n11781 , n3471 , n355 );
    xnor g2086 ( n9320 , n504 , n8915 );
    not g2087 ( n9824 , n2869 );
    xnor g2088 ( n4687 , n7144 , n4713 );
    not g2089 ( n3053 , n3396 );
    not g2090 ( n7424 , n12720 );
    or g2091 ( n5778 , n264 , n3350 );
    nor g2092 ( n11647 , n5882 , n786 );
    or g2093 ( n11864 , n12853 , n9188 );
    not g2094 ( n7731 , n7401 );
    and g2095 ( n3716 , n12501 , n7631 );
    not g2096 ( n4648 , n10167 );
    and g2097 ( n6741 , n5466 , n4578 );
    or g2098 ( n2220 , n876 , n11561 );
    or g2099 ( n5330 , n375 , n11346 );
    xnor g2100 ( n9251 , n12632 , n2990 );
    not g2101 ( n8870 , n7160 );
    or g2102 ( n2261 , n4488 , n11502 );
    not g2103 ( n1164 , n7252 );
    xnor g2104 ( n11227 , n6239 , n8808 );
    or g2105 ( n5554 , n3587 , n2295 );
    and g2106 ( n12219 , n1333 , n6038 );
    xnor g2107 ( n10299 , n7916 , n2642 );
    xnor g2108 ( n12860 , n6635 , n9193 );
    xnor g2109 ( n12055 , n11303 , n1614 );
    or g2110 ( n3821 , n6849 , n10786 );
    and g2111 ( n7198 , n8002 , n8934 );
    or g2112 ( n9472 , n8390 , n2744 );
    xnor g2113 ( n1069 , n7756 , n4681 );
    xnor g2114 ( n9230 , n1260 , n1053 );
    xnor g2115 ( n11383 , n2073 , n8420 );
    or g2116 ( n1154 , n2217 , n5086 );
    xnor g2117 ( n11140 , n5801 , n4160 );
    or g2118 ( n10535 , n10938 , n5356 );
    xnor g2119 ( n7252 , n12268 , n4486 );
    and g2120 ( n113 , n2033 , n8014 );
    nor g2121 ( n11839 , n9324 , n12805 );
    xnor g2122 ( n11454 , n7083 , n12586 );
    or g2123 ( n4089 , n3746 , n12816 );
    xnor g2124 ( n3159 , n8143 , n976 );
    and g2125 ( n903 , n5940 , n6495 );
    xnor g2126 ( n3437 , n12387 , n4258 );
    and g2127 ( n11642 , n12886 , n4117 );
    xnor g2128 ( n8904 , n5428 , n2647 );
    xnor g2129 ( n2492 , n8193 , n4752 );
    not g2130 ( n7351 , n9059 );
    xnor g2131 ( n7415 , n2704 , n6163 );
    xnor g2132 ( n5313 , n11080 , n3441 );
    and g2133 ( n11041 , n8377 , n5770 );
    xnor g2134 ( n5750 , n8736 , n6643 );
    not g2135 ( n6678 , n3910 );
    and g2136 ( n1214 , n5650 , n11675 );
    and g2137 ( n9459 , n12841 , n6563 );
    and g2138 ( n1259 , n4633 , n6062 );
    nor g2139 ( n2835 , n2779 , n8001 );
    xnor g2140 ( n10566 , n2869 , n6292 );
    nor g2141 ( n8168 , n10320 , n2747 );
    not g2142 ( n5479 , n2100 );
    or g2143 ( n2980 , n9370 , n12843 );
    nor g2144 ( n8771 , n5023 , n4063 );
    or g2145 ( n6756 , n2906 , n6213 );
    xnor g2146 ( n2693 , n9778 , n4240 );
    and g2147 ( n10333 , n4469 , n1428 );
    or g2148 ( n12938 , n9563 , n3881 );
    xnor g2149 ( n340 , n8795 , n12151 );
    or g2150 ( n5277 , n9389 , n12328 );
    xnor g2151 ( n1804 , n5122 , n10977 );
    and g2152 ( n4734 , n6770 , n2508 );
    and g2153 ( n936 , n5177 , n10438 );
    xnor g2154 ( n5534 , n7684 , n12162 );
    and g2155 ( n9560 , n673 , n7022 );
    xnor g2156 ( n2310 , n2502 , n11123 );
    not g2157 ( n9680 , n6768 );
    and g2158 ( n1625 , n10612 , n12938 );
    and g2159 ( n4781 , n4212 , n4350 );
    not g2160 ( n11868 , n4991 );
    xnor g2161 ( n8578 , n2945 , n5725 );
    or g2162 ( n7046 , n9043 , n10840 );
    xnor g2163 ( n5581 , n2897 , n12421 );
    or g2164 ( n11816 , n8583 , n12771 );
    or g2165 ( n1241 , n994 , n10419 );
    and g2166 ( n6385 , n9616 , n5262 );
    and g2167 ( n8670 , n1239 , n5737 );
    nor g2168 ( n5510 , n7563 , n9272 );
    xnor g2169 ( n472 , n2761 , n1190 );
    not g2170 ( n220 , n3264 );
    xnor g2171 ( n9641 , n10728 , n8985 );
    xnor g2172 ( n5297 , n12717 , n10156 );
    xnor g2173 ( n3923 , n7310 , n11202 );
    or g2174 ( n2405 , n10339 , n9188 );
    or g2175 ( n12173 , n11259 , n6119 );
    not g2176 ( n2531 , n12276 );
    or g2177 ( n7777 , n752 , n10919 );
    xnor g2178 ( n4379 , n11957 , n7460 );
    not g2179 ( n6071 , n503 );
    xnor g2180 ( n992 , n4977 , n104 );
    xnor g2181 ( n7446 , n11555 , n11609 );
    or g2182 ( n3585 , n7839 , n6169 );
    not g2183 ( n7041 , n7566 );
    nor g2184 ( n10040 , n1810 , n10778 );
    or g2185 ( n7913 , n4992 , n875 );
    xnor g2186 ( n10788 , n7215 , n4269 );
    xnor g2187 ( n2027 , n6567 , n11161 );
    and g2188 ( n3394 , n4675 , n5818 );
    or g2189 ( n5940 , n12467 , n918 );
    xnor g2190 ( n3987 , n9366 , n3063 );
    not g2191 ( n4654 , n405 );
    xnor g2192 ( n3090 , n11221 , n3260 );
    and g2193 ( n12666 , n4180 , n4990 );
    not g2194 ( n8530 , n2342 );
    or g2195 ( n12691 , n6718 , n1047 );
    and g2196 ( n2339 , n12479 , n8174 );
    xnor g2197 ( n11904 , n10118 , n5601 );
    not g2198 ( n10188 , n12637 );
    xnor g2199 ( n11780 , n11241 , n2062 );
    or g2200 ( n8274 , n3127 , n11746 );
    xnor g2201 ( n626 , n12271 , n12707 );
    xnor g2202 ( n4748 , n1872 , n625 );
    nor g2203 ( n8710 , n4239 , n5998 );
    and g2204 ( n12366 , n7071 , n8338 );
    or g2205 ( n10367 , n8870 , n10422 );
    not g2206 ( n6944 , n9487 );
    or g2207 ( n1747 , n349 , n3520 );
    not g2208 ( n4180 , n9869 );
    or g2209 ( n5178 , n4294 , n1120 );
    or g2210 ( n10674 , n4263 , n8131 );
    and g2211 ( n4447 , n5145 , n1247 );
    nor g2212 ( n10219 , n9445 , n651 );
    or g2213 ( n10925 , n6577 , n5012 );
    and g2214 ( n1621 , n5038 , n2570 );
    not g2215 ( n1117 , n3074 );
    xnor g2216 ( n10341 , n10380 , n4609 );
    or g2217 ( n6033 , n11887 , n8740 );
    not g2218 ( n9958 , n6039 );
    or g2219 ( n10509 , n3322 , n9842 );
    not g2220 ( n8695 , n8808 );
    xnor g2221 ( n3004 , n223 , n4172 );
    and g2222 ( n4450 , n1599 , n11816 );
    xnor g2223 ( n9340 , n6952 , n4592 );
    or g2224 ( n1731 , n3747 , n12249 );
    xnor g2225 ( n7278 , n7467 , n1063 );
    xnor g2226 ( n11834 , n812 , n11007 );
    nor g2227 ( n1388 , n9261 , n9726 );
    nor g2228 ( n10092 , n11234 , n12522 );
    xnor g2229 ( n8016 , n6612 , n3069 );
    or g2230 ( n2957 , n11887 , n8655 );
    and g2231 ( n4595 , n11980 , n3142 );
    not g2232 ( n1851 , n12591 );
    or g2233 ( n11498 , n5765 , n795 );
    and g2234 ( n9701 , n11796 , n5093 );
    not g2235 ( n1004 , n11208 );
    or g2236 ( n7612 , n8026 , n3421 );
    and g2237 ( n7566 , n6474 , n10755 );
    or g2238 ( n10477 , n12 , n3805 );
    xnor g2239 ( n7501 , n5742 , n10360 );
    or g2240 ( n10411 , n9365 , n3307 );
    or g2241 ( n12114 , n8552 , n12535 );
    and g2242 ( n3640 , n7038 , n6907 );
    nor g2243 ( n7373 , n4576 , n7365 );
    or g2244 ( n6730 , n4504 , n12036 );
    xnor g2245 ( n4997 , n3577 , n4372 );
    and g2246 ( n12132 , n288 , n11386 );
    or g2247 ( n11008 , n9693 , n8708 );
    xnor g2248 ( n1807 , n3626 , n5062 );
    and g2249 ( n1256 , n1542 , n9639 );
    xnor g2250 ( n2546 , n9677 , n4331 );
    or g2251 ( n8576 , n9370 , n11430 );
    and g2252 ( n3117 , n6407 , n2208 );
    and g2253 ( n506 , n6325 , n12504 );
    or g2254 ( n11417 , n3746 , n10903 );
    and g2255 ( n9500 , n321 , n3426 );
    or g2256 ( n7468 , n989 , n7341 );
    xnor g2257 ( n3610 , n12047 , n4004 );
    xnor g2258 ( n9392 , n1959 , n5349 );
    and g2259 ( n8561 , n10832 , n7421 );
    not g2260 ( n8541 , n8712 );
    or g2261 ( n1421 , n236 , n3770 );
    xnor g2262 ( n6289 , n3208 , n6757 );
    not g2263 ( n3803 , n4004 );
    not g2264 ( n5173 , n5522 );
    nor g2265 ( n7570 , n2318 , n9475 );
    nor g2266 ( n1141 , n2598 , n7576 );
    or g2267 ( n8896 , n5530 , n5781 );
    or g2268 ( n3684 , n8187 , n6402 );
    or g2269 ( n6993 , n7449 , n9280 );
    xnor g2270 ( n11091 , n835 , n7979 );
    xnor g2271 ( n7163 , n4723 , n8905 );
    or g2272 ( n7822 , n3467 , n11304 );
    not g2273 ( n1243 , n833 );
    and g2274 ( n1975 , n6306 , n12452 );
    not g2275 ( n11475 , n1973 );
    or g2276 ( n7416 , n3137 , n1711 );
    not g2277 ( n4793 , n12286 );
    and g2278 ( n832 , n3920 , n4934 );
    or g2279 ( n4612 , n8738 , n4474 );
    xnor g2280 ( n3696 , n11971 , n10228 );
    not g2281 ( n4822 , n3779 );
    and g2282 ( n12202 , n10721 , n8976 );
    and g2283 ( n5353 , n9560 , n12439 );
    xnor g2284 ( n8742 , n716 , n8670 );
    or g2285 ( n7694 , n1941 , n995 );
    not g2286 ( n11379 , n9851 );
    and g2287 ( n21 , n12363 , n9142 );
    or g2288 ( n3527 , n7801 , n6651 );
    or g2289 ( n12117 , n10879 , n12843 );
    and g2290 ( n3006 , n6364 , n8599 );
    and g2291 ( n6710 , n9785 , n574 );
    or g2292 ( n1456 , n8428 , n5538 );
    or g2293 ( n12758 , n337 , n12329 );
    or g2294 ( n10135 , n8583 , n3606 );
    xnor g2295 ( n11646 , n12054 , n2173 );
    and g2296 ( n11166 , n3172 , n7456 );
    xnor g2297 ( n4021 , n11700 , n11456 );
    xnor g2298 ( n8886 , n5466 , n4578 );
    xnor g2299 ( n956 , n12918 , n4606 );
    not g2300 ( n191 , n7862 );
    nor g2301 ( n2355 , n12200 , n6975 );
    or g2302 ( n12180 , n752 , n6084 );
    or g2303 ( n1981 , n8506 , n2381 );
    and g2304 ( n143 , n9250 , n10453 );
    and g2305 ( n10876 , n12955 , n873 );
    and g2306 ( n6369 , n5305 , n6038 );
    or g2307 ( n7567 , n962 , n1047 );
    not g2308 ( n10082 , n1187 );
    or g2309 ( n12051 , n8055 , n3802 );
    or g2310 ( n6439 , n2612 , n10166 );
    xnor g2311 ( n2376 , n9993 , n1281 );
    xnor g2312 ( n12338 , n2263 , n6568 );
    xnor g2313 ( n10828 , n2333 , n9209 );
    and g2314 ( n7536 , n6560 , n3741 );
    nor g2315 ( n1970 , n8663 , n5056 );
    xnor g2316 ( n10544 , n12544 , n9334 );
    xnor g2317 ( n11568 , n6708 , n7781 );
    and g2318 ( n6758 , n6347 , n9890 );
    and g2319 ( n5274 , n7982 , n7184 );
    or g2320 ( n2780 , n4343 , n3224 );
    or g2321 ( n8894 , n7391 , n4400 );
    xnor g2322 ( n2652 , n11120 , n280 );
    not g2323 ( n3868 , n1520 );
    or g2324 ( n9523 , n3746 , n9971 );
    or g2325 ( n8887 , n10992 , n12749 );
    not g2326 ( n1841 , n1511 );
    or g2327 ( n10185 , n11671 , n7681 );
    or g2328 ( n9205 , n10108 , n3911 );
    and g2329 ( n4556 , n5374 , n3182 );
    or g2330 ( n7012 , n3127 , n7703 );
    not g2331 ( n2769 , n1156 );
    xnor g2332 ( n760 , n5000 , n3649 );
    or g2333 ( n3205 , n989 , n10419 );
    nor g2334 ( n9879 , n9909 , n5227 );
    xnor g2335 ( n3239 , n12023 , n7734 );
    and g2336 ( n5208 , n619 , n8257 );
    or g2337 ( n1224 , n6836 , n2004 );
    xnor g2338 ( n8985 , n899 , n4424 );
    not g2339 ( n8478 , n479 );
    xnor g2340 ( n10456 , n363 , n7411 );
    or g2341 ( n438 , n8428 , n6455 );
    xnor g2342 ( n9294 , n1695 , n276 );
    or g2343 ( n7504 , n8026 , n9741 );
    or g2344 ( n11211 , n3188 , n689 );
    or g2345 ( n10361 , n10196 , n9144 );
    and g2346 ( n3026 , n726 , n3800 );
    or g2347 ( n1922 , n7449 , n4474 );
    xnor g2348 ( n1598 , n6201 , n1957 );
    or g2349 ( n12149 , n6069 , n2586 );
    or g2350 ( n1044 , n8583 , n1047 );
    xnor g2351 ( n10450 , n6361 , n4163 );
    xnor g2352 ( n9985 , n6598 , n10704 );
    xnor g2353 ( n6917 , n689 , n12152 );
    xnor g2354 ( n8023 , n841 , n7242 );
    or g2355 ( n51 , n8127 , n1079 );
    nor g2356 ( n10358 , n5646 , n3134 );
    xnor g2357 ( n2280 , n11142 , n10187 );
    not g2358 ( n117 , n9923 );
    xnor g2359 ( n6694 , n5769 , n7239 );
    and g2360 ( n8093 , n629 , n8432 );
    or g2361 ( n4237 , n12237 , n9188 );
    xnor g2362 ( n2294 , n9390 , n9482 );
    and g2363 ( n1518 , n834 , n5431 );
    or g2364 ( n2447 , n5575 , n9741 );
    xnor g2365 ( n5821 , n9103 , n11114 );
    xnor g2366 ( n12492 , n8666 , n10557 );
    not g2367 ( n2719 , n1624 );
    and g2368 ( n5999 , n4366 , n10752 );
    and g2369 ( n12283 , n6697 , n12225 );
    or g2370 ( n1380 , n8183 , n4720 );
    not g2371 ( n10065 , n774 );
    or g2372 ( n9351 , n5945 , n6169 );
    or g2373 ( n3181 , n1183 , n8109 );
    and g2374 ( n5365 , n6570 , n11756 );
    nor g2375 ( n9295 , n8243 , n2510 );
    and g2376 ( n440 , n3796 , n5592 );
    not g2377 ( n8683 , n4307 );
    xnor g2378 ( n6308 , n10056 , n9809 );
    or g2379 ( n255 , n7116 , n10903 );
    and g2380 ( n1507 , n9622 , n2782 );
    nor g2381 ( n9227 , n3116 , n9931 );
    or g2382 ( n11102 , n7116 , n11410 );
    or g2383 ( n12918 , n8187 , n4400 );
    nor g2384 ( n11815 , n2019 , n11218 );
    xnor g2385 ( n4756 , n38 , n6317 );
    or g2386 ( n275 , n2367 , n4527 );
    or g2387 ( n11413 , n4059 , n11827 );
    xnor g2388 ( n5552 , n10846 , n11890 );
    or g2389 ( n5357 , n989 , n4775 );
    or g2390 ( n1724 , n10108 , n4400 );
    xnor g2391 ( n9206 , n9442 , n12158 );
    or g2392 ( n11254 , n4961 , n231 );
    not g2393 ( n11637 , n4684 );
    or g2394 ( n4136 , n4059 , n5497 );
    or g2395 ( n10801 , n3632 , n2416 );
    or g2396 ( n4457 , n8428 , n7558 );
    xnor g2397 ( n6975 , n1586 , n4236 );
    xnor g2398 ( n745 , n845 , n5325 );
    or g2399 ( n11825 , n824 , n261 );
    or g2400 ( n7977 , n10751 , n4114 );
    xnor g2401 ( n10821 , n4124 , n1342 );
    xnor g2402 ( n11021 , n6004 , n7204 );
    xnor g2403 ( n1389 , n7194 , n3514 );
    or g2404 ( n10383 , n813 , n9865 );
    xnor g2405 ( n1029 , n3021 , n7548 );
    not g2406 ( n698 , n5337 );
    and g2407 ( n884 , n5501 , n4792 );
    and g2408 ( n1385 , n8279 , n3861 );
    and g2409 ( n2827 , n8336 , n6703 );
    and g2410 ( n10436 , n1043 , n11532 );
    or g2411 ( n2947 , n9878 , n3924 );
    or g2412 ( n3002 , n1795 , n1748 );
    and g2413 ( n1091 , n8269 , n5528 );
    or g2414 ( n12251 , n7283 , n1162 );
    and g2415 ( n4070 , n9441 , n7837 );
    xnor g2416 ( n7596 , n3829 , n8150 );
    and g2417 ( n6167 , n10075 , n4837 );
    xnor g2418 ( n8975 , n6414 , n4749 );
    not g2419 ( n1200 , n6535 );
    or g2420 ( n9309 , n12429 , n6135 );
    and g2421 ( n2873 , n11641 , n12379 );
    xnor g2422 ( n12258 , n7143 , n1997 );
    not g2423 ( n6340 , n8564 );
    or g2424 ( n8976 , n3215 , n2682 );
    and g2425 ( n2812 , n6859 , n8559 );
    xnor g2426 ( n1786 , n1724 , n3122 );
    xnor g2427 ( n1289 , n2292 , n9276 );
    and g2428 ( n4651 , n1421 , n1254 );
    xnor g2429 ( n12469 , n4167 , n5007 );
    or g2430 ( n9430 , n3405 , n9833 );
    xnor g2431 ( n2820 , n10238 , n3850 );
    xnor g2432 ( n1191 , n10771 , n9904 );
    xnor g2433 ( n6263 , n10745 , n3082 );
    or g2434 ( n161 , n5575 , n12899 );
    and g2435 ( n12321 , n614 , n4443 );
    or g2436 ( n4512 , n12361 , n11122 );
    xnor g2437 ( n8484 , n10 , n11277 );
    or g2438 ( n10842 , n636 , n3924 );
    and g2439 ( n9738 , n4324 , n1085 );
    or g2440 ( n8226 , n7606 , n9822 );
    nor g2441 ( n1626 , n12483 , n3830 );
    nor g2442 ( n8200 , n8806 , n110 );
    nor g2443 ( n9975 , n5709 , n886 );
    or g2444 ( n8752 , n1937 , n6455 );
    xnor g2445 ( n7676 , n4439 , n9375 );
    xnor g2446 ( n11213 , n3762 , n9060 );
    xnor g2447 ( n12634 , n9648 , n5802 );
    nor g2448 ( n2863 , n5607 , n7712 );
    and g2449 ( n10401 , n6616 , n10578 );
    or g2450 ( n8697 , n6265 , n8041 );
    and g2451 ( n8186 , n11588 , n5476 );
    xnor g2452 ( n4131 , n2233 , n1184 );
    or g2453 ( n8299 , n12853 , n530 );
    not g2454 ( n3670 , n6948 );
    or g2455 ( n1287 , n12237 , n4818 );
    xnor g2456 ( n7926 , n3116 , n4061 );
    not g2457 ( n4249 , n1576 );
    or g2458 ( n3772 , n6530 , n3167 );
    or g2459 ( n3338 , n7994 , n7450 );
    or g2460 ( n10079 , n8187 , n5497 );
    or g2461 ( n4754 , n9510 , n11586 );
    nor g2462 ( n12352 , n6268 , n2420 );
    and g2463 ( n9716 , n8406 , n2607 );
    not g2464 ( n11924 , n7097 );
    and g2465 ( n6278 , n6066 , n5292 );
    xnor g2466 ( n11206 , n1012 , n5547 );
    not g2467 ( n4400 , n11407 );
    or g2468 ( n1703 , n11310 , n6964 );
    nor g2469 ( n12095 , n5621 , n4075 );
    xnor g2470 ( n10016 , n8908 , n3736 );
    or g2471 ( n9748 , n994 , n4242 );
    or g2472 ( n3766 , n9748 , n10395 );
    not g2473 ( n8277 , n9319 );
    and g2474 ( n10335 , n10975 , n2152 );
    or g2475 ( n9634 , n5279 , n12258 );
    and g2476 ( n464 , n7396 , n5885 );
    and g2477 ( n8071 , n2215 , n6729 );
    not g2478 ( n12236 , n11545 );
    xnor g2479 ( n3121 , n11177 , n7836 );
    or g2480 ( n505 , n12853 , n8655 );
    or g2481 ( n5465 , n12742 , n11768 );
    or g2482 ( n6663 , n5355 , n9397 );
    xnor g2483 ( n6915 , n4510 , n6410 );
    or g2484 ( n6579 , n10142 , n7881 );
    not g2485 ( n6302 , n12055 );
    and g2486 ( n6064 , n11211 , n3438 );
    and g2487 ( n1320 , n7083 , n672 );
    and g2488 ( n10329 , n5279 , n12258 );
    xnor g2489 ( n11807 , n1542 , n5317 );
    and g2490 ( n7944 , n5923 , n412 );
    or g2491 ( n8785 , n10374 , n3898 );
    xnor g2492 ( n12005 , n9737 , n3263 );
    xnor g2493 ( n6420 , n1628 , n417 );
    xnor g2494 ( n3061 , n1312 , n2518 );
    xnor g2495 ( n9103 , n317 , n4065 );
    nor g2496 ( n4330 , n3362 , n2178 );
    not g2497 ( n10373 , n6086 );
    or g2498 ( n6241 , n7133 , n2395 );
    xnor g2499 ( n12650 , n5899 , n3201 );
    xnor g2500 ( n9621 , n12865 , n6627 );
    nor g2501 ( n11084 , n1371 , n6392 );
    and g2502 ( n7392 , n1908 , n315 );
    or g2503 ( n9519 , n3127 , n1546 );
    not g2504 ( n8297 , n10535 );
    or g2505 ( n2946 , n3603 , n2715 );
    not g2506 ( n880 , n8719 );
    nor g2507 ( n11667 , n8474 , n3774 );
    or g2508 ( n3030 , n11026 , n12120 );
    xnor g2509 ( n5483 , n8668 , n2206 );
    xnor g2510 ( n11641 , n9405 , n1794 );
    not g2511 ( n3079 , n7074 );
    and g2512 ( n5916 , n1777 , n304 );
    xnor g2513 ( n9478 , n2535 , n11416 );
    xnor g2514 ( n10697 , n7612 , n10080 );
    and g2515 ( n3681 , n11550 , n7051 );
    xnor g2516 ( n1818 , n1774 , n3777 );
    or g2517 ( n4885 , n10656 , n7948 );
    xnor g2518 ( n10164 , n7396 , n1995 );
    or g2519 ( n12310 , n3105 , n358 );
    not g2520 ( n310 , n1979 );
    and g2521 ( n7798 , n3742 , n390 );
    and g2522 ( n12506 , n8049 , n12510 );
    nor g2523 ( n6919 , n11879 , n11392 );
    xnor g2524 ( n6148 , n1608 , n9668 );
    and g2525 ( n9086 , n8169 , n6633 );
    xnor g2526 ( n1767 , n1457 , n8297 );
    xnor g2527 ( n4505 , n4210 , n12769 );
    not g2528 ( n7968 , n6289 );
    xnor g2529 ( n3975 , n8454 , n5734 );
    xnor g2530 ( n2283 , n12612 , n5537 );
    nor g2531 ( n12763 , n7630 , n5736 );
    xnor g2532 ( n9839 , n6234 , n11982 );
    not g2533 ( n1643 , n7454 );
    and g2534 ( n10857 , n10902 , n1393 );
    or g2535 ( n4144 , n9370 , n1738 );
    or g2536 ( n9155 , n11026 , n7506 );
    or g2537 ( n10855 , n11076 , n7067 );
    not g2538 ( n5018 , n5976 );
    not g2539 ( n3867 , n3858 );
    not g2540 ( n7834 , n11289 );
    or g2541 ( n6426 , n10835 , n8830 );
    xnor g2542 ( n5033 , n9054 , n1187 );
    nor g2543 ( n489 , n5542 , n7234 );
    nor g2544 ( n7353 , n3510 , n7366 );
    and g2545 ( n5909 , n4134 , n1943 );
    nor g2546 ( n3882 , n9429 , n7092 );
    xnor g2547 ( n11143 , n6246 , n10345 );
    or g2548 ( n1719 , n12853 , n4913 );
    and g2549 ( n8797 , n5730 , n10407 );
    or g2550 ( n1511 , n11474 , n9371 );
    nor g2551 ( n1028 , n11335 , n6518 );
    and g2552 ( n9269 , n12867 , n3434 );
    nor g2553 ( n9011 , n8682 , n1525 );
    or g2554 ( n4107 , n1183 , n1932 );
    not g2555 ( n4557 , n3776 );
    or g2556 ( n10121 , n11682 , n12092 );
    xnor g2557 ( n4663 , n4716 , n7053 );
    or g2558 ( n10572 , n5066 , n3226 );
    nor g2559 ( n9864 , n1074 , n5426 );
    not g2560 ( n11978 , n3877 );
    xnor g2561 ( n10967 , n5491 , n3664 );
    or g2562 ( n7054 , n10108 , n10066 );
    or g2563 ( n11443 , n5530 , n8259 );
    not g2564 ( n3717 , n3565 );
    xnor g2565 ( n8948 , n6122 , n189 );
    or g2566 ( n504 , n11958 , n3356 );
    and g2567 ( n11055 , n7862 , n2879 );
    xnor g2568 ( n4159 , n4766 , n3635 );
    xnor g2569 ( n5295 , n7251 , n4264 );
    xnor g2570 ( n1552 , n10046 , n6927 );
    or g2571 ( n7228 , n10104 , n10498 );
    or g2572 ( n5287 , n10269 , n3308 );
    nor g2573 ( n12832 , n905 , n11505 );
    xnor g2574 ( n6372 , n9708 , n4822 );
    not g2575 ( n9352 , n4948 );
    xnor g2576 ( n11651 , n1611 , n11337 );
    not g2577 ( n6885 , n11373 );
    xnor g2578 ( n2370 , n2244 , n5697 );
    or g2579 ( n1897 , n11890 , n4291 );
    or g2580 ( n7400 , n12361 , n3468 );
    or g2581 ( n5585 , n5889 , n802 );
    or g2582 ( n3895 , n752 , n1413 );
    xnor g2583 ( n8734 , n8124 , n3270 );
    or g2584 ( n5747 , n12565 , n903 );
    xnor g2585 ( n12358 , n3988 , n11105 );
    or g2586 ( n11265 , n8738 , n795 );
    nor g2587 ( n5835 , n1017 , n4853 );
    and g2588 ( n3257 , n8336 , n7500 );
    and g2589 ( n2267 , n11254 , n7847 );
    xnor g2590 ( n12140 , n11462 , n5398 );
    and g2591 ( n5577 , n10641 , n3867 );
    xnor g2592 ( n6079 , n11451 , n6853 );
    or g2593 ( n4564 , n7495 , n12843 );
    or g2594 ( n455 , n8752 , n1918 );
    not g2595 ( n10350 , n2365 );
    not g2596 ( n5419 , n7304 );
    or g2597 ( n4029 , n4380 , n5245 );
    xnor g2598 ( n5795 , n12671 , n1615 );
    or g2599 ( n12151 , n12136 , n9779 );
    xnor g2600 ( n12374 , n9745 , n3112 );
    or g2601 ( n12456 , n12503 , n4875 );
    or g2602 ( n11551 , n12774 , n2423 );
    nor g2603 ( n9936 , n6367 , n987 );
    nor g2604 ( n2779 , n4301 , n2204 );
    and g2605 ( n12652 , n12839 , n1279 );
    or g2606 ( n12731 , n11754 , n3073 );
    or g2607 ( n10513 , n6373 , n8285 );
    and g2608 ( n8089 , n7756 , n4681 );
    not g2609 ( n11552 , n5767 );
    xnor g2610 ( n7616 , n9035 , n4616 );
    xnor g2611 ( n11395 , n11720 , n11089 );
    xnor g2612 ( n9863 , n9247 , n9033 );
    nor g2613 ( n2967 , n1612 , n4673 );
    or g2614 ( n2772 , n12245 , n300 );
    or g2615 ( n2293 , n11928 , n11308 );
    not g2616 ( n11294 , n7658 );
    or g2617 ( n6780 , n8854 , n1035 );
    and g2618 ( n6046 , n12739 , n3108 );
    nor g2619 ( n4951 , n5463 , n12693 );
    and g2620 ( n718 , n7074 , n4105 );
    or g2621 ( n1842 , n6625 , n12959 );
    and g2622 ( n12429 , n7176 , n506 );
    or g2623 ( n5438 , n3127 , n1851 );
    not g2624 ( n8371 , n391 );
    xnor g2625 ( n11312 , n3416 , n4687 );
    not g2626 ( n6036 , n7796 );
    not g2627 ( n1720 , n12693 );
    or g2628 ( n12933 , n7173 , n8125 );
    xnor g2629 ( n8824 , n3405 , n10106 );
    not g2630 ( n11494 , n6338 );
    xnor g2631 ( n2438 , n1124 , n8110 );
    or g2632 ( n5959 , n5355 , n510 );
    not g2633 ( n2579 , n11267 );
    xnor g2634 ( n1614 , n10735 , n4091 );
    xnor g2635 ( n5309 , n3628 , n894 );
    xnor g2636 ( n8989 , n862 , n2668 );
    or g2637 ( n5366 , n1941 , n2815 );
    and g2638 ( n10718 , n12214 , n4423 );
    or g2639 ( n11624 , n6718 , n9521 );
    or g2640 ( n8620 , n12009 , n788 );
    xnor g2641 ( n12162 , n5749 , n8809 );
    and g2642 ( n11492 , n8294 , n6316 );
    xnor g2643 ( n5403 , n1412 , n12957 );
    xnor g2644 ( n4462 , n11824 , n1545 );
    or g2645 ( n10094 , n754 , n624 );
    xnor g2646 ( n3931 , n10215 , n4848 );
    or g2647 ( n6137 , n191 , n9589 );
    and g2648 ( n6319 , n6003 , n11614 );
    xnor g2649 ( n4619 , n5758 , n8210 );
    xnor g2650 ( n8995 , n8972 , n2667 );
    and g2651 ( n9410 , n11879 , n11392 );
    xnor g2652 ( n2965 , n11532 , n1195 );
    or g2653 ( n8327 , n343 , n7278 );
    xnor g2654 ( n3568 , n11053 , n5745 );
    xnor g2655 ( n8022 , n1803 , n6421 );
    xnor g2656 ( n9358 , n11723 , n8487 );
    and g2657 ( n1229 , n10545 , n7733 );
    not g2658 ( n9218 , n669 );
    xnor g2659 ( n3811 , n1707 , n700 );
    not g2660 ( n8624 , n1132 );
    and g2661 ( n4071 , n10698 , n7208 );
    and g2662 ( n11934 , n12814 , n8431 );
    not g2663 ( n12621 , n1410 );
    or g2664 ( n10109 , n10714 , n43 );
    not g2665 ( n2898 , n860 );
    or g2666 ( n3015 , n5575 , n6084 );
    xnor g2667 ( n7062 , n1569 , n7211 );
    nor g2668 ( n3969 , n11042 , n6350 );
    or g2669 ( n3033 , n9286 , n2889 );
    or g2670 ( n12370 , n12393 , n1463 );
    xnor g2671 ( n11835 , n6097 , n4496 );
    or g2672 ( n4446 , n11923 , n1476 );
    or g2673 ( n649 , n191 , n10066 );
    or g2674 ( n11065 , n1699 , n12754 );
    and g2675 ( n3829 , n9003 , n7006 );
    or g2676 ( n8123 , n2099 , n2259 );
    or g2677 ( n11259 , n8870 , n12080 );
    or g2678 ( n4723 , n8870 , n9586 );
    and g2679 ( n4407 , n6720 , n7516 );
    xnor g2680 ( n9095 , n656 , n3516 );
    nor g2681 ( n3400 , n2183 , n5920 );
    and g2682 ( n7901 , n1230 , n811 );
    not g2683 ( n388 , n3646 );
    and g2684 ( n173 , n11222 , n10848 );
    or g2685 ( n1438 , n3127 , n3911 );
    xnor g2686 ( n7866 , n3055 , n10950 );
    xnor g2687 ( n11260 , n5632 , n6483 );
    not g2688 ( n3884 , n9858 );
    xnor g2689 ( n10863 , n6543 , n5480 );
    or g2690 ( n2853 , n8552 , n8740 );
    not g2691 ( n9315 , n11499 );
    xnor g2692 ( n5535 , n9748 , n10395 );
    xnor g2693 ( n1010 , n11088 , n9952 );
    xnor g2694 ( n11629 , n10658 , n10946 );
    xnor g2695 ( n4776 , n6423 , n1125 );
    xnor g2696 ( n8938 , n4446 , n6647 );
    or g2697 ( n1848 , n7564 , n1363 );
    or g2698 ( n5020 , n6470 , n7392 );
    and g2699 ( n6548 , n11691 , n8511 );
    and g2700 ( n2570 , n4831 , n426 );
    nor g2701 ( n10447 , n7762 , n8302 );
    and g2702 ( n1451 , n3926 , n10474 );
    or g2703 ( n11883 , n3088 , n8080 );
    xnor g2704 ( n4334 , n2111 , n7631 );
    or g2705 ( n5087 , n10142 , n5851 );
    and g2706 ( n1532 , n9652 , n9798 );
    and g2707 ( n1349 , n9621 , n1490 );
    not g2708 ( n3199 , n10191 );
    or g2709 ( n10379 , n8738 , n9144 );
    not g2710 ( n916 , n12553 );
    not g2711 ( n2139 , n1451 );
    or g2712 ( n6883 , n6741 , n3136 );
    and g2713 ( n6739 , n6426 , n11009 );
    not g2714 ( n8909 , n4883 );
    not g2715 ( n3080 , n7977 );
    xnor g2716 ( n66 , n12263 , n3569 );
    or g2717 ( n6888 , n7322 , n256 );
    xnor g2718 ( n12035 , n9117 , n3266 );
    not g2719 ( n7710 , n3804 );
    nor g2720 ( n10177 , n1923 , n6640 );
    not g2721 ( n2122 , n8356 );
    and g2722 ( n2788 , n5413 , n10170 );
    or g2723 ( n1186 , n7151 , n7714 );
    xnor g2724 ( n601 , n7488 , n8876 );
    xnor g2725 ( n5390 , n6686 , n7599 );
    or g2726 ( n3755 , n6644 , n2461 );
    or g2727 ( n4244 , n8026 , n184 );
    not g2728 ( n6382 , n1324 );
    and g2729 ( n9236 , n12614 , n1022 );
    or g2730 ( n8736 , n5575 , n9971 );
    or g2731 ( n4920 , n10835 , n9521 );
    xnor g2732 ( n6961 , n4076 , n10213 );
    or g2733 ( n9543 , n6868 , n793 );
    not g2734 ( n12385 , n2350 );
    nor g2735 ( n7225 , n9336 , n11463 );
    and g2736 ( n6680 , n12223 , n7114 );
    or g2737 ( n12019 , n12183 , n10177 );
    nor g2738 ( n6850 , n2664 , n7797 );
    or g2739 ( n6147 , n4387 , n4162 );
    xnor g2740 ( n5720 , n6110 , n4199 );
    and g2741 ( n11480 , n9836 , n8081 );
    or g2742 ( n5371 , n7495 , n10066 );
    xnor g2743 ( n3283 , n4322 , n512 );
    or g2744 ( n6386 , n10744 , n2240 );
    or g2745 ( n5378 , n1003 , n6517 );
    xnor g2746 ( n1499 , n9752 , n7238 );
    nor g2747 ( n9 , n12538 , n10690 );
    xnor g2748 ( n544 , n2249 , n9983 );
    xnor g2749 ( n4353 , n11356 , n5342 );
    not g2750 ( n12686 , n7610 );
    or g2751 ( n3736 , n8959 , n3421 );
    and g2752 ( n9021 , n10018 , n10021 );
    not g2753 ( n11430 , n12000 );
    and g2754 ( n1263 , n1679 , n10359 );
    or g2755 ( n6979 , n289 , n11772 );
    and g2756 ( n805 , n9335 , n11031 );
    nor g2757 ( n9823 , n10195 , n3161 );
    xnor g2758 ( n235 , n4121 , n11975 );
    or g2759 ( n11386 , n8583 , n1509 );
    xnor g2760 ( n4701 , n8030 , n8060 );
    or g2761 ( n8727 , n9504 , n11910 );
    not g2762 ( n7293 , n5898 );
    and g2763 ( n9347 , n12218 , n2632 );
    nor g2764 ( n3228 , n6624 , n10834 );
    xnor g2765 ( n3515 , n5577 , n3204 );
    or g2766 ( n4576 , n5530 , n12124 );
    xor g2767 ( n2183 , n10004 , n6289 );
    xnor g2768 ( n6821 , n6461 , n3211 );
    and g2769 ( n12584 , n81 , n12343 );
    and g2770 ( n1898 , n2003 , n12762 );
    or g2771 ( n7748 , n4059 , n2358 );
    or g2772 ( n12761 , n989 , n5851 );
    or g2773 ( n3105 , n12361 , n9741 );
    xnor g2774 ( n7595 , n12114 , n944 );
    or g2775 ( n11470 , n4120 , n2805 );
    xnor g2776 ( n4270 , n9757 , n5806 );
    or g2777 ( n4129 , n7941 , n9113 );
    xnor g2778 ( n7164 , n5981 , n282 );
    and g2779 ( n6164 , n1073 , n6790 );
    and g2780 ( n10770 , n5860 , n10848 );
    not g2781 ( n3808 , n7405 );
    or g2782 ( n12567 , n2286 , n7581 );
    and g2783 ( n5736 , n7544 , n7228 );
    not g2784 ( n11944 , n12811 );
    not g2785 ( n8959 , n7436 );
    xnor g2786 ( n1466 , n1486 , n4221 );
    and g2787 ( n7178 , n6698 , n2158 );
    xnor g2788 ( n4172 , n1330 , n106 );
    not g2789 ( n486 , n10023 );
    or g2790 ( n4161 , n10750 , n12883 );
    nor g2791 ( n1959 , n12887 , n539 );
    xnor g2792 ( n9555 , n11284 , n5626 );
    xnor g2793 ( n8482 , n3065 , n7032 );
    xnor g2794 ( n7175 , n8776 , n123 );
    or g2795 ( n8404 , n3096 , n11896 );
    or g2796 ( n10354 , n12119 , n7928 );
    xnor g2797 ( n12054 , n10809 , n11107 );
    or g2798 ( n11162 , n6681 , n10894 );
    xnor g2799 ( n11219 , n815 , n11075 );
    and g2800 ( n1372 , n5066 , n3226 );
    or g2801 ( n9318 , n3664 , n6712 );
    xnor g2802 ( n4709 , n2215 , n6729 );
    not g2803 ( n3058 , n4838 );
    xnor g2804 ( n12014 , n2805 , n5521 );
    nor g2805 ( n10991 , n1361 , n8577 );
    or g2806 ( n6654 , n8870 , n7382 );
    not g2807 ( n2689 , n1479 );
    and g2808 ( n8165 , n23 , n7844 );
    nor g2809 ( n825 , n11745 , n2578 );
    not g2810 ( n3229 , n5819 );
    xnor g2811 ( n3391 , n9281 , n8563 );
    xnor g2812 ( n1971 , n7713 , n9343 );
    or g2813 ( n4964 , n10975 , n2152 );
    not g2814 ( n4674 , n4499 );
    xnor g2815 ( n7818 , n705 , n8192 );
    or g2816 ( n10480 , n12361 , n6169 );
    xnor g2817 ( n3354 , n933 , n12666 );
    xnor g2818 ( n9932 , n6222 , n9902 );
    not g2819 ( n4802 , n1880 );
    xnor g2820 ( n2565 , n396 , n8802 );
    xnor g2821 ( n8408 , n11489 , n1403 );
    not g2822 ( n7943 , n12700 );
    and g2823 ( n9169 , n1128 , n6110 );
    xnor g2824 ( n7482 , n2382 , n6633 );
    not g2825 ( n8090 , n8799 );
    xnor g2826 ( n7887 , n3804 , n3531 );
    or g2827 ( n4676 , n8738 , n3606 );
    nor g2828 ( n11721 , n3327 , n11046 );
    not g2829 ( n10982 , n12003 );
    or g2830 ( n243 , n6146 , n6749 );
    or g2831 ( n12856 , n9370 , n1455 );
    or g2832 ( n11547 , n10157 , n8643 );
    not g2833 ( n2790 , n5888 );
    and g2834 ( n2922 , n7012 , n2026 );
    or g2835 ( n10957 , n9193 , n6351 );
    xnor g2836 ( n12097 , n3209 , n8681 );
    or g2837 ( n78 , n5530 , n12080 );
    and g2838 ( n12733 , n11222 , n405 );
    or g2839 ( n770 , n6348 , n10175 );
    or g2840 ( n1053 , n11719 , n12843 );
    not g2841 ( n9536 , n10734 );
    xnor g2842 ( n3689 , n3966 , n11977 );
    or g2843 ( n1266 , n6577 , n2815 );
    and g2844 ( n12693 , n508 , n8530 );
    xnor g2845 ( n1712 , n4542 , n5403 );
    and g2846 ( n8569 , n12127 , n3081 );
    not g2847 ( n10773 , n8900 );
    xnor g2848 ( n7766 , n1787 , n7591 );
    or g2849 ( n11249 , n1539 , n1455 );
    or g2850 ( n4206 , n7283 , n7424 );
    xnor g2851 ( n2296 , n8353 , n1922 );
    or g2852 ( n7108 , n6650 , n5386 );
    xnor g2853 ( n10359 , n3182 , n4082 );
    or g2854 ( n8098 , n6111 , n212 );
    xnor g2855 ( n1485 , n10313 , n6603 );
    not g2856 ( n10910 , n82 );
    or g2857 ( n7465 , n8026 , n11775 );
    and g2858 ( n1736 , n646 , n494 );
    or g2859 ( n7370 , n4204 , n5028 );
    xnor g2860 ( n6023 , n12884 , n4139 );
    or g2861 ( n8847 , n12119 , n2964 );
    not g2862 ( n5462 , n3284 );
    and g2863 ( n6291 , n4811 , n8090 );
    xnor g2864 ( n8138 , n8460 , n5610 );
    xnor g2865 ( n5533 , n11935 , n10821 );
    or g2866 ( n8659 , n4059 , n4775 );
    or g2867 ( n9510 , n4498 , n11827 );
    not g2868 ( n11292 , n3206 );
    not g2869 ( n9335 , n11188 );
    xnor g2870 ( n5831 , n8704 , n11689 );
    or g2871 ( n10808 , n12853 , n7928 );
    not g2872 ( n3682 , n5284 );
    and g2873 ( n5880 , n8587 , n10206 );
    xnor g2874 ( n6702 , n8320 , n6588 );
    not g2875 ( n2804 , n742 );
    xnor g2876 ( n9947 , n9620 , n9238 );
    xnor g2877 ( n2932 , n1356 , n10540 );
    xnor g2878 ( n6533 , n11997 , n930 );
    xnor g2879 ( n8680 , n6073 , n8947 );
    and g2880 ( n5350 , n11841 , n3002 );
    or g2881 ( n10974 , n4628 , n12535 );
    or g2882 ( n8945 , n1051 , n9741 );
    xor g2883 ( n4686 , n1027 , n3950 );
    not g2884 ( n10157 , n3992 );
    nor g2885 ( n7029 , n10878 , n5623 );
    xnor g2886 ( n10559 , n2397 , n12403 );
    or g2887 ( n10587 , n8552 , n7382 );
    or g2888 ( n6701 , n11445 , n247 );
    xnor g2889 ( n985 , n1266 , n6324 );
    or g2890 ( n2672 , n8552 , n8109 );
    xnor g2891 ( n7426 , n5263 , n3657 );
    or g2892 ( n365 , n1699 , n10854 );
    and g2893 ( n10403 , n1594 , n10964 );
    or g2894 ( n5486 , n8583 , n9521 );
    nor g2895 ( n4445 , n3988 , n5039 );
    and g2896 ( n8237 , n10118 , n5887 );
    or g2897 ( n1854 , n11226 , n2658 );
    not g2898 ( n3356 , n8236 );
    nor g2899 ( n1319 , n4718 , n3634 );
    nor g2900 ( n4278 , n7643 , n913 );
    and g2901 ( n7275 , n637 , n5996 );
    and g2902 ( n8878 , n10434 , n9894 );
    and g2903 ( n6024 , n197 , n8330 );
    or g2904 ( n6398 , n3713 , n3227 );
    nor g2905 ( n1323 , n6865 , n9059 );
    not g2906 ( n11119 , n6353 );
    or g2907 ( n6117 , n1856 , n3748 );
    or g2908 ( n6581 , n8354 , n6513 );
    xnor g2909 ( n1177 , n12471 , n535 );
    nor g2910 ( n11035 , n12524 , n8898 );
    and g2911 ( n7067 , n762 , n6312 );
    and g2912 ( n7301 , n2251 , n4277 );
    nor g2913 ( n2196 , n7897 , n4918 );
    xnor g2914 ( n3124 , n12267 , n7399 );
    and g2915 ( n9753 , n9279 , n10331 );
    or g2916 ( n5844 , n11182 , n4200 );
    xnor g2917 ( n600 , n3906 , n11203 );
    xnor g2918 ( n7222 , n1536 , n12651 );
    xnor g2919 ( n11284 , n1347 , n7216 );
    xnor g2920 ( n5517 , n9467 , n9312 );
    or g2921 ( n4856 , n5575 , n8768 );
    or g2922 ( n1639 , n8428 , n12816 );
    not g2923 ( n4348 , n707 );
    and g2924 ( n8844 , n2226 , n2522 );
    not g2925 ( n9586 , n11967 );
    xnor g2926 ( n10711 , n10724 , n10581 );
    or g2927 ( n9887 , n6977 , n9741 );
    and g2928 ( n4919 , n2930 , n4901 );
    or g2929 ( n5251 , n636 , n3224 );
    and g2930 ( n2707 , n12263 , n9203 );
    xnor g2931 ( n10705 , n582 , n11014 );
    xnor g2932 ( n2796 , n3976 , n10429 );
    not g2933 ( n8211 , n7277 );
    not g2934 ( n6182 , n1082 );
    xnor g2935 ( n2320 , n4191 , n6555 );
    xnor g2936 ( n10693 , n3396 , n12700 );
    not g2937 ( n10606 , n10171 );
    nor g2938 ( n12088 , n6894 , n7105 );
    and g2939 ( n12628 , n1842 , n10943 );
    xnor g2940 ( n12058 , n6514 , n5373 );
    xnor g2941 ( n11246 , n4597 , n394 );
    xnor g2942 ( n458 , n1873 , n11223 );
    or g2943 ( n8751 , n10835 , n1739 );
    xnor g2944 ( n1428 , n2274 , n11858 );
    and g2945 ( n6226 , n7243 , n2460 );
    xnor g2946 ( n3869 , n8097 , n4520 );
    xnor g2947 ( n10192 , n3888 , n10029 );
    and g2948 ( n12689 , n116 , n5826 );
    and g2949 ( n7540 , n9656 , n12411 );
    and g2950 ( n10259 , n1951 , n11244 );
    nor g2951 ( n5099 , n9461 , n6363 );
    nor g2952 ( n9962 , n5963 , n4102 );
    xor g2953 ( n112 , n9321 , n3824 );
    xnor g2954 ( n12943 , n8545 , n4824 );
    or g2955 ( n11973 , n9389 , n11430 );
    xnor g2956 ( n4469 , n1949 , n12487 );
    xnor g2957 ( n9405 , n8949 , n6724 );
    and g2958 ( n11263 , n8322 , n6737 );
    nor g2959 ( n12887 , n6751 , n3519 );
    or g2960 ( n1112 , n1051 , n7425 );
    or g2961 ( n4675 , n2613 , n3826 );
    xnor g2962 ( n1118 , n4001 , n592 );
    or g2963 ( n2398 , n4628 , n6513 );
    xnor g2964 ( n5304 , n6728 , n3827 );
    xnor g2965 ( n6938 , n2991 , n8769 );
    nor g2966 ( n540 , n2561 , n6572 );
    xnor g2967 ( n3100 , n9230 , n8689 );
    xnor g2968 ( n6834 , n4437 , n5220 );
    nor g2969 ( n1379 , n1127 , n11848 );
    and g2970 ( n482 , n10697 , n4968 );
    xnor g2971 ( n9613 , n3792 , n1244 );
    xnor g2972 ( n5555 , n7009 , n7664 );
    or g2973 ( n12912 , n11887 , n12080 );
    xnor g2974 ( n6520 , n5334 , n4884 );
    nor g2975 ( n11804 , n5335 , n9207 );
    xnor g2976 ( n3046 , n11960 , n3273 );
    or g2977 ( n2414 , n3145 , n1267 );
    xnor g2978 ( n2584 , n7983 , n2334 );
    xnor g2979 ( n5109 , n4315 , n8832 );
    nor g2980 ( n6037 , n10203 , n7219 );
    xnor g2981 ( n8840 , n5988 , n6856 );
    nor g2982 ( n6341 , n6874 , n10455 );
    xnor g2983 ( n2146 , n8635 , n2698 );
    xnor g2984 ( n8942 , n35 , n9110 );
    xnor g2985 ( n9502 , n9432 , n7226 );
    xnor g2986 ( n7781 , n8319 , n8044 );
    not g2987 ( n2445 , n5371 );
    xnor g2988 ( n11216 , n7230 , n9154 );
    nor g2989 ( n10247 , n8092 , n5459 );
    xnor g2990 ( n12111 , n7708 , n2758 );
    or g2991 ( n4384 , n1288 , n2868 );
    and g2992 ( n10486 , n2854 , n1961 );
    not g2993 ( n9210 , n292 );
    or g2994 ( n9622 , n11228 , n8573 );
    or g2995 ( n6560 , n5765 , n4642 );
    xnor g2996 ( n4024 , n3928 , n9075 );
    xnor g2997 ( n5859 , n8254 , n6490 );
    xnor g2998 ( n4058 , n2975 , n10901 );
    nor g2999 ( n1468 , n3329 , n9053 );
    and g3000 ( n2861 , n7965 , n9763 );
    xnor g3001 ( n4538 , n10048 , n9129 );
    nor g3002 ( n9643 , n3954 , n8955 );
    or g3003 ( n10727 , n346 , n7721 );
    or g3004 ( n11905 , n1937 , n7876 );
    or g3005 ( n8946 , n60 , n11213 );
    or g3006 ( n1267 , n8428 , n5012 );
    or g3007 ( n2893 , n5355 , n7341 );
    nor g3008 ( n5986 , n12870 , n10107 );
    not g3009 ( n3617 , n1199 );
    or g3010 ( n4994 , n994 , n7341 );
    or g3011 ( n2874 , n5575 , n8414 );
    not g3012 ( n2134 , n6946 );
    or g3013 ( n1566 , n10010 , n10815 );
    and g3014 ( n2436 , n8900 , n5531 );
    xnor g3015 ( n5639 , n3653 , n2021 );
    and g3016 ( n7552 , n11317 , n1265 );
    and g3017 ( n8102 , n10464 , n4164 );
    or g3018 ( n1305 , n2064 , n5122 );
    or g3019 ( n11133 , n2619 , n4978 );
    xnor g3020 ( n3785 , n4256 , n5534 );
    not g3021 ( n5006 , n8765 );
    or g3022 ( n1024 , n12119 , n1163 );
    not g3023 ( n6455 , n3719 );
    not g3024 ( n2716 , n8275 );
    or g3025 ( n5589 , n10835 , n4642 );
    or g3026 ( n12090 , n3715 , n9788 );
    or g3027 ( n1695 , n9370 , n7881 );
    or g3028 ( n8981 , n5059 , n11994 );
    xnor g3029 ( n7008 , n110 , n2882 );
    not g3030 ( n269 , n9581 );
    or g3031 ( n8991 , n2850 , n9469 );
    and g3032 ( n11732 , n2408 , n1931 );
    or g3033 ( n10210 , n4778 , n7382 );
    nor g3034 ( n12857 , n9907 , n9927 );
    xnor g3035 ( n8621 , n6085 , n4762 );
    xnor g3036 ( n5997 , n7037 , n8613 );
    or g3037 ( n9196 , n8187 , n3911 );
    nor g3038 ( n7417 , n6165 , n8787 );
    xnor g3039 ( n7039 , n10877 , n4406 );
    and g3040 ( n1531 , n7195 , n7793 );
    xnor g3041 ( n230 , n7457 , n9017 );
    xnor g3042 ( n10724 , n11537 , n11206 );
    nor g3043 ( n8883 , n8750 , n10537 );
    or g3044 ( n4941 , n7503 , n11066 );
    not g3045 ( n5121 , n5590 );
    xnor g3046 ( n5117 , n5969 , n11591 );
    or g3047 ( n7509 , n6577 , n6455 );
    or g3048 ( n7121 , n5765 , n1476 );
    or g3049 ( n5732 , n191 , n1455 );
    xnor g3050 ( n12508 , n12059 , n2796 );
    and g3051 ( n1900 , n6131 , n2060 );
    or g3052 ( n12680 , n8406 , n2607 );
    and g3053 ( n2060 , n3486 , n7825 );
    xnor g3054 ( n8953 , n12761 , n50 );
    xnor g3055 ( n3731 , n10435 , n4895 );
    xnor g3056 ( n9412 , n8750 , n6167 );
    not g3057 ( n5156 , n8289 );
    and g3058 ( n11777 , n9138 , n2135 );
    not g3059 ( n265 , n7576 );
    or g3060 ( n2162 , n5765 , n7921 );
    or g3061 ( n2732 , n7149 , n9026 );
    and g3062 ( n8050 , n12385 , n12353 );
    and g3063 ( n12326 , n4500 , n1483 );
    nor g3064 ( n3763 , n9814 , n9609 );
    and g3065 ( n3321 , n6650 , n5386 );
    or g3066 ( n11169 , n1899 , n5376 );
    or g3067 ( n101 , n1197 , n4827 );
    nor g3068 ( n12238 , n2227 , n9716 );
    or g3069 ( n10542 , n8496 , n4583 );
    not g3070 ( n1047 , n1980 );
    or g3071 ( n1102 , n2363 , n229 );
    nor g3072 ( n12491 , n10346 , n7372 );
    and g3073 ( n8603 , n5077 , n12350 );
    not g3074 ( n10382 , n5029 );
    not g3075 ( n3597 , n11953 );
    not g3076 ( n7634 , n3881 );
    or g3077 ( n4254 , n11958 , n5311 );
    xnor g3078 ( n10654 , n5569 , n1877 );
    xnor g3079 ( n3450 , n9108 , n3983 );
    not g3080 ( n1175 , n11198 );
    or g3081 ( n830 , n6090 , n2811 );
    and g3082 ( n2806 , n9231 , n6051 );
    not g3083 ( n12603 , n11685 );
    not g3084 ( n1575 , n4492 );
    or g3085 ( n5453 , n2217 , n3599 );
    and g3086 ( n9739 , n4805 , n1564 );
    or g3087 ( n5948 , n8026 , n11410 );
    not g3088 ( n8470 , n9842 );
    and g3089 ( n1146 , n9797 , n2900 );
    xnor g3090 ( n3898 , n1037 , n2402 );
    or g3091 ( n10806 , n11239 , n5980 );
    not g3092 ( n6128 , n5673 );
    xnor g3093 ( n9792 , n7827 , n711 );
    or g3094 ( n4289 , n752 , n3468 );
    or g3095 ( n3678 , n11923 , n609 );
    and g3096 ( n10081 , n5995 , n769 );
    nor g3097 ( n3630 , n8817 , n4099 );
    xnor g3098 ( n7259 , n9655 , n865 );
    or g3099 ( n2326 , n7449 , n3606 );
    xnor g3100 ( n170 , n12492 , n425 );
    not g3101 ( n4305 , n3257 );
    not g3102 ( n4973 , n3428 );
    xnor g3103 ( n3676 , n12104 , n11215 );
    or g3104 ( n7334 , n4059 , n6389 );
    not g3105 ( n9726 , n2440 );
    or g3106 ( n7114 , n9389 , n8524 );
    not g3107 ( n1941 , n4187 );
    and g3108 ( n3619 , n12052 , n9818 );
    xnor g3109 ( n1218 , n2268 , n7047 );
    or g3110 ( n11234 , n11552 , n9144 );
    not g3111 ( n7560 , n131 );
    or g3112 ( n11998 , n6577 , n2232 );
    xnor g3113 ( n8979 , n10730 , n4507 );
    not g3114 ( n8375 , n267 );
    or g3115 ( n628 , n3097 , n7281 );
    xnor g3116 ( n2375 , n6326 , n6631 );
    and g3117 ( n4900 , n1814 , n739 );
    not g3118 ( n3280 , n5405 );
    or g3119 ( n8729 , n9976 , n1638 );
    or g3120 ( n9000 , n10835 , n3606 );
    and g3121 ( n4010 , n2562 , n5484 );
    xnor g3122 ( n48 , n11025 , n6958 );
    or g3123 ( n9908 , n2213 , n1443 );
    or g3124 ( n8256 , n973 , n12170 );
    xnor g3125 ( n12048 , n12879 , n10887 );
    xnor g3126 ( n5911 , n54 , n11751 );
    xor g3127 ( n7680 , n250 , n11151 );
    xnor g3128 ( n10599 , n10018 , n10021 );
    and g3129 ( n7205 , n1471 , n8028 );
    and g3130 ( n9367 , n7268 , n1767 );
    and g3131 ( n11252 , n9141 , n5149 );
    not g3132 ( n10827 , n7233 );
    and g3133 ( n449 , n10532 , n7374 );
    and g3134 ( n1232 , n8538 , n1504 );
    or g3135 ( n6244 , n11552 , n3606 );
    and g3136 ( n8919 , n5577 , n7816 );
    xnor g3137 ( n8971 , n4561 , n10280 );
    xnor g3138 ( n12239 , n12775 , n12157 );
    xnor g3139 ( n5133 , n7605 , n3031 );
    and g3140 ( n6631 , n9182 , n6245 );
    or g3141 ( n10309 , n3743 , n8830 );
    and g3142 ( n12435 , n1708 , n12114 );
    or g3143 ( n11621 , n6413 , n166 );
    xor g3144 ( n6742 , n3166 , n3894 );
    nor g3145 ( n6600 , n12129 , n12573 );
    or g3146 ( n3038 , n9370 , n11827 );
    xnor g3147 ( n10567 , n3543 , n4861 );
    or g3148 ( n1166 , n11433 , n12816 );
    xnor g3149 ( n9283 , n2817 , n12589 );
    xnor g3150 ( n6436 , n12370 , n10650 );
    or g3151 ( n1943 , n2118 , n1155 );
    xnor g3152 ( n169 , n11073 , n10424 );
    xnor g3153 ( n3075 , n8054 , n9338 );
    or g3154 ( n385 , n5038 , n2570 );
    not g3155 ( n1996 , n7035 );
    or g3156 ( n1137 , n1233 , n6330 );
    and g3157 ( n10220 , n2536 , n12112 );
    or g3158 ( n5505 , n2067 , n12568 );
    xnor g3159 ( n10481 , n7332 , n6932 );
    or g3160 ( n9308 , n10142 , n2358 );
    or g3161 ( n12350 , n3874 , n6060 );
    or g3162 ( n7128 , n6055 , n6997 );
    or g3163 ( n11293 , n705 , n1310 );
    nor g3164 ( n6868 , n9692 , n4439 );
    not g3165 ( n2046 , n1104 );
    or g3166 ( n2243 , n10390 , n10883 );
    not g3167 ( n10364 , n12949 );
    xnor g3168 ( n10417 , n267 , n3548 );
    xnor g3169 ( n9388 , n1630 , n2046 );
    or g3170 ( n305 , n6977 , n7952 );
    nor g3171 ( n12607 , n6993 , n9915 );
    nor g3172 ( n4235 , n8945 , n1859 );
    or g3173 ( n11382 , n6080 , n2953 );
    xnor g3174 ( n10005 , n6872 , n7751 );
    xnor g3175 ( n11441 , n4728 , n12275 );
    or g3176 ( n11879 , n3743 , n6922 );
    and g3177 ( n11531 , n2593 , n8497 );
    not g3178 ( n3998 , n2209 );
    xnor g3179 ( n8828 , n978 , n977 );
    xnor g3180 ( n4118 , n3372 , n5322 );
    xor g3181 ( n4367 , n8521 , n10445 );
    xnor g3182 ( n3572 , n3302 , n3771 );
    or g3183 ( n7376 , n11958 , n3903 );
    xnor g3184 ( n11897 , n6722 , n8318 );
    or g3185 ( n5988 , n3617 , n826 );
    not g3186 ( n5328 , n9606 );
    or g3187 ( n9793 , n215 , n939 );
    xnor g3188 ( n7779 , n2788 , n12627 );
    or g3189 ( n2556 , n9584 , n9521 );
    or g3190 ( n4627 , n12091 , n2348 );
    xnor g3191 ( n3871 , n11444 , n439 );
    xnor g3192 ( n6469 , n1646 , n11022 );
    nor g3193 ( n3164 , n12421 , n10063 );
    xnor g3194 ( n11888 , n12610 , n10283 );
    or g3195 ( n9326 , n2099 , n12535 );
    nor g3196 ( n12183 , n10100 , n9839 );
    not g3197 ( n351 , n400 );
    not g3198 ( n11860 , n3797 );
    or g3199 ( n5537 , n3746 , n12899 );
    and g3200 ( n2603 , n6027 , n2250 );
    not g3201 ( n9077 , n12952 );
    nor g3202 ( n3702 , n7491 , n10470 );
    or g3203 ( n3271 , n10663 , n8937 );
    or g3204 ( n11290 , n6939 , n208 );
    or g3205 ( n11974 , n8203 , n10722 );
    nor g3206 ( n9750 , n7667 , n9348 );
    xnor g3207 ( n7162 , n3404 , n12828 );
    or g3208 ( n3374 , n1699 , n530 );
    or g3209 ( n8353 , n10835 , n12771 );
    or g3210 ( n3032 , n9048 , n5993 );
    xnor g3211 ( n12854 , n2729 , n647 );
    or g3212 ( n6053 , n5530 , n7928 );
    xnor g3213 ( n11373 , n9084 , n9478 );
    or g3214 ( n4303 , n4059 , n1162 );
    nor g3215 ( n2341 , n3376 , n12134 );
    nor g3216 ( n3135 , n7542 , n12896 );
    not g3217 ( n4498 , n5240 );
    and g3218 ( n4894 , n5779 , n10102 );
    and g3219 ( n473 , n5674 , n11330 );
    xnor g3220 ( n12230 , n7493 , n8075 );
    not g3221 ( n10939 , n3424 );
    or g3222 ( n10269 , n7116 , n2815 );
    or g3223 ( n9306 , n2292 , n662 );
    xnor g3224 ( n4395 , n5364 , n12595 );
    or g3225 ( n588 , n6718 , n8643 );
    not g3226 ( n12859 , n4325 );
    and g3227 ( n10830 , n5967 , n3028 );
    or g3228 ( n9444 , n994 , n1455 );
    not g3229 ( n4474 , n9763 );
    and g3230 ( n7948 , n5441 , n1862 );
    nor g3231 ( n6017 , n3577 , n46 );
    and g3232 ( n7654 , n12310 , n9430 );
    and g3233 ( n1121 , n3133 , n10313 );
    not g3234 ( n10561 , n3769 );
    xnor g3235 ( n6964 , n8547 , n4020 );
    nor g3236 ( n6401 , n7779 , n10248 );
    not g3237 ( n3903 , n6126 );
    xnor g3238 ( n10303 , n12436 , n12389 );
    nor g3239 ( n12635 , n7170 , n9038 );
    nor g3240 ( n9935 , n1537 , n8188 );
    or g3241 ( n2037 , n7313 , n3640 );
    xnor g3242 ( n10651 , n10423 , n4517 );
    or g3243 ( n8441 , n2686 , n10618 );
    and g3244 ( n11273 , n8545 , n12783 );
    not g3245 ( n3924 , n8665 );
    and g3246 ( n819 , n11744 , n2222 );
    and g3247 ( n1472 , n10761 , n3234 );
    or g3248 ( n7629 , n3984 , n3902 );
    not g3249 ( n4014 , n2106 );
    or g3250 ( n3220 , n5116 , n11361 );
    and g3251 ( n3470 , n4299 , n5698 );
    xnor g3252 ( n3122 , n7620 , n1181 );
    not g3253 ( n3658 , n6631 );
    nor g3254 ( n8826 , n3221 , n3314 );
    xnor g3255 ( n11957 , n9162 , n7106 );
    or g3256 ( n2733 , n12818 , n541 );
    or g3257 ( n10266 , n5138 , n8471 );
    not g3258 ( n6084 , n8065 );
    not g3259 ( n9607 , n4659 );
    xnor g3260 ( n2316 , n11439 , n1609 );
    xnor g3261 ( n3471 , n7335 , n8466 );
    xnor g3262 ( n12944 , n4246 , n4265 );
    and g3263 ( n6165 , n8451 , n5430 );
    and g3264 ( n1264 , n12079 , n1704 );
    and g3265 ( n8225 , n5515 , n6683 );
    nor g3266 ( n9286 , n10560 , n5029 );
    or g3267 ( n11 , n4628 , n8259 );
    xnor g3268 ( n10785 , n9844 , n9225 );
    or g3269 ( n357 , n7283 , n7341 );
    and g3270 ( n592 , n9990 , n2840 );
    xnor g3271 ( n495 , n602 , n10024 );
    xnor g3272 ( n2458 , n10289 , n6679 );
    or g3273 ( n633 , n9554 , n8507 );
    xnor g3274 ( n3049 , n12008 , n5555 );
    not g3275 ( n209 , n7936 );
    xnor g3276 ( n833 , n3220 , n5675 );
    not g3277 ( n10442 , n2826 );
    xnor g3278 ( n1986 , n5571 , n537 );
    xnor g3279 ( n57 , n2950 , n7252 );
    and g3280 ( n3673 , n1623 , n7323 );
    or g3281 ( n9541 , n9370 , n1546 );
    or g3282 ( n5416 , n6256 , n7489 );
    and g3283 ( n5815 , n9107 , n2986 );
    not g3284 ( n10729 , n4468 );
    nor g3285 ( n18 , n4514 , n9659 );
    or g3286 ( n11832 , n10945 , n7318 );
    nor g3287 ( n3563 , n5101 , n9206 );
    xnor g3288 ( n7210 , n8273 , n4909 );
    or g3289 ( n2319 , n2217 , n6922 );
    or g3290 ( n7088 , n8870 , n6513 );
    or g3291 ( n10012 , n9170 , n6389 );
    or g3292 ( n11769 , n1075 , n8013 );
    xnor g3293 ( n4151 , n6050 , n3424 );
    and g3294 ( n5368 , n309 , n8529 );
    xnor g3295 ( n7042 , n11443 , n11237 );
    or g3296 ( n5031 , n6718 , n28 );
    not g3297 ( n3760 , n3001 );
    or g3298 ( n12527 , n636 , n8109 );
    xnor g3299 ( n10699 , n3428 , n1166 );
    not g3300 ( n1794 , n11154 );
    nor g3301 ( n6190 , n832 , n3178 );
    and g3302 ( n2684 , n4332 , n9232 );
    or g3303 ( n10199 , n5530 , n4818 );
    xnor g3304 ( n12866 , n8045 , n7557 );
    or g3305 ( n929 , n8127 , n12843 );
    xnor g3306 ( n8658 , n5415 , n4248 );
    nor g3307 ( n2179 , n9064 , n3185 );
    or g3308 ( n1581 , n3976 , n12059 );
    xnor g3309 ( n6711 , n5733 , n1237 );
    not g3310 ( n4636 , n313 );
    not g3311 ( n8280 , n8281 );
    or g3312 ( n2921 , n6948 , n8357 );
    or g3313 ( n10805 , n11061 , n9759 );
    nor g3314 ( n1527 , n6151 , n11219 );
    not g3315 ( n6141 , n6330 );
    and g3316 ( n5424 , n7273 , n5985 );
    and g3317 ( n11792 , n6072 , n891 );
    or g3318 ( n5938 , n3042 , n2965 );
    xnor g3319 ( n6646 , n5865 , n8480 );
    or g3320 ( n276 , n3127 , n5497 );
    xnor g3321 ( n9575 , n1215 , n5055 );
    xnor g3322 ( n9456 , n6516 , n9533 );
    or g3323 ( n2491 , n582 , n11014 );
    xnor g3324 ( n715 , n12912 , n8916 );
    xnor g3325 ( n4372 , n10776 , n4809 );
    or g3326 ( n3078 , n989 , n2358 );
    or g3327 ( n6660 , n8187 , n1546 );
    xnor g3328 ( n5358 , n4917 , n5870 );
    xnor g3329 ( n12851 , n11397 , n5821 );
    xnor g3330 ( n11208 , n2395 , n8893 );
    and g3331 ( n3786 , n5989 , n6704 );
    or g3332 ( n10315 , n11026 , n1509 );
    or g3333 ( n11985 , n3324 , n12771 );
    xnor g3334 ( n845 , n5244 , n5443 );
    or g3335 ( n7865 , n6457 , n12627 );
    and g3336 ( n12448 , n8748 , n4814 );
    or g3337 ( n9287 , n8054 , n3524 );
    and g3338 ( n876 , n11527 , n8072 );
    and g3339 ( n2913 , n4862 , n5230 );
    and g3340 ( n1087 , n9212 , n9932 );
    or g3341 ( n12171 , n5473 , n11792 );
    xnor g3342 ( n11164 , n9910 , n4795 );
    and g3343 ( n3507 , n1695 , n8066 );
    not g3344 ( n1825 , n1697 );
    not g3345 ( n309 , n12348 );
    not g3346 ( n4912 , n9026 );
    or g3347 ( n11764 , n9432 , n7226 );
    and g3348 ( n3088 , n8649 , n9624 );
    xnor g3349 ( n7614 , n5485 , n5083 );
    or g3350 ( n898 , n7701 , n10486 );
    xnor g3351 ( n1662 , n5161 , n4915 );
    or g3352 ( n6293 , n9389 , n11827 );
    and g3353 ( n9598 , n9698 , n665 );
    not g3354 ( n11994 , n4099 );
    and g3355 ( n8193 , n8554 , n10561 );
    or g3356 ( n10862 , n8326 , n10044 );
    xnor g3357 ( n5213 , n438 , n12631 );
    xnor g3358 ( n5963 , n9819 , n10795 );
    xnor g3359 ( n381 , n3941 , n11054 );
    xnor g3360 ( n12836 , n5247 , n9020 );
    xnor g3361 ( n11301 , n4034 , n400 );
    or g3362 ( n4657 , n7687 , n2352 );
    xnor g3363 ( n8884 , n8544 , n5051 );
    nor g3364 ( n10433 , n4500 , n1483 );
    xnor g3365 ( n3880 , n346 , n7721 );
    and g3366 ( n2078 , n1909 , n1773 );
    nor g3367 ( n9249 , n2444 , n1176 );
    not g3368 ( n1442 , n7909 );
    xnor g3369 ( n9253 , n2918 , n10425 );
    and g3370 ( n8097 , n2082 , n7007 );
    nor g3371 ( n205 , n6966 , n11981 );
    not g3372 ( n7336 , n10751 );
    or g3373 ( n637 , n10601 , n3576 );
    or g3374 ( n12877 , n10196 , n8830 );
    or g3375 ( n5430 , n8110 , n2767 );
    and g3376 ( n5912 , n7715 , n3883 );
    or g3377 ( n8564 , n11457 , n4240 );
    not g3378 ( n11122 , n2433 );
    not g3379 ( n12543 , n10998 );
    or g3380 ( n4819 , n4778 , n10854 );
    or g3381 ( n6130 , n8305 , n1667 );
    or g3382 ( n6096 , n9170 , n1162 );
    and g3383 ( n9437 , n6687 , n2879 );
    or g3384 ( n3951 , n3609 , n11286 );
    or g3385 ( n7037 , n3127 , n7424 );
    xnor g3386 ( n9605 , n3474 , n8780 );
    xnor g3387 ( n7000 , n11233 , n3489 );
    nor g3388 ( n7070 , n9179 , n9479 );
    xnor g3389 ( n9847 , n8163 , n4448 );
    xnor g3390 ( n4640 , n9846 , n5409 );
    or g3391 ( n9301 , n7391 , n7341 );
    or g3392 ( n12845 , n11547 , n6832 );
    xnor g3393 ( n2281 , n11390 , n3431 );
    or g3394 ( n167 , n8345 , n2635 );
    not g3395 ( n1987 , n7505 );
    xnor g3396 ( n5124 , n3864 , n10234 );
    not g3397 ( n5765 , n11153 );
    nor g3398 ( n4662 , n4135 , n5339 );
    and g3399 ( n1872 , n2924 , n2141 );
    xnor g3400 ( n3701 , n10332 , n9484 );
    not g3401 ( n3580 , n9194 );
    xnor g3402 ( n2115 , n4480 , n7123 );
    and g3403 ( n4199 , n1972 , n3977 );
    xnor g3404 ( n860 , n469 , n7349 );
    and g3405 ( n12540 , n2537 , n151 );
    not g3406 ( n5616 , n11053 );
    or g3407 ( n12495 , n8792 , n7972 );
    xnor g3408 ( n6421 , n11155 , n3574 );
    xnor g3409 ( n5545 , n10359 , n8424 );
    or g3410 ( n1111 , n3743 , n3606 );
    or g3411 ( n5562 , n12853 , n8740 );
    not g3412 ( n10170 , n10034 );
    xnor g3413 ( n3043 , n2060 , n6131 );
    not g3414 ( n2612 , n12619 );
    or g3415 ( n4625 , n7977 , n755 );
    not g3416 ( n6373 , n11892 );
    or g3417 ( n1246 , n8221 , n11268 );
    and g3418 ( n4833 , n12683 , n6552 );
    not g3419 ( n8354 , n3616 );
    and g3420 ( n2219 , n5708 , n12892 );
    xnor g3421 ( n2908 , n5819 , n1697 );
    xnor g3422 ( n7227 , n4170 , n10599 );
    and g3423 ( n709 , n6628 , n11372 );
    and g3424 ( n6222 , n12087 , n4267 );
    xnor g3425 ( n4857 , n3885 , n11729 );
    not g3426 ( n2202 , n9275 );
    xnor g3427 ( n7193 , n1505 , n4118 );
    xnor g3428 ( n11156 , n4021 , n10654 );
    nor g3429 ( n9044 , n7295 , n2785 );
    nor g3430 ( n9244 , n7316 , n9090 );
    not g3431 ( n8429 , n7824 );
    or g3432 ( n2993 , n12186 , n2815 );
    xnor g3433 ( n2593 , n10028 , n4651 );
    not g3434 ( n2557 , n9982 );
    and g3435 ( n4568 , n10852 , n12019 );
    or g3436 ( n3672 , n24 , n7334 );
    or g3437 ( n5292 , n6718 , n795 );
    or g3438 ( n7352 , n4100 , n9385 );
    not g3439 ( n5042 , n9307 );
    or g3440 ( n1326 , n11552 , n4642 );
    or g3441 ( n5706 , n3820 , n8643 );
    and g3442 ( n1190 , n7788 , n11654 );
    or g3443 ( n4065 , n5858 , n1455 );
    or g3444 ( n6552 , n2478 , n2387 );
    xnor g3445 ( n93 , n6767 , n1508 );
    or g3446 ( n4360 , n4498 , n1455 );
    xnor g3447 ( n6273 , n10382 , n11167 );
    and g3448 ( n5081 , n5964 , n11662 );
    and g3449 ( n9982 , n7124 , n4307 );
    xnor g3450 ( n7408 , n12272 , n6950 );
    and g3451 ( n11730 , n1757 , n303 );
    nor g3452 ( n6805 , n8532 , n442 );
    xnor g3453 ( n10090 , n6995 , n9305 );
    or g3454 ( n12273 , n4856 , n10610 );
    xnor g3455 ( n6356 , n913 , n8493 );
    xor g3456 ( n4442 , n10647 , n10009 );
    and g3457 ( n2428 , n1224 , n8422 );
    and g3458 ( n11463 , n10078 , n8652 );
    xnor g3459 ( n3711 , n6962 , n7049 );
    and g3460 ( n8204 , n6776 , n12145 );
    or g3461 ( n4859 , n2099 , n9586 );
    not g3462 ( n11753 , n3541 );
    or g3463 ( n10667 , n2217 , n8745 );
    xnor g3464 ( n10665 , n8197 , n1098 );
    not g3465 ( n380 , n9698 );
    or g3466 ( n8321 , n10879 , n7424 );
    not g3467 ( n4405 , n4070 );
    and g3468 ( n6802 , n9806 , n8579 );
    nor g3469 ( n10420 , n3365 , n5811 );
    nor g3470 ( n9799 , n9669 , n12196 );
    xnor g3471 ( n9145 , n1622 , n10189 );
    and g3472 ( n1813 , n2102 , n517 );
    xnor g3473 ( n1787 , n7663 , n11886 );
    and g3474 ( n11666 , n6244 , n8180 );
    or g3475 ( n7028 , n2854 , n1961 );
    xor g3476 ( n397 , n649 , n8270 );
    not g3477 ( n12220 , n6553 );
    or g3478 ( n3378 , n4272 , n11833 );
    not g3479 ( n88 , n1795 );
    xnor g3480 ( n9094 , n7254 , n11190 );
    or g3481 ( n4418 , n9528 , n10054 );
    and g3482 ( n3665 , n3819 , n2966 );
    nor g3483 ( n11113 , n4060 , n2225 );
    not g3484 ( n9083 , n4463 );
    not g3485 ( n10553 , n987 );
    xnor g3486 ( n12795 , n1560 , n12697 );
    and g3487 ( n12275 , n2414 , n1920 );
    or g3488 ( n10089 , n8959 , n11122 );
    or g3489 ( n11076 , n12853 , n3224 );
    nor g3490 ( n12062 , n4273 , n11934 );
    not g3491 ( n3361 , n9627 );
    xnor g3492 ( n2021 , n3757 , n10363 );
    and g3493 ( n4976 , n632 , n4881 );
    nor g3494 ( n12685 , n2230 , n7302 );
    xnor g3495 ( n7984 , n5332 , n12952 );
    xnor g3496 ( n6889 , n5380 , n4305 );
    and g3497 ( n3074 , n6509 , n2657 );
    or g3498 ( n4146 , n2872 , n2815 );
    or g3499 ( n5179 , n752 , n11122 );
    xnor g3500 ( n5137 , n7418 , n3061 );
    not g3501 ( n9736 , n5931 );
    or g3502 ( n4202 , n10196 , n9568 );
    or g3503 ( n11928 , n752 , n7395 );
    xnor g3504 ( n5144 , n9 , n12486 );
    not g3505 ( n7129 , n11307 );
    xnor g3506 ( n5702 , n9340 , n263 );
    or g3507 ( n4503 , n9945 , n11486 );
    nor g3508 ( n9097 , n4074 , n5104 );
    or g3509 ( n3750 , n10741 , n10149 );
    and g3510 ( n6364 , n5860 , n10898 );
    xnor g3511 ( n9695 , n3508 , n12096 );
    or g3512 ( n9260 , n11719 , n4400 );
    xnor g3513 ( n815 , n7062 , n145 );
    xnor g3514 ( n2636 , n2098 , n6959 );
    xnor g3515 ( n12762 , n1458 , n3942 );
    nor g3516 ( n6229 , n3228 , n2603 );
    xnor g3517 ( n12563 , n6620 , n11660 );
    or g3518 ( n418 , n5809 , n9188 );
    xnor g3519 ( n11686 , n9905 , n10792 );
    xnor g3520 ( n9537 , n861 , n9545 );
    and g3521 ( n2928 , n2559 , n502 );
    and g3522 ( n15 , n10615 , n4699 );
    xnor g3523 ( n2480 , n4349 , n4927 );
    or g3524 ( n6043 , n5061 , n11720 );
    or g3525 ( n6325 , n3265 , n1454 );
    and g3526 ( n2022 , n8137 , n7076 );
    and g3527 ( n8525 , n2833 , n553 );
    xnor g3528 ( n44 , n12223 , n4389 );
    xnor g3529 ( n9986 , n3464 , n8805 );
    xnor g3530 ( n2255 , n7984 , n6362 );
    nor g3531 ( n10137 , n3233 , n4402 );
    or g3532 ( n10141 , n8552 , n9586 );
    and g3533 ( n1889 , n5084 , n562 );
    xnor g3534 ( n10954 , n9872 , n6941 );
    or g3535 ( n376 , n959 , n5155 );
    or g3536 ( n12344 , n2969 , n11072 );
    or g3537 ( n1009 , n5575 , n2232 );
    or g3538 ( n3491 , n7391 , n4242 );
    xor g3539 ( n5641 , n1548 , n6838 );
    or g3540 ( n6345 , n4178 , n1751 );
    or g3541 ( n10377 , n2099 , n12446 );
    or g3542 ( n5542 , n752 , n184 );
    not g3543 ( n2866 , n6085 );
    xnor g3544 ( n9390 , n5476 , n8360 );
    or g3545 ( n1993 , n11749 , n4165 );
    and g3546 ( n6160 , n11181 , n4268 );
    nor g3547 ( n8212 , n12537 , n11978 );
    or g3548 ( n4178 , n239 , n8788 );
    xnor g3549 ( n10720 , n1059 , n10875 );
    or g3550 ( n11953 , n5032 , n760 );
    nor g3551 ( n11684 , n489 , n10184 );
    xnor g3552 ( n12059 , n366 , n2035 );
    or g3553 ( n8560 , n7539 , n1328 );
    xnor g3554 ( n2003 , n11173 , n8603 );
    not g3555 ( n9743 , n1853 );
    or g3556 ( n3486 , n12033 , n6781 );
    and g3557 ( n11947 , n584 , n8887 );
    not g3558 ( n12687 , n1166 );
    not g3559 ( n4565 , n9993 );
    xnor g3560 ( n12402 , n6125 , n2867 );
    and g3561 ( n4337 , n12837 , n12554 );
    or g3562 ( n396 , n12361 , n3421 );
    or g3563 ( n164 , n11856 , n6911 );
    nor g3564 ( n1290 , n12859 , n2412 );
    and g3565 ( n3070 , n6147 , n9876 );
    nor g3566 ( n2510 , n6551 , n2086 );
    xnor g3567 ( n7020 , n8553 , n5073 );
    or g3568 ( n5228 , n10833 , n7761 );
    nor g3569 ( n1568 , n1424 , n8707 );
    xnor g3570 ( n4971 , n12818 , n11461 );
    xnor g3571 ( n7528 , n11414 , n11375 );
    not g3572 ( n12312 , n7390 );
    not g3573 ( n5013 , n1688 );
    or g3574 ( n6177 , n1699 , n7928 );
    and g3575 ( n6997 , n6795 , n11424 );
    or g3576 ( n8961 , n11421 , n6212 );
    not g3577 ( n10108 , n9080 );
    or g3578 ( n5559 , n2099 , n7136 );
    and g3579 ( n2650 , n5198 , n9111 );
    and g3580 ( n3983 , n839 , n69 );
    not g3581 ( n9188 , n2558 );
    or g3582 ( n8481 , n8026 , n6197 );
    xnor g3583 ( n7831 , n8022 , n724 );
    xnor g3584 ( n2516 , n8449 , n4758 );
    xnor g3585 ( n11824 , n1038 , n3466 );
    xnor g3586 ( n3762 , n11559 , n6978 );
    or g3587 ( n7669 , n5902 , n3911 );
    xnor g3588 ( n7333 , n7021 , n10726 );
    xnor g3589 ( n4688 , n8557 , n7275 );
    or g3590 ( n6175 , n6977 , n7876 );
    xnor g3591 ( n7269 , n4963 , n9362 );
    and g3592 ( n491 , n11200 , n9393 );
    or g3593 ( n1642 , n11958 , n7425 );
    or g3594 ( n5864 , n8354 , n8740 );
    and g3595 ( n514 , n11013 , n1346 );
    not g3596 ( n1780 , n8600 );
    or g3597 ( n6777 , n5355 , n7246 );
    or g3598 ( n10710 , n3324 , n795 );
    xnor g3599 ( n10637 , n9395 , n10386 );
    xnor g3600 ( n11644 , n5438 , n1856 );
    or g3601 ( n3190 , n10882 , n9665 );
    and g3602 ( n12789 , n9433 , n11196 );
    or g3603 ( n8269 , n683 , n12834 );
    and g3604 ( n5335 , n676 , n4331 );
    or g3605 ( n1534 , n8387 , n12856 );
    nor g3606 ( n653 , n1181 , n12808 );
    not g3607 ( n12869 , n4331 );
    xnor g3608 ( n3112 , n987 , n6367 );
    and g3609 ( n6335 , n2505 , n8388 );
    or g3610 ( n9777 , n7176 , n506 );
    or g3611 ( n1126 , n7391 , n10066 );
    or g3612 ( n8589 , n11584 , n4156 );
    or g3613 ( n11634 , n4311 , n2572 );
    and g3614 ( n8307 , n10522 , n2943 );
    and g3615 ( n7295 , n1387 , n2954 );
    not g3616 ( n6775 , n8966 );
    not g3617 ( n6808 , n10658 );
    xnor g3618 ( n1213 , n2519 , n4673 );
    xnor g3619 ( n12234 , n53 , n7541 );
    or g3620 ( n2675 , n5190 , n6371 );
    xnor g3621 ( n11562 , n9381 , n7277 );
    and g3622 ( n8821 , n298 , n8746 );
    xnor g3623 ( n7603 , n12730 , n3123 );
    nor g3624 ( n9759 , n9615 , n5253 );
    nor g3625 ( n4739 , n4451 , n1852 );
    not g3626 ( n6491 , n2721 );
    or g3627 ( n8579 , n8354 , n9188 );
    or g3628 ( n4015 , n11266 , n8286 );
    nor g3629 ( n9554 , n10658 , n2513 );
    xnor g3630 ( n6565 , n4049 , n11554 );
    and g3631 ( n73 , n7884 , n1930 );
    or g3632 ( n4702 , n7470 , n1286 );
    and g3633 ( n6800 , n1311 , n799 );
    xnor g3634 ( n6250 , n6285 , n7515 );
    or g3635 ( n7457 , n2099 , n12883 );
    or g3636 ( n1701 , n7154 , n10837 );
    and g3637 ( n2211 , n8727 , n6756 );
    not g3638 ( n9106 , n253 );
    or g3639 ( n6004 , n5575 , n2754 );
    not g3640 ( n7260 , n5500 );
    or g3641 ( n928 , n10750 , n8740 );
    xnor g3642 ( n7135 , n5137 , n7340 );
    or g3643 ( n4476 , n7709 , n12771 );
    xnor g3644 ( n2064 , n3284 , n5841 );
    or g3645 ( n8395 , n5915 , n6513 );
    and g3646 ( n935 , n4727 , n4140 );
    xnor g3647 ( n6155 , n10843 , n1169 );
    nor g3648 ( n5310 , n1479 , n1088 );
    or g3649 ( n8227 , n3743 , n4864 );
    or g3650 ( n7663 , n2099 , n8259 );
    or g3651 ( n415 , n3776 , n7665 );
    and g3652 ( n7989 , n4576 , n7365 );
    and g3653 ( n2180 , n1684 , n3408 );
    xnor g3654 ( n3656 , n11556 , n6173 );
    and g3655 ( n3158 , n6654 , n8578 );
    xnor g3656 ( n11760 , n12037 , n8968 );
    and g3657 ( n2364 , n8476 , n5645 );
    or g3658 ( n9645 , n5179 , n8417 );
    nor g3659 ( n8873 , n548 , n2184 );
    or g3660 ( n574 , n7709 , n9521 );
    xnor g3661 ( n3206 , n6518 , n9790 );
    xnor g3662 ( n663 , n9678 , n9384 );
    or g3663 ( n3927 , n8443 , n12769 );
    nor g3664 ( n4142 , n11400 , n7590 );
    xnor g3665 ( n402 , n1299 , n11634 );
    xnor g3666 ( n8466 , n6548 , n3910 );
    and g3667 ( n11987 , n8441 , n10645 );
    xnor g3668 ( n1611 , n3213 , n9694 );
    and g3669 ( n11051 , n11764 , n7533 );
    and g3670 ( n757 , n7902 , n10675 );
    and g3671 ( n2090 , n3145 , n1267 );
    xnor g3672 ( n10067 , n8827 , n364 );
    xnor g3673 ( n1365 , n8652 , n5293 );
    xnor g3674 ( n11795 , n9755 , n10274 );
    nor g3675 ( n5246 , n9227 , n11615 );
    nor g3676 ( n10307 , n1142 , n5933 );
    and g3677 ( n5700 , n12659 , n6846 );
    or g3678 ( n5571 , n6577 , n3468 );
    or g3679 ( n2427 , n6577 , n3903 );
    nor g3680 ( n5620 , n4719 , n5723 );
    not g3681 ( n10066 , n6038 );
    or g3682 ( n12914 , n989 , n561 );
    and g3683 ( n1863 , n9465 , n3003 );
    xnor g3684 ( n8242 , n5118 , n4081 );
    or g3685 ( n1593 , n257 , n5333 );
    xnor g3686 ( n10490 , n11400 , n4691 );
    or g3687 ( n4509 , n12177 , n12386 );
    and g3688 ( n5418 , n2564 , n9956 );
    xnor g3689 ( n1573 , n49 , n8775 );
    xnor g3690 ( n7183 , n4699 , n7565 );
    or g3691 ( n3349 , n5470 , n4672 );
    xnor g3692 ( n5037 , n4799 , n4607 );
    or g3693 ( n11773 , n6857 , n4544 );
    xnor g3694 ( n6094 , n9615 , n10981 );
    and g3695 ( n1288 , n9376 , n11160 );
    xnor g3696 ( n3466 , n10530 , n3470 );
    or g3697 ( n10086 , n2832 , n12843 );
    or g3698 ( n9369 , n9170 , n7881 );
    xnor g3699 ( n10617 , n623 , n5157 );
    or g3700 ( n11546 , n9492 , n4420 );
    and g3701 ( n2519 , n10534 , n12546 );
    xnor g3702 ( n1687 , n11231 , n7553 );
    xnor g3703 ( n6895 , n7752 , n9868 );
    xnor g3704 ( n3476 , n5242 , n79 );
    and g3705 ( n6712 , n5491 , n7743 );
    xnor g3706 ( n7142 , n762 , n6312 );
    not g3707 ( n8340 , n203 );
    xnor g3708 ( n10378 , n8912 , n7830 );
    and g3709 ( n3420 , n9895 , n1832 );
    xnor g3710 ( n3533 , n3880 , n9498 );
    not g3711 ( n1840 , n5820 );
    and g3712 ( n1076 , n3291 , n8686 );
    not g3713 ( n8240 , n2680 );
    xnor g3714 ( n11908 , n3038 , n1030 );
    or g3715 ( n6145 , n8959 , n12816 );
    xnor g3716 ( n2955 , n12939 , n6858 );
    not g3717 ( n6759 , n8850 );
    and g3718 ( n2074 , n7822 , n5165 );
    nor g3719 ( n4530 , n11248 , n7525 );
    or g3720 ( n5791 , n5530 , n4249 );
    not g3721 ( n3224 , n1564 );
    and g3722 ( n11943 , n8387 , n12856 );
    nor g3723 ( n12245 , n12367 , n11600 );
    xnor g3724 ( n12926 , n5564 , n7451 );
    xnor g3725 ( n10560 , n4058 , n1554 );
    xnor g3726 ( n7057 , n3016 , n5356 );
    xnor g3727 ( n1949 , n312 , n11600 );
    or g3728 ( n2989 , n10922 , n8021 );
    and g3729 ( n8091 , n10928 , n4141 );
    xnor g3730 ( n3626 , n1786 , n10971 );
    xnor g3731 ( n4279 , n7603 , n11951 );
    nor g3732 ( n1435 , n5346 , n9704 );
    or g3733 ( n3485 , n3765 , n3158 );
    nor g3734 ( n2774 , n7186 , n11809 );
    and g3735 ( n9355 , n8679 , n1360 );
    nor g3736 ( n997 , n8646 , n7314 );
    or g3737 ( n7213 , n11569 , n4115 );
    or g3738 ( n5254 , n618 , n7139 );
    xnor g3739 ( n6355 , n6625 , n7625 );
    and g3740 ( n7525 , n4442 , n4110 );
    and g3741 ( n8222 , n3024 , n7596 );
    not g3742 ( n12909 , n9819 );
    xnor g3743 ( n572 , n12661 , n1211 );
    and g3744 ( n1113 , n12643 , n4537 );
    not g3745 ( n8720 , n11987 );
    xnor g3746 ( n6477 , n9657 , n7969 );
    or g3747 ( n12010 , n8127 , n1851 );
    xnor g3748 ( n1373 , n2150 , n5723 );
    xnor g3749 ( n2617 , n9825 , n9776 );
    or g3750 ( n8988 , n1151 , n4573 );
    xnor g3751 ( n7335 , n7915 , n11435 );
    not g3752 ( n8214 , n9810 );
    xnor g3753 ( n4959 , n7001 , n12897 );
    or g3754 ( n494 , n6718 , n7506 );
    or g3755 ( n12683 , n7831 , n10979 );
    or g3756 ( n10064 , n10018 , n10021 );
    xnor g3757 ( n10563 , n12460 , n360 );
    xnor g3758 ( n2062 , n12930 , n9350 );
    and g3759 ( n11127 , n3131 , n10813 );
    nor g3760 ( n10161 , n1975 , n11606 );
    not g3761 ( n4604 , n4437 );
    or g3762 ( n6204 , n191 , n7703 );
    nor g3763 ( n10796 , n10004 , n7968 );
    or g3764 ( n3024 , n868 , n8323 );
    xnor g3765 ( n6060 , n3791 , n11806 );
    xnor g3766 ( n10526 , n1681 , n7048 );
    xnor g3767 ( n9057 , n4063 , n179 );
    nor g3768 ( n297 , n1830 , n3860 );
    not g3769 ( n1983 , n9567 );
    xnor g3770 ( n8079 , n9928 , n2501 );
    or g3771 ( n5661 , n8187 , n11827 );
    or g3772 ( n6784 , n1315 , n2211 );
    nor g3773 ( n10446 , n1439 , n9427 );
    or g3774 ( n5195 , n3367 , n3056 );
    not g3775 ( n6054 , n6335 );
    xnor g3776 ( n10104 , n8198 , n4403 );
    nor g3777 ( n11697 , n5574 , n9133 );
    or g3778 ( n11695 , n3617 , n4913 );
    or g3779 ( n10363 , n11923 , n1509 );
    xnor g3780 ( n11669 , n7280 , n11909 );
    and g3781 ( n6032 , n12413 , n8866 );
    not g3782 ( n4154 , n12702 );
    and g3783 ( n5597 , n2638 , n8358 );
    not g3784 ( n9952 , n11459 );
    and g3785 ( n6707 , n4560 , n11334 );
    xnor g3786 ( n5998 , n10710 , n10083 );
    xnor g3787 ( n696 , n8174 , n12937 );
    xnor g3788 ( n1223 , n1354 , n9167 );
    xnor g3789 ( n5495 , n5048 , n1159 );
    xnor g3790 ( n707 , n11931 , n4008 );
    and g3791 ( n557 , n12346 , n12083 );
    xnor g3792 ( n11309 , n1352 , n7851 );
    or g3793 ( n5501 , n10142 , n8524 );
    not g3794 ( n10988 , n588 );
    xnor g3795 ( n2781 , n11279 , n11020 );
    not g3796 ( n8856 , n5665 );
    or g3797 ( n2938 , n10132 , n3476 );
    and g3798 ( n843 , n3608 , n3488 );
    or g3799 ( n4465 , n6977 , n2815 );
    xnor g3800 ( n8298 , n4135 , n8076 );
    or g3801 ( n10400 , n3470 , n9175 );
    and g3802 ( n2371 , n5089 , n10823 );
    and g3803 ( n3534 , n3614 , n8539 );
    xnor g3804 ( n7684 , n272 , n3095 );
    nor g3805 ( n4198 , n74 , n7776 );
    or g3806 ( n940 , n10339 , n826 );
    xnor g3807 ( n6487 , n3106 , n1759 );
    and g3808 ( n8838 , n11838 , n7344 );
    or g3809 ( n9395 , n3820 , n1509 );
    or g3810 ( n8761 , n7196 , n4087 );
    and g3811 ( n10622 , n8831 , n3918 );
    or g3812 ( n3328 , n6814 , n2929 );
    or g3813 ( n904 , n10750 , n10422 );
    or g3814 ( n7904 , n4674 , n9188 );
    nor g3815 ( n1778 , n10839 , n5248 );
    not g3816 ( n9632 , n2428 );
    nor g3817 ( n4589 , n1632 , n11730 );
    and g3818 ( n1907 , n8217 , n10941 );
    xnor g3819 ( n12934 , n11327 , n7000 );
    or g3820 ( n10936 , n12119 , n8957 );
    or g3821 ( n816 , n2099 , n3224 );
    xnor g3822 ( n12228 , n4435 , n10033 );
    not g3823 ( n9046 , n11230 );
    xnor g3824 ( n3592 , n6282 , n12279 );
    not g3825 ( n6667 , n7563 );
    xnor g3826 ( n7958 , n7873 , n9771 );
    or g3827 ( n5489 , n7998 , n4153 );
    and g3828 ( n5660 , n5886 , n770 );
    and g3829 ( n8487 , n6275 , n3907 );
    xnor g3830 ( n2690 , n8429 , n7326 );
    not g3831 ( n242 , n8526 );
    not g3832 ( n10234 , n3246 );
    and g3833 ( n10110 , n11490 , n1919 );
    xnor g3834 ( n6344 , n8194 , n4035 );
    and g3835 ( n8477 , n11153 , n7270 );
    or g3836 ( n7551 , n6577 , n6169 );
    or g3837 ( n4134 , n6053 , n5830 );
    xnor g3838 ( n9805 , n12496 , n5124 );
    or g3839 ( n8669 , n11005 , n11297 );
    or g3840 ( n5219 , n2099 , n8655 );
    or g3841 ( n12386 , n8959 , n6169 );
    xnor g3842 ( n5633 , n6350 , n11412 );
    not g3843 ( n7717 , n1882 );
    xnor g3844 ( n10034 , n8395 , n7863 );
    or g3845 ( n4535 , n10157 , n4642 );
    and g3846 ( n6955 , n5054 , n6300 );
    xnor g3847 ( n3294 , n8520 , n7815 );
    and g3848 ( n3212 , n11234 , n12522 );
    xnor g3849 ( n10166 , n2688 , n5315 );
    and g3850 ( n291 , n8194 , n4035 );
    nor g3851 ( n6779 , n5975 , n2362 );
    or g3852 ( n2254 , n1799 , n8544 );
    xnor g3853 ( n2005 , n9304 , n549 );
    or g3854 ( n9329 , n6544 , n6422 );
    or g3855 ( n7176 , n12119 , n9586 );
    xnor g3856 ( n9047 , n11934 , n4273 );
    and g3857 ( n12760 , n6941 , n6764 );
    xnor g3858 ( n7249 , n10153 , n8437 );
    not g3859 ( n918 , n9270 );
    or g3860 ( n5516 , n603 , n12688 );
    or g3861 ( n1145 , n1696 , n3102 );
    not g3862 ( n8414 , n4928 );
    or g3863 ( n10340 , n10732 , n476 );
    or g3864 ( n8499 , n9373 , n5502 );
    and g3865 ( n2962 , n6408 , n5787 );
    nor g3866 ( n6959 , n8141 , n12804 );
    and g3867 ( n5993 , n7108 , n12164 );
    and g3868 ( n5547 , n8411 , n4596 );
    or g3869 ( n4837 , n5398 , n3248 );
    or g3870 ( n2618 , n4911 , n7341 );
    xnor g3871 ( n11437 , n2138 , n723 );
    and g3872 ( n11220 , n585 , n4670 );
    nor g3873 ( n8795 , n9514 , n3751 );
    nor g3874 ( n154 , n9017 , n8199 );
    and g3875 ( n2943 , n6709 , n8356 );
    or g3876 ( n8587 , n11556 , n6173 );
    and g3877 ( n11247 , n3155 , n7213 );
    or g3878 ( n10594 , n4116 , n7188 );
    or g3879 ( n8431 , n11933 , n11322 );
    xnor g3880 ( n8270 , n6520 , n5991 );
    xnor g3881 ( n5756 , n6517 , n10246 );
    and g3882 ( n9215 , n8221 , n11268 );
    or g3883 ( n10754 , n3617 , n5468 );
    or g3884 ( n6227 , n11060 , n11247 );
    or g3885 ( n8814 , n10157 , n1509 );
    and g3886 ( n11243 , n9777 , n9309 );
    nor g3887 ( n10471 , n8518 , n5697 );
    xnor g3888 ( n9375 , n7758 , n793 );
    xnor g3889 ( n7182 , n4395 , n7923 );
    and g3890 ( n9808 , n6142 , n830 );
    xnor g3891 ( n3988 , n9197 , n12110 );
    and g3892 ( n12776 , n2564 , n2585 );
    not g3893 ( n2292 , n3817 );
    xnor g3894 ( n877 , n12178 , n1481 );
    or g3895 ( n5384 , n5355 , n1546 );
    xnor g3896 ( n461 , n2885 , n9715 );
    xnor g3897 ( n8250 , n359 , n9357 );
    not g3898 ( n130 , n2512 );
    xnor g3899 ( n1713 , n2365 , n932 );
    xnor g3900 ( n39 , n10152 , n1693 );
    and g3901 ( n3775 , n3992 , n11876 );
    xnor g3902 ( n536 , n5206 , n2311 );
    xnor g3903 ( n2443 , n2481 , n3504 );
    xnor g3904 ( n480 , n6039 , n10488 );
    xnor g3905 ( n11409 , n11076 , n7142 );
    not g3906 ( n11852 , n4990 );
    xnor g3907 ( n3092 , n10844 , n8471 );
    not g3908 ( n10891 , n9385 );
    xnor g3909 ( n5675 , n7268 , n1767 );
    and g3910 ( n5783 , n8336 , n9640 );
    xnor g3911 ( n3722 , n11352 , n12265 );
    not g3912 ( n3152 , n187 );
    nor g3913 ( n2065 , n3665 , n2452 );
    xnor g3914 ( n654 , n8282 , n12298 );
    nor g3915 ( n3737 , n11405 , n9285 );
    xnor g3916 ( n8061 , n1031 , n9297 );
    xnor g3917 ( n2526 , n10414 , n10369 );
    or g3918 ( n7311 , n10339 , n12535 );
    xnor g3919 ( n10537 , n4829 , n11301 );
    or g3920 ( n7327 , n2217 , n4527 );
    nor g3921 ( n2692 , n7835 , n8885 );
    xnor g3922 ( n6830 , n3108 , n6610 );
    or g3923 ( n354 , n636 , n6513 );
    not g3924 ( n836 , n5418 );
    not g3925 ( n4080 , n5841 );
    not g3926 ( n10386 , n7205 );
    and g3927 ( n8243 , n2792 , n5060 );
    not g3928 ( n2830 , n4017 );
    or g3929 ( n2750 , n6475 , n10867 );
    xnor g3930 ( n7852 , n3826 , n2613 );
    xnor g3931 ( n4072 , n6556 , n6007 );
    nor g3932 ( n7724 , n11128 , n558 );
    or g3933 ( n10614 , n6914 , n4447 );
    not g3934 ( n26 , n7922 );
    xnor g3935 ( n4577 , n985 , n5558 );
    or g3936 ( n11405 , n3324 , n9521 );
    or g3937 ( n6901 , n9792 , n7554 );
    nor g3938 ( n2407 , n1844 , n6094 );
    and g3939 ( n4824 , n11567 , n4209 );
    xnor g3940 ( n4594 , n5001 , n6787 );
    xnor g3941 ( n9866 , n2329 , n8000 );
    or g3942 ( n9758 , n12155 , n6473 );
    or g3943 ( n5989 , n10835 , n4875 );
    or g3944 ( n9687 , n9529 , n7950 );
    not g3945 ( n7601 , n1905 );
    xnor g3946 ( n1274 , n10790 , n11235 );
    and g3947 ( n12244 , n982 , n8230 );
    or g3948 ( n1749 , n10129 , n11946 );
    and g3949 ( n10308 , n4238 , n6304 );
    xnor g3950 ( n11583 , n1459 , n1984 );
    xnor g3951 ( n1771 , n961 , n1359 );
    not g3952 ( n2023 , n8410 );
    and g3953 ( n12547 , n8309 , n10441 );
    xnor g3954 ( n6605 , n8412 , n3429 );
    and g3955 ( n2649 , n10874 , n1300 );
    and g3956 ( n5551 , n8229 , n1276 );
    nor g3957 ( n2911 , n4442 , n4110 );
    and g3958 ( n7668 , n137 , n7610 );
    not g3959 ( n3621 , n4520 );
    xnor g3960 ( n8447 , n4357 , n10299 );
    xnor g3961 ( n4109 , n240 , n1076 );
    xnor g3962 ( n10140 , n5044 , n7639 );
    or g3963 ( n6310 , n10750 , n12446 );
    nor g3964 ( n12509 , n7599 , n8910 );
    xnor g3965 ( n4272 , n2304 , n4839 );
    not g3966 ( n8201 , n11363 );
    xnor g3967 ( n6570 , n12055 , n8246 );
    xnor g3968 ( n2486 , n2838 , n6164 );
    xnor g3969 ( n72 , n10015 , n12517 );
    not g3970 ( n316 , n985 );
    not g3971 ( n2715 , n10443 );
    nor g3972 ( n11218 , n9453 , n9646 );
    and g3973 ( n888 , n610 , n469 );
    not g3974 ( n12585 , n11784 );
    and g3975 ( n9440 , n399 , n7949 );
    and g3976 ( n8349 , n1960 , n1019 );
    not g3977 ( n4376 , n10974 );
    xnor g3978 ( n4417 , n12432 , n6162 );
    xnor g3979 ( n712 , n644 , n9966 );
    not g3980 ( n8185 , n6935 );
    xnor g3981 ( n6083 , n8481 , n1048 );
    and g3982 ( n2006 , n10893 , n9121 );
    or g3983 ( n6237 , n9373 , n4474 );
    or g3984 ( n10487 , n2456 , n12754 );
    and g3985 ( n6559 , n4079 , n150 );
    nor g3986 ( n1788 , n6607 , n10753 );
    or g3987 ( n7027 , n10750 , n12535 );
    xnor g3988 ( n2613 , n685 , n12191 );
    not g3989 ( n5638 , n1637 );
    xnor g3990 ( n9229 , n11171 , n5712 );
    and g3991 ( n9916 , n5794 , n4340 );
    and g3992 ( n5400 , n10057 , n5822 );
    or g3993 ( n11036 , n11958 , n11122 );
    not g3994 ( n12129 , n3467 );
    or g3995 ( n4313 , n7301 , n10158 );
    or g3996 ( n3110 , n9616 , n5262 );
    or g3997 ( n1156 , n2973 , n9613 );
    xnor g3998 ( n6201 , n12180 , n4558 );
    not g3999 ( n3819 , n10414 );
    or g4000 ( n1910 , n5404 , n6823 );
    or g4001 ( n6672 , n11801 , n10413 );
    or g4002 ( n5836 , n4628 , n2964 );
    and g4003 ( n11553 , n10899 , n7532 );
    or g4004 ( n11591 , n11887 , n4913 );
    and g4005 ( n10923 , n6481 , n7437 );
    and g4006 ( n7231 , n2012 , n11497 );
    xnor g4007 ( n11972 , n3067 , n1793 );
    and g4008 ( n11042 , n6945 , n423 );
    xnor g4009 ( n6220 , n6585 , n12534 );
    not g4010 ( n11573 , n3027 );
    xnor g4011 ( n2330 , n10498 , n7857 );
    or g4012 ( n11328 , n5780 , n960 );
    or g4013 ( n6108 , n1621 , n1331 );
    or g4014 ( n8977 , n9784 , n6920 );
    and g4015 ( n7477 , n4567 , n9960 );
    or g4016 ( n12622 , n6577 , n11820 );
    nor g4017 ( n5070 , n3716 , n3586 );
    and g4018 ( n6908 , n7167 , n2477 );
    xnor g4019 ( n4605 , n12231 , n5041 );
    not g4020 ( n7431 , n12166 );
    xnor g4021 ( n6097 , n7073 , n9628 );
    not g4022 ( n4945 , n4851 );
    xnor g4023 ( n5115 , n6497 , n10554 );
    xnor g4024 ( n4927 , n5368 , n11651 );
    xnor g4025 ( n11906 , n4388 , n4898 );
    and g4026 ( n7679 , n7643 , n913 );
    and g4027 ( n7840 , n1854 , n4620 );
    xnor g4028 ( n11400 , n3089 , n3692 );
    not g4029 ( n6314 , n9444 );
    xnor g4030 ( n6063 , n8902 , n12784 );
    and g4031 ( n1408 , n9394 , n6789 );
    or g4032 ( n10117 , n12833 , n984 );
    or g4033 ( n6810 , n4724 , n7896 );
    or g4034 ( n8393 , n11923 , n8285 );
    and g4035 ( n11964 , n10740 , n5703 );
    or g4036 ( n10849 , n3930 , n4483 );
    and g4037 ( n11099 , n1911 , n1004 );
    not g4038 ( n3197 , n9131 );
    xnor g4039 ( n7543 , n7127 , n7774 );
    nor g4040 ( n786 , n95 , n6792 );
    or g4041 ( n392 , n9170 , n7424 );
    or g4042 ( n12874 , n9005 , n1608 );
    and g4043 ( n3709 , n969 , n5046 );
    or g4044 ( n4866 , n9373 , n4527 );
    and g4045 ( n10692 , n5860 , n5760 );
    xnor g4046 ( n11951 , n7502 , n12213 );
    or g4047 ( n1368 , n566 , n5656 );
    or g4048 ( n6669 , n5355 , n4775 );
    xnor g4049 ( n4362 , n2458 , n12238 );
    or g4050 ( n9009 , n9343 , n12425 );
    or g4051 ( n2101 , n2448 , n3799 );
    not g4052 ( n10068 , n11653 );
    and g4053 ( n6504 , n3625 , n9031 );
    or g4054 ( n11128 , n11433 , n5540 );
    xnor g4055 ( n7 , n3476 , n1193 );
    and g4056 ( n12087 , n12069 , n2558 );
    xnor g4057 ( n12240 , n12318 , n6900 );
    xnor g4058 ( n1596 , n10374 , n3898 );
    xor g4059 ( n5899 , n2913 , n368 );
    and g4060 ( n11336 , n7043 , n7190 );
    and g4061 ( n3162 , n10983 , n2817 );
    and g4062 ( n3309 , n11036 , n8030 );
    nor g4063 ( n1140 , n11692 , n12484 );
    xnor g4064 ( n8693 , n9348 , n7667 );
    or g4065 ( n1946 , n10196 , n4642 );
    or g4066 ( n8766 , n9389 , n1738 );
    and g4067 ( n4718 , n1041 , n11364 );
    xnor g4068 ( n4569 , n7726 , n5533 );
    or g4069 ( n7626 , n7874 , n12918 );
    not g4070 ( n8890 , n3163 );
    xnor g4071 ( n5162 , n10960 , n10315 );
    and g4072 ( n1619 , n8743 , n9505 );
    or g4073 ( n4018 , n9884 , n3411 );
    and g4074 ( n682 , n8785 , n6021 );
    not g4075 ( n10123 , n6001 );
    and g4076 ( n3106 , n11070 , n4599 );
    or g4077 ( n5027 , n8412 , n3521 );
    or g4078 ( n10874 , n5530 , n1163 );
    xnor g4079 ( n11702 , n3397 , n6382 );
    or g4080 ( n5341 , n994 , n1546 );
    not g4081 ( n2740 , n9298 );
    and g4082 ( n1722 , n11900 , n8871 );
    xnor g4083 ( n2426 , n7376 , n7465 );
    or g4084 ( n7306 , n8428 , n11896 );
    xnor g4085 ( n9515 , n7585 , n8283 );
    or g4086 ( n9401 , n2917 , n2465 );
    xnor g4087 ( n6008 , n6051 , n9635 );
    nor g4088 ( n12485 , n3712 , n9805 );
    xnor g4089 ( n6210 , n1884 , n3312 );
    not g4090 ( n12735 , n6254 );
    xnor g4091 ( n8075 , n6506 , n12372 );
    or g4092 ( n8737 , n11026 , n1047 );
    xnor g4093 ( n10949 , n948 , n7482 );
    and g4094 ( n6159 , n8418 , n11472 );
    and g4095 ( n10734 , n5215 , n8095 );
    and g4096 ( n11802 , n9970 , n2224 );
    or g4097 ( n6303 , n4604 , n5220 );
    and g4098 ( n6205 , n6995 , n2405 );
    not g4099 ( n3721 , n12757 );
    or g4100 ( n6013 , n8192 , n10193 );
    xnor g4101 ( n6807 , n10610 , n1855 );
    nor g4102 ( n4479 , n2109 , n6274 );
    not g4103 ( n4342 , n11491 );
    or g4104 ( n3265 , n12119 , n12735 );
    or g4105 ( n12549 , n4674 , n826 );
    not g4106 ( n12816 , n12709 );
    and g4107 ( n2298 , n5573 , n7618 );
    nor g4108 ( n2951 , n7732 , n11246 );
    not g4109 ( n2302 , n6015 );
    or g4110 ( n9705 , n10396 , n11491 );
    xnor g4111 ( n2789 , n9515 , n2825 );
    or g4112 ( n12920 , n7283 , n7389 );
    or g4113 ( n1990 , n3743 , n1476 );
    xor g4114 ( n9814 , n395 , n8479 );
    or g4115 ( n7322 , n2217 , n8285 );
    or g4116 ( n5917 , n1446 , n10492 );
    xnor g4117 ( n8077 , n574 , n6427 );
    not g4118 ( n6656 , n4273 );
    not g4119 ( n580 , n6242 );
    xnor g4120 ( n11054 , n8836 , n11376 );
    and g4121 ( n4502 , n2272 , n10258 );
    or g4122 ( n3284 , n8026 , n11122 );
    and g4123 ( n987 , n7617 , n9667 );
    or g4124 ( n2753 , n12644 , n265 );
    or g4125 ( n1247 , n6145 , n3647 );
    or g4126 ( n6195 , n7495 , n3911 );
    or g4127 ( n4613 , n10196 , n1047 );
    xnor g4128 ( n8614 , n11984 , n6460 );
    xnor g4129 ( n6949 , n10155 , n2140 );
    and g4130 ( n6855 , n3627 , n7265 );
    and g4131 ( n8241 , n7965 , n10848 );
    xnor g4132 ( n8490 , n478 , n12475 );
    or g4133 ( n1308 , n686 , n3903 );
    nor g4134 ( n7191 , n11343 , n3499 );
    xor g4135 ( n10851 , n11557 , n12360 );
    or g4136 ( n12195 , n3746 , n995 );
    nor g4137 ( n11683 , n9987 , n2361 );
    xnor g4138 ( n6664 , n8786 , n2419 );
    and g4139 ( n3741 , n5151 , n11670 );
    or g4140 ( n6172 , n4666 , n10863 );
    and g4141 ( n10522 , n6770 , n4370 );
    not g4142 ( n8438 , n12123 );
    or g4143 ( n9314 , n880 , n11758 );
    nor g4144 ( n6940 , n1448 , n5789 );
    xnor g4145 ( n9381 , n11148 , n12140 );
    or g4146 ( n7120 , n2017 , n2883 );
    or g4147 ( n8273 , n2456 , n12735 );
    and g4148 ( n3505 , n10091 , n100 );
    and g4149 ( n12870 , n1717 , n3813 );
    not g4150 ( n9878 , n6294 );
    not g4151 ( n1129 , n1689 );
    or g4152 ( n9859 , n636 , n2964 );
    or g4153 ( n7788 , n2584 , n9258 );
    nor g4154 ( n6047 , n6033 , n214 );
    not g4155 ( n2843 , n9465 );
    and g4156 ( n7224 , n7236 , n8028 );
    and g4157 ( n8 , n3156 , n12008 );
    xnor g4158 ( n2902 , n11187 , n7671 );
    or g4159 ( n1515 , n12007 , n2328 );
    or g4160 ( n9764 , n8552 , n8648 );
    or g4161 ( n2268 , n9389 , n3911 );
    or g4162 ( n10585 , n1051 , n7876 );
    not g4163 ( n4869 , n10399 );
    xnor g4164 ( n11620 , n7898 , n2622 );
    nor g4165 ( n4855 , n7911 , n5323 );
    not g4166 ( n12900 , n85 );
    or g4167 ( n5456 , n5575 , n6197 );
    xnor g4168 ( n3532 , n1409 , n12780 );
    or g4169 ( n2327 , n418 , n7924 );
    nor g4170 ( n2306 , n4781 , n138 );
    or g4171 ( n2970 , n6237 , n9526 );
    xnor g4172 ( n7092 , n11405 , n11665 );
    or g4173 ( n1865 , n12361 , n11896 );
    or g4174 ( n7888 , n5838 , n10892 );
    or g4175 ( n7645 , n1890 , n3343 );
    or g4176 ( n4591 , n5765 , n609 );
    xnor g4177 ( n5804 , n8191 , n11176 );
    not g4178 ( n166 , n12778 );
    xnor g4179 ( n8965 , n10467 , n12288 );
    and g4180 ( n11975 , n11668 , n7538 );
    or g4181 ( n12203 , n191 , n4775 );
    xnor g4182 ( n228 , n3075 , n314 );
    and g4183 ( n11648 , n11856 , n6911 );
    or g4184 ( n2521 , n3026 , n3896 );
    or g4185 ( n3976 , n5355 , n8524 );
    and g4186 ( n1002 , n6894 , n7105 );
    and g4187 ( n3516 , n7044 , n10185 );
    or g4188 ( n2008 , n12361 , n2232 );
    not g4189 ( n6416 , n10466 );
    and g4190 ( n12749 , n4994 , n2980 );
    or g4191 ( n6261 , n8214 , n10857 );
    or g4192 ( n5984 , n6718 , n7921 );
    nor g4193 ( n546 , n10019 , n11667 );
    or g4194 ( n5753 , n3153 , n6982 );
    xnor g4195 ( n4233 , n8378 , n8061 );
    and g4196 ( n5482 , n2067 , n12568 );
    xnor g4197 ( n1855 , n4856 , n3348 );
    not g4198 ( n6755 , n2903 );
    xnor g4199 ( n3960 , n8934 , n10460 );
    and g4200 ( n3410 , n444 , n12829 );
    and g4201 ( n9506 , n3620 , n5718 );
    or g4202 ( n3449 , n3820 , n5258 );
    and g4203 ( n2121 , n11080 , n12597 );
    xnor g4204 ( n9316 , n10059 , n10827 );
    and g4205 ( n10265 , n2226 , n8819 );
    xnor g4206 ( n7385 , n12827 , n1674 );
    xnor g4207 ( n14 , n4994 , n2980 );
    and g4208 ( n1436 , n4644 , n11624 );
    not g4209 ( n12371 , n1322 );
    not g4210 ( n6863 , n3354 );
    or g4211 ( n3905 , n10347 , n12182 );
    or g4212 ( n6391 , n5016 , n12202 );
    or g4213 ( n5441 , n2456 , n3924 );
    not g4214 ( n9625 , n8370 );
    xnor g4215 ( n11530 , n11286 , n12320 );
    and g4216 ( n3388 , n5404 , n6823 );
    or g4217 ( n9588 , n3050 , n11524 );
    xnor g4218 ( n4821 , n7247 , n199 );
    nor g4219 ( n9207 , n1350 , n1912 );
    or g4220 ( n1071 , n7536 , n1191 );
    nor g4221 ( n1754 , n646 , n494 );
    xnor g4222 ( n858 , n1746 , n2404 );
    nor g4223 ( n10320 , n11490 , n1919 );
    nor g4224 ( n3233 , n5969 , n1313 );
    or g4225 ( n10139 , n2217 , n4642 );
    xnor g4226 ( n11391 , n6801 , n6011 );
    not g4227 ( n177 , n9289 );
    or g4228 ( n133 , n10108 , n5497 );
    xnor g4229 ( n11763 , n10587 , n12727 );
    or g4230 ( n7298 , n602 , n10024 );
    xnor g4231 ( n6333 , n8445 , n9766 );
    xnor g4232 ( n871 , n11712 , n9574 );
    xnor g4233 ( n6129 , n3335 , n9062 );
    or g4234 ( n8645 , n2244 , n9402 );
    and g4235 ( n62 , n12324 , n2736 );
    xnor g4236 ( n3143 , n12653 , n5229 );
    or g4237 ( n11244 , n2033 , n8014 );
    or g4238 ( n4432 , n989 , n4400 );
    or g4239 ( n10838 , n10157 , n8830 );
    xnor g4240 ( n644 , n8116 , n9576 );
    and g4241 ( n7002 , n2652 , n3518 );
    xnor g4242 ( n12084 , n2899 , n4182 );
    nor g4243 ( n2098 , n1907 , n12566 );
    xnor g4244 ( n5576 , n5584 , n5672 );
    or g4245 ( n4173 , n2874 , n9587 );
    or g4246 ( n8575 , n12698 , n2298 );
    xnor g4247 ( n446 , n9363 , n4807 );
    xnor g4248 ( n11012 , n10810 , n4144 );
    or g4249 ( n7532 , n884 , n3639 );
    not g4250 ( n11891 , n6439 );
    or g4251 ( n9895 , n3344 , n11086 );
    or g4252 ( n3382 , n10343 , n9535 );
    or g4253 ( n10940 , n9170 , n2358 );
    nor g4254 ( n5367 , n5720 , n6565 );
    and g4255 ( n10501 , n9908 , n12874 );
    or g4256 ( n1947 , n7417 , n2149 );
    not g4257 ( n4452 , n623 );
    not g4258 ( n9373 , n6358 );
    xnor g4259 ( n2759 , n1154 , n10804 );
    or g4260 ( n10997 , n8187 , n12328 );
    and g4261 ( n9665 , n432 , n9549 );
    or g4262 ( n12739 , n3096 , n3903 );
    xnor g4263 ( n6753 , n8580 , n6223 );
    xnor g4264 ( n9293 , n6938 , n5481 );
    xnor g4265 ( n8950 , n880 , n5131 );
    or g4266 ( n5528 , n12953 , n4878 );
    or g4267 ( n1483 , n11719 , n3911 );
    not g4268 ( n12102 , n5901 );
    or g4269 ( n11161 , n6320 , n2821 );
    or g4270 ( n1727 , n2539 , n5910 );
    or g4271 ( n6184 , n9101 , n9516 );
    xnor g4272 ( n11853 , n12200 , n12789 );
    and g4273 ( n10132 , n515 , n5941 );
    xnor g4274 ( n6217 , n4791 , n5925 );
    xnor g4275 ( n1269 , n10631 , n2095 );
    and g4276 ( n55 , n4984 , n9153 );
    xnor g4277 ( n2070 , n646 , n11540 );
    or g4278 ( n6782 , n4498 , n7424 );
    xnor g4279 ( n9819 , n10648 , n8179 );
    xnor g4280 ( n2611 , n1680 , n31 );
    and g4281 ( n335 , n4948 , n12021 );
    or g4282 ( n8462 , n3262 , n4072 );
    nor g4283 ( n11916 , n2713 , n6937 );
    or g4284 ( n5136 , n3617 , n8740 );
    xnor g4285 ( n7268 , n9460 , n6159 );
    and g4286 ( n12690 , n9274 , n10814 );
    nor g4287 ( n4352 , n10279 , n9855 );
    not g4288 ( n11977 , n8051 );
    xnor g4289 ( n10313 , n7650 , n3 );
    not g4290 ( n524 , n2481 );
    or g4291 ( n3107 , n1898 , n3673 );
    or g4292 ( n9807 , n11838 , n7344 );
    or g4293 ( n11722 , n2976 , n11495 );
    xnor g4294 ( n4248 , n10255 , n696 );
    and g4295 ( n8700 , n1598 , n5564 );
    xnor g4296 ( n1885 , n11535 , n8403 );
    and g4297 ( n1048 , n3933 , n3406 );
    or g4298 ( n3648 , n9176 , n12409 );
    not g4299 ( n4285 , n4414 );
    or g4300 ( n11368 , n7709 , n9160 );
    xnor g4301 ( n4349 , n2321 , n5704 );
    or g4302 ( n6473 , n3820 , n9521 );
    nor g4303 ( n6752 , n2319 , n10252 );
    not g4304 ( n2574 , n2761 );
    xnor g4305 ( n199 , n11517 , n5883 );
    or g4306 ( n5749 , n4274 , n11810 );
    xnor g4307 ( n6107 , n3533 , n1284 );
    and g4308 ( n11681 , n4957 , n7771 );
    xnor g4309 ( n10084 , n4747 , n2534 );
    or g4310 ( n4544 , n11026 , n28 );
    and g4311 ( n591 , n11142 , n10187 );
    and g4312 ( n2894 , n10738 , n3150 );
    xnor g4313 ( n12718 , n9853 , n1831 );
    or g4314 ( n2493 , n4657 , n3971 );
    not g4315 ( n4884 , n7224 );
    nor g4316 ( n3427 , n1007 , n10410 );
    not g4317 ( n4350 , n1485 );
    xnor g4318 ( n6841 , n9518 , n5197 );
    not g4319 ( n8326 , n9591 );
    xnor g4320 ( n8565 , n3915 , n11558 );
    and g4321 ( n10237 , n7906 , n9794 );
    xnor g4322 ( n8911 , n457 , n8086 );
    or g4323 ( n6074 , n9170 , n4400 );
    or g4324 ( n5739 , n191 , n2358 );
    and g4325 ( n585 , n6877 , n3602 );
    xnor g4326 ( n7157 , n2352 , n2643 );
    xnor g4327 ( n10970 , n1433 , n5853 );
    or g4328 ( n4716 , n2099 , n8648 );
    or g4329 ( n6498 , n12503 , n4527 );
    nor g4330 ( n12260 , n8608 , n8160 );
    or g4331 ( n11542 , n11641 , n12379 );
    or g4332 ( n6793 , n306 , n40 );
    or g4333 ( n10252 , n11923 , n5502 );
    or g4334 ( n3165 , n4352 , n1388 );
    or g4335 ( n4001 , n989 , n7703 );
    not g4336 ( n1691 , n972 );
    or g4337 ( n2792 , n5235 , n433 );
    or g4338 ( n12155 , n6718 , n4875 );
    or g4339 ( n12289 , n2099 , n6071 );
    nor g4340 ( n4311 , n4224 , n7290 );
    and g4341 ( n7941 , n11324 , n12756 );
    or g4342 ( n9379 , n191 , n510 );
    xnor g4343 ( n2333 , n8499 , n7574 );
    xnor g4344 ( n2095 , n3184 , n11333 );
    or g4345 ( n7707 , n4183 , n3886 );
    xnor g4346 ( n12885 , n6174 , n1885 );
    or g4347 ( n6066 , n3743 , n1047 );
    xnor g4348 ( n11703 , n11713 , n4695 );
    and g4349 ( n3945 , n10845 , n8426 );
    not g4350 ( n4825 , n12398 );
    not g4351 ( n9659 , n10160 );
    xnor g4352 ( n5447 , n11835 , n2891 );
    xnor g4353 ( n8666 , n8439 , n8953 );
    not g4354 ( n8845 , n12455 );
    xnor g4355 ( n10978 , n5739 , n10241 );
    xnor g4356 ( n4409 , n7509 , n9998 );
    or g4357 ( n8180 , n7709 , n2020 );
    not g4358 ( n2217 , n11222 );
    not g4359 ( n10279 , n2569 );
    xnor g4360 ( n5047 , n10434 , n1362 );
    nor g4361 ( n8188 , n8290 , n5095 );
    or g4362 ( n12332 , n2456 , n8259 );
    and g4363 ( n10295 , n5209 , n10312 );
    nor g4364 ( n8635 , n6393 , n1343 );
    not g4365 ( n3950 , n6369 );
    or g4366 ( n9970 , n8002 , n8934 );
    xnor g4367 ( n9660 , n4726 , n8098 );
    and g4368 ( n2257 , n2097 , n3792 );
    and g4369 ( n5665 , n9400 , n7354 );
    or g4370 ( n12721 , n320 , n8869 );
    not g4371 ( n11433 , n10678 );
    nor g4372 ( n5420 , n9980 , n1587 );
    not g4373 ( n5355 , n5305 );
    xnor g4374 ( n7711 , n9701 , n6861 );
    xnor g4375 ( n2828 , n12336 , n3572 );
    not g4376 ( n12662 , n3513 );
    nor g4377 ( n9762 , n2590 , n1544 );
    or g4378 ( n5204 , n7449 , n1047 );
    or g4379 ( n7869 , n5765 , n7506 );
    or g4380 ( n4413 , n7391 , n510 );
    or g4381 ( n4078 , n597 , n5896 );
    or g4382 ( n6827 , n3383 , n2297 );
    not g4383 ( n3746 , n6776 );
    and g4384 ( n6723 , n11893 , n9885 );
    xnor g4385 ( n11772 , n8374 , n3113 );
    xnor g4386 ( n11268 , n2100 , n4650 );
    xnor g4387 ( n10866 , n8847 , n9356 );
    xnor g4388 ( n5500 , n12856 , n7698 );
    not g4389 ( n1437 , n10753 );
    and g4390 ( n10355 , n4535 , n501 );
    xnor g4391 ( n9310 , n1435 , n9040 );
    xnor g4392 ( n5734 , n8954 , n6852 );
    xnor g4393 ( n9026 , n5405 , n8025 );
    not g4394 ( n9934 , n5849 );
    and g4395 ( n2017 , n10614 , n7859 );
    xnor g4396 ( n3809 , n3968 , n11016 );
    nor g4397 ( n4695 , n11419 , n12685 );
    or g4398 ( n246 , n3240 , n8801 );
    or g4399 ( n11593 , n3127 , n10066 );
    xnor g4400 ( n8047 , n2308 , n10415 );
    or g4401 ( n3418 , n12119 , n4249 );
    nor g4402 ( n4027 , n8102 , n5006 );
    and g4403 ( n11366 , n1791 , n5344 );
    not g4404 ( n11422 , n4651 );
    nor g4405 ( n2291 , n11540 , n1736 );
    or g4406 ( n7331 , n3746 , n5538 );
    or g4407 ( n2213 , n10835 , n5258 );
    nor g4408 ( n10349 , n5567 , n7187 );
    or g4409 ( n4510 , n5765 , n5258 );
    xnor g4410 ( n4795 , n9982 , n10923 );
    not g4411 ( n11144 , n9676 );
    and g4412 ( n8851 , n5331 , n5645 );
    not g4413 ( n7810 , n8672 );
    or g4414 ( n10423 , n3838 , n5529 );
    xnor g4415 ( n8249 , n6331 , n1383 );
    and g4416 ( n10850 , n804 , n3714 );
    or g4417 ( n11179 , n9170 , n10066 );
    or g4418 ( n4390 , n7283 , n12328 );
    and g4419 ( n11575 , n1114 , n12030 );
    xnor g4420 ( n2404 , n5475 , n1395 );
    not g4421 ( n6811 , n3821 );
    not g4422 ( n12294 , n12248 );
    nor g4423 ( n4820 , n810 , n2058 );
    not g4424 ( n4719 , n2150 );
    or g4425 ( n4152 , n6910 , n2668 );
    not g4426 ( n7274 , n3601 );
    or g4427 ( n4038 , n12340 , n1385 );
    or g4428 ( n1061 , n1699 , n9586 );
    xnor g4429 ( n3893 , n4119 , n6949 );
    not g4430 ( n2367 , n45 );
    or g4431 ( n6481 , n5730 , n10407 );
    and g4432 ( n10715 , n1402 , n5866 );
    and g4433 ( n7123 , n6784 , n2103 );
    or g4434 ( n127 , n5832 , n6531 );
    xnor g4435 ( n2077 , n5269 , n1535 );
    xnor g4436 ( n2138 , n1694 , n3727 );
    not g4437 ( n11159 , n7954 );
    xnor g4438 ( n4003 , n8799 , n4811 );
    not g4439 ( n8703 , n3588 );
    and g4440 ( n9466 , n7732 , n11246 );
    not g4441 ( n4653 , n6342 );
    or g4442 ( n3395 , n10196 , n5258 );
    xnor g4443 ( n759 , n4036 , n9503 );
    xnor g4444 ( n10044 , n9610 , n8172 );
    or g4445 ( n1560 , n11552 , n795 );
    and g4446 ( n12817 , n3747 , n12249 );
    and g4447 ( n2680 , n12705 , n2879 );
    not g4448 ( n608 , n7039 );
    or g4449 ( n5601 , n11923 , n9160 );
    or g4450 ( n1565 , n4750 , n4652 );
    not g4451 ( n6726 , n8130 );
    and g4452 ( n1577 , n949 , n5917 );
    or g4453 ( n2899 , n5355 , n130 );
    or g4454 ( n5990 , n910 , n9852 );
    xnor g4455 ( n12475 , n4460 , n5272 );
    or g4456 ( n4232 , n2099 , n8957 );
    xnor g4457 ( n70 , n3758 , n7031 );
    or g4458 ( n168 , n11305 , n10501 );
    or g4459 ( n1377 , n6451 , n2894 );
    not g4460 ( n8265 , n1922 );
    or g4461 ( n1254 , n8094 , n12865 );
    or g4462 ( n5395 , n4469 , n1428 );
    not g4463 ( n2506 , n6092 );
    or g4464 ( n6268 , n2099 , n5781 );
    or g4465 ( n7021 , n8552 , n530 );
    xnor g4466 ( n3184 , n5221 , n8032 );
    not g4467 ( n4735 , n8049 );
    xnor g4468 ( n1823 , n7942 , n2484 );
    not g4469 ( n12340 , n6813 );
    or g4470 ( n12043 , n11093 , n9211 );
    not g4471 ( n10600 , n3705 );
    xnor g4472 ( n6266 , n6779 , n4801 );
    or g4473 ( n1601 , n5397 , n9174 );
    not g4474 ( n9582 , n3350 );
    nor g4475 ( n4671 , n3579 , n4342 );
    and g4476 ( n12542 , n2660 , n10205 );
    not g4477 ( n8367 , n1201 );
    xnor g4478 ( n86 , n10964 , n1311 );
    not g4479 ( n7785 , n3968 );
    nor g4480 ( n6965 , n12502 , n11276 );
    or g4481 ( n519 , n1539 , n11827 );
    and g4482 ( n2133 , n2400 , n2705 );
    and g4483 ( n3512 , n4997 , n3937 );
    or g4484 ( n7348 , n752 , n12274 );
    nor g4485 ( n1196 , n2858 , n10188 );
    xnor g4486 ( n6792 , n2373 , n3696 );
    and g4487 ( n9360 , n9826 , n3979 );
    not g4488 ( n6076 , n42 );
    or g4489 ( n9394 , n7037 , n3232 );
    or g4490 ( n12157 , n7391 , n1162 );
    not g4491 ( n9458 , n11086 );
    not g4492 ( n3979 , n6771 );
    and g4493 ( n5519 , n8197 , n1098 );
    or g4494 ( n2979 , n9170 , n1079 );
    not g4495 ( n8685 , n2632 );
    and g4496 ( n9165 , n1277 , n4946 );
    and g4497 ( n10152 , n9377 , n6523 );
    not g4498 ( n5897 , n10558 );
    nor g4499 ( n3925 , n8447 , n203 );
    xnor g4500 ( n9200 , n5231 , n7537 );
    xnor g4501 ( n10387 , n12064 , n11987 );
    xnor g4502 ( n1545 , n5859 , n12038 );
    and g4503 ( n6317 , n3257 , n4096 );
    not g4504 ( n6887 , n3894 );
    or g4505 ( n8313 , n10835 , n8643 );
    not g4506 ( n2256 , n2007 );
    not g4507 ( n995 , n9189 );
    xnor g4508 ( n3360 , n8260 , n12065 );
    xnor g4509 ( n245 , n8362 , n12232 );
    and g4510 ( n1359 , n2524 , n11431 );
    xnor g4511 ( n3189 , n538 , n8465 );
    or g4512 ( n11253 , n11509 , n6804 );
    nor g4513 ( n4890 , n2176 , n8516 );
    not g4514 ( n12601 , n2336 );
    xnor g4515 ( n11774 , n7912 , n4136 );
    xnor g4516 ( n4620 , n6479 , n877 );
    xnor g4517 ( n12292 , n6370 , n5408 );
    xnor g4518 ( n10175 , n5746 , n7472 );
    nor g4519 ( n6183 , n7330 , n11630 );
    xnor g4520 ( n8998 , n4823 , n7140 );
    not g4521 ( n1633 , n10138 );
    xnor g4522 ( n823 , n9438 , n8744 );
    xnor g4523 ( n9135 , n1249 , n7963 );
    xnor g4524 ( n12667 , n4392 , n11710 );
    or g4525 ( n5242 , n5809 , n3224 );
    xnor g4526 ( n1080 , n4732 , n8773 );
    or g4527 ( n4297 , n8567 , n10536 );
    not g4528 ( n5127 , n847 );
    or g4529 ( n9974 , n8187 , n8524 );
    and g4530 ( n5614 , n12648 , n521 );
    or g4531 ( n320 , n6577 , n7952 );
    and g4532 ( n12168 , n3271 , n6179 );
    or g4533 ( n7324 , n7116 , n3421 );
    and g4534 ( n7233 , n2226 , n8595 );
    or g4535 ( n9600 , n10180 , n4234 );
    or g4536 ( n6719 , n2605 , n11921 );
    xnor g4537 ( n730 , n2032 , n1939 );
    not g4538 ( n1387 , n3491 );
    nor g4539 ( n2435 , n888 , n8328 );
    and g4540 ( n4168 , n6687 , n7265 );
    or g4541 ( n7801 , n3746 , n2232 );
    not g4542 ( n12930 , n84 );
    and g4543 ( n9662 , n9645 , n12301 );
    xnor g4544 ( n75 , n5100 , n6264 );
    and g4545 ( n3531 , n3870 , n7120 );
    or g4546 ( n7288 , n5494 , n5401 );
    not g4547 ( n11341 , n6222 );
    or g4548 ( n9648 , n12361 , n3903 );
    xnor g4549 ( n7957 , n4968 , n6992 );
    and g4550 ( n5746 , n9306 , n4078 );
    or g4551 ( n8551 , n11466 , n8222 );
    xnor g4552 ( n1540 , n12823 , n1143 );
    xnor g4553 ( n1849 , n6759 , n11160 );
    not g4554 ( n10767 , n11325 );
    and g4555 ( n5611 , n11723 , n12821 );
    and g4556 ( n3412 , n3020 , n1355 );
    or g4557 ( n10114 , n4589 , n9128 );
    not g4558 ( n140 , n7452 );
    not g4559 ( n6839 , n1702 );
    or g4560 ( n11080 , n752 , n12899 );
    xnor g4561 ( n6865 , n9915 , n1496 );
    not g4562 ( n8496 , n12788 );
    nor g4563 ( n8762 , n6686 , n5407 );
    or g4564 ( n5817 , n12248 , n7723 );
    xnor g4565 ( n2373 , n6308 , n5352 );
    not g4566 ( n264 , n11997 );
    or g4567 ( n12423 , n12119 , n1932 );
    or g4568 ( n10205 , n6095 , n781 );
    and g4569 ( n5164 , n3658 , n10207 );
    and g4570 ( n12110 , n12397 , n11508 );
    or g4571 ( n2862 , n8552 , n4913 );
    xnor g4572 ( n5472 , n8406 , n3783 );
    xnor g4573 ( n10238 , n11312 , n8586 );
    or g4574 ( n9158 , n2516 , n11559 );
    xor g4575 ( n4226 , n6527 , n10214 );
    and g4576 ( n12606 , n3279 , n6871 );
    xnor g4577 ( n4836 , n12552 , n8115 );
    not g4578 ( n7894 , n10152 );
    or g4579 ( n782 , n11476 , n1125 );
    nor g4580 ( n8498 , n7861 , n5327 );
    xnor g4581 ( n1953 , n12224 , n5268 );
    xnor g4582 ( n4165 , n8081 , n11340 );
    not g4583 ( n4628 , n8476 );
    or g4584 ( n11236 , n1937 , n5012 );
    or g4585 ( n9323 , n4784 , n3419 );
    or g4586 ( n3273 , n10108 , n1162 );
    xnor g4587 ( n11198 , n7627 , n12128 );
    or g4588 ( n10696 , n9389 , n561 );
    or g4589 ( n1181 , n8127 , n5497 );
    xnor g4590 ( n781 , n10567 , n2771 );
    xnor g4591 ( n911 , n11756 , n10459 );
    or g4592 ( n3021 , n9373 , n2020 );
    or g4593 ( n890 , n1811 , n829 );
    not g4594 ( n11347 , n7440 );
    or g4595 ( n6763 , n7901 , n5701 );
    xnor g4596 ( n7430 , n9146 , n2453 );
    xnor g4597 ( n10592 , n9565 , n6469 );
    xnor g4598 ( n6639 , n251 , n8980 );
    xnor g4599 ( n11828 , n9310 , n10043 );
    xnor g4600 ( n11819 , n6442 , n3462 );
    nor g4601 ( n3999 , n10887 , n323 );
    and g4602 ( n5061 , n5780 , n960 );
    and g4603 ( n8743 , n8759 , n2024 );
    and g4604 ( n5344 , n2813 , n7613 );
    not g4605 ( n2259 , n5694 );
    or g4606 ( n4511 , n9367 , n7471 );
    not g4607 ( n1729 , n11508 );
    xnor g4608 ( n457 , n10656 , n12903 );
    or g4609 ( n6245 , n8207 , n8650 );
    and g4610 ( n8925 , n3845 , n10733 );
    xnor g4611 ( n5830 , n8468 , n8278 );
    or g4612 ( n9616 , n10750 , n5326 );
    or g4613 ( n3848 , n5219 , n4926 );
    or g4614 ( n11595 , n8026 , n9971 );
    or g4615 ( n2686 , n2099 , n8644 );
    xnor g4616 ( n1964 , n5404 , n6823 );
    and g4617 ( n5646 , n5594 , n11095 );
    and g4618 ( n8199 , n7457 , n872 );
    nor g4619 ( n7606 , n463 , n625 );
    or g4620 ( n12468 , n488 , n10691 );
    or g4621 ( n8852 , n6718 , n8285 );
    not g4622 ( n2971 , n8656 );
    not g4623 ( n7147 , n8266 );
    xnor g4624 ( n8324 , n2467 , n311 );
    or g4625 ( n10656 , n12853 , n826 );
    xnor g4626 ( n247 , n4429 , n4659 );
    not g4627 ( n6412 , n3472 );
    or g4628 ( n11894 , n9837 , n6529 );
    and g4629 ( n10515 , n5681 , n10646 );
    and g4630 ( n7134 , n9688 , n8446 );
    or g4631 ( n7101 , n6577 , n11775 );
    or g4632 ( n2704 , n3743 , n3451 );
    or g4633 ( n11017 , n8127 , n10066 );
    not g4634 ( n7839 , n10510 );
    xnor g4635 ( n10615 , n8009 , n4744 );
    or g4636 ( n10179 , n12800 , n9418 );
    nor g4637 ( n12185 , n9391 , n5302 );
    and g4638 ( n680 , n1557 , n7030 );
    xnor g4639 ( n11089 , n5780 , n960 );
    or g4640 ( n1321 , n1051 , n6197 );
    and g4641 ( n6068 , n11822 , n8382 );
    or g4642 ( n7745 , n10745 , n12072 );
    or g4643 ( n11751 , n8959 , n8768 );
    or g4644 ( n2111 , n8959 , n7558 );
    or g4645 ( n8118 , n7391 , n7424 );
    xnor g4646 ( n2477 , n9360 , n4260 );
    and g4647 ( n1491 , n8550 , n10934 );
    or g4648 ( n6475 , n8187 , n12843 );
    or g4649 ( n4373 , n2217 , n609 );
    or g4650 ( n4789 , n8395 , n10588 );
    and g4651 ( n7950 , n11110 , n10794 );
    xnor g4652 ( n7812 , n7429 , n4344 );
    nor g4653 ( n6923 , n10128 , n6714 );
    and g4654 ( n7625 , n10636 , n367 );
    and g4655 ( n2157 , n7992 , n8569 );
    or g4656 ( n8310 , n8552 , n12080 );
    xnor g4657 ( n11053 , n3987 , n11636 );
    and g4658 ( n6896 , n10466 , n2678 );
    xnor g4659 ( n8283 , n12046 , n1287 );
    or g4660 ( n11829 , n8778 , n12718 );
    or g4661 ( n8550 , n2217 , n5759 );
    not g4662 ( n11287 , n9720 );
    or g4663 ( n11657 , n4205 , n10817 );
    not g4664 ( n8513 , n917 );
    and g4665 ( n12092 , n9661 , n5130 );
    and g4666 ( n4658 , n4788 , n9620 );
    not g4667 ( n12187 , n5622 );
    or g4668 ( n4035 , n10879 , n11746 );
    or g4669 ( n517 , n4179 , n8266 );
    or g4670 ( n548 , n9370 , n8524 );
    xnor g4671 ( n4030 , n7276 , n5974 );
    xnor g4672 ( n9319 , n285 , n180 );
    and g4673 ( n5755 , n1070 , n4306 );
    nor g4674 ( n5868 , n3433 , n1722 );
    or g4675 ( n10078 , n3836 , n12371 );
    xnor g4676 ( n9129 , n5384 , n12652 );
    and g4677 ( n11043 , n1382 , n11657 );
    and g4678 ( n4145 , n10545 , n1512 );
    or g4679 ( n6414 , n12361 , n2815 );
    and g4680 ( n6395 , n10212 , n907 );
    nor g4681 ( n4704 , n1760 , n2859 );
    nor g4682 ( n6336 , n12579 , n6506 );
    and g4683 ( n4747 , n10224 , n11452 );
    nor g4684 ( n11004 , n805 , n7656 );
    xnor g4685 ( n3579 , n3753 , n2941 );
    xnor g4686 ( n6156 , n12870 , n440 );
    nor g4687 ( n9861 , n2947 , n940 );
    xnor g4688 ( n5269 , n10608 , n5950 );
    or g4689 ( n9481 , n4628 , n12446 );
    not g4690 ( n5088 , n11533 );
    or g4691 ( n12052 , n8187 , n1915 );
    xnor g4692 ( n11665 , n10148 , n7996 );
    xnor g4693 ( n5731 , n9626 , n1597 );
    xnor g4694 ( n3459 , n867 , n4731 );
    or g4695 ( n334 , n9878 , n3224 );
    xnor g4696 ( n7692 , n7151 , n1501 );
    and g4697 ( n6039 , n12673 , n10440 );
    or g4698 ( n5125 , n9688 , n8446 );
    not g4699 ( n5439 , n3130 );
    xnor g4700 ( n9686 , n12123 , n9490 );
    not g4701 ( n1741 , n7920 );
    and g4702 ( n11274 , n10124 , n455 );
    xnor g4703 ( n9113 , n4420 , n1603 );
    or g4704 ( n492 , n9370 , n4242 );
    and g4705 ( n3920 , n2845 , n4177 );
    xnor g4706 ( n5556 , n10667 , n8317 );
    or g4707 ( n8251 , n8187 , n6389 );
    or g4708 ( n89 , n3363 , n5509 );
    xnor g4709 ( n7814 , n4524 , n10068 );
    and g4710 ( n6734 , n8193 , n5002 );
    or g4711 ( n9876 , n4894 , n36 );
    xnor g4712 ( n1608 , n9787 , n1904 );
    xnor g4713 ( n10539 , n1705 , n12251 );
    not g4714 ( n8577 , n9550 );
    xnor g4715 ( n5259 , n1112 , n8588 );
    or g4716 ( n10057 , n8870 , n8655 );
    xnor g4717 ( n2897 , n7505 , n3049 );
    xnor g4718 ( n3128 , n9339 , n4763 );
    nor g4719 ( n10184 , n11232 , n8064 );
    xnor g4720 ( n10041 , n349 , n3520 );
    nor g4721 ( n6812 , n8522 , n3882 );
    or g4722 ( n6370 , n12119 , n12535 );
    xnor g4723 ( n9820 , n1264 , n4776 );
    or g4724 ( n4785 , n9379 , n1356 );
    xnor g4725 ( n851 , n12327 , n1660 );
    or g4726 ( n5231 , n8583 , n4875 );
    xnor g4727 ( n812 , n6175 , n11006 );
    not g4728 ( n1562 , n3928 );
    or g4729 ( n2285 , n752 , n9741 );
    or g4730 ( n11245 , n11026 , n3606 );
    xnor g4731 ( n11010 , n7243 , n2460 );
    xnor g4732 ( n7095 , n8904 , n12193 );
    or g4733 ( n9651 , n4911 , n5497 );
    and g4734 ( n11948 , n9029 , n2615 );
    or g4735 ( n6450 , n1016 , n1979 );
    xnor g4736 ( n3375 , n12532 , n1620 );
    not g4737 ( n11896 , n5105 );
    not g4738 ( n7657 , n1216 );
    not g4739 ( n9028 , n9655 );
    xnor g4740 ( n2073 , n4224 , n7155 );
    not g4741 ( n8830 , n7294 );
    xnor g4742 ( n689 , n1255 , n10444 );
    not g4743 ( n3948 , n3519 );
    not g4744 ( n12748 , n11050 );
    or g4745 ( n9732 , n3795 , n10294 );
    xnor g4746 ( n4810 , n1475 , n5414 );
    not g4747 ( n6124 , n1505 );
    xnor g4748 ( n1450 , n9089 , n11980 );
    xnor g4749 ( n7402 , n5832 , n6531 );
    and g4750 ( n10813 , n681 , n10418 );
    not g4751 ( n373 , n3921 );
    xnor g4752 ( n10115 , n1721 , n10114 );
    xnor g4753 ( n12649 , n7375 , n5256 );
    and g4754 ( n917 , n7588 , n9543 );
    not g4755 ( n6234 , n5299 );
    xnor g4756 ( n7075 , n3337 , n3294 );
    and g4757 ( n8042 , n3642 , n10963 );
    xnor g4758 ( n5336 , n5432 , n12292 );
    or g4759 ( n11126 , n8835 , n9595 );
    and g4760 ( n8958 , n7218 , n4313 );
    or g4761 ( n8839 , n11958 , n11410 );
    or g4762 ( n3207 , n6635 , n9863 );
    or g4763 ( n5393 , n11958 , n3468 );
    not g4764 ( n6747 , n11038 );
    nor g4765 ( n8972 , n9988 , n6332 );
    or g4766 ( n6105 , n11953 , n11242 );
    xnor g4767 ( n4741 , n3869 , n6209 );
    nor g4768 ( n11419 , n6374 , n5757 );
    or g4769 ( n6153 , n3096 , n7558 );
    or g4770 ( n11822 , n4480 , n7866 );
    nor g4771 ( n603 , n9499 , n17 );
    nor g4772 ( n1013 , n4142 , n4691 );
    or g4773 ( n10945 , n6718 , n3606 );
    and g4774 ( n2842 , n6786 , n10373 );
    or g4775 ( n12261 , n432 , n9549 );
    xnor g4776 ( n3787 , n2193 , n4708 );
    or g4777 ( n3393 , n5547 , n5810 );
    xnor g4778 ( n8520 , n3883 , n5807 );
    xnor g4779 ( n10769 , n1390 , n1292 );
    or g4780 ( n6021 , n6772 , n1596 );
    and g4781 ( n7701 , n5285 , n6902 );
    and g4782 ( n3991 , n7657 , n9315 );
    nor g4783 ( n2225 , n9164 , n6802 );
    xnor g4784 ( n5784 , n12799 , n12253 );
    and g4785 ( n1956 , n11627 , n7205 );
    nor g4786 ( n575 , n102 , n5875 );
    or g4787 ( n873 , n12090 , n4871 );
    and g4788 ( n12588 , n5319 , n9763 );
    and g4789 ( n12790 , n12115 , n1761 );
    or g4790 ( n11740 , n1419 , n9216 );
    and g4791 ( n214 , n2947 , n940 );
    xnor g4792 ( n841 , n5370 , n339 );
    or g4793 ( n5967 , n11026 , n8643 );
    nor g4794 ( n6657 , n3412 , n12407 );
    or g4795 ( n9212 , n12941 , n1624 );
    or g4796 ( n1663 , n10219 , n7477 );
    xnor g4797 ( n5475 , n11264 , n3744 );
    nor g4798 ( n11466 , n3198 , n12772 );
    or g4799 ( n6851 , n1900 , n9556 );
    and g4800 ( n12698 , n5247 , n9020 );
    and g4801 ( n7993 , n7236 , n9111 );
    xnor g4802 ( n9851 , n6313 , n498 );
    nor g4803 ( n3045 , n12950 , n1381 );
    or g4804 ( n2072 , n97 , n2129 );
    xnor g4805 ( n4975 , n4138 , n9929 );
    and g4806 ( n4724 , n9101 , n9516 );
    or g4807 ( n1654 , n11719 , n1455 );
    nor g4808 ( n2948 , n2075 , n6972 );
    xnor g4809 ( n100 , n11184 , n11018 );
    not g4810 ( n10449 , n6997 );
    xnor g4811 ( n5856 , n5324 , n518 );
    and g4812 ( n4108 , n2069 , n10458 );
    not g4813 ( n2766 , n5627 );
    or g4814 ( n10751 , n1200 , n1482 );
    and g4815 ( n9822 , n3700 , n5294 );
    and g4816 ( n10904 , n6867 , n187 );
    xnor g4817 ( n1694 , n11929 , n6253 );
    or g4818 ( n4966 , n11319 , n4310 );
    xnor g4819 ( n3492 , n5605 , n3745 );
    and g4820 ( n9765 , n8645 , n9594 );
    xnor g4821 ( n3404 , n6576 , n5150 );
    not g4822 ( n4177 , n6705 );
    or g4823 ( n1646 , n8959 , n11896 );
    not g4824 ( n12954 , n11708 );
    or g4825 ( n9090 , n5945 , n11775 );
    or g4826 ( n11060 , n7283 , n1546 );
    or g4827 ( n8916 , n10339 , n5468 );
    or g4828 ( n10136 , n7409 , n1868 );
    or g4829 ( n419 , n12038 , n1913 );
    xnor g4830 ( n5888 , n6070 , n56 );
    not g4831 ( n12771 , n9111 );
    xnor g4832 ( n11676 , n6190 , n11658 );
    xnor g4833 ( n6476 , n4647 , n11236 );
    and g4834 ( n3840 , n12750 , n376 );
    and g4835 ( n7440 , n5916 , n6785 );
    or g4836 ( n5885 , n114 , n6169 );
    and g4837 ( n12343 , n4189 , n4370 );
    xnor g4838 ( n8501 , n737 , n6132 );
    or g4839 ( n8445 , n1316 , n6898 );
    and g4840 ( n2805 , n12135 , n1380 );
    xnor g4841 ( n9366 , n1275 , n8240 );
    and g4842 ( n4437 , n8823 , n2049 );
    xnor g4843 ( n10913 , n10857 , n8385 );
    not g4844 ( n8073 , n6498 );
    xnor g4845 ( n278 , n458 , n2992 );
    xnor g4846 ( n8068 , n3340 , n4228 );
    or g4847 ( n10392 , n8839 , n10927 );
    nor g4848 ( n11283 , n5213 , n12602 );
    or g4849 ( n5512 , n807 , n2232 );
    nor g4850 ( n2315 , n1359 , n6658 );
    xnor g4851 ( n9197 , n3076 , n7402 );
    and g4852 ( n6080 , n2541 , n10427 );
    xnor g4853 ( n1457 , n663 , n9039 );
    nor g4854 ( n11899 , n8165 , n297 );
    not g4855 ( n3571 , n1426 );
    or g4856 ( n1484 , n2967 , n10447 );
    and g4857 ( n2408 , n8759 , n3602 );
    or g4858 ( n3406 , n9538 , n4064 );
    or g4859 ( n7209 , n1741 , n8715 );
    and g4860 ( n9049 , n12388 , n2492 );
    not g4861 ( n10634 , n5336 );
    or g4862 ( n11851 , n7283 , n2358 );
    xnor g4863 ( n11723 , n1518 , n3536 );
    or g4864 ( n8940 , n10247 , n5597 );
    and g4865 ( n9067 , n4255 , n10411 );
    or g4866 ( n5853 , n686 , n7952 );
    xnor g4867 ( n1195 , n1043 , n4780 );
    xnor g4868 ( n9469 , n8752 , n9850 );
    or g4869 ( n9029 , n4639 , n6140 );
    xnor g4870 ( n7697 , n10039 , n5591 );
    xnor g4871 ( n7991 , n12859 , n2652 );
    xnor g4872 ( n4607 , n8266 , n2102 );
    not g4873 ( n6042 , n5533 );
    or g4874 ( n3266 , n3573 , n10624 );
    or g4875 ( n2867 , n11059 , n12300 );
    and g4876 ( n6134 , n10626 , n12317 );
    and g4877 ( n2344 , n621 , n6844 );
    not g4878 ( n6362 , n1541 );
    xnor g4879 ( n10593 , n5603 , n11345 );
    and g4880 ( n10677 , n2534 , n4747 );
    or g4881 ( n8430 , n1465 , n6272 );
    or g4882 ( n7406 , n8136 , n4879 );
    nor g4883 ( n9449 , n3546 , n9225 );
    and g4884 ( n1634 , n5685 , n5658 );
    and g4885 ( n12466 , n11717 , n9120 );
    and g4886 ( n9657 , n7974 , n9532 );
    xor g4887 ( n11248 , n11460 , n39 );
    or g4888 ( n5923 , n5214 , n2616 );
    nor g4889 ( n3587 , n8334 , n6234 );
    or g4890 ( n9431 , n10799 , n917 );
    or g4891 ( n6296 , n10142 , n8735 );
    not g4892 ( n2668 , n8121 );
    or g4893 ( n11487 , n422 , n12482 );
    not g4894 ( n10716 , n146 );
    and g4895 ( n1454 , n1627 , n5813 );
    and g4896 ( n5656 , n2700 , n3268 );
    not g4897 ( n10709 , n9708 );
    and g4898 ( n5126 , n4451 , n1852 );
    nor g4899 ( n7059 , n1477 , n11049 );
    or g4900 ( n5605 , n5530 , n2964 );
    and g4901 ( n7729 , n11305 , n10501 );
    xnor g4902 ( n1031 , n11687 , n6599 );
    xnor g4903 ( n7738 , n12107 , n6632 );
    xnor g4904 ( n12651 , n9985 , n5777 );
    and g4905 ( n7908 , n2564 , n7265 );
    not g4906 ( n4425 , n2973 );
    and g4907 ( n8618 , n3887 , n3583 );
    or g4908 ( n5737 , n6226 , n7666 );
    not g4909 ( n47 , n2085 );
    or g4910 ( n6943 , n7015 , n9959 );
    xnor g4911 ( n12654 , n8510 , n8274 );
    or g4912 ( n9273 , n5341 , n11947 );
    not g4913 ( n1233 , n11280 );
    xnor g4914 ( n8403 , n7299 , n2239 );
    or g4915 ( n12253 , n5945 , n7952 );
    not g4916 ( n10332 , n6379 );
    and g4917 ( n5413 , n9233 , n8244 );
    xnor g4918 ( n12710 , n2014 , n12259 );
    and g4919 ( n2465 , n7376 , n7465 );
    or g4920 ( n12823 , n8738 , n9568 );
    or g4921 ( n5777 , n9507 , n1602 );
    xnor g4922 ( n8861 , n431 , n8546 );
    xnor g4923 ( n11237 , n531 , n1338 );
    and g4924 ( n5895 , n9400 , n12145 );
    not g4925 ( n711 , n12776 );
    xnor g4926 ( n5572 , n4458 , n9783 );
    and g4927 ( n74 , n6465 , n4645 );
    and g4928 ( n4281 , n2699 , n1618 );
    xnor g4929 ( n7635 , n11932 , n8841 );
    or g4930 ( n7851 , n7839 , n2232 );
    and g4931 ( n5399 , n3878 , n1565 );
    nor g4932 ( n5591 , n10291 , n11261 );
    xnor g4933 ( n5122 , n10699 , n5490 );
    or g4934 ( n2726 , n11026 , n9521 );
    or g4935 ( n5848 , n12237 , n12080 );
    nor g4936 ( n8527 , n8149 , n5517 );
    xnor g4937 ( n3483 , n121 , n1389 );
    or g4938 ( n668 , n6339 , n3157 );
    or g4939 ( n1679 , n5673 , n8756 );
    xnor g4940 ( n4240 , n9322 , n3475 );
    and g4941 ( n11796 , n11153 , n159 );
    or g4942 ( n5761 , n3127 , n4400 );
    or g4943 ( n3653 , n8583 , n795 );
    and g4944 ( n2860 , n5340 , n11957 );
    and g4945 ( n756 , n8273 , n4909 );
    not g4946 ( n9237 , n4105 );
    not g4947 ( n1957 , n11358 );
    xnor g4948 ( n4444 , n8535 , n2410 );
    or g4949 ( n12165 , n4778 , n8655 );
    and g4950 ( n2535 , n9880 , n10801 );
    or g4951 ( n116 , n12195 , n4622 );
    or g4952 ( n9073 , n12186 , n7876 );
    or g4953 ( n7479 , n10748 , n2039 );
    or g4954 ( n7702 , n8046 , n4497 );
    xnor g4955 ( n6970 , n4206 , n4303 );
    not g4956 ( n3322 , n7267 );
    and g4957 ( n8973 , n6482 , n4586 );
    and g4958 ( n399 , n5754 , n1983 );
    xnor g4959 ( n11306 , n11718 , n350 );
    and g4960 ( n5301 , n8342 , n4051 );
    and g4961 ( n5930 , n4812 , n2573 );
    and g4962 ( n4906 , n1220 , n12621 );
    or g4963 ( n7363 , n4289 , n3035 );
    not g4964 ( n7397 , n5003 );
    not g4965 ( n2959 , n12178 );
    xnor g4966 ( n2038 , n583 , n6202 );
    xnor g4967 ( n3877 , n7416 , n950 );
    xnor g4968 ( n4174 , n1916 , n655 );
    nor g4969 ( n8448 , n4158 , n4407 );
    nor g4970 ( n9268 , n5728 , n6335 );
    xnor g4971 ( n4761 , n10361 , n12246 );
    nor g4972 ( n12474 , n862 , n8121 );
    and g4973 ( n12031 , n2464 , n8595 );
    nor g4974 ( n1434 , n4577 , n10423 );
    xnor g4975 ( n2776 , n9832 , n8657 );
    and g4976 ( n8238 , n6076 , n5169 );
    nor g4977 ( n7281 , n12871 , n5649 );
    nor g4978 ( n5253 , n5109 , n12295 );
    xnor g4979 ( n3217 , n12639 , n9823 );
    or g4980 ( n11805 , n3931 , n9720 );
    and g4981 ( n12438 , n4624 , n8281 );
    xnor g4982 ( n12641 , n1867 , n8734 );
    and g4983 ( n2105 , n92 , n4789 );
    or g4984 ( n6103 , n10842 , n5823 );
    and g4985 ( n7005 , n3382 , n8620 );
    and g4986 ( n203 , n1910 , n3114 );
    nor g4987 ( n8080 , n6773 , n9419 );
    and g4988 ( n535 , n5771 , n415 );
    and g4989 ( n7196 , n4562 , n12689 );
    xnor g4990 ( n12807 , n310 , n3008 );
    not g4991 ( n5929 , n6136 );
    and g4992 ( n4439 , n1345 , n6887 );
    and g4993 ( n10598 , n12280 , n2937 );
    not g4994 ( n10938 , n3016 );
    or g4995 ( n6795 , n4023 , n1870 );
    xnor g4996 ( n3851 , n8894 , n11774 );
    nor g4997 ( n12639 , n9936 , n2634 );
    nor g4998 ( n12486 , n7798 , n2194 );
    or g4999 ( n9498 , n10862 , n10421 );
    xnor g5000 ( n1268 , n5590 , n12406 );
    xnor g5001 ( n4251 , n8229 , n1276 );
    and g5002 ( n6529 , n7468 , n271 );
    nor g5003 ( n11510 , n6541 , n1219 );
    xnor g5004 ( n5232 , n925 , n10714 );
    xnor g5005 ( n7650 , n10000 , n6912 );
    and g5006 ( n11197 , n12775 , n12913 );
    xnor g5007 ( n10062 , n2602 , n2106 );
    and g5008 ( n7433 , n2483 , n4040 );
    or g5009 ( n11675 , n7449 , n8285 );
    or g5010 ( n7549 , n8583 , n9078 );
    xnor g5011 ( n6236 , n10438 , n12160 );
    or g5012 ( n12518 , n12659 , n6846 );
    or g5013 ( n1684 , n3767 , n7600 );
    and g5014 ( n2460 , n4693 , n5182 );
    xnor g5015 ( n2009 , n7102 , n7017 );
    xnor g5016 ( n10262 , n12747 , n8685 );
    xnor g5017 ( n9187 , n9770 , n2556 );
    and g5018 ( n5531 , n3992 , n10990 );
    xnor g5019 ( n977 , n10367 , n2164 );
    and g5020 ( n190 , n8929 , n11141 );
    xnor g5021 ( n7671 , n10711 , n6094 );
    nor g5022 ( n2362 , n6886 , n8213 );
    xnor g5023 ( n5161 , n9629 , n11870 );
    or g5024 ( n5995 , n10157 , n9280 );
    not g5025 ( n10835 , n7965 );
    and g5026 ( n7240 , n6442 , n10619 );
    and g5027 ( n9924 , n2959 , n1481 );
    xnor g5028 ( n2200 , n5026 , n4539 );
    not g5029 ( n641 , n12071 );
    or g5030 ( n6518 , n6718 , n9078 );
    xnor g5031 ( n10695 , n6665 , n8726 );
    or g5032 ( n2782 , n3402 , n3391 );
    nor g5033 ( n12804 , n12433 , n5417 );
    xnor g5034 ( n8122 , n12242 , n8909 );
    or g5035 ( n7369 , n6022 , n8427 );
    or g5036 ( n10983 , n9370 , n7424 );
    xnor g5037 ( n12939 , n10700 , n7435 );
    or g5038 ( n7145 , n4498 , n7703 );
    nor g5039 ( n6041 , n4635 , n12369 );
    nor g5040 ( n777 , n3726 , n8031 );
    and g5041 ( n12719 , n307 , n3471 );
    or g5042 ( n5407 , n8687 , n9521 );
    xnor g5043 ( n788 , n10343 , n9535 );
    or g5044 ( n925 , n8187 , n1079 );
    or g5045 ( n5826 , n1205 , n4282 );
    xnor g5046 ( n7842 , n12945 , n9859 );
    and g5047 ( n8370 , n7780 , n8901 );
    not g5048 ( n2317 , n8144 );
    xnor g5049 ( n10858 , n10365 , n8512 );
    xnor g5050 ( n9574 , n8130 , n9284 );
    not g5051 ( n7921 , n5814 );
    xnor g5052 ( n4440 , n7188 , n10807 );
    or g5053 ( n2168 , n2326 , n10869 );
    xnor g5054 ( n7911 , n11972 , n11732 );
    xnor g5055 ( n197 , n12012 , n3054 );
    or g5056 ( n7077 , n9900 , n5063 );
    or g5057 ( n5249 , n9844 , n7976 );
    or g5058 ( n10163 , n5372 , n4163 );
    xnor g5059 ( n12152 , n3188 , n5561 );
    not g5060 ( n10270 , n1354 );
    or g5061 ( n12936 , n4126 , n12608 );
    or g5062 ( n8637 , n10715 , n5316 );
    xnor g5063 ( n4133 , n578 , n8938 );
    or g5064 ( n10911 , n5774 , n10011 );
    not g5065 ( n12531 , n1837 );
    or g5066 ( n1495 , n1941 , n7558 );
    and g5067 ( n10498 , n5141 , n545 );
    or g5068 ( n587 , n505 , n12592 );
    or g5069 ( n8411 , n6204 , n11735 );
    and g5070 ( n7494 , n5981 , n5661 );
    and g5071 ( n5327 , n7476 , n10942 );
    not g5072 ( n4059 , n1097 );
    and g5073 ( n12047 , n12297 , n11611 );
    nor g5074 ( n3417 , n8733 , n5632 );
    and g5075 ( n12764 , n8476 , n6806 );
    or g5076 ( n9492 , n6977 , n995 );
    not g5077 ( n81 , n3205 );
    or g5078 ( n4562 , n3746 , n7558 );
    xnor g5079 ( n8275 , n8369 , n4284 );
    not g5080 ( n8629 , n10231 );
    and g5081 ( n2560 , n3352 , n1765 );
    and g5082 ( n8418 , n9996 , n6634 );
    or g5083 ( n5908 , n7709 , n1509 );
    nor g5084 ( n6005 , n10335 , n2378 );
    xnor g5085 ( n7152 , n6003 , n2919 );
    and g5086 ( n11460 , n10045 , n6345 );
    and g5087 ( n1760 , n12067 , n9214 );
    nor g5088 ( n4944 , n7300 , n9252 );
    and g5089 ( n10647 , n5465 , n6783 );
    xnor g5090 ( n11067 , n2877 , n7973 );
    and g5091 ( n23 , n1519 , n564 );
    xnor g5092 ( n801 , n1207 , n10696 );
    xnor g5093 ( n842 , n8998 , n8575 );
    xnor g5094 ( n10028 , n1516 , n2181 );
    and g5095 ( n10546 , n12023 , n7734 );
    xnor g5096 ( n5356 , n12282 , n4631 );
    xnor g5097 ( n2547 , n12728 , n340 );
    or g5098 ( n1276 , n636 , n10854 );
    nor g5099 ( n4033 , n10921 , n7522 );
    or g5100 ( n240 , n2217 , n9078 );
    not g5101 ( n3397 , n7735 );
    or g5102 ( n12626 , n7283 , n6389 );
    or g5103 ( n1605 , n8228 , n956 );
    and g5104 ( n5053 , n8336 , n7946 );
    nor g5105 ( n8017 , n5280 , n1801 );
    xnor g5106 ( n10009 , n3313 , n11809 );
    or g5107 ( n5209 , n1349 , n8258 );
    xnor g5108 ( n6614 , n451 , n9502 );
    nor g5109 ( n8223 , n5148 , n6675 );
    xnor g5110 ( n5934 , n917 , n7262 );
    and g5111 ( n12359 , n8074 , n735 );
    and g5112 ( n1327 , n6674 , n7075 );
    xnor g5113 ( n5052 , n12667 , n11737 );
    xnor g5114 ( n2662 , n1792 , n8636 );
    or g5115 ( n7035 , n12503 , n795 );
    or g5116 ( n7153 , n8764 , n8918 );
    and g5117 ( n9581 , n11473 , n6925 );
    xnor g5118 ( n7201 , n4863 , n7145 );
    nor g5119 ( n11269 , n9746 , n6586 );
    xnor g5120 ( n2540 , n9791 , n7905 );
    or g5121 ( n3791 , n10142 , n7246 );
    and g5122 ( n12421 , n77 , n8056 );
    and g5123 ( n5955 , n3605 , n9888 );
    xnor g5124 ( n4315 , n2586 , n2486 );
    or g5125 ( n9219 , n1076 , n3439 );
    xnor g5126 ( n3982 , n6597 , n6845 );
    and g5127 ( n10883 , n2031 , n650 );
    xnor g5128 ( n10950 , n9656 , n12411 );
    or g5129 ( n10282 , n5769 , n7239 );
    xnor g5130 ( n1555 , n7838 , n9135 );
    or g5131 ( n9100 , n11697 , n2985 );
    not g5132 ( n6718 , n8384 );
    nor g5133 ( n6829 , n9508 , n146 );
    or g5134 ( n183 , n11958 , n7395 );
    xnor g5135 ( n8825 , n6330 , n6996 );
    or g5136 ( n8813 , n7376 , n7465 );
    or g5137 ( n6544 , n9373 , n795 );
    nor g5138 ( n3798 , n12789 , n2355 );
    or g5139 ( n1879 , n11433 , n5012 );
    not g5140 ( n8687 , n5857 );
    xnor g5141 ( n9156 , n3944 , n1719 );
    nor g5142 ( n3052 , n11079 , n3847 );
    not g5143 ( n3501 , n927 );
    xnor g5144 ( n5708 , n290 , n4551 );
    and g5145 ( n8522 , n7778 , n7276 );
    not g5146 ( n8837 , n2921 );
    not g5147 ( n7015 , n6891 );
    or g5148 ( n7195 , n10966 , n7447 );
    not g5149 ( n9015 , n5846 );
    not g5150 ( n8113 , n8556 );
    xnor g5151 ( n7799 , n10912 , n6143 );
    or g5152 ( n10555 , n2217 , n11698 );
    or g5153 ( n10820 , n4778 , n12080 );
    not g5154 ( n9724 , n6343 );
    nor g5155 ( n4077 , n852 , n8335 );
    not g5156 ( n563 , n8927 );
    and g5157 ( n1648 , n3478 , n1104 );
    xnor g5158 ( n10700 , n1307 , n3239 );
    xnor g5159 ( n9209 , n11544 , n5944 );
    or g5160 ( n855 , n7116 , n9741 );
    or g5161 ( n3072 , n636 , n8655 );
    xnor g5162 ( n12387 , n4416 , n4253 );
    not g5163 ( n6197 , n8595 );
    and g5164 ( n7344 , n9066 , n11894 );
    or g5165 ( n7365 , n636 , n7928 );
    nor g5166 ( n9427 , n3222 , n12228 );
    nor g5167 ( n749 , n7253 , n12848 );
    not g5168 ( n11645 , n5808 );
    or g5169 ( n9374 , n11433 , n995 );
    not g5170 ( n10226 , n8851 );
    or g5171 ( n8467 , n8410 , n6101 );
    nor g5172 ( n10233 , n4759 , n1569 );
    and g5173 ( n7364 , n6559 , n2977 );
    and g5174 ( n785 , n3665 , n2452 );
    nor g5175 ( n4402 , n11591 , n9841 );
    or g5176 ( n2987 , n10847 , n12626 );
    nor g5177 ( n2702 , n8381 , n3163 );
    xnor g5178 ( n4273 , n10529 , n626 );
    and g5179 ( n12210 , n5081 , n3953 );
    not g5180 ( n10257 , n3795 );
    and g5181 ( n1407 , n4247 , n554 );
    not g5182 ( n8082 , n1408 );
    and g5183 ( n10921 , n10947 , n11800 );
    or g5184 ( n7618 , n8209 , n160 );
    nor g5185 ( n9969 , n5129 , n11770 );
    and g5186 ( n4062 , n6115 , n1566 );
    xnor g5187 ( n11737 , n10306 , n1042 );
    or g5188 ( n5514 , n4296 , n11865 );
    xnor g5189 ( n4494 , n5567 , n4959 );
    or g5190 ( n7156 , n338 , n11885 );
    xnor g5191 ( n8935 , n333 , n2955 );
    and g5192 ( n12001 , n3627 , n9956 );
    xnor g5193 ( n7047 , n1726 , n3718 );
    and g5194 ( n6109 , n7487 , n7752 );
    xnor g5195 ( n8014 , n8628 , n12625 );
    xnor g5196 ( n12537 , n1837 , n5565 );
    or g5197 ( n12846 , n1699 , n6513 );
    xnor g5198 ( n4999 , n1588 , n12677 );
    xnor g5199 ( n1853 , n3576 , n6403 );
    nor g5200 ( n12196 , n3516 , n11845 );
    not g5201 ( n889 , n4697 );
    or g5202 ( n7588 , n7758 , n1861 );
    xnor g5203 ( n1721 , n6229 , n3473 );
    and g5204 ( n1723 , n3445 , n10261 );
    and g5205 ( n11489 , n10661 , n5276 );
    nor g5206 ( n12109 , n9989 , n10408 );
    or g5207 ( n4950 , n7071 , n8338 );
    xnor g5208 ( n8131 , n11242 , n3597 );
    xnor g5209 ( n2057 , n5987 , n8723 );
    and g5210 ( n10181 , n12335 , n9743 );
    or g5211 ( n10804 , n9584 , n4527 );
    nor g5212 ( n2361 , n4564 , n4487 );
    or g5213 ( n6931 , n5765 , n3606 );
    xnor g5214 ( n12154 , n11219 , n4800 );
    xnor g5215 ( n6459 , n7267 , n11797 );
    xnor g5216 ( n8664 , n2855 , n8874 );
    xnor g5217 ( n9509 , n8208 , n5512 );
    not g5218 ( n9486 , n6423 );
    and g5219 ( n8630 , n2600 , n12332 );
    and g5220 ( n8799 , n9838 , n11645 );
    and g5221 ( n11027 , n8489 , n5696 );
    or g5222 ( n4287 , n7638 , n7419 );
    xnor g5223 ( n2158 , n6896 , n7636 );
    or g5224 ( n412 , n8584 , n12605 );
    xnor g5225 ( n10165 , n6116 , n4188 );
    and g5226 ( n9010 , n3992 , n6611 );
    or g5227 ( n2711 , n12443 , n1734 );
    and g5228 ( n12632 , n7397 , n11166 );
    or g5229 ( n3823 , n7577 , n5796 );
    or g5230 ( n7117 , n6373 , n12771 );
    xnor g5231 ( n4404 , n928 , n3650 );
    and g5232 ( n4135 , n5778 , n1591 );
    xnor g5233 ( n10037 , n12057 , n654 );
    or g5234 ( n404 , n373 , n10191 );
    xnor g5235 ( n11945 , n12854 , n7589 );
    or g5236 ( n8558 , n5951 , n5678 );
    not g5237 ( n9272 , n604 );
    not g5238 ( n12357 , n4190 );
    xnor g5239 ( n3132 , n10864 , n4198 );
    or g5240 ( n4283 , n8428 , n995 );
    or g5241 ( n11250 , n8428 , n3468 );
    xnor g5242 ( n8374 , n12692 , n11882 );
    xnor g5243 ( n2397 , n6561 , n10705 );
    and g5244 ( n3685 , n7393 , n12362 );
    and g5245 ( n1728 , n9792 , n7554 );
    and g5246 ( n12012 , n740 , n406 );
    or g5247 ( n2978 , n5809 , n8740 );
    and g5248 ( n972 , n10928 , n3719 );
    xnor g5249 ( n12159 , n6405 , n7440 );
    and g5250 ( n5170 , n3544 , n4715 );
    or g5251 ( n10652 , n6718 , n1509 );
    or g5252 ( n10896 , n5765 , n1509 );
    nor g5253 ( n10432 , n7457 , n872 );
    or g5254 ( n2482 , n12119 , n10311 );
    and g5255 ( n1845 , n713 , n96 );
    xnor g5256 ( n8667 , n650 , n2031 );
    not g5257 ( n10376 , n12880 );
    xnor g5258 ( n11529 , n10199 , n7637 );
    or g5259 ( n3202 , n10750 , n7928 );
    or g5260 ( n4931 , n8189 , n5797 );
    nor g5261 ( n11359 , n9697 , n1778 );
    xnor g5262 ( n2745 , n5219 , n3461 );
    not g5263 ( n11135 , n8467 );
    or g5264 ( n6284 , n2659 , n3186 );
    and g5265 ( n7023 , n3401 , n1996 );
    nor g5266 ( n9845 , n12760 , n2199 );
    xnor g5267 ( n6447 , n7866 , n2115 );
    xnor g5268 ( n9966 , n9068 , n9871 );
    and g5269 ( n5936 , n12584 , n5733 );
    and g5270 ( n12341 , n8789 , n1733 );
    xnor g5271 ( n10131 , n2172 , n11897 );
    or g5272 ( n11910 , n10750 , n10854 );
    nor g5273 ( n8986 , n8896 , n4710 );
    or g5274 ( n5111 , n697 , n1109 );
    and g5275 ( n5110 , n12380 , n4985 );
    nor g5276 ( n931 , n269 , n10924 );
    not g5277 ( n4104 , n5652 );
    xnor g5278 ( n5921 , n8469 , n2617 );
    xnor g5279 ( n8677 , n11578 , n975 );
    xnor g5280 ( n4399 , n12266 , n2438 );
    or g5281 ( n10771 , n11552 , n4527 );
    or g5282 ( n2896 , n9262 , n2020 );
    or g5283 ( n5183 , n1339 , n8940 );
    not g5284 ( n3213 , n7993 );
    and g5285 ( n10336 , n6358 , n11791 );
    and g5286 ( n9778 , n7993 , n5845 );
    xnor g5287 ( n12788 , n1520 , n8247 );
    and g5288 ( n7074 , n7236 , n10848 );
    not g5289 ( n6922 , n12247 );
    or g5290 ( n9836 , n5575 , n3421 );
    xnor g5291 ( n1770 , n8079 , n741 );
    xnor g5292 ( n1453 , n9555 , n10550 );
    or g5293 ( n4791 , n7283 , n7703 );
    xnor g5294 ( n12676 , n11287 , n11954 );
    or g5295 ( n10565 , n6373 , n9160 );
    xnor g5296 ( n6051 , n12718 , n234 );
    not g5297 ( n11072 , n11783 );
    or g5298 ( n11406 , n12361 , n11775 );
    and g5299 ( n2682 , n3141 , n4721 );
    xnor g5300 ( n1206 , n902 , n5829 );
    and g5301 ( n8672 , n2941 , n1567 );
    xnor g5302 ( n10765 , n11445 , n247 );
    or g5303 ( n3936 , n11026 , n5502 );
    or g5304 ( n6700 , n11607 , n10719 );
    xnor g5305 ( n6423 , n7206 , n11655 );
    xnor g5306 ( n6918 , n6628 , n1424 );
    xnor g5307 ( n5197 , n8996 , n4053 );
    or g5308 ( n10103 , n4791 , n5762 );
    and g5309 ( n9382 , n4411 , n10007 );
    xnor g5310 ( n3850 , n409 , n12094 );
    and g5311 ( n9031 , n12842 , n5654 );
    xnor g5312 ( n8652 , n8979 , n4334 );
    or g5313 ( n3081 , n6695 , n6006 );
    not g5314 ( n1559 , n2752 );
    nor g5315 ( n8012 , n11366 , n7237 );
    nor g5316 ( n5672 , n12024 , n8821 );
    xnor g5317 ( n8602 , n4385 , n7266 );
    or g5318 ( n1773 , n7540 , n3055 );
    or g5319 ( n12730 , n11887 , n7382 );
    nor g5320 ( n612 , n11369 , n2990 );
    not g5321 ( n1171 , n10788 );
    nor g5322 ( n7624 , n5898 , n633 );
    not g5323 ( n10396 , n3579 );
    or g5324 ( n7141 , n1784 , n11355 );
    or g5325 ( n3570 , n5575 , n3356 );
    xnor g5326 ( n532 , n1912 , n2546 );
    not g5327 ( n5044 , n1397 );
    and g5328 ( n960 , n2987 , n6214 );
    not g5329 ( n4924 , n2180 );
    and g5330 ( n12796 , n7316 , n9090 );
    not g5331 ( n17 , n4923 );
    xnor g5332 ( n7332 , n225 , n8039 );
    xnor g5333 ( n12903 , n5441 , n1862 );
    or g5334 ( n4536 , n2456 , n4818 );
    and g5335 ( n1632 , n2532 , n4802 );
    xnor g5336 ( n12884 , n5799 , n801 );
    or g5337 ( n5202 , n6577 , n11410 );
    or g5338 ( n12144 , n5530 , n1932 );
    or g5339 ( n4815 , n9878 , n9188 );
    and g5340 ( n10004 , n10282 , n3409 );
    xnor g5341 ( n12657 , n9029 , n3500 );
    xnor g5342 ( n2746 , n7516 , n3809 );
    and g5343 ( n11040 , n9241 , n6703 );
    or g5344 ( n6981 , n5765 , n11698 );
    or g5345 ( n3631 , n4343 , n826 );
    not g5346 ( n4911 , n12705 );
    xnor g5347 ( n3443 , n11348 , n472 );
    and g5348 ( n3286 , n10365 , n10723 );
    or g5349 ( n2677 , n5575 , n7425 );
    and g5350 ( n9737 , n3325 , n1386 );
    or g5351 ( n432 , n2217 , n4875 );
    or g5352 ( n8882 , n5915 , n10854 );
    nor g5353 ( n4316 , n1256 , n3254 );
    and g5354 ( n12551 , n1403 , n765 );
    xnor g5355 ( n12319 , n5965 , n169 );
    not g5356 ( n12501 , n2111 );
    or g5357 ( n10438 , n7197 , n8069 );
    not g5358 ( n12640 , n3732 );
    or g5359 ( n69 , n1438 , n2409 );
    or g5360 ( n7961 , n4716 , n7 );
    xnor g5361 ( n9423 , n11838 , n7344 );
    or g5362 ( n3810 , n12237 , n7382 );
    and g5363 ( n7945 , n7807 , n1412 );
    not g5364 ( n1612 , n2519 );
    or g5365 ( n10356 , n595 , n9449 );
    or g5366 ( n12053 , n4059 , n7341 );
    or g5367 ( n8452 , n6373 , n9568 );
    xnor g5368 ( n11325 , n4771 , n5082 );
    nor g5369 ( n4765 , n11961 , n1090 );
    or g5370 ( n3967 , n8552 , n826 );
    and g5371 ( n1595 , n10180 , n4234 );
    not g5372 ( n12130 , n6725 );
    or g5373 ( n964 , n8687 , n9160 );
    or g5374 ( n12825 , n11282 , n3517 );
    and g5375 ( n6541 , n1018 , n6093 );
    xnor g5376 ( n12713 , n9115 , n11924 );
    xnor g5377 ( n1202 , n8857 , n7842 );
    nor g5378 ( n7660 , n4819 , n10515 );
    xnor g5379 ( n9264 , n3198 , n7596 );
    not g5380 ( n9142 , n7027 );
    or g5381 ( n7859 , n5971 , n8824 );
    xnor g5382 ( n3149 , n4535 , n501 );
    xnor g5383 ( n1609 , n2109 , n859 );
    not g5384 ( n9327 , n3990 );
    and g5385 ( n3231 , n6130 , n6708 );
    and g5386 ( n10429 , n10673 , n8926 );
    and g5387 ( n12950 , n12210 , n601 );
    or g5388 ( n1874 , n5765 , n4864 );
    xnor g5389 ( n3148 , n10798 , n10707 );
    or g5390 ( n616 , n7284 , n10144 );
    xnor g5391 ( n671 , n10853 , n11300 );
    xnor g5392 ( n2086 , n553 , n4133 );
    or g5393 ( n5024 , n11026 , n4474 );
    nor g5394 ( n11107 , n202 , n9086 );
    or g5395 ( n6869 , n5110 , n2795 );
    or g5396 ( n7584 , n9304 , n8148 );
    or g5397 ( n315 , n5664 , n2145 );
    or g5398 ( n1401 , n2154 , n6459 );
    not g5399 ( n9243 , n11225 );
    or g5400 ( n3861 , n1891 , n11920 );
    or g5401 ( n1212 , n1960 , n1019 );
    or g5402 ( n3297 , n9370 , n6402 );
    or g5403 ( n3300 , n8405 , n9188 );
    or g5404 ( n12046 , n8870 , n8648 );
    or g5405 ( n9496 , n8687 , n4474 );
    or g5406 ( n6471 , n11598 , n5096 );
    or g5407 ( n9681 , n5348 , n581 );
    xnor g5408 ( n4006 , n2937 , n1297 );
    xnor g5409 ( n9338 , n11968 , n6 );
    or g5410 ( n5893 , n6221 , n9851 );
    not g5411 ( n3578 , n3003 );
    not g5412 ( n12745 , n9381 );
    not g5413 ( n10475 , n10394 );
    or g5414 ( n856 , n6977 , n10919 );
    or g5415 ( n12524 , n3617 , n6513 );
    or g5416 ( n3777 , n11032 , n12830 );
    or g5417 ( n9834 , n1937 , n11820 );
    xnor g5418 ( n6502 , n11937 , n1547 );
    xnor g5419 ( n6989 , n100 , n12100 );
    and g5420 ( n4632 , n3494 , n2646 );
    not g5421 ( n8749 , n1304 );
    and g5422 ( n11275 , n9858 , n10972 );
    or g5423 ( n12554 , n5602 , n2463 );
    or g5424 ( n4247 , n7449 , n8830 );
    xnor g5425 ( n5965 , n1010 , n5187 );
    not g5426 ( n8509 , n2533 );
    or g5427 ( n10224 , n4535 , n501 );
    or g5428 ( n9119 , n12324 , n2736 );
    xnor g5429 ( n8402 , n730 , n4345 );
    and g5430 ( n499 , n9093 , n5682 );
    and g5431 ( n7520 , n9886 , n3370 );
    xnor g5432 ( n155 , n2826 , n758 );
    xnor g5433 ( n7515 , n6365 , n9702 );
    nor g5434 ( n9034 , n6512 , n12681 );
    not g5435 ( n4643 , n8580 );
    xnor g5436 ( n9096 , n946 , n3258 );
    xnor g5437 ( n6187 , n8339 , n9540 );
    xnor g5438 ( n225 , n8448 , n10161 );
    not g5439 ( n1700 , n3531 );
    not g5440 ( n2099 , n5331 );
    not g5441 ( n4100 , n12582 );
    not g5442 ( n4853 , n8324 );
    xnor g5443 ( n4009 , n6813 , n4156 );
    or g5444 ( n10504 , n5575 , n7395 );
    or g5445 ( n2525 , n12361 , n12816 );
    or g5446 ( n9048 , n7116 , n7952 );
    and g5447 ( n9907 , n8750 , n10537 );
    not g5448 ( n3115 , n1017 );
    or g5449 ( n5151 , n10118 , n5887 );
    nor g5450 ( n7448 , n8044 , n8319 );
    xnor g5451 ( n6453 , n10008 , n8494 );
    not g5452 ( n3989 , n11563 );
    or g5453 ( n7642 , n2407 , n12137 );
    xnor g5454 ( n5270 , n7953 , n12148 );
    xnor g5455 ( n5078 , n7531 , n9259 );
    or g5456 ( n7414 , n10677 , n5079 );
    or g5457 ( n12390 , n1169 , n4891 );
    or g5458 ( n6062 , n7984 , n1541 );
    xnor g5459 ( n1414 , n5260 , n1108 );
    xnor g5460 ( n2996 , n2120 , n12885 );
    not g5461 ( n5538 , n4141 );
    not g5462 ( n11698 , n4903 );
    and g5463 ( n6460 , n1534 , n8112 );
    not g5464 ( n8951 , n1646 );
    not g5465 ( n4434 , n12723 );
    or g5466 ( n4728 , n5575 , n7558 );
    or g5467 ( n5354 , n4568 , n12558 );
    xnor g5468 ( n11527 , n1456 , n8842 );
    or g5469 ( n3938 , n12633 , n6508 );
    or g5470 ( n326 , n5989 , n6704 );
    nor g5471 ( n6828 , n12430 , n6281 );
    or g5472 ( n8698 , n4422 , n12809 );
    and g5473 ( n11688 , n5619 , n7308 );
    xnor g5474 ( n7048 , n7474 , n7654 );
    xnor g5475 ( n12364 , n2536 , n2670 );
    and g5476 ( n2420 , n2011 , n4899 );
    and g5477 ( n11659 , n8304 , n10469 );
    or g5478 ( n6239 , n11958 , n6455 );
    nor g5479 ( n6399 , n8781 , n4330 );
    and g5480 ( n3254 , n2506 , n11807 );
    or g5481 ( n3583 , n7384 , n2005 );
    not g5482 ( n11976 , n6303 );
    and g5483 ( n105 , n11037 , n10573 );
    and g5484 ( n7795 , n8510 , n8274 );
    and g5485 ( n11420 , n10202 , n9729 );
    and g5486 ( n3834 , n5419 , n11619 );
    and g5487 ( n11656 , n3176 , n8167 );
    xnor g5488 ( n6357 , n9414 , n2038 );
    or g5489 ( n7319 , n9081 , n6258 );
    xnor g5490 ( n12450 , n8304 , n190 );
    or g5491 ( n7780 , n10761 , n3234 );
    or g5492 ( n4585 , n4725 , n12396 );
    or g5493 ( n6924 , n10750 , n7382 );
    not g5494 ( n1344 , n165 );
    xnor g5495 ( n10221 , n8436 , n86 );
    or g5496 ( n4150 , n11694 , n4377 );
    nor g5497 ( n12927 , n6566 , n4542 );
    or g5498 ( n483 , n9621 , n1490 );
    xnor g5499 ( n652 , n4962 , n10016 );
    xnor g5500 ( n642 , n296 , n6837 );
    xnor g5501 ( n952 , n9134 , n5775 );
    xnor g5502 ( n7066 , n6659 , n7524 );
    xnor g5503 ( n10687 , n9445 , n4567 );
    xnor g5504 ( n6400 , n474 , n1556 );
    xnor g5505 ( n3230 , n12359 , n94 );
    and g5506 ( n2231 , n8730 , n5588 );
    xnor g5507 ( n7988 , n5881 , n9979 );
    not g5508 ( n4169 , n11628 );
    or g5509 ( n6295 , n8838 , n8029 );
    or g5510 ( n7770 , n5600 , n2793 );
    nor g5511 ( n984 , n6076 , n5169 );
    not g5512 ( n3712 , n5495 );
    or g5513 ( n4571 , n955 , n5442 );
    and g5514 ( n1828 , n4956 , n5000 );
    or g5515 ( n6352 , n6290 , n11439 );
    nor g5516 ( n3454 , n12422 , n8568 );
    nor g5517 ( n9128 , n2532 , n4802 );
    and g5518 ( n10895 , n3065 , n577 );
    or g5519 ( n2137 , n11417 , n1314 );
    or g5520 ( n11597 , n10101 , n2218 );
    xnor g5521 ( n1858 , n9969 , n7604 );
    not g5522 ( n2815 , n7946 );
    xnor g5523 ( n5332 , n3608 , n11467 );
    or g5524 ( n10626 , n11037 , n10573 );
    or g5525 ( n4548 , n10564 , n9733 );
    or g5526 ( n4560 , n11390 , n3431 );
    xnor g5527 ( n9409 , n4536 , n4220 );
    and g5528 ( n7329 , n7404 , n11438 );
    or g5529 ( n3841 , n5913 , n2751 );
    xnor g5530 ( n11393 , n9942 , n2477 );
    nor g5531 ( n3788 , n8557 , n7653 );
    not g5532 ( n5763 , n12115 );
    not g5533 ( n1122 , n2413 );
    or g5534 ( n1862 , n1699 , n8740 );
    and g5535 ( n2768 , n11621 , n11956 );
    not g5536 ( n1739 , n6431 );
    xnor g5537 ( n4996 , n1960 , n1019 );
    nor g5538 ( n3355 , n11992 , n1293 );
    xnor g5539 ( n2410 , n195 , n12049 );
    not g5540 ( n12878 , n2038 );
    or g5541 ( n131 , n11601 , n10724 );
    and g5542 ( n4482 , n7474 , n1681 );
    and g5543 ( n4398 , n3549 , n98 );
    xnor g5544 ( n6733 , n1804 , n1105 );
    xnor g5545 ( n8381 , n5202 , n12240 );
    not g5546 ( n4423 , n302 );
    not g5547 ( n3714 , n1716 );
    or g5548 ( n4126 , n11958 , n10919 );
    not g5549 ( n5410 , n8940 );
    xnor g5550 ( n12702 , n8864 , n8788 );
    or g5551 ( n3908 , n3891 , n8409 );
    or g5552 ( n11517 , n11958 , n12357 );
    not g5553 ( n2762 , n11553 );
    nor g5554 ( n10149 , n7248 , n12159 );
    or g5555 ( n77 , n8227 , n10209 );
    and g5556 ( n4282 , n12195 , n4622 );
    xnor g5557 ( n1430 , n4910 , n4361 );
    or g5558 ( n2182 , n994 , n2076 );
    or g5559 ( n12015 , n686 , n5012 );
    or g5560 ( n4532 , n2078 , n10596 );
    or g5561 ( n7843 , n12632 , n10244 );
    or g5562 ( n7202 , n2626 , n4041 );
    and g5563 ( n6034 , n2288 , n1145 );
    xnor g5564 ( n10859 , n9744 , n3963 );
    and g5565 ( n8203 , n9748 , n10395 );
    nor g5566 ( n4563 , n3463 , n8178 );
    or g5567 ( n7756 , n4498 , n1851 );
    nor g5568 ( n10277 , n8277 , n12370 );
    or g5569 ( n7168 , n6595 , n6639 );
    xnor g5570 ( n364 , n3551 , n12205 );
    xnor g5571 ( n4227 , n3210 , n11192 );
    xnor g5572 ( n5123 , n2155 , n5786 );
    or g5573 ( n8311 , n4768 , n9619 );
    xnor g5574 ( n2206 , n5618 , n1430 );
    xnor g5575 ( n5762 , n12913 , n12239 );
    nor g5576 ( n11817 , n3106 , n11945 );
    not g5577 ( n8807 , n3465 );
    and g5578 ( n5023 , n674 , n10606 );
    or g5579 ( n401 , n10852 , n12019 );
    or g5580 ( n10162 , n2756 , n327 );
    and g5581 ( n11990 , n8984 , n12268 );
    not g5582 ( n4216 , n4275 );
    or g5583 ( n2041 , n12157 , n11197 );
    not g5584 ( n10514 , n10711 );
    or g5585 ( n7764 , n12503 , n4654 );
    and g5586 ( n7305 , n6242 , n8791 );
    or g5587 ( n8679 , n2526 , n8491 );
    and g5588 ( n10193 , n705 , n1310 );
    xnor g5589 ( n10558 , n12880 , n2690 );
    nor g5590 ( n7848 , n8713 , n6850 );
    and g5591 ( n5792 , n4932 , n12548 );
    xnor g5592 ( n2567 , n2686 , n10618 );
    xnor g5593 ( n8252 , n8011 , n10518 );
    not g5594 ( n1488 , n11227 );
    and g5595 ( n8435 , n4637 , n11288 );
    not g5596 ( n2748 , n5916 );
    nor g5597 ( n6449 , n5177 , n10438 );
    and g5598 ( n10775 , n677 , n7811 );
    xnor g5599 ( n8491 , n6258 , n12412 );
    or g5600 ( n9787 , n11026 , n2020 );
    xnor g5601 ( n2235 , n9109 , n6207 );
    xnor g5602 ( n9084 , n1961 , n6791 );
    not g5603 ( n8796 , n3179 );
    or g5604 ( n1920 , n1266 , n2090 );
    and g5605 ( n8261 , n3126 , n188 );
    and g5606 ( n12905 , n7998 , n4153 );
    not g5607 ( n8722 , n9541 );
    xnor g5608 ( n8593 , n5024 , n5255 );
    and g5609 ( n1489 , n3050 , n11524 );
    xnor g5610 ( n11566 , n7572 , n7394 );
    not g5611 ( n5954 , n5967 );
    xnor g5612 ( n11030 , n7761 , n3259 );
    or g5613 ( n2011 , n4628 , n12754 );
    or g5614 ( n5685 , n3743 , n9144 );
    and g5615 ( n8083 , n1471 , n8433 );
    or g5616 ( n638 , n12119 , n530 );
    or g5617 ( n991 , n5530 , n7382 );
    xnor g5618 ( n4829 , n7148 , n8106 );
    or g5619 ( n12781 , n5575 , n12274 );
    or g5620 ( n4380 , n10142 , n7703 );
    or g5621 ( n913 , n6977 , n11122 );
    xnor g5622 ( n9121 , n597 , n1289 );
    or g5623 ( n12879 , n1051 , n11820 );
    and g5624 ( n4064 , n6534 , n10826 );
    or g5625 ( n11024 , n8127 , n4400 );
    or g5626 ( n12561 , n12669 , n6360 );
    not g5627 ( n12946 , n8353 );
    and g5628 ( n12712 , n996 , n11791 );
    and g5629 ( n10033 , n1727 , n12514 );
    and g5630 ( n796 , n5341 , n11947 );
    or g5631 ( n3550 , n1153 , n55 );
    nor g5632 ( n869 , n3440 , n5755 );
    nor g5633 ( n2998 , n436 , n3299 );
    xnor g5634 ( n6342 , n6293 , n9157 );
    and g5635 ( n1655 , n12110 , n1133 );
    and g5636 ( n2497 , n7864 , n8099 );
    xnor g5637 ( n5487 , n8299 , n10860 );
    xnor g5638 ( n5028 , n9719 , n11529 );
    or g5639 ( n1382 , n12622 , n3919 );
    nor g5640 ( n11584 , n6813 , n10871 );
    and g5641 ( n2309 , n12200 , n6975 );
    xnor g5642 ( n10029 , n12765 , n8664 );
    xnor g5643 ( n12674 , n205 , n11965 );
    or g5644 ( n10869 , n6373 , n28 );
    or g5645 ( n8536 , n191 , n8970 );
    and g5646 ( n8136 , n8423 , n7315 );
    or g5647 ( n5890 , n9222 , n342 );
    xnor g5648 ( n5009 , n9480 , n6956 );
    or g5649 ( n4650 , n11887 , n3224 );
    or g5650 ( n7491 , n12119 , n7136 );
    and g5651 ( n12636 , n4266 , n3626 );
    or g5652 ( n3462 , n7495 , n1162 );
    and g5653 ( n9426 , n1808 , n2210 );
    or g5654 ( n7404 , n8348 , n12282 );
    not g5655 ( n543 , n7530 );
    or g5656 ( n3620 , n4059 , n1079 );
    or g5657 ( n11869 , n383 , n10621 );
    or g5658 ( n3671 , n10339 , n10854 );
    or g5659 ( n10915 , n6461 , n3148 );
    not g5660 ( n6221 , n4868 );
    not g5661 ( n5223 , n2629 );
    nor g5662 ( n10058 , n1061 , n12022 );
    xnor g5663 ( n1296 , n4986 , n4810 );
    not g5664 ( n12138 , n6816 );
    xnor g5665 ( n6716 , n6894 , n1616 );
    nor g5666 ( n11859 , n4389 , n6680 );
    nor g5667 ( n7521 , n5644 , n7220 );
    not g5668 ( n1782 , n12764 );
    or g5669 ( n1405 , n3285 , n2738 );
    xnor g5670 ( n9298 , n3374 , n11789 );
    and g5671 ( n8247 , n4953 , n8301 );
    or g5672 ( n2925 , n11689 , n11058 );
    or g5673 ( n12747 , n3743 , n4654 );
    and g5674 ( n2475 , n7504 , n224 );
    xnor g5675 ( n5822 , n10402 , n3249 );
    and g5676 ( n12616 , n11556 , n6173 );
    xnor g5677 ( n963 , n2893 , n1014 );
    or g5678 ( n8619 , n3804 , n1700 );
    or g5679 ( n10886 , n5945 , n3903 );
    xnor g5680 ( n4017 , n10839 , n600 );
    or g5681 ( n10893 , n6717 , n5867 );
    not g5682 ( n8059 , n4700 );
    xnor g5683 ( n3188 , n12734 , n1283 );
    or g5684 ( n8489 , n9570 , n12050 );
    nor g5685 ( n2148 , n688 , n7853 );
    or g5686 ( n11557 , n5355 , n1455 );
    nor g5687 ( n6198 , n5234 , n9597 );
    not g5688 ( n2380 , n3083 );
    xnor g5689 ( n6612 , n7312 , n8718 );
    or g5690 ( n1606 , n636 , n8259 );
    or g5691 ( n3728 , n1511 , n7602 );
    xnor g5692 ( n6980 , n3005 , n9251 );
    nor g5693 ( n2114 , n3201 , n10782 );
    not g5694 ( n8246 , n9454 );
    or g5695 ( n12433 , n12503 , n12771 );
    xnor g5696 ( n4570 , n10481 , n6480 );
    xnor g5697 ( n11006 , n5064 , n8974 );
    not g5698 ( n3482 , n2871 );
    or g5699 ( n3076 , n12361 , n7876 );
    xnor g5700 ( n4757 , n8573 , n9691 );
    nor g5701 ( n10076 , n5364 , n9781 );
    and g5702 ( n12586 , n2597 , n934 );
    xnor g5703 ( n11270 , n6242 , n2469 );
    not g5704 ( n149 , n2913 );
    and g5705 ( n160 , n5710 , n12926 );
    not g5706 ( n576 , n7726 );
    xnor g5707 ( n9706 , n4427 , n1110 );
    or g5708 ( n7932 , n8545 , n12783 );
    and g5709 ( n9585 , n7662 , n1800 );
    and g5710 ( n330 , n7919 , n5872 );
    or g5711 ( n9976 , n12237 , n6513 );
    or g5712 ( n2714 , n6977 , n11896 );
    and g5713 ( n4618 , n8348 , n12282 );
    or g5714 ( n11782 , n7449 , n5258 );
    not g5715 ( n4518 , n11623 );
    or g5716 ( n7754 , n3746 , n6114 );
    nor g5717 ( n12410 , n10401 , n8771 );
    nor g5718 ( n90 , n5995 , n769 );
    or g5719 ( n4872 , n2089 , n7962 );
    and g5720 ( n3264 , n12025 , n9956 );
    xnor g5721 ( n4345 , n5503 , n12844 );
    and g5722 ( n5596 , n4958 , n5514 );
    or g5723 ( n7112 , n4498 , n3911 );
    or g5724 ( n1803 , n10142 , n11430 );
    xnor g5725 ( n2250 , n6702 , n9901 );
    xnor g5726 ( n3203 , n6582 , n10121 );
    and g5727 ( n9288 , n11294 , n7507 );
    and g5728 ( n8125 , n5377 , n6701 );
    xnor g5729 ( n1431 , n6994 , n1538 );
    not g5730 ( n7742 , n2094 );
    nor g5731 ( n11261 , n9165 , n2729 );
    or g5732 ( n11581 , n11433 , n3903 );
    xnor g5733 ( n11738 , n9699 , n2084 );
    xnor g5734 ( n9679 , n6137 , n3901 );
    nor g5735 ( n11000 , n1177 , n5354 );
    xnor g5736 ( n2752 , n10480 , n1173 );
    and g5737 ( n12198 , n7685 , n3179 );
    not g5738 ( n7007 , n4241 );
    or g5739 ( n3221 , n5355 , n8859 );
    and g5740 ( n3234 , n348 , n5667 );
    not g5741 ( n4925 , n9390 );
    and g5742 ( n3330 , n9070 , n9786 );
    and g5743 ( n4488 , n8291 , n3104 );
    or g5744 ( n453 , n8674 , n5642 );
    or g5745 ( n769 , n6718 , n1476 );
    xnor g5746 ( n8876 , n10443 , n5544 );
    xnor g5747 ( n4905 , n10568 , n133 );
    not g5748 ( n10736 , n3294 );
    xnor g5749 ( n6135 , n12428 , n7210 );
    xnor g5750 ( n11558 , n3684 , n12333 );
    not g5751 ( n8109 , n7159 );
    xnor g5752 ( n6179 , n4468 , n3034 );
    not g5753 ( n6378 , n4953 );
    or g5754 ( n6256 , n4628 , n1163 );
    xnor g5755 ( n6773 , n6688 , n6255 );
    and g5756 ( n3693 , n8692 , n2421 );
    and g5757 ( n2210 , n2786 , n9009 );
    and g5758 ( n9140 , n2584 , n9258 );
    xnor g5759 ( n6262 , n5018 , n12593 );
    and g5760 ( n11649 , n9825 , n8469 );
    xor g5761 ( n10766 , n5209 , n7241 );
    xnor g5762 ( n1167 , n11864 , n11458 );
    and g5763 ( n9615 , n857 , n6691 );
    or g5764 ( n11176 , n4059 , n7246 );
    and g5765 ( n2469 , n1397 , n8359 );
    not g5766 ( n11483 , n9351 );
    or g5767 ( n6801 , n11958 , n9971 );
    not g5768 ( n5086 , n12511 );
    or g5769 ( n9292 , n3567 , n11440 );
    xnor g5770 ( n4954 , n7906 , n4338 );
    or g5771 ( n4183 , n3746 , n5540 );
    or g5772 ( n5466 , n2099 , n4818 );
    not g5773 ( n7573 , n9838 );
    xnor g5774 ( n9361 , n24 , n7334 );
    or g5775 ( n2864 , n5743 , n7840 );
    or g5776 ( n6837 , n7709 , n28 );
    not g5777 ( n2683 , n544 );
    and g5778 ( n3826 , n2137 , n4335 );
    xnor g5779 ( n3475 , n0 , n2127 );
    and g5780 ( n12050 , n1212 , n3039 );
    and g5781 ( n10782 , n5899 , n2928 );
    xnor g5782 ( n10116 , n6935 , n12438 );
    xnor g5783 ( n5062 , n11642 , n8562 );
    xnor g5784 ( n289 , n2714 , n7125 );
    or g5785 ( n8818 , n7084 , n9091 );
    xnor g5786 ( n2673 , n6301 , n2823 );
    and g5787 ( n539 , n4769 , n8956 );
    and g5788 ( n2058 , n3014 , n9939 );
    and g5789 ( n5975 , n9036 , n8225 );
    xnor g5790 ( n5728 , n496 , n2939 );
    xnor g5791 ( n56 , n8342 , n5900 );
    or g5792 ( n11183 , n1054 , n12657 );
    and g5793 ( n324 , n5378 , n8697 );
    or g5794 ( n10323 , n8959 , n1413 );
    xnor g5795 ( n2912 , n12478 , n7759 );
    or g5796 ( n5250 , n8847 , n9356 );
    and g5797 ( n5931 , n5291 , n11040 );
    or g5798 ( n12306 , n1051 , n5540 );
    not g5799 ( n9761 , n2742 );
    or g5800 ( n6666 , n5456 , n87 );
    or g5801 ( n12597 , n12361 , n8768 );
    or g5802 ( n8574 , n969 , n5046 );
    xnor g5803 ( n251 , n11285 , n33 );
    or g5804 ( n1620 , n686 , n9741 );
    or g5805 ( n11691 , n9082 , n10865 );
    nor g5806 ( n6496 , n12318 , n6900 );
    not g5807 ( n11088 , n4145 );
    and g5808 ( n1251 , n10392 , n10911 );
    and g5809 ( n9870 , n1642 , n12325 );
    or g5810 ( n5828 , n5355 , n1915 );
    xnor g5811 ( n12824 , n1418 , n8941 );
    or g5812 ( n7883 , n9370 , n4400 );
    nor g5813 ( n11635 , n12479 , n8174 );
    not g5814 ( n994 , n1333 );
    nor g5815 ( n11092 , n5368 , n2221 );
    and g5816 ( n8943 , n5394 , n5152 );
    nor g5817 ( n5904 , n6149 , n3454 );
    xnor g5818 ( n6419 , n3930 , n4483 );
    or g5819 ( n4116 , n6977 , n3903 );
    or g5820 ( n10352 , n8738 , n1509 );
    or g5821 ( n3461 , n4628 , n10854 );
    xnor g5822 ( n9628 , n4857 , n2310 );
    or g5823 ( n6820 , n636 , n12754 );
    or g5824 ( n5055 , n8187 , n11746 );
    xnor g5825 ( n11986 , n1657 , n9030 );
    nor g5826 ( n6598 , n2783 , n1531 );
    xnor g5827 ( n7412 , n7221 , n10500 );
    not g5828 ( n5296 , n6188 );
    or g5829 ( n11344 , n10953 , n9999 );
    and g5830 ( n9275 , n7431 , n1175 );
    xnor g5831 ( n1063 , n9834 , n11043 );
    and g5832 ( n5188 , n12053 , n4464 );
    not g5833 ( n7789 , n9311 );
    not g5834 ( n3644 , n11908 );
    xnor g5835 ( n8030 , n5805 , n11447 );
    xnor g5836 ( n1814 , n8084 , n11976 );
    xnor g5837 ( n924 , n4272 , n11833 );
    or g5838 ( n8132 , n2472 , n11952 );
    and g5839 ( n3956 , n504 , n3873 );
    not g5840 ( n6270 , n12537 );
    not g5841 ( n10871 , n1385 );
    or g5842 ( n562 , n5982 , n9166 );
    not g5843 ( n6206 , n6748 );
    nor g5844 ( n10680 , n9134 , n10397 );
    or g5845 ( n10912 , n2217 , n10916 );
    and g5846 ( n4091 , n3552 , n7061 );
    or g5847 ( n8474 , n1699 , n8648 );
    xnor g5848 ( n5043 , n8917 , n5487 );
    nor g5849 ( n12082 , n10432 , n154 );
    and g5850 ( n10052 , n7050 , n2106 );
    xnor g5851 ( n3677 , n4720 , n11918 );
    and g5852 ( n7712 , n8308 , n6581 );
    nor g5853 ( n2944 , n384 , n5972 );
    and g5854 ( n9802 , n7493 , n8551 );
    xnor g5855 ( n5768 , n5972 , n384 );
    not g5856 ( n4753 , n4960 );
    nor g5857 ( n4979 , n6951 , n12081 );
    xnor g5858 ( n7857 , n10104 , n4835 );
    xnor g5859 ( n12113 , n12456 , n12743 );
    xnor g5860 ( n11039 , n11351 , n6023 );
    or g5861 ( n1225 , n7551 , n10825 );
    and g5862 ( n640 , n12177 , n12386 );
    or g5863 ( n9727 , n4628 , n9188 );
    or g5864 ( n9122 , n12119 , n8655 );
    or g5865 ( n4755 , n5530 , n10311 );
    not g5866 ( n5530 , n12069 );
    or g5867 ( n497 , n7266 , n4385 );
    xnor g5868 ( n12282 , n3967 , n5927 );
    or g5869 ( n2717 , n3096 , n5012 );
    xnor g5870 ( n7361 , n107 , n11005 );
    xnor g5871 ( n7368 , n9274 , n12513 );
    or g5872 ( n5546 , n3642 , n10963 );
    not g5873 ( n12813 , n3258 );
    or g5874 ( n3629 , n276 , n3507 );
    or g5875 ( n6746 , n7191 , n942 );
    xnor g5876 ( n3613 , n3747 , n1561 );
    nor g5877 ( n8190 , n5202 , n9513 );
    nor g5878 ( n6972 , n6788 , n1214 );
    or g5879 ( n1398 , n8738 , n4875 );
    and g5880 ( n12487 , n507 , n2797 );
    and g5881 ( n3707 , n8390 , n2744 );
    not g5882 ( n6547 , n10531 );
    or g5883 ( n12945 , n10750 , n12124 );
    not g5884 ( n7389 , n9583 );
    or g5885 ( n7140 , n9268 , n11706 );
    or g5886 ( n4336 , n686 , n11820 );
    and g5887 ( n5627 , n4529 , n8749 );
    or g5888 ( n3392 , n9170 , n1546 );
    and g5889 ( n11855 , n11390 , n3431 );
    xnor g5890 ( n1999 , n9931 , n7926 );
    not g5891 ( n1937 , n11311 );
    nor g5892 ( n5678 , n6208 , n5878 );
    xnor g5893 ( n8494 , n2056 , n2595 );
    xnor g5894 ( n8235 , n10421 , n11367 );
    not g5895 ( n5008 , n555 );
    xnor g5896 ( n700 , n1202 , n10115 );
    nor g5897 ( n1006 , n6442 , n10619 );
    xnor g5898 ( n2088 , n3810 , n3181 );
    or g5899 ( n11449 , n4304 , n1117 );
    xnor g5900 ( n5640 , n8296 , n1427 );
    not g5901 ( n7928 , n6016 );
    and g5902 ( n8504 , n2530 , n7610 );
    xnor g5903 ( n4309 , n11039 , n6641 );
    or g5904 ( n8000 , n1699 , n2964 );
    not g5905 ( n6977 , n6986 );
    and g5906 ( n6535 , n393 , n7260 );
    nor g5907 ( n10388 , n7890 , n9162 );
    and g5908 ( n12864 , n5016 , n12202 );
    not g5909 ( n8040 , n308 );
    and g5910 ( n6960 , n5505 , n5009 );
    not g5911 ( n10655 , n8538 );
    or g5912 ( n5681 , n5809 , n8655 );
    or g5913 ( n1919 , n6373 , n9078 );
    xnor g5914 ( n2609 , n4415 , n8175 );
    or g5915 ( n2488 , n7283 , n10419 );
    and g5916 ( n2474 , n10827 , n10944 );
    and g5917 ( n6550 , n453 , n9013 );
    or g5918 ( n5549 , n4911 , n7703 );
    not g5919 ( n12049 , n12256 );
    and g5920 ( n1716 , n6354 , n10952 );
    xnor g5921 ( n12575 , n7850 , n3394 );
    not g5922 ( n9033 , n12001 );
    xnor g5923 ( n7518 , n2003 , n12762 );
    nor g5924 ( n10586 , n10701 , n7148 );
    not g5925 ( n10897 , n4657 );
    not g5926 ( n2658 , n5274 );
    not g5927 ( n2016 , n3064 );
    and g5928 ( n10394 , n3992 , n7270 );
    or g5929 ( n726 , n8452 , n8978 );
    or g5930 ( n2833 , n2050 , n4736 );
    or g5931 ( n1734 , n9370 , n6389 );
    nor g5932 ( n2423 , n10290 , n12640 );
    xnor g5933 ( n4318 , n432 , n10882 );
    or g5934 ( n4322 , n10142 , n1738 );
    and g5935 ( n12133 , n12391 , n4970 );
    not g5936 ( n12124 , n2347 );
    and g5937 ( n4099 , n3912 , n10030 );
    or g5938 ( n11142 , n7449 , n4642 );
    xnor g5939 ( n2331 , n10272 , n3390 );
    not g5940 ( n660 , n6624 );
    or g5941 ( n6574 , n12596 , n3288 );
    or g5942 ( n182 , n5809 , n826 );
    or g5943 ( n1979 , n10298 , n9596 );
    xnor g5944 ( n12658 , n6465 , n8843 );
    not g5945 ( n10534 , n6007 );
    or g5946 ( n6608 , n12454 , n1029 );
    or g5947 ( n9547 , n4498 , n6389 );
    or g5948 ( n7502 , n12853 , n9586 );
    xnor g5949 ( n12444 , n6913 , n11383 );
    xnor g5950 ( n622 , n5366 , n6476 );
    and g5951 ( n2161 , n7319 , n2521 );
    not g5952 ( n8889 , n8373 );
    and g5953 ( n529 , n2887 , n6963 );
    and g5954 ( n10588 , n7407 , n10662 );
    or g5955 ( n5690 , n11923 , n9144 );
    and g5956 ( n5602 , n8135 , n2229 );
    xnor g5957 ( n8184 , n7072 , n12449 );
    xnor g5958 ( n4656 , n6814 , n2929 );
    and g5959 ( n2594 , n9082 , n10865 );
    or g5960 ( n10180 , n191 , n7881 );
    xnor g5961 ( n1410 , n8804 , n8391 );
    nor g5962 ( n12373 , n12713 , n10027 );
    nor g5963 ( n2985 , n2550 , n2422 );
    xnor g5964 ( n11223 , n3226 , n5066 );
    xnor g5965 ( n2440 , n2569 , n9855 );
    and g5966 ( n10010 , n12262 , n8253 );
    xnor g5967 ( n9387 , n739 , n1318 );
    xnor g5968 ( n6585 , n4075 , n3385 );
    and g5969 ( n2415 , n2363 , n229 );
    and g5970 ( n5007 , n10351 , n3629 );
    nor g5971 ( n8994 , n8550 , n10934 );
    or g5972 ( n6953 , n1466 , n7055 );
    or g5973 ( n2403 , n9190 , n8079 );
    not g5974 ( n2513 , n9124 );
    xnor g5975 ( n6026 , n11037 , n1883 );
    or g5976 ( n10887 , n5945 , n1413 );
    or g5977 ( n5511 , n9297 , n10020 );
    or g5978 ( n1718 , n8428 , n3356 );
    xnor g5979 ( n10399 , n2744 , n1553 );
    xnor g5980 ( n3339 , n2412 , n7991 );
    xnor g5981 ( n6576 , n1544 , n9558 );
    not g5982 ( n6402 , n2585 );
    or g5983 ( n4893 , n9389 , n510 );
    nor g5984 ( n7638 , n7882 , n8454 );
    or g5985 ( n8267 , n636 , n7382 );
    and g5986 ( n5401 , n9732 , n3404 );
    or g5987 ( n12096 , n114 , n1413 );
    or g5988 ( n398 , n928 , n6381 );
    or g5989 ( n3169 , n11041 , n7423 );
    not g5990 ( n3713 , n10497 );
    or g5991 ( n6191 , n11415 , n12606 );
    and g5992 ( n8582 , n11425 , n6025 );
    or g5993 ( n8860 , n8582 , n772 );
    xnor g5994 ( n9571 , n767 , n9686 );
    not g5995 ( n7830 , n11055 );
    or g5996 ( n4846 , n10835 , n7921 );
    nor g5997 ( n4588 , n5681 , n10646 );
    xnor g5998 ( n4525 , n546 , n7011 );
    or g5999 ( n1315 , n5530 , n12686 );
    xnor g6000 ( n3018 , n7740 , n12724 );
    or g6001 ( n7461 , n3131 , n10813 );
    not g6002 ( n3421 , n12145 );
    and g6003 ( n3748 , n5438 , n11986 );
    and g6004 ( n9828 , n5543 , n3485 );
    and g6005 ( n6905 , n7690 , n12925 );
    xnor g6006 ( n8563 , n11784 , n5536 );
    xnor g6007 ( n12276 , n858 , n7757 );
    xnor g6008 ( n9926 , n5982 , n3923 );
    or g6009 ( n993 , n11887 , n12535 );
    or g6010 ( n12477 , n6407 , n2208 );
    not g6011 ( n3227 , n1091 );
    and g6012 ( n5004 , n4647 , n11236 );
    or g6013 ( n12027 , n7283 , n11430 );
    or g6014 ( n6899 , n5575 , n5540 );
    xnor g6015 ( n10743 , n11620 , n3100 );
    not g6016 ( n2002 , n11541 );
    nor g6017 ( n6594 , n400 , n4034 );
    or g6018 ( n5861 , n4911 , n11827 );
    and g6019 ( n8806 , n4617 , n9736 );
    nor g6020 ( n3838 , n4349 , n3580 );
    and g6021 ( n4529 , n8247 , n3868 );
    and g6022 ( n6879 , n5666 , n8134 );
    xnor g6023 ( n10300 , n1990 , n8207 );
    and g6024 ( n9526 , n10502 , n6189 );
    or g6025 ( n6967 , n2633 , n11339 );
    not g6026 ( n6615 , n5282 );
    and g6027 ( n4579 , n4561 , n10280 );
    or g6028 ( n7892 , n11127 , n9555 );
    not g6029 ( n810 , n8537 );
    or g6030 ( n3343 , n5312 , n2886 );
    and g6031 ( n3472 , n11478 , n2558 );
    xnor g6032 ( n9125 , n34 , n11214 );
    or g6033 ( n12346 , n2599 , n10681 );
    or g6034 ( n9549 , n11923 , n9521 );
    and g6035 ( n8650 , n1990 , n7635 );
    and g6036 ( n7896 , n4508 , n6184 );
    or g6037 ( n11541 , n7449 , n1476 );
    not g6038 ( n9612 , n7081 );
    xnor g6039 ( n12529 , n12582 , n3893 );
    or g6040 ( n7992 , n752 , n7558 );
    xnor g6041 ( n9708 , n9293 , n4664 );
    or g6042 ( n8139 , n8187 , n10419 );
    xnor g6043 ( n10890 , n6228 , n9525 );
    xnor g6044 ( n1680 , n11505 , n520 );
    not g6045 ( n12464 , n6709 );
    or g6046 ( n5953 , n11719 , n6389 );
    and g6047 ( n552 , n5361 , n6282 );
    not g6048 ( n2026 , n3834 );
    xnor g6049 ( n10589 , n6997 , n5692 );
    or g6050 ( n3939 , n2700 , n3268 );
    nor g6051 ( n4768 , n2504 , n3814 );
    xnor g6052 ( n7272 , n6914 , n4447 );
    or g6053 ( n1250 , n2147 , n10329 );
    and g6054 ( n2150 , n8505 , n11731 );
    xnor g6055 ( n5586 , n11181 , n9803 );
    or g6056 ( n11110 , n4644 , n11624 );
    xnor g6057 ( n12320 , n11851 , n9255 );
    not g6058 ( n1989 , n9358 );
    not g6059 ( n10267 , n3953 );
    or g6060 ( n11334 , n2197 , n11855 );
    or g6061 ( n4907 , n989 , n8859 );
    xnor g6062 ( n9173 , n7812 , n559 );
    or g6063 ( n7137 , n2456 , n8644 );
    xnor g6064 ( n12249 , n7753 , n11771 );
    or g6065 ( n4531 , n5441 , n1862 );
    and g6066 ( n7762 , n8462 , n736 );
    and g6067 ( n7924 , n1811 , n829 );
    and g6068 ( n2184 , n9744 , n3963 );
    xnor g6069 ( n7068 , n1310 , n7818 );
    xnor g6070 ( n3200 , n3056 , n3367 );
    or g6071 ( n4392 , n11958 , n2589 );
    not g6072 ( n973 , n10228 );
    xnor g6073 ( n1590 , n7700 , n9132 );
    and g6074 ( n10051 , n6687 , n2509 );
    and g6075 ( n1271 , n2605 , n11921 );
    or g6076 ( n5926 , n807 , n5540 );
    nor g6077 ( n2391 , n387 , n11859 );
    or g6078 ( n2175 , n11317 , n1265 );
    not g6079 ( n1546 , n3842 );
    xnor g6080 ( n5719 , n10973 , n4399 );
    nor g6081 ( n2399 , n11711 , n4833 );
    nor g6082 ( n5148 , n1392 , n2337 );
    and g6083 ( n656 , n9246 , n3017 );
    xnor g6084 ( n8493 , n7643 , n8232 );
    nor g6085 ( n5875 , n12551 , n8647 );
    or g6086 ( n252 , n8187 , n1162 );
    xnor g6087 ( n11149 , n5075 , n9434 );
    not g6088 ( n8062 , n10640 );
    or g6089 ( n9332 , n2494 , n10775 );
    or g6090 ( n3594 , n11782 , n5114 );
    nor g6091 ( n5382 , n12375 , n7444 );
    or g6092 ( n6650 , n7116 , n5540 );
    xnor g6093 ( n7563 , n3027 , n8459 );
    xnor g6094 ( n12917 , n10502 , n6189 );
    xnor g6095 ( n10809 , n10260 , n9975 );
    not g6096 ( n2872 , n10174 );
    xnor g6097 ( n8638 , n11744 , n499 );
    xnor g6098 ( n10784 , n3126 , n188 );
    xnor g6099 ( n12553 , n3679 , n4494 );
    or g6100 ( n10274 , n1259 , n3778 );
    or g6101 ( n7832 , n41 , n1255 );
    and g6102 ( n5288 , n12617 , n1648 );
    not g6103 ( n895 , n4422 );
    and g6104 ( n11104 , n688 , n7853 );
    or g6105 ( n2340 , n5530 , n8957 );
    or g6106 ( n12889 , n2919 , n6319 );
    or g6107 ( n1808 , n10750 , n4818 );
    not g6108 ( n11719 , n11257 );
    xnor g6109 ( n4601 , n8352 , n9879 );
    xnor g6110 ( n9565 , n3585 , n3554 );
    xnor g6111 ( n1062 , n11295 , n6155 );
    not g6112 ( n3917 , n6621 );
    and g6113 ( n4200 , n164 , n10881 );
    or g6114 ( n9304 , n8552 , n6513 );
    not g6115 ( n9056 , n12031 );
    xnor g6116 ( n9981 , n2828 , n12623 );
    or g6117 ( n11507 , n10750 , n8644 );
    and g6118 ( n1895 , n1827 , n11479 );
    xnor g6119 ( n9152 , n1892 , n481 );
    or g6120 ( n4302 , n1384 , n9194 );
    nor g6121 ( n12136 , n6322 , n8035 );
    and g6122 ( n12915 , n10928 , n6703 );
    nor g6123 ( n5584 , n4767 , n4987 );
    nor g6124 ( n11661 , n8329 , n11063 );
    or g6125 ( n10768 , n994 , n7389 );
    xnor g6126 ( n3806 , n9163 , n402 );
    or g6127 ( n7208 , n3561 , n8312 );
    xnor g6128 ( n9439 , n12084 , n6502 );
    and g6129 ( n5925 , n12330 , n3980 );
    or g6130 ( n3916 , n4796 , n9493 );
    xnor g6131 ( n565 , n10842 , n2123 );
    and g6132 ( n5036 , n12033 , n6781 );
    not g6133 ( n1092 , n3988 );
    or g6134 ( n11535 , n1271 , n12528 );
    and g6135 ( n6209 , n4173 , n7858 );
    and g6136 ( n7664 , n12512 , n7414 );
    and g6137 ( n8792 , n6252 , n7089 );
    or g6138 ( n4582 , n8313 , n879 );
    not g6139 ( n11277 , n5526 );
    nor g6140 ( n7056 , n10776 , n5683 );
    and g6141 ( n9754 , n4121 , n11975 );
    and g6142 ( n11007 , n5783 , n12915 );
    xnor g6143 ( n3398 , n11332 , n2772 );
    xnor g6144 ( n742 , n8927 , n9071 );
    and g6145 ( n12454 , n4777 , n7475 );
    or g6146 ( n1616 , n12503 , n1509 );
    or g6147 ( n3964 , n5355 , n7389 );
    or g6148 ( n10292 , n12503 , n9144 );
    nor g6149 ( n6279 , n4207 , n3371 );
    xnor g6150 ( n6950 , n10379 , n964 );
    xnor g6151 ( n1339 , n6807 , n10465 );
    not g6152 ( n6968 , n6430 );
    and g6153 ( n1683 , n5739 , n10241 );
    or g6154 ( n4831 , n4510 , n6410 );
    nor g6155 ( n12036 , n7766 , n12898 );
    or g6156 ( n1809 , n12237 , n8655 );
    or g6157 ( n1702 , n10750 , n6513 );
    or g6158 ( n8502 , n7718 , n5884 );
    or g6159 ( n8422 , n332 , n3703 );
    and g6160 ( n822 , n5362 , n7725 );
    and g6161 ( n9091 , n11602 , n7707 );
    nor g6162 ( n3191 , n1755 , n6913 );
    not g6163 ( n4720 , n9332 );
    and g6164 ( n5101 , n10797 , n7954 );
    or g6165 ( n8516 , n1141 , n1192 );
    nor g6166 ( n9495 , n7317 , n11492 );
    xnor g6167 ( n2303 , n11885 , n9804 );
    and g6168 ( n8389 , n11150 , n6726 );
    not g6169 ( n2356 , n6786 );
    or g6170 ( n5392 , n8882 , n12435 );
    xnor g6171 ( n280 , n1335 , n10027 );
    and g6172 ( n2392 , n149 , n368 );
    not g6173 ( n6309 , n7458 );
    xnor g6174 ( n3817 , n3247 , n5028 );
    xnor g6175 ( n2091 , n5904 , n1379 );
    not g6176 ( n2964 , n5798 );
    xnor g6177 ( n12714 , n2312 , n3899 );
    or g6178 ( n10672 , n3638 , n7528 );
    xnor g6179 ( n2534 , n11468 , n7789 );
    not g6180 ( n4364 , n8544 );
    xnor g6181 ( n8147 , n12277 , n1769 );
    xnor g6182 ( n5610 , n7405 , n11066 );
    and g6183 ( n6249 , n6881 , n6489 );
    and g6184 ( n9051 , n12561 , n1586 );
    and g6185 ( n9728 , n1471 , n9763 );
    or g6186 ( n4522 , n3734 , n12508 );
    nor g6187 ( n12890 , n4292 , n3690 );
    not g6188 ( n763 , n5128 );
    xnor g6189 ( n194 , n5281 , n8777 );
    or g6190 ( n4780 , n1937 , n2232 );
    nor g6191 ( n6637 , n8719 , n2637 );
    not g6192 ( n3352 , n9341 );
    and g6193 ( n9252 , n708 , n2032 );
    xnor g6194 ( n4241 , n11561 , n4067 );
    and g6195 ( n595 , n9248 , n6592 );
    or g6196 ( n10018 , n2456 , n12686 );
    or g6197 ( n7317 , n8026 , n7395 );
    and g6198 ( n10951 , n5554 , n11625 );
    xnor g6199 ( n3259 , n5828 , n5186 );
    and g6200 ( n11502 , n9943 , n9035 );
    xnor g6201 ( n6282 , n10604 , n7356 );
    and g6202 ( n3831 , n8276 , n11728 );
    xnor g6203 ( n9930 , n1392 , n1992 );
    xnor g6204 ( n2193 , n5345 , n2614 );
    xnor g6205 ( n6264 , n5922 , n9614 );
    not g6206 ( n7343 , n11155 );
    or g6207 ( n2335 , n9370 , n4775 );
    or g6208 ( n8458 , n9370 , n7341 );
    nor g6209 ( n6825 , n9861 , n6047 );
    and g6210 ( n2968 , n1963 , n11769 );
    and g6211 ( n8041 , n1003 , n6517 );
    and g6212 ( n5529 , n4302 , n4927 );
    not g6213 ( n1133 , n9197 );
    not g6214 ( n5396 , n3208 );
    or g6215 ( n2001 , n1170 , n6748 );
    not g6216 ( n1870 , n6745 );
    not g6217 ( n8745 , n10022 );
    xnor g6218 ( n741 , n9190 , n7901 );
    xnor g6219 ( n4752 , n7350 , n454 );
    or g6220 ( n4328 , n8405 , n12535 );
    nor g6221 ( n8263 , n9676 , n1451 );
    and g6222 ( n4685 , n7641 , n9910 );
    xnor g6223 ( n10865 , n9651 , n12543 );
    or g6224 ( n8508 , n5486 , n3557 );
    or g6225 ( n6328 , n962 , n2020 );
    and g6226 ( n8461 , n12284 , n663 );
    or g6227 ( n6020 , n3211 , n8653 );
    or g6228 ( n4290 , n1051 , n6455 );
    or g6229 ( n12847 , n4363 , n6321 );
    or g6230 ( n10080 , n6977 , n7558 );
    and g6231 ( n10250 , n1123 , n396 );
    xnor g6232 ( n7085 , n11905 , n6715 );
    not g6233 ( n7759 , n9102 );
    not g6234 ( n3922 , n4462 );
    xnor g6235 ( n9718 , n11306 , n5381 );
    xnor g6236 ( n6467 , n8350 , n4455 );
    xnor g6237 ( n8032 , n6754 , n6573 );
    or g6238 ( n10281 , n10912 , n6143 );
    not g6239 ( n11914 , n11679 );
    xnor g6240 ( n226 , n5350 , n5175 );
    or g6241 ( n5119 , n4256 , n4467 );
    and g6242 ( n2563 , n2108 , n5590 );
    and g6243 ( n6651 , n2285 , n2525 );
    and g6244 ( n12670 , n1445 , n5727 );
    and g6245 ( n6363 , n4356 , n6210 );
    and g6246 ( n9064 , n2413 , n10802 );
    not g6247 ( n10311 , n4436 );
    xnor g6248 ( n747 , n7772 , n5421 );
    and g6249 ( n10133 , n11266 , n8286 );
    xnor g6250 ( n9945 , n12951 , n12840 );
    xnor g6251 ( n9035 , n10413 , n12254 );
    and g6252 ( n11459 , n7690 , n1564 );
    or g6253 ( n1282 , n6696 , n1938 );
    xnor g6254 ( n9042 , n9328 , n11826 );
    or g6255 ( n11057 , n1903 , n3332 );
    or g6256 ( n12839 , n2893 , n1014 );
    not g6257 ( n4677 , n1500 );
    or g6258 ( n6788 , n6373 , n7506 );
    or g6259 ( n1330 , n10349 , n7328 );
    xnor g6260 ( n721 , n11099 , n3288 );
    nor g6261 ( n11622 , n12088 , n3490 );
    or g6262 ( n6946 , n2456 , n530 );
    nor g6263 ( n2151 , n4365 , n4323 );
    xnor g6264 ( n9606 , n6816 , n7132 );
    or g6265 ( n4355 , n5445 , n9215 );
    xnor g6266 ( n7597 , n9250 , n12117 );
    not g6267 ( n201 , n6239 );
    or g6268 ( n444 , n9122 , n4460 );
    xnor g6269 ( n8654 , n7306 , n10584 );
    or g6270 ( n10791 , n8810 , n318 );
    and g6271 ( n8688 , n5101 , n9206 );
    or g6272 ( n1978 , n7686 , n6074 );
    and g6273 ( n10825 , n7100 , n9714 );
    or g6274 ( n2606 , n7083 , n672 );
    or g6275 ( n1375 , n2285 , n2525 );
    or g6276 ( n3236 , n752 , n3903 );
    or g6277 ( n10609 , n724 , n8022 );
    xnor g6278 ( n8788 , n983 , n4109 );
    or g6279 ( n12365 , n3746 , n3903 );
    and g6280 ( n8907 , n2613 , n3826 );
    or g6281 ( n2123 , n8870 , n8740 );
    and g6282 ( n6693 , n9364 , n1458 );
    or g6283 ( n1473 , n9170 , n4242 );
    and g6284 ( n3604 , n7862 , n3932 );
    not g6285 ( n10007 , n7616 );
    not g6286 ( n2504 , n11754 );
    not g6287 ( n5666 , n11184 );
    or g6288 ( n1354 , n5765 , n9078 );
    xnor g6289 ( n6367 , n7019 , n9666 );
    xor g6290 ( n791 , n3618 , n11585 );
    or g6291 ( n988 , n11531 , n10295 );
    or g6292 ( n10905 , n9021 , n4170 );
    or g6293 ( n7587 , n7283 , n1915 );
    not g6294 ( n4391 , n6905 );
    and g6295 ( n1733 , n4426 , n1225 );
    xnor g6296 ( n12515 , n9179 , n4217 );
    or g6297 ( n6339 , n4059 , n10066 );
    not g6298 ( n8607 , n8634 );
    or g6299 ( n12243 , n10169 , n1411 );
    or g6300 ( n2018 , n7306 , n10584 );
    nor g6301 ( n2248 , n161 , n550 );
    or g6302 ( n12892 , n1814 , n739 );
    xnor g6303 ( n7547 , n6551 , n8243 );
    xnor g6304 ( n5553 , n7569 , n12207 );
    xnor g6305 ( n2554 , n8262 , n11093 );
    xnor g6306 ( n704 , n9201 , n5911 );
    not g6307 ( n1345 , n3166 );
    or g6308 ( n4592 , n1539 , n4400 );
    xnor g6309 ( n1522 , n10417 , n3660 );
    xnor g6310 ( n6936 , n5181 , n3410 );
    nor g6311 ( n3097 , n8983 , n4172 );
    and g6312 ( n1584 , n2650 , n9728 );
    xnor g6313 ( n10427 , n4384 , n6587 );
    and g6314 ( n974 , n7221 , n6453 );
    or g6315 ( n3913 , n1183 , n5468 );
    and g6316 ( n2934 , n1936 , n6723 );
    not g6317 ( n5858 , n10547 );
    xnor g6318 ( n12360 , n3460 , n12229 );
    nor g6319 ( n3380 , n5533 , n7726 );
    not g6320 ( n799 , n10964 );
    or g6321 ( n7651 , n7391 , n12328 );
    or g6322 ( n1172 , n7992 , n8569 );
    and g6323 ( n6151 , n5994 , n8722 );
    or g6324 ( n8322 , n10309 , n11180 );
    or g6325 ( n11015 , n11674 , n2726 );
    or g6326 ( n1529 , n4071 , n5612 );
    or g6327 ( n537 , n1937 , n11122 );
    and g6328 ( n9631 , n7564 , n1363 );
    or g6329 ( n7006 , n5596 , n6829 );
    or g6330 ( n10829 , n9791 , n10393 );
    or g6331 ( n5380 , n8026 , n6169 );
    xnor g6332 ( n5692 , n4806 , n6236 );
    and g6333 ( n8800 , n8020 , n1644 );
    and g6334 ( n12200 , n5507 , n5045 );
    xnor g6335 ( n10099 , n12423 , n7303 );
    xnor g6336 ( n8960 , n12597 , n5313 );
    or g6337 ( n8869 , n1941 , n6169 );
    not g6338 ( n629 , n11913 );
    xnor g6339 ( n10884 , n6830 , n9316 );
    xnor g6340 ( n3222 , n12353 , n2350 );
    or g6341 ( n11177 , n6718 , n2020 );
    xnor g6342 ( n10362 , n6989 , n4836 );
    and g6343 ( n8515 , n7678 , n1526 );
    xnor g6344 ( n12415 , n12466 , n8960 );
    or g6345 ( n1832 , n5120 , n174 );
    not g6346 ( n12328 , n9195 );
    or g6347 ( n5637 , n3453 , n2809 );
    and g6348 ( n3995 , n998 , n4129 );
    or g6349 ( n11330 , n5031 , n6798 );
    nor g6350 ( n11682 , n3058 , n5901 );
    nor g6351 ( n11615 , n4061 , n10437 );
    or g6352 ( n8816 , n1937 , n11896 );
    or g6353 ( n3699 , n4131 , n10190 );
    nor g6354 ( n6452 , n605 , n9288 );
    not g6355 ( n9490 , n9544 );
    xnor g6356 ( n2051 , n8839 , n5774 );
    or g6357 ( n3318 , n855 , n10699 );
    not g6358 ( n12503 , n5319 );
    xnor g6359 ( n5444 , n8315 , n2789 );
    nor g6360 ( n7118 , n6244 , n8180 );
    and g6361 ( n1777 , n5013 , n3588 );
    not g6362 ( n8787 , n10116 );
    not g6363 ( n9618 , n3762 );
    xnor g6364 ( n729 , n11409 , n9032 );
    xnor g6365 ( n1681 , n7458 , n11748 );
    or g6366 ( n7181 , n1249 , n7963 );
    xnor g6367 ( n547 , n2684 , n5103 );
    or g6368 ( n3695 , n4798 , n4368 );
    and g6369 ( n2572 , n4286 , n8472 );
    not g6370 ( n7379 , n8225 );
    xnor g6371 ( n7576 , n8184 , n10655 );
    nor g6372 ( n9296 , n5338 , n8933 );
    or g6373 ( n10119 , n4911 , n2358 );
    not g6374 ( n12899 , n10391 );
    xnor g6375 ( n1294 , n6392 , n4090 );
    xnor g6376 ( n10601 , n6946 , n9104 );
    and g6377 ( n2550 , n12819 , n3379 );
    nor g6378 ( n7098 , n5097 , n9773 );
    nor g6379 ( n7291 , n2148 , n5275 );
    xnor g6380 ( n9501 , n9365 , n3307 );
    and g6381 ( n2900 , n7802 , n7141 );
    or g6382 ( n3756 , n10502 , n6189 );
    xnor g6383 ( n11938 , n11545 , n5067 );
    xnor g6384 ( n4067 , n8072 , n11527 );
    xnor g6385 ( n8400 , n7271 , n11263 );
    xor g6386 ( n1020 , n2177 , n1150 );
    or g6387 ( n9226 , n7116 , n2232 );
    xnor g6388 ( n2222 , n7286 , n7443 );
    not g6389 ( n8718 , n2408 );
    and g6390 ( n448 , n11543 , n3378 );
    not g6391 ( n2052 , n1105 );
    and g6392 ( n11322 , n8118 , n9965 );
    xnor g6393 ( n8351 , n7071 , n8338 );
    xnor g6394 ( n162 , n8835 , n8793 );
    xnor g6395 ( n4590 , n2448 , n12070 );
    xnor g6396 ( n3077 , n11828 , n5133 );
    not g6397 ( n9161 , n9416 );
    and g6398 ( n7575 , n7133 , n2395 );
    not g6399 ( n5991 , n7826 );
    and g6400 ( n11756 , n6352 , n1533 );
    and g6401 ( n7177 , n5767 , n5760 );
    xnor g6402 ( n10285 , n8714 , n10468 );
    not g6403 ( n12453 , n458 );
    not g6404 ( n9185 , n10604 );
    xnor g6405 ( n8723 , n6933 , n3994 );
    not g6406 ( n12772 , n8323 );
    xnor g6407 ( n6112 , n2180 , n927 );
    nor g6408 ( n6971 , n6121 , n5946 );
    not g6409 ( n3862 , n9099 );
    xnor g6410 ( n2094 , n10922 , n11650 );
    and g6411 ( n3376 , n580 , n2469 );
    or g6412 ( n8116 , n8583 , n1476 );
    nor g6413 ( n6393 , n4892 , n583 );
    not g6414 ( n6433 , n535 );
    nor g6415 ( n7819 , n11875 , n1408 );
    or g6416 ( n6561 , n8870 , n9188 );
    or g6417 ( n4246 , n4628 , n12883 );
    or g6418 ( n11528 , n4561 , n10280 );
    xnor g6419 ( n2960 , n2909 , n6280 );
    or g6420 ( n6948 , n2630 , n5324 );
    xnor g6421 ( n9337 , n2405 , n10090 );
    and g6422 ( n719 , n7862 , n4921 );
    xnor g6423 ( n11062 , n5166 , n4285 );
    and g6424 ( n9489 , n2653 , n12359 );
    or g6425 ( n872 , n5915 , n8648 );
    and g6426 ( n10689 , n2293 , n10956 );
    or g6427 ( n706 , n12594 , n5469 );
    nor g6428 ( n2142 , n8473 , n2442 );
    and g6429 ( n8823 , n7578 , n3644 );
    not g6430 ( n9344 , n2047 );
    xnor g6431 ( n456 , n3262 , n4072 );
    not g6432 ( n5307 , n9443 );
    xnor g6433 ( n528 , n4379 , n11693 );
    or g6434 ( n4426 , n7100 , n9714 );
    or g6435 ( n3480 , n2830 , n4405 );
    and g6436 ( n6709 , n9920 , n5212 );
    or g6437 ( n4415 , n11026 , n9160 );
    nor g6438 ( n7192 , n5695 , n6745 );
    nor g6439 ( n11059 , n10996 , n8292 );
    xnor g6440 ( n3910 , n12630 , n5074 );
    and g6441 ( n6670 , n4393 , n4829 );
    and g6442 ( n3825 , n1581 , n437 );
    or g6443 ( n349 , n1699 , n12080 );
    not g6444 ( n3943 , n7831 );
    xnor g6445 ( n7362 , n4019 , n2027 );
    xnor g6446 ( n12949 , n10034 , n5413 );
    or g6447 ( n430 , n2456 , n10854 );
    and g6448 ( n1424 , n1714 , n2592 );
    or g6449 ( n7099 , n3746 , n3356 );
    xnor g6450 ( n8271 , n8166 , n3253 );
    xnor g6451 ( n5980 , n2416 , n9088 );
    or g6452 ( n7078 , n6577 , n7876 );
    or g6453 ( n6044 , n7487 , n7752 );
    and g6454 ( n7043 , n5860 , n9111 );
    xnor g6455 ( n2624 , n651 , n10687 );
    not g6456 ( n4280 , n10178 );
    or g6457 ( n11532 , n1941 , n12816 );
    nor g6458 ( n3596 , n10228 , n11971 );
    or g6459 ( n6677 , n10057 , n5822 );
    or g6460 ( n2963 , n5765 , n12771 );
    and g6461 ( n8773 , n12243 , n11331 );
    xnor g6462 ( n11523 , n3000 , n6639 );
    not g6463 ( n5876 , n7377 );
    not g6464 ( n1781 , n4522 );
    xnor g6465 ( n94 , n10686 , n8935 );
    xnor g6466 ( n369 , n6066 , n8814 );
    xnor g6467 ( n7585 , n4107 , n11695 );
    or g6468 ( n10305 , n2670 , n10220 );
    xnor g6469 ( n7985 , n2216 , n2810 );
    and g6470 ( n10073 , n3433 , n1722 );
    and g6471 ( n508 , n7862 , n11407 );
    xnor g6472 ( n7359 , n10210 , n8366 );
    or g6473 ( n4047 , n10926 , n11396 );
    xnor g6474 ( n12123 , n12379 , n1429 );
    xnor g6475 ( n9676 , n494 , n2070 );
    or g6476 ( n12775 , n4059 , n7424 );
    xnor g6477 ( n475 , n9413 , n9022 );
    xnor g6478 ( n9546 , n11788 , n3641 );
    or g6479 ( n8004 , n744 , n11432 );
    or g6480 ( n2890 , n12503 , n9521 );
    and g6481 ( n7658 , n648 , n6769 );
    or g6482 ( n5102 , n10530 , n1038 );
    xnor g6483 ( n2104 , n10461 , n12523 );
    and g6484 ( n7554 , n2575 , n175 );
    not g6485 ( n423 , n7023 );
    and g6486 ( n9781 , n3954 , n8955 );
    xnor g6487 ( n4930 , n4893 , n5085 );
    and g6488 ( n6787 , n3961 , n9219 );
    or g6489 ( n2995 , n8129 , n12603 );
    xnor g6490 ( n8202 , n3296 , n5557 );
    nor g6491 ( n2794 , n3297 , n12424 );
    not g6492 ( n6288 , n1190 );
    nor g6493 ( n12556 , n2702 , n449 );
    xnor g6494 ( n8362 , n3128 , n12381 );
    xnor g6495 ( n1637 , n10023 , n11085 );
    nor g6496 ( n3545 , n8142 , n6308 );
    not g6497 ( n2578 , n9216 );
    xnor g6498 ( n11983 , n3991 , n12154 );
    xnor g6499 ( n7036 , n4904 , n5493 );
    or g6500 ( n1591 , n10262 , n5630 );
    xnor g6501 ( n12287 , n6544 , n6435 );
    or g6502 ( n1370 , n7839 , n1413 );
    xnor g6503 ( n3559 , n4114 , n7336 );
    and g6504 ( n10348 , n905 , n11505 );
    and g6505 ( n1316 , n2619 , n4978 );
    or g6506 ( n1073 , n8789 , n1733 );
    not g6507 ( n2977 , n9683 );
    not g6508 ( n2582 , n8763 );
    or g6509 ( n10370 , n2911 , n4530 );
    xnor g6510 ( n4809 , n11534 , n9184 );
    or g6511 ( n10385 , n8814 , n6278 );
    nor g6512 ( n3847 , n7157 , n6746 );
    xnor g6513 ( n5112 , n5578 , n780 );
    and g6514 ( n8284 , n6386 , n3841 );
    xnor g6515 ( n1015 , n4566 , n10370 );
    xnor g6516 ( n5175 , n382 , n1060 );
    xnor g6517 ( n8163 , n8239 , n11857 );
    xnor g6518 ( n12572 , n6650 , n305 );
    xnor g6519 ( n2583 , n10269 , n5295 );
    or g6520 ( n7441 , n1051 , n7952 );
    nor g6521 ( n3994 , n10092 , n1666 );
    or g6522 ( n3796 , n12552 , n6989 );
    or g6523 ( n6635 , n8187 , n7341 );
    nor g6524 ( n1299 , n3244 , n6024 );
    or g6525 ( n3409 , n5450 , n6694 );
    xnor g6526 ( n3720 , n10761 , n3234 );
    xnor g6527 ( n12505 , n9572 , n6711 );
    xnor g6528 ( n7824 , n4259 , n10003 );
    not g6529 ( n5434 , n8347 );
    xnor g6530 ( n10459 , n6570 , n8478 );
    xnor g6531 ( n3554 , n7441 , n3009 );
    and g6532 ( n1350 , n9677 , n12869 );
    xnor g6533 ( n9238 , n4788 , n2787 );
    or g6534 ( n10529 , n4059 , n6402 );
    and g6535 ( n4684 , n9299 , n11158 );
    and g6536 ( n7850 , n6002 , n9590 );
    xnor g6537 ( n1948 , n816 , n7530 );
    xnor g6538 ( n579 , n2856 , n3165 );
    or g6539 ( n6894 , n11552 , n1047 );
    xnor g6540 ( n9967 , n3895 , n1729 );
    xnor g6541 ( n6641 , n6488 , n5731 );
    and g6542 ( n5469 , n2249 , n1676 );
    nor g6543 ( n8897 , n12399 , n4889 );
    and g6544 ( n8312 , n12098 , n5499 );
    not g6545 ( n11497 , n4089 );
    nor g6546 ( n34 , n64 , n5143 );
    xnor g6547 ( n11185 , n10575 , n3187 );
    and g6548 ( n8613 , n11616 , n3023 );
    or g6549 ( n2400 , n5355 , n12328 );
    xnor g6550 ( n5451 , n4562 , n12689 );
    xnor g6551 ( n8468 , n4237 , n12852 );
    xnor g6552 ( n7721 , n3858 , n9738 );
    not g6553 ( n6323 , n525 );
    or g6554 ( n4265 , n5915 , n8644 );
    or g6555 ( n9816 , n8206 , n3195 );
    and g6556 ( n5067 , n2816 , n9378 );
    or g6557 ( n5321 , n254 , n7775 );
    or g6558 ( n5484 , n180 , n285 );
    xnor g6559 ( n655 , n6045 , n6432 );
    not g6560 ( n4593 , n2485 );
    and g6561 ( n7736 , n8835 , n9595 );
    and g6562 ( n6898 , n2308 , n11133 );
    xnor g6563 ( n176 , n4620 , n9912 );
    xnor g6564 ( n9594 , n1712 , n11632 );
    not g6565 ( n1667 , n8319 );
    or g6566 ( n12578 , n7111 , n11131 );
    xnor g6567 ( n8836 , n11395 , n4735 );
    or g6568 ( n11690 , n1051 , n7558 );
    xnor g6569 ( n9407 , n8692 , n2421 );
    xnor g6570 ( n1255 , n5808 , n7573 );
    xnor g6571 ( n11342 , n6018 , n5892 );
    xnor g6572 ( n9900 , n2492 , n12099 );
    not g6573 ( n2844 , n10013 );
    xnor g6574 ( n7403 , n2332 , n6034 );
    not g6575 ( n7050 , n2602 );
    not g6576 ( n8539 , n1420 );
    not g6577 ( n7703 , n2508 );
    xnor g6578 ( n4245 , n10838 , n3060 );
    xnor g6579 ( n5670 , n5649 , n3004 );
    nor g6580 ( n6819 , n2073 , n12028 );
    or g6581 ( n4881 , n8705 , n12336 );
    and g6582 ( n1300 , n398 , n2322 );
    and g6583 ( n10344 , n1442 , n3668 );
    or g6584 ( n12514 , n12840 , n12951 );
    nor g6585 ( n1764 , n6612 , n4896 );
    xnor g6586 ( n4477 , n2943 , n11097 );
    or g6587 ( n1014 , n7283 , n12843 );
    or g6588 ( n2591 , n5786 , n9464 );
    xnor g6589 ( n6337 , n4438 , n12498 );
    xnor g6590 ( n3837 , n7507 , n7658 );
    not g6591 ( n7938 , n11526 );
    and g6592 ( n5186 , n10739 , n3938 );
    xnor g6593 ( n3551 , n10249 , n12082 );
    xnor g6594 ( n1419 , n3565 , n1894 );
    or g6595 ( n12379 , n9696 , n6394 );
    and g6596 ( n1516 , n9953 , n6396 );
    and g6597 ( n3060 , n7964 , n9329 );
    or g6598 ( n2573 , n6251 , n3403 );
    xnor g6599 ( n11766 , n2531 , n9945 );
    and g6600 ( n1314 , n2511 , n926 );
    xnor g6601 ( n9943 , n11541 , n4936 );
    or g6602 ( n2503 , n12503 , n1047 );
    not g6603 ( n7949 , n2467 );
    xnor g6604 ( n9460 , n5 , n3720 );
    and g6605 ( n6768 , n7965 , n11876 );
    and g6606 ( n3804 , n2437 , n2085 );
    xnor g6607 ( n11809 , n6424 , n1332 );
    xnor g6608 ( n7867 , n11408 , n12450 );
    xnor g6609 ( n2605 , n7956 , n11251 );
    not g6610 ( n4645 , n8843 );
    and g6611 ( n1638 , n8267 , n11939 );
    or g6612 ( n9714 , n8428 , n5540 );
    xnor g6613 ( n9983 , n7659 , n117 );
    or g6614 ( n1928 , n2267 , n1096 );
    or g6615 ( n10381 , n2456 , n2964 );
    and g6616 ( n2470 , n5305 , n3932 );
    nor g6617 ( n570 , n10071 , n1604 );
    not g6618 ( n12724 , n3728 );
    or g6619 ( n3253 , n8026 , n12899 );
    xnor g6620 ( n3054 , n11715 , n12575 );
    nor g6621 ( n10552 , n4739 , n1846 );
    xnor g6622 ( n59 , n5598 , n11672 );
    and g6623 ( n11034 , n7914 , n4351 );
    nor g6624 ( n4408 , n12513 , n12690 );
    nor g6625 ( n10948 , n9250 , n10453 );
    xnor g6626 ( n2831 , n6381 , n4404 );
    and g6627 ( n4401 , n6660 , n5406 );
    or g6628 ( n10347 , n6977 , n11820 );
    or g6629 ( n10172 , n8552 , n7928 );
    or g6630 ( n646 , n3743 , n6138 );
    and g6631 ( n7060 , n12155 , n6473 );
    or g6632 ( n11196 , n10500 , n974 );
    nor g6633 ( n2265 , n1006 , n9217 );
    xnor g6634 ( n3639 , n8029 , n9423 );
    and g6635 ( n9052 , n3604 , n4421 );
    nor g6636 ( n3503 , n5936 , n2998 );
    or g6637 ( n3311 , n4092 , n5907 );
    not g6638 ( n10780 , n12623 );
    xnor g6639 ( n3771 , n1776 , n9452 );
    or g6640 ( n12281 , n2099 , n10311 );
    xnor g6641 ( n5467 , n9860 , n9100 );
    and g6642 ( n1594 , n2393 , n11791 );
    or g6643 ( n11993 , n6303 , n8084 );
    or g6644 ( n2638 , n11380 , n11115 );
    xnor g6645 ( n7493 , n4171 , n10077 );
    and g6646 ( n7720 , n5961 , n2804 );
    or g6647 ( n9428 , n191 , n7246 );
    xnor g6648 ( n7929 , n1240 , n10183 );
    not g6649 ( n11137 , n11777 );
    xnor g6650 ( n8417 , n8824 , n7272 );
    xnor g6651 ( n3783 , n4718 , n11260 );
    not g6652 ( n6925 , n3633 );
    xnor g6653 ( n3883 , n12291 , n923 );
    and g6654 ( n8355 , n10222 , n3828 );
    or g6655 ( n6003 , n1937 , n3903 );
    nor g6656 ( n9987 , n2618 , n1654 );
    xnor g6657 ( n2757 , n10057 , n5399 );
    not g6658 ( n156 , n9010 );
    xnor g6659 ( n12250 , n7595 , n4709 );
    or g6660 ( n2308 , n2548 , n8435 );
    and g6661 ( n3003 , n186 , n3435 );
    xnor g6662 ( n12381 , n2852 , n1789 );
    xnor g6663 ( n4106 , n11684 , n10731 );
    xnor g6664 ( n2581 , n3945 , n7259 );
    xnor g6665 ( n4708 , n12841 , n6563 );
    not g6666 ( n7800 , n8779 );
    or g6667 ( n10261 , n4185 , n4965 );
    or g6668 ( n5237 , n10079 , n10538 );
    nor g6669 ( n743 , n4211 , n6259 );
    not g6670 ( n7732 , n7814 );
    or g6671 ( n9905 , n10835 , n9568 );
    or g6672 ( n9918 , n4628 , n4913 );
    xnor g6673 ( n3001 , n5872 , n9018 );
    not g6674 ( n10275 , n4034 );
    or g6675 ( n1337 , n1223 , n2892 );
    xnor g6676 ( n2311 , n4899 , n4329 );
    not g6677 ( n2499 , n613 );
    xnor g6678 ( n3035 , n6771 , n9662 );
    or g6679 ( n3114 , n10605 , n3388 );
    xnor g6680 ( n8721 , n70 , n11210 );
    or g6681 ( n10726 , n5809 , n12686 );
    or g6682 ( n5813 , n8822 , n4472 );
    and g6683 ( n2634 , n12708 , n9745 );
    or g6684 ( n12767 , n196 , n11477 );
    xnor g6685 ( n6246 , n12074 , n1540 );
    nor g6686 ( n11087 , n9810 , n11696 );
    xnor g6687 ( n5604 , n11281 , n4629 );
    nor g6688 ( n12066 , n8919 , n1582 );
    xnor g6689 ( n828 , n7400 , n10089 );
    or g6690 ( n7557 , n114 , n11775 );
    xnor g6691 ( n11946 , n3420 , n594 );
    and g6692 ( n10187 , n10088 , n3295 );
    not g6693 ( n3249 , n6884 );
    xnor g6694 ( n7484 , n4630 , n7722 );
    and g6695 ( n11735 , n2042 , n10305 );
    or g6696 ( n96 , n4502 , n9610 );
    or g6697 ( n1627 , n2424 , n12846 );
    or g6698 ( n11452 , n10355 , n5863 );
    xnor g6699 ( n11130 , n8017 , n3364 );
    xnor g6700 ( n2666 , n5756 , n11913 );
    not g6701 ( n9548 , n11934 );
    or g6702 ( n10448 , n10879 , n3911 );
    not g6703 ( n12797 , n7523 );
    xnor g6704 ( n7263 , n6812 , n12018 );
    not g6705 ( n3624 , n933 );
    and g6706 ( n11758 , n8961 , n3193 );
    and g6707 ( n10499 , n2262 , n2066 );
    xnor g6708 ( n6892 , n11289 , n11024 );
    or g6709 ( n2042 , n2536 , n12112 );
    nor g6710 ( n8503 , n7393 , n12362 );
    not g6711 ( n9650 , n1 );
    and g6712 ( n1913 , n5859 , n11824 );
    xnor g6713 ( n8130 , n12409 , n11258 );
    or g6714 ( n5969 , n9878 , n1932 );
    xnor g6715 ( n733 , n5167 , n11781 );
    xnor g6716 ( n768 , n5852 , n4095 );
    xnor g6717 ( n9992 , n683 , n12953 );
    nor g6718 ( n3892 , n5594 , n11095 );
    or g6719 ( n4501 , n1699 , n10422 );
    not g6720 ( n5725 , n11141 );
    xnor g6721 ( n8196 , n3115 , n4853 );
    or g6722 ( n7204 , n114 , n2232 );
    not g6723 ( n299 , n3874 );
    or g6724 ( n11078 , n10194 , n9928 );
    nor g6725 ( n2576 , n1995 , n464 );
    not g6726 ( n4084 , n6174 );
    xnor g6727 ( n12548 , n6272 , n2126 );
    and g6728 ( n12347 , n1122 , n12427 );
    not g6729 ( n10304 , n2924 );
    xnor g6730 ( n7589 , n2871 , n6415 );
    or g6731 ( n10002 , n962 , n3606 );
    or g6732 ( n11668 , n5394 , n5152 );
    nor g6733 ( n5225 , n3420 , n7634 );
    and g6734 ( n669 , n6462 , n7742 );
    not g6735 ( n5871 , n3479 );
    or g6736 ( n12829 , n430 , n10085 );
    and g6737 ( n2671 , n6256 , n7489 );
    not g6738 ( n2730 , n10061 );
    not g6739 ( n311 , n399 );
    nor g6740 ( n6962 , n7594 , n4902 );
    not g6741 ( n12801 , n3087 );
    xnor g6742 ( n10971 , n4697 , n6430 );
    and g6743 ( n10296 , n11449 , n1365 );
    and g6744 ( n5095 , n1809 , n882 );
    or g6745 ( n165 , n10142 , n3911 );
    or g6746 ( n11594 , n12662 , n10491 );
    not g6747 ( n7212 , n5758 );
    or g6748 ( n2354 , n9787 , n7619 );
    or g6749 ( n2068 , n1561 , n12817 );
    xnor g6750 ( n1671 , n8227 , n10209 );
    xnor g6751 ( n38 , n12426 , n12085 );
    not g6752 ( n8114 , n2307 );
    or g6753 ( n7094 , n3413 , n4877 );
    xnor g6754 ( n11157 , n10541 , n8852 );
    not g6755 ( n5961 , n12746 );
    xnor g6756 ( n10431 , n9570 , n12050 );
    and g6757 ( n1418 , n7593 , n3377 );
    and g6758 ( n10719 , n9929 , n4842 );
    xnor g6759 ( n3985 , n6727 , n9439 );
    not g6760 ( n5788 , n7667 );
    xnor g6761 ( n853 , n6773 , n9419 );
    xnor g6762 ( n9984 , n2947 , n6033 );
    xnor g6763 ( n122 , n6825 , n6100 );
    xnor g6764 ( n10800 , n4637 , n4454 );
    and g6765 ( n1404 , n7749 , n8602 );
    not g6766 ( n8622 , n7820 );
    nor g6767 ( n5437 , n10433 , n4485 );
    and g6768 ( n3178 , n8678 , n10154 );
    not g6769 ( n12602 , n11942 );
    and g6770 ( n12476 , n4698 , n3815 );
    or g6771 ( n12784 , n1319 , n3417 );
    xnor g6772 ( n7459 , n6788 , n4495 );
    nor g6773 ( n9477 , n6896 , n9856 );
    or g6774 ( n374 , n1111 , n11177 );
    or g6775 ( n12723 , n9373 , n10916 );
    and g6776 ( n10437 , n3116 , n9931 );
    and g6777 ( n6832 , n5816 , n6522 );
    xnor g6778 ( n7722 , n1415 , n4431 );
    not g6779 ( n9521 , n8433 );
    xnor g6780 ( n110 , n7792 , n12048 );
    xnor g6781 ( n2152 , n8329 , n6434 );
    xnor g6782 ( n5775 , n8896 , n4710 );
    and g6783 ( n7611 , n4380 , n5245 );
    xnor g6784 ( n4669 , n9898 , n1513 );
    xnor g6785 ( n2425 , n85 , n2884 );
    nor g6786 ( n6567 , n3784 , n3317 );
    and g6787 ( n7339 , n6909 , n845 );
    nor g6788 ( n6022 , n11752 , n11781 );
    nor g6789 ( n3562 , n5396 , n6757 );
    xnor g6790 ( n8968 , n356 , n3398 );
    or g6791 ( n4389 , n989 , n1738 );
    or g6792 ( n7900 , n3820 , n10916 );
    or g6793 ( n8268 , n114 , n6455 );
    or g6794 ( n8368 , n7112 , n7795 );
    not g6795 ( n9350 , n6947 );
    not g6796 ( n9741 , n6429 );
    and g6797 ( n9591 , n6317 , n12929 );
    or g6798 ( n5306 , n4059 , n12843 );
    and g6799 ( n5612 , n11801 , n10413 );
    or g6800 ( n6329 , n8598 , n5581 );
    or g6801 ( n1226 , n11867 , n6075 );
    xnor g6802 ( n6120 , n2541 , n10427 );
    or g6803 ( n7864 , n4628 , n5326 );
    not g6804 ( n11165 , n8973 );
    and g6805 ( n10795 , n5250 , n2214 );
    xnor g6806 ( n3854 , n8765 , n29 );
    not g6807 ( n3958 , n5041 );
    xnor g6808 ( n1045 , n2700 , n566 );
    or g6809 ( n7109 , n11652 , n5939 );
    or g6810 ( n8401 , n8687 , n1509 );
    not g6811 ( n5787 , n528 );
    and g6812 ( n1236 , n6294 , n1067 );
    xnor g6813 ( n9832 , n5576 , n4353 );
    not g6814 ( n510 , n11662 );
    not g6815 ( n10755 , n2233 );
    or g6816 ( n11603 , n2123 , n11101 );
    nor g6817 ( n1742 , n9753 , n12671 );
    xnor g6818 ( n1237 , n12584 , n436 );
    not g6819 ( n3242 , n11936 );
    xnor g6820 ( n6838 , n8475 , n12600 );
    xnor g6821 ( n5298 , n9341 , n1765 );
    xnor g6822 ( n5544 , n1334 , n5566 );
    or g6823 ( n9995 , n1183 , n12080 );
    or g6824 ( n3800 , n9530 , n7879 );
    not g6825 ( n3591 , n11875 );
    or g6826 ( n2191 , n4984 , n9153 );
    nor g6827 ( n11770 , n3729 , n10250 );
    or g6828 ( n3084 , n1092 , n3175 );
    not g6829 ( n7649 , n3089 );
    or g6830 ( n2155 , n5355 , n7881 );
    or g6831 ( n9222 , n10196 , n795 );
    or g6832 ( n12156 , n4059 , n11430 );
    xnor g6833 ( n3770 , n5174 , n6068 );
    nor g6834 ( n1381 , n12536 , n883 );
    or g6835 ( n3174 , n8262 , n3085 );
    or g6836 ( n5432 , n5575 , n6455 );
    or g6837 ( n3518 , n4325 , n628 );
    and g6838 ( n4314 , n137 , n11922 );
    xnor g6839 ( n12226 , n3863 , n3293 );
    and g6840 ( n7517 , n5087 , n5357 );
    xnor g6841 ( n6528 , n6662 , n8311 );
    or g6842 ( n8153 , n10844 , n5699 );
    xnor g6843 ( n10271 , n6834 , n2996 );
    xnor g6844 ( n9556 , n10605 , n1964 );
    and g6845 ( n2476 , n10545 , n2498 );
    xnor g6846 ( n915 , n3221 , n7846 );
    not g6847 ( n5372 , n6361 );
    xnor g6848 ( n7758 , n7909 , n4432 );
    xnor g6849 ( n11861 , n10666 , n10431 );
    and g6850 ( n6640 , n3699 , n2733 );
    and g6851 ( n2271 , n9131 , n12463 );
    nor g6852 ( n2286 , n12235 , n12154 );
    xnor g6853 ( n6873 , n4057 , n908 );
    and g6854 ( n10059 , n3053 , n7943 );
    or g6855 ( n6590 , n994 , n1851 );
    nor g6856 ( n11436 , n952 , n9828 );
    not g6857 ( n9818 , n6440 );
    xnor g6858 ( n12471 , n4602 , n6980 );
    xnor g6859 ( n11650 , n78 , n1934 );
    not g6860 ( n5766 , n173 );
    not g6861 ( n12883 , n12044 );
    and g6862 ( n7004 , n11417 , n1314 );
    nor g6863 ( n3341 , n11523 , n7973 );
    and g6864 ( n10701 , n8113 , n8626 );
    not g6865 ( n9877 , n10253 );
    and g6866 ( n10870 , n800 , n2468 );
    or g6867 ( n7286 , n8738 , n4527 );
    xnor g6868 ( n462 , n9453 , n9646 );
    nor g6869 ( n9267 , n5958 , n4765 );
    or g6870 ( n4597 , n5271 , n2006 );
    or g6871 ( n1180 , n11552 , n5258 );
    xnor g6872 ( n8712 , n3093 , n6690 );
    not g6873 ( n7861 , n10378 );
    xnor g6874 ( n12074 , n8751 , n523 );
    not g6875 ( n7973 , n572 );
    xnor g6876 ( n9224 , n7084 , n9091 );
    not g6877 ( n5474 , n3931 );
    or g6878 ( n12530 , n3743 , n8285 );
    or g6879 ( n4638 , n4546 , n7545 );
    xnor g6880 ( n4691 , n3088 , n853 );
    or g6881 ( n6890 , n9878 , n4818 );
    not g6882 ( n12388 , n12099 );
    and g6883 ( n5839 , n573 , n11044 );
    and g6884 ( n2751 , n10744 , n2240 );
    xnor g6885 ( n6415 , n4993 , n6099 );
    and g6886 ( n6864 , n9432 , n7226 );
    or g6887 ( n7105 , n7709 , n795 );
    xnor g6888 ( n12736 , n6145 , n12101 );
    not g6889 ( n8259 , n12826 );
    or g6890 ( n4393 , n351 , n10275 );
    nor g6891 ( n3161 , n7019 , n3782 );
    or g6892 ( n3150 , n1051 , n6169 );
    and g6893 ( n4514 , n4858 , n2243 );
    xnor g6894 ( n3246 , n7652 , n4830 );
    xnor g6895 ( n2457 , n9935 , n9488 );
    xnor g6896 ( n9101 , n8911 , n2734 );
    xnor g6897 ( n4473 , n9900 , n5063 );
    or g6898 ( n12135 , n1768 , n206 );
    xnor g6899 ( n5324 , n5572 , n12908 );
    xnor g6900 ( n4063 , n6210 , n6112 );
    xnor g6901 ( n5074 , n8758 , n12027 );
    xnor g6902 ( n1793 , n3236 , n1057 );
    or g6903 ( n10255 , n6336 , n4077 );
    xnor g6904 ( n8009 , n7078 , n838 );
    and g6905 ( n3904 , n5314 , n217 );
    nor g6906 ( n5143 , n6260 , n2770 );
    and g6907 ( n6831 , n8981 , n4379 );
    not g6908 ( n3768 , n5368 );
    or g6909 ( n279 , n5026 , n9139 );
    nor g6910 ( n9693 , n12555 , n9947 );
    or g6911 ( n2197 , n6977 , n12816 );
    and g6912 ( n7997 , n8855 , n10760 );
    xnor g6913 ( n6101 , n5980 , n3532 );
    xnor g6914 ( n4300 , n9734 , n2857 );
    nor g6915 ( n10204 , n8633 , n5713 );
    nor g6916 ( n219 , n12832 , n4271 );
    or g6917 ( n12414 , n274 , n11815 );
    and g6918 ( n9464 , n2155 , n11112 );
    or g6919 ( n9376 , n8850 , n10805 );
    nor g6920 ( n7937 , n8492 , n6188 );
    xnor g6921 ( n3972 , n8682 , n6736 );
    not g6922 ( n807 , n7320 );
    not g6923 ( n7170 , n7526 );
    or g6924 ( n607 , n5859 , n11824 );
    xnor g6925 ( n6688 , n354 , n12793 );
    and g6926 ( n11329 , n5204 , n283 );
    or g6927 ( n7825 , n5036 , n2991 );
    and g6928 ( n3244 , n12012 , n11889 );
    nor g6929 ( n2856 , n8101 , n10885 );
    xnor g6930 ( n11416 , n866 , n1580 );
    or g6931 ( n2502 , n12361 , n7395 );
    and g6932 ( n10787 , n1867 , n7371 );
    or g6933 ( n9349 , n4465 , n12916 );
    and g6934 ( n8868 , n11074 , n3652 );
    and g6935 ( n12904 , n3256 , n1081 );
    and g6936 ( n1901 , n3210 , n10527 );
    xnor g6937 ( n9473 , n10927 , n2051 );
    or g6938 ( n5710 , n10117 , n5140 );
    and g6939 ( n10748 , n3816 , n5228 );
    not g6940 ( n10469 , n190 );
    not g6941 ( n8217 , n2699 );
    xnor g6942 ( n6085 , n1009 , n1639 );
    and g6943 ( n215 , n8941 , n1418 );
    xnor g6944 ( n12820 , n8308 , n5607 );
    or g6945 ( n273 , n7480 , n1080 );
    nor g6946 ( n9977 , n4914 , n4364 );
    not g6947 ( n4449 , n1229 );
    and g6948 ( n11677 , n6185 , n5017 );
    nor g6949 ( n1537 , n1809 , n882 );
    or g6950 ( n5780 , n5355 , n2358 );
    not g6951 ( n740 , n11802 );
    or g6952 ( n5573 , n5247 , n9020 );
    or g6953 ( n10922 , n636 , n9188 );
    or g6954 ( n9685 , n6579 , n3093 );
    and g6955 ( n1446 , n3698 , n2394 );
    xnor g6956 ( n12581 , n11867 , n6475 );
    or g6957 ( n7847 , n11678 , n5805 );
    or g6958 ( n288 , n11923 , n1047 );
    xnor g6959 ( n4751 , n1296 , n12948 );
    not g6960 ( n6257 , n7869 );
    or g6961 ( n12380 , n10435 , n4895 );
    not g6962 ( n4223 , n11955 );
    xnor g6963 ( n12937 , n2880 , n792 );
    and g6964 ( n3348 , n6666 , n8991 );
    and g6965 ( n2039 , n5959 , n8534 );
    and g6966 ( n7631 , n11577 , n8053 );
    xnor g6967 ( n4621 , n2275 , n4543 );
    and g6968 ( n1508 , n6191 , n8895 );
    nor g6969 ( n6211 , n7396 , n5885 );
    xnor g6970 ( n185 , n6204 , n11735 );
    xnor g6971 ( n2126 , n1465 , n848 );
    not g6972 ( n11077 , n150 );
    xnor g6973 ( n1890 , n755 , n3080 );
    xnor g6974 ( n8820 , n8087 , n10371 );
    or g6975 ( n11538 , n752 , n7425 );
    xnor g6976 ( n1961 , n6454 , n177 );
    not g6977 ( n3383 , n7459 );
    nor g6978 ( n6662 , n3359 , n10047 );
    not g6979 ( n12361 , n12299 );
    xnor g6980 ( n6676 , n11305 , n10501 );
    nor g6981 ( n9217 , n3462 , n7240 );
    or g6982 ( n5299 , n825 , n10284 );
    and g6983 ( n5580 , n11221 , n3260 );
    xnor g6984 ( n384 , n10252 , n8932 );
    not g6985 ( n748 , n9265 );
    xnor g6986 ( n12291 , n2204 , n751 );
    not g6987 ( n9953 , n6068 );
    nor g6988 ( n1763 , n1645 , n11000 );
    xnor g6989 ( n262 , n3723 , n712 );
    or g6990 ( n6673 , n5915 , n10422 );
    nor g6991 ( n1965 , n929 , n11453 );
    or g6992 ( n5040 , n945 , n4521 );
    xnor g6993 ( n2566 , n804 , n1716 );
    or g6994 ( n1230 , n835 , n7979 );
    or g6995 ( n4957 , n8181 , n8485 );
    or g6996 ( n7396 , n1941 , n7952 );
    xnor g6997 ( n33 , n12365 , n11406 );
    not g6998 ( n6577 , n2464 );
    xnor g6999 ( n2975 , n5762 , n6217 );
    nor g7000 ( n5716 , n11138 , n10218 );
    or g7001 ( n864 , n3996 , n1046 );
    or g7002 ( n708 , n8367 , n388 );
    and g7003 ( n12286 , n9843 , n1066 );
    xnor g7004 ( n868 , n9345 , n3167 );
    and g7005 ( n1217 , n2384 , n3852 );
    and g7006 ( n3612 , n3682 , n8958 );
    xnor g7007 ( n5322 , n6010 , n2117 );
    nor g7008 ( n12368 , n9785 , n574 );
    xnor g7009 ( n3109 , n9187 , n12113 );
    or g7010 ( n8594 , n3743 , n5759 );
    and g7011 ( n12071 , n4773 , n403 );
    and g7012 ( n3083 , n938 , n3311 );
    nor g7013 ( n238 , n4799 , n7147 );
    or g7014 ( n11154 , n11878 , n10215 );
    nor g7015 ( n12901 , n5848 , n3913 );
    nor g7016 ( n12656 , n4119 , n378 );
    xnor g7017 ( n5635 , n3667 , n3090 );
    and g7018 ( n7826 , n6877 , n7354 );
    nor g7019 ( n8770 , n12271 , n12707 );
    or g7020 ( n5077 , n3791 , n11806 );
    or g7021 ( n3386 , n5530 , n12446 );
    or g7022 ( n2580 , n10682 , n4011 );
    and g7023 ( n6383 , n7441 , n3009 );
    and g7024 ( n5745 , n10239 , n9325 );
    and g7025 ( n11189 , n6877 , n9640 );
    not g7026 ( n10879 , n3627 );
    xnor g7027 ( n10268 , n6554 , n5201 );
    not g7028 ( n6274 , n11439 );
    or g7029 ( n949 , n638 , n7227 );
    or g7030 ( n2724 , n10955 , n6744 );
    and g7031 ( n1838 , n4683 , n2732 );
    nor g7032 ( n11205 , n9123 , n3969 );
    xnor g7033 ( n7628 , n12520 , n12664 );
    nor g7034 ( n10019 , n144 , n7137 );
    not g7035 ( n8244 , n2398 );
    or g7036 ( n12298 , n7116 , n5538 );
    and g7037 ( n3235 , n1297 , n1391 );
    xnor g7038 ( n5873 , n5553 , n2765 );
    or g7039 ( n12679 , n3076 , n10868 );
    not g7040 ( n8149 , n874 );
    xnor g7041 ( n394 , n8235 , n10175 );
    not g7042 ( n11958 , n8336 );
    or g7043 ( n2562 , n3015 , n2294 );
    and g7044 ( n3133 , n12093 , n10939 );
    xnor g7045 ( n1969 , n10874 , n1300 );
    xnor g7046 ( n12672 , n6270 , n11978 );
    not g7047 ( n5264 , n12133 );
    not g7048 ( n11520 , n11983 );
    or g7049 ( n1272 , n4562 , n12689 );
    xnor g7050 ( n5241 , n353 , n10828 );
    or g7051 ( n775 , n752 , n12357 );
    or g7052 ( n5071 , n3533 , n5660 );
    xnor g7053 ( n8566 , n6399 , n1740 );
    xnor g7054 ( n1610 , n12129 , n5165 );
    and g7055 ( n11049 , n10340 , n1460 );
    xnor g7056 ( n3005 , n11081 , n3086 );
    or g7057 ( n6077 , n7850 , n3566 );
    nor g7058 ( n6259 , n4357 , n3103 );
    and g7059 ( n8124 , n12940 , n4297 );
    or g7060 ( n4506 , n8583 , n2020 );
    and g7061 ( n2742 , n5964 , n6038 );
    xnor g7062 ( n7667 , n4501 , n6334 );
    or g7063 ( n7806 , n10142 , n130 );
    or g7064 ( n907 , n4528 , n6187 );
    or g7065 ( n3718 , n989 , n11746 );
    or g7066 ( n866 , n2456 , n10422 );
    or g7067 ( n6163 , n9262 , n9521 );
    or g7068 ( n3255 , n2099 , n8109 );
    xnor g7069 ( n4031 , n7316 , n9090 );
    xnor g7070 ( n6403 , n10601 , n1802 );
    and g7071 ( n10833 , n5828 , n5186 );
    xnor g7072 ( n5879 , n1688 , n8703 );
    xnor g7073 ( n5852 , n6663 , n8456 );
    xnor g7074 ( n2918 , n672 , n11454 );
    and g7075 ( n4185 , n4582 , n3955 );
    xnor g7076 ( n3633 , n9139 , n2200 );
    or g7077 ( n10186 , n6293 , n11194 );
    xor g7078 ( n4922 , n8831 , n6406 );
    or g7079 ( n6365 , n8959 , n3903 );
    xnor g7080 ( n5015 , n11027 , n3611 );
    xnor g7081 ( n12085 , n58 , n6146 );
    and g7082 ( n8798 , n1375 , n3527 );
    and g7083 ( n10892 , n6283 , n3543 );
    or g7084 ( n8559 , n6554 , n5201 );
    and g7085 ( n9514 , n8951 , n11022 );
    not g7086 ( n10732 , n8960 );
    not g7087 ( n2169 , n5635 );
    and g7088 ( n6921 , n1583 , n7077 );
    and g7089 ( n4351 , n4101 , n9349 );
    not g7090 ( n10207 , n6326 );
    or g7091 ( n12256 , n1078 , n5983 );
    and g7092 ( n9852 , n2696 , n10412 );
    xnor g7093 ( n3637 , n1044 , n5602 );
    nor g7094 ( n5022 , n8826 , n631 );
    not g7095 ( n9170 , n9920 );
    and g7096 ( n11241 , n4038 , n8589 );
    or g7097 ( n5436 , n9000 , n5391 );
    xnor g7098 ( n9979 , n10218 , n11393 );
    and g7099 ( n12520 , n1185 , n7755 );
    xnor g7100 ( n9065 , n3452 , n1370 );
    xnor g7101 ( n7031 , n4195 , n12121 );
    not g7102 ( n8309 , n12904 );
    xnor g7103 ( n2381 , n6777 , n2908 );
    and g7104 ( n4504 , n4511 , n8863 );
    nor g7105 ( n7522 , n3593 , n12291 );
    not g7106 ( n8552 , n12648 );
    xnor g7107 ( n7340 , n6337 , n9447 );
    not g7108 ( n6425 , n12539 );
    or g7109 ( n11940 , n5915 , n8740 );
    nor g7110 ( n5644 , n1415 , n4630 );
    and g7111 ( n8099 , n10725 , n5111 );
    not g7112 ( n2066 , n10959 );
    or g7113 ( n7617 , n11744 , n2222 );
    xnor g7114 ( n3293 , n3625 , n9031 );
    or g7115 ( n10781 , n7405 , n1148 );
    and g7116 ( n12956 , n7427 , n11868 );
    and g7117 ( n6884 , n2515 , n12925 );
    or g7118 ( n6050 , n10157 , n7506 );
    or g7119 ( n12348 , n12119 , n9188 );
    not g7120 ( n6523 , n5001 );
    not g7121 ( n7555 , n8083 );
    and g7122 ( n9005 , n2213 , n1443 );
    xnor g7123 ( n5284 , n9973 , n7180 );
    not g7124 ( n5695 , n4023 );
    xnor g7125 ( n9894 , n6661 , n4493 );
    and g7126 ( n7267 , n4770 , n560 );
    or g7127 ( n8822 , n2456 , n8109 );
    or g7128 ( n253 , n10142 , n1455 );
    or g7129 ( n9837 , n8187 , n1455 );
    xnor g7130 ( n7833 , n10975 , n2152 );
    nor g7131 ( n4485 , n3469 , n12326 );
    or g7132 ( n2592 , n10283 , n4947 );
    or g7133 ( n3875 , n11552 , n2020 );
    nor g7134 ( n4672 , n12625 , n9963 );
    xnor g7135 ( n2109 , n1218 , n4600 );
    and g7136 ( n5901 , n8967 , n1673 );
    and g7137 ( n2295 , n10216 , n2238 );
    or g7138 ( n2797 , n4 , n3283 );
    xnor g7139 ( n1523 , n2262 , n3564 );
    xnor g7140 ( n1050 , n1706 , n313 );
    or g7141 ( n10671 , n2228 , n5286 );
    not g7142 ( n12941 , n4619 );
    and g7143 ( n3401 , n5767 , n10848 );
    and g7144 ( n3000 , n11732 , n5506 );
    not g7145 ( n7854 , n2488 );
    xnor g7146 ( n6822 , n7030 , n10271 );
    or g7147 ( n5758 , n11958 , n5012 );
    and g7148 ( n2081 , n5416 , n7347 );
    and g7149 ( n3248 , n11462 , n11148 );
    or g7150 ( n9798 , n3820 , n4527 );
    nor g7151 ( n5222 , n7082 , n10579 );
    xnor g7152 ( n5405 , n9549 , n4318 );
    and g7153 ( n8671 , n5240 , n3932 );
    xnor g7154 ( n8936 , n2731 , n5702 );
    and g7155 ( n5157 , n4785 , n6869 );
    xnor g7156 ( n8398 , n7997 , n3092 );
    not g7157 ( n4758 , n564 );
    or g7158 ( n12738 , n9388 , n10302 );
    or g7159 ( n11229 , n12569 , n9067 );
    and g7160 ( n610 , n4983 , n9636 );
    and g7161 ( n12953 , n1747 , n8610 );
    xnor g7162 ( n8315 , n6961 , n9019 );
    not g7163 ( n9202 , n9036 );
    nor g7164 ( n12802 , n9527 , n8050 );
    and g7165 ( n8005 , n10587 , n10140 );
    xnor g7166 ( n12865 , n236 , n3770 );
    and g7167 ( n11003 , n4415 , n325 );
    nor g7168 ( n9696 , n5474 , n11287 );
    xnor g7169 ( n6727 , n2372 , n1032 );
    xnor g7170 ( n12697 , n288 , n11386 );
    not g7171 ( n3292 , n9277 );
    xnor g7172 ( n8150 , n5518 , n9327 );
    xnor g7173 ( n7221 , n904 , n7464 );
    or g7174 ( n7572 , n7449 , n5759 );
    or g7175 ( n5818 , n8907 , n10483 );
    and g7176 ( n4960 , n6353 , n3601 );
    not g7177 ( n9346 , n5140 );
    and g7178 ( n4307 , n7891 , n521 );
    or g7179 ( n7064 , n686 , n7876 );
    or g7180 ( n8682 , n2832 , n4400 );
    or g7181 ( n4012 , n8870 , n3224 );
    or g7182 ( n3305 , n12853 , n8648 );
    and g7183 ( n8701 , n5025 , n56 );
    xnor g7184 ( n5869 , n2525 , n7174 );
    not g7185 ( n9160 , n10898 );
    or g7186 ( n477 , n12797 , n6455 );
    or g7187 ( n3710 , n8738 , n9521 );
    or g7188 ( n835 , n5355 , n4242 );
    nor g7189 ( n8662 , n9564 , n706 );
    or g7190 ( n12815 , n925 , n1958 );
    or g7191 ( n9017 , n4628 , n8644 );
    not g7192 ( n1384 , n4349 );
    nor g7193 ( n10836 , n2048 , n8939 );
    and g7194 ( n10408 , n4222 , n11724 );
    xnor g7195 ( n9774 , n2820 , n9672 );
    or g7196 ( n6411 , n3251 , n1274 );
    or g7197 ( n11125 , n12635 , n4988 );
    and g7198 ( n111 , n10849 , n6284 );
    and g7199 ( n1833 , n5181 , n3410 );
    not g7200 ( n5945 , n9241 );
    or g7201 ( n12455 , n11923 , n5258 );
    nor g7202 ( n900 , n7796 , n4348 );
    xnor g7203 ( n3047 , n4162 , n10406 );
    xnor g7204 ( n11448 , n2201 , n12725 );
    or g7205 ( n6381 , n636 , n826 );
    not g7206 ( n8678 , n5955 );
    xnor g7207 ( n6269 , n2055 , n9941 );
    or g7208 ( n3977 , n2921 , n5604 );
    and g7209 ( n8521 , n3797 , n10816 );
    xnor g7210 ( n11664 , n6835 , n11469 );
    xnor g7211 ( n5201 , n1671 , n5862 );
    or g7212 ( n10662 , n4628 , n8109 );
    nor g7213 ( n2773 , n6211 , n2576 );
    or g7214 ( n7407 , n2099 , n7382 );
    xnor g7215 ( n3935 , n9967 , n1893 );
    or g7216 ( n5524 , n1937 , n2815 );
    and g7217 ( n848 , n4046 , n12171 );
    not g7218 ( n3820 , n5198 );
    not g7219 ( n1498 , n993 );
    nor g7220 ( n2192 , n10555 , n7791 );
    or g7221 ( n9892 , n11552 , n10916 );
    and g7222 ( n7537 , n4015 , n4740 );
    or g7223 ( n6407 , n5575 , n3903 );
    not g7224 ( n2450 , n6772 );
    xnor g7225 ( n6202 , n4892 , n4591 );
    or g7226 ( n6542 , n5793 , n798 );
    not g7227 ( n2756 , n2885 );
    nor g7228 ( n814 , n6496 , n8190 );
    xnor g7229 ( n1888 , n7082 , n7845 );
    and g7230 ( n8442 , n2300 , n4130 );
    xnor g7231 ( n10048 , n11569 , n7880 );
    or g7232 ( n4366 , n10750 , n12735 );
    xnor g7233 ( n9675 , n3934 , n8888 );
    not g7234 ( n3566 , n3394 );
    and g7235 ( n1896 , n4536 , n4220 );
    xnor g7236 ( n8780 , n4451 , n1852 );
    xnor g7237 ( n5805 , n5889 , n7103 );
    or g7238 ( n6368 , n1699 , n7382 );
    xnor g7239 ( n6840 , n7207 , n12674 );
    or g7240 ( n12296 , n11026 , n9078 );
    or g7241 ( n6231 , n752 , n5538 );
    not g7242 ( n1699 , n5283 );
    or g7243 ( n9529 , n3743 , n8643 );
    or g7244 ( n5866 , n1982 , n7621 );
    and g7245 ( n202 , n2382 , n948 );
    xnor g7246 ( n3745 , n6705 , n5909 );
    not g7247 ( n3603 , n5544 );
    or g7248 ( n11988 , n10879 , n7881 );
    xnor g7249 ( n3331 , n7462 , n2105 );
    or g7250 ( n2817 , n4498 , n10066 );
    or g7251 ( n1089 , n1024 , n7498 );
    not g7252 ( n3836 , n2565 );
    or g7253 ( n4622 , n12361 , n5012 );
    xnor g7254 ( n7429 , n5453 , n5550 );
    or g7255 ( n9245 , n2872 , n7876 );
    xnor g7256 ( n1193 , n515 , n5941 );
    xnor g7257 ( n429 , n6629 , n8667 );
    and g7258 ( n2030 , n7961 , n10969 );
    or g7259 ( n10761 , n10835 , n5502 );
    xnor g7260 ( n11066 , n8937 , n534 );
    xnor g7261 ( n9733 , n422 , n12482 );
    xnor g7262 ( n11844 , n2760 , n1555 );
    xnor g7263 ( n4406 , n12122 , n11191 );
    nor g7264 ( n5933 , n4501 , n8630 );
    or g7265 ( n1569 , n10108 , n1455 );
    xnor g7266 ( n12004 , n5633 , n9424 );
    not g7267 ( n7829 , n4409 );
    nor g7268 ( n9063 , n621 , n6844 );
    not g7269 ( n3675 , n6251 );
    not g7270 ( n1836 , n10783 );
    xnor g7271 ( n1356 , n12838 , n3450 );
    xnor g7272 ( n10844 , n7309 , n9083 );
    nor g7273 ( n5349 , n90 , n12732 );
    not g7274 ( n2232 , n11728 );
    or g7275 ( n1007 , n989 , n7246 );
    and g7276 ( n8573 , n1944 , n782 );
    or g7277 ( n1279 , n4849 , n1935 );
    nor g7278 ( n300 , n12487 , n1857 );
    or g7279 ( n8732 , n7449 , n795 );
    xnor g7280 ( n11885 , n8848 , n5651 );
    xnor g7281 ( n53 , n7227 , n10494 );
    xnor g7282 ( n1023 , n1034 , n5722 );
    and g7283 ( n4578 , n6241 , n9948 );
    or g7284 ( n6461 , n5765 , n8643 );
    nor g7285 ( n8997 , n5415 , n389 );
    or g7286 ( n5039 , n10679 , n6409 );
    or g7287 ( n7126 , n5575 , n5311 );
    xnor g7288 ( n1328 , n5822 , n2757 );
    not g7289 ( n12741 , n9246 );
    not g7290 ( n11901 , n6521 );
    not g7291 ( n10663 , n6889 );
    or g7292 ( n681 , n2215 , n6729 );
    nor g7293 ( n7034 , n12960 , n10487 );
    and g7294 ( n6563 , n127 , n12679 );
    xnor g7295 ( n1570 , n10720 , n8088 );
    nor g7296 ( n10690 , n7032 , n10895 );
    or g7297 ( n2956 , n9607 , n4429 );
    xnor g7298 ( n227 , n8205 , n6820 );
    xnor g7299 ( n1035 , n5397 , n6346 );
    and g7300 ( n3479 , n4441 , n4854 );
    xnor g7301 ( n12533 , n12701 , n5309 );
    xnor g7302 ( n470 , n6975 , n11853 );
    xnor g7303 ( n8088 , n5643 , n9173 );
    or g7304 ( n1556 , n2367 , n9521 );
    or g7305 ( n11616 , n10983 , n2817 );
    not g7306 ( n8421 , n2831 );
    or g7307 ( n474 , n10835 , n3451 );
    xnor g7308 ( n10444 , n41 , n383 );
    or g7309 ( n2156 , n10518 , n2916 );
    xnor g7310 ( n874 , n2571 , n11342 );
    not g7311 ( n7765 , n10096 );
    or g7312 ( n2010 , n9943 , n9035 );
    xnor g7313 ( n9771 , n8612 , n2335 );
    nor g7314 ( n3407 , n4619 , n2719 );
    or g7315 ( n3918 , n7937 , n11145 );
    nor g7316 ( n6804 , n8003 , n11638 );
    xnor g7317 ( n7648 , n3645 , n3493 );
    not g7318 ( n6926 , n508 );
    or g7319 ( n6571 , n5915 , n4913 );
    or g7320 ( n1352 , n752 , n2754 );
    not g7321 ( n10816 , n6467 );
    xnor g7322 ( n12193 , n7045 , n10937 );
    not g7323 ( n8492 , n12910 );
    and g7324 ( n3952 , n4514 , n9659 );
    xnor g7325 ( n7455 , n1665 , n5196 );
    or g7326 ( n522 , n8738 , n1047 );
    nor g7327 ( n7087 , n6801 , n6011 );
    xor g7328 ( n11079 , n760 , n12835 );
    and g7329 ( n1155 , n6053 , n5830 );
    or g7330 ( n1899 , n9170 , n3911 );
    xnor g7331 ( n7207 , n7288 , n4845 );
    and g7332 ( n9055 , n7527 , n9772 );
    or g7333 ( n10744 , n5575 , n11122 );
    not g7334 ( n11866 , n11022 );
    nor g7335 ( n1903 , n5544 , n10443 );
    or g7336 ( n4298 , n2832 , n11827 );
    and g7337 ( n1982 , n11984 , n6460 );
    or g7338 ( n4167 , n3127 , n7881 );
    nor g7339 ( n1086 , n8776 , n11526 );
    xnor g7340 ( n9447 , n12270 , n11676 );
    xnor g7341 ( n12139 , n7549 , n8096 );
    not g7342 ( n10906 , n9414 );
    and g7343 ( n3574 , n7629 , n2112 );
    not g7344 ( n2832 , n4516 );
    nor g7345 ( n7381 , n9028 , n3945 );
    nor g7346 ( n9860 , n3276 , n10787 );
    and g7347 ( n6025 , n10818 , n9949 );
    and g7348 ( n541 , n4131 , n10190 );
    and g7349 ( n4878 , n683 , n12834 );
    and g7350 ( n2883 , n2834 , n10526 );
    not g7351 ( n8855 , n11557 );
    and g7352 ( n46 , n10776 , n5683 );
    not g7353 ( n5837 , n6855 );
    and g7354 ( n9186 , n12878 , n10906 );
    not g7355 ( n1280 , n8241 );
    and g7356 ( n5114 , n2168 , n2354 );
    or g7357 ( n9281 , n379 , n5193 );
    xnor g7358 ( n1132 , n2659 , n6419 );
    and g7359 ( n6136 , n124 , n11883 );
    or g7360 ( n7899 , n7449 , n9144 );
    xnor g7361 ( n10597 , n37 , n11920 );
    and g7362 ( n7578 , n11055 , n12958 );
    nor g7363 ( n6874 , n10488 , n6039 );
    or g7364 ( n12633 , n7283 , n11746 );
    xnor g7365 ( n2635 , n1866 , n10603 );
    and g7366 ( n6566 , n12957 , n71 );
    or g7367 ( n5107 , n12237 , n3924 );
    xnor g7368 ( n10603 , n9271 , n4185 );
    not g7369 ( n8154 , n1765 );
    not g7370 ( n9959 , n8455 );
    nor g7371 ( n2216 , n8288 , n3999 );
    xnor g7372 ( n4410 , n420 , n10308 );
    not g7373 ( n11970 , n8122 );
    or g7374 ( n11969 , n9887 , n9226 );
    or g7375 ( n1656 , n5902 , n1455 );
    not g7376 ( n8345 , n1232 );
    xnor g7377 ( n3270 , n5720 , n6565 );
    and g7378 ( n8359 , n7690 , n12489 );
    or g7379 ( n4022 , n5491 , n7743 );
    or g7380 ( n5855 , n1072 , n2975 );
    or g7381 ( n7608 , n3743 , n1739 );
    not g7382 ( n9364 , n2345 );
    or g7383 ( n1649 , n1231 , n10446 );
    or g7384 ( n7316 , n1051 , n3903 );
    or g7385 ( n4358 , n191 , n8524 );
    and g7386 ( n7427 , n2470 , n1994 );
    nor g7387 ( n9596 , n2653 , n12359 );
    nor g7388 ( n12891 , n7894 , n1693 );
    nor g7389 ( n3586 , n8829 , n8979 );
    not g7390 ( n7881 , n11877 );
    xnor g7391 ( n4268 , n10929 , n6328 );
    or g7392 ( n118 , n8481 , n1048 );
    not g7393 ( n2598 , n12644 );
    or g7394 ( n2170 , n10846 , n5525 );
    xnor g7395 ( n7942 , n10405 , n11004 );
    not g7396 ( n2877 , n11523 );
    or g7397 ( n8912 , n994 , n11827 );
    and g7398 ( n1640 , n3196 , n2274 );
    and g7399 ( n10097 , n4929 , n6833 );
    and g7400 ( n4056 , n10051 , n1836 );
    nor g7401 ( n3946 , n11069 , n10056 );
    nor g7402 ( n8999 , n9604 , n1743 );
    xnor g7403 ( n5874 , n11265 , n957 );
    and g7404 ( n7716 , n7731 , n3472 );
    and g7405 ( n11132 , n4973 , n12687 );
    or g7406 ( n3251 , n8870 , n1932 );
    or g7407 ( n2876 , n4539 , n893 );
    or g7408 ( n10541 , n10157 , n6138 );
    xnor g7409 ( n12057 , n8404 , n11739 );
    or g7410 ( n6437 , n11341 , n8484 );
    nor g7411 ( n4294 , n12788 , n11907 );
    not g7412 ( n9517 , n1820 );
    and g7413 ( n2793 , n10926 , n11396 );
    and g7414 ( n10159 , n10377 , n6673 );
    xnor g7415 ( n11537 , n9283 , n9623 );
    or g7416 ( n128 , n12119 , n4818 );
    or g7417 ( n12288 , n5915 , n2964 );
    not g7418 ( n11235 , n2537 );
    and g7419 ( n1231 , n3222 , n12228 );
    not g7420 ( n4661 , n7720 );
    and g7421 ( n10702 , n7965 , n10990 );
    or g7422 ( n7827 , n9389 , n7703 );
    xnor g7423 ( n498 , n6944 , n3897 );
    not g7424 ( n5759 , n11296 );
    xnor g7425 ( n978 , n8386 , n5136 );
    or g7426 ( n9656 , n10750 , n12686 );
    or g7427 ( n12955 , n12858 , n8742 );
    or g7428 ( n5373 , n3324 , n9160 );
    and g7429 ( n4967 , n2515 , n5645 );
    and g7430 ( n9036 , n6358 , n2749 );
    nor g7431 ( n9024 , n2979 , n4298 );
    and g7432 ( n6292 , n2287 , n12313 );
    xnor g7433 ( n2238 , n6810 , n635 );
    and g7434 ( n3703 , n6836 , n2004 );
    or g7435 ( n3878 , n3072 , n8111 );
    xnor g7436 ( n3744 , n9240 , n11671 );
    xnor g7437 ( n9623 , n9884 , n3411 );
    xnor g7438 ( n4852 , n370 , n2780 );
    xnor g7439 ( n4711 , n7322 , n256 );
    xnor g7440 ( n8604 , n11526 , n7175 );
    or g7441 ( n9339 , n11887 , n3924 );
    not g7442 ( n3856 , n1994 );
    xnor g7443 ( n9363 , n4563 , n8007 );
    nor g7444 ( n12896 , n2981 , n6444 );
    not g7445 ( n71 , n1412 );
    xnor g7446 ( n4191 , n7848 , n10574 );
    xnor g7447 ( n3460 , n9326 , n4920 );
    or g7448 ( n4608 , n1896 , n1135 );
    and g7449 ( n3219 , n6358 , n7294 );
    or g7450 ( n24 , n7283 , n1079 );
    and g7451 ( n8815 , n4613 , n4098 );
    not g7452 ( n11820 , n3022 );
    or g7453 ( n970 , n8295 , n5242 );
    and g7454 ( n5919 , n10417 , n10146 );
    and g7455 ( n11685 , n12468 , n1749 );
    and g7456 ( n6440 , n11038 , n12451 );
    or g7457 ( n9043 , n636 , n12080 );
    or g7458 ( n2272 , n11958 , n11896 );
    xnor g7459 ( n6935 , n7409 , n10099 );
    nor g7460 ( n11432 , n4468 , n7508 );
    or g7461 ( n10001 , n1407 , n4886 );
    and g7462 ( n3020 , n137 , n521 );
    xnor g7463 ( n7488 , n6937 , n12257 );
    xnor g7464 ( n6757 , n12374 , n7179 );
    nor g7465 ( n7444 , n9776 , n11649 );
    or g7466 ( n12447 , n1937 , n5540 );
    and g7467 ( n9829 , n5631 , n5068 );
    or g7468 ( n12262 , n8428 , n10903 );
    not g7469 ( n4481 , n5732 );
    and g7470 ( n961 , n953 , n10528 );
    not g7471 ( n1504 , n8184 );
    xnor g7472 ( n9359 , n7539 , n2078 );
    not g7473 ( n11403 , n7168 );
    or g7474 ( n189 , n1937 , n8768 );
    and g7475 ( n7001 , n1470 , n1917 );
    and g7476 ( n3296 , n4168 , n4572 );
    and g7477 ( n7214 , n6924 , n12527 );
    and g7478 ( n11201 , n1097 , n3842 );
    not g7479 ( n10919 , n12221 );
    xnor g7480 ( n5268 , n12781 , n3843 );
    xnor g7481 ( n1460 , n8341 , n8747 );
    xnor g7482 ( n7665 , n1462 , n10617 );
    xnor g7483 ( n1312 , n11589 , n9892 );
    xnor g7484 ( n3635 , n9346 , n12926 );
    not g7485 ( n3897 , n8783 );
    or g7486 ( n468 , n10097 , n2415 );
    or g7487 ( n7641 , n9982 , n2386 );
    xnor g7488 ( n9398 , n2449 , n5721 );
    and g7489 ( n12105 , n8164 , n4762 );
    or g7490 ( n8394 , n10196 , n10916 );
    or g7491 ( n8085 , n114 , n2815 );
    and g7492 ( n5838 , n10281 , n9087 );
    not g7493 ( n3142 , n9089 );
    or g7494 ( n1883 , n636 , n1932 );
    or g7495 ( n10783 , n989 , n10066 );
    and g7496 ( n8115 , n6391 , n5824 );
    xnor g7497 ( n8106 , n12794 , n8113 );
    xnor g7498 ( n1310 , n2203 , n6915 );
    or g7499 ( n9749 , n3127 , n12328 );
    or g7500 ( n589 , n10142 , n1546 );
    xnor g7501 ( n9968 , n5043 , n2237 );
    not g7502 ( n12013 , n5742 );
    or g7503 ( n8915 , n8026 , n8414 );
    xnor g7504 ( n1188 , n7528 , n12216 );
    and g7505 ( n5729 , n349 , n3520 );
    xnor g7506 ( n2054 , n6843 , n12156 );
    and g7507 ( n5789 , n2324 , n3730 );
    not g7508 ( n11488 , n11577 );
    or g7509 ( n9085 , n5172 , n3111 );
    or g7510 ( n8369 , n9370 , n3911 );
    xnor g7511 ( n6638 , n12098 , n3561 );
    xnor g7512 ( n11590 , n1157 , n12418 );
    or g7513 ( n8967 , n4213 , n6233 );
    xnor g7514 ( n7093 , n10060 , n11229 );
    xnor g7515 ( n366 , n7378 , n2914 );
    or g7516 ( n9087 , n3607 , n4794 );
    or g7517 ( n3725 , n6561 , n8008 );
    xnor g7518 ( n11797 , n9842 , n7080 );
    or g7519 ( n2167 , n10091 , n100 );
    not g7520 ( n11207 , n6990 );
    not g7521 ( n6286 , n12516 );
    nor g7522 ( n387 , n12223 , n7114 );
    and g7523 ( n2108 , n7160 , n7610 );
    and g7524 ( n1624 , n5053 , n12655 );
    nor g7525 ( n3481 , n2710 , n4982 );
    and g7526 ( n9734 , n6538 , n10035 );
    not g7527 ( n11493 , n9342 );
    xnor g7528 ( n11549 , n2036 , n2853 );
    xnor g7529 ( n6207 , n6426 , n11009 );
    xnor g7530 ( n7297 , n12857 , n2212 );
    xnor g7531 ( n2731 , n10544 , n3315 );
    or g7532 ( n148 , n10569 , n3479 );
    or g7533 ( n8304 , n8870 , n12735 );
    not g7534 ( n4179 , n4799 );
    and g7535 ( n2080 , n284 , n10693 );
    or g7536 ( n12696 , n7757 , n858 );
    or g7537 ( n11123 , n8959 , n11410 );
    or g7538 ( n7620 , n4498 , n7881 );
    or g7539 ( n12330 , n4206 , n4303 );
    xnor g7540 ( n10932 , n7415 , n1499 );
    xnor g7541 ( n2895 , n11373 , n9883 );
    or g7542 ( n9922 , n191 , n9397 );
    or g7543 ( n5582 , n11958 , n11775 );
    and g7544 ( n3016 , n10404 , n8624 );
    nor g7545 ( n9117 , n6930 , n8873 );
    and g7546 ( n4224 , n4287 , n12376 );
    xnor g7547 ( n10240 , n1783 , n906 );
    and g7548 ( n4895 , n3688 , n12045 );
    nor g7549 ( n4559 , n12309 , n4593 );
    or g7550 ( n11204 , n58 , n12426 );
    xnor g7551 ( n11314 , n11861 , n4410 );
    xnor g7552 ( n5799 , n10420 , n1875 );
    or g7553 ( n8387 , n191 , n7341 );
    and g7554 ( n7741 , n6996 , n1137 );
    xnor g7555 ( n4969 , n4508 , n8495 );
    and g7556 ( n8663 , n380 , n12540 );
    and g7557 ( n7300 , n8367 , n388 );
    nor g7558 ( n10203 , n6137 , n9404 );
    or g7559 ( n11349 , n11433 , n11820 );
    and g7560 ( n3521 , n1824 , n5011 );
    or g7561 ( n11305 , n10835 , n7506 );
    xnor g7562 ( n10460 , n8002 , n1494 );
    xnor g7563 ( n9891 , n2799 , n7711 );
    xnor g7564 ( n8581 , n12296 , n12877 );
    or g7565 ( n10148 , n3820 , n4875 );
    nor g7566 ( n119 , n5563 , n5749 );
    and g7567 ( n2479 , n1222 , n9417 );
    xnor g7568 ( n3990 , n2235 , n5763 );
    and g7569 ( n11061 , n5109 , n12295 );
    and g7570 ( n6213 , n9504 , n11910 );
    xnor g7571 ( n3657 , n12642 , n1589 );
    xnor g7572 ( n3287 , n6443 , n8820 );
    or g7573 ( n1500 , n3743 , n2020 );
    and g7574 ( n9633 , n6827 , n10221 );
    xnor g7575 ( n7592 , n7893 , n6344 );
    nor g7576 ( n7828 , n11068 , n7813 );
    xnor g7577 ( n3204 , n6792 , n6315 );
    not g7578 ( n10649 , n1088 );
    not g7579 ( n12871 , n223 );
    xnor g7580 ( n5536 , n6165 , n3663 );
    xnor g7581 ( n10853 , n10819 , n2776 );
    nor g7582 ( n450 , n1797 , n8525 );
    nor g7583 ( n10249 , n5139 , n5385 );
    not g7584 ( n5239 , n7428 );
    xnor g7585 ( n12637 , n7042 , n10717 );
    xnor g7586 ( n647 , n12315 , n1277 );
    not g7587 ( n6617 , n10163 );
    not g7588 ( n1128 , n4199 );
    not g7589 ( n11481 , n6688 );
    and g7590 ( n10867 , n11867 , n6075 );
    or g7591 ( n11271 , n8114 , n12902 );
    xnor g7592 ( n12020 , n467 , n10549 );
    xnor g7593 ( n5872 , n7308 , n12751 );
    nor g7594 ( n6679 , n3010 , n3702 );
    xnor g7595 ( n1912 , n4980 , n6139 );
    or g7596 ( n3335 , n6577 , n5538 );
    xnor g7597 ( n4470 , n4880 , n7931 );
    not g7598 ( n1261 , n9592 );
    xnor g7599 ( n8358 , n10740 , n4444 );
    nor g7600 ( n11548 , n10615 , n4699 );
    not g7601 ( n1022 , n10643 );
    and g7602 ( n2083 , n3862 , n57 );
    or g7603 ( n10173 , n7078 , n12905 );
    or g7604 ( n7804 , n12878 , n10906 );
    and g7605 ( n3519 , n5125 , n7598 );
    nor g7606 ( n2234 , n4278 , n9769 );
    not g7607 ( n12119 , n4805 );
    or g7608 ( n3123 , n10339 , n8109 );
    not g7609 ( n9644 , n9482 );
    not g7610 ( n1070 , n2968 );
    xnor g7611 ( n11217 , n4613 , n10352 );
    or g7612 ( n6088 , n11193 , n5636 );
    or g7613 ( n2822 , n6036 , n707 );
    or g7614 ( n9664 , n11849 , n7971 );
    or g7615 ( n5957 , n784 , n4440 );
    xnor g7616 ( n8385 , n9810 , n7183 );
    or g7617 ( n5152 , n1699 , n5468 );
    xor g7618 ( n12372 , n852 , n9711 );
    not g7619 ( n10 , n10987 );
    and g7620 ( n2537 , n4828 , n1512 );
    not g7621 ( n4343 , n4938 );
    and g7622 ( n4850 , n12241 , n9235 );
    or g7623 ( n8786 , n12119 , n12441 );
    nor g7624 ( n10071 , n10377 , n6673 );
    or g7625 ( n7872 , n6486 , n1464 );
    or g7626 ( n2681 , n5010 , n2080 );
    not g7627 ( n3370 , n12106 );
    or g7628 ( n12301 , n529 , n8272 );
    or g7629 ( n3698 , n5181 , n3410 );
    nor g7630 ( n2886 , n2997 , n6848 );
    nor g7631 ( n4737 , n547 , n2487 );
    and g7632 ( n1762 , n889 , n6430 );
    and g7633 ( n953 , n2564 , n11662 );
    not g7634 ( n8982 , n3517 );
    or g7635 ( n3506 , n386 , n9354 );
    xnor g7636 ( n7102 , n7769 , n1970 );
    xnor g7637 ( n4269 , n10139 , n3615 );
    and g7638 ( n4838 , n9010 , n10988 );
    and g7639 ( n5236 , n6877 , n2024 );
    and g7640 ( n1820 , n9372 , n3358 );
    or g7641 ( n4814 , n8512 , n3286 );
    or g7642 ( n4508 , n18 , n9599 );
    or g7643 ( n737 , n10196 , n3606 );
    or g7644 ( n3807 , n2217 , n4474 );
    or g7645 ( n6133 , n10750 , n7136 );
    not g7646 ( n1297 , n12280 );
    xnor g7647 ( n927 , n6673 , n12863 );
    not g7648 ( n12821 , n8487 );
    or g7649 ( n5458 , n252 , n3957 );
    not g7650 ( n2020 , n10990 );
    not g7651 ( n403 , n7748 );
    nor g7652 ( n3138 , n8548 , n6380 );
    not g7653 ( n10996 , n9263 );
    and g7654 ( n8450 , n890 , n2327 );
    nor g7655 ( n2160 , n9699 , n4684 );
    xnor g7656 ( n9655 , n5207 , n7367 );
    not g7657 ( n1834 , n5614 );
    or g7658 ( n12604 , n3743 , n3599 );
    or g7659 ( n11450 , n8870 , n7928 );
    xnor g7660 ( n7737 , n9922 , n7669 );
    or g7661 ( n4790 , n4778 , n1932 );
    or g7662 ( n6652 , n11433 , n11775 );
    nor g7663 ( n4575 , n12949 , n8289 );
    not g7664 ( n12579 , n9711 );
    or g7665 ( n10955 , n7116 , n6169 );
    nor g7666 ( n10060 , n12663 , n593 );
    or g7667 ( n7469 , n3127 , n2358 );
    xnor g7668 ( n2903 , n8542 , n8434 );
    xnor g7669 ( n12562 , n8862 , n6630 );
    and g7670 ( n12722 , n1177 , n5354 );
    xnor g7671 ( n4325 , n1596 , n2450 );
    and g7672 ( n10112 , n12303 , n1394 );
    xnor g7673 ( n12517 , n10552 , n11925 );
    xnor g7674 ( n7419 , n4511 , n2623 );
    and g7675 ( n11022 , n684 , n11483 );
    or g7676 ( n11181 , n9373 , n3606 );
    not g7677 ( n2334 , n2851 );
    xor g7678 ( n3071 , n12746 , n742 );
    xnor g7679 ( n944 , n1708 , n8882 );
    or g7680 ( n10937 , n1323 , n11688 );
    and g7681 ( n3651 , n147 , n12571 );
    or g7682 ( n3687 , n9917 , n9958 );
    and g7683 ( n10931 , n1449 , n1174 );
    and g7684 ( n9059 , n6672 , n1529 );
    or g7685 ( n12033 , n989 , n4242 );
    or g7686 ( n6789 , n8613 , n5943 );
    xnor g7687 ( n6992 , n10697 , n3995 );
    not g7688 ( n7371 , n8734 );
    or g7689 ( n11044 , n989 , n12843 );
    nor g7690 ( n5903 , n8605 , n2161 );
    and g7691 ( n11618 , n7485 , n6576 );
    nor g7692 ( n611 , n11109 , n80 );
    xnor g7693 ( n9919 , n12448 , n4930 );
    or g7694 ( n9108 , n994 , n1915 );
    or g7695 ( n4863 , n3127 , n6402 );
    xnor g7696 ( n9415 , n8361 , n9641 );
    xnor g7697 ( n4543 , n8147 , n5270 );
    or g7698 ( n5677 , n7526 , n790 );
    nor g7699 ( n6082 , n4738 , n2794 );
    and g7700 ( n2106 , n8600 , n2445 );
    and g7701 ( n3830 , n4995 , n1652 );
    xnor g7702 ( n7296 , n5967 , n7486 );
    xnor g7703 ( n9242 , n301 , n10285 );
    or g7704 ( n11121 , n10822 , n4711 );
    and g7705 ( n8176 , n5434 , n11354 );
    or g7706 ( n4382 , n1867 , n7371 );
    not g7707 ( n4262 , n2387 );
    or g7708 ( n2258 , n365 , n5457 );
    and g7709 ( n11810 , n6313 , n4816 );
    or g7710 ( n11767 , n7299 , n2239 );
    nor g7711 ( n6984 , n4147 , n9011 );
    not g7712 ( n6306 , n2116 );
    and g7713 ( n10293 , n7978 , n9566 );
    xnor g7714 ( n6771 , n10526 , n3458 );
    or g7715 ( n5769 , n10835 , n4864 );
    not g7716 ( n5025 , n6070 );
    xnor g7717 ( n11025 , n7098 , n2391 );
    not g7718 ( n2813 , n7244 );
    or g7719 ( n9800 , n12417 , n11590 );
    or g7720 ( n1673 , n986 , n11426 );
    xnor g7721 ( n6300 , n6408 , n528 );
    or g7722 ( n2539 , n2099 , n12754 );
    or g7723 ( n6486 , n7449 , n10916 );
    not g7724 ( n9172 , n11672 );
    and g7725 ( n7226 , n11384 , n668 );
    or g7726 ( n12271 , n5355 , n2076 );
    xnor g7727 ( n1588 , n7600 , n8463 );
    xnor g7728 ( n9467 , n8593 , n6511 );
    or g7729 ( n5569 , n8870 , n530 );
    not g7730 ( n11736 , n2402 );
    or g7731 ( n693 , n897 , n4850 );
    nor g7732 ( n9488 , n2563 , n2196 );
    or g7733 ( n4054 , n9500 , n9964 );
    xnor g7734 ( n10580 , n10221 , n5461 );
    or g7735 ( n10398 , n6078 , n2672 );
    or g7736 ( n4854 , n4979 , n8884 );
    xnor g7737 ( n2153 , n6731 , n2283 );
    xnor g7738 ( n8726 , n12248 , n1573 );
    and g7739 ( n11426 , n4213 , n6233 );
    and g7740 ( n12131 , n95 , n6792 );
    nor g7741 ( n3363 , n981 , n3296 );
    xnor g7742 ( n9630 , n6560 , n3741 );
    and g7743 ( n875 , n7874 , n12918 );
    and g7744 ( n1463 , n5183 , n6299 );
    or g7745 ( n2195 , n9648 , n5802 );
    nor g7746 ( n485 , n12670 , n8341 );
    nor g7747 ( n3373 , n7919 , n5872 );
    and g7748 ( n10500 , n11580 , n3823 );
    or g7749 ( n2329 , n2456 , n12124 );
    not g7750 ( n9276 , n662 );
    or g7751 ( n7686 , n9389 , n7881 );
    or g7752 ( n303 , n1404 , n10558 );
    or g7753 ( n5698 , n10771 , n11045 );
    xnor g7754 ( n8170 , n2161 , n8605 );
    xnor g7755 ( n3416 , n10288 , n7900 );
    xnor g7756 ( n8719 , n1152 , n10123 );
    xnor g7757 ( n10618 , n12319 , n2030 );
    or g7758 ( n5808 , n686 , n2815 );
    xnor g7759 ( n3812 , n9026 , n4683 );
    xnor g7760 ( n6835 , n9229 , n6762 );
    or g7761 ( n5408 , n3743 , n9521 );
    and g7762 ( n5608 , n2167 , n8413 );
    xnor g7763 ( n4137 , n5254 , n8264 );
    or g7764 ( n5887 , n8583 , n4527 );
    and g7765 ( n11927 , n10915 , n6020 );
    and g7766 ( n11194 , n2976 , n11495 );
    xnor g7767 ( n12498 , n11450 , n10908 );
    and g7768 ( n1105 , n5134 , n5477 );
    xnor g7769 ( n5566 , n3964 , n2981 );
    xnor g7770 ( n10819 , n2119 , n2264 );
    not g7771 ( n795 , n8028 );
    or g7772 ( n5802 , n8959 , n11775 );
    xnor g7773 ( n2859 , n9204 , n8693 );
    or g7774 ( n762 , n2456 , n1932 );
    or g7775 ( n7188 , n3096 , n6455 );
    or g7776 ( n6203 , n4059 , n4242 );
    not g7777 ( n8285 , n6441 );
    xnor g7778 ( n3727 , n2029 , n8500 );
    xnor g7779 ( n1544 , n10128 , n2451 );
    or g7780 ( n1909 , n9656 , n12411 );
    or g7781 ( n12880 , n9812 , n10836 );
    or g7782 ( n10740 , n4662 , n8987 );
    not g7783 ( n304 , n4484 );
    and g7784 ( n4317 , n4547 , n7335 );
    xnor g7785 ( n8390 , n7200 , n7499 );
    and g7786 ( n8526 , n4772 , n9470 );
    or g7787 ( n8908 , n12361 , n10919 );
    xnor g7788 ( n6624 , n7365 , n1753 );
    not g7789 ( n1861 , n4439 );
    and g7790 ( n10624 , n12344 , n815 );
    or g7791 ( n9682 , n2367 , n795 );
    or g7792 ( n7688 , n4628 , n12686 );
    not g7793 ( n8859 , n1835 );
    or g7794 ( n10216 , n8159 , n5299 );
    xnor g7795 ( n82 , n12348 , n9399 );
    xnor g7796 ( n746 , n3437 , n12075 );
    xnor g7797 ( n2775 , n12052 , n6440 );
    xnor g7798 ( n7308 , n1631 , n7296 );
    or g7799 ( n9531 , n10157 , n4654 );
    nor g7800 ( n4147 , n9369 , n2952 );
    xnor g7801 ( n11588 , n11262 , n9056 );
    or g7802 ( n7244 , n11552 , n4654 );
    or g7803 ( n8120 , n5504 , n9925 );
    and g7804 ( n3186 , n3930 , n4483 );
    and g7805 ( n12024 , n9827 , n11599 );
    xnor g7806 ( n657 , n7662 , n1800 );
    not g7807 ( n9856 , n1050 );
    nor g7808 ( n5854 , n6472 , n2174 );
    or g7809 ( n2629 , n5945 , n6455 );
    xnor g7810 ( n3384 , n7520 , n9133 );
    xnor g7811 ( n8391 , n1151 , n6998 );
    or g7812 ( n5662 , n9498 , n3880 );
    xnor g7813 ( n2449 , n9155 , n3395 );
    xnor g7814 ( n6591 , n7790 , n6416 );
    or g7815 ( n2251 , n6667 , n604 );
    xnor g7816 ( n3839 , n12443 , n1734 );
    not g7817 ( n4896 , n4850 );
    nor g7818 ( n4211 , n7916 , n2642 );
    not g7819 ( n12199 , n1456 );
    nor g7820 ( n4036 , n4588 , n7660 );
    xnor g7821 ( n9136 , n1228 , n7560 );
    or g7822 ( n10338 , n2217 , n8643 );
    or g7823 ( n3997 , n5809 , n4818 );
    xnor g7824 ( n9722 , n8617 , n2375 );
    or g7825 ( n2159 , n6924 , n12527 );
    or g7826 ( n1052 , n7024 , n4661 );
    not g7827 ( n2994 , n3734 );
    or g7828 ( n1696 , n8583 , n4474 );
    xnor g7829 ( n5509 , n1624 , n6194 );
    xnor g7830 ( n1954 , n5825 , n12620 );
    not g7831 ( n4085 , n8760 );
    or g7832 ( n9061 , n11714 , n5551 );
    not g7833 ( n9772 , n5344 );
    or g7834 ( n11704 , n191 , n130 );
    not g7835 ( n11193 , n7416 );
    or g7836 ( n5285 , n8416 , n2933 );
    or g7837 ( n8790 , n752 , n2232 );
    not g7838 ( n1790 , n8204 );
    xnor g7839 ( n9072 , n12287 , n241 );
    xnor g7840 ( n10779 , n10038 , n9451 );
    not g7841 ( n6627 , n8094 );
    or g7842 ( n9150 , n6577 , n12816 );
    not g7843 ( n7683 , n11243 );
    or g7844 ( n8045 , n5575 , n12357 );
    or g7845 ( n3761 , n3127 , n12843 );
    and g7846 ( n2149 , n4679 , n1668 );
    xnor g7847 ( n4486 , n12611 , n10753 );
    not g7848 ( n10479 , n10402 );
    or g7849 ( n11931 , n9171 , n9221 );
    xnor g7850 ( n2365 , n4991 , n7427 );
    xnor g7851 ( n9810 , n8275 , n9052 );
    xnor g7852 ( n12552 , n5948 , n233 );
    and g7853 ( n7979 , n11255 , n2591 );
    xnor g7854 ( n5742 , n4465 , n475 );
    xnor g7855 ( n8350 , n5486 , n3662 );
    or g7856 ( n11878 , n10611 , n7249 );
    or g7857 ( n4546 , n7116 , n5012 );
    xnor g7858 ( n1301 , n262 , n5634 );
    and g7859 ( n4057 , n5233 , n11201 );
    or g7860 ( n11687 , n989 , n8524 );
    or g7861 ( n12041 , n6042 , n576 );
    xor g7862 ( n635 , n3018 , n11831 );
    and g7863 ( n7158 , n3976 , n12059 );
    nor g7864 ( n3195 , n4908 , n6596 );
    xnor g7865 ( n7605 , n6153 , n9374 );
    not g7866 ( n7273 , n3020 );
    or g7867 ( n12398 , n7420 , n12475 );
    xnor g7868 ( n1492 , n12324 , n2736 );
    xnor g7869 ( n12911 , n4148 , n8399 );
    and g7870 ( n2871 , n9634 , n1250 );
    not g7871 ( n1641 , n633 );
    or g7872 ( n8332 , n7052 , n1864 );
    not g7873 ( n8363 , n9757 );
    xor g7874 ( n7253 , n1951 , n3432 );
    or g7875 ( n2270 , n6516 , n4321 );
    xnor g7876 ( n360 , n178 , n5387 );
    not g7877 ( n4624 , n1826 );
    or g7878 ( n1706 , n2217 , n28 );
    not g7879 ( n2384 , n6661 );
    nor g7880 ( n11991 , n4595 , n5624 );
    or g7881 ( n6058 , n6977 , n3468 );
    or g7882 ( n3029 , n8354 , n4913 );
    and g7883 ( n36 , n4387 , n4162 );
    or g7884 ( n5600 , n7391 , n11746 );
    nor g7885 ( n8036 , n4906 , n9830 );
    not g7886 ( n4527 , n11876 );
    xnor g7887 ( n7877 , n4283 , n10925 );
    or g7888 ( n2274 , n6017 , n7056 );
    xnor g7889 ( n9567 , n9203 , n66 );
    xnor g7890 ( n5693 , n6640 , n9463 );
    or g7891 ( n6783 , n10749 , n7229 );
    not g7892 ( n4327 , n6129 );
    and g7893 ( n6745 , n6369 , n3522 );
    nor g7894 ( n3365 , n8194 , n4035 );
    xnor g7895 ( n207 , n1811 , n829 );
    and g7896 ( n9123 , n294 , n7023 );
    xnor g7897 ( n11209 , n1809 , n8290 );
    nor g7898 ( n593 , n3441 , n2121 );
    xnor g7899 ( n12921 , n7189 , n3107 );
    or g7900 ( n8901 , n1472 , n5 );
    and g7901 ( n1322 , n5425 , n2245 );
    or g7902 ( n10956 , n525 , n8058 );
    nor g7903 ( n12500 , n9014 , n10933 );
    nor g7904 ( n7972 , n9708 , n3779 );
    or g7905 ( n9933 , n8267 , n11939 );
    not g7906 ( n5388 , n2166 );
    or g7907 ( n7089 , n5919 , n9242 );
    or g7908 ( n8189 , n994 , n7424 );
    xnor g7909 ( n1027 , n9307 , n1948 );
    xnor g7910 ( n5041 , n6704 , n6428 );
    xnor g7911 ( n2032 , n8647 , n8408 );
    and g7912 ( n8376 , n5205 , n1662 );
    xnor g7913 ( n8715 , n9469 , n10314 );
    xnor g7914 ( n8300 , n5323 , n9025 );
    xnor g7915 ( n8914 , n10483 , n7852 );
    or g7916 ( n1275 , n7495 , n11827 );
    xnor g7917 ( n4705 , n5279 , n2147 );
    not g7918 ( n9710 , n12089 );
    xnor g7919 ( n751 , n4301 , n11741 );
    and g7920 ( n11813 , n5614 , n12895 );
    or g7921 ( n7462 , n2099 , n12735 );
    or g7922 ( n7251 , n8026 , n995 );
    or g7923 ( n7084 , n752 , n11896 );
    and g7924 ( n6067 , n7233 , n10059 );
    and g7925 ( n3615 , n1514 , n1149 );
    and g7926 ( n7919 , n2002 , n12342 );
    xnor g7927 ( n2836 , n196 , n11477 );
    not g7928 ( n1923 , n7342 );
    or g7929 ( n7256 , n9110 , n10628 );
    xnor g7930 ( n5381 , n2142 , n6216 );
    not g7931 ( n518 , n2630 );
    nor g7932 ( n6009 , n885 , n5836 );
    or g7933 ( n8692 , n5765 , n8830 );
    or g7934 ( n7071 , n10142 , n6402 );
    and g7935 ( n2986 , n2982 , n4319 );
    or g7936 ( n1260 , n7495 , n7341 );
    and g7937 ( n8865 , n8295 , n5242 );
    xnor g7938 ( n8706 , n9450 , n11002 );
    or g7939 ( n11533 , n10750 , n9586 );
    or g7940 ( n8978 , n11026 , n12771 );
    or g7941 ( n6251 , n2171 , n10445 );
    or g7942 ( n7661 , n1598 , n5564 );
    or g7943 ( n2112 , n12116 , n6938 );
    xnor g7944 ( n7255 , n9595 , n162 );
    xnor g7945 ( n6427 , n9785 , n7764 );
    xnor g7946 ( n1479 , n2542 , n12206 );
    and g7947 ( n4883 , n7388 , n11876 );
    and g7948 ( n1748 , n639 , n1669 );
    xnor g7949 ( n7868 , n5508 , n3349 );
    and g7950 ( n11971 , n3032 , n281 );
    or g7951 ( n5323 , n1764 , n3495 );
    and g7952 ( n3157 , n1705 , n12251 );
    and g7953 ( n11446 , n11416 , n2535 );
    not g7954 ( n2189 , n2181 );
    or g7955 ( n8286 , n8583 , n4654 );
    nor g7956 ( n9988 , n3706 , n10461 );
    not g7957 ( n4193 , n2858 );
    and g7958 ( n1710 , n505 , n12592 );
    nor g7959 ( n883 , n12210 , n601 );
    xnor g7960 ( n11160 , n1988 , n4194 );
    xnor g7961 ( n1040 , n6782 , n1503 );
    xnor g7962 ( n1003 , n8347 , n8488 );
    or g7963 ( n5203 , n10697 , n4968 );
    not g7964 ( n3488 , n11467 );
    and g7965 ( n7905 , n5663 , n11387 );
    and g7966 ( n9883 , n2466 , n10806 );
    not g7967 ( n3451 , n1357 );
    xnor g7968 ( n10371 , n10563 , n7222 );
    not g7969 ( n12349 , n11040 );
    and g7970 ( n5622 , n11478 , n12925 );
    or g7971 ( n9076 , n12227 , n11940 );
    not g7972 ( n8305 , n8044 );
    not g7973 ( n11731 , n1750 );
    or g7974 ( n8866 , n282 , n7494 );
    xnor g7975 ( n10713 , n10381 , n2837 );
    and g7976 ( n1106 , n12552 , n6989 );
    or g7977 ( n8778 , n8583 , n9568 );
    not g7978 ( n6847 , n9450 );
    not g7979 ( n4573 , n6998 );
    xnor g7980 ( n2299 , n1223 , n9500 );
    not g7981 ( n12028 , n8420 );
    not g7982 ( n2242 , n12915 );
    nor g7983 ( n10201 , n9476 , n10602 );
    xnor g7984 ( n9201 , n1321 , n10886 );
    xnor g7985 ( n7524 , n1921 , n12402 );
    or g7986 ( n10038 , n191 , n6524 );
    nor g7987 ( n2747 , n10318 , n10110 );
    xnor g7988 ( n5286 , n7616 , n1723 );
    and g7989 ( n10025 , n8310 , n2912 );
    or g7990 ( n8456 , n5858 , n3911 );
    not g7991 ( n184 , n11423 );
    xnor g7992 ( n9438 , n2305 , n10643 );
    xnor g7993 ( n9557 , n4174 , n4470 );
    or g7994 ( n8063 , n1699 , n8259 );
    and g7995 ( n8772 , n10928 , n7946 );
    xnor g7996 ( n933 , n11413 , n5653 );
    xnor g7997 ( n3805 , n11637 , n11738 );
    xnor g7998 ( n12671 , n7311 , n10151 );
    xnor g7999 ( n1332 , n2842 , n6260 );
    nor g8000 ( n12007 , n4154 , n5746 );
    or g8001 ( n11495 , n989 , n6389 );
    and g8002 ( n7995 , n6943 , n7182 );
    and g8003 ( n3608 , n8622 , n6200 );
    not g8004 ( n4050 , n1021 );
    and g8005 ( n554 , n10774 , n6765 );
    or g8006 ( n9353 , n10750 , n3224 );
    not g8007 ( n7246 , n4005 );
    xnor g8008 ( n7496 , n551 , n7975 );
    or g8009 ( n9735 , n4628 , n6071 );
    xnor g8010 ( n9487 , n12619 , n10166 );
    xnor g8011 ( n4603 , n2878 , n10786 );
    not g8012 ( n3864 , n4678 );
    and g8013 ( n5711 , n6740 , n9524 );
    xnor g8014 ( n9784 , n7331 , n1865 );
    not g8015 ( n7149 , n6954 );
    not g8016 ( n5574 , n7520 );
    nor g8017 ( n3784 , n3659 , n4993 );
    or g8018 ( n11307 , n1882 , n2043 );
    or g8019 ( n1887 , n4647 , n11236 );
    not g8020 ( n11811 , n7289 );
    xnor g8021 ( n10495 , n255 , n6879 );
    or g8022 ( n3494 , n7662 , n1800 );
    and g8023 ( n9827 , n10780 , n12942 );
    or g8024 ( n7914 , n11958 , n7558 );
    xnor g8025 ( n2514 , n11664 , n8314 );
    or g8026 ( n966 , n994 , n12843 );
    or g8027 ( n5282 , n11433 , n2815 );
    nor g8028 ( n11332 , n8376 , n1378 );
    and g8029 ( n5076 , n11451 , n6466 );
    not g8030 ( n824 , n6322 );
    xnor g8031 ( n8472 , n6730 , n7510 );
    xnor g8032 ( n4435 , n9263 , n8292 );
    xnor g8033 ( n865 , n10191 , n9654 );
    and g8034 ( n8983 , n12871 , n5649 );
    and g8035 ( n7384 , n7462 , n2105 );
    and g8036 ( n5360 , n10381 , n6177 );
    not g8037 ( n11696 , n10857 );
    or g8038 ( n1960 , n989 , n1851 );
    xnor g8039 ( n5568 , n7020 , n5668 );
    or g8040 ( n9341 , n3127 , n1915 );
    xnor g8041 ( n5942 , n11488 , n192 );
    or g8042 ( n891 , n3820 , n4474 );
    or g8043 ( n2430 , n12361 , n5540 );
    or g8044 ( n10798 , n11552 , n9521 );
    or g8045 ( n2363 , n191 , n12328 );
    or g8046 ( n11867 , n9389 , n7341 );
    nor g8047 ( n2328 , n8592 , n5609 );
    not g8048 ( n1915 , n7456 );
    or g8049 ( n1249 , n191 , n4242 );
    xnor g8050 ( n7602 , n8333 , n5446 );
    and g8051 ( n3011 , n4805 , n1067 );
    xnor g8052 ( n6708 , n5035 , n4003 );
    or g8053 ( n5922 , n11958 , n12274 );
    and g8054 ( n8258 , n11534 , n483 );
    or g8055 ( n9013 , n10389 , n9041 );
    xnor g8056 ( n840 , n11086 , n5120 );
    not g8057 ( n4320 , n12733 );
    nor g8058 ( n8713 , n9849 , n8268 );
    or g8059 ( n9372 , n2312 , n3899 );
    or g8060 ( n9232 , n12715 , n7065 );
    xnor g8061 ( n5907 , n4491 , n235 );
    xnor g8062 ( n5083 , n7899 , n10565 );
    not g8063 ( n2637 , n11758 );
    xnor g8064 ( n8899 , n5894 , n9436 );
    or g8065 ( n2359 , n12503 , n9160 );
    and g8066 ( n11170 , n3464 , n8805 );
    xnor g8067 ( n3456 , n8160 , n7692 );
    or g8068 ( n9742 , n6758 , n3387 );
    or g8069 ( n7983 , n2456 , n9586 );
    xnor g8070 ( n10519 , n5888 , n12923 );
    or g8071 ( n4127 , n10960 , n10315 );
    not g8072 ( n2969 , n2 );
    or g8073 ( n2230 , n994 , n561 );
    or g8074 ( n4277 , n5510 , n6609 );
    not g8075 ( n10611 , n5606 );
    or g8076 ( n2915 , n4674 , n12535 );
    xnor g8077 ( n10357 , n6012 , n5440 );
    not g8078 ( n3095 , n11594 );
    nor g8079 ( n12876 , n6009 , n1613 );
    or g8080 ( n8195 , n11887 , n8109 );
    xnor g8081 ( n912 , n10768 , n328 );
    xnor g8082 ( n1033 , n8146 , n5613 );
    xnor g8083 ( n1753 , n4576 , n8052 );
    or g8084 ( n6162 , n3724 , n53 );
    and g8085 ( n7994 , n11850 , n5458 );
    not g8086 ( n9835 , n250 );
    xnor g8087 ( n8081 , n622 , n7987 );
    xnor g8088 ( n774 , n6316 , n210 );
    xnor g8089 ( n2176 , n2635 , n1232 );
    or g8090 ( n9946 , n1699 , n8644 );
    not g8091 ( n8774 , n6867 );
    nor g8092 ( n7026 , n10052 , n7353 );
    or g8093 ( n9303 , n6373 , n4864 );
    nor g8094 ( n1234 , n5067 , n12236 );
    not g8095 ( n11304 , n12573 );
    or g8096 ( n11203 , n994 , n4775 );
    xnor g8097 ( n7151 , n8634 , n11370 );
    xnor g8098 ( n2891 , n5873 , n8867 );
    not g8099 ( n2034 , n7983 );
    nor g8100 ( n6862 , n7845 , n5222 );
    or g8101 ( n7184 , n12244 , n9425 );
    nor g8102 ( n4081 , n6919 , n4935 );
    nor g8103 ( n3496 , n3585 , n6383 );
    or g8104 ( n5491 , n7116 , n995 );
    or g8105 ( n9441 , n8920 , n8547 );
    or g8106 ( n857 , n6331 , n9550 );
    not g8107 ( n2135 , n531 );
    nor g8108 ( n3241 , n4806 , n10449 );
    or g8109 ( n4740 , n10798 , n10133 );
    not g8110 ( n12924 , n12266 );
    xnor g8111 ( n4230 , n5447 , n4621 );
    not g8112 ( n11421 , n1810 );
    not g8113 ( n2927 , n10834 );
    xnor g8114 ( n9578 , n1669 , n5142 );
    xnor g8115 ( n10345 , n12204 , n1858 );
    not g8116 ( n10301 , n2321 );
    xnor g8117 ( n35 , n5570 , n8963 );
    or g8118 ( n3408 , n8601 , n2737 );
    xnor g8119 ( n3514 , n2190 , n2663 );
    xnor g8120 ( n9491 , n12377 , n8881 );
    nor g8121 ( n9511 , n10830 , n1631 );
    or g8122 ( n9785 , n11552 , n4875 );
    or g8123 ( n6583 , n9751 , n10758 );
    xnor g8124 ( n1124 , n1826 , n8280 );
    and g8125 ( n10648 , n2380 , n8177 );
    or g8126 ( n10717 , n10163 , n10321 );
    not g8127 ( n9694 , n5845 );
    not g8128 ( n11316 , n5978 );
    xnor g8129 ( n9109 , n1715 , n2961 );
    not g8130 ( n12655 , n7442 );
    xnor g8131 ( n2029 , n3180 , n10086 );
    not g8132 ( n11082 , n167 );
    and g8133 ( n6186 , n8480 , n5865 );
    xnor g8134 ( n9901 , n4948 , n11275 );
    or g8135 ( n6230 , n10424 , n7245 );
    not g8136 ( n834 , n990 );
    or g8137 ( n8694 , n7449 , n5502 );
    or g8138 ( n7185 , n12119 , n8259 );
    nor g8139 ( n3573 , n2 , n11783 );
    or g8140 ( n10818 , n12263 , n9203 );
    xnor g8141 ( n12919 , n2570 , n5038 );
    xnor g8142 ( n7535 , n12286 , n11836 );
    and g8143 ( n10191 , n9730 , n3306 );
    xnor g8144 ( n6580 , n10324 , n7333 );
    or g8145 ( n6790 , n12341 , n3075 );
    and g8146 ( n2739 , n12199 , n4028 );
    and g8147 ( n8750 , n10762 , n11365 );
    and g8148 ( n630 , n8598 , n5581 );
    or g8149 ( n10790 , n1183 , n3224 );
    and g8150 ( n10280 , n3066 , n8669 );
    or g8151 ( n8549 , n2791 , n278 );
    and g8152 ( n12396 , n11245 , n2673 );
    and g8153 ( n3560 , n3905 , n2270 );
    or g8154 ( n7655 , n10157 , n4864 );
    or g8155 ( n8143 , n4916 , n1263 );
    xnor g8156 ( n5 , n11790 , n2280 );
    or g8157 ( n11324 , n8026 , n7558 );
    or g8158 ( n6661 , n1941 , n5540 );
    or g8159 ( n6704 , n6373 , n9521 );
    and g8160 ( n6749 , n58 , n12426 );
    xnor g8161 ( n12224 , n11721 , n4146 );
    and g8162 ( n3056 , n5990 , n11078 );
    or g8163 ( n3340 , n11026 , n1476 );
    not g8164 ( n5781 , n1353 );
    and g8165 ( n5048 , n10360 , n12013 );
    not g8166 ( n6170 , n1306 );
    not g8167 ( n11655 , n12219 );
    not g8168 ( n5773 , n12520 );
    or g8169 ( n4948 , n8870 , n5326 );
    not g8170 ( n12384 , n11884 );
    not g8171 ( n5974 , n7778 );
    or g8172 ( n11387 , n9426 , n5790 );
    not g8173 ( n651 , n8048 );
    not g8174 ( n8608 , n7151 );
    or g8175 ( n10993 , n6671 , n4526 );
    xnor g8176 ( n6188 , n8013 , n1075 );
    nor g8177 ( n8037 , n8162 , n9845 );
    not g8178 ( n3679 , n7187 );
    or g8179 ( n12023 , n752 , n3421 );
    and g8180 ( n11997 , n1796 , n10623 );
    xnor g8181 ( n12445 , n3794 , n12285 );
    and g8182 ( n8342 , n2052 , n1367 );
    not g8183 ( n4288 , n6879 );
    and g8184 ( n3957 , n6738 , n11179 );
    xnor g8185 ( n5968 , n11182 , n4200 );
    or g8186 ( n12061 , n1699 , n8109 );
    xnor g8187 ( n2471 , n1991 , n6692 );
    xnor g8188 ( n3281 , n8602 , n5897 );
    and g8189 ( n2569 , n11511 , n6885 );
    xor g8190 ( n1645 , n12647 , n10665 );
    xnor g8191 ( n7229 , n12742 , n11768 );
    xnor g8192 ( n12353 , n8515 , n6760 );
    or g8193 ( n5564 , n3892 , n10358 );
    and g8194 ( n1502 , n11528 , n2654 );
    xnor g8195 ( n12309 , n11908 , n7578 );
    nor g8196 ( n6927 , n8155 , n4408 );
    xnor g8197 ( n12751 , n9059 , n6865 );
    and g8198 ( n11267 , n4056 , n2169 );
    xnor g8199 ( n11585 , n3837 , n9096 );
    and g8200 ( n11840 , n10670 , n5488 );
    or g8201 ( n4596 , n1100 , n7763 );
    and g8202 ( n11785 , n7688 , n11465 );
    or g8203 ( n11567 , n7587 , n2343 );
    and g8204 ( n12830 , n2697 , n11348 );
    not g8205 ( n11411 , n2470 );
    xnor g8206 ( n11073 , n1782 , n12598 );
    not g8207 ( n12172 , n6660 );
    nor g8208 ( n3225 , n10909 , n3496 );
    xnor g8209 ( n9577 , n1956 , n8570 );
    or g8210 ( n3907 , n1993 , n5090 );
    or g8211 ( n11747 , n5840 , n6614 );
    or g8212 ( n5134 , n11036 , n8030 );
    xnor g8213 ( n11210 , n4489 , n7013 );
    not g8214 ( n12598 , n4834 );
    or g8215 ( n11037 , n8870 , n4913 );
    and g8216 ( n2811 , n1653 , n10896 );
    not g8217 ( n12030 , n4999 );
    or g8218 ( n12324 , n11958 , n8768 );
    and g8219 ( n5973 , n7889 , n11993 );
    xnor g8220 ( n5421 , n9764 , n3997 );
    and g8221 ( n555 , n3011 , n8660 );
    nor g8222 ( n10054 , n3369 , n9471 );
    not g8223 ( n7422 , n10009 );
    and g8224 ( n3308 , n7251 , n4264 );
    and g8225 ( n12417 , n2045 , n11274 );
    or g8226 ( n1521 , n4696 , n2475 );
    not g8227 ( n6048 , n3824 );
    xnor g8228 ( n2729 , n9522 , n2205 );
    or g8229 ( n1021 , n11283 , n12773 );
    or g8230 ( n4205 , n1941 , n7876 );
    xnor g8231 ( n11167 , n10560 , n2889 );
    xnor g8232 ( n7018 , n4942 , n7580 );
    or g8233 ( n1746 , n10835 , n8285 );
    and g8234 ( n4834 , n2530 , n2802 );
    not g8235 ( n5523 , n5291 );
    or g8236 ( n5786 , n7283 , n5497 );
    xnor g8237 ( n8696 , n11029 , n10800 );
    or g8238 ( n8590 , n8687 , n28 );
    not g8239 ( n1163 , n11922 );
    nor g8240 ( n10298 , n9489 , n8935 );
    or g8241 ( n4295 , n167 , n408 );
    or g8242 ( n6592 , n2025 , n5322 );
    or g8243 ( n6115 , n12262 , n8253 );
    not g8244 ( n3025 , n5728 );
    not g8245 ( n3759 , n2714 );
    or g8246 ( n12819 , n8949 , n6724 );
    not g8247 ( n12297 , n7331 );
    or g8248 ( n2214 , n8332 , n10866 );
    or g8249 ( n7014 , n11550 , n7051 );
    nor g8250 ( n5494 , n10257 , n8868 );
    xnor g8251 ( n4049 , n4212 , n1485 );
    or g8252 ( n4769 , n4176 , n3948 );
    xnor g8253 ( n11442 , n6464 , n9143 );
    or g8254 ( n7473 , n8848 , n1008 );
    or g8255 ( n9322 , n6718 , n4474 );
    and g8256 ( n794 , n2950 , n1164 );
    xnor g8257 ( n11555 , n12445 , n1351 );
    not g8258 ( n8842 , n4028 );
    not g8259 ( n375 , n11834 );
    or g8260 ( n2127 , n10157 , n12771 );
    not g8261 ( n3556 , n625 );
    xnor g8262 ( n336 , n7978 , n4997 );
    and g8263 ( n7954 , n5283 , n521 );
    xnor g8264 ( n950 , n6221 , n11379 );
    or g8265 ( n11184 , n3096 , n1413 );
    and g8266 ( n43 , n925 , n1958 );
    or g8267 ( n10902 , n9655 , n12580 );
    not g8268 ( n6526 , n10243 );
    not g8269 ( n11923 , n5314 );
    not g8270 ( n3548 , n1822 );
    and g8271 ( n12541 , n9400 , n10439 );
    or g8272 ( n10527 , n3324 , n4527 );
    or g8273 ( n8949 , n5575 , n3468 );
    xnor g8274 ( n1535 , n6954 , n3812 );
    xnor g8275 ( n8110 , n3079 , n9237 );
    not g8276 ( n1600 , n1294 );
    or g8277 ( n11856 , n8428 , n9741 );
    and g8278 ( n8101 , n1760 , n2859 );
    xnor g8279 ( n11188 , n5277 , n6240 );
    xnor g8280 ( n3723 , n12354 , n7165 );
    or g8281 ( n3873 , n6977 , n5538 );
    and g8282 ( n11225 , n12069 , n1512 );
    and g8283 ( n102 , n4734 , n11489 );
    or g8284 ( n6318 , n1941 , n1413 );
    xnor g8285 ( n8993 , n10945 , n5348 );
    not g8286 ( n5631 , n2030 );
    and g8287 ( n10443 , n4150 , n4627 );
    nor g8288 ( n11903 , n11831 , n12798 );
    not g8289 ( n1253 , n812 );
    xnor g8290 ( n11146 , n12935 , n9808 );
    and g8291 ( n8455 , n6411 , n4132 );
    or g8292 ( n2905 , n8026 , n6114 );
    xnor g8293 ( n7072 , n2726 , n3289 );
    or g8294 ( n12862 , n10712 , n5583 );
    and g8295 ( n9193 , n1226 , n2750 );
    or g8296 ( n1962 , n10135 , n9854 );
    and g8297 ( n11321 , n4120 , n2805 );
    or g8298 ( n9674 , n191 , n1738 );
    xnor g8299 ( n7132 , n3387 , n12334 );
    xnor g8300 ( n8174 , n2567 , n2455 );
    xnor g8301 ( n3371 , n2928 , n12650 );
    not g8302 ( n11619 , n11017 );
    not g8303 ( n1391 , n2937 );
    and g8304 ( n11230 , n10772 , n10793 );
    xnor g8305 ( n10273 , n10997 , n10940 );
    xnor g8306 ( n6500 , n3936 , n1946 );
    xnor g8307 ( n10264 , n8176 , n324 );
    xnor g8308 ( n3802 , n10722 , n5535 );
    and g8309 ( n2633 , n7084 , n9091 );
    or g8310 ( n10929 , n3820 , n28 );
    and g8311 ( n4581 , n3316 , n7888 );
    or g8312 ( n11255 , n2155 , n11112 );
    not g8313 ( n4204 , n3247 );
    and g8314 ( n9038 , n2718 , n4611 );
    or g8315 ( n577 , n8354 , n826 );
    xnor g8316 ( n103 , n3130 , n7555 );
    not g8317 ( n4365 , n5263 );
    or g8318 ( n10778 , n4383 , n6297 );
    or g8319 ( n4812 , n10590 , n7821 );
    or g8320 ( n1829 , n6373 , n7921 );
    xnor g8321 ( n1517 , n3970 , n7091 );
    nor g8322 ( n12663 , n11080 , n12597 );
    not g8323 ( n11473 , n3825 );
    not g8324 ( n12957 , n7807 );
    nor g8325 ( n1208 , n4788 , n9620 );
    xnor g8326 ( n5987 , n5492 , n10072 );
    xnor g8327 ( n6495 , n5921 , n7360 );
    not g8328 ( n7476 , n6527 );
    not g8329 ( n9074 , n5582 );
    xnor g8330 ( n7934 , n2993 , n6468 );
    or g8331 ( n12539 , n7116 , n11896 );
    xnor g8332 ( n4163 , n9926 , n1969 );
    nor g8333 ( n7372 , n9305 , n6205 );
    and g8334 ( n5233 , n5964 , n2577 );
    or g8335 ( n3659 , n5575 , n6114 );
    not g8336 ( n11228 , n2443 );
    and g8337 ( n12070 , n6893 , n1068 );
    xnor g8338 ( n6240 , n5087 , n5357 );
    or g8339 ( n8779 , n8026 , n12816 );
    xnor g8340 ( n11445 , n9613 , n4425 );
    and g8341 ( n9465 , n4312 , n7456 );
    or g8342 ( n9413 , n11958 , n995 );
    xnor g8343 ( n1203 , n10703 , n12311 );
    nor g8344 ( n7197 , n9438 , n8982 );
    xnor g8345 ( n4076 , n12176 , n7150 );
    or g8346 ( n11392 , n6718 , n5502 );
    xnor g8347 ( n12852 , n9043 , n10840 );
    and g8348 ( n6729 , n3848 , n4974 );
    nor g8349 ( n7769 , n9643 , n10076 );
    or g8350 ( n8054 , n1937 , n6169 );
    and g8351 ( n10868 , n5832 , n6531 );
    xnor g8352 ( n6815 , n6341 , n4419 );
    or g8353 ( n6463 , n3007 , n8561 );
    or g8354 ( n60 , n11958 , n6084 );
    and g8355 ( n478 , n8337 , n5622 );
    xnor g8356 ( n2884 , n10918 , n6420 );
    xnor g8357 ( n8361 , n9392 , n7263 );
    and g8358 ( n9964 , n1223 , n2892 );
    not g8359 ( n11638 , n12564 );
    or g8360 ( n4699 , n11572 , n3192 );
    or g8361 ( n10518 , n6718 , n9160 );
    not g8362 ( n7687 , n2643 );
    not g8363 ( n692 , n8694 );
    not g8364 ( n5402 , n1481 );
    not g8365 ( n12079 , n649 );
    or g8366 ( n6853 , n962 , n28 );
    not g8367 ( n9589 , n9725 );
    or g8368 ( n5797 , n9370 , n1162 );
    and g8369 ( n5971 , n6914 , n4447 );
    xnor g8370 ( n1056 , n2763 , n12633 );
    or g8371 ( n11456 , n3617 , n10854 );
    xnor g8372 ( n2685 , n12960 , n10487 );
    xnor g8373 ( n3680 , n9722 , n3739 );
    and g8374 ( n8156 , n9360 , n7633 );
    and g8375 ( n2247 , n4859 , n2263 );
    xnor g8376 ( n7565 , n10615 , n4523 );
    and g8377 ( n9331 , n7872 , n9468 );
    or g8378 ( n2846 , n2099 , n4249 );
    and g8379 ( n2461 , n8737 , n5874 );
    xnor g8380 ( n12715 , n10866 , n8332 );
    not g8381 ( n10760 , n12360 );
    xnor g8382 ( n6330 , n12533 , n9996 );
    xnor g8383 ( n7556 , n1642 , n6707 );
    nor g8384 ( n3334 , n5301 , n8701 );
    xnor g8385 ( n1553 , n8390 , n757 );
    not g8386 ( n6636 , n11844 );
    and g8387 ( n4196 , n12146 , n10609 );
    xnor g8388 ( n1615 , n9130 , n9279 );
    or g8389 ( n10467 , n4628 , n12124 );
    xnor g8390 ( n10272 , n10769 , n2241 );
    or g8391 ( n7886 , n10108 , n11746 );
    xnor g8392 ( n3055 , n8111 , n9012 );
    xnor g8393 ( n10000 , n6466 , n6079 );
    not g8394 ( n12078 , n8913 );
    not g8395 ( n12442 , n10560 );
    or g8396 ( n348 , n5589 , n11291 );
    or g8397 ( n6766 , n12256 , n195 );
    xor g8398 ( n6406 , n2968 , n4306 );
    not g8399 ( n3540 , n382 );
    or g8400 ( n9913 , n636 , n6071 );
    and g8401 ( n5398 , n3389 , n10001 );
    or g8402 ( n11281 , n12119 , n12754 );
    or g8403 ( n7998 , n5575 , n11820 );
    and g8404 ( n12267 , n9705 , n971 );
    not g8405 ( n11410 , n10451 );
    xnor g8406 ( n5676 , n4500 , n3469 );
    xnor g8407 ( n10245 , n1331 , n12919 );
    xnor g8408 ( n4020 , n8920 , n295 );
    xnor g8409 ( n12459 , n7176 , n506 );
    or g8410 ( n10156 , n7986 , n968 );
    xnor g8411 ( n234 , n8778 , n955 );
    not g8412 ( n8010 , n83 );
    xnor g8413 ( n4000 , n10808 , n2529 );
    and g8414 ( n2055 , n5876 , n5307 );
    xnor g8415 ( n10406 , n4387 , n4894 );
    nor g8416 ( n7689 , n84 , n9350 );
    xnor g8417 ( n5900 , n1364 , n1517 );
    xnor g8418 ( n9747 , n885 , n5836 );
    xnor g8419 ( n2028 , n7672 , n220 );
    or g8420 ( n792 , n7090 , n7255 );
    nor g8421 ( n7104 , n1863 , n11916 );
    xnor g8422 ( n8657 , n10143 , n909 );
    xnor g8423 ( n3879 , n5736 , n9955 );
    xnor g8424 ( n9493 , n7088 , n2926 );
    xnor g8425 ( n8076 , n7775 , n8490 );
    nor g8426 ( n12483 , n774 , n5608 );
    or g8427 ( n12599 , n9389 , n7246 );
    not g8428 ( n6607 , n12611 );
    and g8429 ( n2244 , n1144 , n5210 );
    not g8430 ( n4773 , n4390 );
    and g8431 ( n12766 , n7169 , n1238 );
    or g8432 ( n1026 , n1215 , n5055 );
    not g8433 ( n11599 , n12893 );
    or g8434 ( n2040 , n6073 , n8947 );
    or g8435 ( n894 , n7449 , n9160 );
    xnor g8436 ( n4680 , n7355 , n5444 );
    nor g8437 ( n12233 , n324 , n5686 );
    or g8438 ( n6606 , n12361 , n8414 );
    or g8439 ( n3277 , n11241 , n7689 );
    and g8440 ( n2824 , n4805 , n5645 );
    xnor g8441 ( n6517 , n11268 , n3525 );
    xnor g8442 ( n6443 , n4570 , n9874 );
    and g8443 ( n9593 , n6231 , n3444 );
    not g8444 ( n4835 , n7784 );
    nor g8445 ( n174 , n6575 , n9458 );
    or g8446 ( n12146 , n1803 , n6421 );
    or g8447 ( n2424 , n12119 , n7382 );
    xnor g8448 ( n5315 , n1315 , n2211 );
    xnor g8449 ( n12838 , n7112 , n12654 );
    or g8450 ( n6564 , n3743 , n8745 );
    xnor g8451 ( n7936 , n4409 , n11220 );
    or g8452 ( n10458 , n994 , n11746 );
    and g8453 ( n1563 , n9519 , n9023 );
    or g8454 ( n2453 , n4737 , n5932 );
    xnor g8455 ( n1698 , n1653 , n10896 );
    and g8456 ( n11363 , n2072 , n3908 );
    not g8457 ( n10426 , n12452 );
    or g8458 ( n9476 , n10879 , n6389 );
    and g8459 ( n8380 , n4697 , n6968 );
    or g8460 ( n5032 , n6418 , n729 );
    nor g8461 ( n1711 , n11056 , n1535 );
    nor g8462 ( n10999 , n5194 , n8710 );
    not g8463 ( n11843 , n12052 );
    or g8464 ( n804 , n1937 , n10903 );
    and g8465 ( n4463 , n5964 , n9956 );
    or g8466 ( n9780 , n3995 , n482 );
    not g8467 ( n8523 , n5353 );
    not g8468 ( n1455 , n9956 );
    not g8469 ( n4456 , n758 );
    and g8470 ( n5754 , n6307 , n4636 );
    nor g8471 ( n9324 , n11836 , n12286 );
    xnor g8472 ( n1390 , n10307 , n999 );
    and g8473 ( n1235 , n4892 , n583 );
    xnor g8474 ( n11108 , n2640 , n12181 );
    xnor g8475 ( n7878 , n7130 , n11464 );
    or g8476 ( n8325 , n3820 , n8830 );
    xnor g8477 ( n5648 , n386 , n9354 );
    or g8478 ( n386 , n8026 , n7952 );
    and g8479 ( n3646 , n1701 , n3338 );
    or g8480 ( n11431 , n9180 , n11564 );
    or g8481 ( n236 , n5530 , n6071 );
    xnor g8482 ( n5498 , n5608 , n774 );
    xnor g8483 ( n11915 , n2363 , n10097 );
    and g8484 ( n6408 , n9644 , n4925 );
    nor g8485 ( n10372 , n12737 , n1742 );
    xnor g8486 ( n946 , n4808 , n2166 );
    and g8487 ( n2851 , n5283 , n6254 );
    or g8488 ( n621 , n9878 , n8655 );
    and g8489 ( n4977 , n7203 , n3304 );
    and g8490 ( n83 , n6706 , n10702 );
    not g8491 ( n5506 , n11972 );
    xnor g8492 ( n8425 , n3203 , n9601 );
    nor g8493 ( n10543 , n3733 , n8200 );
    and g8494 ( n4947 , n12610 , n7794 );
    or g8495 ( n9328 , n10879 , n1851 );
    not g8496 ( n561 , n10327 );
    xnor g8497 ( n9116 , n1082 , n11336 );
    or g8498 ( n10206 , n12616 , n10627 );
    xnor g8499 ( n7981 , n11730 , n6215 );
    or g8500 ( n12362 , n636 , n8648 );
    xnor g8501 ( n844 , n2607 , n5472 );
    and g8502 ( n10584 , n5211 , n9287 );
    or g8503 ( n7434 , n2456 , n12446 );
    xnor g8504 ( n327 , n788 , n12009 );
    and g8505 ( n10334 , n12496 , n10286 );
    not g8506 ( n8454 , n10870 );
    xnor g8507 ( n292 , n433 , n11705 );
    xnor g8508 ( n658 , n10146 , n1522 );
    xnor g8509 ( n1248 , n5382 , n2905 );
    or g8510 ( n8066 , n4498 , n4400 );
    or g8511 ( n6470 , n5530 , n12735 );
    nor g8512 ( n5104 , n2922 , n5244 );
    xnor g8513 ( n1942 , n9124 , n11629 );
    xnor g8514 ( n6324 , n3145 , n1267 );
    not g8515 ( n114 , n12753 );
    not g8516 ( n9445 , n12562 );
    or g8517 ( n2907 , n12061 , n10900 );
    xnor g8518 ( n5849 , n7762 , n1213 );
    nor g8519 ( n10405 , n643 , n11979 );
    or g8520 ( n11579 , n2313 , n2669 );
    xnor g8521 ( n5578 , n5021 , n1414 );
    or g8522 ( n10660 , n3947 , n172 );
    xnor g8523 ( n9041 , n891 , n4598 );
    or g8524 ( n1839 , n11245 , n2673 );
    or g8525 ( n1776 , n9370 , n7703 );
    or g8526 ( n12470 , n1941 , n10903 );
    or g8527 ( n8880 , n10139 , n3615 );
    not g8528 ( n7714 , n8160 );
    or g8529 ( n10731 , n7337 , n3400 );
    and g8530 ( n12569 , n9365 , n3307 );
    or g8531 ( n439 , n596 , n5716 );
    and g8532 ( n9551 , n5503 , n730 );
    xnor g8533 ( n7644 , n5214 , n2616 );
    and g8534 ( n3852 , n4203 , n7354 );
    not g8535 ( n5468 , n2498 );
    or g8536 ( n7562 , n6003 , n11614 );
    or g8537 ( n4940 , n6385 , n8468 );
    or g8538 ( n10030 , n9112 , n8186 );
    not g8539 ( n11472 , n7531 );
    and g8540 ( n12422 , n1082 , n919 );
    xnor g8541 ( n11600 , n1662 , n6713 );
    xnor g8542 ( n433 , n5217 , n9200 );
    xnor g8543 ( n932 , n5039 , n12358 );
    xnor g8544 ( n2688 , n11714 , n4251 );
    xor g8545 ( n11831 , n6101 , n2023 );
    or g8546 ( n11569 , n7391 , n1455 );
    xnor g8547 ( n7472 , n6584 , n12702 );
    xnor g8548 ( n11427 , n5685 , n5658 );
    xnor g8549 ( n7838 , n5761 , n5831 );
    not g8550 ( n5199 , n2436 );
    xnor g8551 ( n8457 , n161 , n550 );
    xnor g8552 ( n6891 , n12362 , n9811 );
    or g8553 ( n7409 , n1699 , n3224 );
    xnor g8554 ( n11550 , n6060 , n299 );
    xnor g8555 ( n12609 , n11633 , n9647 );
    not g8556 ( n5738 , n8906 );
    and g8557 ( n3970 , n5462 , n4080 );
    xnor g8558 ( n7923 , n9698 , n12540 );
    or g8559 ( n12742 , n5530 , n8644 );
    and g8560 ( n9311 , n3992 , n159 );
    nor g8561 ( n9002 , n5899 , n2928 );
    not g8562 ( n2935 , n2943 );
    xnor g8563 ( n6061 , n1750 , n2500 );
    and g8564 ( n4877 , n4872 , n12374 );
    and g8565 ( n12773 , n947 , n6533 );
    xnor g8566 ( n2416 , n2933 , n9760 );
    xnor g8567 ( n12428 , n1309 , n9602 );
    or g8568 ( n9357 , n11626 , n12763 );
    and g8569 ( n10979 , n12495 , n4729 );
    xnor g8570 ( n7761 , n5525 , n5552 );
    or g8571 ( n7458 , n5945 , n12816 );
    or g8572 ( n1548 , n5355 , n3911 );
    or g8573 ( n11710 , n807 , n1413 );
    and g8574 ( n12099 , n3872 , n2814 );
    not g8575 ( n11980 , n4314 );
    xnor g8576 ( n3547 , n3790 , n4106 );
    and g8577 ( n1412 , n6091 , n6855 );
    xnor g8578 ( n11094 , n10493 , n9947 );
    xnor g8579 ( n4616 , n9943 , n4488 );
    and g8580 ( n5701 , n9190 , n8079 );
    or g8581 ( n7250 , n6525 , n2860 );
    or g8582 ( n9182 , n1990 , n7635 );
    not g8583 ( n11168 , n3401 );
    or g8584 ( n8343 , n9373 , n1476 );
    nor g8585 ( n12732 , n8594 , n10081 );
    or g8586 ( n9846 , n5355 , n8735 );
    or g8587 ( n12302 , n7709 , n4474 );
    and g8588 ( n9499 , n6876 , n6818 );
    or g8589 ( n6515 , n8187 , n510 );
    or g8590 ( n12284 , n2099 , n10422 );
    and g8591 ( n11933 , n3974 , n2041 );
    nor g8592 ( n7817 , n3210 , n10527 );
    or g8593 ( n11846 , n7449 , n9568 );
    and g8594 ( n10194 , n910 , n9852 );
    or g8595 ( n4225 , n9002 , n2114 );
    xnor g8596 ( n2383 , n8811 , n9774 );
    not g8597 ( n3735 , n8235 );
    or g8598 ( n12462 , n4911 , n1546 );
    nor g8599 ( n7065 , n1878 , n11494 );
    or g8600 ( n6196 , n12447 , n4665 );
    and g8601 ( n6706 , n5331 , n12489 );
    and g8602 ( n1265 , n10542 , n5178 );
    not g8603 ( n11519 , n12505 );
    xnor g8604 ( n12108 , n2482 , n2163 );
    or g8605 ( n6313 , n11808 , n1838 );
    not g8606 ( n6154 , n12448 );
    or g8607 ( n1215 , n9389 , n1851 );
    nor g8608 ( n9789 , n12368 , n7583 );
    not g8609 ( n6969 , n11173 );
    and g8610 ( n12404 , n11375 , n6144 );
    not g8611 ( n3813 , n233 );
    xnor g8612 ( n8862 , n4002 , n6061 );
    xnor g8613 ( n2385 , n613 , n836 );
    xnor g8614 ( n11545 , n5164 , n513 );
    nor g8615 ( n8166 , n434 , n11871 );
    or g8616 ( n10532 , n5724 , n8890 );
    or g8617 ( n11842 , n5530 , n10854 );
    or g8618 ( n3940 , n12289 , n9253 );
    not g8619 ( n4493 , n3852 );
    or g8620 ( n10474 , n9803 , n6160 );
    or g8621 ( n2697 , n2761 , n6288 );
    not g8622 ( n3690 , n12480 );
    or g8623 ( n10102 , n6249 , n251 );
    and g8624 ( n2350 , n9208 , n12696 );
    not g8625 ( n7659 , n10450 );
    not g8626 ( n11793 , n10845 );
    xnor g8627 ( n9790 , n11335 , n12278 );
    not g8628 ( n732 , n49 );
    and g8629 ( n1192 , n12661 , n2753 );
    not g8630 ( n3590 , n6974 );
    xnor g8631 ( n7751 , n3176 , n10322 );
    xnor g8632 ( n152 , n7446 , n1023 );
    or g8633 ( n12118 , n5915 , n12735 );
    xnor g8634 ( n11784 , n11482 , n10635 );
    nor g8635 ( n7045 , n12607 , n10204 );
    or g8636 ( n515 , n4628 , n4818 );
    or g8637 ( n8963 , n6577 , n7425 );
    or g8638 ( n10169 , n10835 , n12120 );
    or g8639 ( n6275 , n8103 , n5741 );
    xnor g8640 ( n6647 , n8550 , n10934 );
    and g8641 ( n4744 , n11189 , n7922 );
    not g8642 ( n2538 , n12122 );
    xnor g8643 ( n6731 , n7059 , n3835 );
    not g8644 ( n734 , n10972 );
    and g8645 ( n7682 , n3188 , n689 );
    not g8646 ( n8944 , n3904 );
    not g8647 ( n12577 , n1275 );
    or g8648 ( n7790 , n2217 , n2020 );
    xnor g8649 ( n1692 , n6231 , n12103 );
    xnor g8650 ( n5120 , n10773 , n490 );
    xnor g8651 ( n12828 , n3795 , n8868 );
    xnor g8652 ( n2834 , n6539 , n47 );
    xnor g8653 ( n12420 , n3301 , n691 );
    xnor g8654 ( n7784 , n12933 , n8989 );
    xnor g8655 ( n6503 , n3544 , n3414 );
    not g8656 ( n10337 , n1124 );
    or g8657 ( n11539 , n5231 , n5217 );
    xnor g8658 ( n9865 , n8869 , n12806 );
    not g8659 ( n12614 , n2305 );
    xnor g8660 ( n12627 , n2005 , n3331 );
    or g8661 ( n11171 , n3096 , n7425 );
    and g8662 ( n3495 , n693 , n3069 );
    and g8663 ( n3439 , n240 , n983 );
    or g8664 ( n3780 , n9098 , n2812 );
    xnor g8665 ( n3914 , n9198 , n8640 );
    xnor g8666 ( n4917 , n9479 , n12515 );
    or g8667 ( n3906 , n191 , n5851 );
    xnor g8668 ( n4139 , n9042 , n11399 );
    or g8669 ( n4637 , n5225 , n1625 );
    or g8670 ( n4201 , n12284 , n663 );
    not g8671 ( n685 , n6002 );
    and g8672 ( n5659 , n11060 , n11247 );
    xnor g8673 ( n9075 , n11842 , n7027 );
    and g8674 ( n12461 , n148 , n3927 );
    xnor g8675 ( n2467 , n772 , n2645 );
    nor g8676 ( n6870 , n6800 , n8436 );
    and g8677 ( n393 , n719 , n6314 );
    nor g8678 ( n10129 , n8015 , n12716 );
    xnor g8679 ( n6435 , n2136 , n10652 );
    nor g8680 ( n12800 , n8444 , n6693 );
    xnor g8681 ( n6545 , n6805 , n869 );
    xnor g8682 ( n5615 , n7122 , n746 );
    or g8683 ( n3980 , n1126 , n4143 );
    nor g8684 ( n5118 , n11240 , n3993 );
    and g8685 ( n6260 , n10829 , n3589 );
    or g8686 ( n3523 , n10835 , n3599 );
    xnor g8687 ( n4385 , n6939 , n208 );
    xnor g8688 ( n10676 , n203 , n8447 );
    xnor g8689 ( n531 , n6453 , n7412 );
    not g8690 ( n120 , n8093 );
    xnor g8691 ( n7907 , n7567 , n11794 );
    and g8692 ( n604 , n19 , n4533 );
    and g8693 ( n11145 , n2014 , n9821 );
    or g8694 ( n11601 , n4223 , n1819 );
    and g8695 ( n2760 , n8459 , n11573 );
    or g8696 ( n4644 , n3743 , n4875 );
    not g8697 ( n10098 , n12047 );
    xnor g8698 ( n7467 , n6318 , n7064 );
    nor g8699 ( n4982 , n11514 , n3012 );
    or g8700 ( n9198 , n12485 , n7670 );
    xnor g8701 ( n6554 , n8231 , n11135 );
    and g8702 ( n945 , n11195 , n9292 );
    or g8703 ( n8317 , n9584 , n2020 );
    or g8704 ( n3256 , n4846 , n11562 );
    not g8705 ( n4736 , n578 );
    xnor g8706 ( n11408 , n12524 , n2088 );
    xnor g8707 ( n9542 , n12309 , n10651 );
    and g8708 ( n10511 , n2170 , n1897 );
    or g8709 ( n5712 , n11433 , n9741 );
    xnor g8710 ( n672 , n1346 , n5163 );
    or g8711 ( n9940 , n10879 , n1162 );
    xnor g8712 ( n11559 , n10693 , n8709 );
    xnor g8713 ( n11929 , n9897 , n979 );
    nor g8714 ( n11476 , n9486 , n1264 );
    or g8715 ( n8449 , n8026 , n8768 );
    xnor g8716 ( n10959 , n7075 , n4746 );
    xnor g8717 ( n6713 , n5205 , n3949 );
    or g8718 ( n6599 , n9389 , n1546 );
    or g8719 ( n1878 , n11560 , n9658 );
    and g8720 ( n12528 , n5516 , n6719 );
    xnor g8721 ( n7978 , n3283 , n2849 );
    nor g8722 ( n6125 , n709 , n1568 );
    or g8723 ( n2374 , n2832 , n5497 );
    or g8724 ( n12668 , n7449 , n5914 );
    and g8725 ( n9102 , n7690 , n2558 );
    nor g8726 ( n6397 , n1028 , n5924 );
    and g8727 ( n7345 , n8256 , n2373 );
    xnor g8728 ( n11798 , n11669 , n652 );
    xnor g8729 ( n8436 , n5532 , n8501 );
    xnor g8730 ( n8647 , n11514 , n7727 );
    or g8731 ( n10144 , n12853 , n12535 );
    or g8732 ( n9990 , n1475 , n4986 );
    xnor g8733 ( n5094 , n11491 , n12222 );
    or g8734 ( n8294 , n11958 , n184 );
    or g8735 ( n4132 , n6134 , n12401 );
    nor g8736 ( n6685 , n3354 , n7607 );
    not g8737 ( n7841 , n7631 );
    or g8738 ( n5824 , n12864 , n9456 );
    and g8739 ( n3524 , n11968 , n6 );
    or g8740 ( n7200 , n989 , n12328 );
    and g8741 ( n12727 , n10398 , n1601 );
    xnor g8742 ( n11636 , n722 , n10325 );
    xnor g8743 ( n10556 , n5079 , n10084 );
    or g8744 ( n11598 , n7449 , n28 );
    and g8745 ( n4028 , n2464 , n5105 );
    and g8746 ( n2839 , n6782 , n7054 );
    not g8747 ( n9815 , n820 );
    xnor g8748 ( n4507 , n688 , n7853 );
    xnor g8749 ( n6253 , n4907 , n8766 );
    and g8750 ( n581 , n10945 , n7318 );
    and g8751 ( n9909 , n9382 , n3760 );
    or g8752 ( n9307 , n752 , n6169 );
    or g8753 ( n10847 , n5355 , n1079 );
    and g8754 ( n1324 , n8476 , n1564 );
    nor g8755 ( n4889 , n6861 , n10985 );
    and g8756 ( n4804 , n9313 , n190 );
    xor g8757 ( n4397 , n165 , n6990 );
    or g8758 ( n9266 , n4628 , n12080 );
    xnor g8759 ( n12215 , n12603 , n8696 );
    or g8760 ( n1677 , n8996 , n9518 );
    xnor g8761 ( n923 , n11800 , n7358 );
    or g8762 ( n3279 , n12365 , n11406 );
    not g8763 ( n3599 , n1906 );
    or g8764 ( n11402 , n11493 , n8122 );
    xnor g8765 ( n1589 , n9391 , n5302 );
    xnor g8766 ( n7194 , n9114 , n11581 );
    xnor g8767 ( n8245 , n1205 , n5617 );
    and g8768 ( n10284 , n11740 , n4969 );
    xnor g8769 ( n5730 , n3202 , n8683 );
    xnor g8770 ( n8598 , n2440 , n9261 );
    and g8771 ( n11310 , n3243 , n5880 );
    and g8772 ( n10963 , n1282 , n12458 );
    xnor g8773 ( n1586 , n8840 , n11315 );
    or g8774 ( n7884 , n6656 , n9548 );
    and g8775 ( n3504 , n7398 , n12219 );
    or g8776 ( n12246 , n8738 , n9160 );
    nor g8777 ( n2212 , n10112 , n12547 );
    not g8778 ( n11746 , n3932 );
    not g8779 ( n2171 , n8521 );
    xnor g8780 ( n9001 , n418 , n207 );
    nor g8781 ( n11808 , n6954 , n4912 );
    and g8782 ( n9261 , n12194 , n2351 );
    or g8783 ( n5650 , n10835 , n6138 );
    xnor g8784 ( n7387 , n8737 , n6644 );
    or g8785 ( n6522 , n6271 , n11420 );
    or g8786 ( n5387 , n5858 , n4400 );
    and g8787 ( n10211 , n10387 , n3019 );
    and g8788 ( n10756 , n2010 , n2261 );
    xnor g8789 ( n9929 , n3694 , n1849 );
    xnor g8790 ( n7815 , n12071 , n11230 );
    xnor g8791 ( n9257 , n12177 , n2430 );
    not g8792 ( n8592 , n6584 );
    not g8793 ( n6490 , n5093 );
    or g8794 ( n1095 , n12701 , n6897 );
    and g8795 ( n10208 , n11547 , n6832 );
    and g8796 ( n8910 , n6686 , n5407 );
    and g8797 ( n2118 , n11162 , n1302 );
    and g8798 ( n9403 , n11936 , n3346 );
    and g8799 ( n8281 , n11478 , n1564 );
    and g8800 ( n1109 , n9266 , n8711 );
    and g8801 ( n8233 , n2319 , n10252 );
    and g8802 ( n12166 , n4950 , n2596 );
    xnor g8803 ( n11872 , n8892 , n8906 );
    not g8804 ( n7673 , n9348 );
    xor g8805 ( n6587 , n4741 , n7253 );
    and g8806 ( n1147 , n12438 , n8185 );
    xnor g8807 ( n10989 , n10880 , n7361 );
    xnor g8808 ( n12519 , n7248 , n12159 );
    xor g8809 ( n3134 , n8516 , n4682 );
    and g8810 ( n2571 , n7166 , n11163 );
    or g8811 ( n5422 , n8010 , n12089 );
    not g8812 ( n7607 , n4427 );
    or g8813 ( n413 , n3381 , n10811 );
    not g8814 ( n12427 , n10802 );
    and g8815 ( n3643 , n8816 , n1084 );
    or g8816 ( n12142 , n2456 , n7382 );
    or g8817 ( n3508 , n5575 , n2589 );
    or g8818 ( n1174 , n8959 , n5012 );
    xnor g8819 ( n7507 , n8389 , n10747 );
    xnor g8820 ( n5628 , n6008 , n4581 );
    or g8821 ( n677 , n7452 , n8615 );
    and g8822 ( n12729 , n443 , n10200 );
    and g8823 ( n10508 , n7911 , n5323 );
    nor g8824 ( n3860 , n23 , n7844 );
    xnor g8825 ( n8591 , n1438 , n6778 );
    or g8826 ( n3843 , n114 , n5012 );
    nor g8827 ( n5375 , n7230 , n11019 );
    and g8828 ( n4092 , n10354 , n1502 );
    or g8829 ( n3520 , n12853 , n5468 );
    or g8830 ( n9164 , n4778 , n5468 );
    or g8831 ( n6844 , n11887 , n10854 );
    not g8832 ( n673 , n1317 );
    and g8833 ( n8937 , n12220 , n6388 );
    or g8834 ( n4346 , n1941 , n6197 );
    or g8835 ( n1444 , n11851 , n9255 );
    not g8836 ( n11346 , n12355 );
    nor g8837 ( n5097 , n2411 , n8486 );
    not g8838 ( n11759 , n4930 );
    or g8839 ( n7590 , n6971 , n7178 );
    xnor g8840 ( n8872 , n6581 , n12820 );
    xnor g8841 ( n9663 , n11988 , n2374 );
    nor g8842 ( n1797 , n8938 , n578 );
    and g8843 ( n7423 , n4457 , n622 );
    not g8844 ( n8921 , n2760 );
    xnor g8845 ( n5894 , n3481 , n575 );
    not g8846 ( n4611 , n6838 );
    or g8847 ( n1012 , n191 , n6402 );
    xnor g8848 ( n12923 , n2019 , n462 );
    xnor g8849 ( n193 , n8452 , n8978 );
    or g8850 ( n4219 , n1449 , n1174 );
    xnor g8851 ( n5184 , n11442 , n728 );
    or g8852 ( n7325 , n9373 , n9078 );
    nor g8853 ( n11995 , n6594 , n6670 );
    xnor g8854 ( n1411 , n1924 , n10014 );
    xnor g8855 ( n5075 , n9718 , n3738 );
    xnor g8856 ( n7559 , n7325 , n8325 );
    and g8857 ( n11671 , n3594 , n7156 );
    xnor g8858 ( n7016 , n3483 , n12894 );
    and g8859 ( n10659 , n9421 , n1885 );
    or g8860 ( n437 , n10429 , n7158 );
    and g8861 ( n1802 , n10064 , n10905 );
    or g8862 ( n7445 , n7537 , n4803 );
    and g8863 ( n2421 , n5800 , n738 );
    xnor g8864 ( n10227 , n12198 , n4024 );
    or g8865 ( n5570 , n8428 , n11122 );
    not g8866 ( n8740 , n1067 );
    or g8867 ( n11714 , n8870 , n12535 );
    or g8868 ( n6738 , n9389 , n7424 );
    or g8869 ( n3065 , n5809 , n3924 );
    xnor g8870 ( n11755 , n5327 , n11912 );
    xnor g8871 ( n6494 , n12895 , n1834 );
    or g8872 ( n1882 , n3717 , n1894 );
    not g8873 ( n4764 , n9072 );
    xnor g8874 ( n703 , n5049 , n958 );
    xnor g8875 ( n11315 , n3346 , n3242 );
    or g8876 ( n6072 , n6718 , n9568 );
    or g8877 ( n1740 , n8428 , n6114 );
    and g8878 ( n12141 , n10512 , n2742 );
    not g8879 ( n10986 , n9805 );
    or g8880 ( n9939 , n6136 , n5835 );
    xnor g8881 ( n4326 , n5978 , n10597 );
    or g8882 ( n7809 , n3628 , n894 );
    and g8883 ( n3782 , n2608 , n4615 );
    xnor g8884 ( n12383 , n9258 , n2584 );
    xnor g8885 ( n12615 , n11490 , n10318 );
    not g8886 ( n6493 , n9467 );
    not g8887 ( n12080 , n5579 );
    not g8888 ( n10330 , n1984 );
    xnor g8889 ( n9508 , n11208 , n1911 );
    and g8890 ( n8532 , n1371 , n6392 );
    xnor g8891 ( n10061 , n11955 , n1819 );
    not g8892 ( n4242 , n4370 );
    not g8893 ( n7398 , n7206 );
    or g8894 ( n4195 , n12186 , n6455 );
    or g8895 ( n11563 , n10835 , n4654 );
    not g8896 ( n362 , n3715 );
    nor g8897 ( n754 , n10582 , n6998 );
    and g8898 ( n1837 , n7773 , n1633 );
    xnor g8899 ( n6754 , n3711 , n912 );
    and g8900 ( n12875 , n3240 , n8801 );
    or g8901 ( n11221 , n10142 , n7424 );
    xnor g8902 ( n4156 , n1021 , n3502 );
    xnor g8903 ( n6555 , n1258 , n7250 );
    and g8904 ( n12266 , n9739 , n7224 );
    or g8905 ( n10725 , n9266 , n8711 );
    or g8906 ( n1806 , n7839 , n5012 );
    not g8907 ( n1796 , n6370 );
    not g8908 ( n11863 , n12292 );
    xnor g8909 ( n2869 , n11575 , n9057 );
    or g8910 ( n1783 , n12891 , n11506 );
    or g8911 ( n2763 , n5355 , n1851 );
    not g8912 ( n5311 , n783 );
    not g8913 ( n11857 , n11271 );
    or g8914 ( n271 , n9389 , n12843 );
    or g8915 ( n8055 , n191 , n10419 );
    or g8916 ( n3180 , n10879 , n7341 );
    and g8917 ( n11787 , n12525 , n3298 );
    and g8918 ( n4851 , n8327 , n2701 );
    and g8919 ( n9454 , n4600 , n410 );
    or g8920 ( n5397 , n5809 , n6513 );
    and g8921 ( n10047 , n8720 , n12064 );
    xnor g8922 ( n10126 , n7653 , n4688 );
    or g8923 ( n12661 , n914 , n2429 );
    xnor g8924 ( n12951 , n2539 , n5910 );
    and g8925 ( n4953 , n5305 , n5212 );
    and g8926 ( n6007 , n12051 , n3091 );
    or g8927 ( n10899 , n5501 , n4792 );
    or g8928 ( n3422 , n12070 , n2621 );
    or g8929 ( n1988 , n6158 , n3052 );
    and g8930 ( n3896 , n9081 , n6258 );
    or g8931 ( n998 , n11324 , n12756 );
    xnor g8932 ( n11372 , n7793 , n536 );
    or g8933 ( n12840 , n7865 , n12338 );
    nor g8934 ( n319 , n9455 , n513 );
    xnor g8935 ( n7990 , n2058 , n4218 );
    and g8936 ( n7699 , n12063 , n12149 );
    xnor g8937 ( n10328 , n1810 , n7990 );
    xnor g8938 ( n6996 , n10404 , n1132 );
    xnor g8939 ( n2588 , n9270 , n6356 );
    and g8940 ( n1524 , n1516 , n2189 );
    xnor g8941 ( n4090 , n1371 , n690 );
    not g8942 ( n10629 , n6760 );
    not g8943 ( n10316 , n3094 );
    or g8944 ( n6695 , n3746 , n5012 );
    and g8945 ( n9757 , n12936 , n6796 );
    xnor g8946 ( n1603 , n9492 , n4546 );
    not g8947 ( n6999 , n9167 );
    not g8948 ( n9709 , n2089 );
    xnor g8949 ( n6056 , n1947 , n3151 );
    or g8950 ( n12716 , n10093 , n12105 );
    nor g8951 ( n4840 , n12198 , n1562 );
    or g8952 ( n2324 , n6767 , n6250 );
    nor g8953 ( n7744 , n6853 , n5076 );
    xnor g8954 ( n12482 , n9443 , n7377 );
    or g8955 ( n2626 , n8428 , n11820 );
    xnor g8956 ( n1864 , n5907 , n5343 );
    not g8957 ( n10070 , n10844 );
    or g8958 ( n4266 , n1549 , n10856 );
    xnor g8959 ( n9163 , n3135 , n11057 );
    xnor g8960 ( n8728 , n2071 , n10323 );
    or g8961 ( n12278 , n10157 , n7921 );
    and g8962 ( n12115 , n9707 , n6526 );
    or g8963 ( n11658 , n1779 , n4685 );
    xnor g8964 ( n4497 , n5661 , n7164 );
    and g8965 ( n390 , n10962 , n9333 );
    and g8966 ( n2178 , n1341 , n9522 );
    xnor g8967 ( n9809 , n11069 , n11128 );
    not g8968 ( n9505 , n1240 );
    or g8969 ( n12743 , n7709 , n4654 );
    or g8970 ( n1493 , n9370 , n2358 );
    nor g8971 ( n867 , n12269 , n7003 );
    not g8972 ( n3347 , n10648 );
    or g8973 ( n12045 , n8369 , n4108 );
    or g8974 ( n9518 , n1699 , n826 );
    xnor g8975 ( n793 , n935 , n606 );
    or g8976 ( n820 , n994 , n4400 );
    or g8977 ( n11778 , n4237 , n10229 );
    xnor g8978 ( n3167 , n11339 , n9224 );
    not g8979 ( n2067 , n20 );
    or g8980 ( n4255 , n9037 , n448 );
    or g8981 ( n11451 , n3820 , n3606 );
    nor g8982 ( n7594 , n7756 , n4681 );
    and g8983 ( n5205 , n8755 , n6648 );
    xnor g8984 ( n11921 , n12226 , n6340 );
    and g8985 ( n11365 , n11892 , n7294 );
    nor g8986 ( n2651 , n3353 , n5545 );
    and g8987 ( n1994 , n5964 , n1798 );
    xnor g8988 ( n10703 , n11704 , n2368 );
    not g8989 ( n9917 , n10488 );
    xnor g8990 ( n4743 , n8828 , n4123 );
    or g8991 ( n4261 , n4911 , n4242 );
    not g8992 ( n7356 , n3250 );
    or g8993 ( n7421 , n4360 , n8396 );
    and g8994 ( n7925 , n2186 , n12453 );
    xnor g8995 ( n10043 , n63 , n11595 );
    and g8996 ( n12681 , n3480 , n2611 );
    and g8997 ( n12756 , n1107 , n5287 );
    xnor g8998 ( n3288 , n3136 , n8886 );
    or g8999 ( n107 , n12119 , n12080 );
    and g9000 ( n7146 , n10520 , n543 );
    xnor g9001 ( n8775 , n7929 , n5588 );
    nor g9002 ( n10523 , n2934 , n2353 );
    or g9003 ( n4870 , n420 , n10308 );
    xnor g9004 ( n7763 , n11593 , n4128 );
    not g9005 ( n9484 , n12934 );
    nor g9006 ( n4419 , n7034 , n10058 );
    not g9007 ( n1079 , n10223 );
    and g9008 ( n2910 , n1465 , n6272 );
    xnor g9009 ( n12592 , n10231 , n993 );
    and g9010 ( n4257 , n1246 , n4355 );
    and g9011 ( n10920 , n7383 , n4893 );
    or g9012 ( n9068 , n5765 , n5759 );
    or g9013 ( n11717 , n6365 , n6285 );
    xnor g9014 ( n4655 , n9684 , n6936 );
    not g9015 ( n12437 , n3011 );
    or g9016 ( n9880 , n12208 , n10017 );
    or g9017 ( n12550 , n2456 , n12883 );
    and g9018 ( n12116 , n3984 , n3902 );
    or g9019 ( n8295 , n5915 , n1932 );
    not g9020 ( n3468 , n8717 );
    or g9021 ( n3890 , n6707 , n9870 );
    xnor g9022 ( n8104 , n7348 , n1806 );
    xnor g9023 ( n8833 , n2773 , n1718 );
    or g9024 ( n12178 , n7391 , n1546 );
    or g9025 ( n7871 , n3127 , n510 );
    not g9026 ( n2483 , n3742 );
    nor g9027 ( n8716 , n4804 , n9957 );
    xnor g9028 ( n1725 , n8903 , n5834 );
    not g9029 ( n1403 , n4734 );
    or g9030 ( n1800 , n8583 , n28 );
    xnor g9031 ( n12378 , n23 , n1830 );
    xnor g9032 ( n5668 , n3676 , n3173 );
    not g9033 ( n12929 , n38 );
    and g9034 ( n3664 , n11546 , n4638 );
    xnor g9035 ( n32 , n7559 , n4712 );
    or g9036 ( n6010 , n1406 , n12168 );
    xnor g9037 ( n2173 , n445 , n9866 );
    xnor g9038 ( n7836 , n1111 , n7959 );
    nor g9039 ( n4987 , n4976 , n5657 );
    not g9040 ( n1704 , n8270 );
    or g9041 ( n1149 , n11147 , n12290 );
    xnor g9042 ( n10889 , n9965 , n6803 );
    xnor g9043 ( n4683 , n21 , n3705 );
    and g9044 ( n7963 , n9600 , n7860 );
    and g9045 ( n6854 , n3837 , n9096 );
    and g9046 ( n7807 , n6770 , n4634 );
    nor g9047 ( n10536 , n8445 , n8754 );
    nor g9048 ( n1892 , n12770 , n8877 );
    xnor g9049 ( n3387 , n3215 , n567 );
    xnor g9050 ( n11707 , n6942 , n10303 );
    or g9051 ( n6569 , n7839 , n6455 );
    and g9052 ( n11491 , n8153 , n10266 );
    or g9053 ( n7574 , n3820 , n4642 );
    or g9054 ( n8229 , n10750 , n8655 );
    nor g9055 ( n7583 , n7764 , n6710 );
    and g9056 ( n10947 , n4312 , n4634 );
    or g9057 ( n3153 , n10750 , n4913 );
    not g9058 ( n8626 , n12794 );
    xnor g9059 ( n2541 , n298 , n4919 );
    xnor g9060 ( n10686 , n12506 , n2489 );
    nor g9061 ( n1774 , n9269 , n9169 );
    not g9062 ( n2974 , n10993 );
    or g9063 ( n5364 , n3617 , n3224 );
    or g9064 ( n10053 , n3667 , n5580 );
    not g9065 ( n6169 , n7354 );
    and g9066 ( n4796 , n6470 , n7392 );
    xnor g9067 ( n5898 , n5869 , n7231 );
    xnor g9068 ( n1363 , n6895 , n414 );
    or g9069 ( n9003 , n3818 , n10716 );
    xnor g9070 ( n6920 , n3268 , n1045 );
    or g9071 ( n3023 , n91 , n3162 );
    or g9072 ( n2847 , n630 , n12394 );
    not g9073 ( n3859 , n8573 );
    and g9074 ( n1505 , n10781 , n4941 );
    not g9075 ( n8803 , n8477 );
    xnor g9076 ( n10694 , n8161 , n8218 );
    xnor g9077 ( n1536 , n10984 , n11643 );
    xnor g9078 ( n5481 , n3984 , n3902 );
    or g9079 ( n3628 , n10835 , n9144 );
    not g9080 ( n10712 , n8605 );
    not g9081 ( n25 , n12201 );
    or g9082 ( n1533 , n4479 , n859 );
    not g9083 ( n3962 , n7309 );
    and g9084 ( n231 , n10049 , n1521 );
    or g9085 ( n12167 , n7283 , n4775 );
    or g9086 ( n1715 , n11026 , n795 );
    not g9087 ( n636 , n7891 );
    not g9088 ( n6596 , n2296 );
    nor g9089 ( n10577 , n5928 , n3511 );
    not g9090 ( n9233 , n3255 );
    xnor g9091 ( n12325 , n4696 , n416 );
    and g9092 ( n1815 , n9657 , n1807 );
    not g9093 ( n7124 , n3202 );
    or g9094 ( n124 , n10055 , n12613 );
    and g9095 ( n10602 , n2979 , n4298 );
    or g9096 ( n8475 , n752 , n7876 );
    and g9097 ( n11726 , n9179 , n9479 );
    or g9098 ( n10735 , n10142 , n1915 );
    or g9099 ( n2559 , n4193 , n12637 );
    and g9100 ( n9289 , n6797 , n5645 );
    and g9101 ( n11434 , n2677 , n9579 );
    xnor g9102 ( n12311 , n8036 , n10094 );
    and g9103 ( n10512 , n5305 , n2509 );
    or g9104 ( n9167 , n11923 , n8830 );
    or g9105 ( n3974 , n12775 , n12913 );
    or g9106 ( n4182 , n5858 , n11827 );
    or g9107 ( n2721 , n5575 , n12816 );
    and g9108 ( n8676 , n4741 , n4384 );
    and g9109 ( n4110 , n11597 , n9573 );
    xnor g9110 ( n7727 , n392 , n9940 );
    xnor g9111 ( n5723 , n9553 , n1771 );
    and g9112 ( n232 , n5848 , n3913 );
    xnor g9113 ( n3307 , n10473 , n10167 );
    or g9114 ( n2505 , n11013 , n1346 );
    xnor g9115 ( n6232 , n6053 , n2118 );
    xnor g9116 ( n11837 , n10562 , n8250 );
    xnor g9117 ( n8239 , n1363 , n6438 );
    and g9118 ( n8512 , n1026 , n11169 );
    or g9119 ( n2687 , n183 , n10638 );
    or g9120 ( n11826 , n2832 , n11746 );
    xnor g9121 ( n5669 , n7029 , n9249 );
    not g9122 ( n790 , n9038 );
    nor g9123 ( n5508 , n6384 , n12233 );
    not g9124 ( n6785 , n6148 );
    or g9125 ( n12701 , n6373 , n4527 );
    xnor g9126 ( n1108 , n12668 , n10462 );
    not g9127 ( n10027 , n1440 );
    not g9128 ( n11233 , n7057 );
    xnor g9129 ( n6099 , n3659 , n11250 );
    or g9130 ( n12376 , n8954 , n10870 );
    nor g9131 ( n1127 , n4202 , n9496 );
    not g9132 ( n10294 , n8868 );
    and g9133 ( n12081 , n9106 , n1488 );
    xnor g9134 ( n8086 , n1024 , n7498 );
    or g9135 ( n1 , n2346 , n6228 );
    xnor g9136 ( n8465 , n8181 , n8485 );
    xnor g9137 ( n10503 , n6534 , n10826 );
    xnor g9138 ( n7179 , n2089 , n2015 );
    xnor g9139 ( n10416 , n2199 , n10954 );
    nor g9140 ( n11572 , n3921 , n3199 );
    and g9141 ( n2924 , n8476 , n6016 );
    xnor g9142 ( n9912 , n5274 , n2418 );
    xnor g9143 ( n10815 , n4205 , n8931 );
    and g9144 ( n4767 , n8117 , n745 );
    nor g9145 ( n9213 , n2144 , n2392 );
    xnor g9146 ( n4208 , n2479 , n8144 );
    or g9147 ( n12107 , n12186 , n12816 );
    or g9148 ( n10516 , n6577 , n10919 );
    or g9149 ( n427 , n4338 , n10237 );
    xnor g9150 ( n11912 , n10378 , n7279 );
    or g9151 ( n8996 , n12119 , n3924 );
    not g9152 ( n5809 , n10545 );
    not g9153 ( n8738 , n3986 );
    or g9154 ( n8810 , n5765 , n4875 );
    and g9155 ( n5146 , n3328 , n10633 );
    or g9156 ( n3358 , n10637 , n3057 );
    xnor g9157 ( n9760 , n8416 , n5562 );
    xnor g9158 ( n12861 , n7521 , n4244 );
    and g9159 ( n7505 , n12312 , n7063 );
    xnor g9160 ( n84 , n6535 , n1482 );
    not g9161 ( n10077 , n3772 );
    and g9162 ( n1447 , n4301 , n2204 );
    or g9163 ( n12708 , n5383 , n10553 );
    or g9164 ( n3909 , n11401 , n2666 );
    and g9165 ( n578 , n11539 , n7445 );
    and g9166 ( n5976 , n10095 , n6546 );
    nor g9167 ( n11046 , n6064 , n7069 );
    or g9168 ( n8748 , n10365 , n10723 );
    or g9169 ( n602 , n752 , n8414 );
    and g9170 ( n2019 , n10162 , n1558 );
    or g9171 ( n12189 , n12503 , n9568 );
    xnor g9172 ( n8013 , n4373 , n5628 );
    or g9173 ( n11331 , n2473 , n7782 );
    and g9174 ( n4652 , n3072 , n8111 );
    xnor g9175 ( n29 , n7490 , n10974 );
    or g9176 ( n4443 , n8964 , n5839 );
    xnor g9177 ( n6343 , n3726 , n277 );
    nor g9178 ( n8902 , n2962 , n6955 );
    or g9179 ( n3625 , n3743 , n10916 );
    or g9180 ( n11490 , n10835 , n11698 );
    or g9181 ( n6104 , n2656 , n5536 );
    not g9182 ( n5671 , n11178 );
    or g9183 ( n648 , n11712 , n9574 );
    nor g9184 ( n2674 , n6041 , n6923 );
    not g9185 ( n1738 , n9637 );
    or g9186 ( n4121 , n2456 , n5326 );
    and g9187 ( n8793 , n3261 , n11673 );
    xnor g9188 ( n7083 , n5652 , n12768 );
    and g9189 ( n720 , n5452 , n6117 );
    nor g9190 ( n3317 , n11250 , n5379 );
    or g9191 ( n705 , n2217 , n7506 );
    xnor g9192 ( n5776 , n8133 , n10317 );
    and g9193 ( n3600 , n2001 , n8698 );
    or g9194 ( n10343 , n5530 , n12754 );
    or g9195 ( n2657 , n6186 , n4998 );
    not g9196 ( n7709 , n9457 );
    xnor g9197 ( n2418 , n3314 , n915 );
    or g9198 ( n4760 , n4366 , n10752 );
    xnor g9199 ( n7355 , n361 , n7728 );
    or g9200 ( n2981 , n7283 , n561 );
    or g9201 ( n12065 , n4498 , n1546 );
    not g9202 ( n609 , n5153 );
    not g9203 ( n6928 , n2141 );
    xnor g9204 ( n9666 , n2608 , n4615 );
    and g9205 ( n1935 , n2893 , n1014 );
    and g9206 ( n7835 , n4808 , n5388 );
    nor g9207 ( n9580 , n7311 , n2344 );
    and g9208 ( n2919 , n9058 , n4197 );
    or g9209 ( n7203 , n6270 , n3877 );
    or g9210 ( n11112 , n4059 , n4400 );
    or g9211 ( n8051 , n1685 , n11030 );
    or g9212 ( n6774 , n4674 , n3224 );
    and g9213 ( n9416 , n4702 , n3750 );
    or g9214 ( n296 , n12503 , n3606 );
    or g9215 ( n8175 , n6373 , n9144 );
    nor g9216 ( n1170 , n895 , n290 );
    or g9217 ( n12194 , n7185 , n2895 );
    or g9218 ( n10777 , n4628 , n10422 );
    not g9219 ( n9225 , n7976 );
    xnor g9220 ( n4495 , n5650 , n11675 );
    and g9221 ( n9707 , n8241 , n8962 );
    not g9222 ( n1997 , n12163 );
    and g9223 ( n11038 , n9920 , n3932 );
    and g9224 ( n3886 , n8216 , n10480 );
    and g9225 ( n12315 , n12163 , n8684 );
    or g9226 ( n5265 , n9734 , n900 );
    or g9227 ( n3141 , n8026 , n11820 );
    not g9228 ( n1058 , n2918 );
    xnor g9229 ( n459 , n1495 , n1506 );
    or g9230 ( n6540 , n3310 , n2706 );
    or g9231 ( n2923 , n10434 , n9894 );
    not g9232 ( n5210 , n7499 );
    xnor g9233 ( n9904 , n5690 , n1607 );
    nor g9234 ( n12565 , n6356 , n9270 );
    xnor g9235 ( n3044 , n9398 , n446 );
    xnor g9236 ( n1159 , n2583 , n954 );
    or g9237 ( n6643 , n8428 , n10919 );
    or g9238 ( n4483 , n4628 , n8740 );
    not g9239 ( n9262 , n4722 );
    xnor g9240 ( n4861 , n6283 , n5838 );
    or g9241 ( n6242 , n8552 , n12735 );
    or g9242 ( n550 , n8428 , n6084 );
    and g9243 ( n920 , n2056 , n10008 );
    xnor g9244 ( n4430 , n9267 , n9044 );
    or g9245 ( n12750 , n8070 , n473 );
    and g9246 ( n8415 , n8920 , n8547 );
    or g9247 ( n8323 , n936 , n5520 );
    xnor g9248 ( n9300 , n4852 , n7868 );
    or g9249 ( n50 , n9389 , n4775 );
    xnor g9250 ( n9137 , n12081 , n153 );
    or g9251 ( n6514 , n962 , n9144 );
    nor g9252 ( n10006 , n4084 , n2120 );
    or g9253 ( n2976 , n10142 , n1079 );
    or g9254 ( n12063 , n2838 , n6164 );
    nor g9255 ( n11240 , n9647 , n11633 );
    or g9256 ( n10832 , n8458 , n3761 );
    nor g9257 ( n1635 , n7275 , n3788 );
    not g9258 ( n2718 , n1548 );
    and g9259 ( n2047 , n5082 , n8365 );
    or g9260 ( n11285 , n8959 , n6455 );
    not g9261 ( n3425 , n8776 );
    nor g9262 ( n3889 , n11507 , n3685 );
    or g9263 ( n12121 , n6940 , n7615 );
    xnor g9264 ( n6387 , n12703 , n8033 );
    not g9265 ( n3489 , n5078 );
    and g9266 ( n5744 , n6377 , n12854 );
    nor g9267 ( n1572 , n7824 , n12880 );
    or g9268 ( n2338 , n8687 , n4654 );
    and g9269 ( n4490 , n1839 , n4585 );
    xnor g9270 ( n10015 , n12556 , n997 );
    not g9271 ( n4381 , n11189 );
    xnor g9272 ( n8990 , n820 , n12499 );
    or g9273 ( n3866 , n3414 , n5170 );
    xnor g9274 ( n218 , n4112 , n2282 );
    nor g9275 ( n8209 , n4766 , n9346 );
    xnor g9276 ( n12412 , n9081 , n3026 );
    or g9277 ( n5050 , n10211 , n8355 );
    xnor g9278 ( n3089 , n2197 , n2281 );
    and g9279 ( n694 , n2191 , n3550 );
    or g9280 ( n1205 , n8959 , n2815 );
    or g9281 ( n9274 , n10835 , n5914 );
    xnor g9282 ( n8811 , n11149 , n7385 );
    xnor g9283 ( n12255 , n12550 , n9946 );
    or g9284 ( n10035 , n2639 , n6420 );
    not g9285 ( n8817 , n5059 );
    nor g9286 ( n12544 , n2271 , n2399 );
    and g9287 ( n6867 , n6776 , n10439 );
    or g9288 ( n2401 , n989 , n9589 );
    or g9289 ( n2511 , n6740 , n9524 );
    or g9290 ( n2852 , n12853 , n10422 );
    or g9291 ( n4667 , n6570 , n11756 );
    not g9292 ( n5867 , n11840 );
    or g9293 ( n6451 , n8959 , n5540 );
    or g9294 ( n3116 , n5530 , n7136 );
    xnor g9295 ( n538 , n5386 , n12572 );
    and g9296 ( n1868 , n12423 , n7303 );
    not g9297 ( n8756 , n8784 );
    or g9298 ( n2116 , n8959 , n7425 );
    or g9299 ( n3441 , n3746 , n6084 );
    xnor g9300 ( n8331 , n7 , n4663 );
    and g9301 ( n4783 , n3242 , n6957 );
    xnor g9302 ( n2889 , n8551 , n12230 );
    not g9303 ( n12439 , n10841 );
    xnor g9304 ( n11360 , n12040 , n11349 );
    and g9305 ( n717 , n9077 , n5332 );
    nor g9306 ( n11692 , n758 , n2826 );
    or g9307 ( n882 , n3617 , n12535 );
    or g9308 ( n3874 , n11653 , n4524 );
    xnor g9309 ( n10031 , n6037 , n5347 );
    or g9310 ( n8758 , n5355 , n9589 );
    xnor g9311 ( n9516 , n7602 , n1841 );
    xnor g9312 ( n3008 , n7115 , n2330 );
    nor g9313 ( n11506 , n11460 , n12888 );
    or g9314 ( n11962 , n8220 , n7838 );
    xnor g9315 ( n12222 , n3579 , n8300 );
    xnor g9316 ( n5163 , n11013 , n2022 );
    xnor g9317 ( n3500 , n8149 , n109 );
    or g9318 ( n6027 , n660 , n2927 );
    not g9319 ( n7856 , n953 );
    nor g9320 ( n7918 , n9606 , n679 );
    xnor g9321 ( n9131 , n666 , n10519 );
    and g9322 ( n4492 , n7854 , n4952 );
    nor g9323 ( n596 , n5881 , n10150 );
    and g9324 ( n8556 , n2393 , n7294 );
    not g9325 ( n12478 , n2476 );
    xnor g9326 ( n5176 , n5660 , n6107 );
    xnor g9327 ( n1221 , n5898 , n3139 );
    xnor g9328 ( n702 , n8458 , n3761 );
    or g9329 ( n6796 , n5369 , n4259 );
    xnor g9330 ( n7299 , n1864 , n10145 );
    nor g9331 ( n5171 , n3910 , n6548 );
    xnor g9332 ( n11308 , n8914 , n11802 );
    or g9333 ( n1705 , n5355 , n7424 );
    and g9334 ( n1426 , n1848 , n1374 );
    xnor g9335 ( n3372 , n5635 , n4056 );
    xnor g9336 ( n10723 , n10448 , n6747 );
    and g9337 ( n10668 , n6681 , n10894 );
    and g9338 ( n10933 , n7765 , n4208 );
    xnor g9339 ( n1751 , n2459 , n4594 );
    or g9340 ( n7499 , n9389 , n2358 );
    and g9341 ( n6988 , n5283 , n7610 );
    not g9342 ( n12229 , n12241 );
    or g9343 ( n8871 , n8429 , n10376 );
    or g9344 ( n5404 , n8187 , n7881 );
    nor g9345 ( n9957 , n11659 , n11408 );
    or g9346 ( n11605 , n5765 , n6922 );
    not g9347 ( n12211 , n7850 );
    not g9348 ( n8330 , n10689 );
    or g9349 ( n9120 , n9702 , n4844 );
    xnor g9350 ( n5352 , n12539 , n10409 );
    or g9351 ( n9325 , n2133 , n11530 );
    not g9352 ( n767 , n9882 );
    not g9353 ( n2653 , n10686 );
    or g9354 ( n10840 , n8870 , n5468 );
    not g9355 ( n9279 , n7668 );
    not g9356 ( n5518 , n721 );
    not g9357 ( n1476 , n6611 );
    or g9358 ( n7903 , n5366 , n5004 );
    xor g9359 ( n8640 , n5108 , n8939 );
    or g9360 ( n7111 , n6373 , n4654 );
    or g9361 ( n4324 , n6098 , n1845 );
    or g9362 ( n11613 , n3820 , n1047 );
    and g9363 ( n8207 , n9687 , n11344 );
    xnor g9364 ( n5443 , n7012 , n3834 );
    not g9365 ( n6510 , n7929 );
    or g9366 ( n9239 , n7268 , n1767 );
    not g9367 ( n10942 , n10214 );
    or g9368 ( n282 , n9389 , n6389 );
    not g9369 ( n4207 , n11323 );
    xnor g9370 ( n1977 , n10834 , n6624 );
    xnor g9371 ( n8562 , n9404 , n9679 );
    not g9372 ( n8655 , n4826 );
    xnor g9373 ( n10484 , n7284 , n365 );
    or g9374 ( n10881 , n11998 , n11648 );
    xnor g9375 ( n2888 , n4023 , n7696 );
    or g9376 ( n6073 , n10142 , n4242 );
    nor g9377 ( n5657 , n8117 , n745 );
    xnor g9378 ( n5906 , n9627 , n833 );
    or g9379 ( n5525 , n7391 , n3911 );
    not g9380 ( n11199 , n7370 );
    xnor g9381 ( n11776 , n11754 , n3814 );
    and g9382 ( n7890 , n10531 , n1467 );
    or g9383 ( n4995 , n10065 , n198 );
    xnor g9384 ( n9788 , n7666 , n11010 );
    or g9385 ( n10576 , n5495 , n10986 );
    xnor g9386 ( n11640 , n12500 , n2829 );
    not g9387 ( n10623 , n5408 );
    xnor g9388 ( n11693 , n5059 , n4099 );
    or g9389 ( n2390 , n1064 , n4813 );
    xnor g9390 ( n1030 , n3381 , n10811 );
    nor g9391 ( n5470 , n120 , n65 );
    nor g9392 ( n487 , n12939 , n6858 );
    or g9393 ( n443 , n6368 , n1309 );
    nor g9394 ( n6721 , n7680 , n8662 );
    xnor g9395 ( n12003 , n822 , n7162 );
    or g9396 ( n8905 , n12237 , n12735 );
    and g9397 ( n11500 , n2997 , n6848 );
    or g9398 ( n8145 , n9373 , n7506 );
    and g9399 ( n7735 , n5331 , n1512 );
    or g9400 ( n6218 , n8011 , n4866 );
    or g9401 ( n9843 , n8310 , n2912 );
    or g9402 ( n3155 , n357 , n5306 );
    xnor g9403 ( n395 , n7635 , n10300 );
    not g9404 ( n1799 , n4914 );
    or g9405 ( n1182 , n62 , n377 );
    or g9406 ( n12673 , n5361 , n6282 );
    nor g9407 ( n12137 , n10514 , n11187 );
    nor g9408 ( n12434 , n4779 , n4890 );
    xnor g9409 ( n7122 , n7622 , n10067 );
    xnor g9410 ( n4253 , n7675 , n6828 );
    and g9411 ( n2941 , n3962 , n4463 );
    xnor g9412 ( n780 , n5707 , n9944 );
    or g9413 ( n6161 , n989 , n2076 );
    xnor g9414 ( n3827 , n6882 , n6622 );
    not g9415 ( n10055 , n6773 );
    xnor g9416 ( n11870 , n6660 , n7096 );
    nor g9417 ( n3402 , n2443 , n3859 );
    and g9418 ( n142 , n5621 , n4075 );
    and g9419 ( n6413 , n12133 , n6866 );
    and g9420 ( n4256 , n5893 , n6088 );
    xnor g9421 ( n5565 , n1046 , n3683 );
    not g9422 ( n919 , n11336 );
    and g9423 ( n5278 , n5527 , n1217 );
    or g9424 ( n11518 , n8273 , n4909 );
    not g9425 ( n526 , n4292 );
    or g9426 ( n9570 , n989 , n1915 );
    not g9427 ( n261 , n8035 );
    xnor g9428 ( n7531 , n7614 , n471 );
    or g9429 ( n8674 , n10157 , n10916 );
    and g9430 ( n2500 , n4870 , n500 );
    xnor g9431 ( n5030 , n4323 , n7426 );
    and g9432 ( n11187 , n2520 , n1745 );
    nor g9433 ( n10235 , n8596 , n3584 );
    xnor g9434 ( n3086 , n720 , n12516 );
    xnor g9435 ( n2343 , n11396 , n4847 );
    not g9436 ( n6630 , n6059 );
    xnor g9437 ( n11789 , n1461 , n7491 );
    nor g9438 ( n2865 , n5715 , n7720 );
    or g9439 ( n2607 , n1469 , n10489 );
    or g9440 ( n4777 , n3743 , n5258 );
    or g9441 ( n8112 , n966 , n11943 );
    or g9442 ( n5982 , n8870 , n826 );
    or g9443 ( n54 , n12361 , n6084 );
    nor g9444 ( n12898 , n4511 , n8863 );
    xnor g9445 ( n11224 , n8267 , n11939 );
    not g9446 ( n6991 , n12215 );
    or g9447 ( n11370 , n989 , n3911 );
    or g9448 ( n12858 , n3743 , n609 );
    xnor g9449 ( n9115 , n4289 , n3035 );
    xnor g9450 ( n9941 , n601 , n3269 );
    xnor g9451 ( n1884 , n577 , n8482 );
    and g9452 ( n12560 , n4263 , n8131 );
    xnor g9453 ( n9539 , n8293 , n12519 );
    or g9454 ( n7996 , n962 , n4654 );
    and g9455 ( n6029 , n12443 , n1734 );
    or g9456 ( n7564 , n10142 , n12328 );
    not g9457 ( n7186 , n3313 );
    and g9458 ( n5082 , n173 , n3686 );
    xnor g9459 ( n1034 , n10031 , n5467 );
    or g9460 ( n5532 , n8687 , n2020 );
    not g9461 ( n12235 , n3991 );
    or g9462 ( n2282 , n11923 , n12771 );
    or g9463 ( n8848 , n10196 , n2020 );
    or g9464 ( n12913 , n4911 , n10066 );
    and g9465 ( n10517 , n11311 , n2522 );
    not g9466 ( n530 , n4970 );
    xnor g9467 ( n3432 , n2033 , n8014 );
    and g9468 ( n3593 , n7358 , n466 );
    xnor g9469 ( n4542 , n4298 , n1001 );
    or g9470 ( n2722 , n12423 , n7303 );
    and g9471 ( n6243 , n1415 , n4630 );
    not g9472 ( n7138 , n6121 );
    xnor g9473 ( n1346 , n4449 , n4391 );
    xnor g9474 ( n6860 , n12693 , n10616 );
    and g9475 ( n5172 , n3533 , n5660 );
    not g9476 ( n8031 , n4417 );
    and g9477 ( n1697 , n5855 , n3487 );
    or g9478 ( n3474 , n114 , n7876 );
    not g9479 ( n4267 , n3807 );
    or g9480 ( n3487 , n11051 , n9731 );
    or g9481 ( n2524 , n3611 , n11027 );
    xnor g9482 ( n7242 , n3305 , n6890 );
    xnor g9483 ( n8399 , n10873 , n1950 );
    or g9484 ( n6509 , n8480 , n5865 );
    xnor g9485 ( n11565 , n4442 , n11248 );
    or g9486 ( n1157 , n1941 , n6455 );
    and g9487 ( n10878 , n5363 , n3006 );
    xnor g9488 ( n8605 , n10814 , n7368 );
    or g9489 ( n8423 , n11958 , n6197 );
    and g9490 ( n4045 , n8557 , n7653 );
    xnor g9491 ( n3641 , n2061 , n1158 );
    xnor g9492 ( n2855 , n4755 , n11338 );
    not g9493 ( n8615 , n9737 );
    not g9494 ( n10464 , n9326 );
    xnor g9495 ( n6653 , n7480 , n1080 );
    xnor g9496 ( n8044 , n12526 , n5750 );
    or g9497 ( n2858 , n6298 , n6721 );
    and g9498 ( n10872 , n6077 , n11715 );
    and g9499 ( n6111 , n3106 , n11945 );
    xnor g9500 ( n2803 , n2284 , n11102 );
    nor g9501 ( n7220 , n4431 , n6243 );
    not g9502 ( n11026 , n2393 );
    xnor g9503 ( n2961 , n5204 , n283 );
    xnor g9504 ( n9804 , n11782 , n5114 );
    not g9505 ( n12218 , n12747 );
    not g9506 ( n7558 , n2522 );
    or g9507 ( n11425 , n2217 , n5258 );
    nor g9508 ( n4614 , n8503 , n3889 );
    xnor g9509 ( n5733 , n10452 , n10676 );
    or g9510 ( n11192 , n962 , n9160 );
    xnor g9511 ( n9133 , n11945 , n6487 );
    not g9512 ( n8714 , n4603 );
    not g9513 ( n2931 , n7490 );
    xnor g9514 ( n7693 , n129 , n9330 );
    and g9515 ( n9702 , n2195 , n1101 );
    nor g9516 ( n6525 , n391 , n1821 );
    xnor g9517 ( n10914 , n1644 , n11612 );
    nor g9518 ( n9183 , n5503 , n730 );
    not g9519 ( n7970 , n9727 );
    not g9520 ( n679 , n7647 );
    xnor g9521 ( n8333 , n4866 , n8252 );
    not g9522 ( n7739 , n11575 );
    xnor g9523 ( n4880 , n12305 , n3223 );
    or g9524 ( n3700 , n1872 , n3556 );
    or g9525 ( n11352 , n5575 , n7876 );
    or g9526 ( n6235 , n4053 , n10130 );
    nor g9527 ( n1578 , n1879 , n142 );
    or g9528 ( n358 , n8959 , n2232 );
    not g9529 ( n7090 , n12790 );
    or g9530 ( n2625 , n10157 , n609 );
    xnor g9531 ( n1032 , n4690 , n8965 );
    and g9532 ( n3163 , n7432 , n5058 );
    xnor g9533 ( n11300 , n9557 , n4574 );
    and g9534 ( n3692 , n11475 , n7800 );
    nor g9535 ( n3463 , n737 , n6132 );
    and g9536 ( n7734 , n1172 , n3669 );
    not g9537 ( n3818 , n9508 );
    xnor g9538 ( n8360 , n11588 , n9112 );
    not g9539 ( n5389 , n1062 );
    and g9540 ( n9050 , n11542 , n6333 );
    not g9541 ( n7755 , n8533 );
    and g9542 ( n5010 , n10594 , n6540 );
    xnor g9543 ( n1158 , n7297 , n7935 );
    or g9544 ( n6224 , n10108 , n12843 );
    or g9545 ( n12659 , n3743 , n5502 );
    or g9546 ( n8215 , n11753 , n3341 );
    or g9547 ( n2204 , n11719 , n11827 );
    and g9548 ( n7321 , n8430 , n1452 );
    not g9549 ( n1148 , n8460 );
    or g9550 ( n7967 , n12023 , n7734 );
    nor g9551 ( n3857 , n2881 , n7744 );
    and g9552 ( n4799 , n6437 , n12847 );
    xnor g9553 ( n5587 , n1355 , n7273 );
    or g9554 ( n5944 , n6718 , n4864 );
    xnor g9555 ( n345 , n6931 , n1197 );
    or g9556 ( n9058 , n2427 , n1157 );
    or g9557 ( n9248 , n7586 , n1505 );
    not g9558 ( n211 , n3536 );
    xnor g9559 ( n11414 , n1784 , n11686 );
    xnor g9560 ( n3611 , n7856 , n2798 );
    or g9561 ( n1393 , n7381 , n865 );
    xnor g9562 ( n12806 , n320 , n12447 );
    xnor g9563 ( n7917 , n11360 , n2803 );
    and g9564 ( n1338 , n2101 , n3422 );
    nor g9565 ( n11056 , n5269 , n12488 );
    or g9566 ( n1066 , n8450 , n10025 );
    not g9567 ( n1843 , n7652 );
    and g9568 ( n5445 , n664 , n9991 );
    or g9569 ( n6312 , n1699 , n4913 );
    or g9570 ( n9884 , n994 , n7703 );
    or g9571 ( n3145 , n5575 , n995 );
    not g9572 ( n126 , n5789 );
    xnor g9573 ( n3139 , n849 , n329 );
    xnor g9574 ( n12908 , n3265 , n1454 );
    or g9575 ( n11592 , n5393 , n6733 );
    xnor g9576 ( n8609 , n10516 , n778 );
    or g9577 ( n5485 , n11026 , n4527 );
    xnor g9578 ( n11264 , n2673 , n2648 );
    xnor g9579 ( n8278 , n9616 , n5262 );
    or g9580 ( n6030 , n3544 , n4715 );
    not g9581 ( n6852 , n7419 );
    or g9582 ( n12318 , n5575 , n184 );
    or g9583 ( n5619 , n6171 , n7351 );
    xnor g9584 ( n9654 , n3921 , n429 );
    xnor g9585 ( n4344 , n2503 , n5908 );
    xnor g9586 ( n2264 , n8023 , n9300 );
    nor g9587 ( n11761 , n2162 , n7307 );
    not g9588 ( n2079 , n11633 );
    and g9589 ( n4882 , n4791 , n5762 );
    not g9590 ( n2386 , n10923 );
    or g9591 ( n3130 , n3820 , n4654 );
    and g9592 ( n147 , n12648 , n2802 );
    xnor g9593 ( n7700 , n10958 , n540 );
    and g9594 ( n6982 , n12144 , n5251 );
    nor g9595 ( n5290 , n2309 , n3798 );
    xnor g9596 ( n7621 , n10992 , n14 );
    xnor g9597 ( n9840 , n248 , n11837 );
    not g9598 ( n6200 , n10457 );
    not g9599 ( n1160 , n822 );
    xnor g9600 ( n5705 , n9481 , n12507 );
    nor g9601 ( n63 , n12095 , n1578 );
    xnor g9602 ( n6428 , n5989 , n3457 );
    not g9603 ( n3674 , n10877 );
    or g9604 ( n11762 , n7329 , n8461 );
    or g9605 ( n9016 , n12119 , n8109 );
    xnor g9606 ( n606 , n6121 , n2158 );
    xnor g9607 ( n1420 , n7278 , n598 );
    not g9608 ( n8611 , n12628 );
    or g9609 ( n1374 , n8019 , n9631 );
    or g9610 ( n12497 , n209 , n4050 );
    and g9611 ( n3773 , n10309 , n11180 );
    or g9612 ( n9504 , n5530 , n8655 );
    and g9613 ( n7960 , n810 , n2058 );
    not g9614 ( n4983 , n7612 );
    and g9615 ( n2966 , n11892 , n806 );
    and g9616 ( n1178 , n4097 , n11394 );
    and g9617 ( n9830 , n6478 , n3855 );
    or g9618 ( n4112 , n5765 , n9568 );
    or g9619 ( n10091 , n7116 , n11820 );
    xnor g9620 ( n1905 , n2858 , n5772 );
    not g9621 ( n1277 , n2784 );
    xnor g9622 ( n10861 , n12715 , n11494 );
    not g9623 ( n9751 , n5688 );
    not g9624 ( n5502 , n159 );
    or g9625 ( n257 , n11594 , n272 );
    or g9626 ( n10688 , n5700 , n2958 );
    not g9627 ( n2412 , n628 );
    or g9628 ( n614 , n573 , n11044 );
    and g9629 ( n10802 , n5479 , n8519 );
    xnor g9630 ( n1860 , n8070 , n473 );
    xnor g9631 ( n6767 , n8774 , n3152 );
    xnor g9632 ( n6705 , n10407 , n2755 );
    nor g9633 ( n10864 , n11734 , n6862 );
    not g9634 ( n11251 , n9007 );
    xnor g9635 ( n12279 , n5361 , n12729 );
    not g9636 ( n5507 , n904 );
    or g9637 ( n5658 , n10157 , n9160 );
    and g9638 ( n1039 , n1518 , n211 );
    or g9639 ( n5718 , n7391 , n6389 );
    xnor g9640 ( n11279 , n12782 , n2379 );
    xnor g9641 ( n1707 , n6536 , n6532 );
    and g9642 ( n2999 , n255 , n4288 );
    or g9643 ( n1123 , n752 , n9971 );
    or g9644 ( n9256 , n3348 , n67 );
    or g9645 ( n8881 , n5620 , n9864 );
    nor g9646 ( n11032 , n2574 , n1190 );
    and g9647 ( n4545 , n4214 , n7650 );
    and g9648 ( n7879 , n8452 , n8978 );
    not g9649 ( n4448 , n3914 );
    not g9650 ( n962 , n1471 );
    xnor g9651 ( n4454 , n5856 , n10890 );
    or g9652 ( n2288 , n4112 , n2282 );
    xnor g9653 ( n11134 , n5554 , n12161 );
    not g9654 ( n4873 , n12939 );
    or g9655 ( n9299 , n3160 , n1116 );
    xnor g9656 ( n5090 , n8103 , n5741 );
    nor g9657 ( n2601 , n3235 , n407 );
    or g9658 ( n6214 , n11413 , n937 );
    xnor g9659 ( n1037 , n6987 , n3200 );
    and g9660 ( n6521 , n5195 , n4478 );
    not g9661 ( n4766 , n10117 );
    and g9662 ( n4331 , n9185 , n3250 );
    and g9663 ( n1036 , n8453 , n4625 );
    xnor g9664 ( n343 , n11119 , n7274 );
    and g9665 ( n942 , n1947 , n11587 );
    and g9666 ( n7245 , n11073 , n5965 );
    xnor g9667 ( n11323 , n10096 , n4208 );
    or g9668 ( n2100 , n9878 , n4913 );
    or g9669 ( n7604 , n6854 , n2439 );
    or g9670 ( n10050 , n612 , n9775 );
    and g9671 ( n10521 , n10242 , n12660 );
    xnor g9672 ( n6937 , n1483 , n5676 );
    or g9673 ( n1131 , n2456 , n7928 );
    or g9674 ( n800 , n3361 , n1243 );
    xnor g9675 ( n6610 , n12739 , n6652 );
    not g9676 ( n11823 , n4435 );
    nor g9677 ( n12018 , n9899 , n3737 );
    xnor g9678 ( n9127 , n10738 , n6451 );
    not g9679 ( n3686 , n11498 );
    and g9680 ( n10817 , n12622 , n3919 );
    or g9681 ( n9744 , n191 , n8859 );
    not g9682 ( n5567 , n2376 );
    not g9683 ( n12147 , n10918 );
    or g9684 ( n2190 , n6977 , n6084 );
    not g9685 ( n2823 , n1210 );
    xnor g9686 ( n4374 , n6557 , n11804 );
    xnor g9687 ( n7793 , n8872 , n11270 );
    nor g9688 ( n2025 , n3372 , n6124 );
    xnor g9689 ( n2929 , n3633 , n3825 );
    or g9690 ( n5289 , n9448 , n4181 );
    xnor g9691 ( n9848 , n11727 , n1119 );
    nor g9692 ( n7055 , n9342 , n11970 );
    or g9693 ( n5477 , n5252 , n3309 );
    not g9694 ( n10750 , n12391 );
    xnor g9695 ( n68 , n7016 , n11437 );
    nor g9696 ( n11845 , n656 , n10580 );
    xnor g9697 ( n5478 , n5243 , n11640 );
    and g9698 ( n7511 , n8549 , n2493 );
    or g9699 ( n11743 , n9054 , n10082 );
    xnor g9700 ( n9855 , n2859 , n2949 );
    or g9701 ( n11689 , n9370 , n5497 );
    and g9702 ( n4375 , n2254 , n10227 );
    xnor g9703 ( n7211 , n4759 , n929 );
    or g9704 ( n9871 , n11923 , n9280 );
    or g9705 ( n1973 , n11958 , n2232 );
    or g9706 ( n3377 , n591 , n11790 );
    xnor g9707 ( n6315 , n95 , n5882 );
    xnor g9708 ( n6809 , n6700 , n6120 );
    xnor g9709 ( n3779 , n6212 , n10328 );
    and g9710 ( n1362 , n12721 , n6196 );
    nor g9711 ( n12931 , n8294 , n6316 );
    and g9712 ( n6897 , n3628 , n894 );
    nor g9713 ( n12430 , n4613 , n4098 );
    not g9714 ( n10468 , n9608 );
    xnor g9715 ( n2942 , n8816 , n1217 );
    xor g9716 ( n5189 , n8928 , n2974 );
    or g9717 ( n3544 , n11958 , n3421 );
    nor g9718 ( n11486 , n9161 , n2531 );
    and g9719 ( n6665 , n3998 , n608 );
    xnor g9720 ( n1211 , n2598 , n265 );
    nor g9721 ( n3329 , n6782 , n7054 );
    xnor g9722 ( n567 , n3141 , n4721 );
    xnor g9723 ( n10232 , n6738 , n252 );
    or g9724 ( n4458 , n12853 , n6513 );
    xnor g9725 ( n3385 , n5621 , n1879 );
    and g9726 ( n4700 , n2923 , n7999 );
    or g9727 ( n8641 , n1642 , n12325 );
    xnor g9728 ( n2958 , n5863 , n3149 );
    and g9729 ( n11477 , n12758 , n7584 );
    xnor g9730 ( n7811 , n6750 , n3701 );
    not g9731 ( n5727 , n3815 );
    not g9732 ( n7443 , n6364 );
    or g9733 ( n7052 , n9007 , n7956 );
    and g9734 ( n8140 , n9105 , n1981 );
    and g9735 ( n12573 , n7128 , n6684 );
    nor g9736 ( n4359 , n12117 , n143 );
    and g9737 ( n274 , n9453 , n9646 );
    and g9738 ( n5180 , n7694 , n12015 );
    or g9739 ( n4460 , n1699 , n12535 );
    or g9740 ( n3108 , n807 , n6455 );
    xnor g9741 ( n7366 , n10619 , n11819 );
    and g9742 ( n9833 , n3105 , n358 );
    not g9743 ( n5699 , n7997 );
    not g9744 ( n239 , n8864 );
    xnor g9745 ( n6488 , n5080 , n7917 );
    xnor g9746 ( n6912 , n11677 , n1025 );
    or g9747 ( n697 , n8552 , n9188 );
    not g9748 ( n2107 , n1113 );
    or g9749 ( n8221 , n12853 , n1932 );
    not g9750 ( n8970 , n11536 );
    and g9751 ( n344 , n204 , n6608 );
    and g9752 ( n4428 , n3110 , n4940 );
    and g9753 ( n3211 , n10791 , n8508 );
    and g9754 ( n4602 , n8858 , n4452 );
    or g9755 ( n347 , n5685 , n5658 );
    and g9756 ( n3513 , n5950 , n5359 );
    not g9757 ( n10248 , n4181 );
    not g9758 ( n1486 , n3326 );
    or g9759 ( n9066 , n7468 , n271 );
    nor g9760 ( n10093 , n6085 , n12029 );
    or g9761 ( n2933 , n9878 , n826 );
    and g9762 ( n4175 , n1024 , n7498 );
    xnor g9763 ( n1482 , n7621 , n8614 );
    not g9764 ( n5937 , n11136 );
    and g9765 ( n12780 , n1089 , n10310 );
    or g9766 ( n4016 , n6637 , n461 );
    or g9767 ( n11673 , n6739 , n9109 );
    or g9768 ( n10846 , n7283 , n1851 );
    xnor g9769 ( n2622 , n9290 , n6049 );
    not g9770 ( n2437 , n6539 );
    or g9771 ( n8410 , n8702 , n8911 );
    and g9772 ( n2357 , n2176 , n8516 );
    and g9773 ( n1416 , n5158 , n7751 );
    or g9774 ( n6122 , n6577 , n6084 );
    xnor g9775 ( n5563 , n6447 , n11891 );
    or g9776 ( n7927 , n5671 , n1134 );
    not g9777 ( n10607 , n8445 );
    and g9778 ( n9180 , n3611 , n11027 );
    and g9779 ( n9285 , n10148 , n7996 );
    nor g9780 ( n4649 , n7493 , n8551 );
    xnor g9781 ( n10069 , n6470 , n7392 );
    xnor g9782 ( n5221 , n4981 , n12209 );
    or g9783 ( n1334 , n4059 , n510 );
    not g9784 ( n4843 , n11388 );
    and g9785 ( n10130 , n8996 , n9518 );
    xnor g9786 ( n5825 , n12545 , n1180 );
    nor g9787 ( n9008 , n10225 , n3598 );
    not g9788 ( n10422 , n2551 );
    xnor g9789 ( n10213 , n11205 , n11622 );
    or g9790 ( n8094 , n6439 , n6447 );
    not g9791 ( n3530 , n3170 );
    xnor g9792 ( n9371 , n7380 , n11427 );
    or g9793 ( n1668 , n3740 , n10116 );
    nor g9794 ( n9951 , n8879 , n7199 );
    and g9795 ( n7647 , n5330 , n1401 );
    and g9796 ( n3941 , n11709 , n831 );
    or g9797 ( n3926 , n11181 , n4268 );
    nor g9798 ( n9503 , n10598 , n2601 );
    and g9799 ( n11239 , n1409 , n12780 );
    xnor g9800 ( n5557 , n1629 , n5509 );
    xnor g9801 ( n98 , n7910 , n8706 );
    not g9802 ( n6674 , n4746 );
    or g9803 ( n6952 , n10142 , n6524 );
    nor g9804 ( n8781 , n1341 , n9522 );
    nor g9805 ( n2194 , n7433 , n1884 );
    or g9806 ( n4424 , n6718 , n9280 );
    not g9807 ( n9247 , n10742 );
    xnor g9808 ( n9558 , n12723 , n1584 );
    or g9809 ( n11674 , n7449 , n4875 );
    nor g9810 ( n803 , n3925 , n4797 );
    nor g9811 ( n10158 , n11844 , n6991 );
    and g9812 ( n11577 , n8276 , n2024 );
    xnor g9813 ( n5927 , n12227 , n11940 );
    xnor g9814 ( n1950 , n1530 , n1115 );
    or g9815 ( n337 , n4628 , n7382 );
    and g9816 ( n8335 , n12579 , n6506 );
    and g9817 ( n9993 , n7231 , n6505 );
    or g9818 ( n11935 , n11923 , n7506 );
    xnor g9819 ( n9069 , n9848 , n2568 );
    or g9820 ( n2520 , n2730 , n3094 );
    or g9821 ( n2490 , n4343 , n9188 );
    xnor g9822 ( n5155 , n7318 , n8993 );
    and g9823 ( n1525 , n9369 , n2952 );
    or g9824 ( n12734 , n6577 , n7558 );
    or g9825 ( n2660 , n6181 , n10334 );
    xnor g9826 ( n744 , n9353 , n9243 );
    and g9827 ( n11098 , n961 , n9553 );
    or g9828 ( n7019 , n6373 , n5502 );
    nor g9829 ( n1772 , n9735 , n12481 );
    or g9830 ( n325 , n10196 , n4527 );
    or g9831 ( n8764 , n9277 , n9473 );
    xnor g9832 ( n11075 , n11783 , n2 );
    xnor g9833 ( n9811 , n7393 , n11507 );
    xnor g9834 ( n1925 , n10169 , n2473 );
    not g9835 ( n9333 , n6507 );
    and g9836 ( n12179 , n885 , n5836 );
    nor g9837 ( n618 , n5773 , n12664 );
    xnor g9838 ( n5992 , n8417 , n9857 );
    or g9839 ( n7771 , n12150 , n538 );
    and g9840 ( n12664 , n10763 , n11582 );
    and g9841 ( n4813 , n2516 , n11559 );
    not g9842 ( n8746 , n4919 );
    xnor g9843 ( n8314 , n675 , n2290 );
    or g9844 ( n1653 , n2217 , n1047 );
    or g9845 ( n2496 , n2252 , n8340 );
    not g9846 ( n11111 , n10702 );
    or g9847 ( n2901 , n515 , n5941 );
    xnor g9848 ( n8517 , n2605 , n11921 );
    or g9849 ( n317 , n5355 , n8970 );
    xnor g9850 ( n5244 , n7054 , n1040 );
    xnor g9851 ( n210 , n8294 , n7317 );
    or g9852 ( n11749 , n7512 , n12181 );
    xnor g9853 ( n12534 , n302 , n12214 );
    and g9854 ( n11560 , n7299 , n2239 );
    and g9855 ( n8338 , n4029 , n8834 );
    xnor g9856 ( n11643 , n11212 , n12002 );
    and g9857 ( n8069 , n12825 , n8744 );
    and g9858 ( n3192 , n404 , n429 );
    or g9859 ( n10056 , n807 , n6169 );
    not g9860 ( n12356 , n8823 );
    and g9861 ( n690 , n7947 , n493 );
    not g9862 ( n1078 , n9347 );
    or g9863 ( n7051 , n6602 , n2951 );
    xnor g9864 ( n1991 , n10254 , n8833 );
    xnor g9865 ( n4236 , n3330 , n7693 );
    or g9866 ( n2983 , n5915 , n6071 );
    xnor g9867 ( n10927 , n9456 , n3101 );
    or g9868 ( n2466 , n1409 , n12780 );
    nor g9869 ( n5238 , n8380 , n1786 );
    or g9870 ( n1506 , n686 , n995 );
    and g9871 ( n8220 , n1249 , n7963 );
    xnor g9872 ( n2777 , n4007 , n7095 );
    or g9873 ( n1678 , n4643 , n8913 );
    or g9874 ( n5679 , n2217 , n9568 );
    or g9875 ( n7959 , n10157 , n28 );
    xnor g9876 ( n8146 , n8741 , n2942 );
    or g9877 ( n2838 , n5575 , n5538 );
    xnor g9878 ( n4293 , n11317 , n916 );
    and g9879 ( n4321 , n10347 , n12182 );
    or g9880 ( n10414 , n7449 , n12120 );
    xnor g9881 ( n11348 , n532 , n480 );
    not g9882 ( n410 , n1218 );
    not g9883 ( n9399 , n8529 );
    or g9884 ( n5207 , n994 , n3911 );
    or g9885 ( n9849 , n1941 , n3903 );
    xnor g9886 ( n6035 , n9141 , n901 );
    and g9887 ( n3226 , n586 , n6172 );
    nor g9888 ( n1417 , n372 , n1060 );
    and g9889 ( n12678 , n12471 , n6433 );
    xnor g9890 ( n8087 , n3044 , n7066 );
    not g9891 ( n7420 , n478 );
    xnor g9892 ( n12490 , n2277 , n4865 );
    not g9893 ( n2358 , n4634 );
    not g9894 ( n8858 , n5157 );
    or g9895 ( n8702 , n5008 , n6841 );
    xnor g9896 ( n5035 , n8085 , n11814 );
    and g9897 ( n9411 , n12870 , n10107 );
    xnor g9898 ( n10106 , n3105 , n358 );
    not g9899 ( n8733 , n6483 );
    or g9900 ( n2904 , n3457 , n3786 );
    or g9901 ( n4184 , n4457 , n622 );
    and g9902 ( n1659 , n4001 , n592 );
    or g9903 ( n10613 , n2217 , n1739 );
    nor g9904 ( n3473 , n7373 , n1340 );
    not g9905 ( n7875 , n12653 );
    xnor g9906 ( n1916 , n8992 , n5106 );
    not g9907 ( n5497 , n5212 );
    not g9908 ( n6648 , n6599 );
    not g9909 ( n1636 , n4406 );
    or g9910 ( n10772 , n722 , n3987 );
    nor g9911 ( n3183 , n5208 , n4917 );
    or g9912 ( n3887 , n7462 , n2105 );
    not g9913 ( n1519 , n8449 );
    or g9914 ( n12208 , n2456 , n1163 );
    or g9915 ( n3007 , n3127 , n7341 );
    and g9916 ( n8760 , n11293 , n6013 );
    nor g9917 ( n8218 , n5288 , n3040 );
    not g9918 ( n115 , n9512 );
    nor g9919 ( n5271 , n331 , n11840 );
    xnor g9920 ( n12389 , n11798 , n11143 );
    or g9921 ( n10793 , n10325 , n10127 );
    and g9922 ( n5248 , n3906 , n11203 );
    nor g9923 ( n2819 , n9551 , n4044 );
    or g9924 ( n582 , n10750 , n12080 );
    xnor g9925 ( n7935 , n9559 , n5050 );
    and g9926 ( n3953 , n1097 , n7456 );
    not g9927 ( n12754 , n447 );
    and g9928 ( n10342 , n11812 , n6879 );
    nor g9929 ( n5267 , n135 , n11786 );
    xnor g9930 ( n4095 , n3045 , n8558 );
    xnor g9931 ( n10549 , n10551 , n7988 );
    xnor g9932 ( n145 , n9519 , n1648 );
    or g9933 ( n10645 , n2455 , n2567 );
    or g9934 ( n2700 , n8959 , n7952 );
    not g9935 ( n1881 , n6415 );
    or g9936 ( n1041 , n10277 , n6343 );
    xnor g9937 ( n4690 , n11113 , n1005 );
    or g9938 ( n7131 , n686 , n6455 );
    xnor g9939 ( n7569 , n5437 , n7104 );
    xnor g9940 ( n7548 , n8757 , n5031 );
    nor g9941 ( n9897 , n10948 , n4359 );
    xnor g9942 ( n10612 , n11050 , n1336 );
    nor g9943 ( n8877 , n7091 , n5427 );
    xnor g9944 ( n8888 , n6880 , n12440 );
    and g9945 ( n11141 , n2515 , n12489 );
    xor g9946 ( n11326 , n3722 , n11793 );
    xnor g9947 ( n3403 , n10590 , n7821 );
    and g9948 ( n2089 , n692 , n8763 );
    xnor g9949 ( n3649 , n4956 , n10521 );
    xnor g9950 ( n3934 , n12470 , n4336 );
    xnor g9951 ( n6558 , n7791 , n1227 );
    nor g9952 ( n7003 , n3335 , n5740 );
    or g9953 ( n3961 , n240 , n983 );
    not g9954 ( n11827 , n7265 );
    not g9955 ( n4670 , n438 );
    xnor g9956 ( n513 , n5130 , n9831 );
    not g9957 ( n1936 , n7469 );
    or g9958 ( n1886 , n9050 , n2873 );
    xnor g9959 ( n6511 , n9797 , n2900 );
    and g9960 ( n5810 , n1012 , n11537 );
    and g9961 ( n3440 , n1543 , n1600 );
    or g9962 ( n2103 , n1752 , n2688 );
    xnor g9963 ( n7898 , n11683 , n7110 );
    or g9964 ( n12002 , n5915 , n12754 );
    or g9965 ( n10943 , n7625 , n2709 );
    or g9966 ( n11338 , n8405 , n6513 );
    or g9967 ( n2917 , n6977 , n6455 );
    xnor g9968 ( n5000 , n1135 , n9409 );
    or g9969 ( n8984 , n12611 , n1437 );
    nor g9970 ( n4060 , n9806 , n8579 );
    not g9971 ( n1526 , n5475 );
    and g9972 ( n5882 , n6979 , n6404 );
    xnor g9973 ( n6089 , n7301 , n3237 );
    not g9974 ( n7534 , n9647 );
    xnor g9975 ( n9857 , n5179 , n529 );
    and g9976 ( n10410 , n8596 , n3584 );
    or g9977 ( n8205 , n10750 , n5781 );
    not g9978 ( n11752 , n5167 );
    xnor g9979 ( n5038 , n7869 , n12455 );
    xnor g9980 ( n4962 , n11690 , n1914 );
    not g9981 ( n2798 , n10528 );
    or g9982 ( n12526 , n6577 , n3421 );
    nor g9983 ( n7870 , n11174 , n2863 );
    or g9984 ( n9093 , n4415 , n325 );
    nor g9985 ( n8288 , n12879 , n7792 );
    or g9986 ( n7058 , n9107 , n2986 );
    xnor g9987 ( n11919 , n7081 , n1713 );
    or g9988 ( n11014 , n636 , n5468 );
    or g9989 ( n10794 , n9531 , n1436 );
    nor g9990 ( n2279 , n4235 , n7828 );
    not g9991 ( n4073 , n1821 );
    and g9992 ( n2377 , n4167 , n6892 );
    xnor g9993 ( n4120 , n9733 , n10564 );
    not g9994 ( n6331 , n1361 );
    xnor g9995 ( n7418 , n2146 , n2636 );
    and g9996 ( n9838 , n4187 , n2024 );
    xnor g9997 ( n10630 , n1626 , n1376 );
    or g9998 ( n7380 , n6718 , n4527 );
    and g9999 ( n135 , n10831 , n10959 );
    and g10000 ( n5493 , n428 , n244 );
    and g10001 ( n3978 , n10727 , n5662 );
    or g10002 ( n12624 , n1335 , n1440 );
    or g10003 ( n6698 , n7138 , n935 );
    or g10004 ( n1115 , n8263 , n4545 );
    and g10005 ( n2761 , n2034 , n2851 );
    not g10006 ( n10369 , n2966 );
    and g10007 ( n5252 , n8641 , n3890 );
    xnor g10008 ( n6728 , n12831 , n2915 );
    not g10009 ( n1367 , n1804 );
    and g10010 ( n5160 , n9884 , n3411 );
    xnor g10011 ( n4567 , n10963 , n465 );
    not g10012 ( n11716 , n6159 );
    or g10013 ( n9179 , n5809 , n1932 );
    and g10014 ( n2548 , n5856 , n10890 );
    nor g10015 ( n7069 , n8555 , n11568 );
    and g10016 ( n9037 , n4272 , n11833 );
    or g10017 ( n9079 , n752 , n995 );
    or g10018 ( n12940 , n10607 , n341 );
    nor g10019 ( n8708 , n7005 , n1291 );
    nor g10020 ( n1875 , n6903 , n8419 );
    or g10021 ( n2448 , n5530 , n10422 );
    or g10022 ( n5391 , n6373 , n2020 );
    xnor g10023 ( n10125 , n11834 , n6459 );
    and g10024 ( n3801 , n3078 , n6895 );
    or g10025 ( n1402 , n11984 , n6460 );
    nor g10026 ( n10571 , n4217 , n11726 );
    xnor g10027 ( n298 , n9827 , n12893 );
    xnor g10028 ( n1110 , n3354 , n8604 );
    xnor g10029 ( n9025 , n7911 , n6753 );
    and g10030 ( n11019 , n808 , n9934 );
    nor g10031 ( n4039 , n6291 , n5035 );
    and g10032 ( n2826 , n7745 , n11854 );
    and g10033 ( n1074 , n9881 , n9474 );
    and g10034 ( n3655 , n9437 , n7908 );
    nor g10035 ( n9282 , n504 , n3873 );
    not g10036 ( n8334 , n8159 );
    or g10037 ( n12329 , n5915 , n8109 );
    xnor g10038 ( n2517 , n6133 , n9913 );
    or g10039 ( n12197 , n4358 , n10165 );
    or g10040 ( n10877 , n752 , n2815 );
    nor g10041 ( n3835 , n12476 , n485 );
    not g10042 ( n2678 , n7790 );
    or g10043 ( n3156 , n7009 , n4534 );
    and g10044 ( n8529 , n7236 , n9763 );
    or g10045 ( n11195 , n2124 , n3553 );
    or g10046 ( n12643 , n4859 , n2263 );
    or g10047 ( n7154 , n8187 , n7424 );
    or g10048 ( n301 , n7232 , n1013 );
    and g10049 ( n1966 , n10104 , n10498 );
    xnor g10050 ( n11333 , n3876 , n10111 );
    not g10051 ( n4229 , n3017 );
    or g10052 ( n196 , n4628 , n12735 );
    xnor g10053 ( n6856 , n5107 , n258 );
    nor g10054 ( n9221 , n1816 , n5037 );
    or g10055 ( n10463 , n3622 , n7803 );
    xnor g10056 ( n6722 , n5099 , n570 );
    or g10057 ( n5342 , n5902 , n10066 );
    and g10058 ( n6002 , n6776 , n10451 );
    or g10059 ( n4464 , n7391 , n12843 );
    not g10060 ( n10797 , n1131 );
    or g10061 ( n527 , n5655 , n2296 );
    xnor g10062 ( n11458 , n5394 , n5152 );
    or g10063 ( n2053 , n9914 , n1573 );
    nor g10064 ( n9755 , n843 , n717 );
    xnor g10065 ( n7966 , n5615 , n5717 );
    and g10066 ( n7302 , n6374 , n5757 );
    or g10067 ( n11623 , n3691 , n4315 );
    nor g10068 ( n8879 , n3464 , n8805 );
    and g10069 ( n1459 , n3571 , n4869 );
    or g10070 ( n2743 , n11846 , n7117 );
    or g10071 ( n4888 , n636 , n8644 );
    not g10072 ( n12191 , n9590 );
    not g10073 ( n7447 , n5206 );
    or g10074 ( n2287 , n7663 , n11886 );
    not g10075 ( n8957 , n10685 );
    nor g10076 ( n4354 , n1160 , n7162 );
    or g10077 ( n12333 , n9170 , n7703 );
    or g10078 ( n725 , n4327 , n8059 );
    and g10079 ( n295 , n1303 , n4754 );
    or g10080 ( n12188 , n6286 , n424 );
    or g10081 ( n6902 , n5562 , n4550 );
    not g10082 ( n3175 , n5039 );
    and g10083 ( n4004 , n8977 , n5040 );
    xnor g10084 ( n12201 , n7519 , n9371 );
    or g10085 ( n7955 , n3038 , n11124 );
    or g10086 ( n11679 , n5530 , n8109 );
    and g10087 ( n8947 , n9685 , n1926 );
    not g10088 ( n12237 , n4828 );
    or g10089 ( n12317 , n1883 , n105 );
    not g10090 ( n1162 , n2509 );
    xnor g10091 ( n8537 , n9440 , n7068 );
    or g10092 ( n4787 , n10750 , n1163 );
    xnor g10093 ( n9867 , n7100 , n9714 );
    xnor g10094 ( n208 , n10399 , n1426 );
    and g10095 ( n11095 , n4549 , n8215 );
    xnor g10096 ( n4904 , n1131 , n11159 );
    xnor g10097 ( n8927 , n8171 , n11111 );
    and g10098 ( n4521 , n9784 , n6920 );
    xnor g10099 ( n5108 , n12405 , n3415 );
    or g10100 ( n11396 , n4911 , n3911 );
    and g10101 ( n4275 , n1333 , n9195 );
    not g10102 ( n11262 , n12541 );
    xnor g10103 ( n861 , n51 , n3764 );
    xnor g10104 ( n3894 , n6591 , n10653 );
    nor g10105 ( n99 , n4658 , n2723 );
    and g10106 ( n12808 , n7620 , n1724 );
    or g10107 ( n9107 , n2099 , n5326 );
    xnor g10108 ( n10430 , n10135 , n4632 );
    and g10109 ( n2990 , n2848 , n3695 );
    xnor g10110 ( n6813 , n5500 , n393 );
    xnor g10111 ( n10209 , n10556 , n7390 );
    xnor g10112 ( n4673 , n1807 , n6477 );
    or g10113 ( n9624 , n2544 , n9477 );
    and g10114 ( n9550 , n12026 , n6104 );
    and g10115 ( n8024 , n10135 , n9854 );
    xnor g10116 ( n1244 , n2097 , n8794 );
    or g10117 ( n8318 , n6819 , n3191 );
    xnor g10118 ( n8709 , n284 , n5010 );
    or g10119 ( n8038 , n4403 , n8198 );
    and g10120 ( n11779 , n9632 , n9210 );
    nor g10121 ( n3789 , n5189 , n7960 );
    xnor g10122 ( n9999 , n9729 , n1690 );
    or g10123 ( n1119 , n7839 , n5540 );
    or g10124 ( n11214 , n2774 , n1617 );
    or g10125 ( n10620 , n5328 , n7647 );
    and g10126 ( n7330 , n9352 , n11275 );
    xnor g10127 ( n6907 , n10592 , n216 );
    nor g10128 ( n9893 , n1672 , n8513 );
    and g10129 ( n8117 , n3833 , n11418 );
    xnor g10130 ( n9791 , n6086 , n2356 );
    xnor g10131 ( n6842 , n10387 , n3019 );
    or g10132 ( n5621 , n3096 , n995 );
    and g10133 ( n8160 , n1344 , n11207 );
    and g10134 ( n4212 , n9536 , n6755 );
    xnor g10135 ( n10151 , n621 , n6844 );
    or g10136 ( n2229 , n1560 , n12132 );
    or g10137 ( n258 , n1183 , n8740 );
    or g10138 ( n9617 , n7914 , n4351 );
    or g10139 ( n10440 , n12729 , n552 );
    xnor g10140 ( n3484 , n4644 , n9531 );
    xnor g10141 ( n7956 , n1167 , n8971 );
    not g10142 ( n5131 , n461 );
    and g10143 ( n3947 , n5014 , n11938 );
    xnor g10144 ( n4019 , n7808 , n2306 );
    and g10145 ( n10409 , n10122 , n11428 );
    and g10146 ( n150 , n11153 , n9763 );
    not g10147 ( n7382 , n12777 );
    or g10148 ( n8546 , n5809 , n1163 );
    xnor g10149 ( n980 , n4932 , n6550 );
    not g10150 ( n2446 , n5363 );
    xnor g10151 ( n9480 , n1313 , n5117 );
    and g10152 ( n5385 , n7927 , n5358 );
    xnor g10153 ( n9683 , n7718 , n1933 );
    and g10154 ( n1210 , n3986 , n10990 );
    or g10155 ( n7312 , n3746 , n6455 );
    or g10156 ( n9451 , n5902 , n4400 );
    and g10157 ( n7082 , n6257 , n8845 );
    not g10158 ( n11150 , n9284 );
    nor g10159 ( n5427 , n3970 , n1364 );
    xnor g10160 ( n11672 , n11109 , n11391 );
    or g10161 ( n11069 , n3096 , n7952 );
    xnor g10162 ( n11151 , n2129 , n7529 );
    or g10163 ( n339 , n10339 , n4913 );
    or g10164 ( n8366 , n8354 , n8109 );
    or g10165 ( n157 , n2160 , n8725 );
    not g10166 ( n4778 , n7690 );
    not g10167 ( n2260 , n7783 );
    or g10168 ( n5084 , n7310 , n11202 );
    nor g10169 ( n12252 , n5014 , n11938 );
    xnor g10170 ( n12264 , n12010 , n7886 );
    not g10171 ( n10854 , n7733 );
    and g10172 ( n7969 , n3174 , n12043 );
    or g10173 ( n7490 , n2099 , n10854 );
    or g10174 ( n11596 , n4778 , n3924 );
    or g10175 ( n9740 , n5159 , n2304 );
    xnor g10176 ( n8179 , n9206 , n293 );
    xnor g10177 ( n2084 , n5516 , n8517 );
    not g10178 ( n2845 , n5909 );
    not g10179 ( n4471 , n7276 );
    or g10180 ( n10434 , n1937 , n7952 );
    and g10181 ( n6575 , n8040 , n4677 );
    and g10182 ( n12778 , n8560 , n4532 );
    not g10183 ( n4642 , n2749 );
    xnor g10184 ( n9691 , n2443 , n3391 );
    and g10185 ( n4666 , n10838 , n3060 );
    and g10186 ( n849 , n5422 , n7885 );
    or g10187 ( n1908 , n991 , n354 );
    xnor g10188 ( n1497 , n6452 , n8226 );
    or g10189 ( n11090 , n7474 , n1681 );
    and g10190 ( n4665 , n320 , n8869 );
    or g10191 ( n6482 , n10504 , n6682 );
    or g10192 ( n5889 , n3096 , n12816 );
    or g10193 ( n11729 , n5945 , n11820 );
    or g10194 ( n3452 , n752 , n2589 );
    or g10195 ( n8584 , n4911 , n4400 );
    xnor g10196 ( n6725 , n5639 , n11146 );
    or g10197 ( n1580 , n1699 , n1163 );
    or g10198 ( n1811 , n5915 , n12080 );
    nor g10199 ( n6930 , n9744 , n3963 );
    not g10200 ( n8673 , n9199 );
    or g10201 ( n76 , n6669 , n3568 );
    or g10202 ( n321 , n8692 , n2421 );
    xnor g10203 ( n12077 , n3559 , n11725 );
    and g10204 ( n5941 , n12752 , n1425 );
    and g10205 ( n5193 , n4660 , n4399 );
    xnor g10206 ( n10287 , n2526 , n9331 );
    not g10207 ( n9699 , n11108 );
    or g10208 ( n3669 , n2157 , n8245 );
    not g10209 ( n9078 , n12704 );
    and g10210 ( n1185 , n5964 , n2585 );
    not g10211 ( n3013 , n2771 );
    or g10212 ( n7401 , n12119 , n5468 );
    nor g10213 ( n10812 , n6415 , n2871 );
    or g10214 ( n10745 , n8959 , n11820 );
    or g10215 ( n1107 , n7251 , n4264 );
    not g10216 ( n12559 , n9353 );
    or g10217 ( n9997 , n989 , n5497 );
    xnor g10218 ( n10496 , n12463 , n3197 );
    or g10219 ( n6189 , n6718 , n12771 );
    xnor g10220 ( n6549 , n3334 , n2580 );
    not g10221 ( n6138 , n11999 );
    and g10222 ( n955 , n2727 , n2735 );
    not g10223 ( n7704 , n384 );
    xnor g10224 ( n941 , n289 , n11681 );
    xnor g10225 ( n6081 , n8213 , n12073 );
    or g10226 ( n7530 , n10835 , n795 );
    xnor g10227 ( n9552 , n11702 , n4296 );
    nor g10228 ( n5623 , n11362 , n2314 );
    or g10229 ( n7439 , n3620 , n5718 );
    xnor g10230 ( n1904 , n2326 , n10869 );
    not g10231 ( n476 , n12466 );
    or g10232 ( n5452 , n5438 , n11986 );
    or g10233 ( n6516 , n3096 , n7876 );
    or g10234 ( n7513 , n4498 , n2358 );
    and g10235 ( n1088 , n8574 , n8739 );
    xnor g10236 ( n1940 , n5830 , n6232 );
    xnor g10237 ( n11215 , n3844 , n3360 );
    not g10238 ( n12510 , n11395 );
    and g10239 ( n1752 , n1315 , n2211 );
    and g10240 ( n10167 , n10671 , n4295 );
    and g10241 ( n5338 , n1686 , n2898 );
    xnor g10242 ( n10583 , n8117 , n4976 );
    or g10243 ( n4635 , n3820 , n9568 );
    xnor g10244 ( n2619 , n8357 , n3670 );
    xnor g10245 ( n3502 , n7936 , n8298 );
    and g10246 ( n7619 , n2326 , n10869 );
    not g10247 ( n3306 , n12265 );
    and g10248 ( n2640 , n5558 , n316 );
    nor g10249 ( n10507 , n1815 , n6225 );
    xnor g10250 ( n1098 , n3780 , n11357 );
    xnor g10251 ( n1880 , n3170 , n11583 );
    xnor g10252 ( n2117 , n4756 , n2323 );
    or g10253 ( n9524 , n12361 , n1413 );
    or g10254 ( n632 , n3771 , n3302 );
    and g10255 ( n9270 , n3318 , n2675 );
    and g10256 ( n6422 , n2136 , n10652 );
    not g10257 ( n1932 , n533 );
    not g10258 ( n9639 , n5317 );
    and g10259 ( n2485 , n12786 , n5687 );
    xnor g10260 ( n8471 , n4850 , n8016 );
    xnor g10261 ( n1501 , n9385 , n12529 );
    or g10262 ( n11540 , n10157 , n8285 );
    or g10263 ( n5279 , n1937 , n9741 );
    or g10264 ( n11158 , n1434 , n4887 );
    nor g10265 ( n4066 , n4753 , n4851 );
    xnor g10266 ( n4259 , n4126 , n12608 );
    and g10267 ( n1822 , n10344 , n8541 );
    or g10268 ( n3605 , n5605 , n3745 );
    xnor g10269 ( n2143 , n5880 , n3243 );
    xnor g10270 ( n5255 , n11846 , n7117 );
    or g10271 ( n4641 , n12322 , n10872 );
    not g10272 ( n12631 , n585 );
    and g10273 ( n12493 , n4692 , n4977 );
    and g10274 ( n1252 , n1646 , n11866 );
    xnor g10275 ( n4496 , n7408 , n3547 );
    or g10276 ( n6691 , n10991 , n6056 );
    nor g10277 ( n11100 , n4783 , n8840 );
    and g10278 ( n12038 , n3822 , n1071 );
    xnor g10279 ( n3928 , n4320 , n1840 );
    xnor g10280 ( n863 , n2514 , n12097 );
    xnor g10281 ( n2275 , n768 , n10131 );
    or g10282 ( n12521 , n8251 , n6109 );
    or g10283 ( n1068 , n2649 , n9926 );
    xnor g10284 ( n2140 , n1317 , n4386 );
    or g10285 ( n1341 , n1941 , n9741 );
    or g10286 ( n4387 , n752 , n8768 );
    or g10287 ( n1011 , n589 , n12321 );
    not g10288 ( n827 , n7672 );
    xnor g10289 ( n6956 , n10802 , n1122 );
    xnor g10290 ( n7740 , n2958 , n11663 );
    or g10291 ( n12675 , n9544 , n9882 );
    xnor g10292 ( n5741 , n6917 , n990 );
    xnor g10293 ( n6536 , n7806 , n519 );
    xnor g10294 ( n10554 , n10548 , n1579 );
    not g10295 ( n7723 , n6665 );
    xnor g10296 ( n6717 , n9591 , n10044 );
    nor g10297 ( n6446 , n2248 , n5854 );
    or g10298 ( n5949 , n10338 , n6123 );
    xnor g10299 ( n11564 , n10723 , n10858 );
    xnor g10300 ( n11909 , n7291 , n9523 );
    and g10301 ( n10733 , n4219 , n1817 );
    not g10302 ( n7586 , n3372 );
    and g10303 ( n4580 , n3534 , n11350 );
    xnor g10304 ( n8547 , n9547 , n3194 );
    not g10305 ( n7357 , n4554 );
    or g10306 ( n7453 , n6231 , n3444 );
    not g10307 ( n5583 , n2161 );
    and g10308 ( n9385 , n2827 , n6170 );
    or g10309 ( n1475 , n9389 , n1162 );
    or g10310 ( n7860 , n7883 , n1595 );
    or g10311 ( n6732 , n11087 , n7183 );
    xnor g10312 ( n9435 , n6178 , n6494 );
    xnor g10313 ( n2 , n548 , n10859 );
    or g10314 ( n8388 , n2022 , n514 );
    or g10315 ( n4217 , n4778 , n4913 );
    or g10316 ( n4586 , n11307 , n1550 );
    nor g10317 ( n5951 , n8853 , n9941 );
    and g10318 ( n12225 , n347 , n5560 );
    not g10319 ( n5158 , n6872 );
    or g10320 ( n9141 , n752 , n3356 );
    not g10321 ( n8791 , n2469 );
    and g10322 ( n10395 , n3345 , n2925 );
    xnor g10323 ( n3243 , n1493 , n4216 );
    or g10324 ( n6098 , n11958 , n5538 );
    or g10325 ( n2164 , n12237 , n1163 );
    xnor g10326 ( n11806 , n11198 , n12166 );
    xnor g10327 ( n11404 , n9652 , n1766 );
    nor g10328 ( n7581 , n1036 , n11520 );
    not g10329 ( n1222 , n1251 );
    xnor g10330 ( n11504 , n7434 , n8063 );
    not g10331 ( n8187 , n6770 );
    or g10332 ( n3730 , n1508 , n9862 );
    not g10333 ( n511 , n2128 );
    xnor g10334 ( n9703 , n11512 , n5065 );
    xnor g10335 ( n4679 , n718 , n7454 );
    xnor g10336 ( n4083 , n7171 , n1999 );
    and g10337 ( n12484 , n1955 , n7008 );
    or g10338 ( n9408 , n10506 , n7060 );
    xnor g10339 ( n10154 , n3920 , n11164 );
    not g10340 ( n12067 , n866 );
    nor g10341 ( n10346 , n6995 , n2405 );
    and g10342 ( n1945 , n11097 , n2935 );
    or g10343 ( n9661 , n4838 , n12102 );
    and g10344 ( n8008 , n582 , n11014 );
    or g10345 ( n6686 , n10196 , n4875 );
    and g10346 ( n8157 , n5235 , n433 );
    or g10347 ( n2699 , n8583 , n10916 );
    or g10348 ( n3147 , n4632 , n8024 );
    nor g10349 ( n9927 , n6167 , n8883 );
    not g10350 ( n9584 , n4817 );
    and g10351 ( n9513 , n12318 , n6900 );
    xnor g10352 ( n3289 , n11674 , n7111 );
    and g10353 ( n11439 , n1186 , n12849 );
    nor g10354 ( n7542 , n3964 , n1334 );
    xnor g10355 ( n10368 , n4362 , n5115 );
    or g10356 ( n9483 , n12395 , n11818 );
    or g10357 ( n958 , n1539 , n3911 );
    or g10358 ( n3168 , n8127 , n6389 );
    xnor g10359 ( n9254 , n12262 , n8253 );
    not g10360 ( n1422 , n9891 );
    or g10361 ( n9825 , n3096 , n9741 );
    and g10362 ( n3607 , n10912 , n6143 );
    xnor g10363 ( n10540 , n9379 , n5110 );
    nor g10364 ( n11992 , n7383 , n4893 );
    or g10365 ( n5833 , n8026 , n3356 );
    nor g10366 ( n11937 , n5318 , n1327 );
    and g10367 ( n1096 , n2064 , n5122 );
    xnor g10368 ( n9854 , n2695 , n9302 );
    or g10369 ( n9022 , n8026 , n5012 );
    or g10370 ( n525 , n8966 , n3960 );
    or g10371 ( n1789 , n9878 , n1163 );
    not g10372 ( n9030 , n9485 );
    and g10373 ( n11354 , n5283 , n2802 );
    xnor g10374 ( n9463 , n7342 , n9839 );
    not g10375 ( n6031 , n1655 );
    xnor g10376 ( n10669 , n9849 , n2664 );
    and g10377 ( n7726 , n1962 , n3147 );
    xnor g10378 ( n7289 , n6339 , n10539 );
    or g10379 ( n9007 , n7933 , n10989 );
    or g10380 ( n4042 , n12503 , n28 );
    not g10381 ( n11949 , n5598 );
    or g10382 ( n3091 , n8344 , n1756 );
    xnor g10383 ( n11724 , n7592 , n2775 );
    not g10384 ( n1278 , n7685 );
    or g10385 ( n2165 , n2862 , n8865 );
    or g10386 ( n11106 , n9370 , n7246 );
    or g10387 ( n12458 , n12642 , n12185 );
    or g10388 ( n9250 , n9170 , n7341 );
    xnor g10389 ( n10415 , n2619 , n4978 );
    xnor g10390 ( n3661 , n7051 , n12323 );
    and g10391 ( n3891 , n8880 , n12629 );
    or g10392 ( n481 , n12797 , n12816 );
    not g10393 ( n5724 , n8381 );
    xnor g10394 ( n352 , n3534 , n10914 );
    nor g10395 ( n12907 , n8562 , n11642 );
    or g10396 ( n12841 , n752 , n10903 );
    not g10397 ( n7876 , n6703 );
    or g10398 ( n4858 , n2031 , n650 );
    xnor g10399 ( n11317 , n1304 , n7767 );
    not g10400 ( n5515 , n1139 );
    xnor g10401 ( n7399 , n526 , n3690 );
    xnor g10402 ( n4123 , n9317 , n12645 );
    and g10403 ( n1759 , n5599 , n7256 );
    nor g10404 ( n1617 , n10647 , n7422 );
    or g10405 ( n11744 , n11026 , n9144 );
    and g10406 ( n4746 , n76 , n9323 );
    and g10407 ( n6150 , n200 , n6906 );
    xnor g10408 ( n4949 , n701 , n7036 );
    or g10409 ( n8634 , n10142 , n11746 );
    not g10410 ( n2349 , n10762 );
    not g10411 ( n5979 , n12657 );
    or g10412 ( n12263 , n2217 , n3606 );
    or g10413 ( n2130 , n12186 , n6169 );
    xnor g10414 ( n7079 , n8606 , n170 );
    xnor g10415 ( n4918 , n882 , n11209 );
    xnor g10416 ( n1810 , n4701 , n6811 );
    and g10417 ( n188 , n11015 , n12578 );
    not g10418 ( n6941 , n12712 );
    not g10419 ( n8426 , n3722 );
    xnor g10420 ( n263 , n3503 , n11139 );
    or g10421 ( n4901 , n131 , n1228 );
    or g10422 ( n11202 , n636 , n8740 );
    not g10423 ( n11163 , n7878 );
    xnor g10424 ( n2452 , n5595 , n8170 );
    or g10425 ( n10351 , n1695 , n8066 );
    or g10426 ( n3067 , n12361 , n6455 );
    xnor g10427 ( n821 , n4257 , n20 );
    xnor g10428 ( n12153 , n2730 , n10316 );
    xnor g10429 ( n2181 , n11956 , n1168 );
    or g10430 ( n4153 , n8428 , n1413 );
    not g10431 ( n765 , n11489 );
    or g10432 ( n3726 , n7410 , n3763 );
    xnor g10433 ( n12570 , n144 , n7137 );
    or g10434 ( n10088 , n7899 , n5485 );
    or g10435 ( n2694 , n4498 , n4242 );
    or g10436 ( n10353 , n749 , n8676 );
    or g10437 ( n4721 , n6977 , n1413 );
    or g10438 ( n4166 , n7391 , n10419 );
    xnor g10439 ( n5293 , n1322 , n2565 );
    xnor g10440 ( n5910 , n7428 , n1113 );
    or g10441 ( n10318 , n7449 , n7921 );
    xnor g10442 ( n7405 , n10783 , n12039 );
    not g10443 ( n3614 , n557 );
    not g10444 ( n1025 , n10336 );
    not g10445 ( n5258 , n11791 );
    or g10446 ( n4101 , n9413 , n9022 );
    not g10447 ( n5575 , n6877 );
    nor g10448 ( n3539 , n1945 , n3972 );
    not g10449 ( n11115 , n5459 );
    or g10450 ( n2800 , n182 , n6267 );
    xnor g10451 ( n2246 , n797 , n12169 );
    xnor g10452 ( n5863 , n9798 , n11404 );
    xnor g10453 ( n10375 , n5681 , n4819 );
    or g10454 ( n5377 , n8527 , n11948 );
    xnor g10455 ( n1867 , n3384 , n2550 );
    xnor g10456 ( n1480 , n10172 , n8119 );
    xnor g10457 ( n7516 , n3752 , n2920 );
    or g10458 ( n3870 , n2834 , n10526 );
    xnor g10459 ( n7880 , n357 , n5306 );
    and g10460 ( n8660 , n11478 , n5645 );
    xnor g10461 ( n9240 , n12741 , n4229 );
    or g10462 ( n10739 , n2763 , n789 );
    and g10463 ( n2736 , n8514 , n7406 );
    nor g10464 ( n12375 , n9825 , n8469 );
    or g10465 ( n4209 , n10511 , n484 );
    xnor g10466 ( n10393 , n1274 , n6492 );
    not g10467 ( n200 , n10265 );
    or g10468 ( n8347 , n2456 , n8648 );
    xnor g10469 ( n12523 , n3706 , n2625 );
    not g10470 ( n3344 , n6575 );
    xnor g10471 ( n2218 , n1751 , n4178 );
    or g10472 ( n1238 , n11446 , n9084 );
    nor g10473 ( n2767 , n12266 , n10337 );
    xnor g10474 ( n12910 , n3492 , n698 );
    or g10475 ( n1817 , n9228 , n10931 );
    or g10476 ( n1992 , n8026 , n6084 );
    xnor g10477 ( n1513 , n1675 , n344 );
    nor g10478 ( n12300 , n10033 , n11823 );
    or g10479 ( n4500 , n4911 , n1851 );
    and g10480 ( n4583 , n1052 , n266 );
    xnor g10481 ( n5653 , n10847 , n12626 );
    or g10482 ( n11335 , n3743 , n11698 );
    or g10483 ( n5816 , n10202 , n9729 );
    not g10484 ( n8479 , n6766 );
    not g10485 ( n9963 , n8628 );
    xnor g10486 ( n8198 , n7777 , n11872 );
    nor g10487 ( n5843 , n12516 , n720 );
    or g10488 ( n4660 , n2552 , n6974 );
    xnor g10489 ( n9766 , n8567 , n341 );
    or g10490 ( n9720 , n12755 , n9954 );
    xnor g10491 ( n7931 , n3046 , n7201 );
    and g10492 ( n4468 , n4414 , n3781 );
    xnor g10493 ( n9898 , n5155 , n1860 );
    not g10494 ( n424 , n720 );
    not g10495 ( n2552 , n10973 );
    and g10496 ( n9130 , n8629 , n1498 );
    xnor g10497 ( n465 , n3642 , n7601 );
    xnor g10498 ( n5085 , n7383 , n12914 );
    not g10499 ( n4040 , n390 );
    xnor g10500 ( n11256 , n2110 , n11776 );
    xnor g10501 ( n620 , n3442 , n2694 );
    or g10502 ( n11013 , n8552 , n8655 );
    and g10503 ( n8580 , n3303 , n1744 );
    or g10504 ( n8955 , n1183 , n4913 );
    xnor g10505 ( n8802 , n1123 , n3729 );
    or g10506 ( n10506 , n9373 , n4654 );
    and g10507 ( n9166 , n7310 , n11202 );
    xnor g10508 ( n12128 , n7554 , n9792 );
    or g10509 ( n12488 , n9977 , n4375 );
    and g10510 ( n9779 , n11825 , n10592 );
    and g10511 ( n7053 , n11902 , n6883 );
    nor g10512 ( n818 , n4401 , n9629 );
    not g10513 ( n9259 , n8418 );
    not g10514 ( n10419 , n5320 );
    and g10515 ( n6070 , n11592 , n12419 );
    and g10516 ( n3208 , n9625 , n5937 );
    or g10517 ( n6247 , n5423 , n1528 );
    nor g10518 ( n979 , n7940 , n818 );
    and g10519 ( n7773 , n2499 , n5418 );
    or g10520 ( n4561 , n12119 , n5326 );
    or g10521 ( n3497 , n4694 , n2768 );
    or g10522 ( n1859 , n7839 , n12816 );
    nor g10523 ( n7314 , n10850 , n9605 );
    xnor g10524 ( n722 , n4390 , n7748 );
    and g10525 ( n3601 , n2464 , n11023 );
    or g10526 ( n7218 , n6636 , n12215 );
    and g10527 ( n11297 , n107 , n10880 );
    or g10528 ( n4845 , n4354 , n11639 );
    or g10529 ( n11854 , n3082 , n2875 );
    and g10530 ( n3509 , n527 , n9816 );
    xnor g10531 ( n8931 , n12622 , n3919 );
    xnor g10532 ( n4886 , n9222 , n5162 );
    or g10533 ( n6546 , n1086 , n123 );
    and g10534 ( n6848 , n2236 , n3277 );
    or g10535 ( n5607 , n4778 , n8109 );
    or g10536 ( n2848 , n7774 , n7127 );
    and g10537 ( n383 , n1887 , n7903 );
    not g10538 ( n7190 , n4612 );
    and g10539 ( n9669 , n656 , n10580 );
    xnor g10540 ( n4631 , n8348 , n111 );
    or g10541 ( n678 , n3243 , n5880 );
    and g10542 ( n9194 , n6621 , n10910 );
    or g10543 ( n4433 , n284 , n10693 );
    xnor g10544 ( n3094 , n8577 , n8249 );
    and g10545 ( n12 , n8412 , n3521 );
    xnor g10546 ( n723 , n4821 , n48 );
    xnor g10547 ( n12336 , n3232 , n5997 );
    nor g10548 ( n12134 , n7305 , n8872 );
    not g10549 ( n125 , n1948 );
    xnor g10550 ( n3663 , n10116 , n4679 );
    not g10551 ( n8768 , n10439 );
    xnor g10552 ( n764 , n634 , n11178 );
    or g10553 ( n4707 , n3772 , n4171 );
    xnor g10554 ( n10321 , n3799 , n4590 );
    xnor g10555 ( n9928 , n8584 , n7644 );
    xnor g10556 ( n9406 , n11839 , n12876 );
    xnor g10557 ( n5905 , n8455 , n6891 );
    not g10558 ( n7962 , n2015 );
    or g10559 ( n2930 , n9428 , n9981 );
    and g10560 ( n3042 , n11182 , n4200 );
    xnor g10561 ( n3697 , n2819 , n11830 );
    nor g10562 ( n2723 , n2787 , n1208 );
    or g10563 ( n1972 , n11281 , n4629 );
    or g10564 ( n5345 , n8959 , n7876 );
    xnor g10565 ( n12405 , n4715 , n6503 );
    and g10566 ( n6683 , n1471 , n11876 );
    or g10567 ( n6934 , n10738 , n3150 );
    or g10568 ( n4926 , n5915 , n12535 );
    xor g10569 ( n12314 , n9564 , n7680 );
    or g10570 ( n2125 , n6697 , n12225 );
    xnor g10571 ( n9157 , n2976 , n11495 );
    and g10572 ( n2473 , n2188 , n8006 );
    or g10573 ( n5064 , n11958 , n11820 );
    not g10574 ( n12768 , n8504 );
    or g10575 ( n7383 , n10142 , n7389 );
    nor g10576 ( n5139 , n11178 , n634 );
    and g10577 ( n1153 , n9273 , n11048 );
    and g10578 ( n12605 , n5214 , n2616 );
    xnor g10579 ( n7695 , n12144 , n3153 );
    and g10580 ( n7561 , n11165 , n352 );
    xnor g10581 ( n10786 , n12325 , n7556 );
    or g10582 ( n3345 , n8704 , n5761 );
    xnor g10583 ( n10143 , n5412 , n12255 );
    or g10584 ( n10200 , n12416 , n9961 );
    not g10585 ( n6106 , n3499 );
    and g10586 ( n879 , n326 , n2904 );
    xnor g10587 ( n9923 , n10788 , n8523 );
    and g10588 ( n4323 , n4667 , n6199 );
    xnor g10589 ( n8379 , n4984 , n1153 );
    xnor g10590 ( n223 , n5627 , n1770 );
    not g10591 ( n11226 , n2418 );
    nor g10592 ( n6100 , n11378 , n11991 );
    or g10593 ( n441 , n12267 , n12890 );
    nor g10594 ( n1585 , n3386 , n129 );
    not g10595 ( n9853 , n6618 );
    or g10596 ( n3691 , n8699 , n228 );
    and g10597 ( n7328 , n6219 , n4959 );
    or g10598 ( n10197 , n1539 , n10066 );
    xnor g10599 ( n9027 , n10777 , n10171 );
    xnor g10600 ( n3769 , n6250 , n93 );
    xnor g10601 ( n10452 , n3972 , n4477 );
    or g10602 ( n10803 , n4911 , n1915 );
    xnor g10603 ( n9419 , n9567 , n5754 );
    and g10604 ( n8548 , n10265 , n11132 );
    xnor g10605 ( n6432 , n12618 , n10353 );
    xnor g10606 ( n8129 , n5606 , n7249 );
    or g10607 ( n0 , n3743 , n9568 );
    or g10608 ( n6484 , n5815 , n6018 );
    or g10609 ( n11083 , n1474 , n9633 );
    or g10610 ( n1081 , n792 , n2880 );
    nor g10611 ( n12618 , n10917 , n6238 );
    or g10612 ( n4441 , n2385 , n5803 );
    or g10613 ( n4356 , n3501 , n4924 );
    not g10614 ( n6524 , n6604 );
    not g10615 ( n2422 , n3384 );
    or g10616 ( n4867 , n12494 , n12719 );
    not g10617 ( n10625 , n2104 );
    or g10618 ( n5369 , n773 , n12405 );
    and g10619 ( n8025 , n12733 , n5820 );
    or g10620 ( n3140 , n191 , n2076 );
    or g10621 ( n11302 , n7918 , n544 );
    nor g10622 ( n434 , n12739 , n3108 );
    and g10623 ( n11375 , n12946 , n8265 );
    not g10624 ( n4140 , n6591 );
    or g10625 ( n1688 , n10835 , n28 );
    and g10626 ( n6255 , n11914 , n6839 );
    or g10627 ( n9134 , n636 , n9586 );
    xnor g10628 ( n5014 , n12564 , n8003 );
    or g10629 ( n426 , n3118 , n2203 );
    not g10630 ( n6388 , n11062 );
    xnor g10631 ( n5632 , n8442 , n4745 );
    or g10632 ( n3912 , n11588 , n5476 );
    and g10633 ( n3252 , n6095 , n781 );
    xnor g10634 ( n8043 , n6981 , n9149 );
    xnor g10635 ( n1046 , n9837 , n12126 );
    xnor g10636 ( n4260 , n2746 , n7887 );
    xnor g10637 ( n356 , n12882 , n11249 );
    not g10638 ( n12335 , n1577 );
    or g10639 ( n11739 , n11433 , n7952 );
    not g10640 ( n10962 , n2978 );
    not g10641 ( n9452 , n3833 );
    or g10642 ( n6001 , n3821 , n4701 );
    or g10643 ( n6078 , n5915 , n7382 );
    xnor g10644 ( n4438 , n9995 , n10754 );
    not g10645 ( n9148 , n3726 );
    and g10646 ( n11862 , n2071 , n10323 );
    xnor g10647 ( n272 , n377 , n1492 );
    not g10648 ( n5496 , n9016 );
    and g10649 ( n2878 , n3692 , n7649 );
    xnor g10650 ( n12620 , n61 , n8393 );
    xnor g10651 ( n4306 , n1543 , n1294 );
    not g10652 ( n4617 , n2665 );
    and g10653 ( n3968 , n11090 , n7010 );
    or g10654 ( n6468 , n4396 , n10296 );
    not g10655 ( n8432 , n5756 );
    or g10656 ( n6347 , n11958 , n10903 );
    xnor g10657 ( n4712 , n5812 , n5984 );
    and g10658 ( n12653 , n4433 , n2681 );
    and g10659 ( n8053 , n9241 , n7946 );
    nor g10660 ( n5958 , n158 , n9260 );
    xnor g10661 ( n7386 , n407 , n4006 );
    or g10662 ( n5414 , n989 , n7424 );
    xnor g10663 ( n5490 , n855 , n5190 );
    or g10664 ( n2322 , n3650 , n1285 );
    xnor g10665 ( n8495 , n9101 , n9516 );
    or g10666 ( n1877 , n12237 , n12686 );
    or g10667 ( n8686 , n5748 , n5639 );
    and g10668 ( n3558 , n5563 , n5749 );
    and g10669 ( n4554 , n4111 , n4215 );
    xnor g10670 ( n5169 , n11095 , n10087 );
    not g10671 ( n5415 , n5504 );
    and g10672 ( n9342 , n8851 , n6768 );
    nor g10673 ( n9146 , n1039 , n5611 );
    xnor g10674 ( n8545 , n7338 , n10267 );
    not g10675 ( n1077 , n9281 );
    xnor g10676 ( n10557 , n10230 , n10273 );
    or g10677 ( n3747 , n5530 , n9586 );
    xnor g10678 ( n11020 , n4254 , n5926 );
    nor g10679 ( n5847 , n8509 , n3099 );
    not g10680 ( n5431 , n6917 );
    xor g10681 ( n1055 , n4270 , n7579 );
    xnor g10682 ( n10789 , n3343 , n7849 );
    and g10683 ( n2771 , n7364 , n1843 );
    or g10684 ( n1325 , n4707 , n495 );
    xnor g10685 ( n9831 , n4838 , n5901 );
    and g10686 ( n9284 , n7768 , n2631 );
    and g10687 ( n4725 , n11773 , n7473 );
    xnor g10688 ( n2396 , n3050 , n11524 );
    xnor g10689 ( n4517 , n4577 , n4887 );
    and g10690 ( n436 , n1664 , n6851 );
    not g10691 ( n6055 , n4806 );
    xnor g10692 ( n1016 , n3419 , n4610 );
    or g10693 ( n10578 , n2081 , n4068 );
    or g10694 ( n11471 , n9170 , n1915 );
    and g10695 ( n7497 , n4124 , n11935 );
    and g10696 ( n2318 , n11779 , n2256 );
    xnor g10697 ( n10160 , n555 , n6841 );
    or g10698 ( n7752 , n9170 , n11827 );
    and g10699 ( n4600 , n8607 , n371 );
    or g10700 ( n789 , n4059 , n3911 );
    nor g10701 ( n12143 , n1651 , n12695 );
    xnor g10702 ( n10650 , n8277 , n9724 );
    not g10703 ( n8543 , n2954 );
    xnor g10704 ( n5300 , n12293 , n5833 );
    and g10705 ( n6913 , n11470 , n7264 );
    and g10706 ( n333 , n1099 , n11183 );
    and g10707 ( n5688 , n1619 , n3477 );
    or g10708 ( n8739 , n9366 , n3709 );
    or g10709 ( n11580 , n4787 , n1889 );
    and g10710 ( n5234 , n6151 , n11219 );
    and g10711 ( n11362 , n2446 , n11631 );
    not g10712 ( n7952 , n1209 );
    or g10713 ( n6049 , n4059 , n1738 );
    nor g10714 ( n8707 , n6628 , n11372 );
    nor g10715 ( n1474 , n7459 , n4490 );
    or g10716 ( n11033 , n7777 , n11872 );
    xnor g10717 ( n6424 , n7182 , n5905 );
    or g10718 ( n3776 , n7041 , n2932 );
    xnor g10719 ( n6987 , n10865 , n8849 );
    and g10720 ( n11058 , n8704 , n5761 );
    or g10721 ( n9801 , n1937 , n11775 );
    nor g10722 ( n1801 , n12027 , n10176 );
    and g10723 ( n2044 , n11846 , n7117 );
    or g10724 ( n1257 , n4552 , n12184 );
    and g10725 ( n3332 , n2946 , n7488 );
    xnor g10726 ( n11464 , n5089 , n10823 );
    and g10727 ( n7545 , n9492 , n4420 );
    nor g10728 ( n2075 , n5650 , n11675 );
    nor g10729 ( n136 , n8140 , n9877 );
    xnor g10730 ( n1427 , n8531 , n11985 );
    or g10731 ( n3963 , n994 , n1738 );
    xnor g10732 ( n4263 , n3971 , n10897 );
    xnor g10733 ( n1136 , n4587 , n4975 );
    xnor g10734 ( n6947 , n11115 , n3320 );
    xnor g10735 ( n1597 , n11052 , n7719 );
    not g10736 ( n12120 , n7270 );
    and g10737 ( n3902 , n2040 , n1605 );
    xnor g10738 ( n1792 , n7609 , n7907 );
    or g10739 ( n12638 , n1728 , n7627 );
    not g10740 ( n7338 , n5081 );
    nor g10741 ( n4383 , n8714 , n9608 );
    xnor g10742 ( n4732 , n8491 , n10287 );
    and g10743 ( n7498 , n1677 , n6235 );
    and g10744 ( n7337 , n10566 , n6730 );
    not g10745 ( n5266 , n2650 );
    or g10746 ( n1386 , n5448 , n932 );
    not g10747 ( n11750 , n5233 );
    or g10748 ( n9271 , n10835 , n1476 );
    or g10749 ( n2720 , n8354 , n10854 );
    or g10750 ( n4420 , n3096 , n2815 );
    nor g10751 ( n8224 , n237 , n4556 );
    xnor g10752 ( n4329 , n2011 , n6268 );
    not g10753 ( n11742 , n2571 );
    xnor g10754 ( n2323 , n4552 , n12011 );
    xnor g10755 ( n12209 , n9695 , n10708 );
    and g10756 ( n302 , n967 , n6615 );
    xnor g10757 ( n4484 , n5391 , n11320 );
    not g10758 ( n5691 , n1878 );
    not g10759 ( n8554 , n3070 );
    nor g10760 ( n2821 , n8124 , n5367 );
    or g10761 ( n12522 , n7709 , n4527 );
    or g10762 ( n6765 , n1715 , n11329 );
    or g10763 ( n1574 , n2071 , n10323 );
    or g10764 ( n6075 , n9170 , n1455 );
    not g10765 ( n6290 , n2109 );
    nor g10766 ( n10679 , n9967 , n7357 );
    nor g10767 ( n5056 , n9598 , n4395 );
    or g10768 ( n10992 , n3127 , n1455 );
    xnor g10769 ( n2481 , n12112 , n12364 );
    and g10770 ( n6140 , n12216 , n10672 );
    or g10771 ( n7747 , n4728 , n10505 );
    and g10772 ( n12337 , n12271 , n12707 );
    or g10773 ( n831 , n6685 , n8604 );
    not g10774 ( n7508 , n8018 );
    xnor g10775 ( n9443 , n12783 , n12943 );
    xnor g10776 ( n772 , n4506 , n345 );
    xnor g10777 ( n10476 , n12573 , n1610 );
    xnor g10778 ( n7013 , n2641 , n11574 );
    not g10779 ( n665 , n12540 );
    xnor g10780 ( n7248 , n12338 , n2528 );
    xnor g10781 ( n8206 , n10178 , n9727 );
    and g10782 ( n10013 , n587 , n12665 );
    or g10783 ( n3901 , n994 , n11430 );
    not g10784 ( n11138 , n11393 );
    not g10785 ( n8755 , n11687 );
    or g10786 ( n12700 , n11433 , n6455 );
    xnor g10787 ( n2553 , n7590 , n10490 );
    not g10788 ( n569 , n1037 );
    xnor g10789 ( n5476 , n11614 , n7152 );
    xnor g10790 ( n8934 , n3319 , n516 );
    or g10791 ( n5141 , n4873 , n11880 );
    xnor g10792 ( n12564 , n10181 , n10126 );
    or g10793 ( n7855 , n10471 , n9765 );
    xnor g10794 ( n4069 , n11001 , n6528 );
    nor g10795 ( n1927 , n4367 , n119 );
    or g10796 ( n6697 , n3743 , n4642 );
    or g10797 ( n10960 , n6373 , n1047 );
    and g10798 ( n2015 , n4466 , n9793 );
    nor g10799 ( n8155 , n9274 , n10814 );
    and g10800 ( n7486 , n2260 , n2454 );
    xnor g10801 ( n10994 , n11879 , n7655 );
    xnor g10802 ( n662 , n6725 , n9344 );
    or g10803 ( n7939 , n2456 , n5781 );
    or g10804 ( n5200 , n8552 , n1932 );
    and g10805 ( n10998 , n12025 , n11407 );
    not g10806 ( n9455 , n5164 );
    and g10807 ( n3414 , n9617 , n139 );
    or g10808 ( n11524 , n7449 , n1509 );
    xnor g10809 ( n5333 , n60 , n11213 );
    not g10810 ( n8127 , n11821 );
    and g10811 ( n2413 , n137 , n2802 );
    or g10812 ( n926 , n5345 , n5711 );
    xnor g10813 ( n7849 , n1890 , n6436 );
    nor g10814 ( n10930 , n4855 , n6753 );
    and g10815 ( n8675 , n6551 , n2086 );
    not g10816 ( n1383 , n6056 );
    xnor g10817 ( n6609 , n12716 , n10524 );
    xnor g10818 ( n9629 , n10453 , n7597 );
    not g10819 ( n1509 , n10848 );
    xnor g10820 ( n8843 , n10579 , n1888 );
    or g10821 ( n4750 , n8870 , n10854 );
    or g10822 ( n10564 , n8051 , n3966 );
    not g10823 ( n9885 , n3194 );
    or g10824 ( n1952 , n3512 , n10293 );
    xnor g10825 ( n12793 , n991 , n5664 );
    and g10826 ( n9961 , n6368 , n1309 );
    xnor g10827 ( n9635 , n9231 , n6395 );
    and g10828 ( n3557 , n8810 , n318 );
    xnor g10829 ( n9424 , n4337 , n6558 );
    or g10830 ( n2529 , n9878 , n5326 );
    nor g10831 ( n2628 , n10756 , n3373 );
    xnor g10832 ( n10120 , n573 , n11044 );
    nor g10833 ( n9609 , n12234 , n7292 );
    nor g10834 ( n12590 , n3810 , n3181 );
    or g10835 ( n10882 , n5765 , n4654 );
    and g10836 ( n3949 , n11571 , n5511 );
    and g10837 ( n4539 , n6227 , n11129 );
    xnor g10838 ( n12011 , n1637 , n11325 );
    and g10839 ( n8600 , n12705 , n2509 );
    not g10840 ( n12406 , n2108 );
    nor g10841 ( n5005 , n680 , n2996 );
    nor g10842 ( n10046 , n5903 , n7119 );
    and g10843 ( n12757 , n8476 , n11967 );
    not g10844 ( n1831 , n12588 );
    xnor g10845 ( n400 , n1919 , n12615 );
    and g10846 ( n6157 , n4365 , n4323 );
    xnor g10847 ( n6174 , n4165 , n6878 );
    not g10848 ( n10856 , n11642 );
    xnor g10849 ( n5411 , n604 , n1329 );
    not g10850 ( n4308 , n11365 );
    xnor g10851 ( n2166 , n2452 , n11298 );
    and g10852 ( n342 , n10960 , n10315 );
    or g10853 ( n8002 , n752 , n11410 );
    not g10854 ( n4221 , n2364 );
    xnor g10855 ( n6751 , n769 , n3129 );
    and g10856 ( n4808 , n4841 , n6456 );
    and g10857 ( n6537 , n12365 , n11406 );
    xnor g10858 ( n9434 , n5640 , n6840 );
    or g10859 ( n6015 , n6718 , n8830 );
    xnor g10860 ( n11725 , n5410 , n460 );
    and g10861 ( n8049 , n12666 , n3624 );
    or g10862 ( n4647 , n6577 , n995 );
    and g10863 ( n9258 , n11518 , n878 );
    not g10864 ( n6634 , n12533 );
    and g10865 ( n10455 , n3687 , n532 );
    xnor g10866 ( n12354 , n450 , n11516 );
    and g10867 ( n5226 , n7630 , n5736 );
    or g10868 ( n12646 , n8405 , n3224 );
    xnor g10869 ( n1873 , n10637 , n12714 );
    or g10870 ( n12886 , n4167 , n6892 );
    xnor g10871 ( n248 , n8104 , n7934 );
    not g10872 ( n1189 , n4707 );
    and g10873 ( n8898 , n3810 , n3181 );
    or g10874 ( n284 , n7116 , n3903 );
    and g10875 ( n6872 , n11033 , n8038 );
    or g10876 ( n975 , n11719 , n5497 );
    xnor g10877 ( n5521 , n4120 , n10032 );
    or g10878 ( n11968 , n8428 , n7952 );
    or g10879 ( n6737 , n3773 , n12287 );
    and g10880 ( n10489 , n6436 , n7645 );
    or g10881 ( n10531 , n1937 , n6197 );
    xnor g10882 ( n10441 , n12303 , n6904 );
    xnor g10883 ( n285 , n3015 , n2294 );
    or g10884 ( n8377 , n4283 , n5524 );
    xnor g10885 ( n11632 , n11501 , n11188 );
    nor g10886 ( n9053 , n1503 , n2839 );
    not g10887 ( n3855 , n5973 );
    or g10888 ( n11625 , n5794 , n4340 );
    xnor g10889 ( n11705 , n5235 , n11927 );
    xnor g10890 ( n7568 , n1952 , n2092 );
    and g10891 ( n7009 , n9311 , n9534 );
    xnor g10892 ( n11614 , n7131 , n8807 );
    not g10893 ( n12304 , n8952 );
    not g10894 ( n4310 , n8486 );
    and g10895 ( n2144 , n1571 , n1422 );
    xnor g10896 ( n8928 , n12249 , n3613 );
    not g10897 ( n8644 , n5069 );
    xnor g10898 ( n6584 , n3125 , n11199 );
    not g10899 ( n9730 , n11352 );
    and g10900 ( n5684 , n8759 , n12709 );
    not g10901 ( n10122 , n12692 );
    and g10902 ( n10127 , n722 , n3987 );
    not g10903 ( n4113 , n1639 );
    xnor g10904 ( n3525 , n8221 , n5445 );
    xnor g10905 ( n1850 , n667 , n10978 );
    nor g10906 ( n6321 , n6222 , n3323 );
    or g10907 ( n6880 , n6577 , n7395 );
    xnor g10908 ( n7805 , n3163 , n8381 );
    xnor g10909 ( n8262 , n1241 , n492 );
    nor g10910 ( n5709 , n10381 , n6177 );
    or g10911 ( n3009 , n5945 , n5540 );
    xnor g10912 ( n2627 , n5776 , n10454 );
    not g10913 ( n9470 , n6799 );
    or g10914 ( n8924 , n9262 , n4527 );
    not g10915 ( n11429 , n10512 );
    nor g10916 ( n12695 , n12167 , n4774 );
    or g10917 ( n7713 , n10750 , n1932 );
    or g10918 ( n10502 , n10157 , n9568 );
    xnor g10919 ( n5947 , n5992 , n12384 );
    and g10920 ( n1464 , n2743 , n8597 );
    xnor g10921 ( n1933 , n5679 , n2963 );
    not g10922 ( n1938 , n5302 );
    or g10923 ( n10095 , n3425 , n7938 );
    or g10924 ( n7323 , n3681 , n7492 );
    not g10925 ( n10944 , n10059 );
    xnor g10926 ( n10852 , n7665 , n4557 );
    not g10927 ( n488 , n8015 );
    or g10928 ( n11700 , n1183 , n8655 );
    or g10929 ( n2459 , n2217 , n7921 );
    xnor g10930 ( n11096 , n4923 , n2693 );
    nor g10931 ( n9649 , n6649 , n542 );
    xnor g10932 ( n7360 , n11132 , n200 );
    or g10933 ( n2664 , n686 , n11775 );
    xnor g10934 ( n7454 , n5292 , n369 );
    or g10935 ( n9149 , n11923 , n7921 );
    nor g10936 ( n5629 , n12590 , n11035 );
    nor g10937 ( n7503 , n3808 , n8460 );
    or g10938 ( n5823 , n12237 , n826 );
    or g10939 ( n6772 , n2766 , n1770 );
    xor g10940 ( n3201 , n10290 , n3732 );
    xnor g10941 ( n10973 , n6899 , n8856 );
    xnor g10942 ( n2033 , n9712 , n7511 );
    or g10943 ( n507 , n4322 , n512 );
    not g10944 ( n5012 , n2024 );
    xnor g10945 ( n2432 , n12530 , n12779 );
    xnor g10946 ( n2382 , n6478 , n5973 );
    nor g10947 ( n2543 , n8307 , n3539 );
    or g10948 ( n431 , n8552 , n10422 );
    xnor g10949 ( n12181 , n10505 , n11441 );
    and g10950 ( n10493 , n11944 , n5389 );
    and g10951 ( n2706 , n4116 , n7188 );
    or g10952 ( n12725 , n1937 , n5538 );
    nor g10953 ( n9004 , n1987 , n3049 );
    nor g10954 ( n3490 , n1616 , n1002 );
    xnor g10955 ( n7600 , n2978 , n6507 );
    or g10956 ( n9520 , n11120 , n12373 );
    not g10957 ( n4623 , n10409 );
    or g10958 ( n8320 , n3617 , n9188 );
    or g10959 ( n738 , n3653 , n5764 );
    and g10960 ( n1755 , n2073 , n12028 );
    not g10961 ( n3353 , n7925 );
    xnor g10962 ( n6299 , n7292 , n4786 );
    or g10963 ( n6472 , n6577 , n8768 );
    or g10964 ( n4717 , n11552 , n9568 );
    not g10965 ( n8524 , n2577 );
    or g10966 ( n1347 , n5809 , n12535 );
    xnor g10967 ( n12060 , n9663 , n6623 );
    and g10968 ( n10283 , n12767 , n6780 );
    xnor g10969 ( n6492 , n3251 , n6134 );
    not g10970 ( n5915 , n2530 );
    or g10971 ( n9305 , n11887 , n5468 );
    or g10972 ( n3455 , n1708 , n12114 );
    or g10973 ( n5801 , n1183 , n7382 );
    xnor g10974 ( n11836 , n9223 , n9747 );
    and g10975 ( n2604 , n737 , n6132 );
    nor g10976 ( n11174 , n8308 , n6581 );
    xnor g10977 ( n3223 , n2182 , n11106 );
    or g10978 ( n3039 , n9196 , n8349 );
    and g10979 ( n1093 , n6398 , n9442 );
    not g10980 ( n3144 , n7327 );
    not g10981 ( n192 , n8053 );
    and g10982 ( n11050 , n5496 , n9603 );
    or g10983 ( n1242 , n7283 , n4400 );
    nor g10984 ( n4738 , n3140 , n3447 );
    or g10985 ( n8623 , n7293 , n1641 );
    and g10986 ( n4943 , n6098 , n1845 );
    and g10987 ( n2737 , n3767 , n7600 );
    xnor g10988 ( n9626 , n2759 , n16 );
    xnor g10989 ( n8121 , n6653 , n2956 );
    and g10990 ( n11849 , n1737 , n11299 );
    xnor g10991 ( n9569 , n8483 , n2495 );
    or g10992 ( n3549 , n7704 , n9671 );
    not g10993 ( n8643 , n217 );
    and g10994 ( n5093 , n5314 , n2749 );
    not g10995 ( n6457 , n2788 );
    nor g10996 ( n2841 , n9024 , n10201 );
    and g10997 ( n10834 , n12173 , n1405 );
    xnor g10998 ( n11628 , n308 , n1500 );
    not g10999 ( n331 , n6717 );
    or g11000 ( n4097 , n4904 , n701 );
    and g11001 ( n7276 , n5439 , n8083 );
    and g11002 ( n9255 , n3672 , n8255 );
    not g11003 ( n11880 , n6858 );
    or g11004 ( n11071 , n7839 , n11775 );
    xor g11005 ( n9955 , n10005 , n791 );
    xnor g11006 ( n1125 , n6974 , n5719 );
    and g11007 ( n3996 , n589 , n12321 );
    xnor g11008 ( n2177 , n7442 , n568 );
    not g11009 ( n12568 , n4257 );
    or g11010 ( n9538 , n7116 , n6455 );
    xnor g11011 ( n12834 , n5522 , n115 );
    nor g11012 ( n5743 , n2418 , n5274 );
    xnor g11013 ( n6978 , n2516 , n1064 );
    or g11014 ( n7292 , n627 , n11964 );
    or g11015 ( n12223 , n10142 , n8859 );
    not g11016 ( n1685 , n12956 );
    or g11017 ( n1963 , n4373 , n5628 );
    not g11018 ( n9653 , n12198 );
    not g11019 ( n897 , n6612 );
    and g11020 ( n7410 , n12234 , n7292 );
    not g11021 ( n8853 , n2055 );
    not g11022 ( n10520 , n816 );
    xor g11023 ( n4779 , n1453 , n1000 );
    or g11024 ( n8181 , n8026 , n11896 );
    xnor g11025 ( n5051 , n4914 , n10227 );
    or g11026 ( n9677 , n12853 , n12735 );
    not g11027 ( n7180 , n10642 );
    xnor g11028 ( n30 , n12089 , n5879 );
    and g11029 ( n3258 , n273 , n9126 );
    and g11030 ( n7171 , n6677 , n12175 );
    or g11031 ( n10738 , n12361 , n7952 );
    or g11032 ( n4726 , n2872 , n12816 );
    xnor g11033 ( n4609 , n2699 , n10941 );
    or g11034 ( n108 , n12062 , n73 );
    and g11035 ( n12394 , n3780 , n6329 );
    or g11036 ( n2207 , n2740 , n2844 );
    xnor g11037 ( n2555 , n12866 , n194 );
    not g11038 ( n22 , n5947 );
    xnor g11039 ( n10111 , n3448 , n12744 );
    and g11040 ( n10147 , n9108 , n3983 );
    or g11041 ( n7783 , n10196 , n4654 );
    xnor g11042 ( n4806 , n7289 , n12141 );
    not g11043 ( n7639 , n8359 );
    or g11044 ( n10242 , n128 , n5460 );
    or g11045 ( n10212 , n2332 , n6034 );
    xnor g11046 ( n7976 , n5867 , n11522 );
    not g11047 ( n3668 , n4432 );
    not g11048 ( n2676 , n6980 );
    xnor g11049 ( n6626 , n1147 , n729 );
    xnor g11050 ( n7375 , n11309 , n7738 );
    xnor g11051 ( n3973 , n2578 , n5842 );
    or g11052 ( n7885 , n5879 , n2940 );
    nor g11053 ( n12293 , n3946 , n7724 );
    xnor g11054 ( n3099 , n11117 , n7628 );
    or g11055 ( n4338 , n12853 , n10854 );
    xnor g11056 ( n5827 , n814 , n2847 );
    xnor g11057 ( n10505 , n5524 , n7877 );
    or g11058 ( n7802 , n9905 , n10792 );
    xnor g11059 ( n10276 , n5539 , n7430 );
    xnor g11060 ( n10488 , n1061 , n2685 );
    xnor g11061 ( n10413 , n7783 , n3710 );
    or g11062 ( n8835 , n10835 , n9078 );
    and g11063 ( n2463 , n1044 , n6668 );
    or g11064 ( n346 , n11958 , n8414 );
    xnor g11065 ( n5243 , n12109 , n3355 );
    or g11066 ( n948 , n4900 , n2219 );
    nor g11067 ( n3299 , n12584 , n5733 );
    nor g11068 ( n2442 , n8085 , n5180 );
    xnor g11069 ( n5461 , n4490 , n7459 );
    not g11070 ( n8364 , n11024 );
    or g11071 ( n10826 , n6977 , n11775 );
    or g11072 ( n2097 , n2099 , n7928 );
    xnor g11073 ( n5065 , n7651 , n10119 );
    xnor g11074 ( n2431 , n7618 , n12836 );
    not g11075 ( n1291 , n11094 );
    xnor g11076 ( n1306 , n7327 , n2971 );
    and g11077 ( n10683 , n11415 , n12606 );
    xnor g11078 ( n2102 , n6462 , n2094 );
    xnor g11079 ( n1060 , n4633 , n2255 );
    or g11080 ( n10604 , n9878 , n8109 );
    xnor g11081 ( n10107 , n1652 , n5498 );
    nor g11082 ( n6248 , n1524 , n8540 );
    and g11083 ( n4990 , n5964 , n7265 );
    xnor g11084 ( n2920 , n2116 , n12452 );
    or g11085 ( n3210 , n3820 , n9144 );
    or g11086 ( n9915 , n6373 , n1476 );
    xnor g11087 ( n9088 , n12208 , n10017 );
    not g11088 ( n10326 , n9060 );
    or g11089 ( n12313 , n7591 , n1787 );
    xnor g11090 ( n5080 , n10630 , n12861 );
    or g11091 ( n7097 , n11884 , n5992 );
    or g11092 ( n233 , n6977 , n10903 );
    xnor g11093 ( n11357 , n8598 , n5581 );
    or g11094 ( n3316 , n6283 , n3543 );
    or g11095 ( n9190 , n5355 , n10419 );
    nor g11096 ( n2641 , n6734 , n9049 );
    or g11097 ( n3933 , n6534 , n10826 );
    or g11098 ( n1709 , n7552 , n12553 );
    xnor g11099 ( n8480 , n1790 , n2016 );
    or g11100 ( n8891 , n6162 , n12432 );
    or g11101 ( n3298 , n8552 , n3224 );
    xnor g11102 ( n5066 , n6015 , n8673 );
    or g11103 ( n8386 , n1183 , n3924 );
    and g11104 ( n6621 , n6877 , n7946 );
    xnor g11105 ( n10616 , n8990 , n11496 );
    and g11106 ( n7172 , n7804 , n10341 );
    not g11107 ( n10799 , n1672 );
    or g11108 ( n2587 , n3324 , n28 );
    xnor g11109 ( n3350 , n8585 , n12187 );
    and g11110 ( n9980 , n1459 , n10330 );
    xnor g11111 ( n256 , n10245 , n8760 );
    and g11112 ( n4792 , n1011 , n864 );
    not g11113 ( n7678 , n1395 );
    not g11114 ( n2528 , n7865 );
    or g11115 ( n5664 , n10750 , n8109 );
    and g11116 ( n4528 , n2332 , n6034 );
    or g11117 ( n1207 , n989 , n7389 );
    or g11118 ( n9178 , n7509 , n3117 );
    or g11119 ( n5182 , n6504 , n3863 );
    and g11120 ( n7489 , n9076 , n4032 );
    xnor g11121 ( n3467 , n6824 , n6614 );
    and g11122 ( n3326 , n5331 , n1067 );
    or g11123 ( n10880 , n1699 , n9188 );
    xnor g11124 ( n377 , n4440 , n6083 );
    or g11125 ( n6818 , n11337 , n11092 );
    not g11126 ( n9280 , n6359 );
    or g11127 ( n870 , n5638 , n10767 );
    and g11128 ( n5962 , n343 , n7278 );
    and g11129 ( n6102 , n2330 , n6450 );
    not g11130 ( n1183 , n2515 );
    or g11131 ( n11587 , n6626 , n6106 );
    xnor g11132 ( n3027 , n7883 , n4341 );
    xnor g11133 ( n7216 , n5850 , n3218 );
    xnor g11134 ( n11435 , n3491 , n2954 );
    xnor g11135 ( n4188 , n5341 , n11947 );
    not g11136 ( n6171 , n6865 );
    and g11137 ( n2728 , n289 , n11772 );
    and g11138 ( n4909 , n3282 , n2907 );
    xnor g11139 ( n5247 , n7463 , n5146 );
    or g11140 ( n7715 , n2689 , n10649 );
    or g11141 ( n11526 , n12392 , n2231 );
    or g11142 ( n1676 , n10450 , n117 );
    or g11143 ( n8095 , n5329 , n9898 );
    not g11144 ( n6376 , n3574 );
    and g11145 ( n11085 , n11225 , n12559 );
    nor g11146 ( n1378 , n3949 , n5935 );
    or g11147 ( n1465 , n9373 , n9568 );
    or g11148 ( n3325 , n10350 , n7081 );
    xnor g11149 ( n2031 , n12437 , n11238 );
    and g11150 ( n6586 , n3386 , n129 );
    xnor g11151 ( n8636 , n3159 , n3459 );
    not g11152 ( n7506 , n12947 );
    or g11153 ( n1599 , n11923 , n9568 );
    or g11154 ( n11961 , n7495 , n5497 );
    and g11155 ( n766 , n3944 , n334 );
    and g11156 ( n4797 , n2496 , n10452 );
    or g11157 ( n9888 , n5337 , n3492 );
    or g11158 ( n8339 , n11552 , n4474 );
    not g11159 ( n3606 , n1478 );
    or g11160 ( n4759 , n4498 , n7341 );
    xnor g11161 ( n11715 , n7008 , n155 );
    and g11162 ( n12625 , n3909 , n6105 );
    not g11163 ( n11175 , n12895 );
    xnor g11164 ( n12277 , n3217 , n5669 );
    and g11165 ( n2402 , n2403 , n6763 );
    not g11166 ( n3477 , n8975 );
    xnor g11167 ( n4715 , n9113 , n12032 );
    or g11168 ( n3261 , n6426 , n11009 );
    xnor g11169 ( n6045 , n12016 , n6082 );
    or g11170 ( n4234 , n994 , n5497 );
    nor g11171 ( n2881 , n11451 , n6466 );
    or g11172 ( n901 , n3746 , n8414 );
    not g11173 ( n7413 , n9651 );
    xnor g11174 ( n1644 , n7374 , n7805 );
    not g11175 ( n12835 , n5032 );
    not g11176 ( n8832 , n3691 );
    or g11177 ( n910 , n7283 , n4242 );
    xnor g11178 ( n2434 , n1507 , n12153 );
    nor g11179 ( n1651 , n4972 , n2542 );
    xnor g11180 ( n329 , n12949 , n8289 );
    and g11181 ( n10113 , n9648 , n5802 );
    xnor g11182 ( n9181 , n9094 , n5113 );
    xnor g11183 ( n667 , n11608 , n3839 );
    not g11184 ( n4698 , n1445 );
    xnor g11185 ( n6724 , n12106 , n8284 );
    and g11186 ( n2665 , n7436 , n11023 );
    or g11187 ( n10670 , n8969 , n10961 );
    and g11188 ( n12916 , n9413 , n9022 );
    nor g11189 ( n11509 , n3059 , n10126 );
    or g11190 ( n5003 , n994 , n510 );
    not g11191 ( n7571 , n186 );
    not g11192 ( n684 , n12306 );
    xnor g11193 ( n7774 , n5003 , n892 );
    xnor g11194 ( n4915 , n8486 , n2411 );
    or g11195 ( n8469 , n807 , n12816 );
    and g11196 ( n8875 , n9383 , n8195 );
    and g11197 ( n9731 , n1072 , n2975 );
    and g11198 ( n501 , n6218 , n2156 );
    nor g11199 ( n12331 , n5350 , n3540 );
    not g11200 ( n1791 , n7527 );
    or g11201 ( n5181 , n12119 , n12686 );
    or g11202 ( n3828 , n10387 , n3019 );
    and g11203 ( n4989 , n718 , n1643 );
    or g11204 ( n12629 , n7951 , n7215 );
    xnor g11205 ( n1369 , n4166 , n4261 );
    or g11206 ( n3764 , n10108 , n6389 );
    or g11207 ( n3396 , n3096 , n11775 );
    not g11208 ( n11701 , n7321 );
    and g11209 ( n12411 , n2187 , n9061 );
    nor g11210 ( n2940 , n83 , n9710 );
    xnor g11211 ( n12894 , n3109 , n1103 );
    not g11212 ( n8254 , n11796 );
    or g11213 ( n1675 , n3743 , n7506 );
    not g11214 ( n9291 , n719 );
    or g11215 ( n1042 , n9411 , n12408 );
    xnor g11216 ( n8831 , n10154 , n5955 );
    or g11217 ( n6507 , n4778 , n826 );
    nor g11218 ( n132 , n4026 , n12410 );
    and g11219 ( n5649 , n2175 , n1709 );
    xnor g11220 ( n451 , n1126 , n6970 );
    xnor g11221 ( n1541 , n10222 , n6842 );
    nor g11222 ( n7237 , n9055 , n8077 );
    nor g11223 ( n9697 , n3906 , n11203 );
    or g11224 ( n1240 , n3746 , n2815 );
    xnor g11225 ( n11461 , n4131 , n3973 );
    not g11226 ( n10916 , n806 );
    or g11227 ( n7640 , n6373 , n795 );
    or g11228 ( n1075 , n3013 , n10567 );
    nor g11229 ( n8234 , n4692 , n4977 );
    xnor g11230 ( n7609 , n12604 , n11118 );
    and g11231 ( n564 , n6986 , n8595 );
    or g11232 ( n12175 , n5399 , n5400 );
    xnor g11233 ( n2451 , n4635 , n12369 );
    not g11234 ( n3240 , n6558 );
    or g11235 ( n11272 , n12530 , n12779 );
    xnor g11236 ( n4340 , n6859 , n10268 );
    and g11237 ( n11955 , n3504 , n524 );
    not g11238 ( n9214 , n1580 );
    xnor g11239 ( n8128 , n2124 , n3553 );
    and g11240 ( n11063 , n4207 , n3371 );
    not g11241 ( n9071 , n5684 );
    xnor g11242 ( n11875 , n3297 , n10757 );
    not g11243 ( n9313 , n8304 );
    not g11244 ( n4933 , n11677 );
    or g11245 ( n556 , n5200 , n1010 );
    not g11246 ( n7541 , n3724 );
    nor g11247 ( n5275 , n10730 , n11104 );
    or g11248 ( n3381 , n191 , n1079 );
    xnor g11249 ( n520 , n905 , n3168 );
    and g11250 ( n4252 , n12041 , n10416 );
    or g11251 ( n5423 , n9373 , n9144 );
    nor g11252 ( n7986 , n3347 , n8179 );
    xnor g11253 ( n4082 , n1820 , n3206 );
    nor g11254 ( n4125 , n2202 , n8402 );
    nor g11255 ( n1258 , n11503 , n10388 );
    xnor g11256 ( n11956 , n11479 , n4083 );
    or g11257 ( n3493 , n5519 , n1441 );
    or g11258 ( n1914 , n5945 , n995 );
    or g11259 ( n5667 , n11455 , n7614 );
    xnor g11260 ( n3125 , n12959 , n6355 );
    nor g11261 ( n12269 , n3570 , n9972 );
    or g11262 ( n12127 , n9079 , n6414 );
    not g11263 ( n10903 , n11023 );
    xnor g11264 ( n9608 , n5929 , n8196 );
    or g11265 ( n829 , n8552 , n5468 );
    nor g11266 ( n11116 , n12056 , n12678 );
    or g11267 ( n1998 , n7534 , n2079 );
    not g11268 ( n2366 , n7957 );
    not g11269 ( n11963 , n7463 );
    or g11270 ( n12507 , n5915 , n8259 );
    xnor g11271 ( n6478 , n1220 , n1410 );
    xnor g11272 ( n10228 , n3873 , n9320 );
    or g11273 ( n8074 , n8836 , n3941 );
    not g11274 ( n4830 , n7364 );
    xnor g11275 ( n12305 , n1468 , n9097 );
    and g11276 ( n2013 , n4151 , n3840 );
    xnor g11277 ( n6689 , n7720 , n1732 );
    and g11278 ( n6629 , n2824 , n10042 );
    xnor g11279 ( n5643 , n6983 , n10037 );
    not g11280 ( n12574 , n4989 );
    and g11281 ( n9124 , n5684 , n563 );
    xnor g11282 ( n2799 , n98 , n5768 );
    xnor g11283 ( n1152 , n5393 , n6733 );
    xnor g11284 ( n8553 , n12932 , n2320 );
    and g11285 ( n5503 , n12776 , n12587 );
    xnor g11286 ( n2240 , n2965 , n5968 );
    or g11287 ( n12694 , n3025 , n6054 );
    not g11288 ( n8648 , n6806 );
    and g11289 ( n10762 , n7388 , n12704 );
    xnor g11290 ( n4102 , n12003 , n10876 );
    or g11291 ( n10595 , n7959 , n2725 );
    not g11292 ( n12467 , n6356 );
    and g11293 ( n10596 , n7539 , n1328 );
    and g11294 ( n3929 , n6137 , n9404 );
    xnor g11295 ( n9756 , n3479 , n4505 );
    or g11296 ( n8413 , n3560 , n3505 );
    nor g11297 ( n3453 , n7739 , n9057 );
    xnor g11298 ( n6958 , n4316 , n943 );
    xnor g11299 ( n10841 , n11147 , n12850 );
    or g11300 ( n6769 , n1156 , n871 );
    or g11301 ( n7999 , n1362 , n8878 );
    not g11302 ( n6454 , n1236 );
    xnor g11303 ( n6366 , n11172 , n4832 );
    xnor g11304 ( n9850 , n4250 , n7101 );
    not g11305 ( n11097 , n10522 );
    xnor g11306 ( n8867 , n12785 , n3806 );
    xnor g11307 ( n1930 , n7366 , n10062 );
    xnor g11308 ( n549 , n337 , n12329 );
    not g11309 ( n896 , n4119 );
    or g11310 ( n5337 , n8373 , n1940 );
    not g11311 ( n11745 , n1419 );
    or g11312 ( n10823 , n4628 , n5468 );
    xnor g11313 ( n5079 , n1528 , n2273 );
    and g11314 ( n8046 , n9308 , n9562 );
    xnor g11315 ( n2290 , n3132 , n435 );
    xnor g11316 ( n8850 , n7632 , n4518 );
    xnor g11317 ( n7254 , n7697 , n8566 );
    nor g11318 ( n1604 , n11 , n10159 );
    not g11319 ( n10190 , n3973 );
    nor g11320 ( n6348 , n8235 , n4597 );
    xnor g11321 ( n571 , n6654 , n3765 );
    xnor g11322 ( n10023 , n5251 , n7695 );
    xnor g11323 ( n2645 , n11425 , n6025 );
    not g11324 ( n3435 , n6195 );
    nor g11325 ( n5492 , n2944 , n4398 );
    or g11326 ( n713 , n2272 , n10258 );
    xnor g11327 ( n2518 , n6180 , n3678 );
    or g11328 ( n8216 , n752 , n7952 );
    xnor g11329 ( n12334 , n6347 , n9890 );
    and g11330 ( n8656 , n12069 , n5645 );
    or g11331 ( n971 , n4671 , n8300 );
    nor g11332 ( n3542 , n8831 , n3918 );
    not g11333 ( n11941 , n11836 );
    and g11334 ( n67 , n4856 , n10610 );
    and g11335 ( n1065 , n10517 , n8799 );
    xnor g11336 ( n9973 , n3802 , n8151 );
    and g11337 ( n10100 , n1923 , n6640 );
    xnor g11338 ( n9544 , n456 , n779 );
    xnor g11339 ( n3881 , n3121 , n2436 );
    and g11340 ( n2875 , n10745 , n12072 );
    xnor g11341 ( n954 , n7914 , n4351 );
    or g11342 ( n5450 , n11716 , n9460 );
    or g11343 ( n1452 , n848 , n2910 );
    xnor g11344 ( n3824 , n6553 , n11062 );
    and g11345 ( n11586 , n12327 , n1660 );
    not g11346 ( n7613 , n2890 );
    xnor g11347 ( n1631 , n5407 , n5390 );
    nor g11348 ( n6019 , n1515 , n4832 );
    and g11349 ( n6750 , n3084 , n2801 );
    and g11350 ( n3609 , n11851 , n9255 );
    not g11351 ( n3965 , n6413 );
    and g11352 ( n3647 , n3959 , n2008 );
    xnor g11353 ( n2818 , n6745 , n2888 );
    xnor g11354 ( n7148 , n4098 , n11217 );
    xnor g11355 ( n5714 , n1140 , n10543 );
    not g11356 ( n4832 , n2218 );
    xnor g11357 ( n1135 , n334 , n9156 );
    nor g11358 ( n12717 , n8688 , n7086 );
    xnor g11359 ( n1318 , n1814 , n5708 );
    not g11360 ( n1084 , n1217 );
    xnor g11361 ( n10901 , n1072 , n11051 );
    xnor g11362 ( n6215 , n2532 , n1880 );
    xnor g11363 ( n5717 , n9546 , n5184 );
    xnor g11364 ( n10314 , n5456 , n87 );
    xnor g11365 ( n12684 , n6296 , n10197 );
    xnor g11366 ( n7239 , n11136 , n8370 );
    or g11367 ( n10482 , n3682 , n8958 );
    xnor g11368 ( n7241 , n2593 , n8497 );
    or g11369 ( n7474 , n8959 , n9741 );
    and g11370 ( n332 , n5949 , n661 );
    not g11371 ( n11319 , n2411 );
    and g11372 ( n6394 , n11805 , n8047 );
    xnor g11373 ( n2857 , n6036 , n4348 );
    or g11374 ( n1558 , n12855 , n9717 );
    nor g11375 ( n6966 , n8736 , n12526 );
    or g11376 ( n12525 , n4628 , n1932 );
    xnor g11377 ( n12073 , n8225 , n9202 );
    nor g11378 ( n359 , n11656 , n1416 );
    xnor g11379 ( n10758 , n8245 , n8464 );
    xnor g11380 ( n4626 , n5596 , n9906 );
    not g11381 ( n1114 , n4897 );
    not g11382 ( n3120 , n7908 );
    or g11383 ( n2735 , n8339 , n4450 );
    or g11384 ( n5230 , n9151 , n951 );
    xnor g11385 ( n2096 , n9038 , n7623 );
    nor g11386 ( n6845 , n1585 , n11269 );
    or g11387 ( n9869 , n5355 , n6389 );
    nor g11388 ( n8105 , n8320 , n232 );
    or g11389 ( n1415 , n3096 , n11820 );
    xnor g11390 ( n2527 , n4290 , n12634 );
    or g11391 ( n3291 , n12935 , n9808 );
    xnor g11392 ( n4286 , n197 , n10689 );
    xnor g11393 ( n553 , n8077 , n3575 );
    xnor g11394 ( n11612 , n4960 , n4851 );
    xnor g11395 ( n4088 , n2485 , n9542 );
    or g11396 ( n11712 , n2099 , n2964 );
    nor g11397 ( n4011 , n2790 , n666 );
    or g11398 ( n12355 , n8642 , n259 );
    not g11399 ( n8599 , n7286 );
    or g11400 ( n10222 , n11635 , n3037 );
    not g11401 ( n12446 , n4094 );
    and g11402 ( n8003 , n6542 , n8891 );
    xnor g11403 ( n1307 , n4087 , n5451 );
    and g11404 ( n4371 , n6458 , n9204 );
    and g11405 ( n6158 , n7157 , n6746 );
    nor g11406 ( n11981 , n6643 , n9092 );
    and g11407 ( n3478 , n5240 , n4921 );
    xnor g11408 ( n2301 , n1663 , n7833 );
    nor g11409 ( n1176 , n12246 , n287 );
    xnor g11410 ( n2035 , n11060 , n11247 );
    or g11411 ( n1985 , n3236 , n3067 );
    and g11412 ( n9092 , n8736 , n12526 );
    and g11413 ( n10628 , n35 , n887 );
    and g11414 ( n12086 , n4728 , n10505 );
    not g11415 ( n151 , n10790 );
    not g11416 ( n8067 , n11002 );
    and g11417 ( n5820 , n11153 , n8433 );
    not g11418 ( n8735 , n615 );
    xnor g11419 ( n6346 , n6078 , n2672 );
    nor g11420 ( n2698 , n9186 , n7172 );
    or g11421 ( n11741 , n7495 , n6389 );
    xnor g11422 ( n2129 , n1191 , n9630 );
    xnor g11423 ( n12339 , n8945 , n11068 );
    xnor g11424 ( n6194 , n4619 , n9932 );
    not g11425 ( n9397 , n753 );
    xnor g11426 ( n3849 , n1265 , n4293 );
    not g11427 ( n12669 , n7693 );
    or g11428 ( n12112 , n9370 , n10066 );
    or g11429 ( n4899 , n5915 , n9586 );
    or g11430 ( n11727 , n752 , n5311 );
    not g11431 ( n957 , n10770 );
    or g11432 ( n12960 , n12119 , n5781 );
    or g11433 ( n6271 , n6718 , n4654 );
    nor g11434 ( n9559 , n2972 , n10888 );
    nor g11435 ( n12782 , n12131 , n11647 );
    and g11436 ( n12811 , n1731 , n2068 );
    and g11437 ( n5442 , n8778 , n12718 );
    not g11438 ( n8026 , n10928 );
    and g11439 ( n1090 , n158 , n9260 );
    xnor g11440 ( n5103 , n5963 , n4102 );
    nor g11441 ( n3177 , n9355 , n2065 );
    not g11442 ( n6530 , n9345 );
    and g11443 ( n9528 , n2739 , n1033 );
    xnor g11444 ( n4703 , n4232 , n12549 );
    or g11445 ( n9700 , n4540 , n4448 );
    xnor g11446 ( n3068 , n11318 , n8924 );
    xnor g11447 ( n1902 , n10507 , n1484 );
    or g11448 ( n2786 , n7713 , n4012 );
    xnor g11449 ( n6258 , n4612 , n2417 );
    or g11450 ( n11485 , n12586 , n1320 );
    or g11451 ( n8777 , n3630 , n6831 );
    nor g11452 ( n2783 , n2311 , n5206 );
    or g11453 ( n2224 , n1494 , n7198 );
    nor g11454 ( n11626 , n791 , n5226 );
    and g11455 ( n11361 , n11327 , n599 );
    xnor g11456 ( n5272 , n9122 , n430 );
    or g11457 ( n5593 , n2036 , n2853 );
    xnor g11458 ( n4745 , n5014 , n11938 );
    and g11459 ( n9527 , n8515 , n10629 );
    xnor g11460 ( n12922 , n3519 , n6751 );
    nor g11461 ( n8642 , n12582 , n10891 );
    or g11462 ( n1470 , n10364 , n5156 );
    and g11463 ( n986 , n12845 , n260 );
    xor g11464 ( n7510 , n10566 , n2183 );
    or g11465 ( n2642 , n989 , n11430 );
    or g11466 ( n1664 , n6131 , n2060 );
    not g11467 ( n7495 , n12025 );
    xnor g11468 ( n5263 , n11388 , n11314 );
    or g11469 ( n9931 , n636 , n530 );
    not g11470 ( n28 , n5760 );
    or g11471 ( n3282 , n12142 , n4458 );
    and g11472 ( n9723 , n11538 , n8798 );
    or g11473 ( n5543 , n6654 , n8578 );
    and g11474 ( n4646 , n2207 , n5795 );
    xnor g11475 ( n391 , n6472 , n8457 );
    xnor g11476 ( n6916 , n6310 , n1606 );
    xnor g11477 ( n9715 , n12855 , n11989 );
    and g11478 ( n10302 , n3007 , n8561 );
    nor g11479 ( n1974 , n8986 , n10680 );
    xnor g11480 ( n4368 , n11986 , n11644 );
    nor g11481 ( n3051 , n4756 , n6010 );
    xnor g11482 ( n1775 , n4202 , n9497 );
    nor g11483 ( n7313 , n10098 , n4004 );
    not g11484 ( n11457 , n9778 );
    not g11485 ( n10196 , n5860 );
    xnor g11486 ( n4932 , n10475 , n748 );
    or g11487 ( n5361 , n12853 , n7382 );
    xnor g11488 ( n847 , n9150 , n5308 );
    or g11489 ( n3959 , n3746 , n9741 );
    xnor g11490 ( n7987 , n4457 , n11041 );
    not g11491 ( n5878 , n6269 );
    xnor g11492 ( n4361 , n4601 , n7093 );
    xnor g11493 ( n7106 , n10531 , n670 );
    not g11494 ( n2472 , n952 );
    or g11495 ( n8633 , n10835 , n5759 );
    not g11496 ( n2186 , n2992 );
    and g11497 ( n4844 , n6365 , n6285 );
    and g11498 ( n250 , n5353 , n1171 );
    or g11499 ( n1139 , n3820 , n9160 );
    and g11500 ( n7637 , n2523 , n5753 );
    nor g11501 ( n10168 , n1999 , n7171 );
    and g11502 ( n2269 , n3367 , n3056 );
    or g11503 ( n3715 , n8564 , n12226 );
    xnor g11504 ( n4181 , n6148 , n2748 );
    xnor g11505 ( n9906 , n9508 , n146 );
    or g11506 ( n4972 , n5355 , n5851 );
    nor g11507 ( n902 , n3596 , n7345 );
    and g11508 ( n7760 , n7271 , n11263 );
    xnor g11509 ( n7155 , n4286 , n8472 );
    and g11510 ( n8057 , n12227 , n11940 );
    xnor g11511 ( n10631 , n4513 , n2331 );
    xnor g11512 ( n7746 , n2057 , n1431 );
    or g11513 ( n9729 , n9373 , n9521 );
    not g11514 ( n3666 , n9440 );
    not g11515 ( n1657 , n8671 );
    and g11516 ( n2174 , n161 , n550 );
    xnor g11517 ( n5001 , n2892 , n2299 );
    not g11518 ( n8177 , n4949 );
    and g11519 ( n8601 , n5593 , n2800 );
    and g11520 ( n1008 , n6857 , n4544 );
    or g11521 ( n9614 , n807 , n5012 );
    and g11522 ( n12872 , n8556 , n12794 );
    xnor g11523 ( n5726 , n6374 , n2230 );
    and g11524 ( n6508 , n2763 , n789 );
    xnor g11525 ( n6532 , n5420 , n7855 );
    nor g11526 ( n9599 , n25 , n3952 );
    xnor g11527 ( n1894 , n7085 , n1725 );
    xnor g11528 ( n6139 , n9383 , n8195 );
    or g11529 ( n4892 , n2217 , n5914 );
    not g11530 ( n6849 , n2878 );
    or g11531 ( n5347 , n12907 , n12636 );
    xnor g11532 ( n5806 , n1686 , n860 );
    xnor g11533 ( n5063 , n4255 , n9501 );
    xnor g11534 ( n6603 , n3133 , n6541 );
    and g11535 ( n12536 , n7932 , n6065 );
    nor g11536 ( n12408 , n440 , n5986 );
    and g11537 ( n4377 , n4047 , n7770 );
    not g11538 ( n27 , n6896 );
    xnor g11539 ( n12254 , n11801 , n4071 );
    or g11540 ( n8834 , n7611 , n1296 );
    not g11541 ( n1929 , n12309 );
    not g11542 ( n4572 , n2177 );
    not g11543 ( n12535 , n12925 );
    and g11544 ( n3795 , n10394 , n9265 );
    and g11545 ( n6238 , n11011 , n3869 );
    not g11546 ( n6418 , n1147 );
    or g11547 ( n11048 , n796 , n6116 );
    xnor g11548 ( n20 , n8474 , n12570 );
    xnor g11549 ( n229 , n10627 , n3656 );
    or g11550 ( n1409 , n12119 , n10422 );
    or g11551 ( n11514 , n2832 , n10066 );
    not g11552 ( n10145 , n7052 );
    not g11553 ( n9642 , n8892 );
    xnor g11554 ( n6087 , n3047 , n11403 );
    xnor g11555 ( n5794 , n1550 , n7129 );
    or g11556 ( n4961 , n8026 , n7425 );
    and g11557 ( n5019 , n4904 , n701 );
    xnor g11558 ( n6645 , n10525 , n1245 );
    not g11559 ( n10339 , n3146 );
    or g11560 ( n11925 , n8428 , n184 );
    or g11561 ( n8704 , n994 , n7881 );
    or g11562 ( n4710 , n10750 , n12754 );
    nor g11563 ( n5636 , n4868 , n11379 );
    xor g11564 ( n5191 , n2342 , n6926 );
    nor g11565 ( n8248 , n10529 , n12337 );
    or g11566 ( n1392 , n11958 , n12899 );
    and g11567 ( n10229 , n9043 , n10840 );
    and g11568 ( n3632 , n12208 , n10017 );
    xnor g11569 ( n11440 , n3150 , n9127 );
    xnor g11570 ( n11178 , n872 , n230 );
    and g11571 ( n11942 , n7705 , n11863 );
    xnor g11572 ( n2892 , n6668 , n3637 );
    or g11573 ( n10792 , n7449 , n12771 );
    and g11574 ( n6462 , n10987 , n5526 );
    xnor g11575 ( n1924 , n9530 , n193 );
    xnor g11576 ( n6350 , n7105 , n6716 );
    or g11577 ( n12630 , n4059 , n10419 );
    xnor g11578 ( n10918 , n6342 , n3655 );
    xnor g11579 ( n7666 , n9041 , n6276 );
    or g11580 ( n6442 , n4911 , n7424 );
    xor g11581 ( n8809 , n5563 , n4367 );
    xnor g11582 ( n8846 , n8555 , n6064 );
    xnor g11583 ( n2744 , n1958 , n5232 );
    xnor g11584 ( n551 , n3982 , n6005 );
    xnor g11585 ( n6012 , n10368 , n7269 );
    nor g11586 ( n172 , n8442 , n12252 );
    or g11587 ( n10698 , n12098 , n5499 );
    and g11588 ( n8396 , n8458 , n3761 );
    xnor g11589 ( n5618 , n2153 , n704 );
    not g11590 ( n5977 , n804 );
    not g11591 ( n4946 , n12315 );
    not g11592 ( n3127 , n11757 );
    not g11593 ( n3073 , n3814 );
    nor g11594 ( n3528 , n10235 , n3427 );
    or g11595 ( n308 , n12119 , n6513 );
    xnor g11596 ( n7580 , n4374 , n3595 );
    xnor g11597 ( n951 , n695 , n2389 );
    or g11598 ( n5386 , n3096 , n6169 );
    nor g11599 ( n12382 , n2999 , n7484 );
    xnor g11600 ( n3069 , n8102 , n3854 );
    or g11601 ( n2208 , n8428 , n11775 );
    xnor g11602 ( n11173 , n9275 , n8402 );
    nor g11603 ( n12322 , n12211 , n3394 );
    or g11604 ( n1303 , n12327 , n1660 );
    and g11605 ( n12399 , n9701 , n2799 );
    not g11606 ( n12868 , n9728 );
    xnor g11607 ( n2314 , n6305 , n4761 );
    or g11608 ( n11571 , n1031 , n8378 );
    not g11609 ( n11907 , n4583 );
    not g11610 ( n7125 , n8091 );
    or g11611 ( n778 , n1937 , n3421 );
    xnor g11612 ( n594 , n3881 , n10612 );
    xnor g11613 ( n10153 , n6911 , n52 );
    xnor g11614 ( n8849 , n9082 , n7944 );
    or g11615 ( n982 , n12053 , n4464 );
    or g11616 ( n7061 , n2268 , n3351 );
    xnor g11617 ( n11814 , n7694 , n12015 );
    xnor g11618 ( n3753 , n4849 , n963 );
    or g11619 ( n6404 , n11681 , n2728 );
    xnor g11620 ( n3390 , n7737 , n2000 );
    and g11621 ( n10425 , n7461 , n7892 );
    and g11622 ( n4955 , n3221 , n3314 );
    or g11623 ( n2394 , n1833 , n9684 );
    or g11624 ( n7706 , n10585 , n11862 );
    xnor g11625 ( n6762 , n6058 , n10182 );
    xnor g11626 ( n3526 , n3036 , n6549 );
    xnor g11627 ( n12948 , n4380 , n5245 );
    xnor g11628 ( n3499 , n9072 , n12574 );
    not g11629 ( n3198 , n868 );
    xnor g11630 ( n2648 , n11245 , n4725 );
    xnor g11631 ( n4860 , n2846 , n7904 );
    or g11632 ( n1827 , n10478 , n4055 );
    xnor g11633 ( n12257 , n3003 , n2843 );
    xnor g11634 ( n5634 , n11156 , n11906 );
    or g11635 ( n4537 , n8618 , n2247 );
    nor g11636 ( n4935 , n7655 , n9410 );
    not g11637 ( n1567 , n3753 );
    xnor g11638 ( n5952 , n12525 , n6571 );
    nor g11639 ( n1054 , n5128 , n5018 );
    or g11640 ( n5812 , n10157 , n11698 );
    or g11641 ( n1934 , n10750 , n5468 );
    and g11642 ( n12818 , n6261 , n6732 );
    or g11643 ( n3582 , n8959 , n5538 );
    or g11644 ( n3561 , n11026 , n4654 );
    nor g11645 ( n2063 , n7087 , n611 );
    or g11646 ( n1449 , n12361 , n995 );
    xnor g11647 ( n4388 , n3399 , n4328 );
    xnor g11648 ( n1984 , n9594 , n2370 );
    or g11649 ( n2542 , n4059 , n12328 );
    xnor g11650 ( n6276 , n8674 , n5642 );
    not g11651 ( n7283 , n5964 );
    or g11652 ( n9354 , n6977 , n5540 );
    or g11653 ( n2124 , n3746 , n11896 );
    nor g11654 ( n2647 , n2661 , n9511 );
    not g11655 ( n4775 , n2253 );
    xnor g11656 ( n414 , n3078 , n6032 );
    not g11657 ( n10661 , n6096 );
    or g11658 ( n6616 , n9027 , n1588 );
    and g11659 ( n10256 , n7912 , n4136 );
    not g11660 ( n11029 , n8129 );
    and g11661 ( n1395 , n168 , n6761 );
    not g11662 ( n11484 , n10747 );
    xnor g11663 ( n5073 , n10932 , n8425 );
    and g11664 ( n8646 , n5977 , n1716 );
    and g11665 ( n7315 , n8813 , n9401 );
    xnor g11666 ( n3732 , n11777 , n470 );
    or g11667 ( n11139 , n9713 , n9873 );
    xnor g11668 ( n7915 , n9260 , n3981 );
    xnor g11669 ( n9540 , n1599 , n11816 );
    and g11670 ( n11503 , n6547 , n670 );
    and g11671 ( n187 , n12299 , n8595 );
    and g11672 ( n5966 , n2790 , n666 );
    xnor g11673 ( n5034 , n6390 , n322 );
    or g11674 ( n1744 , n29 , n4027 );
    or g11675 ( n3650 , n5530 , n3924 );
    xnor g11676 ( n2198 , n4279 , n3446 );
    and g11677 ( n8632 , n8132 , n7867 );
    nor g11678 ( n7011 , n5482 , n6960 );
    and g11679 ( n8544 , n201 , n8695 );
    and g11680 ( n2713 , n2843 , n3578 );
    not g11681 ( n5985 , n1355 );
    xnor g11682 ( n10757 , n3140 , n3447 );
    not g11683 ( n6417 , n2827 );
    and g11684 ( n95 , n8091 , n3759 );
    not g11685 ( n11889 , n3054 );
    or g11686 ( n6973 , n9921 , n10533 );
    xnor g11687 ( n6910 , n871 , n2769 );
    not g11688 ( n9563 , n3420 );
    xnor g11689 ( n6932 , n5259 , n828 );
    not g11690 ( n6327 , n8392 );
    not g11691 ( n12214 , n8844 );
    or g11692 ( n1944 , n6423 , n7786 );
    and g11693 ( n1100 , n6204 , n11735 );
    and g11694 ( n8019 , n5429 , n7702 );
    xnor g11695 ( n4794 , n1696 , n218 );
    or g11696 ( n2701 , n4062 , n5962 );
    xnor g11697 ( n5130 , n8956 , n12922 );
    nor g11698 ( n1613 , n9223 , n12179 );
    or g11699 ( n6305 , n8687 , n4527 );
    xnor g11700 ( n12345 , n2296 , n8206 );
    or g11701 ( n12792 , n11527 , n8072 );
    and g11702 ( n4304 , n8204 , n3064 );
    or g11703 ( n8383 , n4066 , n8800 );
    and g11704 ( n10759 , n1475 , n4986 );
    and g11705 ( n959 , n8070 , n473 );
    or g11706 ( n7480 , n10835 , n609 );
    or g11707 ( n4729 , n10709 , n4822 );
    nor g11708 ( n11630 , n335 , n6702 );
    and g11709 ( n4788 , n5088 , n3636 );
    or g11710 ( n2419 , n4343 , n12535 );
    or g11711 ( n5147 , n7495 , n1851 );
    xnor g11712 ( n1658 , n11966 , n9847 );
    and g11713 ( n11120 , n4519 , n7109 );
    not g11714 ( n10952 , n7064 );
    or g11715 ( n6543 , n3820 , n795 );
    not g11716 ( n7115 , n1016 );
    xnor g11717 ( n12473 , n5499 , n6638 );
    not g11718 ( n12170 , n11971 );
    xnor g11719 ( n6434 , n3371 , n11323 );
    xnor g11720 ( n11231 , n3639 , n6499 );
    or g11721 ( n10814 , n6373 , n12120 );
    xnor g11722 ( n2203 , n3875 , n657 );
    nor g11723 ( n5273 , n8770 , n8248 );
    not g11724 ( n4111 , n8475 );
    or g11725 ( n13 , n2832 , n1162 );
    and g11726 ( n666 , n4016 , n9314 );
    or g11727 ( n7533 , n6864 , n451 );
    nor g11728 ( n4093 , n4042 , n11666 );
    xnor g11729 ( n11895 , n8145 , n3449 );
    and g11730 ( n9110 , n5844 , n5938 );
    not g11731 ( n5002 , n4752 );
    xnor g11732 ( n8932 , n2319 , n1874 );
    or g11733 ( n2615 , n874 , n109 );
    nor g11734 ( n7086 , n1178 , n3563 );
    and g11735 ( n9211 , n8262 , n3085 );
    xnor g11736 ( n9533 , n10347 , n12182 );
    xnor g11737 ( n675 , n5556 , n642 );
    xnor g11738 ( n4007 , n8068 , n11566 );
    or g11739 ( n11390 , n11958 , n9741 );
    or g11740 ( n7238 , n3324 , n4654 );
    xnor g11741 ( n6272 , n5266 , n12868 );
    or g11742 ( n12426 , n6977 , n6169 );
    not g11743 ( n3160 , n4577 );
    nor g11744 ( n7219 , n3901 , n3929 );
    not g11745 ( n10026 , n9603 );
    or g11746 ( n5029 , n6600 , n2074 );
    and g11747 ( n6644 , n4127 , n5890 );
    or g11748 ( n7889 , n12203 , n10593 );
    and g11749 ( n4220 , n1812 , n10855 );
    not g11750 ( n9568 , n3342 );
    and g11751 ( n10987 , n12069 , n2498 );
    and g11752 ( n259 , n7352 , n3893 );
    and g11753 ( n5224 , n835 , n7979 );
    or g11754 ( n5689 , n5518 , n3990 );
    or g11755 ( n943 , n1165 , n1640 );
    nor g11756 ( n11607 , n4138 , n4587 );
    xnor g11757 ( n9396 , n2401 , n11973 );
    xnor g11758 ( n750 , n8936 , n10192 );
    and g11759 ( n1298 , n10735 , n4091 );
    not g11760 ( n6185 , n10929 );
    xnor g11761 ( n4551 , n895 , n6206 );
    or g11762 ( n3424 , n6718 , n5258 );
    xnor g11763 ( n12207 , n12920 , n2113 );
    not g11764 ( n1283 , n5895 );
    or g11765 ( n5886 , n3735 , n2325 );
    and g11766 ( n1587 , n3530 , n11583 );
    or g11767 ( n6252 , n10417 , n10146 );
    xnor g11768 ( n4378 , n12787 , n2960 );
    xnor g11769 ( n6682 , n1420 , n557 );
    and g11770 ( n1371 , n8477 , n8952 );
    and g11771 ( n8316 , n5064 , n8974 );
    nor g11772 ( n8219 , n181 , n5375 );
    xnor g11773 ( n8144 , n10107 , n6156 );
    or g11774 ( n573 , n10142 , n7341 );
    xnor g11775 ( n6121 , n1973 , n8779 );
    or g11776 ( n9380 , n3728 , n7740 );
    or g11777 ( n10198 , n699 , n7085 );
    and g11778 ( n5764 , n3757 , n10363 );
    and g11779 ( n1481 , n827 , n3264 );
    xnor g11780 ( n838 , n7998 , n4153 );
    and g11781 ( n1830 , n9158 , n2390 );
    and g11782 ( n8027 , n10635 , n8078 );
    not g11783 ( n8337 , n8585 );
    or g11784 ( n11960 , n8127 , n7424 );
    or g11785 ( n6311 , n12275 , n12086 );
    xnor g11786 ( n8341 , n6569 , n4031 );
    nor g11787 ( n6658 , n961 , n9553 );
    and g11788 ( n1592 , n2526 , n8491 );
    xnor g11789 ( n2000 , n11116 , n10050 );
    and g11790 ( n9199 , n3992 , n12704 );
    or g11791 ( n1396 , n6808 , n9124 );
    and g11792 ( n11280 , n11402 , n6953 );
    and g11793 ( n2643 , n4989 , n4764 );
    or g11794 ( n12799 , n1051 , n11896 );
    and g11795 ( n1669 , n3033 , n1049 );
    or g11796 ( n12882 , n10142 , n8970 );
    and g11797 ( n8409 , n97 , n2129 );
    or g11798 ( n10574 , n8428 , n12899 );
    or g11799 ( n12842 , n0 , n9322 );
    or g11800 ( n3215 , n7116 , n7876 );
    or g11801 ( n11401 , n12119 , n8644 );
    xnor g11802 ( n4162 , n2527 , n7257 );
    and g11803 ( n3833 , n1333 , n2585 );
    xnor g11804 ( n9998 , n6407 , n2208 );
    xnor g11805 ( n2263 , n1035 , n2836 );
    nor g11806 ( n5280 , n8758 , n12630 );
    or g11807 ( n7285 , n11552 , n9160 );
    and g11808 ( n8344 , n7181 , n11962 );
    or g11809 ( n2069 , n191 , n1851 );
    xnor g11810 ( n5140 , n4656 , n1781 );
    nor g11811 ( n10682 , n12923 , n5966 );
    not g11812 ( n9692 , n7758 );
    xnor g11813 ( n12125 , n6448 , n7570 );
    nor g11814 ( n5448 , n2365 , n9612 );
    not g11815 ( n7341 , n11917 );
    and g11816 ( n854 , n5449 , n427 );
    or g11817 ( n1607 , n8583 , n9160 );
    and g11818 ( n5609 , n4154 , n5746 );
    or g11819 ( n1826 , n12119 , n4913 );
    xnor g11820 ( n1351 , n12316 , n8576 );
    and g11821 ( n5713 , n6993 , n9915 );
    xnor g11822 ( n1173 , n8216 , n4183 );
    xnor g11823 ( n5440 , n9415 , n9968 );
    and g11824 ( n87 , n12477 , n9178 );
    xnor g11825 ( n12959 , n5790 , n12174 );
    and g11826 ( n4874 , n3706 , n10461 );
    xnor g11827 ( n10215 , n2240 , n6127 );
    xnor g11828 ( n4800 , n6151 , n694 );
    or g11829 ( n6316 , n6977 , n11410 );
    nor g11830 ( n4694 , n3965 , n12778 );
    and g11831 ( n9890 , n7282 , n11604 );
    xnor g11832 ( n10246 , n1003 , n6265 );
    xnor g11833 ( n10608 , n2917 , n2426 );
    not g11834 ( n3062 , n5783 );
    or g11835 ( n3368 , n8583 , n5502 );
    and g11836 ( n6613 , n2599 , n10681 );
    xnor g11837 ( n9673 , n4787 , n1889 );
    xnor g11838 ( n11570 , n132 , n5637 );
    and g11839 ( n7235 , n9048 , n5993 );
    or g11840 ( n8533 , n4059 , n7703 );
    xnor g11841 ( n3187 , n4339 , n5246 );
    or g11842 ( n11939 , n8870 , n8109 );
    not g11843 ( n3429 , n3805 );
    or g11844 ( n5832 , n752 , n11820 );
    and g11845 ( n6149 , n6182 , n11336 );
    nor g11846 ( n9704 , n10718 , n6585 );
    or g11847 ( n5779 , n6881 , n6489 );
    or g11848 ( n3314 , n4059 , n8524 );
    or g11849 ( n6632 , n5548 , n9768 );
    xnor g11850 ( n9143 , n6387 , n1487 );
    not g11851 ( n9782 , n5229 );
    xnor g11852 ( n4598 , n6072 , n5473 );
    xnor g11853 ( n8980 , n6881 , n6489 );
    xnor g11854 ( n9386 , n10002 , n2587 );
    not g11855 ( n7633 , n4260 );
    xnor g11856 ( n9176 , n10304 , n6928 );
    or g11857 ( n4533 , n4951 , n11496 );
    xnor g11858 ( n5412 , n10137 , n2179 );
    and g11859 ( n5227 , n4648 , n10473 );
    and g11860 ( n5590 , n10479 , n6884 );
    not g11861 ( n6301 , n10692 );
    and g11862 ( n10360 , n7212 , n8772 );
    or g11863 ( n4053 , n2456 , n8740 );
    xnor g11864 ( n7953 , n6562 , n8861 );
    or g11865 ( n4332 , n5691 , n6338 );
    or g11866 ( n11576 , n9335 , n11031 );
    or g11867 ( n4515 , n9172 , n11949 );
    or g11868 ( n7538 , n11864 , n8943 );
    xnor g11869 ( n5072 , n710 , n12851 );
    nor g11870 ( n922 , n3643 , n8741 );
    xnor g11871 ( n8497 , n5752 , n5930 );
    xnor g11872 ( n5626 , n7688 , n11465 );
    not g11873 ( n10032 , n3975 );
    nor g11874 ( n1735 , n5146 , n11963 );
    and g11875 ( n8460 , n3498 , n6048 );
    xnor g11876 ( n9018 , n7919 , n10756 );
    and g11877 ( n3012 , n392 , n9940 );
    and g11878 ( n11101 , n10842 , n5823 );
    and g11879 ( n8725 , n10485 , n2084 );
    or g11880 ( n739 , n5005 , n1968 );
    or g11881 ( n12164 , n305 , n3321 );
    xnor g11882 ( n10975 , n1373 , n1074 );
    xnor g11883 ( n10483 , n12072 , n6263 );
    or g11884 ( n12413 , n5981 , n5661 );
    and g11885 ( n10657 , n420 , n10308 );
    xnor g11886 ( n8231 , n7185 , n2895 );
    nor g11887 ( n2561 , n4124 , n11935 );
    xnor g11888 ( n1440 , n9161 , n11766 );
    or g11889 ( n8612 , n994 , n5851 );
    or g11890 ( n4681 , n8127 , n11746 );
    xor g11891 ( n852 , n12790 , n7255 );
    xnor g11892 ( n12418 , n2427 , n9801 );
    not g11893 ( n12699 , n1009 );
    nor g11894 ( n5920 , n10566 , n6730 );
    or g11895 ( n11288 , n5856 , n10890 );
    xnor g11896 ( n10407 , n3285 , n5513 );
    nor g11897 ( n12494 , n1575 , n6521 );
    xnor g11898 ( n8372 , n10820 , n10737 );
    or g11899 ( n467 , n1290 , n7002 );
    xnor g11900 ( n8918 , n183 , n10638 );
    and g11901 ( n11009 , n9588 , n3832 );
    xnor g11902 ( n2043 , n10681 , n5433 );
    xnor g11903 ( n8018 , n11498 , n5766 );
    or g11904 ( n5471 , n1766 , n1532 );
    and g11905 ( n2595 , n6103 , n11603 );
    nor g11906 ( n7290 , n4286 , n8472 );
    or g11907 ( n12881 , n9782 , n7875 );
    or g11908 ( n3767 , n8552 , n3924 );
    xnor g11909 ( n1893 , n9342 , n6052 );
    or g11910 ( n3552 , n1726 , n3718 );
    or g11911 ( n283 , n6373 , n1509 );
    xnor g11912 ( n10946 , n83 , n30 );
    or g11913 ( n2646 , n3875 , n9585 );
    xnor g11914 ( n12812 , n6095 , n781 );
    nor g11915 ( n4158 , n11016 , n3968 );
    not g11916 ( n7691 , n11702 );
    not g11917 ( n2754 , n1198 );
    xnor g11918 ( n8808 , n1278 , n8796 );
    and g11919 ( n6618 , n5767 , n9111 );
    not g11920 ( n3059 , n10181 );
    or g11921 ( n2228 , n10835 , n9280 );
    or g11922 ( n7874 , n989 , n7881 );
    not g11923 ( n12093 , n6050 );
    xnor g11924 ( n4762 , n6575 , n840 );
    and g11925 ( n9841 , n5969 , n1313 );
    nor g11926 ( n10289 , n6113 , n4646 );
    or g11927 ( n7144 , n10157 , n5914 );
    xnor g11928 ( n37 , n9444 , n9291 );
    xnor g11929 ( n9062 , n3570 , n9972 );
    or g11930 ( n8510 , n9370 , n1851 );
    or g11931 ( n2313 , n8428 , n2232 );
    and g11932 ( n5460 , n2722 , n10136 );
    xnor g11933 ( n9012 , n3072 , n4750 );
    nor g11934 ( n1343 , n4591 , n1235 );
    xnor g11935 ( n9204 , n5624 , n1450 );
    and g11936 ( n1844 , n10514 , n11187 );
    or g11937 ( n1514 , n9368 , n809 );
    not g11938 ( n7425 , n8819 );
    or g11939 ( n8514 , n8423 , n7315 );
    or g11940 ( n10908 , n12237 , n5326 );
    xnor g11941 ( n6338 , n4871 , n12090 );
    or g11942 ( n8103 , n5575 , n10919 );
    xnor g11943 ( n4037 , n8596 , n1007 );
    or g11944 ( n9321 , n10142 , n10066 );
    or g11945 ( n9991 , n1719 , n766 );
    xnor g11946 ( n7526 , n11411 , n3856 );
    or g11947 ( n583 , n11923 , n12120 );
    or g11948 ( n9462 , n757 , n3707 );
    xnor g11949 ( n1204 , n8223 , n988 );
    or g11950 ( n1628 , n3407 , n1087 );
    or g11951 ( n422 , n5355 , n561 );
    xnor g11952 ( n6990 , n1306 , n6417 );
    nor g11953 ( n5924 , n12278 , n3853 );
    xnor g11954 ( n8841 , n11547 , n6832 );
    or g11955 ( n4130 , n3680 , n777 );
    xnor g11956 ( n4574 , n2471 , n2662 );
    and g11957 ( n7166 , n4280 , n7970 );
    or g11958 ( n7038 , n12047 , n3803 );
    xnor g11959 ( n10764 , n759 , n10907 );
    xnor g11960 ( n241 , n10309 , n11180 );
    or g11961 ( n3399 , n5530 , n12441 );
    not g11962 ( n862 , n6910 );
    or g11963 ( n6277 , n8510 , n8274 );
    xnor g11964 ( n9564 , n10321 , n6617 );
    or g11965 ( n7909 , n10142 , n5497 );
    nor g11966 ( n9006 , n9627 , n833 );
    xnor g11967 ( n5174 , n1328 , n9359 );
    not g11968 ( n5326 , n521 );
    xnor g11969 ( n4981 , n11703 , n7648 );
    and g11970 ( n5881 , n9520 , n12624 );
    or g11971 ( n2536 , n191 , n7424 );
    or g11972 ( n10297 , n4628 , n7136 );
    or g11973 ( n2741 , n1372 , n1873 );
    and g11974 ( n1756 , n8055 , n3802 );
    and g11975 ( n6208 , n11487 , n4548 );
    and g11976 ( n10236 , n12188 , n11081 );
    and g11977 ( n10640 , n8276 , n3602 );
    not g11978 ( n4936 , n12342 );
    nor g11979 ( n9713 , n3098 , n6711 );
    or g11980 ( n3438 , n5561 , n7682 );
    or g11981 ( n7304 , n4498 , n1162 );
    or g11982 ( n771 , n7449 , n11698 );
    or g11983 ( n5409 , n5858 , n10066 );
    and g11984 ( n7475 , n374 , n10595 );
    and g11985 ( n9175 , n10530 , n1038 );
    or g11986 ( n5981 , n989 , n1079 );
    or g11987 ( n2368 , n5902 , n11827 );
    or g11988 ( n7930 , n2430 , n640 );
    xnor g11989 ( n9384 , n6256 , n7489 );
    or g11990 ( n2602 , n7391 , n7703 );
    not g11991 ( n846 , n1956 );
    or g11992 ( n97 , n2217 , n5502 );
    and g11993 ( n2954 , n7413 , n10998 );
    or g11994 ( n9960 , n12562 , n8048 );
    xnor g11995 ( n3129 , n5995 , n8594 );
    xnor g11996 ( n12593 , n763 , n5979 );
    xnor g11997 ( n12432 , n5793 , n798 );
    or g11998 ( n5599 , n35 , n887 );
    or g11999 ( n3262 , n191 , n11430 );
    or g12000 ( n7394 , n6373 , n9280 );
    xnor g12001 ( n12089 , n3255 , n2398 );
    or g12002 ( n6833 , n1683 , n667 );
    not g12003 ( n10569 , n4210 );
    not g12004 ( n389 , n9925 );
    and g12005 ( n3553 , n4509 , n7930 );
    or g12006 ( n11118 , n9262 , n795 );
    not g12007 ( n1150 , n4168 );
    not g12008 ( n12853 , n137 );
    or g12009 ( n7264 , n3975 , n11321 );
    xnor g12010 ( n5752 , n11779 , n2007 );
    or g12011 ( n11900 , n1572 , n12710 );
    or g12012 ( n11890 , n4059 , n11746 );
    and g12013 ( n8253 , n7202 , n4103 );
    or g12014 ( n9393 , n6750 , n8346 );
    not g12015 ( n752 , n8759 );
    not g12016 ( n12472 , n12343 );
    not g12017 ( n1284 , n3111 );
    xnor g12018 ( n3642 , n8918 , n8764 );
    not g12019 ( n4138 , n9136 );
    and g12020 ( n2953 , n2870 , n6700 );
    not g12021 ( n11652 , n1330 );
    xnor g12022 ( n6095 , n1940 , n8889 );
    xnor g12023 ( n12744 , n6655 , n5827 );
    xnor g12024 ( n4923 , n10989 , n7716 );
    not g12025 ( n10063 , n2897 );
    xnor g12026 ( n3366 , n12066 , n10179 );
    or g12027 ( n8974 , n8026 , n1413 );
    or g12028 ( n3066 , n107 , n10880 );
    and g12029 ( n8142 , n12539 , n4623 );
    xnor g12030 ( n9842 , n10841 , n9560 );
    and g12031 ( n4239 , n8570 , n846 );
    or g12032 ( n12822 , n7088 , n7214 );
    xnor g12033 ( n11242 , n11401 , n2666 );
    and g12034 ( n40 , n12691 , n6543 );
    xnor g12035 ( n12787 , n152 , n9181 );
    and g12036 ( n6123 , n12261 , n3190 );
    or g12037 ( n2887 , n11538 , n8798 );
    and g12038 ( n12280 , n12648 , n7610 );
    or g12039 ( n3362 , n686 , n2232 );
    xnor g12040 ( n808 , n1886 , n12641 );
    or g12041 ( n5425 , n3845 , n10733 );
    xnor g12042 ( n11286 , n5861 , n9994 );
    or g12043 ( n12803 , n12520 , n12307 );
    xnor g12044 ( n8534 , n2343 , n8930 );
    xnor g12045 ( n3981 , n158 , n11961 );
    or g12046 ( n4547 , n6678 , n3267 );
    not g12047 ( n3323 , n8484 );
    not g12048 ( n10003 , n5369 );
    and g12049 ( n1104 , n11821 , n9956 );
    or g12050 ( n2289 , n2677 , n9579 );
    nor g12051 ( n5630 , n11997 , n9582 );
    xnor g12052 ( n4148 , n11895 , n11157 );
    nor g12053 ( n5896 , n3817 , n9276 );
    xnor g12054 ( n3858 , n11772 , n941 );
    xnor g12055 ( n6699 , n9504 , n11910 );
    xnor g12056 ( n11790 , n325 , n2609 );
    or g12057 ( n9343 , n636 , n4913 );
    xnor g12058 ( n11295 , n8578 , n571 );
    or g12059 ( n11005 , n2456 , n5468 );
    xnor g12060 ( n10591 , n6606 , n3582 );
    and g12061 ( n11291 , n7809 , n1095 );
    or g12062 ( n11841 , n639 , n1669 );
    and g12063 ( n9414 , n11829 , n4571 );
    and g12064 ( n9721 , n9834 , n7467 );
    and g12065 ( n990 , n7107 , n12400 );
    and g12066 ( n9089 , n1236 , n9289 );
    xnor g12067 ( n5132 , n4833 , n10496 );
    or g12068 ( n9404 , n9370 , n10419 );
    or g12069 ( n6995 , n9878 , n12080 );
    nor g12070 ( n3529 , n5988 , n10706 );
    and g12071 ( n5845 , n3992 , n9763 );
    xnor g12072 ( n16 , n10292 , n11368 );
    not g12073 ( n8167 , n10322 );
    or g12074 ( n5303 , n1012 , n11537 );
    or g12075 ( n1503 , n8127 , n1162 );
    or g12076 ( n8531 , n962 , n9568 );
    not g12077 ( n1618 , n10941 );
    nor g12078 ( n1376 , n10342 , n12382 );
    or g12079 ( n9566 , n7025 , n8234 );
    xnor g12080 ( n2991 , n6074 , n1400 );
    xnor g12081 ( n12104 , n10694 , n11012 );
    xnor g12082 ( n3792 , n9001 , n1650 );
    or g12083 ( n10548 , n2456 , n7136 );
    nor g12084 ( n6181 , n3864 , n3246 );
    xnor g12085 ( n10445 , n2004 , n11398 );
    and g12086 ( n10538 , n7686 , n6074 );
    not g12087 ( n11989 , n327 );
    or g12088 ( n7487 , n9389 , n1079 );
    and g12089 ( n6353 , n9400 , n10451 );
    or g12090 ( n6743 , n9416 , n12276 );
    xnor g12091 ( n12403 , n6681 , n10894 );
    xnor g12092 ( n11064 , n3845 , n10733 );
    or g12093 ( n5499 , n10196 , n9521 );
    and g12094 ( n850 , n7080 , n10509 );
    xnor g12095 ( n8689 , n1358 , n12462 );
    and g12096 ( n10466 , n12069 , n12489 );
    or g12097 ( n664 , n3944 , n334 );
    and g12098 ( n10972 , n2515 , n2558 );
    and g12099 ( n4291 , n10846 , n5525 );
    xnor g12100 ( n731 , n9308 , n9562 );
    not g12101 ( n3498 , n9321 );
    xnor g12102 ( n361 , n12684 , n3697 );
    xnor g12103 ( n3036 , n803 , n743 );
    xnor g12104 ( n3876 , n72 , n9675 );
    xnor g12105 ( n6131 , n3205 , n12472 );
    xnor g12106 ( n12932 , n3423 , n8948 );
    or g12107 ( n328 , n9370 , n561 );
    xnor g12108 ( n701 , n12834 , n9992 );
    and g12109 ( n10074 , n4480 , n7866 );
    and g12110 ( n12431 , n9791 , n10393 );
    xnor g12111 ( n12460 , n7369 , n4867 );
    not g12112 ( n10581 , n11601 );
    and g12113 ( n11800 , n2680 , n12577 );
    or g12114 ( n4480 , n5530 , n530 );
    or g12115 ( n934 , n11785 , n11284 );
    or g12116 ( n4357 , n9389 , n10419 );
    and g12117 ( n3733 , n2665 , n5931 );
    or g12118 ( n4386 , n5765 , n4527 );
    or g12119 ( n2885 , n4820 , n3789 );
    and g12120 ( n12424 , n3140 , n3447 );
    or g12121 ( n6622 , n1788 , n11990 );
    xnor g12122 ( n12677 , n9027 , n2081 );
    and g12123 ( n11818 , n5200 , n1010 );
    or g12124 ( n8052 , n10750 , n2964 );
    or g12125 ( n9383 , n9878 , n7382 );
    or g12126 ( n4862 , n695 , n2389 );
    not g12127 ( n8092 , n11380 );
    nor g12128 ( n237 , n3206 , n1820 );
    and g12129 ( n5918 , n128 , n5460 );
    nor g12130 ( n4339 , n10168 , n1895 );
    and g12131 ( n2549 , n7469 , n12465 );
    xnor g12132 ( n8439 , n2841 , n7582 );
    or g12133 ( n10575 , n12583 , n10333 );
    or g12134 ( n213 , n1 , n4669 );
    or g12135 ( n11830 , n4125 , n2655 );
    or g12136 ( n8572 , n2447 , n9150 );
    xnor g12137 ( n1364 , n6495 , n2588 );
    xnor g12138 ( n10138 , n8964 , n10120 );
    and g12139 ( n2725 , n1111 , n11177 );
    and g12140 ( n5245 , n11881 , n10053 );
    xnor g12141 ( n7478 , n9529 , n7950 );
    xor g12142 ( n3119 , n7157 , n11079 );
    or g12143 ( n139 , n11034 , n2583 );
    nor g12144 ( n10072 , n6752 , n12017 );
    or g12145 ( n1812 , n762 , n6312 );
    nor g12146 ( n6882 , n794 , n2083 );
    not g12147 ( n10664 , n5603 );
    or g12148 ( n7206 , n191 , n1162 );
    not g12149 ( n686 , n4203 );
    xnor g12150 ( n6379 , n1655 , n3787 );
    not g12151 ( n7161 , n8102 );
    and g12152 ( n7615 , n2984 , n7350 );
    xnor g12153 ( n6736 , n9369 , n2952 );
    and g12154 ( n11045 , n5690 , n1607 );
    xnor g12155 ( n9019 , n12139 , n8043 );
    or g12156 ( n8588 , n5945 , n9741 );
    xnor g12157 ( n3232 , n7304 , n11017 );
    xnor g12158 ( n9678 , n182 , n11549 );
    xnor g12159 ( n11462 , n2349 , n4308 );
    or g12160 ( n8805 , n3746 , n3468 );
    or g12161 ( n2829 , n11661 , n6279 );
    or g12162 ( n11574 , n6921 , n8812 );
    not g12163 ( n9978 , n12506 );
    or g12164 ( n12906 , n10879 , n1079 );
    nor g12165 ( n11444 , n8156 , n6908 );
    or g12166 ( n1197 , n11923 , n28 );
    and g12167 ( n287 , n10361 , n6305 );
    or g12168 ( n4117 , n5007 , n2377 );
    nor g12169 ( n5216 , n11873 , n1758 );
    or g12170 ( n1423 , n9652 , n9798 );
    and g12171 ( n5972 , n5102 , n10400 );
    xnor g12172 ( n9601 , n6446 , n10660 );
    and g12173 ( n5262 , n2491 , n3725 );
    xnor g12174 ( n3799 , n5796 , n9673 );
    xnor g12175 ( n10457 , n6920 , n1262 );
    not g12176 ( n1630 , n3478 );
    not g12177 ( n8173 , n7012 );
    not g12178 ( n674 , n10777 );
    nor g12179 ( n9873 , n4196 , n11519 );
    or g12180 ( n3445 , n9271 , n1866 );
    xnor g12181 ( n5142 , n639 , n88 );
    or g12182 ( n12707 , n7283 , n7246 );
    xnor g12183 ( n728 , n9069 , n5785 );
    or g12184 ( n5996 , n1802 , n1869 );
    xnor g12185 ( n12457 , n3528 , n4944 );
    xnor g12186 ( n10551 , n733 , n682 );
    not g12187 ( n7167 , n9942 );
    xnor g12188 ( n12855 , n4711 , n10822 );
    or g12189 ( n11654 , n9140 , n3592 );
    not g12190 ( n4934 , n11164 );
    not g12191 ( n11367 , n10862 );
    not g12192 ( n12596 , n11099 );
    or g12193 ( n7464 , n636 , n1163 );
    xnor g12194 ( n4292 , n8672 , n4538 );
    or g12195 ( n5149 , n12361 , n5538 );
    not g12196 ( n4913 , n1512 );
    or g12197 ( n452 , n5530 , n2259 );
    or g12198 ( n8056 , n9380 , n1671 );
    and g12199 ( n3517 , n5042 , n125 );
    xor g12200 ( n4786 , n12234 , n9814 );
    not g12201 ( n8753 , n5930 );
    xor g12202 ( n4218 , n5189 , n8537 );
    or g12203 ( n6 , n6577 , n5540 );
    or g12204 ( n4431 , n11433 , n1413 );
    not g12205 ( n5751 , n12370 );
    not g12206 ( n1432 , n9499 );
    not g12207 ( n2997 , n3559 );
    and g12208 ( n7670 , n11931 , n10576 );
    xnor g12209 ( n9039 , n12284 , n7329 );
    and g12210 ( n8485 , n3506 , n2724 );
    or g12211 ( n12026 , n12585 , n1077 );
    not g12212 ( n2049 , n1850 );
    xnor g12213 ( n8627 , n3708 , n11253 );
    nor g12214 ( n8922 , n9611 , n6178 );
    xnor g12215 ( n3915 , n8321 , n13 );
    nor g12216 ( n4566 , n9282 , n5464 );
    xnor g12217 ( n5796 , n5823 , n565 );
    xnor g12218 ( n5187 , n5200 , n12395 );
    xnor g12219 ( n1647 , n9806 , n9164 );
    not g12220 ( n6906 , n11132 );
    xnor g12221 ( n6280 , n7018 , n6735 );
    nor g12222 ( n11848 , n9497 , n10472 );
    and g12223 ( n9768 , n8619 , n2746 );
    not g12224 ( n8954 , n7882 );
    nor g12225 ( n379 , n10973 , n3590 );
    xnor g12226 ( n10155 , n3087 , n511 );
    and g12227 ( n4143 , n4206 , n4303 );
    or g12228 ( n12040 , n3096 , n10903 );
    xnor g12229 ( n7374 , n9605 , n2566 );
    or g12230 ( n3930 , n2099 , n3924 );
    or g12231 ( n12692 , n3096 , n5540 );
    xnor g12232 ( n3446 , n12108 , n1818 );
    nor g12233 ( n3778 , n11926 , n6362 );
    and g12234 ( n10894 , n3290 , n2989 );
    not g12235 ( n8428 , n9400 );
    not g12236 ( n5914 , n2507 );
    or g12237 ( n735 , n11699 , n6262 );
    and g12238 ( n1458 , n9085 , n5071 );
    and g12239 ( n4487 , n2618 , n1654 );
    nor g12240 ( n4541 , n6891 , n8455 );
    nor g12241 ( n5428 , n8762 , n12509 );
    and g12242 ( n7450 , n7154 , n10837 );
    xnor g12243 ( n471 , n5589 , n11291 );
    or g12244 ( n2337 , n6977 , n8768 );
    xnor g12245 ( n12436 , n9840 , n3238 );
    and g12246 ( n8021 , n78 , n1934 );
    not g12247 ( n2406 , n7285 );
    xnor g12248 ( n11920 , n11942 , n11765 );
    or g12249 ( n6146 , n8026 , n5540 );
    xnor g12250 ( n12516 , n5757 , n5726 );
    or g12251 ( n7310 , n10750 , n3924 );
    xnor g12252 ( n4968 , n7743 , n10967 );
    and g12253 ( n11996 , n4515 , n6220 );
    xor g12254 ( n4155 , n2209 , n7039 );
    xnor g12255 ( n8039 , n2279 , n7754 );
    not g12256 ( n11511 , n9883 );
    or g12257 ( n3126 , n7449 , n8643 );
    xnor g12258 ( n5790 , n10573 , n6026 );
    and g12259 ( n3336 , n2116 , n10426 );
    nor g12260 ( n9899 , n10148 , n7996 );
    or g12261 ( n8033 , n11719 , n1162 );
    xnor g12262 ( n7539 , n5264 , n11803 );
    or g12263 ( n11604 , n6175 , n8316 );
    xnor g12264 ( n11351 , n5052 , n5478 );
    and g12265 ( n4427 , n5817 , n2053 );
    or g12266 ( n11047 , n5959 , n8534 );
    not g12267 ( n1413 , n9640 );
    xnor g12268 ( n9587 , n4241 , n7699 );
    not g12269 ( n294 , n6945 );
    xnor g12270 ( n10728 , n8343 , n5706 );
    or g12271 ( n5211 , n11968 , n6 );
    not g12272 ( n11374 , n12734 );
    or g12273 ( n3447 , n994 , n7246 );
    and g12274 ( n1083 , n2936 , n10198 );
    or g12275 ( n9468 , n11898 , n1924 );
    or g12276 ( n1018 , n4151 , n3840 );
    xnor g12277 ( n3312 , n390 , n2483 );
    xnor g12278 ( n7073 , n5714 , n7985 );
    xnor g12279 ( n10610 , n11590 , n2778 );
    and g12280 ( n3171 , n2128 , n12801 );
    or g12281 ( n509 , n6066 , n5292 );
    xnor g12282 ( n9627 , n3960 , n6775 );
    xnor g12283 ( n4871 , n12858 , n8742 );
    and g12284 ( n8557 , n2134 , n6988 );
    nor g12285 ( n5686 , n8176 , n2388 );
    xnor g12286 ( n7165 , n8012 , n9789 );
    xnor g12287 ( n617 , n2739 , n3369 );
    or g12288 ( n7598 , n103 , n7134 );
    not g12289 ( n9144 , n3754 );
    nor g12290 ( n10824 , n641 , n11230 );
    and g12291 ( n8829 , n2111 , n7841 );
    xnor g12292 ( n5343 , n10354 , n1502 );
    xnor g12293 ( n3921 , n4381 , n26 );
    or g12294 ( n9746 , n10750 , n8259 );
    xnor g12295 ( n277 , n3680 , n8031 );
    xnor g12296 ( n2614 , n6740 , n9524 );
    xnor g12297 ( n10428 , n505 , n854 );
    or g12298 ( n9378 , n3739 , n9722 );
    not g12299 ( n3324 , n7646 );
    xnor g12300 ( n12351 , n2265 , n7026 );
    xnor g12301 ( n11148 , n5874 , n7387 );
    xnor g12302 ( n9610 , n10955 , n5648 );
    or g12303 ( n6553 , n11958 , n6169 );
    nor g12304 ( n4916 , n6128 , n8784 );
    xnor g12305 ( n9391 , n9473 , n3292 );
    and g12306 ( n10011 , n8839 , n10927 );
    and g12307 ( n5647 , n5203 , n9780 );
    and g12308 ( n3411 , n4931 , n4459 );
    not g12309 ( n965 , n6008 );
    or g12310 ( n5394 , n2456 , n12080 );
    not g12311 ( n10691 , n12716 );
    xnor g12312 ( n9334 , n8767 , n1974 );
    or g12313 ( n178 , n5355 , n6524 );
    and g12314 ( n6410 , n8108 , n101 );
    not g12315 ( n4839 , n5159 );
    or g12316 ( n4956 , n12119 , n8648 );
    or g12317 ( n11556 , n994 , n2358 );
    not g12318 ( n11070 , n5570 );
    nor g12319 ( n5312 , n11500 , n11725 );
    and g12320 ( n6265 , n12217 , n4608 );
    not g12321 ( n7630 , n10005 );
    not g12322 ( n4215 , n12600 );
    or g12323 ( n6761 , n7729 , n2303 );
    and g12324 ( n10525 , n5249 , n10356 );
    nor g12325 ( n3037 , n12937 , n2339 );
    and g12326 ( n7519 , n2336 , n3775 );
    xnor g12327 ( n363 , n8224 , n6397 );
    or g12328 ( n10684 , n7097 , n9115 );
    xnor g12329 ( n559 , n1015 , n10240 );
    and g12330 ( n8731 , n1665 , n10889 );
    or g12331 ( n8070 , n10157 , n5258 );
    nor g12332 ( n9336 , n2565 , n1322 );
    or g12333 ( n1824 , n1929 , n2485 );
    xnor g12334 ( n12897 , n9448 , n10248 );
    xnor g12335 ( n9365 , n57 , n9099 );
    or g12336 ( n10171 , n5915 , n1163 );
    xnor g12337 ( n2239 , n9788 , n362 );
    not g12338 ( n3781 , n5166 );
    nor g12339 ( n10039 , n10812 , n5744 );
    and g12340 ( n3313 , n8611 , n9015 );
    xnor g12341 ( n9903 , n9177 , n9386 );
    not g12342 ( n8488 , n11354 );
    xnor g12343 ( n12259 , n8492 , n5296 );
    or g12344 ( n2245 , n5942 , n8925 );
    xnor g12345 ( n1273 , n9688 , n8446 );
    xnor g12346 ( n12608 , n7957 , n9592 );
    not g12347 ( n10390 , n6629 );
    and g12348 ( n9562 , n11722 , n10186 );
    xnor g12349 ( n1304 , n3851 , n11091 );
    and g12350 ( n8192 , n7287 , n8860 );
    and g12351 ( n6320 , n5720 , n6565 );
    not g12352 ( n7435 , n6583 );
    or g12353 ( n11313 , n8197 , n1098 );
    or g12354 ( n6876 , n3768 , n1611 );
    and g12355 ( n2937 , n1229 , n6905 );
    nor g12356 ( n8161 , n10233 , n1965 );
    or g12357 ( n421 , n9893 , n2553 );
    xnor g12358 ( n3444 , n11440 , n8128 );
    or g12359 ( n9474 , n6059 , n8862 );
    and g12360 ( n3567 , n2124 , n3553 );
    or g12361 ( n11152 , n3612 , n12676 );
    nor g12362 ( n5464 , n8915 , n3956 );
    xnor g12363 ( n8992 , n7126 , n5154 );
    or g12364 ( n8291 , n3126 , n188 );
    xnor g12365 ( n5294 , n9435 , n7535 );
    and g12366 ( n12805 , n6028 , n9435 );
    or g12367 ( n8164 , n2866 , n4742 );
    nor g12368 ( n6675 , n1992 , n12212 );
    xnor g12369 ( n3245 , n9301 , n12244 );
    or g12370 ( n12083 , n1083 , n6613 );
    xnor g12371 ( n2939 , n5559 , n9735 );
    and g12372 ( n10325 , n1444 , n3951 );
    not g12373 ( n11733 , n5450 );
    or g12374 ( n10239 , n2400 , n2705 );
    and g12375 ( n12952 , n7298 , n1325 );
    xnor g12376 ( n153 , n2385 , n8884 );
    or g12377 ( n11799 , n5679 , n2963 );
    not g12378 ( n3660 , n9242 );
    xnor g12379 ( n4210 , n10138 , n7773 );
    and g12380 ( n627 , n8535 , n2410 );
    nor g12381 ( n3010 , n1461 , n3374 );
    nor g12382 ( n10885 , n12766 , n4704 );
    not g12383 ( n9191 , n5276 );
    nor g12384 ( n11516 , n8994 , n3041 );
    nor g12385 ( n8126 , n785 , n3177 );
    xnor g12386 ( n5256 , n11130 , n3871 );
    and g12387 ( n7922 , n9400 , n6703 );
    not g12388 ( n5054 , n4010 );
    or g12389 ( n4335 , n7004 , n3319 );
    xnor g12390 ( n10707 , n11266 , n8286 );
    xnor g12391 ( n10837 , n6096 , n9191 );
    xnor g12392 ( n65 , n2388 , n10264 );
    or g12393 ( n12647 , n10951 , n9916 );
    xnor g12394 ( n2411 , n7114 , n44 );
    xnor g12395 ( n11954 , n3931 , n8047 );
    xnor g12396 ( n10380 , n12302 , n2462 );
    or g12397 ( n4222 , n11759 , n6154 );
    or g12398 ( n817 , n7391 , n11827 );
    xnor g12399 ( n930 , n3350 , n10262 );
    xnor g12400 ( n9362 , n6198 , n12567 );
    xnor g12401 ( n787 , n9689 , n7040 );
    nor g12402 ( n9418 , n9364 , n1458 );
    xor g12403 ( n8939 , n2660 , n12812 );
    or g12404 ( n8230 , n7378 , n5188 );
    or g12405 ( n12532 , n1941 , n7425 );
    or g12406 ( n11424 , n7192 , n7696 );
    xnor g12407 ( n598 , n343 , n4062 );
    or g12408 ( n12006 , n7495 , n1079 );
    or g12409 ( n3919 , n1937 , n1413 );
    nor g12410 ( n7049 , n2560 , n6965 );
    xnor g12411 ( n10984 , n7870 , n2341 );
    or g12412 ( n502 , n8287 , n1196 );
    and g12413 ( n4706 , n11743 , n12004 );
    or g12414 ( n2284 , n6977 , n7395 );
    xnor g12415 ( n1921 , n12281 , n4939 );
    xor g12416 ( n6014 , n1177 , n1645 );
    not g12417 ( n619 , n147 );
    xnor g12418 ( n2501 , n910 , n9852 );
    or g12419 ( n1766 , n9373 , n9160 );
    and g12420 ( n8885 , n12813 , n946 );
    or g12421 ( n11415 , n3746 , n6197 );
    xnor g12422 ( n7280 , n7225 , n5070 );
    or g12423 ( n4633 , n5168 , n8997 );
    not g12424 ( n3638 , n3509 );
    not g12425 ( n2456 , n11478 );
    xnor g12426 ( n12204 , n8126 , n2692 );
    or g12427 ( n3431 , n8026 , n2232 );
    or g12428 ( n8416 , n1699 , n3924 );
    nor g12429 ( n11713 , n5843 , n10236 );
    xnor g12430 ( n623 , n4368 , n7543 );
    or g12431 ( n11965 , n714 , n3537 );
    and g12432 ( n8923 , n5219 , n4926 );
    xnor g12433 ( n4114 , n10165 , n2276 );
    or g12434 ( n8895 , n10683 , n2527 );
    xnor g12435 ( n12645 , n5290 , n11551 );
    xnor g12436 ( n8661 , n10852 , n11134 );
    or g12437 ( n4041 , n6577 , n1413 );
    not g12438 ( n5540 , n7500 );
    or g12439 ( n7438 , n10717 , n7042 );
    xnor g12440 ( n11932 , n6473 , n1194 );
    nor g12441 ( n2494 , n140 , n9737 );
    or g12442 ( n2596 , n12366 , n1366 );
    or g12443 ( n8597 , n5024 , n2044 );
    not g12444 ( n981 , n1629 );
    and g12445 ( n9611 , n1834 , n11175 );
    or g12446 ( n12752 , n12525 , n3298 );
    nor g12447 ( n2444 , n10361 , n6305 );
    nor g12448 ( n10260 , n163 , n1093 );
    xnor g12449 ( n7460 , n1821 , n391 );
    xnor g12450 ( n12232 , n3430 , n579 );
    and g12451 ( n645 , n6847 , n11002 );
    not g12452 ( n8171 , n6706 );
    or g12453 ( n3469 , n7495 , n11746 );
    xnor g12454 ( n7350 , n1460 , n12415 );
    and g12455 ( n8162 , n12712 , n9872 );
    or g12456 ( n2608 , n10835 , n6922 );
    and g12457 ( n11911 , n4283 , n5524 );
    or g12458 ( n7792 , n7839 , n7876 );
    or g12459 ( n4549 , n2877 , n572 );
    or g12460 ( n11318 , n3743 , n5086 );
    or g12461 ( n2136 , n10157 , n1047 );
    or g12462 ( n7010 , n7654 , n4482 );
    xnor g12463 ( n11339 , n12386 , n9257 );
    xnor g12464 ( n797 , n12557 , n1270 );
    xnor g12465 ( n1336 , n12846 , n7514 );
    xnor g12466 ( n5128 , n5688 , n10758 );
    or g12467 ( n3955 , n1805 , n7072 );
    nor g12468 ( n12566 , n4281 , n10380 );
    and g12469 ( n5417 , n4717 , n12302 );
    or g12470 ( n10721 , n3141 , n4721 );
    or g12471 ( n1309 , n9878 , n6513 );
    xnor g12472 ( n12101 , n3959 , n2008 );
    or g12473 ( n5049 , n10142 , n9397 );
    and g12474 ( n7685 , n12069 , n12925 );
    xnor g12475 ( n8747 , n1445 , n3815 );
    not g12476 ( n2325 , n4597 );
    xnor g12477 ( n31 , n7469 , n6723 );
    xnor g12478 ( n9767 , n12420 , n4309 );
    or g12479 ( n11881 , n11221 , n3260 );
    or g12480 ( n9223 , n5915 , n7928 );
    not g12481 ( n4051 , n5900 );
    xnor g12482 ( n3430 , n10936 , n3631 );
    xnor g12483 ( n9231 , n8803 , n12304 );
    nor g12484 ( n7582 , n7945 , n12927 );
    xnor g12485 ( n4455 , n10338 , n6123 );
    xnor g12486 ( n2495 , n9951 , n1649 );
    nor g12487 ( n12726 , n5278 , n922 );
    nor g12488 ( n659 , n6157 , n3657 );
    xnor g12489 ( n12463 , n12505 , n4196 );
    xnor g12490 ( n939 , n2222 , n8638 );
    not g12491 ( n12367 , n312 );
    not g12492 ( n7470 , n7248 );
    and g12493 ( n6744 , n386 , n9354 );
    or g12494 ( n11582 , n5196 , n8731 );
    xnor g12495 ( n716 , n12548 , n980 );
    nor g12496 ( n8473 , n7694 , n12015 );
    xnor g12497 ( n8287 , n951 , n9151 );
    and g12498 ( n605 , n8389 , n11484 );
    and g12499 ( n1918 , n4250 , n7101 );
    or g12500 ( n3104 , n8261 , n12473 );
    and g12501 ( n11754 , n12764 , n4834 );
    or g12502 ( n4160 , n3617 , n8109 );
    not g12503 ( n1051 , n8276 );
    xnor g12504 ( n1550 , n10504 , n6682 );
    or g12505 ( n7593 , n11142 , n10187 );
    and g12506 ( n11783 , n6463 , n12738 );
    or g12507 ( n7133 , n2099 , n1932 );
    or g12508 ( n2059 , n12103 , n9593 );
    xnor g12509 ( n6620 , n2835 , n4033 );
    not g12510 ( n6456 , n4732 );
    xnor g12511 ( n4412 , n3222 , n12228 );
    xnor g12512 ( n1017 , n10976 , n4526 );
    not g12513 ( n3028 , n7486 );
    xnor g12514 ( n7017 , n4161 , n4888 );
    and g12515 ( n3057 , n2312 , n3899 );
    and g12516 ( n12103 , n8818 , n6967 );
    nor g12517 ( n5939 , n5947 , n9539 );
    and g12518 ( n8134 , n10678 , n6703 );
    xnor g12519 ( n10491 , n4879 , n4157 );
    xor g12520 ( n7579 , n3918 , n4922 );
    or g12521 ( n58 , n11958 , n7952 );
    or g12522 ( n12217 , n4536 , n4220 );
    and g12523 ( n12619 , n21 , n10600 );
    and g12524 ( n3137 , n5269 , n12488 );
    xnor g12525 ( n3654 , n1570 , n4680 );
    not g12526 ( n8078 , n11482 );
    and g12527 ( n3634 , n8733 , n5632 );
    not g12528 ( n2297 , n4490 );
    or g12529 ( n1462 , n191 , n561 );
    or g12530 ( n318 , n11923 , n4654 );
    or g12531 ( n2610 , n994 , n8524 );
    or g12532 ( n5154 , n114 , n5540 );
    xnor g12533 ( n5892 , n9107 , n2986 );
    or g12534 ( n10178 , n2099 , n5468 );
    or g12535 ( n6086 , n636 , n4818 );
    not g12536 ( n5655 , n4908 );
    or g12537 ( n10763 , n1665 , n10889 );
    xnor g12538 ( n3790 , n7094 , n3900 );
    or g12539 ( n1689 , n12237 , n8740 );
    xnor g12540 ( n12248 , n9869 , n11852 );
    xnor g12541 ( n11765 , n5213 , n6533 );
    not g12542 ( n12587 , n7827 );
    nor g12543 ( n914 , n8580 , n12078 );
    or g12544 ( n2906 , n636 , n12535 );
    and g12545 ( n7492 , n7014 , n5176 );
    not g12546 ( n6671 , n10976 );
    or g12547 ( n12440 , n1937 , n11410 );
    or g12548 ( n5089 , n2099 , n12080 );
    and g12549 ( n6040 , n1988 , n10674 );
    or g12550 ( n2837 , n12119 , n12124 );
    and g12551 ( n4115 , n357 , n5306 );
    and g12552 ( n2661 , n5954 , n7486 );
    or g12553 ( n5891 , n5861 , n9506 );
    or g12554 ( n1313 , n10339 , n3224 );
    not g12555 ( n8583 , n996 );
    and g12556 ( n10021 , n616 , n2258 );
    or g12557 ( n6180 , n5765 , n5914 );
    or g12558 ( n9522 , n114 , n12816 );
    not g12559 ( n6513 , n12489 );
    or g12560 ( n3667 , n9389 , n10066 );
    not g12561 ( n3096 , n1094 );
    not g12562 ( n1761 , n2235 );
    or g12563 ( n5145 , n3959 , n2008 );
    and g12564 ( n9425 , n9301 , n2028 );
    xnor g12565 ( n5785 , n3535 , n11795 );
    and g12566 ( n3742 , n12648 , n11922 );
    xnor g12567 ( n2926 , n6924 , n12527 );
    xnor g12568 ( n6573 , n12264 , n11385 );
    or g12569 ( n420 , n10142 , n510 );
    and g12570 ( n2992 , n8782 , n4555 );
    xnor g12571 ( n12206 , n4972 , n12167 );
    or g12572 ( n7485 , n10625 , n11701 );
    and g12573 ( n10241 , n413 , n7955 );
    and g12574 ( n10976 , n6255 , n11481 );
    and g12575 ( n11180 , n509 , n10385 );
    and g12576 ( n6267 , n2036 , n2853 );
    xnor g12577 ( n3576 , n12592 , n10428 );
    or g12578 ( n3845 , n8959 , n995 );
    xnor g12579 ( n2755 , n5730 , n4428 );
    xnor g12580 ( n8568 , n9496 , n1775 );
    nor g12581 ( n2266 , n2104 , n7321 );
    and g12582 ( n3588 , n7388 , n10990 );
    and g12583 ( n7749 , n8397 , n9700 );
    nor g12584 ( n2868 , n6759 , n3694 );
    and g12585 ( n7845 , n385 , n6108 );
    and g12586 ( n714 , n5963 , n4102 );
    and g12587 ( n4664 , n1822 , n8375 );
    not g12588 ( n12711 , n9712 );
    and g12589 ( n11898 , n6486 , n1464 );
    nor g12590 ( n9118 , n11192 , n1901 );
    xnor g12591 ( n10524 , n8015 , n11946 );
    or g12592 ( n3464 , n752 , n6114 );
    or g12593 ( n10969 , n7053 , n7346 );
    xnor g12594 ( n121 , n11515 , n8271 );
    and g12595 ( n8072 , n2018 , n10383 );
    or g12596 ( n1951 , n12560 , n6040 );
    and g12597 ( n1805 , n8313 , n879 );
    and g12598 ( n5363 , n2393 , n2749 );
    nor g12599 ( n631 , n7846 , n4955 );
    and g12600 ( n624 , n8988 , n8804 );
    and g12601 ( n11699 , n8836 , n3941 );
    and g12602 ( n9429 , n5974 , n4471 );
    not g12603 ( n568 , n5053 );
    and g12604 ( n11186 , n2626 , n4041 );
    not g12605 ( n1554 , n11747 );
    and g12606 ( n4026 , n5023 , n4063 );
    nor g12607 ( n9461 , n927 , n2180 );
    and g12608 ( n1869 , n10601 , n3576 );
    or g12609 ( n4214 , n11144 , n2139 );
    and g12610 ( n3179 , n11222 , n8433 );
    xnor g12611 ( n10322 , n1365 , n7787 );
    xnor g12612 ( n776 , n1449 , n1174 );
    or g12613 ( n1143 , n8687 , n12771 );
    or g12614 ( n6152 , n8405 , n826 );
    nor g12615 ( n1219 , n3133 , n10313 );
    not g12616 ( n371 , n11370 );
    not g12617 ( n10478 , n1999 );
    or g12618 ( n7044 , n9240 , n11264 );
    nor g12619 ( n12393 , n5185 , n5410 );
    xnor g12620 ( n7529 , n97 , n3891 );
    or g12621 ( n222 , n6347 , n9890 );
    xnor g12622 ( n3136 , n3298 , n5952 );
    xnor g12623 ( n6018 , n697 , n1295 );
    or g12624 ( n5674 , n8757 , n3021 );
    not g12625 ( n9671 , n5972 );
    xnor g12626 ( n1665 , n8533 , n6193 );
    xnor g12627 ( n12076 , n8958 , n1551 );
    and g12628 ( n3346 , n1129 , n4967 );
    xnor g12629 ( n8941 , n8694 , n2582 );
    not g12630 ( n5680 , n12242 );
    xnor g12631 ( n11513 , n4213 , n986 );
    or g12632 ( n7662 , n11923 , n3606 );
    nor g12633 ( n6380 , n6150 , n5921 );
    not g12634 ( n9561 , n7146 );
    and g12635 ( n6816 , n11007 , n1253 );
    or g12636 ( n7858 , n11623 , n7632 );
    xnor g12637 ( n10230 , n12906 , n9889 );
    not g12638 ( n10244 , n2990 );
    not g12639 ( n12039 , n10051 );
    and g12640 ( n11453 , n4759 , n1569 );
    not g12641 ( n8518 , n2244 );
    xnor g12642 ( n4008 , n3712 , n10986 );
    nor g12643 ( n7675 , n12872 , n10586 );
    and g12644 ( n3247 , n11085 , n486 );
    nor g12645 ( n7025 , n12493 , n3785 );
    xnor g12646 ( n11617 , n10863 , n4245 );
    and g12647 ( n1543 , n1399 , n965 );
    xnor g12648 ( n293 , n5101 , n1178 );
    or g12649 ( n4985 , n3623 , n8591 );
    not g12650 ( n3694 , n10805 );
    xnor g12651 ( n6778 , n6590 , n11930 );
    xnor g12652 ( n6593 , n1682 , n9303 );
    xnor g12653 ( n4171 , n3444 , n1692 );
    or g12654 ( n6519 , n7391 , n6402 );
    or g12655 ( n12496 , n238 , n1813 );
    xnor g12656 ( n11155 , n9556 , n3043 );
    nor g12657 ( n8767 , n11436 , n8632 );
    xnor g12658 ( n10807 , n4116 , n3310 );
    and g12659 ( n12163 , n4187 , n11728 );
    and g12660 ( n1571 , n8201 , n3922 );
    not g12661 ( n9813 , n1493 );
    not g12662 ( n6091 , n10012 );
    or g12663 ( n7258 , n10587 , n10140 );
    and g12664 ( n10150 , n11138 , n10218 );
    not g12665 ( n9971 , n10217 );
    or g12666 ( n6090 , n11923 , n795 );
    or g12667 ( n2312 , n9373 , n1047 );
    or g12668 ( n4301 , n4911 , n1079 );
    and g12669 ( n249 , n7747 , n6311 );
    and g12670 ( n9099 , n3940 , n9740 );
    or g12671 ( n6466 , n3324 , n2020 );
    xnor g12672 ( n2131 , n6848 , n12077 );
    xnor g12673 ( n8616 , n10141 , n2223 );
    xnor g12674 ( n12037 , n10366 , n11185 );
    and g12675 ( n2439 , n3618 , n3793 );
    xnor g12676 ( n758 , n7234 , n9234 );
    or g12677 ( n6374 , n191 , n7389 );
    or g12678 ( n2346 , n5199 , n3121 );
    nor g12679 ( n4865 , n9403 , n11100 );
    and g12680 ( n12395 , n970 , n2165 );
    or g12681 ( n9698 , n8870 , n4818 );
    and g12682 ( n7471 , n3220 , n9239 );
    xnor g12683 ( n407 , n10646 , n10375 );
    not g12684 ( n6057 , n12463 );
    or g12685 ( n9290 , n7283 , n8859 );
    and g12686 ( n4742 , n6491 , n4169 );
    xnor g12687 ( n2304 , n12289 , n9253 );
    not g12688 ( n6957 , n3346 );
    and g12689 ( n2850 , n5456 , n87 );
    xnor g12690 ( n3196 , n11807 , n6092 );
    xnor g12691 ( n8913 , n6799 , n4772 );
    not g12692 ( n11952 , n9828 );
    and g12693 ( n9896 , n7862 , n5212 );
    xnor g12694 ( n5100 , n2435 , n10995 );
    and g12695 ( n1765 , n8671 , n9485 );
    and g12696 ( n9098 , n6554 , n5201 );
    xnor g12697 ( n12161 , n5794 , n4340 );
    or g12698 ( n6216 , n8428 , n9971 );
    not g12699 ( n8699 , n8027 );
    or g12700 ( n11670 , n5601 , n8237 );
    not g12701 ( n11018 , n8134 );
    and g12702 ( n4552 , n7750 , n8004 );
    or g12703 ( n736 , n779 , n456 );
    or g12704 ( n11578 , n7495 , n7881 );
endmodule
