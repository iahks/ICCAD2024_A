// Benchmark "top_809568696_809776567_809698999_863110837_1234615" written by ABC on Mon Aug 19 00:27:34 2024

module top_809568696_809776567_809698999_863110837_1234615 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128;
  wire new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1910, new_n1911, new_n1912,
    new_n1913, new_n1914, new_n1915, new_n1916, new_n1917, new_n1918,
    new_n1919, new_n1920, new_n1921, new_n1922, new_n1923, new_n1924,
    new_n1925, new_n1926, new_n1927, new_n1928, new_n1929, new_n1930,
    new_n1931, new_n1932, new_n1933, new_n1934, new_n1935, new_n1936,
    new_n1937, new_n1938, new_n1939, new_n1940, new_n1941, new_n1942,
    new_n1943, new_n1944, new_n1945, new_n1946, new_n1947, new_n1948,
    new_n1949, new_n1950, new_n1951, new_n1952, new_n1953, new_n1954,
    new_n1955, new_n1957, new_n1958, new_n1959, new_n1960, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2093, new_n2094, new_n2095, new_n2096,
    new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102,
    new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132,
    new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144,
    new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150,
    new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2156,
    new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2281, new_n2282, new_n2283, new_n2284,
    new_n2285, new_n2286, new_n2287, new_n2288, new_n2289, new_n2290,
    new_n2291, new_n2292, new_n2293, new_n2294, new_n2295, new_n2296,
    new_n2297, new_n2298, new_n2299, new_n2300, new_n2301, new_n2302,
    new_n2303, new_n2304, new_n2305, new_n2307, new_n2308, new_n2309,
    new_n2310, new_n2311, new_n2312, new_n2313, new_n2314, new_n2315,
    new_n2316, new_n2317, new_n2318, new_n2319, new_n2320, new_n2321,
    new_n2322, new_n2323, new_n2324, new_n2325, new_n2326, new_n2327,
    new_n2328, new_n2329, new_n2330, new_n2331, new_n2332, new_n2333,
    new_n2334, new_n2335, new_n2336, new_n2337, new_n2338, new_n2339,
    new_n2340, new_n2341, new_n2342, new_n2343, new_n2344, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2423, new_n2424, new_n2425, new_n2426, new_n2427, new_n2428,
    new_n2429, new_n2430, new_n2431, new_n2432, new_n2433, new_n2434,
    new_n2435, new_n2436, new_n2438, new_n2439, new_n2440, new_n2441,
    new_n2442, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460,
    new_n2461, new_n2462, new_n2463, new_n2465, new_n2466, new_n2468,
    new_n2469, new_n2470, new_n2472, new_n2474, new_n2475, new_n2476,
    new_n2477, new_n2478, new_n2479, new_n2480, new_n2481, new_n2482,
    new_n2484, new_n2485, new_n2486, new_n2487, new_n2488, new_n2489,
    new_n2491, new_n2492, new_n2493, new_n2494, new_n2496, new_n2497,
    new_n2498, new_n2499, new_n2500, new_n2501, new_n2502, new_n2503,
    new_n2504, new_n2505, new_n2506, new_n2507, new_n2508, new_n2509,
    new_n2510, new_n2511, new_n2512, new_n2513, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2552, new_n2553, new_n2554,
    new_n2555, new_n2557, new_n2558, new_n2559, new_n2562, new_n2563,
    new_n2564, new_n2565, new_n2566, new_n2568, new_n2570, new_n2571,
    new_n2573, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578,
    new_n2579, new_n2580, new_n2581, new_n2582, new_n2583, new_n2584,
    new_n2585, new_n2586, new_n2587, new_n2588, new_n2589, new_n2590,
    new_n2591, new_n2592, new_n2594, new_n2595, new_n2597, new_n2598,
    new_n2599, new_n2600, new_n2601, new_n2603, new_n2604, new_n2605,
    new_n2606, new_n2607, new_n2608, new_n2609, new_n2610, new_n2611,
    new_n2612, new_n2613, new_n2614, new_n2615, new_n2616, new_n2617,
    new_n2618, new_n2619, new_n2620, new_n2622, new_n2623, new_n2624,
    new_n2626, new_n2627, new_n2629, new_n2630, new_n2631, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2646,
    new_n2647, new_n2648, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2674, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679,
    new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685,
    new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2692,
    new_n2693, new_n2694, new_n2697, new_n2698, new_n2699, new_n2700,
    new_n2701, new_n2702, new_n2703, new_n2704, new_n2705, new_n2706,
    new_n2707, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2719, new_n2720, new_n2721,
    new_n2722, new_n2723, new_n2724, new_n2725, new_n2726, new_n2727,
    new_n2728, new_n2729, new_n2730, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2738, new_n2739, new_n2740, new_n2742,
    new_n2743, new_n2744, new_n2746, new_n2747, new_n2749, new_n2750,
    new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2783,
    new_n2784, new_n2785, new_n2787, new_n2788, new_n2790, new_n2791,
    new_n2793, new_n2794, new_n2795, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2813, new_n2814,
    new_n2815, new_n2816, new_n2817, new_n2818, new_n2819, new_n2821,
    new_n2823, new_n2825, new_n2826, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2841, new_n2842, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2854, new_n2855, new_n2856, new_n2859,
    new_n2860, new_n2862, new_n2863, new_n2864, new_n2866, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2873, new_n2874, new_n2877,
    new_n2878, new_n2880, new_n2882, new_n2884, new_n2886, new_n2887,
    new_n2889, new_n2890, new_n2892, new_n2893, new_n2894, new_n2895,
    new_n2897, new_n2899, new_n2900, new_n2903, new_n2904, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2911, new_n2912, new_n2915,
    new_n2916, new_n2918, new_n2919, new_n2921, new_n2923, new_n2924,
    new_n2925, new_n2928, new_n2929, new_n2931, new_n2932, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2940, new_n2941,
    new_n2943, new_n2945, new_n2946, new_n2947, new_n2949, new_n2951,
    new_n2952, new_n2954, new_n2956, new_n2958, new_n2959, new_n2961,
    new_n2962, new_n2965, new_n2966, new_n2967, new_n2969, new_n2970,
    new_n2971, new_n2973, new_n2974, new_n2977, new_n2980, new_n2981,
    new_n2985, new_n2986, new_n2990, new_n2992, new_n2993, new_n2995,
    new_n2996, new_n2997, new_n2998;
  nand g0000 ( new_n386 , pi238 , pi238 );
  nand g0001 ( new_n387 , pi060 , pi060 );
  nand g0002 ( new_n388 , pi200 , pi200 );
  nand     g0003 ( new_n389 , new_n387 , new_n388 );
  nand g0004 ( new_n390 , new_n389 , new_n389 );
  nand g0005 ( new_n391 , pi094 , pi094 );
  nand g0006 ( new_n392 , pi146 , pi146 );
  nand     g0007 ( new_n393 , pi128 , new_n392 );
  nand     g0008 ( new_n394 , new_n391 , new_n393 );
  nand g0009 ( new_n395 , new_n394 , new_n394 );
  nand     g0010 ( new_n396 , new_n390 , new_n395 );
  nand g0011 ( new_n397 , new_n396 , new_n396 );
  nand g0012 ( new_n398 , pi246 , pi246 );
  nand     g0013 ( new_n399 , new_n392 , new_n398 );
  nand g0014 ( new_n400 , new_n399 , new_n399 );
  nand     g0015 ( new_n401 , pi117 , new_n400 );
  nand     g0016 ( new_n402 , new_n397 , new_n401 );
  nand g0017 ( new_n403 , pi171 , pi171 );
  nand     g0018 ( new_n404 , new_n388 , pi226 );
  nand     g0019 ( new_n405 , new_n403 , new_n404 );
  nand g0020 ( new_n406 , new_n405 , new_n405 );
  nand     g0021 ( new_n407 , new_n402 , new_n406 );
  nand g0022 ( new_n408 , pi144 , pi144 );
  nand g0023 ( new_n409 , pi077 , pi077 );
  nand g0024 ( new_n410 , pi090 , pi090 );
  nand     g0025 ( new_n411 , new_n409 , new_n410 );
  nand g0026 ( new_n412 , new_n411 , new_n411 );
  nand     g0027 ( new_n413 , new_n408 , new_n412 );
  nand g0028 ( new_n414 , pi182 , pi182 );
  or       g0029 ( new_n415 , pi103 , pi153 );
  nand g0030 ( new_n416 , pi021 , pi021 );
  nand     g0031 ( new_n417 , new_n416 , new_n387 );
  nor      g0032 ( new_n418 , new_n415 , new_n417 );
  nand     g0033 ( new_n419 , new_n414 , new_n418 );
  nor      g0034 ( new_n420 , new_n413 , new_n419 );
  nand     g0035 ( new_n421 , new_n407 , new_n420 );
  nand g0036 ( new_n422 , new_n421 , new_n421 );
  nor      g0037 ( new_n423 , pi069 , pi098 );
  nand g0038 ( new_n424 , pi223 , pi223 );
  nand g0039 ( new_n425 , pi220 , pi220 );
  or       g0040 ( new_n426 , pi069 , new_n425 );
  nand     g0041 ( new_n427 , new_n424 , new_n426 );
  nor      g0042 ( new_n428 , new_n423 , new_n427 );
  nor      g0043 ( new_n429 , pi120 , new_n428 );
  nand g0044 ( new_n430 , pi156 , pi156 );
  nor      g0045 ( new_n431 , pi049 , pi076 );
  nand     g0046 ( new_n432 , new_n430 , new_n431 );
  nand g0047 ( new_n433 , pi239 , pi239 );
  nand g0048 ( new_n434 , pi010 , pi010 );
  or       g0049 ( new_n435 , new_n434 , pi204 );
  nand     g0050 ( new_n436 , new_n433 , new_n435 );
  nand g0051 ( new_n437 , new_n436 , new_n436 );
  or       g0052 ( new_n438 , new_n432 , new_n437 );
  nand g0053 ( new_n439 , pi237 , pi237 );
  nor      g0054 ( new_n440 , pi049 , new_n439 );
  nor      g0055 ( new_n441 , pi030 , new_n440 );
  nor      g0056 ( new_n442 , pi156 , new_n441 );
  nor      g0057 ( new_n443 , pi159 , pi220 );
  nand     g0058 ( new_n444 , new_n424 , new_n443 );
  nor      g0059 ( new_n445 , new_n442 , new_n444 );
  nand     g0060 ( new_n446 , new_n438 , new_n445 );
  nand     g0061 ( new_n447 , new_n429 , new_n446 );
  nand g0062 ( new_n448 , pi016 , pi016 );
  nand g0063 ( new_n449 , pi056 , pi056 );
  nand     g0064 ( new_n450 , new_n448 , new_n449 );
  nand g0065 ( new_n451 , pi139 , pi139 );
  nand g0066 ( new_n452 , pi232 , pi232 );
  nand     g0067 ( new_n453 , new_n451 , new_n452 );
  or       g0068 ( new_n454 , pi126 , new_n453 );
  nor      g0069 ( new_n455 , new_n450 , new_n454 );
  nand     g0070 ( new_n456 , new_n447 , new_n455 );
  nand g0071 ( new_n457 , pi178 , pi178 );
  nor      g0072 ( new_n458 , new_n457 , new_n453 );
  nand g0073 ( new_n459 , pi012 , pi012 );
  nand     g0074 ( new_n460 , new_n451 , pi207 );
  nand     g0075 ( new_n461 , new_n459 , new_n460 );
  nor      g0076 ( new_n462 , new_n458 , new_n461 );
  nor      g0077 ( new_n463 , new_n450 , new_n462 );
  nand g0078 ( new_n464 , pi082 , pi082 );
  or       g0079 ( new_n465 , pi011 , new_n449 );
  nor      g0080 ( new_n466 , pi011 , pi152 );
  nand g0081 ( new_n467 , new_n466 , new_n466 );
  nand     g0082 ( new_n468 , new_n465 , new_n467 );
  nand     g0083 ( new_n469 , new_n464 , new_n468 );
  nor      g0084 ( new_n470 , new_n463 , new_n469 );
  nand     g0085 ( new_n471 , new_n456 , new_n470 );
  nand g0086 ( new_n472 , pi227 , pi227 );
  nand g0087 ( new_n473 , pi253 , pi253 );
  nand     g0088 ( new_n474 , new_n472 , new_n473 );
  nand g0089 ( new_n475 , new_n474 , new_n474 );
  nand g0090 ( new_n476 , pi255 , pi255 );
  nand     g0091 ( new_n477 , pi252 , new_n476 );
  nand g0092 ( new_n478 , pi125 , pi125 );
  nand g0093 ( new_n479 , pi251 , pi251 );
  nand     g0094 ( new_n480 , new_n478 , new_n479 );
  nand g0095 ( new_n481 , new_n480 , new_n480 );
  nand     g0096 ( new_n482 , new_n477 , new_n481 );
  nor      g0097 ( new_n483 , pi176 , new_n482 );
  nand     g0098 ( new_n484 , new_n475 , new_n483 );
  nand g0099 ( new_n485 , pi007 , pi007 );
  nor      g0100 ( new_n486 , pi025 , pi190 );
  nand g0101 ( new_n487 , new_n486 , new_n486 );
  nand g0102 ( new_n488 , pi165 , pi165 );
  nor      g0103 ( new_n489 , new_n488 , pi190 );
  nand g0104 ( new_n490 , new_n489 , new_n489 );
  nand     g0105 ( new_n491 , new_n487 , new_n490 );
  nand     g0106 ( new_n492 , new_n485 , new_n491 );
  nand g0107 ( new_n493 , new_n492 , new_n492 );
  nand g0108 ( new_n494 , pi155 , pi155 );
  nor      g0109 ( new_n495 , pi047 , pi141 );
  nand     g0110 ( new_n496 , new_n494 , new_n495 );
  nand     g0111 ( new_n497 , pi198 , new_n495 );
  nand     g0112 ( new_n498 , new_n496 , new_n497 );
  nand     g0113 ( new_n499 , new_n493 , new_n498 );
  nand g0114 ( new_n500 , pi143 , pi143 );
  nand     g0115 ( new_n501 , new_n500 , new_n488 );
  nand     g0116 ( new_n502 , new_n493 , new_n501 );
  nand g0117 ( new_n503 , new_n502 , new_n502 );
  nand g0118 ( new_n504 , pi066 , pi066 );
  nand     g0119 ( new_n505 , new_n485 , pi199 );
  nand     g0120 ( new_n506 , new_n504 , new_n505 );
  nor      g0121 ( new_n507 , new_n503 , new_n506 );
  nand g0122 ( new_n508 , new_n507 , new_n507 );
  nand g0123 ( new_n509 , pi092 , pi092 );
  nor      g0124 ( new_n510 , new_n509 , pi141 );
  nand     g0125 ( new_n511 , new_n493 , new_n510 );
  nor      g0126 ( new_n512 , pi041 , pi215 );
  nand g0127 ( new_n513 , pi050 , pi050 );
  nand g0128 ( new_n514 , pi079 , pi079 );
  nand     g0129 ( new_n515 , new_n513 , new_n514 );
  nand g0130 ( new_n516 , new_n515 , new_n515 );
  nand     g0131 ( new_n517 , new_n512 , new_n516 );
  nand g0132 ( new_n518 , new_n517 , new_n517 );
  nand     g0133 ( new_n519 , new_n511 , new_n518 );
  nor      g0134 ( new_n520 , new_n508 , new_n519 );
  nand     g0135 ( new_n521 , new_n499 , new_n520 );
  or       g0136 ( new_n522 , new_n484 , new_n521 );
  nand g0137 ( new_n523 , pi067 , pi067 );
  nand     g0138 ( new_n524 , new_n523 , pi079 );
  nand g0139 ( new_n525 , pi109 , pi109 );
  nand     g0140 ( new_n526 , new_n523 , new_n525 );
  nand     g0141 ( new_n527 , new_n524 , new_n526 );
  nand     g0142 ( new_n528 , new_n476 , new_n527 );
  nand g0143 ( new_n529 , new_n512 , new_n512 );
  nand g0144 ( new_n530 , pi228 , pi228 );
  nor      g0145 ( new_n531 , pi215 , new_n530 );
  nor      g0146 ( new_n532 , pi105 , new_n531 );
  nand     g0147 ( new_n533 , new_n529 , new_n532 );
  nand     g0148 ( new_n534 , new_n516 , new_n533 );
  nand g0149 ( new_n535 , pi183 , pi183 );
  nand     g0150 ( new_n536 , new_n535 , new_n530 );
  or       g0151 ( new_n537 , pi105 , new_n536 );
  nand g0152 ( new_n538 , new_n537 , new_n537 );
  nor      g0153 ( new_n539 , new_n534 , new_n538 );
  nor      g0154 ( new_n540 , new_n528 , new_n539 );
  nor      g0155 ( new_n541 , new_n484 , new_n540 );
  nand     g0156 ( new_n542 , new_n430 , new_n423 );
  nand g0157 ( new_n543 , new_n542 , new_n542 );
  nand     g0158 ( new_n544 , new_n431 , new_n543 );
  nor      g0159 ( new_n545 , pi120 , new_n544 );
  nand g0160 ( new_n546 , new_n545 , new_n545 );
  nor      g0161 ( new_n547 , pi138 , pi210 );
  nand g0162 ( new_n548 , new_n547 , new_n547 );
  nor      g0163 ( new_n549 , pi242 , new_n548 );
  nand g0164 ( new_n550 , new_n549 , new_n549 );
  nand     g0165 ( new_n551 , pi125 , new_n547 );
  nand g0166 ( new_n552 , new_n551 , new_n551 );
  nand g0167 ( new_n553 , pi176 , pi176 );
  nor      g0168 ( new_n554 , pi138 , new_n553 );
  nand g0169 ( new_n555 , new_n554 , new_n554 );
  nand     g0170 ( new_n556 , new_n475 , new_n555 );
  nor      g0171 ( new_n557 , new_n552 , new_n556 );
  nand     g0172 ( new_n558 , new_n550 , new_n557 );
  nand g0173 ( new_n559 , pi115 , pi115 );
  nand     g0174 ( new_n560 , pi214 , new_n472 );
  nand     g0175 ( new_n561 , new_n559 , new_n560 );
  nor      g0176 ( new_n562 , pi204 , new_n561 );
  nand     g0177 ( new_n563 , new_n558 , new_n562 );
  nor      g0178 ( new_n564 , new_n546 , new_n563 );
  nand     g0179 ( new_n565 , new_n470 , new_n564 );
  nor      g0180 ( new_n566 , new_n541 , new_n565 );
  nand     g0181 ( new_n567 , new_n522 , new_n566 );
  nand g0182 ( new_n568 , new_n567 , new_n567 );
  nand g0183 ( new_n569 , pi219 , pi219 );
  nand g0184 ( new_n570 , pi163 , pi163 );
  nand g0185 ( new_n571 , pi248 , pi248 );
  nand     g0186 ( new_n572 , new_n570 , new_n571 );
  nand g0187 ( new_n573 , new_n572 , new_n572 );
  nand     g0188 ( new_n574 , new_n569 , new_n573 );
  nand g0189 ( new_n575 , pi136 , pi136 );
  nand g0190 ( new_n576 , pi166 , pi166 );
  nand g0191 ( new_n577 , pi187 , pi187 );
  or       g0192 ( new_n578 , pi123 , new_n577 );
  nand     g0193 ( new_n579 , new_n576 , new_n578 );
  nand g0194 ( new_n580 , new_n579 , new_n579 );
  nand g0195 ( new_n581 , pi129 , pi129 );
  nand g0196 ( new_n582 , pi189 , pi189 );
  nand     g0197 ( new_n583 , new_n581 , new_n582 );
  nand g0198 ( new_n584 , new_n583 , new_n583 );
  nor      g0199 ( new_n585 , pi057 , pi123 );
  nand     g0200 ( new_n586 , new_n581 , pi194 );
  nand     g0201 ( new_n587 , new_n585 , new_n586 );
  nor      g0202 ( new_n588 , new_n584 , new_n587 );
  nand g0203 ( new_n589 , new_n588 , new_n588 );
  nand     g0204 ( new_n590 , new_n580 , new_n589 );
  nand g0205 ( new_n591 , new_n590 , new_n590 );
  nand     g0206 ( new_n592 , new_n575 , new_n591 );
  nand g0207 ( new_n593 , new_n592 , new_n592 );
  nand g0208 ( new_n594 , pi164 , pi164 );
  nand g0209 ( new_n595 , pi194 , pi194 );
  nand     g0210 ( new_n596 , new_n594 , new_n595 );
  nand g0211 ( new_n597 , new_n596 , new_n596 );
  nand     g0212 ( new_n598 , new_n585 , new_n597 );
  nand g0213 ( new_n599 , new_n598 , new_n598 );
  nor      g0214 ( new_n600 , pi111 , pi224 );
  nand g0215 ( new_n601 , pi108 , pi108 );
  nand g0216 ( new_n602 , pi185 , pi185 );
  nor      g0217 ( new_n603 , pi111 , new_n602 );
  nand g0218 ( new_n604 , new_n603 , new_n603 );
  nand     g0219 ( new_n605 , new_n601 , new_n604 );
  or       g0220 ( new_n606 , new_n600 , new_n605 );
  nand     g0221 ( new_n607 , new_n599 , new_n606 );
  nand     g0222 ( new_n608 , new_n593 , new_n607 );
  nor      g0223 ( new_n609 , new_n574 , new_n608 );
  nand g0224 ( new_n610 , pi089 , pi089 );
  nor      g0225 ( new_n611 , pi042 , pi102 );
  nand g0226 ( new_n612 , new_n611 , new_n611 );
  nor      g0227 ( new_n613 , pi042 , new_n575 );
  nand g0228 ( new_n614 , new_n613 , new_n613 );
  nand     g0229 ( new_n615 , new_n612 , new_n614 );
  nand     g0230 ( new_n616 , new_n610 , new_n615 );
  nand g0231 ( new_n617 , new_n616 , new_n616 );
  nand     g0232 ( new_n618 , new_n610 , pi219 );
  nand     g0233 ( new_n619 , new_n573 , new_n618 );
  nor      g0234 ( new_n620 , new_n617 , new_n619 );
  nand g0235 ( new_n621 , pi169 , pi169 );
  nand g0236 ( new_n622 , pi118 , pi118 );
  or       g0237 ( new_n623 , new_n622 , pi192 );
  nor      g0238 ( new_n624 , pi192 , pi217 );
  nand g0239 ( new_n625 , new_n624 , new_n624 );
  nand     g0240 ( new_n626 , new_n623 , new_n625 );
  nand     g0241 ( new_n627 , new_n621 , new_n626 );
  nand g0242 ( new_n628 , new_n627 , new_n627 );
  nand g0243 ( new_n629 , pi100 , pi100 );
  nor      g0244 ( new_n630 , pi017 , pi167 );
  nor      g0245 ( new_n631 , pi068 , pi113 );
  nand     g0246 ( new_n632 , new_n630 , new_n631 );
  nand g0247 ( new_n633 , new_n632 , new_n632 );
  nand     g0248 ( new_n634 , new_n629 , new_n633 );
  nand g0249 ( new_n635 , new_n634 , new_n634 );
  nand     g0250 ( new_n636 , pi026 , new_n571 );
  nand     g0251 ( new_n637 , new_n635 , new_n636 );
  nand g0252 ( new_n638 , new_n637 , new_n637 );
  nand     g0253 ( new_n639 , new_n628 , new_n638 );
  nor      g0254 ( new_n640 , new_n620 , new_n639 );
  nand g0255 ( new_n641 , new_n640 , new_n640 );
  nor      g0256 ( new_n642 , new_n609 , new_n641 );
  nand g0257 ( new_n643 , pi221 , pi221 );
  nand g0258 ( new_n644 , pi062 , pi062 );
  nand g0259 ( new_n645 , pi071 , pi071 );
  nand g0260 ( new_n646 , pi172 , pi172 );
  nand     g0261 ( new_n647 , new_n646 , pi181 );
  nand     g0262 ( new_n648 , new_n645 , new_n647 );
  nand     g0263 ( new_n649 , new_n644 , new_n648 );
  nand     g0264 ( new_n650 , new_n643 , new_n649 );
  nand     g0265 ( new_n651 , new_n644 , new_n646 );
  nor      g0266 ( new_n652 , pi247 , new_n651 );
  nand g0267 ( new_n653 , new_n652 , new_n652 );
  nand g0268 ( new_n654 , pi196 , pi196 );
  nand     g0269 ( new_n655 , pi078 , new_n654 );
  nand g0270 ( new_n656 , pi201 , pi201 );
  nand     g0271 ( new_n657 , new_n654 , new_n656 );
  nand     g0272 ( new_n658 , new_n655 , new_n657 );
  nor      g0273 ( new_n659 , new_n653 , new_n658 );
  nand     g0274 ( new_n660 , new_n601 , new_n602 );
  nand g0275 ( new_n661 , new_n660 , new_n660 );
  nand     g0276 ( new_n662 , new_n576 , new_n577 );
  nor      g0277 ( new_n663 , new_n583 , new_n662 );
  nand     g0278 ( new_n664 , new_n661 , new_n663 );
  nand g0279 ( new_n665 , new_n664 , new_n664 );
  nand     g0280 ( new_n666 , new_n575 , new_n665 );
  or       g0281 ( new_n667 , new_n659 , new_n666 );
  or       g0282 ( new_n668 , new_n650 , new_n667 );
  nand g0283 ( new_n669 , new_n574 , new_n574 );
  nand     g0284 ( new_n670 , new_n600 , new_n652 );
  nand g0285 ( new_n671 , new_n670 , new_n670 );
  nand     g0286 ( new_n672 , new_n599 , new_n671 );
  nand g0287 ( new_n673 , new_n672 , new_n672 );
  nand g0288 ( new_n674 , pi039 , pi039 );
  nor      g0289 ( new_n675 , pi078 , pi195 );
  nand     g0290 ( new_n676 , new_n674 , new_n675 );
  nand     g0291 ( new_n677 , pi104 , new_n675 );
  nand     g0292 ( new_n678 , new_n676 , new_n677 );
  nand     g0293 ( new_n679 , new_n673 , new_n678 );
  nand     g0294 ( new_n680 , new_n669 , new_n679 );
  nor      g0295 ( new_n681 , new_n668 , new_n680 );
  nand g0296 ( new_n682 , pi013 , pi013 );
  nand g0297 ( new_n683 , pi168 , pi168 );
  nand     g0298 ( new_n684 , new_n682 , new_n683 );
  nor      g0299 ( new_n685 , pi070 , new_n684 );
  nand g0300 ( new_n686 , new_n685 , new_n685 );
  nand g0301 ( new_n687 , pi051 , pi051 );
  nand     g0302 ( new_n688 , new_n682 , pi074 );
  nand     g0303 ( new_n689 , new_n687 , new_n688 );
  nand     g0304 ( new_n690 , new_n683 , new_n689 );
  nand g0305 ( new_n691 , new_n690 , new_n690 );
  nand g0306 ( new_n692 , pi114 , pi114 );
  nand g0307 ( new_n693 , pi179 , pi179 );
  nand     g0308 ( new_n694 , new_n692 , new_n693 );
  nor      g0309 ( new_n695 , new_n691 , new_n694 );
  nand     g0310 ( new_n696 , new_n686 , new_n695 );
  nand g0311 ( new_n697 , pi147 , pi147 );
  nand     g0312 ( new_n698 , pi009 , new_n697 );
  or       g0313 ( new_n699 , pi051 , pi074 );
  nand g0314 ( new_n700 , pi240 , pi240 );
  nand     g0315 ( new_n701 , new_n693 , new_n700 );
  nor      g0316 ( new_n702 , new_n699 , new_n701 );
  nand     g0317 ( new_n703 , new_n692 , new_n702 );
  nand g0318 ( new_n704 , new_n703 , new_n703 );
  nand     g0319 ( new_n705 , new_n698 , new_n704 );
  nand     g0320 ( new_n706 , new_n696 , new_n705 );
  nand g0321 ( new_n707 , new_n706 , new_n706 );
  nor      g0322 ( new_n708 , new_n681 , new_n707 );
  nand     g0323 ( new_n709 , new_n642 , new_n708 );
  nand g0324 ( new_n710 , pi154 , pi154 );
  nand     g0325 ( new_n711 , pi055 , new_n710 );
  nand g0326 ( new_n712 , new_n711 , new_n711 );
  or       g0327 ( new_n713 , pi035 , pi132 );
  nor      g0328 ( new_n714 , new_n712 , new_n713 );
  nand g0329 ( new_n715 , pi083 , pi083 );
  nand g0330 ( new_n716 , pi145 , pi145 );
  nand     g0331 ( new_n717 , new_n715 , new_n716 );
  nor      g0332 ( new_n718 , pi243 , new_n717 );
  nor      g0333 ( new_n719 , pi059 , pi208 );
  nand     g0334 ( new_n720 , new_n718 , new_n719 );
  nand g0335 ( new_n721 , pi001 , pi001 );
  nand g0336 ( new_n722 , pi151 , pi151 );
  nand     g0337 ( new_n723 , new_n721 , new_n722 );
  nand g0338 ( new_n724 , new_n723 , new_n723 );
  nor      g0339 ( new_n725 , pi061 , pi173 );
  nand     g0340 ( new_n726 , new_n724 , new_n725 );
  nor      g0341 ( new_n727 , new_n720 , new_n726 );
  nand     g0342 ( new_n728 , new_n714 , new_n727 );
  nand g0343 ( new_n729 , new_n728 , new_n728 );
  nand g0344 ( new_n730 , pi188 , pi188 );
  nand     g0345 ( new_n731 , pi084 , new_n730 );
  nand g0346 ( new_n732 , new_n731 , new_n731 );
  nand g0347 ( new_n733 , pi048 , pi048 );
  nand g0348 ( new_n734 , pi052 , pi052 );
  nand     g0349 ( new_n735 , new_n733 , new_n734 );
  nor      g0350 ( new_n736 , new_n732 , new_n735 );
  nand g0351 ( new_n737 , pi015 , pi015 );
  nand     g0352 ( new_n738 , new_n734 , pi235 );
  nand     g0353 ( new_n739 , new_n737 , new_n738 );
  nor      g0354 ( new_n740 , new_n736 , new_n739 );
  nor      g0355 ( new_n741 , pi148 , new_n740 );
  nor      g0356 ( new_n742 , pi086 , new_n741 );
  nand g0357 ( new_n743 , pi091 , pi091 );
  nand g0358 ( new_n744 , pi142 , pi142 );
  nand     g0359 ( new_n745 , new_n743 , new_n744 );
  nor      g0360 ( new_n746 , new_n742 , new_n745 );
  nand g0361 ( new_n747 , pi216 , pi216 );
  nor      g0362 ( new_n748 , pi045 , pi058 );
  nand     g0363 ( new_n749 , new_n747 , new_n748 );
  nand g0364 ( new_n750 , new_n748 , new_n748 );
  nand g0365 ( new_n751 , pi058 , pi058 );
  nand     g0366 ( new_n752 , new_n751 , pi064 );
  and      g0367 ( new_n753 , new_n750 , new_n752 );
  nor      g0368 ( new_n754 , pi064 , pi191 );
  nor      g0369 ( new_n755 , new_n753 , new_n754 );
  nand g0370 ( new_n756 , pi046 , pi046 );
  nand g0371 ( new_n757 , pi112 , pi112 );
  nand     g0372 ( new_n758 , new_n756 , new_n757 );
  nor      g0373 ( new_n759 , new_n755 , new_n758 );
  nand     g0374 ( new_n760 , new_n749 , new_n759 );
  nand g0375 ( new_n761 , pi222 , pi222 );
  nand     g0376 ( new_n762 , new_n761 , new_n754 );
  nand g0377 ( new_n763 , new_n762 , new_n762 );
  nand g0378 ( new_n764 , pi004 , pi004 );
  nand     g0379 ( new_n765 , new_n764 , pi150 );
  nand g0380 ( new_n766 , new_n765 , new_n765 );
  nor      g0381 ( new_n767 , new_n758 , new_n766 );
  nand     g0382 ( new_n768 , new_n763 , new_n767 );
  nand     g0383 ( new_n769 , new_n760 , new_n768 );
  nand g0384 ( new_n770 , pi133 , pi133 );
  nand g0385 ( new_n771 , pi175 , pi175 );
  nand     g0386 ( new_n772 , new_n770 , new_n771 );
  nand g0387 ( new_n773 , new_n772 , new_n772 );
  nand g0388 ( new_n774 , pi053 , pi053 );
  nand     g0389 ( new_n775 , new_n774 , pi184 );
  nand     g0390 ( new_n776 , new_n773 , new_n775 );
  nand g0391 ( new_n777 , pi110 , pi110 );
  nand g0392 ( new_n778 , pi093 , pi093 );
  nand     g0393 ( new_n779 , new_n778 , pi244 );
  nand     g0394 ( new_n780 , new_n777 , new_n779 );
  nor      g0395 ( new_n781 , pi053 , new_n780 );
  nor      g0396 ( new_n782 , new_n776 , new_n781 );
  nand g0397 ( new_n783 , pi229 , pi229 );
  nand     g0398 ( new_n784 , pi124 , new_n770 );
  nand     g0399 ( new_n785 , new_n783 , new_n784 );
  nor      g0400 ( new_n786 , pi008 , new_n785 );
  nand g0401 ( new_n787 , new_n786 , new_n786 );
  nor      g0402 ( new_n788 , new_n782 , new_n787 );
  and      g0403 ( new_n789 , new_n769 , new_n788 );
  nand     g0404 ( new_n790 , new_n746 , new_n789 );
  nor      g0405 ( new_n791 , pi160 , pi209 );
  nand g0406 ( new_n792 , new_n791 , new_n791 );
  nand g0407 ( new_n793 , pi008 , pi008 );
  or       g0408 ( new_n794 , new_n793 , pi160 );
  nand     g0409 ( new_n795 , new_n792 , new_n794 );
  nand     g0410 ( new_n796 , new_n764 , new_n795 );
  or       g0411 ( new_n797 , new_n749 , new_n796 );
  nand     g0412 ( new_n798 , new_n769 , new_n797 );
  nand g0413 ( new_n799 , new_n798 , new_n798 );
  or       g0414 ( new_n800 , new_n789 , new_n799 );
  nor      g0415 ( new_n801 , new_n776 , new_n797 );
  or       g0416 ( new_n802 , pi031 , pi093 );
  nand g0417 ( new_n803 , pi249 , pi249 );
  nor      g0418 ( new_n804 , pi091 , new_n803 );
  nor      g0419 ( new_n805 , new_n802 , new_n804 );
  nand     g0420 ( new_n806 , new_n801 , new_n805 );
  nand     g0421 ( new_n807 , new_n800 , new_n806 );
  nand     g0422 ( new_n808 , new_n790 , new_n807 );
  nand     g0423 ( new_n809 , new_n729 , new_n808 );
  nor      g0424 ( new_n810 , pi135 , pi203 );
  nor      g0425 ( new_n811 , pi087 , pi177 );
  nand g0426 ( new_n812 , new_n811 , new_n811 );
  nand g0427 ( new_n813 , pi059 , pi059 );
  nor      g0428 ( new_n814 , new_n813 , pi177 );
  nor      g0429 ( new_n815 , pi208 , new_n814 );
  nand     g0430 ( new_n816 , new_n812 , new_n815 );
  nand     g0431 ( new_n817 , new_n810 , new_n816 );
  nand g0432 ( new_n818 , pi173 , pi173 );
  nand g0433 ( new_n819 , pi061 , pi061 );
  nor      g0434 ( new_n820 , new_n819 , pi203 );
  nand g0435 ( new_n821 , new_n820 , new_n820 );
  nand     g0436 ( new_n822 , new_n818 , new_n821 );
  nand g0437 ( new_n823 , new_n822 , new_n822 );
  nand     g0438 ( new_n824 , new_n817 , new_n823 );
  nand g0439 ( new_n825 , pi211 , pi211 );
  nand g0440 ( new_n826 , pi225 , pi225 );
  nand     g0441 ( new_n827 , new_n825 , new_n826 );
  nand g0442 ( new_n828 , new_n827 , new_n827 );
  nand     g0443 ( new_n829 , new_n824 , new_n828 );
  or       g0444 ( new_n830 , pi024 , pi040 );
  nor      g0445 ( new_n831 , pi024 , new_n716 );
  nor      g0446 ( new_n832 , pi243 , new_n831 );
  nand     g0447 ( new_n833 , new_n830 , new_n832 );
  nand     g0448 ( new_n834 , new_n811 , new_n833 );
  nor      g0449 ( new_n835 , new_n718 , new_n834 );
  nand     g0450 ( new_n836 , new_n819 , new_n815 );
  nor      g0451 ( new_n837 , new_n835 , new_n836 );
  nand     g0452 ( new_n838 , new_n818 , new_n837 );
  nand g0453 ( new_n839 , pi014 , pi014 );
  nand     g0454 ( new_n840 , pi001 , new_n839 );
  nand g0455 ( new_n841 , new_n840 , new_n840 );
  nand g0456 ( new_n842 , pi140 , pi140 );
  nand     g0457 ( new_n843 , new_n839 , new_n842 );
  nand g0458 ( new_n844 , pi250 , pi250 );
  nor      g0459 ( new_n845 , pi132 , new_n844 );
  nor      g0460 ( new_n846 , pi134 , new_n845 );
  nor      g0461 ( new_n847 , pi151 , new_n846 );
  nor      g0462 ( new_n848 , new_n843 , new_n847 );
  nor      g0463 ( new_n849 , new_n841 , new_n848 );
  nor      g0464 ( new_n850 , new_n830 , new_n849 );
  nor      g0465 ( new_n851 , new_n838 , new_n850 );
  nor      g0466 ( new_n852 , new_n829 , new_n851 );
  nand     g0467 ( new_n853 , new_n728 , new_n852 );
  nor      g0468 ( new_n854 , new_n676 , new_n853 );
  nand g0469 ( new_n855 , new_n676 , new_n676 );
  nand     g0470 ( new_n856 , new_n855 , new_n828 );
  nor      g0471 ( new_n857 , new_n812 , new_n830 );
  nand g0472 ( new_n858 , new_n857 , new_n857 );
  nand g0473 ( new_n859 , pi134 , pi134 );
  nand     g0474 ( new_n860 , new_n859 , new_n844 );
  or       g0475 ( new_n861 , new_n843 , new_n860 );
  nor      g0476 ( new_n862 , new_n858 , new_n861 );
  nand g0477 ( new_n863 , new_n862 , new_n862 );
  nand g0478 ( new_n864 , pi197 , pi197 );
  nand     g0479 ( new_n865 , pi006 , new_n757 );
  nand     g0480 ( new_n866 , new_n864 , new_n865 );
  nor      g0481 ( new_n867 , pi154 , new_n866 );
  nand     g0482 ( new_n868 , new_n810 , new_n867 );
  nor      g0483 ( new_n869 , new_n863 , new_n868 );
  nand g0484 ( new_n870 , new_n869 , new_n869 );
  nor      g0485 ( new_n871 , new_n856 , new_n870 );
  nor      g0486 ( new_n872 , new_n854 , new_n871 );
  nand     g0487 ( new_n873 , new_n594 , new_n671 );
  nor      g0488 ( new_n874 , new_n872 , new_n873 );
  nand     g0489 ( new_n875 , new_n809 , new_n874 );
  nand g0490 ( new_n876 , new_n605 , new_n605 );
  nand     g0491 ( new_n877 , new_n600 , new_n650 );
  nand     g0492 ( new_n878 , new_n876 , new_n877 );
  nand g0493 ( new_n879 , new_n878 , new_n878 );
  nand     g0494 ( new_n880 , new_n670 , new_n879 );
  nand     g0495 ( new_n881 , new_n594 , new_n880 );
  nand     g0496 ( new_n882 , new_n584 , new_n881 );
  nand     g0497 ( new_n883 , new_n658 , new_n677 );
  nand g0498 ( new_n884 , pi054 , pi054 );
  nand     g0499 ( new_n885 , new_n884 , pi211 );
  nand     g0500 ( new_n886 , new_n855 , new_n885 );
  nand g0501 ( new_n887 , new_n886 , new_n886 );
  nor      g0502 ( new_n888 , new_n883 , new_n887 );
  nand g0503 ( new_n889 , new_n888 , new_n888 );
  nand g0504 ( new_n890 , new_n657 , new_n657 );
  nand g0505 ( new_n891 , pi104 , pi104 );
  nand g0506 ( new_n892 , pi158 , pi158 );
  nand     g0507 ( new_n893 , new_n884 , new_n892 );
  nand g0508 ( new_n894 , new_n893 , new_n893 );
  nand     g0509 ( new_n895 , new_n891 , new_n894 );
  nand g0510 ( new_n896 , new_n895 , new_n895 );
  nand     g0511 ( new_n897 , new_n890 , new_n896 );
  nand     g0512 ( new_n898 , new_n889 , new_n897 );
  nand     g0513 ( new_n899 , pi221 , new_n600 );
  nand     g0514 ( new_n900 , new_n876 , new_n899 );
  nand g0515 ( new_n901 , pi181 , pi181 );
  nand     g0516 ( new_n902 , new_n645 , new_n901 );
  nand g0517 ( new_n903 , new_n902 , new_n902 );
  nand     g0518 ( new_n904 , new_n584 , new_n903 );
  nor      g0519 ( new_n905 , new_n900 , new_n904 );
  nand     g0520 ( new_n906 , new_n898 , new_n905 );
  nand     g0521 ( new_n907 , new_n882 , new_n906 );
  nand     g0522 ( new_n908 , new_n875 , new_n907 );
  nand g0523 ( new_n909 , new_n788 , new_n788 );
  nand g0524 ( new_n910 , new_n802 , new_n802 );
  nand     g0525 ( new_n911 , pi142 , new_n803 );
  nand     g0526 ( new_n912 , new_n743 , new_n911 );
  nand g0527 ( new_n913 , new_n912 , new_n912 );
  nor      g0528 ( new_n914 , pi086 , pi249 );
  nand     g0529 ( new_n915 , pi148 , new_n914 );
  nand     g0530 ( new_n916 , new_n913 , new_n915 );
  nand     g0531 ( new_n917 , new_n910 , new_n916 );
  nand g0532 ( new_n918 , new_n917 , new_n917 );
  nand     g0533 ( new_n919 , new_n737 , new_n914 );
  nand     g0534 ( new_n920 , new_n738 , new_n910 );
  nor      g0535 ( new_n921 , new_n919 , new_n920 );
  or       g0536 ( new_n922 , new_n918 , new_n921 );
  nand g0537 ( new_n923 , new_n922 , new_n922 );
  nor      g0538 ( new_n924 , new_n776 , new_n923 );
  nor      g0539 ( new_n925 , new_n909 , new_n924 );
  nor      g0540 ( new_n926 , new_n796 , new_n925 );
  nand     g0541 ( new_n927 , new_n760 , new_n869 );
  nor      g0542 ( new_n928 , new_n829 , new_n927 );
  nand     g0543 ( new_n929 , new_n926 , new_n928 );
  nand g0544 ( new_n930 , pi193 , pi193 );
  nor      g0545 ( new_n931 , pi096 , pi162 );
  nand g0546 ( new_n932 , pi002 , pi002 );
  nand g0547 ( new_n933 , pi095 , pi095 );
  nand     g0548 ( new_n934 , pi034 , new_n933 );
  nand     g0549 ( new_n935 , new_n932 , new_n934 );
  nand     g0550 ( new_n936 , new_n931 , new_n935 );
  nand g0551 ( new_n937 , pi044 , pi044 );
  nor      g0552 ( new_n938 , new_n937 , pi162 );
  nor      g0553 ( new_n939 , pi205 , new_n938 );
  nand     g0554 ( new_n940 , new_n936 , new_n939 );
  nand     g0555 ( new_n941 , new_n930 , new_n940 );
  nor      g0556 ( new_n942 , pi084 , pi116 );
  nand     g0557 ( new_n943 , new_n941 , new_n942 );
  nand g0558 ( new_n944 , pi245 , pi245 );
  nand     g0559 ( new_n945 , pi023 , new_n944 );
  nor      g0560 ( new_n946 , pi095 , pi101 );
  nand     g0561 ( new_n947 , new_n945 , new_n946 );
  nand     g0562 ( new_n948 , new_n930 , new_n931 );
  nor      g0563 ( new_n949 , new_n947 , new_n948 );
  nor      g0564 ( new_n950 , new_n943 , new_n949 );
  nand g0565 ( new_n951 , pi130 , pi130 );
  nor      g0566 ( new_n952 , pi084 , new_n951 );
  nand g0567 ( new_n953 , pi235 , pi235 );
  nand     g0568 ( new_n954 , new_n730 , new_n953 );
  nor      g0569 ( new_n955 , new_n952 , new_n954 );
  nand g0570 ( new_n956 , new_n955 , new_n955 );
  nor      g0571 ( new_n957 , new_n950 , new_n956 );
  nand g0572 ( new_n958 , new_n957 , new_n957 );
  or       g0573 ( new_n959 , new_n929 , new_n958 );
  nand     g0574 ( new_n960 , new_n575 , new_n669 );
  nand g0575 ( new_n961 , new_n960 , new_n960 );
  nand     g0576 ( new_n962 , new_n580 , new_n961 );
  nand g0577 ( new_n963 , new_n962 , new_n962 );
  nand     g0578 ( new_n964 , new_n959 , new_n963 );
  nor      g0579 ( new_n965 , new_n908 , new_n964 );
  nor      g0580 ( new_n966 , new_n709 , new_n965 );
  nand g0581 ( new_n967 , pi174 , pi174 );
  nand g0582 ( new_n968 , pi180 , pi180 );
  nor      g0583 ( new_n969 , pi068 , new_n968 );
  nand g0584 ( new_n970 , new_n969 , new_n969 );
  nand     g0585 ( new_n971 , new_n967 , new_n970 );
  nand     g0586 ( new_n972 , new_n630 , new_n971 );
  nand g0587 ( new_n973 , pi005 , pi005 );
  nor      g0588 ( new_n974 , new_n973 , pi167 );
  or       g0589 ( new_n975 , pi107 , new_n974 );
  nand g0590 ( new_n976 , new_n975 , new_n975 );
  nand     g0591 ( new_n977 , new_n972 , new_n976 );
  nand g0592 ( new_n978 , new_n977 , new_n977 );
  nand     g0593 ( new_n979 , pi063 , new_n633 );
  nand     g0594 ( new_n980 , new_n978 , new_n979 );
  nor      g0595 ( new_n981 , pi118 , new_n980 );
  nand g0596 ( new_n982 , new_n981 , new_n981 );
  nand     g0597 ( new_n983 , new_n628 , new_n982 );
  nand     g0598 ( new_n984 , pi019 , new_n621 );
  nand g0599 ( new_n985 , new_n984 , new_n984 );
  nand g0600 ( new_n986 , pi037 , pi037 );
  nand     g0601 ( new_n987 , new_n986 , new_n697 );
  nor      g0602 ( new_n988 , new_n985 , new_n987 );
  nand     g0603 ( new_n989 , new_n685 , new_n988 );
  nand g0604 ( new_n990 , new_n989 , new_n989 );
  nand     g0605 ( new_n991 , new_n983 , new_n990 );
  nand     g0606 ( new_n992 , new_n706 , new_n991 );
  nand g0607 ( new_n993 , new_n484 , new_n484 );
  nand g0608 ( new_n994 , pi043 , pi043 );
  nand g0609 ( new_n995 , pi198 , pi198 );
  nand     g0610 ( new_n996 , new_n509 , new_n995 );
  nand g0611 ( new_n997 , new_n996 , new_n996 );
  nand     g0612 ( new_n998 , new_n994 , new_n997 );
  nand g0613 ( new_n999 , new_n501 , new_n501 );
  nor      g0614 ( new_n1000 , pi066 , pi199 );
  nand     g0615 ( new_n1001 , new_n999 , new_n1000 );
  nor      g0616 ( new_n1002 , new_n998 , new_n1001 );
  nand g0617 ( new_n1003 , new_n1002 , new_n1002 );
  nand     g0618 ( new_n1004 , pi106 , new_n692 );
  nand     g0619 ( new_n1005 , new_n518 , new_n1004 );
  nor      g0620 ( new_n1006 , new_n1003 , new_n1005 );
  and      g0621 ( new_n1007 , new_n993 , new_n1006 );
  nand     g0622 ( new_n1008 , new_n992 , new_n1007 );
  or       g0623 ( new_n1009 , new_n966 , new_n1008 );
  nand     g0624 ( new_n1010 , new_n568 , new_n1009 );
  nand     g0625 ( new_n1011 , new_n471 , new_n1010 );
  nand     g0626 ( new_n1012 , new_n422 , new_n1011 );
  nor      g0627 ( new_n1013 , pi184 , new_n802 );
  nand g0628 ( new_n1014 , new_n1013 , new_n1013 );
  nand     g0629 ( new_n1015 , new_n771 , new_n914 );
  nor      g0630 ( new_n1016 , new_n1014 , new_n1015 );
  nand g0631 ( new_n1017 , new_n1016 , new_n1016 );
  nand     g0632 ( new_n1018 , new_n931 , new_n946 );
  nand g0633 ( new_n1019 , new_n1018 , new_n1018 );
  nor      g0634 ( new_n1020 , new_n940 , new_n1019 );
  nand g0635 ( new_n1021 , pi034 , pi034 );
  nand     g0636 ( new_n1022 , new_n932 , new_n1021 );
  nand g0637 ( new_n1023 , pi205 , pi205 );
  nand     g0638 ( new_n1024 , new_n937 , new_n1023 );
  or       g0639 ( new_n1025 , pi245 , new_n1024 );
  nor      g0640 ( new_n1026 , new_n1022 , new_n1025 );
  nor      g0641 ( new_n1027 , new_n1020 , new_n1026 );
  or       g0642 ( new_n1028 , pi116 , new_n1027 );
  nor      g0643 ( new_n1029 , pi085 , pi170 );
  nand g0644 ( new_n1030 , pi233 , pi233 );
  nand     g0645 ( new_n1031 , pi119 , new_n1030 );
  nor      g0646 ( new_n1032 , pi157 , pi233 );
  nor      g0647 ( new_n1033 , pi202 , new_n1032 );
  nand     g0648 ( new_n1034 , new_n1031 , new_n1033 );
  and      g0649 ( new_n1035 , new_n1029 , new_n1034 );
  nand g0650 ( new_n1036 , pi023 , pi023 );
  nand g0651 ( new_n1037 , pi170 , pi170 );
  nand     g0652 ( new_n1038 , pi137 , new_n1037 );
  nand     g0653 ( new_n1039 , new_n1036 , new_n1038 );
  nor      g0654 ( new_n1040 , new_n1035 , new_n1039 );
  nand g0655 ( new_n1041 , pi119 , pi119 );
  nand g0656 ( new_n1042 , pi234 , pi234 );
  nand     g0657 ( new_n1043 , new_n1041 , new_n1042 );
  nor      g0658 ( new_n1044 , pi137 , pi202 );
  nand     g0659 ( new_n1045 , new_n1036 , new_n1044 );
  nor      g0660 ( new_n1046 , new_n1043 , new_n1045 );
  nand g0661 ( new_n1047 , new_n1046 , new_n1046 );
  nand     g0662 ( new_n1048 , new_n944 , new_n1047 );
  nor      g0663 ( new_n1049 , new_n1040 , new_n1048 );
  nor      g0664 ( new_n1050 , new_n1018 , new_n1049 );
  nor      g0665 ( new_n1051 , new_n1028 , new_n1050 );
  nor      g0666 ( new_n1052 , pi000 , pi231 );
  nand g0667 ( new_n1053 , pi161 , pi161 );
  nor      g0668 ( new_n1054 , new_n1053 , pi231 );
  or       g0669 ( new_n1055 , new_n1052 , new_n1054 );
  nand     g0670 ( new_n1056 , new_n1035 , new_n1055 );
  or       g0671 ( new_n1057 , new_n1028 , new_n1056 );
  nand     g0672 ( new_n1058 , new_n951 , new_n930 );
  nand     g0673 ( new_n1059 , pi116 , new_n951 );
  and      g0674 ( new_n1060 , new_n1058 , new_n1059 );
  nand g0675 ( new_n1061 , new_n954 , new_n954 );
  nor      g0676 ( new_n1062 , pi015 , pi086 );
  nand     g0677 ( new_n1063 , new_n1061 , new_n1062 );
  nor      g0678 ( new_n1064 , new_n1060 , new_n1063 );
  nand     g0679 ( new_n1065 , new_n1057 , new_n1064 );
  nor      g0680 ( new_n1066 , new_n1051 , new_n1065 );
  nand g0681 ( new_n1067 , new_n740 , new_n740 );
  nand g0682 ( new_n1068 , pi073 , pi073 );
  nand     g0683 ( new_n1069 , new_n1068 , new_n1053 );
  nand g0684 ( new_n1070 , new_n1069 , new_n1069 );
  nand g0685 ( new_n1071 , pi065 , pi065 );
  nand     g0686 ( new_n1072 , new_n1071 , pi072 );
  nand     g0687 ( new_n1073 , new_n1070 , new_n1072 );
  nand g0688 ( new_n1074 , new_n1073 , new_n1073 );
  nand     g0689 ( new_n1075 , new_n1019 , new_n1074 );
  nor      g0690 ( new_n1076 , new_n1047 , new_n1075 );
  nand     g0691 ( new_n1077 , new_n1064 , new_n1076 );
  nand     g0692 ( new_n1078 , new_n1067 , new_n1077 );
  nor      g0693 ( new_n1079 , new_n1066 , new_n1078 );
  nor      g0694 ( new_n1080 , new_n1017 , new_n1079 );
  nor      g0695 ( new_n1081 , pi124 , pi229 );
  nand     g0696 ( new_n1082 , new_n915 , new_n919 );
  nand     g0697 ( new_n1083 , new_n1013 , new_n1082 );
  nor      g0698 ( new_n1084 , pi052 , pi148 );
  nor      g0699 ( new_n1085 , new_n1083 , new_n1084 );
  nand g0700 ( new_n1086 , pi184 , pi184 );
  nand     g0701 ( new_n1087 , new_n1086 , new_n780 );
  nand     g0702 ( new_n1088 , new_n912 , new_n1013 );
  nand     g0703 ( new_n1089 , new_n1087 , new_n1088 );
  nor      g0704 ( new_n1090 , new_n1085 , new_n1089 );
  nand     g0705 ( new_n1091 , new_n774 , new_n1090 );
  nand     g0706 ( new_n1092 , new_n771 , new_n1091 );
  nand     g0707 ( new_n1093 , new_n1081 , new_n1092 );
  nor      g0708 ( new_n1094 , new_n1080 , new_n1093 );
  nor      g0709 ( new_n1095 , new_n770 , pi229 );
  nand     g0710 ( new_n1096 , new_n747 , pi222 );
  nand     g0711 ( new_n1097 , new_n764 , new_n747 );
  nand     g0712 ( new_n1098 , new_n1096 , new_n1097 );
  nand     g0713 ( new_n1099 , new_n710 , new_n864 );
  nand g0714 ( new_n1100 , pi006 , pi006 );
  nand     g0715 ( new_n1101 , new_n1100 , new_n748 );
  nor      g0716 ( new_n1102 , new_n1099 , new_n1101 );
  nand     g0717 ( new_n1103 , new_n1098 , new_n1102 );
  nand g0718 ( new_n1104 , new_n1103 , new_n1103 );
  nand     g0719 ( new_n1105 , new_n862 , new_n1104 );
  nand g0720 ( new_n1106 , new_n1105 , new_n1105 );
  nand     g0721 ( new_n1107 , new_n791 , new_n1106 );
  nor      g0722 ( new_n1108 , new_n1095 , new_n1107 );
  nand g0723 ( new_n1109 , new_n1108 , new_n1108 );
  nor      g0724 ( new_n1110 , new_n1094 , new_n1109 );
  nand g0725 ( new_n1111 , new_n936 , new_n936 );
  nor      g0726 ( new_n1112 , new_n1111 , new_n1050 );
  nand g0727 ( new_n1113 , new_n1112 , new_n1112 );
  nor      g0728 ( new_n1114 , pi188 , new_n1060 );
  nand     g0729 ( new_n1115 , new_n1113 , new_n1114 );
  nand g0730 ( new_n1116 , new_n1115 , new_n1115 );
  nand g0731 ( new_n1117 , pi072 , pi072 );
  nand     g0732 ( new_n1118 , new_n1117 , pi080 );
  nand     g0733 ( new_n1119 , new_n1071 , new_n1118 );
  nand     g0734 ( new_n1120 , new_n1070 , new_n1119 );
  nand     g0735 ( new_n1121 , new_n1055 , new_n1120 );
  nand g0736 ( new_n1122 , new_n1121 , new_n1121 );
  nand     g0737 ( new_n1123 , new_n1117 , new_n1070 );
  nand g0738 ( new_n1124 , pi213 , pi213 );
  nand     g0739 ( new_n1125 , pi027 , new_n1124 );
  or       g0740 ( new_n1126 , new_n1123 , new_n1125 );
  nand g0741 ( new_n1127 , new_n1126 , new_n1126 );
  nand     g0742 ( new_n1128 , new_n944 , new_n1029 );
  nand g0743 ( new_n1129 , new_n1128 , new_n1128 );
  nand g0744 ( new_n1130 , new_n1032 , new_n1032 );
  nor      g0745 ( new_n1131 , new_n1022 , new_n1130 );
  nand     g0746 ( new_n1132 , new_n1129 , new_n1131 );
  nor      g0747 ( new_n1133 , new_n1127 , new_n1132 );
  nand     g0748 ( new_n1134 , new_n1122 , new_n1133 );
  nand g0749 ( new_n1135 , new_n1134 , new_n1134 );
  nand g0750 ( new_n1136 , new_n1123 , new_n1123 );
  nor      g0751 ( new_n1137 , pi097 , pi213 );
  nand     g0752 ( new_n1138 , pi236 , new_n1137 );
  nand g0753 ( new_n1139 , pi036 , pi036 );
  nand     g0754 ( new_n1140 , new_n1139 , new_n1137 );
  nand     g0755 ( new_n1141 , new_n1138 , new_n1140 );
  nand     g0756 ( new_n1142 , new_n1136 , new_n1141 );
  nand     g0757 ( new_n1143 , new_n1135 , new_n1142 );
  nand     g0758 ( new_n1144 , new_n1116 , new_n1143 );
  nand g0759 ( new_n1145 , new_n746 , new_n746 );
  nand g0760 ( new_n1146 , new_n1026 , new_n1026 );
  nor      g0761 ( new_n1147 , new_n1146 , new_n1040 );
  nand     g0762 ( new_n1148 , new_n733 , new_n942 );
  nand g0763 ( new_n1149 , new_n1148 , new_n1148 );
  nand     g0764 ( new_n1150 , new_n1147 , new_n1149 );
  nor      g0765 ( new_n1151 , new_n1145 , new_n1150 );
  nand     g0766 ( new_n1152 , new_n1144 , new_n1151 );
  nand     g0767 ( new_n1153 , new_n1110 , new_n1152 );
  nand g0768 ( new_n1154 , new_n867 , new_n867 );
  nor      g0769 ( new_n1155 , new_n800 , new_n1154 );
  nand g0770 ( new_n1156 , new_n620 , new_n620 );
  nand     g0771 ( new_n1157 , new_n1156 , new_n962 );
  nand g0772 ( new_n1158 , new_n1157 , new_n1157 );
  nand     g0773 ( new_n1159 , new_n638 , new_n1158 );
  nand     g0774 ( new_n1160 , new_n981 , new_n1159 );
  nand     g0775 ( new_n1161 , new_n990 , new_n1006 );
  nor      g0776 ( new_n1162 , new_n1160 , new_n1161 );
  nand g0777 ( new_n1163 , new_n1162 , new_n1162 );
  nand g0778 ( new_n1164 , new_n906 , new_n906 );
  nand     g0779 ( new_n1165 , new_n729 , new_n1164 );
  nor      g0780 ( new_n1166 , new_n1163 , new_n1165 );
  nand g0781 ( new_n1167 , new_n1166 , new_n1166 );
  nor      g0782 ( new_n1168 , new_n1155 , new_n1167 );
  nand     g0783 ( new_n1169 , new_n1153 , new_n1168 );
  nand     g0784 ( new_n1170 , new_n856 , new_n1164 );
  nand     g0785 ( new_n1171 , new_n599 , new_n880 );
  nand     g0786 ( new_n1172 , new_n589 , new_n1171 );
  nand g0787 ( new_n1173 , new_n1172 , new_n1172 );
  nand     g0788 ( new_n1174 , new_n617 , new_n638 );
  nor      g0789 ( new_n1175 , new_n1173 , new_n1174 );
  nand     g0790 ( new_n1176 , new_n1170 , new_n1175 );
  nand     g0791 ( new_n1177 , new_n1162 , new_n1176 );
  nand     g0792 ( new_n1178 , new_n815 , new_n834 );
  nand     g0793 ( new_n1179 , new_n810 , new_n1178 );
  nand g0794 ( new_n1180 , new_n1179 , new_n1179 );
  or       g0795 ( new_n1181 , new_n720 , new_n841 );
  nand     g0796 ( new_n1182 , new_n1180 , new_n1181 );
  nand g0797 ( new_n1183 , new_n843 , new_n843 );
  nand     g0798 ( new_n1184 , pi134 , new_n722 );
  nand     g0799 ( new_n1185 , new_n1183 , new_n1184 );
  nand g0800 ( new_n1186 , new_n1185 , new_n1185 );
  nand     g0801 ( new_n1187 , new_n1180 , new_n1186 );
  nand     g0802 ( new_n1188 , pi035 , new_n844 );
  nand g0803 ( new_n1189 , new_n1188 , new_n1188 );
  or       g0804 ( new_n1190 , pi132 , pi151 );
  nor      g0805 ( new_n1191 , new_n1189 , new_n1190 );
  or       g0806 ( new_n1192 , new_n1187 , new_n1191 );
  nand     g0807 ( new_n1193 , new_n1182 , new_n1192 );
  nand     g0808 ( new_n1194 , new_n823 , new_n1164 );
  nor      g0809 ( new_n1195 , new_n1193 , new_n1194 );
  nand g0810 ( new_n1196 , new_n1195 , new_n1195 );
  nand g0811 ( new_n1197 , new_n1187 , new_n1187 );
  nand     g0812 ( new_n1198 , new_n711 , new_n1099 );
  nand     g0813 ( new_n1199 , new_n844 , new_n1198 );
  nand g0814 ( new_n1200 , new_n1199 , new_n1199 );
  nand     g0815 ( new_n1201 , new_n1197 , new_n1200 );
  nand     g0816 ( new_n1202 , new_n1162 , new_n1201 );
  nor      g0817 ( new_n1203 , new_n1196 , new_n1202 );
  nor      g0818 ( new_n1204 , new_n499 , new_n536 );
  nand g0819 ( new_n1205 , new_n696 , new_n696 );
  nand     g0820 ( new_n1206 , new_n627 , new_n988 );
  nand g0821 ( new_n1207 , new_n1206 , new_n1206 );
  nor      g0822 ( new_n1208 , new_n705 , new_n1207 );
  or       g0823 ( new_n1209 , new_n1205 , new_n1208 );
  nand     g0824 ( new_n1210 , new_n1204 , new_n1209 );
  nor      g0825 ( new_n1211 , new_n539 , new_n1006 );
  nand     g0826 ( new_n1212 , new_n521 , new_n1211 );
  nand     g0827 ( new_n1213 , new_n1210 , new_n1212 );
  nand g0828 ( new_n1214 , new_n1213 , new_n1213 );
  nor      g0829 ( new_n1215 , new_n1203 , new_n1214 );
  nand     g0830 ( new_n1216 , new_n1177 , new_n1215 );
  nand g0831 ( new_n1217 , new_n1216 , new_n1216 );
  and      g0832 ( new_n1218 , new_n1169 , new_n1217 );
  nand g0833 ( new_n1219 , new_n1168 , new_n1168 );
  nand g0834 ( new_n1220 , pi186 , pi186 );
  nand     g0835 ( new_n1221 , new_n1220 , pi230 );
  nand g0836 ( new_n1222 , new_n1221 , new_n1221 );
  nand g0837 ( new_n1223 , pi122 , pi122 );
  nand g0838 ( new_n1224 , pi236 , pi236 );
  nand     g0839 ( new_n1225 , new_n1223 , new_n1224 );
  nor      g0840 ( new_n1226 , new_n1222 , new_n1225 );
  nand g0841 ( new_n1227 , new_n1226 , new_n1226 );
  nand     g0842 ( new_n1228 , new_n1141 , new_n1227 );
  nand g0843 ( new_n1229 , new_n1228 , new_n1228 );
  nor      g0844 ( new_n1230 , pi065 , pi080 );
  nand     g0845 ( new_n1231 , new_n1125 , new_n1230 );
  nor      g0846 ( new_n1232 , new_n1229 , new_n1231 );
  nand g0847 ( new_n1233 , new_n1232 , new_n1232 );
  nand     g0848 ( new_n1234 , new_n1074 , new_n1233 );
  nand     g0849 ( new_n1235 , new_n746 , new_n1234 );
  or       g0850 ( new_n1236 , new_n1057 , new_n1235 );
  nor      g0851 ( new_n1237 , new_n1219 , new_n1236 );
  nand     g0852 ( new_n1238 , new_n1042 , new_n1121 );
  nand     g0853 ( new_n1239 , new_n1032 , new_n1238 );
  nand g0854 ( new_n1240 , new_n1239 , new_n1239 );
  nand g0855 ( new_n1241 , pi206 , pi206 );
  nand g0856 ( new_n1242 , pi020 , pi020 );
  nand g0857 ( new_n1243 , pi028 , pi028 );
  nand     g0858 ( new_n1244 , new_n1242 , new_n1243 );
  nor      g0859 ( new_n1245 , pi127 , new_n1244 );
  nand     g0860 ( new_n1246 , new_n1241 , new_n1245 );
  nand g0861 ( new_n1247 , new_n1246 , new_n1246 );
  nand g0862 ( new_n1248 , pi099 , pi099 );
  or       g0863 ( new_n1249 , pi029 , new_n1248 );
  and      g0864 ( new_n1250 , new_n1247 , new_n1249 );
  nand g0865 ( new_n1251 , pi230 , pi230 );
  nand     g0866 ( new_n1252 , new_n1223 , new_n1251 );
  nand g0867 ( new_n1253 , pi027 , pi027 );
  nand     g0868 ( new_n1254 , new_n1253 , new_n1224 );
  nor      g0869 ( new_n1255 , new_n1252 , new_n1254 );
  nand     g0870 ( new_n1256 , new_n1250 , new_n1255 );
  nand g0871 ( new_n1257 , new_n1256 , new_n1256 );
  nor      g0872 ( new_n1258 , pi029 , pi032 );
  nand g0873 ( new_n1259 , pi033 , pi033 );
  nand     g0874 ( new_n1260 , new_n1259 , pi131 );
  nand     g0875 ( new_n1261 , new_n1258 , new_n1260 );
  nand     g0876 ( new_n1262 , new_n1257 , new_n1261 );
  nand     g0877 ( new_n1263 , new_n1125 , new_n1138 );
  nand     g0878 ( new_n1264 , new_n1117 , new_n1263 );
  nand g0879 ( new_n1265 , new_n1252 , new_n1252 );
  nand     g0880 ( new_n1266 , pi018 , new_n1245 );
  nand g0881 ( new_n1267 , new_n1266 , new_n1266 );
  nand     g0882 ( new_n1268 , new_n1265 , new_n1267 );
  nand g0883 ( new_n1269 , pi254 , pi254 );
  nand g0884 ( new_n1270 , pi241 , pi241 );
  nand     g0885 ( new_n1271 , pi127 , new_n1270 );
  nand g0886 ( new_n1272 , new_n1271 , new_n1271 );
  nor      g0887 ( new_n1273 , pi212 , pi241 );
  nand g0888 ( new_n1274 , new_n1273 , new_n1273 );
  nand     g0889 ( new_n1275 , new_n1243 , new_n1274 );
  nor      g0890 ( new_n1276 , new_n1272 , new_n1275 );
  nand g0891 ( new_n1277 , new_n1276 , new_n1276 );
  nand     g0892 ( new_n1278 , new_n1269 , new_n1277 );
  nand     g0893 ( new_n1279 , new_n1265 , new_n1278 );
  nand g0894 ( new_n1280 , new_n1279 , new_n1279 );
  nor      g0895 ( new_n1281 , pi072 , new_n1140 );
  nand     g0896 ( new_n1282 , new_n1223 , pi186 );
  nand     g0897 ( new_n1283 , new_n1281 , new_n1282 );
  nor      g0898 ( new_n1284 , new_n1280 , new_n1283 );
  nand     g0899 ( new_n1285 , new_n1268 , new_n1284 );
  nand     g0900 ( new_n1286 , new_n1264 , new_n1285 );
  nand     g0901 ( new_n1287 , new_n1042 , new_n1070 );
  nand g0902 ( new_n1288 , new_n1287 , new_n1287 );
  nand     g0903 ( new_n1289 , new_n1286 , new_n1288 );
  nand g0904 ( new_n1290 , new_n1289 , new_n1289 );
  nand     g0905 ( new_n1291 , new_n1262 , new_n1290 );
  nand     g0906 ( new_n1292 , new_n1240 , new_n1291 );
  nand g0907 ( new_n1293 , new_n1292 , new_n1292 );
  nand     g0908 ( new_n1294 , new_n1237 , new_n1293 );
  nand     g0909 ( new_n1295 , new_n1218 , new_n1294 );
  or       g0910 ( new_n1296 , new_n1012 , new_n1295 );
  or       g0911 ( new_n1297 , new_n456 , new_n484 );
  nor      g0912 ( new_n1298 , new_n456 , new_n564 );
  nand     g0913 ( new_n1299 , new_n422 , new_n470 );
  nor      g0914 ( new_n1300 , new_n1298 , new_n1299 );
  nand     g0915 ( new_n1301 , new_n1297 , new_n1300 );
  nand g0916 ( new_n1302 , new_n1301 , new_n1301 );
  nand     g0917 ( new_n1303 , new_n410 , pi218 );
  nand     g0918 ( new_n1304 , new_n411 , new_n1303 );
  nand     g0919 ( new_n1305 , new_n414 , new_n1304 );
  nand g0920 ( new_n1306 , new_n1305 , new_n1305 );
  nand g0921 ( new_n1307 , pi153 , pi153 );
  nand g0922 ( new_n1308 , pi003 , pi003 );
  nand     g0923 ( new_n1309 , new_n1308 , pi103 );
  nand     g0924 ( new_n1310 , new_n1307 , new_n1309 );
  nand g0925 ( new_n1311 , new_n1310 , new_n1310 );
  nand     g0926 ( new_n1312 , new_n416 , new_n1311 );
  nand g0927 ( new_n1313 , new_n1312 , new_n1312 );
  nand g0928 ( new_n1314 , pi081 , pi081 );
  nand     g0929 ( new_n1315 , new_n1308 , new_n1314 );
  nand     g0930 ( new_n1316 , new_n1313 , new_n1315 );
  or       g0931 ( new_n1317 , pi144 , new_n1316 );
  nand g0932 ( new_n1318 , new_n1317 , new_n1317 );
  nand g0933 ( new_n1319 , pi149 , pi149 );
  nor      g0934 ( new_n1320 , pi022 , pi075 );
  nor      g0935 ( new_n1321 , new_n416 , pi075 );
  nor      g0936 ( new_n1322 , pi144 , new_n1321 );
  nand g0937 ( new_n1323 , new_n1322 , new_n1322 );
  or       g0938 ( new_n1324 , new_n1320 , new_n1323 );
  nand     g0939 ( new_n1325 , new_n1319 , new_n1324 );
  or       g0940 ( new_n1326 , pi218 , new_n1325 );
  nor      g0941 ( new_n1327 , new_n1318 , new_n1326 );
  nand g0942 ( new_n1328 , new_n1327 , new_n1327 );
  nand     g0943 ( new_n1329 , new_n1306 , new_n1328 );
  nand     g0944 ( new_n1330 , new_n421 , new_n1329 );
  nand g0945 ( new_n1331 , new_n1330 , new_n1330 );
  nand     g0946 ( new_n1332 , new_n392 , new_n403 );
  nor      g0947 ( new_n1333 , pi226 , new_n1332 );
  nand     g0948 ( new_n1334 , new_n464 , pi088 );
  nand g0949 ( new_n1335 , pi121 , pi121 );
  nand     g0950 ( new_n1336 , new_n1335 , new_n398 );
  nand g0951 ( new_n1337 , new_n1336 , new_n1336 );
  nand     g0952 ( new_n1338 , new_n1334 , new_n1337 );
  nand g0953 ( new_n1339 , new_n1338 , new_n1338 );
  nand     g0954 ( new_n1340 , new_n1333 , new_n1339 );
  nor      g0955 ( new_n1341 , new_n1328 , new_n1340 );
  nor      g0956 ( new_n1342 , new_n1331 , new_n1341 );
  nor      g0957 ( new_n1343 , new_n1302 , new_n1342 );
  nand     g0958 ( new_n1344 , pi038 , new_n414 );
  nand     g0959 ( new_n1345 , new_n1343 , new_n1344 );
  nand g0960 ( new_n1346 , new_n1345 , new_n1345 );
  nand     g0961 ( new_n1347 , new_n1296 , new_n1346 );
  nor      g0962 ( po000 , new_n386 , new_n1347 );
  nand     g0963 ( new_n1349 , new_n781 , new_n917 );
  nand     g0964 ( new_n1350 , new_n801 , new_n867 );
  nand g0965 ( new_n1351 , new_n1350 , new_n1350 );
  and      g0966 ( new_n1352 , new_n1349 , new_n1351 );
  nand     g0967 ( new_n1353 , new_n769 , new_n786 );
  nor      g0968 ( new_n1354 , new_n799 , new_n1154 );
  nand     g0969 ( new_n1355 , new_n1353 , new_n1354 );
  nand     g0970 ( new_n1356 , new_n714 , new_n1355 );
  nor      g0971 ( new_n1357 , new_n1352 , new_n1356 );
  and      g0972 ( new_n1358 , new_n727 , new_n896 );
  nand     g0973 ( new_n1359 , new_n1357 , new_n1358 );
  nand     g0974 ( new_n1360 , new_n823 , new_n896 );
  nand     g0975 ( new_n1361 , new_n892 , pi225 );
  nand     g0976 ( new_n1362 , new_n825 , new_n1361 );
  nor      g0977 ( new_n1363 , pi039 , new_n1362 );
  nand     g0978 ( new_n1364 , new_n674 , pi054 );
  nand     g0979 ( new_n1365 , new_n891 , new_n1364 );
  nor      g0980 ( new_n1366 , new_n1363 , new_n1365 );
  nand g0981 ( new_n1367 , new_n1366 , new_n1366 );
  nand     g0982 ( new_n1368 , new_n1360 , new_n1367 );
  nand g0983 ( new_n1369 , new_n1368 , new_n1368 );
  nor      g0984 ( new_n1370 , new_n852 , new_n1369 );
  nor      g0985 ( new_n1371 , new_n679 , new_n1370 );
  nand     g0986 ( new_n1372 , new_n1359 , new_n1371 );
  nand     g0987 ( new_n1373 , new_n608 , new_n668 );
  nand     g0988 ( new_n1374 , new_n1372 , new_n1373 );
  nand g0989 ( new_n1375 , new_n736 , new_n736 );
  nand g0990 ( new_n1376 , new_n1114 , new_n1114 );
  nand g0991 ( new_n1377 , new_n939 , new_n939 );
  nor      g0992 ( new_n1378 , pi116 , new_n1377 );
  nor      g0993 ( new_n1379 , new_n1376 , new_n1378 );
  nor      g0994 ( new_n1380 , new_n1375 , new_n1379 );
  nand     g0995 ( new_n1381 , new_n1115 , new_n1380 );
  nand g0996 ( new_n1382 , new_n1381 , new_n1381 );
  nand     g0997 ( new_n1383 , new_n921 , new_n1351 );
  nor      g0998 ( new_n1384 , new_n1382 , new_n1383 );
  nand     g0999 ( new_n1385 , new_n1371 , new_n1384 );
  nand g1000 ( new_n1386 , pi131 , pi131 );
  nand     g1001 ( new_n1387 , new_n1386 , new_n414 );
  nand g1002 ( new_n1388 , new_n1387 , new_n1387 );
  nand g1003 ( new_n1389 , new_n1258 , new_n1258 );
  nor      g1004 ( new_n1390 , pi018 , new_n1389 );
  nand     g1005 ( new_n1391 , new_n1273 , new_n1390 );
  nand g1006 ( new_n1392 , new_n1391 , new_n1391 );
  nand     g1007 ( new_n1393 , new_n1388 , new_n1392 );
  nor      g1008 ( new_n1394 , new_n1250 , new_n1267 );
  nand g1009 ( new_n1395 , new_n1394 , new_n1394 );
  nand     g1010 ( new_n1396 , new_n1259 , new_n386 );
  nand     g1011 ( new_n1397 , new_n1260 , new_n1396 );
  nand g1012 ( new_n1398 , new_n1397 , new_n1397 );
  nand     g1013 ( new_n1399 , new_n1390 , new_n1398 );
  and      g1014 ( new_n1400 , new_n1395 , new_n1399 );
  nand     g1015 ( new_n1401 , new_n1393 , new_n1400 );
  nand     g1016 ( new_n1402 , new_n1220 , new_n1269 );
  nor      g1017 ( new_n1403 , new_n1276 , new_n1402 );
  nand     g1018 ( new_n1404 , new_n1401 , new_n1403 );
  nand g1019 ( new_n1405 , pi038 , pi038 );
  nand     g1020 ( new_n1406 , new_n1405 , new_n1303 );
  nor      g1021 ( new_n1407 , new_n1396 , new_n1406 );
  nand     g1022 ( new_n1408 , new_n1250 , new_n1407 );
  nand g1023 ( new_n1409 , new_n1408 , new_n1408 );
  nor      g1024 ( new_n1410 , new_n1404 , new_n1409 );
  nor      g1025 ( new_n1411 , new_n1227 , new_n1410 );
  or       g1026 ( new_n1412 , new_n1142 , new_n1411 );
  nand g1027 ( new_n1413 , new_n1412 , new_n1412 );
  nand     g1028 ( new_n1414 , new_n1135 , new_n1380 );
  nor      g1029 ( new_n1415 , new_n1413 , new_n1414 );
  nor      g1030 ( new_n1416 , new_n1385 , new_n1415 );
  nor      g1031 ( new_n1417 , new_n1374 , new_n1416 );
  nand g1032 ( new_n1418 , new_n630 , new_n630 );
  nand     g1033 ( new_n1419 , new_n1418 , new_n976 );
  nand g1034 ( new_n1420 , new_n1419 , new_n1419 );
  nor      g1035 ( new_n1421 , pi019 , pi037 );
  nand g1036 ( new_n1422 , new_n1421 , new_n1421 );
  nand     g1037 ( new_n1423 , new_n622 , new_n697 );
  nor      g1038 ( new_n1424 , new_n1422 , new_n1423 );
  nand     g1039 ( new_n1425 , new_n1420 , new_n1424 );
  nand     g1040 ( new_n1426 , new_n1208 , new_n1425 );
  nand g1041 ( new_n1427 , new_n470 , new_n470 );
  nand g1042 ( new_n1428 , new_n455 , new_n455 );
  nor      g1043 ( new_n1429 , new_n429 , new_n1428 );
  nor      g1044 ( new_n1430 , new_n1427 , new_n1429 );
  nor      g1045 ( new_n1431 , new_n1338 , new_n1430 );
  nand g1046 ( new_n1432 , pi088 , pi088 );
  nand     g1047 ( new_n1433 , new_n1432 , new_n455 );
  nand g1048 ( new_n1434 , new_n444 , new_n444 );
  nand     g1049 ( new_n1435 , new_n1434 , new_n1337 );
  nor      g1050 ( new_n1436 , new_n1433 , new_n1435 );
  nand g1051 ( new_n1437 , new_n1436 , new_n1436 );
  nand g1052 ( new_n1438 , new_n442 , new_n442 );
  nand     g1053 ( new_n1439 , new_n432 , new_n1438 );
  nor      g1054 ( new_n1440 , new_n1437 , new_n1439 );
  nor      g1055 ( new_n1441 , new_n1431 , new_n1440 );
  nand g1056 ( new_n1442 , new_n1441 , new_n1441 );
  nand     g1057 ( new_n1443 , new_n474 , new_n562 );
  nand     g1058 ( new_n1444 , new_n437 , new_n1443 );
  nand g1059 ( new_n1445 , new_n1444 , new_n1444 );
  nand g1060 ( new_n1446 , pi214 , pi214 );
  nand     g1061 ( new_n1447 , new_n559 , new_n1446 );
  nor      g1062 ( new_n1448 , pi204 , new_n1447 );
  nand     g1063 ( new_n1449 , new_n554 , new_n1448 );
  nand     g1064 ( new_n1450 , new_n1445 , new_n1449 );
  nor      g1065 ( new_n1451 , pi030 , pi237 );
  nand     g1066 ( new_n1452 , new_n1436 , new_n1451 );
  nor      g1067 ( new_n1453 , new_n1450 , new_n1452 );
  nor      g1068 ( new_n1454 , new_n1442 , new_n1453 );
  nand g1069 ( new_n1455 , new_n1315 , new_n1315 );
  nand     g1070 ( new_n1456 , new_n387 , new_n405 );
  nand     g1071 ( new_n1457 , new_n1455 , new_n1456 );
  nand     g1072 ( new_n1458 , new_n1319 , new_n1320 );
  nand g1073 ( new_n1459 , new_n1396 , new_n1396 );
  nand g1074 ( new_n1460 , pi218 , pi218 );
  nand     g1075 ( new_n1461 , new_n1405 , new_n1460 );
  nand g1076 ( new_n1462 , new_n1461 , new_n1461 );
  nand     g1077 ( new_n1463 , new_n1459 , new_n1462 );
  nor      g1078 ( new_n1464 , new_n1458 , new_n1463 );
  nand     g1079 ( new_n1465 , new_n392 , new_n1464 );
  nor      g1080 ( new_n1466 , new_n1457 , new_n1465 );
  nand g1081 ( new_n1467 , new_n1466 , new_n1466 );
  nor      g1082 ( new_n1468 , new_n1454 , new_n1467 );
  nand g1083 ( new_n1469 , pi252 , pi252 );
  nand     g1084 ( new_n1470 , new_n1469 , new_n481 );
  nand g1085 ( new_n1471 , new_n1470 , new_n1470 );
  nand     g1086 ( new_n1472 , new_n1006 , new_n1471 );
  nor      g1087 ( new_n1473 , new_n1205 , new_n1472 );
  nand     g1088 ( new_n1474 , new_n1468 , new_n1473 );
  nand g1089 ( new_n1475 , new_n1474 , new_n1474 );
  nand     g1090 ( new_n1476 , new_n1426 , new_n1475 );
  nand     g1091 ( new_n1477 , new_n567 , new_n1468 );
  nand     g1092 ( new_n1478 , new_n1344 , new_n1459 );
  nor      g1093 ( new_n1479 , new_n1330 , new_n1478 );
  nand g1094 ( new_n1480 , new_n1479 , new_n1479 );
  nand g1095 ( new_n1481 , new_n1281 , new_n1281 );
  nand     g1096 ( new_n1482 , new_n1221 , new_n1402 );
  nand     g1097 ( new_n1483 , new_n1288 , new_n1482 );
  nor      g1098 ( new_n1484 , new_n1481 , new_n1483 );
  nand g1099 ( new_n1485 , new_n1484 , new_n1484 );
  nand     g1100 ( new_n1486 , new_n1260 , new_n1392 );
  nor      g1101 ( new_n1487 , new_n1485 , new_n1486 );
  nand g1102 ( new_n1488 , new_n1487 , new_n1487 );
  nand     g1103 ( new_n1489 , new_n1041 , new_n1044 );
  nor      g1104 ( new_n1490 , new_n1488 , new_n1489 );
  and      g1105 ( new_n1491 , new_n1480 , new_n1490 );
  nand     g1106 ( new_n1492 , new_n1477 , new_n1491 );
  nand g1107 ( new_n1493 , new_n1492 , new_n1492 );
  nand     g1108 ( new_n1494 , new_n1476 , new_n1493 );
  nand     g1109 ( new_n1495 , new_n1417 , new_n1494 );
  nand g1110 ( new_n1496 , pi026 , pi026 );
  nand     g1111 ( new_n1497 , new_n1496 , new_n610 );
  nand g1112 ( new_n1498 , new_n1497 , new_n1497 );
  nand     g1113 ( new_n1499 , new_n611 , new_n1498 );
  nor      g1114 ( new_n1500 , new_n856 , new_n1499 );
  nand     g1115 ( new_n1501 , new_n673 , new_n1500 );
  nor      g1116 ( new_n1502 , new_n1201 , new_n1501 );
  nand g1117 ( new_n1503 , new_n1502 , new_n1502 );
  nand g1118 ( new_n1504 , new_n943 , new_n943 );
  nand g1119 ( new_n1505 , pi137 , pi137 );
  nand     g1120 ( new_n1506 , pi085 , new_n1505 );
  nand g1121 ( new_n1507 , new_n1506 , new_n1506 );
  nand     g1122 ( new_n1508 , new_n1037 , new_n944 );
  nor      g1123 ( new_n1509 , new_n1507 , new_n1508 );
  nand g1124 ( new_n1510 , new_n1509 , new_n1509 );
  nand     g1125 ( new_n1511 , new_n1031 , new_n1044 );
  nand     g1126 ( new_n1512 , pi122 , new_n1281 );
  nand     g1127 ( new_n1513 , new_n1264 , new_n1512 );
  nand     g1128 ( new_n1514 , new_n1288 , new_n1513 );
  nand g1129 ( new_n1515 , new_n1514 , new_n1514 );
  nand     g1130 ( new_n1516 , new_n1240 , new_n1485 );
  nor      g1131 ( new_n1517 , new_n1515 , new_n1516 );
  nor      g1132 ( new_n1518 , new_n1511 , new_n1517 );
  nor      g1133 ( new_n1519 , new_n1510 , new_n1518 );
  nand     g1134 ( new_n1520 , new_n1277 , new_n1394 );
  nand g1135 ( new_n1521 , new_n1520 , new_n1520 );
  nand     g1136 ( new_n1522 , new_n1052 , new_n1230 );
  nor      g1137 ( new_n1523 , new_n1130 , new_n1522 );
  nand g1138 ( new_n1524 , new_n1523 , new_n1523 );
  nand     g1139 ( new_n1525 , new_n1129 , new_n1265 );
  nor      g1140 ( new_n1526 , new_n1524 , new_n1525 );
  nand     g1141 ( new_n1527 , new_n1264 , new_n1526 );
  nor      g1142 ( new_n1528 , new_n1521 , new_n1527 );
  nor      g1143 ( new_n1529 , new_n1519 , new_n1528 );
  nand g1144 ( new_n1530 , new_n1529 , new_n1529 );
  nand     g1145 ( new_n1531 , new_n1504 , new_n1530 );
  nand     g1146 ( new_n1532 , new_n1068 , new_n1284 );
  or       g1147 ( new_n1533 , new_n1252 , new_n1390 );
  nor      g1148 ( new_n1534 , new_n1394 , new_n1533 );
  nor      g1149 ( new_n1535 , new_n1532 , new_n1534 );
  nand g1150 ( new_n1536 , new_n1535 , new_n1535 );
  nand     g1151 ( new_n1537 , new_n1405 , pi090 );
  nand     g1152 ( new_n1538 , new_n1388 , new_n1537 );
  nand g1153 ( new_n1539 , new_n1538 , new_n1538 );
  nand     g1154 ( new_n1540 , new_n409 , new_n1322 );
  nand g1155 ( new_n1541 , new_n1540 , new_n1540 );
  nand     g1156 ( new_n1542 , new_n1539 , new_n1541 );
  nand     g1157 ( new_n1543 , new_n409 , pi149 );
  nand     g1158 ( new_n1544 , new_n1462 , new_n1543 );
  nand     g1159 ( new_n1545 , new_n1539 , new_n1544 );
  nand g1160 ( new_n1546 , new_n1545 , new_n1545 );
  nand     g1161 ( new_n1547 , new_n1248 , new_n1265 );
  nor      g1162 ( new_n1548 , new_n1398 , new_n1547 );
  nand     g1163 ( new_n1549 , new_n1247 , new_n1548 );
  nor      g1164 ( new_n1550 , new_n1546 , new_n1549 );
  nand     g1165 ( new_n1551 , new_n1542 , new_n1550 );
  nor      g1166 ( new_n1552 , new_n1018 , new_n1058 );
  nand g1167 ( new_n1553 , new_n1552 , new_n1552 );
  nand     g1168 ( new_n1554 , new_n1053 , new_n1046 );
  nor      g1169 ( new_n1555 , new_n1553 , new_n1554 );
  nand     g1170 ( new_n1556 , new_n1551 , new_n1555 );
  nor      g1171 ( new_n1557 , new_n1536 , new_n1556 );
  nor      g1172 ( new_n1558 , new_n1531 , new_n1557 );
  nand     g1173 ( new_n1559 , new_n1036 , new_n1061 );
  nor      g1174 ( new_n1560 , new_n1511 , new_n1559 );
  nand     g1175 ( new_n1561 , new_n1552 , new_n1560 );
  nand     g1176 ( new_n1562 , new_n1504 , new_n1509 );
  nand     g1177 ( new_n1563 , new_n957 , new_n1562 );
  nand g1178 ( new_n1564 , new_n1563 , new_n1563 );
  nand     g1179 ( new_n1565 , pi048 , new_n953 );
  nand     g1180 ( new_n1566 , new_n1084 , new_n1565 );
  nor      g1181 ( new_n1567 , new_n1564 , new_n1566 );
  nand     g1182 ( new_n1568 , new_n1561 , new_n1567 );
  nor      g1183 ( new_n1569 , pi006 , new_n753 );
  nand g1184 ( new_n1570 , pi150 , pi150 );
  nand     g1185 ( new_n1571 , new_n1570 , pi160 );
  nand g1186 ( new_n1572 , new_n1571 , new_n1571 );
  nor      g1187 ( new_n1573 , new_n1097 , new_n1572 );
  nand     g1188 ( new_n1574 , new_n1569 , new_n1573 );
  nand g1189 ( new_n1575 , new_n1083 , new_n1083 );
  nor      g1190 ( new_n1576 , pi209 , new_n772 );
  nand     g1191 ( new_n1577 , new_n1575 , new_n1576 );
  nor      g1192 ( new_n1578 , new_n1574 , new_n1577 );
  nand     g1193 ( new_n1579 , new_n1568 , new_n1578 );
  nor      g1194 ( new_n1580 , new_n1558 , new_n1579 );
  nand     g1195 ( new_n1581 , new_n754 , new_n1096 );
  nand     g1196 ( new_n1582 , new_n1569 , new_n1581 );
  nand     g1197 ( new_n1583 , new_n1100 , pi046 );
  nand g1198 ( new_n1584 , new_n1583 , new_n1583 );
  nand g1199 ( new_n1585 , pi055 , pi055 );
  nand     g1200 ( new_n1586 , new_n1585 , new_n757 );
  nor      g1201 ( new_n1587 , new_n1584 , new_n1586 );
  nand     g1202 ( new_n1588 , new_n1582 , new_n1587 );
  nand     g1203 ( new_n1589 , new_n787 , new_n795 );
  nor      g1204 ( new_n1590 , pi150 , new_n1576 );
  nand     g1205 ( new_n1591 , new_n1589 , new_n1590 );
  nand g1206 ( new_n1592 , new_n1591 , new_n1591 );
  nor      g1207 ( new_n1593 , new_n1574 , new_n1592 );
  nand g1208 ( new_n1594 , new_n1593 , new_n1593 );
  nand g1209 ( new_n1595 , new_n1090 , new_n1090 );
  nand     g1210 ( new_n1596 , new_n793 , new_n774 );
  nor      g1211 ( new_n1597 , pi150 , new_n1596 );
  nand     g1212 ( new_n1598 , new_n1081 , new_n1597 );
  nand g1213 ( new_n1599 , new_n1598 , new_n1598 );
  or       g1214 ( new_n1600 , new_n1083 , new_n1565 );
  nand     g1215 ( new_n1601 , new_n1599 , new_n1600 );
  nor      g1216 ( new_n1602 , new_n1595 , new_n1601 );
  nor      g1217 ( new_n1603 , new_n1594 , new_n1602 );
  nor      g1218 ( new_n1604 , new_n1588 , new_n1603 );
  nand g1219 ( new_n1605 , new_n1604 , new_n1604 );
  nor      g1220 ( new_n1606 , new_n1580 , new_n1605 );
  nor      g1221 ( new_n1607 , new_n1503 , new_n1606 );
  and      g1222 ( new_n1608 , new_n1495 , new_n1607 );
  nand     g1223 ( new_n1609 , new_n655 , new_n671 );
  nand     g1224 ( new_n1610 , new_n879 , new_n1609 );
  or       g1225 ( new_n1611 , pi195 , new_n1366 );
  nand     g1226 ( new_n1612 , new_n643 , new_n903 );
  nand     g1227 ( new_n1613 , new_n890 , new_n661 );
  nor      g1228 ( new_n1614 , new_n1612 , new_n1613 );
  nand     g1229 ( new_n1615 , new_n1611 , new_n1614 );
  and      g1230 ( new_n1616 , new_n597 , new_n1615 );
  and      g1231 ( new_n1617 , new_n1610 , new_n1616 );
  nand     g1232 ( new_n1618 , new_n585 , new_n1617 );
  nand     g1233 ( new_n1619 , new_n589 , new_n1618 );
  nor      g1234 ( new_n1620 , new_n1195 , new_n1499 );
  nand     g1235 ( new_n1621 , new_n1619 , new_n1620 );
  nand g1236 ( new_n1622 , pi063 , pi063 );
  nand     g1237 ( new_n1623 , new_n1622 , new_n571 );
  nor      g1238 ( new_n1624 , pi026 , new_n1157 );
  nor      g1239 ( new_n1625 , new_n1623 , new_n1624 );
  nand     g1240 ( new_n1626 , new_n1621 , new_n1625 );
  nor      g1241 ( new_n1627 , new_n1608 , new_n1626 );
  nand     g1242 ( new_n1628 , new_n1622 , pi100 );
  nand     g1243 ( new_n1629 , new_n631 , new_n1628 );
  nor      g1244 ( new_n1630 , new_n1627 , new_n1629 );
  nand     g1245 ( new_n1631 , pi174 , new_n970 );
  nor      g1246 ( po001 , new_n1630 , new_n1631 );
  nand     g1247 ( new_n1633 , new_n1582 , new_n1594 );
  nand     g1248 ( new_n1634 , new_n763 , new_n1599 );
  nor      g1249 ( new_n1635 , new_n1089 , new_n1634 );
  nand g1250 ( new_n1636 , new_n1635 , new_n1635 );
  nand     g1251 ( new_n1637 , new_n1633 , new_n1636 );
  nand     g1252 ( new_n1638 , new_n1587 , new_n1637 );
  nand     g1253 ( new_n1639 , new_n1200 , new_n1638 );
  nand     g1254 ( new_n1640 , new_n1191 , new_n1639 );
  nand g1255 ( new_n1641 , new_n1177 , new_n1177 );
  or       g1256 ( new_n1642 , new_n1641 , new_n1494 );
  nor      g1257 ( new_n1643 , new_n1343 , new_n1488 );
  nand g1258 ( new_n1644 , new_n1478 , new_n1478 );
  nor      g1259 ( new_n1645 , new_n1261 , new_n1644 );
  nor      g1260 ( new_n1646 , new_n1256 , new_n1645 );
  nand g1261 ( new_n1647 , new_n1646 , new_n1646 );
  nand     g1262 ( new_n1648 , new_n1290 , new_n1647 );
  nand g1263 ( new_n1649 , new_n1648 , new_n1648 );
  nand     g1264 ( new_n1650 , new_n1029 , new_n1084 );
  nor      g1265 ( new_n1651 , new_n1148 , new_n1650 );
  nand     g1266 ( new_n1652 , new_n1026 , new_n1651 );
  or       g1267 ( new_n1653 , new_n1239 , new_n1652 );
  nor      g1268 ( new_n1654 , new_n1649 , new_n1653 );
  nand g1269 ( new_n1655 , new_n1654 , new_n1654 );
  nor      g1270 ( new_n1656 , new_n1643 , new_n1655 );
  and      g1271 ( new_n1657 , new_n1642 , new_n1656 );
  nand g1272 ( new_n1658 , new_n1579 , new_n1579 );
  nand     g1273 ( new_n1659 , new_n1200 , new_n1658 );
  nor      g1274 ( new_n1660 , new_n1657 , new_n1659 );
  nor      g1275 ( new_n1661 , new_n1640 , new_n1660 );
  or       g1276 ( new_n1662 , new_n1187 , new_n1661 );
  nand     g1277 ( new_n1663 , new_n1182 , new_n1662 );
  nand     g1278 ( new_n1664 , new_n892 , new_n823 );
  nor      g1279 ( new_n1665 , new_n1663 , new_n1664 );
  nor      g1280 ( new_n1666 , new_n1362 , new_n1665 );
  nor      g1281 ( po002 , new_n884 , new_n1666 );
  nand g1282 ( new_n1668 , new_n832 , new_n832 );
  nand g1283 ( new_n1669 , pi040 , pi040 );
  nand g1284 ( new_n1670 , pi107 , pi107 );
  nand     g1285 ( new_n1671 , new_n973 , new_n1670 );
  nand g1286 ( new_n1672 , new_n1671 , new_n1671 );
  nand     g1287 ( new_n1673 , new_n1622 , new_n967 );
  nor      g1288 ( new_n1674 , pi180 , new_n1673 );
  nand     g1289 ( new_n1675 , new_n1672 , new_n1674 );
  nand     g1290 ( new_n1676 , new_n622 , new_n990 );
  nor      g1291 ( new_n1677 , new_n1675 , new_n1676 );
  nand     g1292 ( new_n1678 , new_n963 , new_n1677 );
  nor      g1293 ( new_n1679 , new_n1194 , new_n1678 );
  nand     g1294 ( new_n1680 , new_n1212 , new_n1679 );
  nor      g1295 ( new_n1681 , new_n1640 , new_n1680 );
  nand     g1296 ( new_n1682 , new_n1656 , new_n1681 );
  nand     g1297 ( new_n1683 , new_n1186 , new_n1682 );
  nor      g1298 ( new_n1684 , new_n1661 , new_n1683 );
  nand     g1299 ( new_n1685 , new_n840 , new_n1662 );
  nor      g1300 ( new_n1686 , new_n1684 , new_n1685 );
  nand     g1301 ( new_n1687 , new_n715 , new_n1686 );
  nand     g1302 ( new_n1688 , new_n1669 , new_n1687 );
  nor      g1303 ( new_n1689 , pi024 , new_n1688 );
  nor      g1304 ( new_n1690 , new_n1668 , new_n1689 );
  nor      g1305 ( new_n1691 , pi087 , new_n1690 );
  nor      g1306 ( po003 , new_n813 , new_n1691 );
  nand g1307 ( new_n1693 , pi215 , pi215 );
  nand     g1308 ( new_n1694 , pi041 , new_n530 );
  nand g1309 ( new_n1695 , new_n510 , new_n510 );
  nand     g1310 ( new_n1696 , new_n497 , new_n1695 );
  nand g1311 ( new_n1697 , new_n1696 , new_n1696 );
  nand     g1312 ( new_n1698 , new_n999 , new_n1697 );
  nand     g1313 ( new_n1699 , new_n491 , new_n1698 );
  nand     g1314 ( new_n1700 , new_n1000 , new_n1699 );
  nand g1315 ( new_n1701 , new_n1700 , new_n1700 );
  nand g1316 ( new_n1702 , pi106 , pi106 );
  nand     g1317 ( new_n1703 , new_n1702 , new_n685 );
  nand g1318 ( new_n1704 , new_n1703 , new_n1703 );
  nand     g1319 ( new_n1705 , new_n697 , new_n1704 );
  nand g1320 ( new_n1706 , new_n1705 , new_n1705 );
  nand     g1321 ( new_n1707 , new_n994 , new_n1706 );
  nand g1322 ( new_n1708 , new_n1707 , new_n1707 );
  nand g1323 ( new_n1709 , new_n1629 , new_n1629 );
  nand     g1324 ( new_n1710 , new_n1623 , new_n1709 );
  nand g1325 ( new_n1711 , new_n1710 , new_n1710 );
  nor      g1326 ( new_n1712 , new_n971 , new_n1711 );
  nand     g1327 ( new_n1713 , new_n1672 , new_n1712 );
  nand g1328 ( new_n1714 , new_n1713 , new_n1713 );
  nand     g1329 ( new_n1715 , new_n624 , new_n1419 );
  nor      g1330 ( new_n1716 , new_n1714 , new_n1715 );
  nand     g1331 ( new_n1717 , new_n623 , new_n1421 );
  nand     g1332 ( new_n1718 , new_n1496 , pi163 );
  nand     g1333 ( new_n1719 , new_n1497 , new_n1718 );
  nand     g1334 ( new_n1720 , new_n624 , new_n1719 );
  nor      g1335 ( new_n1721 , new_n634 , new_n1720 );
  nand g1336 ( new_n1722 , new_n1721 , new_n1721 );
  nand     g1337 ( new_n1723 , new_n570 , new_n569 );
  nor      g1338 ( new_n1724 , new_n613 , new_n1723 );
  nor      g1339 ( new_n1725 , new_n1722 , new_n1724 );
  nor      g1340 ( new_n1726 , new_n1717 , new_n1725 );
  nand g1341 ( new_n1727 , new_n1726 , new_n1726 );
  nor      g1342 ( new_n1728 , new_n1716 , new_n1727 );
  nand     g1343 ( new_n1729 , new_n1708 , new_n1728 );
  nand g1344 ( new_n1730 , new_n1729 , new_n1729 );
  nand     g1345 ( new_n1731 , new_n1701 , new_n1730 );
  nand     g1346 ( new_n1732 , new_n1570 , new_n761 );
  nand g1347 ( new_n1733 , new_n1732 , new_n1732 );
  nand     g1348 ( new_n1734 , new_n1589 , new_n1733 );
  nand     g1349 ( new_n1735 , new_n770 , new_n791 );
  nor      g1350 ( new_n1736 , new_n1092 , new_n1735 );
  nor      g1351 ( new_n1737 , new_n1734 , new_n1736 );
  nand     g1352 ( new_n1738 , new_n954 , new_n1565 );
  nor      g1353 ( new_n1739 , pi015 , new_n1735 );
  nand     g1354 ( new_n1740 , new_n1738 , new_n1739 );
  nor      g1355 ( new_n1741 , new_n1017 , new_n1740 );
  nand g1356 ( new_n1742 , new_n1741 , new_n1741 );
  nand     g1357 ( new_n1743 , new_n1737 , new_n1742 );
  nor      g1358 ( new_n1744 , new_n810 , new_n820 );
  nor      g1359 ( new_n1745 , pi225 , new_n1744 );
  nand g1360 ( new_n1746 , new_n1745 , new_n1745 );
  nor      g1361 ( new_n1747 , new_n1105 , new_n1746 );
  nand     g1362 ( new_n1748 , new_n1743 , new_n1747 );
  or       g1363 ( new_n1749 , new_n1734 , new_n1736 );
  nor      g1364 ( new_n1750 , pi048 , new_n957 );
  or       g1365 ( new_n1751 , new_n1047 , new_n1054 );
  nand g1366 ( new_n1752 , new_n1751 , new_n1751 );
  or       g1367 ( new_n1753 , new_n1150 , new_n1752 );
  nand     g1368 ( new_n1754 , new_n1741 , new_n1753 );
  nor      g1369 ( new_n1755 , new_n1750 , new_n1754 );
  nor      g1370 ( new_n1756 , new_n1749 , new_n1755 );
  nor      g1371 ( new_n1757 , new_n1748 , new_n1756 );
  nand g1372 ( new_n1758 , new_n1264 , new_n1264 );
  or       g1373 ( new_n1759 , new_n1119 , new_n1758 );
  nand     g1374 ( new_n1760 , new_n1068 , new_n1759 );
  nand     g1375 ( new_n1761 , new_n1052 , new_n1760 );
  nor      g1376 ( new_n1762 , new_n1150 , new_n1761 );
  nand     g1377 ( new_n1763 , new_n1737 , new_n1762 );
  nand     g1378 ( new_n1764 , new_n1757 , new_n1763 );
  nand     g1379 ( new_n1765 , new_n836 , new_n1745 );
  nand g1380 ( new_n1766 , new_n1765 , new_n1765 );
  nand     g1381 ( new_n1767 , pi173 , new_n826 );
  nand     g1382 ( new_n1768 , new_n894 , new_n1767 );
  nor      g1383 ( new_n1769 , new_n1766 , new_n1768 );
  nand     g1384 ( new_n1770 , new_n1764 , new_n1769 );
  nand g1385 ( new_n1771 , new_n718 , new_n718 );
  or       g1386 ( new_n1772 , new_n759 , new_n1154 );
  nand g1387 ( new_n1773 , new_n1772 , new_n1772 );
  nand     g1388 ( new_n1774 , new_n714 , new_n724 );
  nor      g1389 ( new_n1775 , new_n1773 , new_n1774 );
  nor      g1390 ( new_n1776 , new_n849 , new_n1775 );
  nor      g1391 ( new_n1777 , new_n1771 , new_n1776 );
  or       g1392 ( new_n1778 , new_n834 , new_n1777 );
  nor      g1393 ( new_n1779 , new_n1746 , new_n1778 );
  nor      g1394 ( new_n1780 , new_n1770 , new_n1779 );
  nor      g1395 ( new_n1781 , new_n883 , new_n1612 );
  nand     g1396 ( new_n1782 , new_n665 , new_n1781 );
  nand g1397 ( new_n1783 , new_n1782 , new_n1782 );
  nand     g1398 ( new_n1784 , new_n1780 , new_n1783 );
  or       g1399 ( new_n1785 , new_n1731 , new_n1784 );
  nand g1400 ( new_n1786 , new_n1785 , new_n1785 );
  nand g1401 ( new_n1787 , new_n1748 , new_n1748 );
  nand     g1402 ( new_n1788 , new_n1557 , new_n1787 );
  nand g1403 ( new_n1789 , new_n1788 , new_n1788 );
  nand     g1404 ( new_n1790 , new_n1247 , new_n1523 );
  nand g1405 ( new_n1791 , new_n1790 , new_n1790 );
  nand     g1406 ( new_n1792 , new_n1248 , new_n1255 );
  nor      g1407 ( new_n1793 , new_n1478 , new_n1792 );
  nand     g1408 ( new_n1794 , new_n1791 , new_n1793 );
  nor      g1409 ( new_n1795 , new_n1342 , new_n1794 );
  nand g1410 ( new_n1796 , new_n1795 , new_n1795 );
  nor      g1411 ( new_n1797 , new_n1300 , new_n1796 );
  nor      g1412 ( new_n1798 , new_n919 , new_n1561 );
  nand     g1413 ( new_n1799 , new_n1292 , new_n1798 );
  nor      g1414 ( new_n1800 , new_n1797 , new_n1799 );
  nor      g1415 ( new_n1801 , new_n428 , new_n1434 );
  nor      g1416 ( new_n1802 , pi126 , new_n1801 );
  nand g1417 ( new_n1803 , pi126 , pi126 );
  nand     g1418 ( new_n1804 , pi120 , new_n1803 );
  nand     g1419 ( new_n1805 , new_n457 , new_n1804 );
  nor      g1420 ( new_n1806 , new_n1802 , new_n1805 );
  nand g1421 ( new_n1807 , new_n1806 , new_n1806 );
  nor      g1422 ( new_n1808 , new_n396 , new_n415 );
  nand g1423 ( new_n1809 , pi207 , pi207 );
  nand     g1424 ( new_n1810 , new_n459 , new_n1809 );
  nand g1425 ( new_n1811 , new_n1810 , new_n1810 );
  nand g1426 ( new_n1812 , pi117 , pi117 );
  nand     g1427 ( new_n1813 , new_n464 , new_n1812 );
  nand g1428 ( new_n1814 , new_n1813 , new_n1813 );
  nand     g1429 ( new_n1815 , new_n466 , new_n1814 );
  nand g1430 ( new_n1816 , new_n1815 , new_n1815 );
  nand     g1431 ( new_n1817 , new_n1811 , new_n1816 );
  nand g1432 ( new_n1818 , new_n1817 , new_n1817 );
  nand     g1433 ( new_n1819 , new_n1808 , new_n1818 );
  nor      g1434 ( new_n1820 , new_n1807 , new_n1819 );
  nand g1435 ( new_n1821 , new_n1820 , new_n1820 );
  nand     g1436 ( new_n1822 , new_n1311 , new_n1457 );
  nand     g1437 ( new_n1823 , new_n1320 , new_n1822 );
  nand g1438 ( new_n1824 , new_n1823 , new_n1823 );
  nand     g1439 ( new_n1825 , new_n1812 , pi121 );
  nand     g1440 ( new_n1826 , new_n400 , new_n1825 );
  nand     g1441 ( new_n1827 , new_n1808 , new_n1826 );
  nand     g1442 ( new_n1828 , new_n1824 , new_n1827 );
  nand     g1443 ( new_n1829 , new_n1432 , new_n465 );
  nand g1444 ( new_n1830 , new_n1829 , new_n1829 );
  nand     g1445 ( new_n1831 , new_n1809 , pi232 );
  nand     g1446 ( new_n1832 , new_n451 , new_n1831 );
  or       g1447 ( new_n1833 , pi016 , new_n1832 );
  nand     g1448 ( new_n1834 , pi012 , new_n448 );
  nand     g1449 ( new_n1835 , new_n466 , new_n1834 );
  nand g1450 ( new_n1836 , new_n1835 , new_n1835 );
  nand     g1451 ( new_n1837 , new_n1833 , new_n1836 );
  nand     g1452 ( new_n1838 , new_n1830 , new_n1837 );
  nand g1453 ( new_n1839 , new_n1838 , new_n1838 );
  nand     g1454 ( new_n1840 , new_n1808 , new_n1814 );
  nor      g1455 ( new_n1841 , new_n1839 , new_n1840 );
  nor      g1456 ( new_n1842 , new_n1828 , new_n1841 );
  nand     g1457 ( new_n1843 , new_n1821 , new_n1842 );
  nand     g1458 ( new_n1844 , new_n434 , new_n433 );
  nand     g1459 ( new_n1845 , new_n475 , new_n1451 );
  nor      g1460 ( new_n1846 , new_n1844 , new_n1845 );
  nand     g1461 ( new_n1847 , new_n1550 , new_n1846 );
  or       g1462 ( new_n1848 , new_n1843 , new_n1847 );
  nor      g1463 ( new_n1849 , pi105 , new_n526 );
  nand     g1464 ( new_n1850 , new_n431 , new_n1448 );
  nand     g1465 ( new_n1851 , new_n479 , pi255 );
  nand     g1466 ( new_n1852 , new_n549 , new_n1851 );
  nor      g1467 ( new_n1853 , new_n1850 , new_n1852 );
  nand     g1468 ( new_n1854 , new_n1849 , new_n1853 );
  nand g1469 ( new_n1855 , new_n482 , new_n482 );
  or       g1470 ( new_n1856 , new_n516 , new_n528 );
  nand     g1471 ( new_n1857 , new_n1855 , new_n1856 );
  nand     g1472 ( new_n1858 , new_n550 , new_n551 );
  nand     g1473 ( new_n1859 , new_n1857 , new_n1858 );
  nand     g1474 ( new_n1860 , new_n555 , new_n1859 );
  nand     g1475 ( new_n1861 , new_n1446 , new_n1860 );
  nand     g1476 ( new_n1862 , new_n1854 , new_n1861 );
  or       g1477 ( new_n1863 , new_n1848 , new_n1862 );
  and      g1478 ( new_n1864 , new_n1800 , new_n1863 );
  nand     g1479 ( new_n1865 , new_n1789 , new_n1864 );
  nand     g1480 ( new_n1866 , new_n1786 , new_n1865 );
  nand     g1481 ( new_n1867 , new_n671 , new_n889 );
  nand     g1482 ( new_n1868 , new_n877 , new_n1867 );
  nand     g1483 ( new_n1869 , new_n599 , new_n611 );
  nand     g1484 ( new_n1870 , new_n592 , new_n615 );
  nand     g1485 ( new_n1871 , new_n569 , new_n1870 );
  nand g1486 ( new_n1872 , new_n1871 , new_n1871 );
  and      g1487 ( new_n1873 , new_n1869 , new_n1872 );
  nand g1488 ( new_n1874 , pi009 , pi009 );
  nand     g1489 ( new_n1875 , new_n1874 , new_n621 );
  nor      g1490 ( new_n1876 , new_n625 , new_n1875 );
  nand g1491 ( new_n1877 , new_n1876 , new_n1876 );
  nand     g1492 ( new_n1878 , new_n630 , new_n1709 );
  nor      g1493 ( new_n1879 , new_n1877 , new_n1878 );
  nand     g1494 ( new_n1880 , new_n1498 , new_n1879 );
  nor      g1495 ( new_n1881 , new_n1873 , new_n1880 );
  nand     g1496 ( new_n1882 , new_n1868 , new_n1881 );
  nand     g1497 ( new_n1883 , new_n599 , new_n605 );
  nand     g1498 ( new_n1884 , new_n591 , new_n1883 );
  nand g1499 ( new_n1885 , new_n1884 , new_n1884 );
  nand     g1500 ( new_n1886 , new_n611 , new_n1721 );
  nor      g1501 ( new_n1887 , new_n1885 , new_n1886 );
  nor      g1502 ( new_n1888 , new_n1731 , new_n1887 );
  nand     g1503 ( new_n1889 , new_n1882 , new_n1888 );
  nand g1504 ( new_n1890 , new_n1889 , new_n1889 );
  nand g1505 ( new_n1891 , new_n496 , new_n496 );
  nand     g1506 ( new_n1892 , new_n1891 , new_n706 );
  nand     g1507 ( new_n1893 , new_n994 , new_n1004 );
  nand     g1508 ( new_n1894 , new_n1891 , new_n1893 );
  nand     g1509 ( new_n1895 , new_n1892 , new_n1894 );
  nand     g1510 ( new_n1896 , new_n486 , new_n1895 );
  nand     g1511 ( new_n1897 , new_n986 , pi169 );
  or       g1512 ( new_n1898 , new_n1707 , new_n1897 );
  nand g1513 ( new_n1899 , new_n1898 , new_n1898 );
  nor      g1514 ( new_n1900 , new_n1896 , new_n1899 );
  nor      g1515 ( new_n1901 , new_n1700 , new_n1900 );
  nand g1516 ( new_n1902 , new_n536 , new_n536 );
  nand     g1517 ( new_n1903 , pi007 , new_n504 );
  nand     g1518 ( new_n1904 , new_n1902 , new_n1903 );
  or       g1519 ( new_n1905 , new_n1901 , new_n1904 );
  nor      g1520 ( new_n1906 , new_n1890 , new_n1905 );
  nand     g1521 ( new_n1907 , new_n1866 , new_n1906 );
  nand     g1522 ( new_n1908 , new_n1694 , new_n1907 );
  nor      g1523 ( po004 , new_n1693 , new_n1908 );
  nand g1524 ( new_n1910 , new_n431 , new_n431 );
  or       g1525 ( new_n1911 , new_n993 , new_n563 );
  nand g1526 ( new_n1912 , new_n1561 , new_n1561 );
  nand     g1527 ( new_n1913 , new_n1306 , new_n1487 );
  nand     g1528 ( new_n1914 , new_n1648 , new_n1913 );
  nand     g1529 ( new_n1915 , new_n1912 , new_n1914 );
  nand     g1530 ( new_n1916 , new_n1237 , new_n1915 );
  nand g1531 ( new_n1917 , new_n1448 , new_n1448 );
  nand g1532 ( new_n1918 , new_n1858 , new_n1858 );
  nand g1533 ( new_n1919 , new_n540 , new_n540 );
  nor      g1534 ( new_n1920 , new_n520 , new_n1919 );
  nor      g1535 ( new_n1921 , new_n482 , new_n1920 );
  nor      g1536 ( new_n1922 , new_n1918 , new_n1921 );
  nand g1537 ( new_n1923 , new_n1204 , new_n1204 );
  nand     g1538 ( new_n1924 , new_n476 , new_n549 );
  nand g1539 ( new_n1925 , new_n1924 , new_n1924 );
  nand     g1540 ( new_n1926 , new_n1849 , new_n1925 );
  nor      g1541 ( new_n1927 , new_n1923 , new_n1926 );
  nor      g1542 ( new_n1928 , new_n1922 , new_n1927 );
  nor      g1543 ( new_n1929 , new_n1917 , new_n1928 );
  nand     g1544 ( new_n1930 , new_n1916 , new_n1929 );
  nor      g1545 ( new_n1931 , new_n1295 , new_n1930 );
  nor      g1546 ( new_n1932 , new_n1814 , new_n1826 );
  nor      g1547 ( new_n1933 , new_n396 , new_n1932 );
  nor      g1548 ( new_n1934 , new_n1457 , new_n1933 );
  or       g1549 ( new_n1935 , new_n413 , new_n1312 );
  nor      g1550 ( new_n1936 , new_n1934 , new_n1935 );
  and      g1551 ( new_n1937 , new_n1441 , new_n1936 );
  nand     g1552 ( new_n1938 , new_n412 , new_n1325 );
  nand     g1553 ( new_n1939 , new_n1409 , new_n1938 );
  nor      g1554 ( new_n1940 , new_n1233 , new_n1939 );
  nand     g1555 ( new_n1941 , new_n1455 , new_n1333 );
  nand g1556 ( new_n1942 , new_n1941 , new_n1941 );
  nand     g1557 ( new_n1943 , new_n1337 , new_n1942 );
  nor      g1558 ( new_n1944 , new_n1838 , new_n1943 );
  nand g1559 ( new_n1945 , new_n1944 , new_n1944 );
  nand     g1560 ( new_n1946 , new_n1936 , new_n1945 );
  nand     g1561 ( new_n1947 , new_n1940 , new_n1946 );
  nor      g1562 ( new_n1948 , new_n1937 , new_n1947 );
  nand     g1563 ( new_n1949 , new_n1237 , new_n1948 );
  nand     g1564 ( new_n1950 , new_n1931 , new_n1949 );
  nand     g1565 ( new_n1951 , new_n1911 , new_n1950 );
  nor      g1566 ( new_n1952 , new_n436 , new_n1951 );
  nor      g1567 ( new_n1953 , new_n1910 , new_n1952 );
  nand g1568 ( new_n1954 , new_n440 , new_n440 );
  nand     g1569 ( new_n1955 , pi030 , new_n1954 );
  nor      g1570 ( po005 , new_n1953 , new_n1955 );
  nand     g1571 ( new_n1957 , new_n1386 , new_n1347 );
  nand     g1572 ( new_n1958 , new_n1397 , new_n1957 );
  nand     g1573 ( new_n1959 , new_n1258 , new_n1958 );
  nand     g1574 ( new_n1960 , new_n1249 , new_n1959 );
  nor      g1575 ( po006 , new_n1241 , new_n1960 );
  nand     g1576 ( new_n1962 , pi189 , new_n595 );
  nor      g1577 ( new_n1963 , new_n585 , new_n1678 );
  nand g1578 ( new_n1964 , new_n991 , new_n991 );
  nand     g1579 ( new_n1965 , new_n641 , new_n1964 );
  nand     g1580 ( new_n1966 , new_n493 , new_n540 );
  nor      g1581 ( new_n1967 , new_n1892 , new_n1966 );
  nand     g1582 ( new_n1968 , new_n1965 , new_n1967 );
  or       g1583 ( new_n1969 , new_n1963 , new_n1968 );
  nor      g1584 ( new_n1970 , new_n528 , new_n1212 );
  nand     g1585 ( new_n1971 , new_n1434 , new_n1846 );
  nand     g1586 ( new_n1972 , new_n455 , new_n483 );
  nor      g1587 ( new_n1973 , new_n1971 , new_n1972 );
  nand g1588 ( new_n1974 , new_n1973 , new_n1973 );
  nor      g1589 ( new_n1975 , new_n1970 , new_n1974 );
  nand     g1590 ( new_n1976 , new_n1795 , new_n1975 );
  nand g1591 ( new_n1977 , new_n1976 , new_n1976 );
  nand     g1592 ( new_n1978 , new_n1969 , new_n1977 );
  nand     g1593 ( new_n1979 , new_n1800 , new_n1978 );
  nand g1594 ( new_n1980 , new_n1567 , new_n1567 );
  nand     g1595 ( new_n1981 , new_n1082 , new_n1980 );
  and      g1596 ( new_n1982 , new_n1635 , new_n1981 );
  nand     g1597 ( new_n1983 , new_n1979 , new_n1982 );
  nand g1598 ( new_n1984 , new_n1633 , new_n1633 );
  nand     g1599 ( new_n1985 , new_n1014 , new_n1087 );
  nor      g1600 ( new_n1986 , new_n1634 , new_n1985 );
  nor      g1601 ( new_n1987 , new_n1984 , new_n1986 );
  nand g1602 ( new_n1988 , new_n1987 , new_n1987 );
  nor      g1603 ( new_n1989 , new_n1201 , new_n1988 );
  nand     g1604 ( new_n1990 , new_n1983 , new_n1989 );
  nor      g1605 ( new_n1991 , new_n1201 , new_n1587 );
  nor      g1606 ( new_n1992 , new_n1193 , new_n1991 );
  nand g1607 ( new_n1993 , new_n1992 , new_n1992 );
  nand g1608 ( new_n1994 , new_n1360 , new_n1360 );
  nand     g1609 ( new_n1995 , new_n1994 , new_n1614 );
  nor      g1610 ( new_n1996 , new_n1993 , new_n1995 );
  nand     g1611 ( new_n1997 , new_n1990 , new_n1996 );
  nand     g1612 ( new_n1998 , new_n1617 , new_n1997 );
  nand     g1613 ( new_n1999 , new_n1962 , new_n1998 );
  nor      g1614 ( new_n2000 , pi129 , new_n1999 );
  nor      g1615 ( new_n2001 , pi057 , new_n2000 );
  nor      g1616 ( po007 , new_n577 , new_n2001 );
  nor      g1617 ( new_n2003 , new_n1588 , new_n1787 );
  nor      g1618 ( new_n2004 , new_n1503 , new_n2003 );
  and      g1619 ( new_n2005 , new_n1424 , new_n1704 );
  nand     g1620 ( new_n2006 , new_n978 , new_n2005 );
  nor      g1621 ( new_n2007 , new_n1626 , new_n2006 );
  nand g1622 ( new_n2008 , new_n2007 , new_n2007 );
  nor      g1623 ( new_n2009 , new_n2004 , new_n2008 );
  nand g1624 ( new_n2010 , new_n1879 , new_n1879 );
  nand     g1625 ( new_n2011 , new_n1874 , new_n1897 );
  nand g1626 ( new_n2012 , new_n2011 , new_n2011 );
  nand g1627 ( new_n2013 , new_n1717 , new_n1717 );
  nand     g1628 ( new_n2014 , new_n624 , new_n977 );
  nand     g1629 ( new_n2015 , new_n2013 , new_n2014 );
  nand     g1630 ( new_n2016 , new_n2012 , new_n2015 );
  nand     g1631 ( new_n2017 , new_n1706 , new_n2016 );
  nand g1632 ( new_n2018 , new_n2017 , new_n2017 );
  nand     g1633 ( new_n2019 , new_n2010 , new_n2018 );
  nand g1634 ( new_n2020 , new_n2019 , new_n2019 );
  nand     g1635 ( new_n2021 , new_n485 , new_n486 );
  nor      g1636 ( new_n2022 , new_n495 , new_n510 );
  nor      g1637 ( new_n2023 , new_n2021 , new_n2022 );
  nand g1638 ( new_n2024 , new_n2023 , new_n2023 );
  nand     g1639 ( new_n2025 , new_n525 , new_n538 );
  nor      g1640 ( new_n2026 , new_n2024 , new_n2025 );
  nand     g1641 ( new_n2027 , new_n692 , new_n494 );
  nand g1642 ( new_n2028 , new_n2027 , new_n2027 );
  nor      g1643 ( new_n2029 , pi106 , new_n702 );
  nand     g1644 ( new_n2030 , new_n696 , new_n2029 );
  nand     g1645 ( new_n2031 , new_n2028 , new_n2030 );
  nand g1646 ( new_n2032 , new_n2031 , new_n2031 );
  nand     g1647 ( new_n2033 , new_n2026 , new_n2032 );
  nor      g1648 ( new_n2034 , new_n2020 , new_n2033 );
  nand g1649 ( new_n2035 , new_n2034 , new_n2034 );
  nor      g1650 ( new_n2036 , new_n2009 , new_n2035 );
  nor      g1651 ( new_n2037 , new_n1540 , new_n1840 );
  nand     g1652 ( new_n2038 , new_n1428 , new_n470 );
  nand     g1653 ( new_n2039 , new_n1432 , new_n2038 );
  nand     g1654 ( new_n2040 , new_n2037 , new_n2039 );
  nand     g1655 ( new_n2041 , new_n1541 , new_n1828 );
  nand g1656 ( new_n2042 , new_n2041 , new_n2041 );
  nor      g1657 ( new_n2043 , new_n1544 , new_n2042 );
  nand     g1658 ( new_n2044 , new_n2040 , new_n2043 );
  nor      g1659 ( new_n2045 , pi183 , new_n507 );
  nand g1660 ( new_n2046 , new_n2045 , new_n2045 );
  nand     g1661 ( new_n2047 , new_n512 , new_n2046 );
  nand     g1662 ( new_n2048 , new_n525 , new_n532 );
  nand g1663 ( new_n2049 , new_n2048 , new_n2048 );
  nand     g1664 ( new_n2050 , new_n2047 , new_n2049 );
  nand g1665 ( new_n2051 , new_n2050 , new_n2050 );
  nand     g1666 ( new_n2052 , pi043 , new_n494 );
  nand     g1667 ( new_n2053 , new_n997 , new_n2052 );
  nand     g1668 ( new_n2054 , new_n2026 , new_n2053 );
  nand g1669 ( new_n2055 , new_n2054 , new_n2054 );
  nor      g1670 ( new_n2056 , new_n1971 , new_n2055 );
  nand     g1671 ( new_n2057 , new_n1861 , new_n2056 );
  nor      g1672 ( new_n2058 , new_n2051 , new_n2057 );
  nand g1673 ( new_n2059 , new_n2058 , new_n2058 );
  or       g1674 ( new_n2060 , new_n2044 , new_n2059 );
  nor      g1675 ( new_n2061 , new_n2036 , new_n2060 );
  nand g1676 ( new_n2062 , new_n2037 , new_n2037 );
  nor      g1677 ( new_n2063 , pi120 , pi178 );
  nand     g1678 ( new_n2064 , new_n543 , new_n2063 );
  nor      g1679 ( new_n2065 , new_n1850 , new_n2064 );
  nand g1680 ( new_n2066 , new_n2065 , new_n2065 );
  nand     g1681 ( new_n2067 , new_n523 , new_n1925 );
  nor      g1682 ( new_n2068 , new_n2066 , new_n2067 );
  nand     g1683 ( new_n2069 , new_n1811 , new_n2068 );
  nor      g1684 ( new_n2070 , new_n463 , new_n1298 );
  nand     g1685 ( new_n2071 , new_n1297 , new_n2070 );
  nand     g1686 ( new_n2072 , new_n2069 , new_n2071 );
  nand     g1687 ( new_n2073 , new_n468 , new_n2072 );
  nor      g1688 ( new_n2074 , new_n2062 , new_n2073 );
  nor      g1689 ( new_n2075 , new_n2044 , new_n2074 );
  nand     g1690 ( new_n2076 , new_n1390 , new_n1539 );
  or       g1691 ( new_n2077 , new_n2075 , new_n2076 );
  nor      g1692 ( new_n2078 , new_n2061 , new_n2077 );
  nand     g1693 ( new_n2079 , new_n1255 , new_n1400 );
  nand g1694 ( new_n2080 , new_n2079 , new_n2079 );
  nor      g1695 ( new_n2081 , new_n1024 , new_n1134 );
  nand     g1696 ( new_n2082 , new_n2080 , new_n2081 );
  nor      g1697 ( new_n2083 , new_n2078 , new_n2082 );
  nand g1698 ( new_n2084 , new_n1532 , new_n1532 );
  or       g1699 ( new_n2085 , new_n2084 , new_n1761 );
  nand     g1700 ( new_n2086 , new_n1752 , new_n2085 );
  nand     g1701 ( new_n2087 , new_n1147 , new_n2086 );
  nor      g1702 ( new_n2088 , new_n1020 , new_n1058 );
  nand     g1703 ( new_n2089 , new_n2087 , new_n2088 );
  nor      g1704 ( new_n2090 , new_n2083 , new_n2089 );
  nand     g1705 ( new_n2091 , pi084 , new_n1059 );
  nor      g1706 ( po008 , new_n2090 , new_n2091 );
  nand g1707 ( new_n2093 , new_n1141 , new_n1141 );
  nand g1708 ( new_n2094 , new_n1411 , new_n1411 );
  nor      g1709 ( new_n2095 , new_n2032 , new_n2053 );
  nand g1710 ( new_n2096 , new_n2095 , new_n2095 );
  nand g1711 ( new_n2097 , new_n1718 , new_n1718 );
  nor      g1712 ( new_n2098 , new_n1623 , new_n2097 );
  nor      g1713 ( new_n2099 , new_n2010 , new_n2098 );
  nor      g1714 ( new_n2100 , new_n998 , new_n2099 );
  nand     g1715 ( new_n2101 , new_n2018 , new_n2100 );
  nand     g1716 ( new_n2102 , new_n2096 , new_n2101 );
  nand     g1717 ( new_n2103 , new_n553 , new_n518 );
  nor      g1718 ( new_n2104 , new_n1470 , new_n2103 );
  nand g1719 ( new_n2105 , new_n2104 , new_n2104 );
  nor      g1720 ( new_n2106 , new_n2045 , new_n2105 );
  nand     g1721 ( new_n2107 , new_n2102 , new_n2106 );
  nand     g1722 ( new_n2108 , new_n1368 , new_n1614 );
  nand g1723 ( new_n2109 , new_n2108 , new_n2108 );
  nand     g1724 ( new_n2110 , new_n1746 , new_n2109 );
  nand     g1725 ( new_n2111 , new_n1868 , new_n2110 );
  nand     g1726 ( new_n2112 , new_n663 , new_n961 );
  nor      g1727 ( new_n2113 , new_n1675 , new_n2112 );
  nand     g1728 ( new_n2114 , new_n879 , new_n2113 );
  nand g1729 ( new_n2115 , new_n2114 , new_n2114 );
  nand     g1730 ( new_n2116 , new_n2111 , new_n2115 );
  nor      g1731 ( new_n2117 , new_n1722 , new_n1873 );
  nand     g1732 ( new_n2118 , new_n2116 , new_n2117 );
  nand g1733 ( new_n2119 , new_n1159 , new_n1159 );
  nor      g1734 ( new_n2120 , new_n2119 , new_n1175 );
  nand     g1735 ( new_n2121 , new_n1891 , new_n1876 );
  nor      g1736 ( new_n2122 , new_n703 , new_n2121 );
  nand g1737 ( new_n2123 , new_n2122 , new_n2122 );
  nor      g1738 ( new_n2124 , new_n2120 , new_n2123 );
  nand g1739 ( new_n2125 , new_n2124 , new_n2124 );
  nor      g1740 ( new_n2126 , new_n2118 , new_n2125 );
  nor      g1741 ( new_n2127 , new_n2107 , new_n2126 );
  nand g1742 ( new_n2128 , pi226 , pi226 );
  nand     g1743 ( new_n2129 , new_n1814 , new_n1829 );
  nand g1744 ( new_n2130 , new_n2129 , new_n2129 );
  nor      g1745 ( new_n2131 , new_n1826 , new_n2130 );
  nand g1746 ( new_n2132 , new_n2131 , new_n2131 );
  nand     g1747 ( new_n2133 , new_n393 , new_n2132 );
  nand     g1748 ( new_n2134 , new_n2128 , new_n2133 );
  nand g1749 ( new_n2135 , new_n2134 , new_n2134 );
  nor      g1750 ( new_n2136 , pi207 , new_n1805 );
  nand g1751 ( new_n2137 , new_n2136 , new_n2136 );
  nor      g1752 ( new_n2138 , pi126 , new_n427 );
  nor      g1753 ( new_n2139 , new_n2137 , new_n2138 );
  nor      g1754 ( new_n2140 , new_n1833 , new_n2139 );
  nand     g1755 ( new_n2141 , new_n2135 , new_n2140 );
  nand     g1756 ( new_n2142 , pi171 , new_n418 );
  nand     g1757 ( new_n2143 , new_n1316 , new_n2142 );
  nor      g1758 ( new_n2144 , new_n1458 , new_n2143 );
  nand g1759 ( new_n2145 , new_n2144 , new_n2144 );
  nand g1760 ( new_n2146 , pi159 , pi159 );
  nand     g1761 ( new_n2147 , new_n2146 , new_n441 );
  or       g1762 ( new_n2148 , new_n2145 , new_n2147 );
  or       g1763 ( new_n2149 , new_n2141 , new_n2148 );
  nand g1764 ( new_n2150 , new_n557 , new_n557 );
  nand     g1765 ( new_n2151 , new_n2150 , new_n562 );
  nand     g1766 ( new_n2152 , new_n437 , new_n2151 );
  nand     g1767 ( new_n2153 , new_n431 , new_n2152 );
  nand     g1768 ( new_n2154 , new_n479 , new_n1469 );
  nand g1769 ( new_n2155 , new_n2154 , new_n2154 );
  nand     g1770 ( new_n2156 , new_n524 , new_n2155 );
  nand     g1771 ( new_n2157 , new_n1853 , new_n2156 );
  nand     g1772 ( new_n2158 , new_n2153 , new_n2157 );
  nor      g1773 ( new_n2159 , new_n2149 , new_n2158 );
  nand g1774 ( new_n2160 , new_n2159 , new_n2159 );
  nand     g1775 ( new_n2161 , pi147 , new_n700 );
  nand     g1776 ( new_n2162 , new_n1002 , new_n2161 );
  nor      g1777 ( new_n2163 , new_n1703 , new_n2162 );
  nand     g1778 ( new_n2164 , new_n700 , new_n2012 );
  or       g1779 ( new_n2165 , new_n2013 , new_n2164 );
  nand g1780 ( new_n2166 , new_n2165 , new_n2165 );
  nand     g1781 ( new_n2167 , new_n513 , new_n512 );
  nor      g1782 ( new_n2168 , new_n2166 , new_n2167 );
  nand     g1783 ( new_n2169 , new_n2163 , new_n2168 );
  nor      g1784 ( new_n2170 , new_n2160 , new_n2169 );
  nand     g1785 ( new_n2171 , new_n2127 , new_n2170 );
  nand g1786 ( new_n2172 , new_n2106 , new_n2106 );
  nand     g1787 ( new_n2173 , new_n1891 , new_n695 );
  nand g1788 ( new_n2174 , new_n2173 , new_n2173 );
  nand     g1789 ( new_n2175 , new_n1697 , new_n1894 );
  nor      g1790 ( new_n2176 , new_n2174 , new_n2175 );
  nor      g1791 ( new_n2177 , new_n2021 , new_n2176 );
  nor      g1792 ( new_n2178 , new_n2172 , new_n2177 );
  nand     g1793 ( new_n2179 , new_n1860 , new_n2065 );
  nand     g1794 ( new_n2180 , new_n2049 , new_n2068 );
  nand     g1795 ( new_n2181 , new_n2179 , new_n2180 );
  nand g1796 ( new_n2182 , new_n2181 , new_n2181 );
  nand     g1797 ( new_n2183 , new_n535 , new_n2023 );
  nand     g1798 ( new_n2184 , new_n2106 , new_n2183 );
  nand     g1799 ( new_n2185 , new_n1818 , new_n2184 );
  nor      g1800 ( new_n2186 , new_n2182 , new_n2185 );
  nand g1801 ( new_n2187 , new_n2186 , new_n2186 );
  or       g1802 ( new_n2188 , new_n2178 , new_n2187 );
  nand     g1803 ( new_n2189 , new_n2159 , new_n2188 );
  nor      g1804 ( new_n2190 , pi128 , new_n1813 );
  nand     g1805 ( new_n2191 , new_n1836 , new_n2190 );
  nand     g1806 ( new_n2192 , new_n2135 , new_n2191 );
  nand     g1807 ( new_n2193 , pi094 , new_n2128 );
  nand     g1808 ( new_n2194 , new_n390 , new_n2193 );
  nor      g1809 ( new_n2195 , new_n1312 , new_n2194 );
  nand     g1810 ( new_n2196 , new_n2192 , new_n2195 );
  nand     g1811 ( new_n2197 , pi156 , new_n2146 );
  nand     g1812 ( new_n2198 , new_n423 , new_n2197 );
  nor      g1813 ( new_n2199 , new_n2137 , new_n2198 );
  nor      g1814 ( new_n2200 , new_n2141 , new_n2199 );
  nor      g1815 ( new_n2201 , new_n2196 , new_n2200 );
  nor      g1816 ( new_n2202 , new_n2143 , new_n2201 );
  nor      g1817 ( new_n2203 , new_n413 , new_n2202 );
  nand g1818 ( new_n2204 , new_n2203 , new_n2203 );
  nand     g1819 ( new_n2205 , new_n1938 , new_n2204 );
  and      g1820 ( new_n2206 , new_n2189 , new_n2205 );
  nor      g1821 ( new_n2207 , new_n1393 , new_n1402 );
  and      g1822 ( new_n2208 , new_n2206 , new_n2207 );
  nand     g1823 ( new_n2209 , new_n2171 , new_n2208 );
  nand     g1824 ( new_n2210 , new_n794 , new_n1733 );
  nand     g1825 ( new_n2211 , new_n1104 , new_n2210 );
  nand     g1826 ( new_n2212 , new_n1775 , new_n2211 );
  nand g1827 ( new_n2213 , new_n2212 , new_n2212 );
  or       g1828 ( new_n2214 , new_n849 , new_n858 );
  nor      g1829 ( new_n2215 , new_n2213 , new_n2214 );
  nor      g1830 ( new_n2216 , new_n1110 , new_n2215 );
  nand g1831 ( new_n2217 , new_n2216 , new_n2216 );
  nor      g1832 ( new_n2218 , new_n838 , new_n897 );
  nand     g1833 ( new_n2219 , new_n2115 , new_n2218 );
  nand g1834 ( new_n2220 , new_n2219 , new_n2219 );
  nand     g1835 ( new_n2221 , new_n2170 , new_n2220 );
  nor      g1836 ( new_n2222 , new_n2217 , new_n2221 );
  nor      g1837 ( new_n2223 , new_n2209 , new_n2222 );
  nor      g1838 ( new_n2224 , new_n2094 , new_n2223 );
  nor      g1839 ( new_n2225 , new_n2093 , new_n2224 );
  nand     g1840 ( new_n2226 , pi080 , new_n1125 );
  nor      g1841 ( po009 , new_n2225 , new_n2226 );
  nand g1842 ( new_n2228 , new_n1400 , new_n1400 );
  nor      g1843 ( new_n2229 , new_n2043 , new_n2076 );
  nor      g1844 ( new_n2230 , new_n2228 , new_n2229 );
  nand     g1845 ( new_n2231 , new_n1265 , new_n2230 );
  nand g1846 ( new_n2232 , new_n2231 , new_n2231 );
  nand     g1847 ( new_n2233 , new_n527 , new_n534 );
  nand     g1848 ( new_n2234 , new_n2155 , new_n2233 );
  nand g1849 ( new_n2235 , new_n2234 , new_n2234 );
  nor      g1850 ( new_n2236 , new_n2150 , new_n1844 );
  nand     g1851 ( new_n2237 , new_n2235 , new_n2236 );
  nor      g1852 ( new_n2238 , new_n1700 , new_n2237 );
  nand g1853 ( new_n2239 , new_n2237 , new_n2237 );
  nand g1854 ( new_n2240 , new_n1904 , new_n1904 );
  nand     g1855 ( new_n2241 , new_n1849 , new_n2240 );
  nand     g1856 ( new_n2242 , new_n2239 , new_n2241 );
  nand g1857 ( new_n2243 , new_n1853 , new_n1853 );
  nand     g1858 ( new_n2244 , new_n2243 , new_n2153 );
  nand     g1859 ( new_n2245 , new_n543 , new_n2244 );
  nor      g1860 ( new_n2246 , pi094 , pi128 );
  nand     g1861 ( new_n2247 , new_n390 , new_n2246 );
  nor      g1862 ( new_n2248 , new_n1805 , new_n2247 );
  nand     g1863 ( new_n2249 , new_n1818 , new_n2248 );
  nor      g1864 ( new_n2250 , new_n2245 , new_n2249 );
  nand     g1865 ( new_n2251 , new_n2242 , new_n2250 );
  nor      g1866 ( new_n2252 , new_n2238 , new_n2251 );
  nor      g1867 ( new_n2253 , new_n544 , new_n1445 );
  nand g1868 ( new_n2254 , new_n441 , new_n441 );
  nand     g1869 ( new_n2255 , new_n2254 , new_n543 );
  nand     g1870 ( new_n2256 , new_n1802 , new_n2255 );
  nor      g1871 ( new_n2257 , new_n2253 , new_n2256 );
  nor      g1872 ( new_n2258 , new_n1805 , new_n2257 );
  nor      g1873 ( new_n2259 , new_n453 , new_n2258 );
  nand g1874 ( new_n2260 , new_n2259 , new_n2259 );
  nor      g1875 ( new_n2261 , new_n461 , new_n1815 );
  nand     g1876 ( new_n2262 , new_n2260 , new_n2261 );
  nand     g1877 ( new_n2263 , new_n1944 , new_n2262 );
  nor      g1878 ( new_n2264 , new_n2252 , new_n2263 );
  nor      g1879 ( new_n2265 , new_n1934 , new_n2264 );
  nand g1880 ( new_n2266 , new_n2101 , new_n2101 );
  nand     g1881 ( new_n2267 , new_n1872 , new_n2266 );
  or       g1882 ( new_n2268 , new_n1755 , new_n2267 );
  or       g1883 ( new_n2269 , new_n2265 , new_n2268 );
  or       g1884 ( new_n2270 , new_n908 , new_n2269 );
  nand     g1885 ( new_n2271 , new_n2078 , new_n2270 );
  nand     g1886 ( new_n2272 , new_n2232 , new_n2271 );
  and      g1887 ( new_n2273 , new_n2084 , new_n2272 );
  nor      g1888 ( new_n2274 , new_n1761 , new_n2273 );
  nor      g1889 ( new_n2275 , new_n1043 , new_n1054 );
  nand g1890 ( new_n2276 , new_n2275 , new_n2275 );
  nor      g1891 ( new_n2277 , new_n2274 , new_n2276 );
  nand     g1892 ( new_n2278 , new_n1041 , pi157 );
  nand     g1893 ( new_n2279 , pi233 , new_n2278 );
  nor      g1894 ( po010 , new_n2277 , new_n2279 );
  nand g1895 ( new_n2281 , new_n1303 , new_n1303 );
  nor      g1896 ( new_n2282 , new_n2281 , new_n2206 );
  nand g1897 ( new_n2283 , new_n1940 , new_n1940 );
  nor      g1898 ( new_n2284 , new_n1480 , new_n2283 );
  nor      g1899 ( new_n2285 , new_n2093 , new_n1404 );
  or       g1900 ( new_n2286 , new_n1233 , new_n2285 );
  nand     g1901 ( new_n2287 , new_n807 , new_n871 );
  nor      g1902 ( new_n2288 , new_n1077 , new_n2287 );
  nand     g1903 ( new_n2289 , new_n2286 , new_n2288 );
  nor      g1904 ( new_n2290 , new_n2284 , new_n2289 );
  nor      g1905 ( new_n2291 , new_n790 , new_n1066 );
  nor      g1906 ( new_n2292 , new_n2287 , new_n2291 );
  nor      g1907 ( new_n2293 , new_n854 , new_n2292 );
  nor      g1908 ( new_n2294 , new_n906 , new_n1158 );
  nand     g1909 ( new_n2295 , new_n2293 , new_n2294 );
  nor      g1910 ( new_n2296 , new_n2290 , new_n2295 );
  nor      g1911 ( new_n2297 , new_n2125 , new_n2296 );
  or       g1912 ( new_n2298 , new_n496 , new_n992 );
  nor      g1913 ( new_n2299 , new_n501 , new_n2175 );
  nand     g1914 ( new_n2300 , new_n2298 , new_n2299 );
  nor      g1915 ( new_n2301 , new_n2297 , new_n2300 );
  nand g1916 ( new_n2302 , new_n2301 , new_n2301 );
  nand     g1917 ( new_n2303 , new_n1460 , new_n2170 );
  nor      g1918 ( new_n2304 , new_n2302 , new_n2303 );
  nor      g1919 ( new_n2305 , new_n2282 , new_n2304 );
  nor      g1920 ( po011 , new_n1405 , new_n2305 );
  nor      g1921 ( new_n2307 , new_n1536 , new_n1550 );
  nor      g1922 ( new_n2308 , new_n1763 , new_n2307 );
  nand g1923 ( new_n2309 , new_n2308 , new_n2308 );
  nand g1924 ( new_n2310 , new_n2179 , new_n2179 );
  nand     g1925 ( new_n2311 , pi016 , new_n1816 );
  nand     g1926 ( new_n2312 , new_n2131 , new_n2311 );
  nand g1927 ( new_n2313 , new_n2312 , new_n2312 );
  nand     g1928 ( new_n2314 , new_n1824 , new_n2313 );
  nor      g1929 ( new_n2315 , new_n2310 , new_n2314 );
  nand     g1930 ( new_n2316 , new_n2259 , new_n2315 );
  nor      g1931 ( new_n2317 , new_n2309 , new_n2316 );
  nand g1932 ( new_n2318 , new_n2317 , new_n2317 );
  nor      g1933 ( new_n2319 , new_n2047 , new_n2318 );
  nand g1934 ( new_n2320 , new_n2319 , new_n2319 );
  nor      g1935 ( new_n2321 , new_n2095 , new_n2183 );
  nor      g1936 ( new_n2322 , new_n2320 , new_n2321 );
  nand     g1937 ( new_n2323 , new_n2180 , new_n2317 );
  nand g1938 ( new_n2324 , new_n2323 , new_n2323 );
  nand g1939 ( new_n2325 , new_n1756 , new_n1756 );
  nand g1940 ( new_n2326 , new_n2196 , new_n2196 );
  nand     g1941 ( new_n2327 , new_n1431 , new_n2135 );
  nand     g1942 ( new_n2328 , new_n2326 , new_n2327 );
  nand     g1943 ( new_n2329 , new_n2144 , new_n2328 );
  nand     g1944 ( new_n2330 , new_n1557 , new_n2329 );
  nand     g1945 ( new_n2331 , new_n2308 , new_n2330 );
  nand     g1946 ( new_n2332 , new_n2325 , new_n2331 );
  nor      g1947 ( new_n2333 , new_n2324 , new_n2332 );
  nand g1948 ( new_n2334 , new_n2333 , new_n2333 );
  nor      g1949 ( new_n2335 , new_n2322 , new_n2334 );
  nand     g1950 ( new_n2336 , new_n2266 , new_n2319 );
  nor      g1951 ( new_n2337 , new_n1881 , new_n2336 );
  nor      g1952 ( new_n2338 , new_n1748 , new_n2337 );
  nand     g1953 ( new_n2339 , new_n2335 , new_n2338 );
  nand     g1954 ( new_n2340 , new_n1769 , new_n1781 );
  nor      g1955 ( new_n2341 , new_n1779 , new_n2340 );
  nand     g1956 ( new_n2342 , new_n2339 , new_n2341 );
  and      g1957 ( new_n2343 , new_n1868 , new_n2342 );
  nand     g1958 ( new_n2344 , pi108 , new_n604 );
  nor      g1959 ( po012 , new_n2343 , new_n2344 );
  nand g1960 ( new_n2346 , new_n2071 , new_n2071 );
  nor      g1961 ( new_n2347 , new_n1931 , new_n2346 );
  nand     g1962 ( new_n2348 , new_n471 , new_n1334 );
  nor      g1963 ( new_n2349 , new_n566 , new_n2348 );
  nand g1964 ( new_n2350 , new_n2349 , new_n2349 );
  nand g1965 ( new_n2351 , new_n1808 , new_n1808 );
  nor      g1966 ( new_n2352 , pi117 , new_n2351 );
  nand     g1967 ( new_n2353 , new_n2350 , new_n2352 );
  nor      g1968 ( new_n2354 , new_n2347 , new_n2353 );
  nor      g1969 ( new_n2355 , new_n1843 , new_n2354 );
  nor      g1970 ( new_n2356 , new_n1540 , new_n2355 );
  nand     g1971 ( new_n2357 , pi218 , new_n1543 );
  nor      g1972 ( po013 , new_n2356 , new_n2357 );
  nand     g1973 ( new_n2359 , new_n619 , new_n638 );
  nand     g1974 ( new_n2360 , new_n1964 , new_n2359 );
  nand     g1975 ( new_n2361 , new_n1208 , new_n2360 );
  nand     g1976 ( new_n2362 , new_n1475 , new_n2361 );
  nand     g1977 ( new_n2363 , new_n931 , new_n1114 );
  and      g1978 ( new_n2364 , new_n1380 , new_n2363 );
  nor      g1979 ( new_n2365 , new_n929 , new_n2364 );
  nor      g1980 ( new_n2366 , new_n1374 , new_n2365 );
  nor      g1981 ( new_n2367 , new_n709 , new_n2366 );
  or       g1982 ( new_n2368 , new_n2362 , new_n2367 );
  nand     g1983 ( new_n2369 , new_n1493 , new_n2368 );
  nand     g1984 ( new_n2370 , new_n1530 , new_n2369 );
  nand g1985 ( new_n2371 , new_n2370 , new_n2370 );
  or       g1986 ( new_n2372 , new_n947 , new_n2371 );
  nand     g1987 ( new_n2373 , new_n934 , new_n2372 );
  nor      g1988 ( po014 , new_n932 , new_n2373 );
  nand     g1989 ( new_n2375 , new_n1363 , new_n1993 );
  nand     g1990 ( new_n2376 , new_n569 , new_n593 );
  nor      g1991 ( new_n2377 , new_n2108 , new_n2376 );
  nand     g1992 ( new_n2378 , new_n2375 , new_n2377 );
  nand g1993 ( new_n2379 , new_n2378 , new_n2378 );
  nand     g1994 ( new_n2380 , new_n1239 , new_n1912 );
  nand     g1995 ( new_n2381 , new_n1635 , new_n2380 );
  nor      g1996 ( new_n2382 , new_n1980 , new_n2381 );
  nand     g1997 ( new_n2383 , new_n2379 , new_n2382 );
  nand g1998 ( new_n2384 , new_n2383 , new_n2383 );
  nand     g1999 ( new_n2385 , new_n1915 , new_n2384 );
  nand     g2000 ( new_n2386 , new_n1083 , new_n1635 );
  nand     g2001 ( new_n2387 , new_n1200 , new_n2386 );
  nor      g2002 ( new_n2388 , new_n1984 , new_n2387 );
  nand     g2003 ( new_n2389 , new_n1371 , new_n2388 );
  nand     g2004 ( new_n2390 , new_n2379 , new_n2389 );
  nand     g2005 ( new_n2391 , pi195 , new_n1614 );
  nand     g2006 ( new_n2392 , new_n1610 , new_n2391 );
  nand     g2007 ( new_n2393 , new_n1872 , new_n2392 );
  nand     g2008 ( new_n2394 , new_n1881 , new_n2393 );
  nand     g2009 ( new_n2395 , new_n702 , new_n2028 );
  nor      g2010 ( new_n2396 , new_n2394 , new_n2395 );
  nand     g2011 ( new_n2397 , new_n2390 , new_n2396 );
  nand g2012 ( new_n2398 , new_n2397 , new_n2397 );
  nand     g2013 ( new_n2399 , new_n2385 , new_n2398 );
  nor      g2014 ( new_n2400 , new_n420 , new_n1328 );
  nand     g2015 ( new_n2401 , new_n1646 , new_n2400 );
  nor      g2016 ( new_n2402 , new_n2383 , new_n2401 );
  nor      g2017 ( new_n2403 , new_n2399 , new_n2402 );
  nor      g2018 ( new_n2404 , new_n2107 , new_n2403 );
  nor      g2019 ( new_n2405 , new_n2187 , new_n2404 );
  nand     g2020 ( new_n2406 , new_n2262 , new_n2313 );
  nor      g2021 ( new_n2407 , new_n2405 , new_n2406 );
  nor      g2022 ( new_n2408 , new_n2351 , new_n2407 );
  nand     g2023 ( new_n2409 , pi022 , new_n1822 );
  nor      g2024 ( po015 , new_n2408 , new_n2409 );
  nand g2025 ( new_n2411 , new_n815 , new_n815 );
  nand     g2026 ( new_n2412 , new_n1106 , new_n1734 );
  nand     g2027 ( new_n2413 , new_n1778 , new_n2412 );
  nand g2028 ( new_n2414 , new_n2413 , new_n2413 );
  or       g2029 ( new_n2415 , new_n1657 , new_n1659 );
  nor      g2030 ( new_n2416 , new_n2415 , new_n2127 );
  or       g2031 ( new_n2417 , new_n1684 , new_n2416 );
  nand     g2032 ( new_n2418 , new_n1106 , new_n2417 );
  nand     g2033 ( new_n2419 , new_n2414 , new_n2418 );
  nor      g2034 ( new_n2420 , new_n2411 , new_n2419 );
  nor      g2035 ( new_n2421 , pi135 , new_n2420 );
  nor      g2036 ( po016 , new_n819 , new_n2421 );
  nand g2037 ( new_n2423 , new_n1929 , new_n1929 );
  nand g2038 ( new_n2424 , new_n2126 , new_n2126 );
  nor      g2039 ( new_n2425 , new_n1776 , new_n2331 );
  nor      g2040 ( new_n2426 , new_n2216 , new_n2425 );
  nor      g2041 ( new_n2427 , new_n2219 , new_n2426 );
  nor      g2042 ( new_n2428 , new_n2424 , new_n2427 );
  nor      g2043 ( new_n2429 , new_n2107 , new_n2428 );
  nor      g2044 ( new_n2430 , new_n2423 , new_n2429 );
  nor      g2045 ( new_n2431 , new_n1450 , new_n2430 );
  nor      g2046 ( new_n2432 , new_n432 , new_n2431 );
  nor      g2047 ( new_n2433 , new_n442 , new_n2432 );
  nand g2048 ( new_n2434 , new_n2433 , new_n2433 );
  nor      g2049 ( new_n2435 , pi159 , new_n2434 );
  nor      g2050 ( new_n2436 , pi098 , new_n2435 );
  nor      g2051 ( po017 , new_n425 , new_n2436 );
  nand g2052 ( new_n2438 , new_n2407 , new_n2407 );
  nand     g2053 ( new_n2439 , new_n397 , new_n2438 );
  nand     g2054 ( new_n2440 , new_n1456 , new_n2439 );
  nor      g2055 ( new_n2441 , pi081 , new_n2440 );
  nor      g2056 ( new_n2442 , pi103 , new_n2441 );
  nor      g2057 ( po018 , new_n1308 , new_n2442 );
  nand g2058 ( new_n2444 , new_n2161 , new_n2161 );
  nand g2059 ( new_n2445 , new_n2177 , new_n2177 );
  or       g2060 ( new_n2446 , new_n1848 , new_n2172 );
  nor      g2061 ( new_n2447 , new_n1784 , new_n2446 );
  and      g2062 ( new_n2448 , new_n2445 , new_n2447 );
  nand g2063 ( new_n2449 , new_n2256 , new_n2256 );
  nand     g2064 ( new_n2450 , new_n2245 , new_n2449 );
  nor      g2065 ( new_n2451 , new_n1935 , new_n2249 );
  nand     g2066 ( new_n2452 , new_n2450 , new_n2451 );
  nor      g2067 ( new_n2453 , new_n2349 , new_n2452 );
  nor      g2068 ( new_n2454 , new_n1947 , new_n2453 );
  nor      g2069 ( new_n2455 , new_n2289 , new_n2454 );
  nor      g2070 ( new_n2456 , new_n2295 , new_n2455 );
  or       g2071 ( new_n2457 , new_n2118 , new_n2456 );
  or       g2072 ( new_n2458 , new_n2448 , new_n2457 );
  and      g2073 ( new_n2459 , new_n1728 , new_n2458 );
  nor      g2074 ( new_n2460 , new_n2164 , new_n2459 );
  or       g2075 ( new_n2461 , new_n2444 , new_n2460 );
  nor      g2076 ( new_n2462 , pi070 , new_n2461 );
  nor      g2077 ( new_n2463 , pi074 , new_n2462 );
  nor      g2078 ( po019 , new_n682 , new_n2463 );
  nor      g2079 ( new_n2465 , new_n1627 , new_n2010 );
  nand     g2080 ( new_n2466 , pi147 , new_n2016 );
  nor      g2081 ( po020 , new_n2465 , new_n2466 );
  nand     g2082 ( new_n2468 , new_n395 , new_n2438 );
  nor      g2083 ( new_n2469 , pi200 , new_n2468 );
  nand     g2084 ( new_n2470 , pi171 , new_n404 );
  nor      g2085 ( po021 , new_n2469 , new_n2470 );
  nand g2086 ( new_n2472 , pi070 , pi070 );
  nor      g2087 ( po022 , new_n2472 , new_n2461 );
  nor      g2088 ( new_n2474 , new_n1607 , new_n2008 );
  or       g2089 ( new_n2475 , new_n2035 , new_n2474 );
  nor      g2090 ( new_n2476 , new_n1433 , new_n2059 );
  and      g2091 ( new_n2477 , new_n2475 , new_n2476 );
  nor      g2092 ( new_n2478 , new_n2251 , new_n2477 );
  nor      g2093 ( new_n2479 , new_n2265 , new_n2478 );
  nor      g2094 ( new_n2480 , new_n1312 , new_n2479 );
  nand     g2095 ( new_n2481 , new_n416 , pi022 );
  nand     g2096 ( new_n2482 , pi075 , new_n2481 );
  nor      g2097 ( po023 , new_n2480 , new_n2482 );
  nand     g2098 ( new_n2484 , new_n1012 , new_n1795 );
  nor      g2099 ( new_n2485 , new_n1293 , new_n1511 );
  nand     g2100 ( new_n2486 , new_n2484 , new_n2485 );
  nand     g2101 ( new_n2487 , new_n1506 , new_n2486 );
  nor      g2102 ( new_n2488 , pi170 , new_n2487 );
  nor      g2103 ( new_n2489 , pi023 , new_n2488 );
  nor      g2104 ( po024 , new_n944 , new_n2489 );
  nor      g2105 ( new_n2491 , new_n2125 , new_n2456 );
  nor      g2106 ( new_n2492 , new_n2300 , new_n2491 );
  nor      g2107 ( new_n2493 , new_n492 , new_n2492 );
  nand     g2108 ( new_n2494 , pi066 , new_n505 );
  nor      g2109 ( po025 , new_n2493 , new_n2494 );
  nand g2110 ( new_n2496 , new_n853 , new_n853 );
  nor      g2111 ( new_n2497 , new_n2496 , new_n928 );
  nor      g2112 ( new_n2498 , new_n679 , new_n2497 );
  nand     g2113 ( new_n2499 , new_n906 , new_n1172 );
  nand g2114 ( new_n2500 , new_n2499 , new_n2499 );
  nor      g2115 ( new_n2501 , new_n1678 , new_n2500 );
  nand g2116 ( new_n2502 , new_n2501 , new_n2501 );
  nor      g2117 ( new_n2503 , new_n2498 , new_n2502 );
  nor      g2118 ( new_n2504 , new_n1968 , new_n2503 );
  or       g2119 ( new_n2505 , new_n728 , new_n768 );
  nor      g2120 ( new_n2506 , new_n2502 , new_n2505 );
  nand     g2121 ( new_n2507 , new_n1988 , new_n2506 );
  nand     g2122 ( new_n2508 , new_n2504 , new_n2507 );
  nand     g2123 ( new_n2509 , new_n1977 , new_n2508 );
  nand     g2124 ( new_n2510 , new_n1800 , new_n2509 );
  nand     g2125 ( new_n2511 , new_n1981 , new_n2510 );
  and      g2126 ( new_n2512 , new_n1013 , new_n2511 );
  nand     g2127 ( new_n2513 , pi053 , new_n1090 );
  nor      g2128 ( po026 , new_n2512 , new_n2513 );
  nand     g2129 ( new_n2515 , new_n1144 , new_n1380 );
  nand g2130 ( new_n2516 , new_n2515 , new_n2515 );
  and      g2131 ( new_n2517 , new_n2283 , new_n2286 );
  or       g2132 ( new_n2518 , new_n1057 , new_n2517 );
  nor      g2133 ( new_n2519 , new_n1375 , new_n2518 );
  nor      g2134 ( new_n2520 , new_n2516 , new_n2519 );
  nand g2135 ( new_n2521 , pi148 , pi148 );
  nand g2136 ( new_n2522 , new_n745 , new_n745 );
  nand     g2137 ( new_n2523 , new_n2521 , new_n2522 );
  nor      g2138 ( new_n2524 , new_n2520 , new_n2523 );
  nor      g2139 ( new_n2525 , new_n909 , new_n1800 );
  nand     g2140 ( new_n2526 , new_n2524 , new_n2525 );
  nand     g2141 ( new_n2527 , new_n926 , new_n2526 );
  nand     g2142 ( new_n2528 , new_n2506 , new_n2527 );
  nand     g2143 ( new_n2529 , new_n2504 , new_n2528 );
  nand g2144 ( new_n2530 , new_n477 , new_n477 );
  nor      g2145 ( new_n2531 , new_n2530 , new_n1970 );
  nand     g2146 ( new_n2532 , new_n2529 , new_n2531 );
  nor      g2147 ( new_n2533 , pi251 , new_n2532 );
  nor      g2148 ( new_n2534 , pi242 , new_n2533 );
  nor      g2149 ( new_n2535 , pi125 , new_n2534 );
  nor      g2150 ( new_n2536 , pi210 , new_n2535 );
  nor      g2151 ( po027 , new_n553 , new_n2536 );
  nand g2152 ( new_n2538 , new_n1415 , new_n1415 );
  nand g2153 ( new_n2539 , new_n2215 , new_n2215 );
  nand     g2154 ( new_n2540 , new_n1107 , new_n2539 );
  nor      g2155 ( new_n2541 , new_n2221 , new_n2540 );
  nor      g2156 ( new_n2542 , new_n2209 , new_n2541 );
  nor      g2157 ( new_n2543 , new_n2538 , new_n2542 );
  nand     g2158 ( new_n2544 , new_n921 , new_n2515 );
  nor      g2159 ( new_n2545 , new_n2543 , new_n2544 );
  nor      g2160 ( new_n2546 , new_n1349 , new_n2545 );
  nor      g2161 ( new_n2547 , new_n776 , new_n2546 );
  nor      g2162 ( new_n2548 , new_n785 , new_n2547 );
  or       g2163 ( new_n2549 , new_n792 , new_n2548 );
  nand     g2164 ( new_n2550 , new_n794 , new_n2549 );
  nor      g2165 ( po028 , new_n1570 , new_n2550 );
  nor      g2166 ( new_n2552 , pi206 , new_n1960 );
  nor      g2167 ( new_n2553 , pi018 , new_n2552 );
  nor      g2168 ( new_n2554 , pi020 , new_n2553 );
  or       g2169 ( new_n2555 , pi212 , new_n2554 );
  and      g2170 ( po029 , pi127 , new_n2555 );
  nor      g2171 ( new_n2557 , new_n989 , new_n2460 );
  nor      g2172 ( new_n2558 , new_n707 , new_n2557 );
  nand     g2173 ( new_n2559 , pi043 , new_n1004 );
  nor      g2174 ( po030 , new_n2558 , new_n2559 );
  nor      g2175 ( po031 , new_n1037 , new_n2487 );
  nand     g2176 ( new_n2562 , new_n1217 , new_n1493 );
  nand     g2177 ( new_n2563 , new_n1656 , new_n2562 );
  nand     g2178 ( new_n2564 , new_n1658 , new_n2563 );
  nand     g2179 ( new_n2565 , new_n1637 , new_n2564 );
  nand     g2180 ( new_n2566 , pi112 , new_n1583 );
  nor      g2181 ( po032 , new_n2565 , new_n2566 );
  nor      g2182 ( new_n2568 , pi209 , new_n2548 );
  nor      g2183 ( po033 , new_n793 , new_n2568 );
  nand g2184 ( new_n2570 , new_n1958 , new_n1958 );
  nor      g2185 ( new_n2571 , pi032 , new_n2570 );
  nor      g2186 ( po034 , new_n1248 , new_n2571 );
  nand g2187 ( new_n2573 , new_n2113 , new_n2113 );
  nand     g2188 ( new_n2574 , new_n1614 , new_n1846 );
  nor      g2189 ( new_n2575 , new_n1792 , new_n2574 );
  nand     g2190 ( new_n2576 , new_n1358 , new_n2575 );
  nor      g2191 ( new_n2577 , new_n2573 , new_n2576 );
  nand     g2192 ( new_n2578 , new_n1436 , new_n1942 );
  nand     g2193 ( new_n2579 , new_n1791 , new_n2005 );
  nor      g2194 ( new_n2580 , new_n2105 , new_n2579 );
  nand g2195 ( new_n2581 , pi244 , pi244 );
  nor      g2196 ( new_n2582 , pi055 , pi110 );
  nand     g2197 ( new_n2583 , new_n2581 , new_n2582 );
  nor      g2198 ( new_n2584 , new_n713 , new_n758 );
  nand     g2199 ( new_n2585 , new_n2522 , new_n2584 );
  or       g2200 ( new_n2586 , new_n2583 , new_n2585 );
  nand     g2201 ( new_n2587 , new_n1002 , new_n1464 );
  or       g2202 ( new_n2588 , new_n2586 , new_n2587 );
  or       g2203 ( new_n2589 , new_n1634 , new_n1652 );
  nor      g2204 ( new_n2590 , new_n2588 , new_n2589 );
  nand     g2205 ( new_n2591 , new_n2580 , new_n2590 );
  nor      g2206 ( new_n2592 , new_n2578 , new_n2591 );
  nand     g2207 ( po035 , new_n2577 , new_n2592 );
  nor      g2208 ( new_n2594 , new_n2183 , new_n2492 );
  nand     g2209 ( new_n2595 , pi041 , new_n2046 );
  nor      g2210 ( po036 , new_n2594 , new_n2595 );
  nor      g2211 ( new_n2597 , new_n2362 , new_n2398 );
  nor      g2212 ( new_n2598 , new_n1492 , new_n2597 );
  nor      g2213 ( new_n2599 , new_n1531 , new_n2598 );
  nor      g2214 ( new_n2600 , new_n958 , new_n2599 );
  nand     g2215 ( new_n2601 , pi052 , new_n1565 );
  nor      g2216 ( po037 , new_n2600 , new_n2601 );
  nand g2217 ( new_n2603 , new_n1888 , new_n1888 );
  nor      g2218 ( new_n2604 , new_n642 , new_n2603 );
  nor      g2219 ( new_n2605 , new_n1901 , new_n2241 );
  nand g2220 ( new_n2606 , new_n2605 , new_n2605 );
  nor      g2221 ( new_n2607 , new_n2604 , new_n2606 );
  nand     g2222 ( new_n2608 , new_n2239 , new_n2449 );
  nor      g2223 ( new_n2609 , new_n2607 , new_n2608 );
  nor      g2224 ( new_n2610 , new_n2452 , new_n2609 );
  nor      g2225 ( new_n2611 , new_n1947 , new_n2610 );
  nor      g2226 ( new_n2612 , new_n2289 , new_n2611 );
  and      g2227 ( new_n2613 , new_n901 , new_n898 );
  nand     g2228 ( new_n2614 , new_n2293 , new_n2613 );
  nor      g2229 ( new_n2615 , new_n2612 , new_n2614 );
  nand     g2230 ( new_n2616 , new_n901 , pi247 );
  nand     g2231 ( new_n2617 , new_n646 , new_n2616 );
  nor      g2232 ( new_n2618 , new_n2615 , new_n2617 );
  nor      g2233 ( new_n2619 , pi071 , new_n2618 );
  nor      g2234 ( new_n2620 , pi062 , new_n2619 );
  nor      g2235 ( po038 , new_n643 , new_n2620 );
  nand g2236 ( new_n2622 , new_n1712 , new_n1712 );
  nor      g2237 ( new_n2623 , new_n1630 , new_n2622 );
  nor      g2238 ( new_n2624 , pi017 , new_n2623 );
  nor      g2239 ( po039 , new_n973 , new_n2624 );
  nor      g2240 ( new_n2626 , new_n900 , new_n2343 );
  nor      g2241 ( new_n2627 , pi164 , new_n2626 );
  nor      g2242 ( po040 , new_n582 , new_n2627 );
  nor      g2243 ( new_n2629 , new_n758 , new_n2565 );
  nor      g2244 ( new_n2630 , new_n1154 , new_n2629 );
  nand     g2245 ( new_n2631 , pi035 , new_n711 );
  nor      g2246 ( po041 , new_n2630 , new_n2631 );
  nor      g2247 ( new_n2633 , new_n1896 , new_n2251 );
  nor      g2248 ( new_n2634 , new_n2265 , new_n2633 );
  nor      g2249 ( new_n2635 , new_n1935 , new_n2634 );
  nor      g2250 ( new_n2636 , new_n1939 , new_n2635 );
  nor      g2251 ( new_n2637 , new_n1915 , new_n2636 );
  or       g2252 ( new_n2638 , new_n1236 , new_n2637 );
  and      g2253 ( new_n2639 , new_n1757 , new_n2638 );
  nor      g2254 ( new_n2640 , new_n908 , new_n2639 );
  nor      g2255 ( new_n2641 , new_n1176 , new_n2640 );
  nor      g2256 ( new_n2642 , new_n1160 , new_n2641 );
  nor      g2257 ( new_n2643 , new_n627 , new_n2642 );
  nand     g2258 ( new_n2644 , pi037 , new_n984 );
  nor      g2259 ( po042 , new_n2643 , new_n2644 );
  nor      g2260 ( new_n2646 , new_n1588 , new_n2565 );
  nor      g2261 ( new_n2647 , new_n1199 , new_n2646 );
  nand     g2262 ( new_n2648 , pi132 , new_n1188 );
  nor      g2263 ( po043 , new_n2647 , new_n2648 );
  and      g2264 ( po044 , pi083 , new_n1686 );
  nand g2265 ( new_n2651 , new_n1854 , new_n1854 );
  nand     g2266 ( new_n2652 , new_n1213 , new_n2651 );
  nand     g2267 ( new_n2653 , new_n1853 , new_n2234 );
  nand     g2268 ( new_n2654 , new_n2153 , new_n2653 );
  nand g2269 ( new_n2655 , new_n2654 , new_n2654 );
  nor      g2270 ( new_n2656 , new_n2254 , new_n2578 );
  nand     g2271 ( new_n2657 , new_n2655 , new_n2656 );
  nand g2272 ( new_n2658 , new_n2657 , new_n2657 );
  nand     g2273 ( new_n2659 , new_n2652 , new_n2658 );
  nand     g2274 ( new_n2660 , new_n2203 , new_n2659 );
  nand g2275 ( new_n2661 , new_n2660 , new_n2660 );
  nand     g2276 ( new_n2662 , new_n2285 , new_n2661 );
  nand     g2277 ( new_n2663 , new_n641 , new_n1730 );
  nor      g2278 ( new_n2664 , new_n2265 , new_n2663 );
  nor      g2279 ( new_n2665 , new_n2662 , new_n2664 );
  nor      g2280 ( new_n2666 , new_n2518 , new_n2665 );
  nand     g2281 ( new_n2667 , new_n874 , new_n2217 );
  nor      g2282 ( new_n2668 , new_n2666 , new_n2667 );
  nor      g2283 ( new_n2669 , new_n908 , new_n2668 );
  nor      g2284 ( new_n2670 , new_n587 , new_n2669 );
  nor      g2285 ( new_n2671 , new_n579 , new_n2670 );
  nor      g2286 ( new_n2672 , pi102 , new_n2671 );
  nor      g2287 ( po045 , new_n575 , new_n2672 );
  or       g2288 ( new_n2674 , new_n1142 , new_n1385 );
  and      g2289 ( new_n2675 , new_n431 , new_n562 );
  or       g2290 ( new_n2676 , new_n446 , new_n2675 );
  or       g2291 ( new_n2677 , new_n2149 , new_n2676 );
  and      g2292 ( new_n2678 , new_n2207 , new_n2677 );
  nand     g2293 ( new_n2679 , new_n2205 , new_n2678 );
  nor      g2294 ( new_n2680 , new_n2674 , new_n2679 );
  nor      g2295 ( new_n2681 , new_n2603 , new_n2680 );
  nand     g2296 ( new_n2682 , new_n1417 , new_n2681 );
  nand g2297 ( new_n2683 , new_n2682 , new_n2682 );
  nand     g2298 ( new_n2684 , new_n1925 , new_n2607 );
  nor      g2299 ( new_n2685 , new_n2683 , new_n2684 );
  nor      g2300 ( new_n2686 , new_n1922 , new_n2685 );
  nor      g2301 ( new_n2687 , pi214 , new_n2686 );
  nor      g2302 ( new_n2688 , pi214 , new_n473 );
  nor      g2303 ( new_n2689 , new_n472 , new_n2688 );
  nand     g2304 ( new_n2690 , new_n1861 , new_n2689 );
  nor      g2305 ( po046 , new_n2687 , new_n2690 );
  nor      g2306 ( new_n2692 , new_n1028 , new_n2090 );
  nor      g2307 ( new_n2693 , new_n1376 , new_n2692 );
  nand     g2308 ( new_n2694 , pi048 , new_n731 );
  nor      g2309 ( po047 , new_n2693 , new_n2694 );
  nor      g2310 ( po048 , new_n1242 , new_n2553 );
  nand     g2311 ( new_n2697 , new_n637 , new_n981 );
  nor      g2312 ( new_n2698 , pi240 , new_n1877 );
  nand     g2313 ( new_n2699 , new_n2697 , new_n2698 );
  and      g2314 ( new_n2700 , new_n2170 , new_n2699 );
  nor      g2315 ( new_n2701 , new_n2674 , new_n2700 );
  nand     g2316 ( new_n2702 , new_n2208 , new_n2701 );
  nand     g2317 ( new_n2703 , new_n1417 , new_n2702 );
  nand     g2318 ( new_n2704 , new_n617 , new_n2703 );
  nand     g2319 ( new_n2705 , new_n618 , new_n2704 );
  nand     g2320 ( new_n2706 , new_n1496 , new_n2705 );
  nand     g2321 ( new_n2707 , new_n1718 , new_n2706 );
  nor      g2322 ( po049 , new_n571 , new_n2707 );
  nor      g2323 ( po050 , new_n1314 , new_n2440 );
  nor      g2324 ( new_n2710 , pi013 , new_n2463 );
  nor      g2325 ( new_n2711 , pi051 , new_n2710 );
  nor      g2326 ( new_n2712 , pi168 , new_n2711 );
  nor      g2327 ( new_n2713 , pi179 , new_n2712 );
  nor      g2328 ( new_n2714 , pi106 , new_n2713 );
  nor      g2329 ( new_n2715 , new_n2027 , new_n2714 );
  nor      g2330 ( new_n2716 , new_n2053 , new_n2715 );
  nor      g2331 ( new_n2717 , new_n2022 , new_n2716 );
  nor      g2332 ( po051 , new_n500 , new_n2717 );
  nor      g2333 ( new_n2719 , new_n918 , new_n2545 );
  nand g2334 ( new_n2720 , new_n2524 , new_n2524 );
  nor      g2335 ( new_n2721 , new_n801 , new_n1884 );
  nand     g2336 ( new_n2722 , new_n2163 , new_n2721 );
  nor      g2337 ( new_n2723 , new_n2340 , new_n2722 );
  nand     g2338 ( new_n2724 , new_n1728 , new_n2723 );
  nor      g2339 ( new_n2725 , new_n2657 , new_n2724 );
  nand     g2340 ( new_n2726 , new_n2414 , new_n2725 );
  nor      g2341 ( new_n2727 , new_n2720 , new_n2726 );
  nor      g2342 ( new_n2728 , new_n2719 , new_n2727 );
  and      g2343 ( new_n2729 , new_n1016 , new_n2728 );
  nand     g2344 ( new_n2730 , pi124 , new_n1092 );
  nor      g2345 ( po052 , new_n2729 , new_n2730 );
  nand     g2346 ( new_n2732 , new_n493 , new_n2302 );
  nand     g2347 ( new_n2733 , new_n2476 , new_n2732 );
  nand     g2348 ( new_n2734 , new_n2350 , new_n2733 );
  nand     g2349 ( new_n2735 , new_n1335 , new_n2734 );
  and      g2350 ( new_n2736 , new_n1812 , new_n2735 );
  nor      g2351 ( po053 , new_n398 , new_n2736 );
  nand g2352 ( new_n2738 , new_n2510 , new_n2510 );
  or       g2353 ( new_n2739 , new_n2738 , new_n2614 );
  nand     g2354 ( new_n2740 , new_n2618 , new_n2739 );
  and      g2355 ( po054 , pi071 , new_n2740 );
  nand g2356 ( new_n2742 , new_n2277 , new_n2277 );
  nor      g2357 ( new_n2743 , pi202 , new_n2742 );
  nand     g2358 ( new_n2744 , pi085 , new_n1034 );
  nor      g2359 ( po055 , new_n2743 , new_n2744 );
  nor      g2360 ( new_n2746 , pi215 , new_n1908 );
  nor      g2361 ( new_n2747 , pi105 , new_n2746 );
  nor      g2362 ( po056 , new_n513 , new_n2747 );
  nor      g2363 ( new_n2749 , new_n2150 , new_n2687 );
  nor      g2364 ( new_n2750 , new_n561 , new_n2749 );
  nor      g2365 ( po057 , new_n434 , new_n2750 );
  nand     g2366 ( new_n2752 , new_n2447 , new_n2662 );
  nand     g2367 ( new_n2753 , new_n2641 , new_n2752 );
  nand     g2368 ( new_n2754 , new_n1159 , new_n2753 );
  nor      g2369 ( new_n2755 , new_n980 , new_n2754 );
  nor      g2370 ( new_n2756 , pi217 , new_n2755 );
  nor      g2371 ( po058 , new_n622 , new_n2756 );
  nand g2372 ( new_n2758 , new_n2335 , new_n2335 );
  nand g2373 ( new_n2759 , new_n837 , new_n837 );
  nand     g2374 ( new_n2760 , new_n840 , new_n843 );
  nor      g2375 ( new_n2761 , new_n2759 , new_n2760 );
  nand     g2376 ( new_n2762 , new_n1180 , new_n1363 );
  nor      g2377 ( new_n2763 , new_n2761 , new_n2762 );
  nand     g2378 ( new_n2764 , new_n1872 , new_n2109 );
  nor      g2379 ( new_n2765 , new_n2763 , new_n2764 );
  nor      g2380 ( new_n2766 , new_n2394 , new_n2765 );
  nor      g2381 ( new_n2767 , new_n2336 , new_n2766 );
  nor      g2382 ( new_n2768 , new_n2758 , new_n2767 );
  nand g2383 ( new_n2769 , new_n1098 , new_n1098 );
  nor      g2384 ( new_n2770 , new_n2336 , new_n2378 );
  nor      g2385 ( new_n2771 , new_n2769 , new_n2770 );
  nand     g2386 ( new_n2772 , new_n2768 , new_n2771 );
  nand g2387 ( new_n2773 , new_n2772 , new_n2772 );
  nor      g2388 ( new_n2774 , pi191 , new_n2773 );
  nor      g2389 ( new_n2775 , pi045 , new_n2774 );
  nor      g2390 ( new_n2776 , new_n860 , new_n1103 );
  nand     g2391 ( new_n2777 , new_n2776 , new_n2768 );
  nand g2392 ( new_n2778 , new_n2777 , new_n2777 );
  nor      g2393 ( new_n2779 , new_n2775 , new_n2778 );
  nor      g2394 ( new_n2780 , pi058 , new_n2779 );
  nand     g2395 ( new_n2781 , pi046 , new_n752 );
  nor      g2396 ( po059 , new_n2780 , new_n2781 );
  nor      g2397 ( new_n2783 , new_n1670 , new_n974 );
  and      g2398 ( new_n2784 , new_n979 , new_n2783 );
  nand     g2399 ( new_n2785 , new_n972 , new_n2784 );
  nor      g2400 ( po060 , new_n2754 , new_n2785 );
  nand g2401 ( new_n2787 , new_n814 , new_n814 );
  nand     g2402 ( new_n2788 , pi208 , new_n2787 );
  nor      g2403 ( po061 , new_n2419 , new_n2788 );
  or       g2404 ( new_n2790 , new_n2027 , new_n2714 );
  nand     g2405 ( new_n2791 , new_n2052 , new_n2790 );
  nor      g2406 ( po062 , new_n995 , new_n2791 );
  nor      g2407 ( new_n2793 , pi000 , new_n2273 );
  nor      g2408 ( new_n2794 , pi161 , new_n2793 );
  nand     g2409 ( new_n2795 , pi231 , new_n1234 );
  nor      g2410 ( po063 , new_n2794 , new_n2795 );
  and      g2411 ( po064 , pi145 , new_n1688 );
  nand g2412 ( new_n2798 , new_n2026 , new_n2026 );
  nand g2413 ( new_n2799 , new_n2102 , new_n2102 );
  nand g2414 ( new_n2800 , new_n2075 , new_n2075 );
  nand     g2415 ( new_n2801 , new_n2080 , new_n2384 );
  nor      g2416 ( new_n2802 , new_n2800 , new_n2801 );
  nor      g2417 ( new_n2803 , new_n2399 , new_n2802 );
  nor      g2418 ( new_n2804 , new_n2799 , new_n2803 );
  nor      g2419 ( new_n2805 , new_n2798 , new_n2804 );
  nand     g2420 ( new_n2806 , pi050 , new_n525 );
  nand     g2421 ( new_n2807 , new_n2050 , new_n2806 );
  nor      g2422 ( new_n2808 , new_n2805 , new_n2807 );
  nor      g2423 ( new_n2809 , pi067 , new_n2808 );
  nand     g2424 ( new_n2810 , pi252 , new_n524 );
  nor      g2425 ( po065 , new_n2809 , new_n2810 );
  and      g2426 ( po066 , pi079 , new_n2808 );
  nor      g2427 ( new_n2813 , new_n1610 , new_n2573 );
  nand     g2428 ( new_n2814 , new_n2266 , new_n2813 );
  nor      g2429 ( new_n2815 , new_n2446 , new_n2814 );
  nor      g2430 ( new_n2816 , new_n2339 , new_n2815 );
  nand     g2431 ( new_n2817 , new_n891 , new_n1780 );
  nor      g2432 ( new_n2818 , new_n2816 , new_n2817 );
  nor      g2433 ( new_n2819 , new_n1611 , new_n2818 );
  nor      g2434 ( po067 , new_n656 , new_n2819 );
  nand     g2435 ( new_n2821 , pi166 , new_n578 );
  nor      g2436 ( po068 , new_n2670 , new_n2821 );
  nand     g2437 ( new_n2823 , pi229 , new_n784 );
  nor      g2438 ( po069 , new_n2547 , new_n2823 );
  nor      g2439 ( new_n2825 , new_n1274 , new_n2554 );
  nand     g2440 ( new_n2826 , pi028 , new_n1271 );
  nor      g2441 ( po070 , new_n2825 , new_n2826 );
  nand     g2442 ( new_n2828 , new_n2196 , new_n2232 );
  nand     g2443 ( new_n2829 , new_n1789 , new_n2828 );
  nand     g2444 ( new_n2830 , new_n1786 , new_n2829 );
  nand g2445 ( new_n2831 , new_n2830 , new_n2830 );
  nand     g2446 ( new_n2832 , new_n2651 , new_n1906 );
  nor      g2447 ( new_n2833 , new_n2831 , new_n2832 );
  nor      g2448 ( new_n2834 , new_n2654 , new_n2833 );
  nor      g2449 ( new_n2835 , new_n542 , new_n2834 );
  nor      g2450 ( new_n2836 , new_n2256 , new_n2835 );
  nor      g2451 ( new_n2837 , new_n2137 , new_n2836 );
  nor      g2452 ( new_n2838 , new_n1832 , new_n2837 );
  nor      g2453 ( new_n2839 , pi012 , new_n2838 );
  nor      g2454 ( po071 , new_n448 , new_n2839 );
  nor      g2455 ( new_n2841 , new_n912 , new_n2511 );
  nor      g2456 ( new_n2842 , pi031 , new_n2841 );
  nor      g2457 ( po072 , new_n2581 , new_n2842 );
  nor      g2458 ( new_n2844 , new_n1218 , new_n2657 );
  nor      g2459 ( new_n2845 , new_n2660 , new_n2844 );
  nor      g2460 ( new_n2846 , new_n1939 , new_n2845 );
  nor      g2461 ( new_n2847 , new_n1404 , new_n2846 );
  nor      g2462 ( new_n2848 , new_n1252 , new_n2847 );
  nand     g2463 ( new_n2849 , new_n1139 , new_n1282 );
  nor      g2464 ( new_n2850 , new_n2848 , new_n2849 );
  nor      g2465 ( new_n2851 , pi236 , new_n2850 );
  nor      g2466 ( new_n2852 , pi097 , new_n2851 );
  nor      g2467 ( po073 , new_n1253 , new_n2852 );
  nor      g2468 ( new_n2854 , pi143 , new_n2717 );
  nor      g2469 ( new_n2855 , new_n487 , new_n2854 );
  nand     g2470 ( new_n2856 , pi199 , new_n490 );
  nor      g2471 ( po074 , new_n2855 , new_n2856 );
  nor      g2472 ( po075 , new_n1224 , new_n2850 );
  nand     g2473 ( new_n2859 , new_n846 , new_n1356 );
  nand     g2474 ( new_n2860 , pi151 , new_n2859 );
  nor      g2475 ( po076 , new_n2778 , new_n2860 );
  nor      g2476 ( new_n2862 , new_n2759 , new_n1663 );
  nor      g2477 ( new_n2863 , new_n1746 , new_n2862 );
  nand     g2478 ( new_n2864 , pi158 , new_n1767 );
  nor      g2479 ( po077 , new_n2863 , new_n2864 );
  nor      g2480 ( new_n2866 , new_n1323 , new_n2355 );
  nor      g2481 ( po078 , new_n1319 , new_n2866 );
  nor      g2482 ( new_n2868 , pi201 , new_n2819 );
  nor      g2483 ( new_n2869 , pi078 , new_n2868 );
  nor      g2484 ( new_n2870 , pi196 , new_n2869 );
  nor      g2485 ( new_n2871 , pi247 , new_n2870 );
  nor      g2486 ( po079 , new_n901 , new_n2871 );
  nor      g2487 ( new_n2873 , new_n625 , new_n2755 );
  nand     g2488 ( new_n2874 , pi019 , new_n623 );
  nor      g2489 ( po080 , new_n2873 , new_n2874 );
  nor      g2490 ( po081 , new_n570 , new_n2705 );
  nor      g2491 ( new_n2877 , pi198 , new_n2791 );
  nor      g2492 ( new_n2878 , pi047 , new_n2877 );
  nor      g2493 ( po082 , new_n509 , new_n2878 );
  nor      g2494 ( new_n2880 , pi025 , new_n2854 );
  nor      g2495 ( po083 , new_n488 , new_n2880 );
  nand     g2496 ( new_n2882 , pi110 , new_n779 );
  nor      g2497 ( po084 , new_n2728 , new_n2882 );
  nand     g2498 ( new_n2884 , pi139 , new_n1831 );
  nor      g2499 ( po085 , new_n2837 , new_n2884 );
  nor      g2500 ( new_n2886 , pi150 , new_n2550 );
  nor      g2501 ( new_n2887 , pi004 , new_n2886 );
  nor      g2502 ( po086 , new_n761 , new_n2887 );
  nor      g2503 ( new_n2889 , pi220 , new_n2436 );
  nor      g2504 ( new_n2890 , pi069 , new_n2889 );
  nor      g2505 ( po087 , new_n424 , new_n2890 );
  nand g2506 ( new_n2892 , new_n2225 , new_n2225 );
  nand     g2507 ( new_n2893 , new_n1646 , new_n2892 );
  and      g2508 ( new_n2894 , new_n1286 , new_n2893 );
  nand     g2509 ( new_n2895 , pi065 , new_n1118 );
  nor      g2510 ( po088 , new_n2894 , new_n2895 );
  nand     g2511 ( new_n2897 , pi239 , new_n435 );
  nor      g2512 ( po089 , new_n1951 , new_n2897 );
  and      g2513 ( new_n2899 , new_n949 , new_n2370 );
  nand     g2514 ( new_n2900 , pi116 , new_n941 );
  nor      g2515 ( po090 , new_n2899 , new_n2900 );
  and      g2516 ( po091 , pi064 , new_n2779 );
  nor      g2517 ( new_n2903 , pi016 , new_n2839 );
  nor      g2518 ( new_n2904 , pi152 , new_n2903 );
  nor      g2519 ( po092 , new_n449 , new_n2904 );
  nor      g2520 ( new_n2906 , pi248 , new_n2707 );
  nor      g2521 ( new_n2907 , pi100 , new_n2906 );
  nor      g2522 ( new_n2908 , pi063 , new_n2907 );
  nor      g2523 ( new_n2909 , pi113 , new_n2908 );
  nor      g2524 ( po093 , new_n968 , new_n2909 );
  nor      g2525 ( new_n2911 , new_n2064 , new_n2433 );
  nand     g2526 ( new_n2912 , pi232 , new_n1807 );
  nor      g2527 ( po094 , new_n2911 , new_n2912 );
  nor      g2528 ( po095 , new_n478 , new_n2534 );
  nor      g2529 ( new_n2915 , pi246 , new_n2736 );
  nor      g2530 ( new_n2916 , pi128 , new_n2915 );
  nor      g2531 ( po096 , new_n392 , new_n2916 );
  nor      g2532 ( new_n2918 , new_n546 , new_n2431 );
  nand     g2533 ( new_n2919 , pi126 , new_n447 );
  nor      g2534 ( po097 , new_n2918 , new_n2919 );
  nor      g2535 ( new_n2921 , pi076 , new_n1952 );
  nor      g2536 ( po098 , new_n439 , new_n2921 );
  or       g2537 ( new_n2923 , new_n1663 , new_n1770 );
  and      g2538 ( new_n2924 , new_n1363 , new_n2923 );
  nand     g2539 ( new_n2925 , pi104 , new_n1364 );
  nor      g2540 ( po099 , new_n2924 , new_n2925 );
  nor      g2541 ( po100 , new_n2146 , new_n2434 );
  nand g2542 ( new_n2928 , new_n831 , new_n831 );
  nand     g2543 ( new_n2929 , pi243 , new_n2928 );
  nor      g2544 ( po101 , new_n1689 , new_n2929 );
  nand     g2545 ( new_n2931 , new_n737 , new_n2600 );
  nand     g2546 ( new_n2932 , new_n1067 , new_n2931 );
  nor      g2547 ( po102 , new_n2521 , new_n2932 );
  and      g2548 ( new_n2934 , new_n1384 , new_n2768 );
  nand     g2549 ( new_n2935 , new_n722 , new_n1357 );
  nor      g2550 ( new_n2936 , new_n2934 , new_n2935 );
  or       g2551 ( new_n2937 , pi140 , new_n847 );
  nor      g2552 ( new_n2938 , new_n2936 , new_n2937 );
  nor      g2553 ( po103 , new_n721 , new_n2938 );
  nor      g2554 ( new_n2940 , pi148 , new_n2932 );
  nor      g2555 ( new_n2941 , pi086 , new_n2940 );
  nor      g2556 ( po104 , new_n744 , new_n2941 );
  nand     g2557 ( new_n2943 , pi122 , new_n1221 );
  nor      g2558 ( po105 , new_n2847 , new_n2943 );
  or       g2559 ( new_n2945 , new_n2271 , new_n2734 );
  and      g2560 ( new_n2946 , new_n2230 , new_n2945 );
  nor      g2561 ( new_n2947 , new_n1278 , new_n2946 );
  nor      g2562 ( po106 , new_n1251 , new_n2947 );
  nor      g2563 ( new_n2949 , new_n473 , new_n554 );
  and      g2564 ( po107 , new_n2686 , new_n2949 );
  nor      g2565 ( new_n2951 , pi131 , new_n386 );
  nor      g2566 ( new_n2952 , new_n1259 , new_n2951 );
  and      g2567 ( po108 , new_n1957 , new_n2952 );
  nor      g2568 ( new_n2954 , new_n866 , new_n2629 );
  nor      g2569 ( po109 , new_n1585 , new_n2954 );
  nand     g2570 ( new_n2956 , pi173 , new_n821 );
  nor      g2571 ( po110 , new_n1663 , new_n2956 );
  nor      g2572 ( new_n2958 , new_n612 , new_n2671 );
  nand     g2573 ( new_n2959 , pi219 , new_n614 );
  nor      g2574 ( po111 , new_n2958 , new_n2959 );
  nor      g2575 ( new_n2961 , pi221 , new_n2620 );
  nor      g2576 ( new_n2962 , pi224 , new_n2961 );
  nor      g2577 ( po112 , new_n602 , new_n2962 );
  nor      g2578 ( po113 , new_n1622 , new_n2907 );
  nand g2579 ( new_n2965 , new_n2838 , new_n2838 );
  nor      g2580 ( new_n2966 , new_n450 , new_n2965 );
  nor      g2581 ( new_n2967 , new_n2073 , new_n2966 );
  nor      g2582 ( po114 , new_n1432 , new_n2967 );
  nor      g2583 ( new_n2969 , new_n1485 , new_n2892 );
  nand     g2584 ( new_n2970 , pi157 , new_n1238 );
  or       g2585 ( new_n2971 , new_n1515 , new_n2970 );
  nor      g2586 ( po115 , new_n2969 , new_n2971 );
  nor      g2587 ( new_n2973 , new_n399 , new_n2735 );
  nor      g2588 ( new_n2974 , new_n2468 , new_n2973 );
  nor      g2589 ( po116 , new_n2128 , new_n2974 );
  and      g2590 ( po117 , pi121 , new_n2734 );
  nand     g2591 ( new_n2977 , pi000 , new_n1760 );
  nor      g2592 ( po118 , new_n2273 , new_n2977 );
  nor      g2593 ( po119 , new_n683 , new_n2711 );
  nor      g2594 ( new_n2980 , pi002 , new_n2373 );
  nor      g2595 ( new_n2981 , pi096 , new_n2980 );
  nor      g2596 ( po120 , new_n937 , new_n2981 );
  nor      g2597 ( po121 , new_n581 , new_n1999 );
  nor      g2598 ( po122 , new_n654 , new_n2869 );
  nor      g2599 ( new_n2985 , pi245 , new_n2489 );
  nor      g2600 ( new_n2986 , pi101 , new_n2985 );
  nor      g2601 ( po123 , new_n1021 , new_n2986 );
  nor      g2602 ( po124 , new_n479 , new_n2532 );
  nor      g2603 ( po125 , new_n1702 , new_n2713 );
  nand     g2604 ( new_n2990 , pi091 , new_n911 );
  nor      g2605 ( po126 , new_n2511 , new_n2990 );
  nor      g2606 ( new_n2992 , new_n1097 , new_n2886 );
  nand     g2607 ( new_n2993 , pi191 , new_n1096 );
  nor      g2608 ( po127 , new_n2992 , new_n2993 );
  nor      g2609 ( new_n2995 , new_n938 , new_n1113 );
  and      g2610 ( new_n2996 , new_n937 , new_n1133 );
  and      g2611 ( new_n2997 , new_n2486 , new_n2996 );
  nor      g2612 ( new_n2998 , new_n2995 , new_n2997 );
  nor      g2613 ( po128 , new_n1023 , new_n2998 );
endmodule


