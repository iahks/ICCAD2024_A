 module top_809960632_810038711_1598227639_893650103 (a, b, o);

      input a, b; output o; nand_3 g0(a,b,o); endmodule