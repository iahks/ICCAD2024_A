// Benchmark "top_810222779_843330999_776144567_776418743_1234615" written by ABC on Wed Aug 14 20:29:23 2024

module top_810222779_843330999_776144567_776418743_1234615 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107;
  wire new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n548, new_n549,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n974, new_n975, new_n976, new_n977, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1017,
    new_n1022, new_n1023, new_n1024, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1303, new_n1306, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332;
  not_3  g0000(.A(pi153), .Y(new_n316));
  nand_5 g0001(.A(pi123), .B(pi000), .Y(new_n317));
  not_3  g0002(.A(new_n317), .Y(new_n318));
  not_3  g0003(.A(pi150), .Y(new_n319));
  nor_5  g0004(.A(new_n319), .B(pi026), .Y(new_n320));
  nor_5  g0005(.A(new_n320), .B(new_n318), .Y(new_n321));
  xor_4  g0006(.A(new_n321), .B(new_n316), .Y(new_n322));
  or_6   g0007(.A(new_n319), .B(pi054), .Y(new_n323));
  nand_5 g0008(.A(new_n323), .B(new_n317), .Y(new_n324));
  nand_5 g0009(.A(new_n324), .B(pi050), .Y(new_n325));
  not_3  g0010(.A(new_n325), .Y(new_n326));
  or_6   g0011(.A(new_n319), .B(pi115), .Y(new_n327));
  nand_5 g0012(.A(new_n327), .B(new_n317), .Y(new_n328));
  nand_5 g0013(.A(new_n328), .B(pi056), .Y(new_n329));
  not_3  g0014(.A(new_n329), .Y(new_n330));
  not_3  g0015(.A(pi122), .Y(new_n331));
  nor_5  g0016(.A(pi154), .B(new_n319), .Y(new_n332));
  nor_5  g0017(.A(new_n332), .B(new_n318), .Y(new_n333));
  nand_5 g0018(.A(new_n333), .B(new_n331), .Y(new_n334));
  xor_4  g0019(.A(new_n333), .B(new_n331), .Y(new_n335));
  not_3  g0020(.A(pi047), .Y(new_n336));
  nor_5  g0021(.A(pi175), .B(new_n319), .Y(new_n337));
  nor_5  g0022(.A(new_n337), .B(new_n318), .Y(new_n338));
  nand_5 g0023(.A(new_n338), .B(new_n336), .Y(new_n339));
  xor_4  g0024(.A(new_n338), .B(new_n336), .Y(new_n340));
  nor_5  g0025(.A(pi186), .B(pi150), .Y(new_n341));
  nor_5  g0026(.A(pi182), .B(new_n319), .Y(new_n342));
  nor_5  g0027(.A(new_n342), .B(new_n341), .Y(new_n343));
  not_3  g0028(.A(new_n343), .Y(new_n344));
  nand_5 g0029(.A(new_n344), .B(pi196), .Y(new_n345));
  not_3  g0030(.A(new_n345), .Y(new_n346));
  nor_5  g0031(.A(new_n344), .B(pi196), .Y(new_n347));
  not_3  g0032(.A(pi199), .Y(new_n348));
  nand_5 g0033(.A(pi150), .B(pi009), .Y(new_n349));
  nand_5 g0034(.A(pi177), .B(new_n319), .Y(new_n350));
  nand_5 g0035(.A(new_n350), .B(new_n349), .Y(new_n351));
  nand_5 g0036(.A(new_n351), .B(new_n348), .Y(new_n352));
  xor_4  g0037(.A(new_n351), .B(new_n348), .Y(new_n353));
  not_3  g0038(.A(pi178), .Y(new_n354));
  nand_5 g0039(.A(pi150), .B(pi080), .Y(new_n355));
  nand_5 g0040(.A(pi203), .B(new_n319), .Y(new_n356));
  nand_5 g0041(.A(new_n356), .B(new_n355), .Y(new_n357));
  nand_5 g0042(.A(new_n357), .B(new_n354), .Y(new_n358));
  or_6   g0043(.A(new_n357), .B(new_n354), .Y(new_n359));
  not_3  g0044(.A(pi162), .Y(new_n360));
  nand_5 g0045(.A(pi151), .B(new_n319), .Y(new_n361));
  nand_5 g0046(.A(pi172), .B(pi150), .Y(new_n362));
  nand_5 g0047(.A(new_n362), .B(new_n361), .Y(new_n363));
  nand_5 g0048(.A(new_n363), .B(new_n360), .Y(new_n364));
  xor_4  g0049(.A(new_n363), .B(new_n360), .Y(new_n365));
  not_3  g0050(.A(pi160), .Y(new_n366));
  not_3  g0051(.A(pi034), .Y(new_n367));
  nand_5 g0052(.A(new_n319), .B(new_n367), .Y(new_n368));
  not_3  g0053(.A(new_n368), .Y(new_n369));
  nor_5  g0054(.A(pi164), .B(new_n319), .Y(new_n370));
  nor_5  g0055(.A(new_n370), .B(new_n369), .Y(new_n371));
  nand_5 g0056(.A(new_n371), .B(new_n366), .Y(new_n372));
  xor_4  g0057(.A(new_n371), .B(new_n366), .Y(new_n373));
  not_3  g0058(.A(pi192), .Y(new_n374));
  nand_5 g0059(.A(new_n319), .B(pi139), .Y(new_n375));
  nand_5 g0060(.A(pi150), .B(pi090), .Y(new_n376));
  nand_5 g0061(.A(new_n376), .B(new_n375), .Y(new_n377));
  nor_5  g0062(.A(new_n377), .B(new_n374), .Y(new_n378));
  xor_4  g0063(.A(new_n377), .B(new_n374), .Y(new_n379));
  not_3  g0064(.A(new_n379), .Y(new_n380));
  not_3  g0065(.A(pi116), .Y(new_n381));
  nand_5 g0066(.A(pi158), .B(pi150), .Y(new_n382));
  nand_5 g0067(.A(new_n319), .B(pi146), .Y(new_n383));
  nand_5 g0068(.A(new_n383), .B(new_n382), .Y(new_n384));
  nand_5 g0069(.A(new_n384), .B(new_n381), .Y(new_n385));
  or_6   g0070(.A(new_n384), .B(new_n381), .Y(new_n386));
  not_3  g0071(.A(pi039), .Y(new_n387));
  nand_5 g0072(.A(new_n319), .B(pi086), .Y(new_n388));
  nand_5 g0073(.A(pi150), .B(pi030), .Y(new_n389));
  nand_5 g0074(.A(new_n389), .B(new_n388), .Y(new_n390));
  nand_5 g0075(.A(new_n390), .B(new_n387), .Y(new_n391));
  not_3  g0076(.A(pi057), .Y(new_n392));
  nand_5 g0077(.A(new_n319), .B(pi142), .Y(new_n393));
  nand_5 g0078(.A(pi150), .B(pi032), .Y(new_n394));
  nand_5 g0079(.A(new_n394), .B(new_n393), .Y(new_n395));
  nor_5  g0080(.A(new_n395), .B(new_n392), .Y(new_n396));
  xor_4  g0081(.A(new_n395), .B(new_n392), .Y(new_n397));
  not_3  g0082(.A(new_n397), .Y(new_n398));
  not_3  g0083(.A(pi183), .Y(new_n399));
  not_3  g0084(.A(pi107), .Y(new_n400));
  nand_5 g0085(.A(pi189), .B(new_n319), .Y(new_n401));
  nand_5 g0086(.A(pi150), .B(pi106), .Y(new_n402));
  nand_5 g0087(.A(new_n402), .B(new_n401), .Y(new_n403));
  nor_5  g0088(.A(new_n403), .B(new_n400), .Y(new_n404));
  xor_4  g0089(.A(new_n403), .B(new_n400), .Y(new_n405));
  not_3  g0090(.A(new_n405), .Y(new_n406));
  not_3  g0091(.A(pi020), .Y(new_n407));
  nand_5 g0092(.A(pi194), .B(pi150), .Y(new_n408));
  nand_5 g0093(.A(pi156), .B(new_n319), .Y(new_n409));
  nand_5 g0094(.A(new_n409), .B(new_n408), .Y(new_n410));
  nand_5 g0095(.A(new_n410), .B(new_n407), .Y(new_n411));
  or_6   g0096(.A(new_n410), .B(new_n407), .Y(new_n412));
  not_3  g0097(.A(pi170), .Y(new_n413));
  nand_5 g0098(.A(pi150), .B(pi012), .Y(new_n414));
  nand_5 g0099(.A(new_n319), .B(pi131), .Y(new_n415));
  nand_5 g0100(.A(new_n415), .B(new_n414), .Y(new_n416));
  nor_5  g0101(.A(new_n416), .B(new_n413), .Y(new_n417));
  not_3  g0102(.A(pi051), .Y(new_n418));
  nand_5 g0103(.A(pi150), .B(pi087), .Y(new_n419));
  nand_5 g0104(.A(new_n319), .B(pi014), .Y(new_n420));
  nand_5 g0105(.A(new_n420), .B(new_n419), .Y(new_n421));
  nor_5  g0106(.A(new_n421), .B(new_n418), .Y(new_n422));
  not_3  g0107(.A(pi074), .Y(new_n423));
  not_3  g0108(.A(pi180), .Y(new_n424));
  nand_5 g0109(.A(pi169), .B(pi150), .Y(new_n425));
  nand_5 g0110(.A(new_n319), .B(pi033), .Y(new_n426));
  nand_5 g0111(.A(new_n426), .B(new_n425), .Y(new_n427));
  nand_5 g0112(.A(new_n427), .B(new_n424), .Y(new_n428));
  xor_4  g0113(.A(new_n427), .B(new_n424), .Y(new_n429));
  not_3  g0114(.A(pi027), .Y(new_n430));
  nand_5 g0115(.A(new_n319), .B(pi042), .Y(new_n431));
  nand_5 g0116(.A(pi150), .B(pi044), .Y(new_n432));
  nand_5 g0117(.A(new_n432), .B(new_n431), .Y(new_n433));
  nand_5 g0118(.A(new_n433), .B(new_n430), .Y(new_n434));
  not_3  g0119(.A(pi083), .Y(new_n435));
  nand_5 g0120(.A(new_n319), .B(pi007), .Y(new_n436));
  nand_5 g0121(.A(pi197), .B(pi150), .Y(new_n437));
  nand_5 g0122(.A(new_n437), .B(new_n436), .Y(new_n438));
  nand_5 g0123(.A(new_n438), .B(new_n435), .Y(new_n439));
  not_3  g0124(.A(pi132), .Y(new_n440));
  nand_5 g0125(.A(new_n319), .B(pi143), .Y(new_n441));
  nand_5 g0126(.A(pi150), .B(pi043), .Y(new_n442));
  nand_5 g0127(.A(new_n442), .B(new_n441), .Y(new_n443));
  nand_5 g0128(.A(new_n443), .B(new_n440), .Y(new_n444));
  not_3  g0129(.A(pi004), .Y(new_n445));
  nand_5 g0130(.A(new_n319), .B(pi058), .Y(new_n446));
  nand_5 g0131(.A(pi150), .B(pi025), .Y(new_n447));
  nand_5 g0132(.A(new_n447), .B(new_n446), .Y(new_n448));
  nand_5 g0133(.A(new_n448), .B(new_n445), .Y(new_n449));
  not_3  g0134(.A(pi092), .Y(new_n450));
  nand_5 g0135(.A(pi193), .B(pi150), .Y(new_n451));
  nand_5 g0136(.A(pi152), .B(new_n319), .Y(new_n452));
  nand_5 g0137(.A(new_n452), .B(new_n451), .Y(new_n453));
  nand_5 g0138(.A(new_n453), .B(new_n450), .Y(new_n454));
  not_3  g0139(.A(pi070), .Y(new_n455));
  or_6   g0140(.A(pi147), .B(pi069), .Y(new_n456));
  and_6  g0141(.A(pi147), .B(pi069), .Y(new_n457));
  nor_5  g0142(.A(new_n457), .B(pi150), .Y(new_n458));
  and_6  g0143(.A(new_n458), .B(new_n456), .Y(new_n459));
  nor_5  g0144(.A(new_n459), .B(new_n455), .Y(new_n460));
  and_6  g0145(.A(new_n458), .B(pi069), .Y(new_n461));
  or_6   g0146(.A(new_n461), .B(new_n460), .Y(new_n462));
  xor_4  g0147(.A(new_n453), .B(new_n450), .Y(new_n463));
  nand_5 g0148(.A(new_n463), .B(new_n462), .Y(new_n464));
  nand_5 g0149(.A(new_n464), .B(new_n454), .Y(new_n465));
  nand_5 g0150(.A(new_n448), .B(pi004), .Y(new_n466));
  or_6   g0151(.A(new_n448), .B(pi004), .Y(new_n467));
  nand_5 g0152(.A(new_n467), .B(new_n466), .Y(new_n468));
  nand_5 g0153(.A(new_n468), .B(new_n465), .Y(new_n469));
  nand_5 g0154(.A(new_n469), .B(new_n449), .Y(new_n470));
  xor_4  g0155(.A(new_n443), .B(pi132), .Y(new_n471));
  not_3  g0156(.A(new_n471), .Y(new_n472));
  nand_5 g0157(.A(new_n472), .B(new_n470), .Y(new_n473));
  nand_5 g0158(.A(new_n473), .B(new_n444), .Y(new_n474));
  nor_5  g0159(.A(new_n438), .B(new_n435), .Y(new_n475));
  not_3  g0160(.A(new_n475), .Y(new_n476));
  nand_5 g0161(.A(new_n476), .B(new_n439), .Y(new_n477));
  not_3  g0162(.A(new_n477), .Y(new_n478));
  nand_5 g0163(.A(new_n478), .B(new_n474), .Y(new_n479));
  nand_5 g0164(.A(new_n479), .B(new_n439), .Y(new_n480));
  xor_4  g0165(.A(new_n433), .B(new_n430), .Y(new_n481));
  nand_5 g0166(.A(new_n481), .B(new_n480), .Y(new_n482));
  nand_5 g0167(.A(new_n482), .B(new_n434), .Y(new_n483));
  nand_5 g0168(.A(new_n483), .B(new_n429), .Y(new_n484));
  nand_5 g0169(.A(new_n484), .B(new_n428), .Y(new_n485));
  nor_5  g0170(.A(new_n485), .B(new_n423), .Y(new_n486));
  nand_5 g0171(.A(new_n319), .B(pi081), .Y(new_n487));
  nand_5 g0172(.A(pi150), .B(pi035), .Y(new_n488));
  nand_5 g0173(.A(new_n488), .B(new_n487), .Y(new_n489));
  xor_4  g0174(.A(new_n485), .B(pi074), .Y(new_n490));
  nor_5  g0175(.A(new_n490), .B(new_n489), .Y(new_n491));
  nor_5  g0176(.A(new_n491), .B(new_n486), .Y(new_n492));
  not_3  g0177(.A(new_n422), .Y(new_n493));
  nand_5 g0178(.A(new_n421), .B(new_n418), .Y(new_n494));
  and_6  g0179(.A(new_n494), .B(new_n493), .Y(new_n495));
  not_3  g0180(.A(new_n495), .Y(new_n496));
  nor_5  g0181(.A(new_n496), .B(new_n492), .Y(new_n497));
  nor_5  g0182(.A(new_n497), .B(new_n422), .Y(new_n498));
  xor_4  g0183(.A(new_n416), .B(pi170), .Y(new_n499));
  nor_5  g0184(.A(new_n499), .B(new_n498), .Y(new_n500));
  nor_5  g0185(.A(new_n500), .B(new_n417), .Y(new_n501));
  nand_5 g0186(.A(new_n501), .B(new_n412), .Y(new_n502));
  nand_5 g0187(.A(new_n502), .B(new_n411), .Y(new_n503));
  nor_5  g0188(.A(new_n503), .B(new_n406), .Y(new_n504));
  nor_5  g0189(.A(new_n504), .B(new_n404), .Y(new_n505));
  nor_5  g0190(.A(new_n505), .B(new_n399), .Y(new_n506));
  xor_4  g0191(.A(new_n505), .B(pi183), .Y(new_n507));
  nand_5 g0192(.A(pi187), .B(pi150), .Y(new_n508));
  nand_5 g0193(.A(new_n319), .B(pi094), .Y(new_n509));
  nand_5 g0194(.A(new_n509), .B(new_n508), .Y(new_n510));
  nor_5  g0195(.A(new_n510), .B(new_n507), .Y(new_n511));
  nor_5  g0196(.A(new_n511), .B(new_n506), .Y(new_n512));
  nor_5  g0197(.A(new_n512), .B(new_n398), .Y(new_n513));
  nor_5  g0198(.A(new_n513), .B(new_n396), .Y(new_n514));
  xor_4  g0199(.A(new_n390), .B(new_n387), .Y(new_n515));
  nand_5 g0200(.A(new_n515), .B(new_n514), .Y(new_n516));
  nand_5 g0201(.A(new_n516), .B(new_n391), .Y(new_n517));
  nand_5 g0202(.A(new_n517), .B(new_n386), .Y(new_n518));
  nand_5 g0203(.A(new_n518), .B(new_n385), .Y(new_n519));
  nor_5  g0204(.A(new_n519), .B(new_n380), .Y(new_n520));
  nor_5  g0205(.A(new_n520), .B(new_n378), .Y(new_n521));
  nand_5 g0206(.A(new_n521), .B(new_n373), .Y(new_n522));
  nand_5 g0207(.A(new_n522), .B(new_n372), .Y(new_n523));
  nand_5 g0208(.A(new_n523), .B(new_n365), .Y(new_n524));
  nand_5 g0209(.A(new_n524), .B(new_n364), .Y(new_n525));
  nand_5 g0210(.A(new_n525), .B(new_n359), .Y(new_n526));
  nand_5 g0211(.A(new_n526), .B(new_n358), .Y(new_n527));
  nand_5 g0212(.A(new_n527), .B(new_n353), .Y(new_n528));
  nand_5 g0213(.A(new_n528), .B(new_n352), .Y(new_n529));
  nor_5  g0214(.A(new_n529), .B(new_n347), .Y(new_n530));
  nor_5  g0215(.A(new_n530), .B(new_n346), .Y(new_n531));
  nand_5 g0216(.A(new_n531), .B(new_n340), .Y(new_n532));
  nand_5 g0217(.A(new_n532), .B(new_n339), .Y(new_n533));
  nand_5 g0218(.A(new_n533), .B(new_n335), .Y(new_n534));
  nand_5 g0219(.A(new_n534), .B(new_n334), .Y(new_n535));
  not_3  g0220(.A(pi056), .Y(new_n536));
  xor_4  g0221(.A(new_n328), .B(new_n536), .Y(new_n537));
  nor_5  g0222(.A(new_n537), .B(new_n535), .Y(new_n538));
  nor_5  g0223(.A(new_n538), .B(new_n330), .Y(new_n539));
  or_6   g0224(.A(new_n324), .B(pi050), .Y(new_n540));
  nand_5 g0225(.A(new_n540), .B(new_n325), .Y(new_n541));
  nor_5  g0226(.A(new_n541), .B(new_n539), .Y(new_n542));
  nor_5  g0227(.A(new_n542), .B(new_n326), .Y(new_n543));
  xor_4  g0228(.A(new_n543), .B(new_n322), .Y(po000));
  not_3  g0229(.A(pi165), .Y(new_n545));
  nand_5 g0230(.A(pi167), .B(new_n545), .Y(po003));
  xor_4  g0231(.A(new_n515), .B(new_n514), .Y(po005));
  nand_5 g0232(.A(pi075), .B(pi037), .Y(new_n548));
  nand_5 g0233(.A(pi198), .B(pi188), .Y(new_n549));
  or_6   g0234(.A(new_n549), .B(new_n548), .Y(po006));
  nor_5  g0235(.A(new_n319), .B(pi028), .Y(new_n551));
  not_3  g0236(.A(new_n551), .Y(new_n552));
  nand_5 g0237(.A(new_n552), .B(new_n317), .Y(new_n553));
  or_6   g0238(.A(pi150), .B(pi041), .Y(new_n554));
  nand_5 g0239(.A(pi181), .B(pi150), .Y(new_n555));
  nand_5 g0240(.A(new_n555), .B(new_n554), .Y(new_n556));
  and_6  g0241(.A(new_n556), .B(new_n553), .Y(new_n557));
  nand_5 g0242(.A(pi203), .B(pi140), .Y(new_n558));
  and_6  g0243(.A(pi177), .B(pi173), .Y(new_n559));
  nand_5 g0244(.A(pi186), .B(pi161), .Y(new_n560));
  nand_5 g0245(.A(new_n560), .B(new_n319), .Y(new_n561));
  nor_5  g0246(.A(new_n561), .B(new_n559), .Y(new_n562));
  nand_5 g0247(.A(new_n562), .B(new_n558), .Y(new_n563));
  and_6  g0248(.A(new_n317), .B(pi110), .Y(new_n564));
  nand_5 g0249(.A(new_n564), .B(new_n336), .Y(new_n565));
  not_3  g0250(.A(pi196), .Y(new_n566));
  nand_5 g0251(.A(new_n566), .B(pi119), .Y(new_n567));
  and_6  g0252(.A(new_n567), .B(pi150), .Y(new_n568));
  nand_5 g0253(.A(new_n568), .B(new_n565), .Y(new_n569));
  nand_5 g0254(.A(new_n354), .B(pi174), .Y(new_n570));
  nand_5 g0255(.A(new_n348), .B(pi006), .Y(new_n571));
  nand_5 g0256(.A(new_n571), .B(new_n570), .Y(new_n572));
  or_6   g0257(.A(new_n572), .B(new_n569), .Y(new_n573));
  nand_5 g0258(.A(new_n573), .B(new_n563), .Y(new_n574));
  nand_5 g0259(.A(new_n445), .B(pi002), .Y(new_n575));
  nand_5 g0260(.A(pi103), .B(pi091), .Y(new_n576));
  nand_5 g0261(.A(new_n576), .B(pi092), .Y(new_n577));
  or_6   g0262(.A(pi103), .B(pi091), .Y(new_n578));
  nand_5 g0263(.A(new_n578), .B(new_n577), .Y(new_n579));
  nand_5 g0264(.A(new_n579), .B(new_n575), .Y(new_n580));
  nor_5  g0265(.A(new_n440), .B(pi089), .Y(new_n581));
  nor_5  g0266(.A(new_n445), .B(pi002), .Y(new_n582));
  nor_5  g0267(.A(new_n582), .B(new_n581), .Y(new_n583));
  and_6  g0268(.A(new_n583), .B(new_n580), .Y(new_n584));
  nand_5 g0269(.A(new_n435), .B(pi055), .Y(new_n585));
  nand_5 g0270(.A(new_n440), .B(pi089), .Y(new_n586));
  nand_5 g0271(.A(new_n586), .B(new_n585), .Y(new_n587));
  nor_5  g0272(.A(new_n587), .B(new_n584), .Y(new_n588));
  nor_5  g0273(.A(pi067), .B(new_n430), .Y(new_n589));
  nor_5  g0274(.A(new_n435), .B(pi055), .Y(new_n590));
  or_6   g0275(.A(new_n590), .B(new_n589), .Y(new_n591));
  nor_5  g0276(.A(new_n591), .B(new_n588), .Y(new_n592));
  nand_5 g0277(.A(new_n424), .B(pi059), .Y(new_n593));
  nand_5 g0278(.A(pi067), .B(new_n430), .Y(new_n594));
  nand_5 g0279(.A(new_n594), .B(new_n593), .Y(new_n595));
  nor_5  g0280(.A(new_n595), .B(new_n592), .Y(new_n596));
  not_3  g0281(.A(pi059), .Y(new_n597));
  nand_5 g0282(.A(pi180), .B(new_n597), .Y(new_n598));
  or_6   g0283(.A(new_n423), .B(pi038), .Y(new_n599));
  nand_5 g0284(.A(new_n599), .B(new_n598), .Y(new_n600));
  nor_5  g0285(.A(new_n600), .B(new_n596), .Y(new_n601));
  nand_5 g0286(.A(new_n423), .B(pi038), .Y(new_n602));
  nand_5 g0287(.A(pi206), .B(new_n418), .Y(new_n603));
  nand_5 g0288(.A(new_n603), .B(new_n602), .Y(new_n604));
  nor_5  g0289(.A(new_n604), .B(new_n601), .Y(new_n605));
  not_3  g0290(.A(pi049), .Y(new_n606));
  nand_5 g0291(.A(pi170), .B(new_n606), .Y(new_n607));
  or_6   g0292(.A(pi206), .B(new_n418), .Y(new_n608));
  nand_5 g0293(.A(new_n608), .B(new_n607), .Y(new_n609));
  nor_5  g0294(.A(new_n609), .B(new_n605), .Y(new_n610));
  nand_5 g0295(.A(pi135), .B(new_n407), .Y(new_n611));
  nand_5 g0296(.A(new_n413), .B(pi049), .Y(new_n612));
  nand_5 g0297(.A(new_n612), .B(new_n611), .Y(new_n613));
  nor_5  g0298(.A(new_n613), .B(new_n610), .Y(new_n614));
  nor_5  g0299(.A(pi135), .B(new_n407), .Y(new_n615));
  nor_5  g0300(.A(new_n400), .B(pi011), .Y(new_n616));
  or_6   g0301(.A(new_n616), .B(new_n615), .Y(new_n617));
  nor_5  g0302(.A(new_n617), .B(new_n614), .Y(new_n618));
  nand_5 g0303(.A(pi195), .B(new_n399), .Y(new_n619));
  nand_5 g0304(.A(new_n400), .B(pi011), .Y(new_n620));
  nand_5 g0305(.A(new_n620), .B(new_n619), .Y(new_n621));
  nor_5  g0306(.A(new_n621), .B(new_n618), .Y(new_n622));
  or_6   g0307(.A(pi195), .B(new_n399), .Y(new_n623));
  not_3  g0308(.A(pi097), .Y(new_n624));
  nand_5 g0309(.A(new_n624), .B(pi057), .Y(new_n625));
  nand_5 g0310(.A(new_n625), .B(new_n623), .Y(new_n626));
  nor_5  g0311(.A(new_n626), .B(new_n622), .Y(new_n627));
  nand_5 g0312(.A(new_n387), .B(pi005), .Y(new_n628));
  nand_5 g0313(.A(pi097), .B(new_n392), .Y(new_n629));
  nand_5 g0314(.A(new_n629), .B(new_n628), .Y(new_n630));
  nor_5  g0315(.A(new_n630), .B(new_n627), .Y(new_n631));
  or_6   g0316(.A(new_n381), .B(pi114), .Y(new_n632));
  not_3  g0317(.A(pi005), .Y(new_n633));
  nand_5 g0318(.A(pi039), .B(new_n633), .Y(new_n634));
  nand_5 g0319(.A(new_n634), .B(new_n632), .Y(new_n635));
  nor_5  g0320(.A(new_n635), .B(new_n631), .Y(new_n636));
  nand_5 g0321(.A(new_n374), .B(pi036), .Y(new_n637));
  nand_5 g0322(.A(new_n381), .B(pi114), .Y(new_n638));
  nand_5 g0323(.A(new_n638), .B(new_n637), .Y(new_n639));
  nor_5  g0324(.A(new_n639), .B(new_n636), .Y(new_n640));
  nor_5  g0325(.A(new_n366), .B(pi052), .Y(new_n641));
  nor_5  g0326(.A(new_n374), .B(pi036), .Y(new_n642));
  or_6   g0327(.A(new_n642), .B(new_n641), .Y(new_n643));
  nor_5  g0328(.A(new_n643), .B(new_n640), .Y(new_n644));
  nand_5 g0329(.A(new_n366), .B(pi052), .Y(new_n645));
  nand_5 g0330(.A(new_n645), .B(pi150), .Y(new_n646));
  nor_5  g0331(.A(new_n646), .B(new_n644), .Y(new_n647));
  or_6   g0332(.A(pi091), .B(pi069), .Y(new_n648));
  and_6  g0333(.A(new_n648), .B(pi096), .Y(new_n649));
  nand_5 g0334(.A(pi152), .B(pi066), .Y(new_n650));
  nand_5 g0335(.A(pi091), .B(pi069), .Y(new_n651));
  nand_5 g0336(.A(new_n651), .B(new_n650), .Y(new_n652));
  nor_5  g0337(.A(new_n652), .B(new_n649), .Y(new_n653));
  nor_5  g0338(.A(pi152), .B(pi066), .Y(new_n654));
  nor_5  g0339(.A(pi111), .B(pi058), .Y(new_n655));
  or_6   g0340(.A(new_n655), .B(new_n654), .Y(new_n656));
  nor_5  g0341(.A(new_n656), .B(new_n653), .Y(new_n657));
  nand_5 g0342(.A(pi111), .B(pi058), .Y(new_n658));
  nand_5 g0343(.A(pi143), .B(pi048), .Y(new_n659));
  nand_5 g0344(.A(new_n659), .B(new_n658), .Y(new_n660));
  nor_5  g0345(.A(new_n660), .B(new_n657), .Y(new_n661));
  nor_5  g0346(.A(pi098), .B(pi007), .Y(new_n662));
  nor_5  g0347(.A(pi143), .B(pi048), .Y(new_n663));
  or_6   g0348(.A(new_n663), .B(new_n662), .Y(new_n664));
  nor_5  g0349(.A(new_n664), .B(new_n661), .Y(new_n665));
  nand_5 g0350(.A(pi042), .B(pi029), .Y(new_n666));
  nand_5 g0351(.A(pi098), .B(pi007), .Y(new_n667));
  nand_5 g0352(.A(new_n667), .B(new_n666), .Y(new_n668));
  nor_5  g0353(.A(new_n668), .B(new_n665), .Y(new_n669));
  nor_5  g0354(.A(pi033), .B(pi023), .Y(new_n670));
  nor_5  g0355(.A(pi042), .B(pi029), .Y(new_n671));
  or_6   g0356(.A(new_n671), .B(new_n670), .Y(new_n672));
  nor_5  g0357(.A(new_n672), .B(new_n669), .Y(new_n673));
  nand_5 g0358(.A(pi117), .B(pi081), .Y(new_n674));
  nand_5 g0359(.A(pi033), .B(pi023), .Y(new_n675));
  nand_5 g0360(.A(new_n675), .B(new_n674), .Y(new_n676));
  nor_5  g0361(.A(new_n676), .B(new_n673), .Y(new_n677));
  nor_5  g0362(.A(pi117), .B(pi081), .Y(new_n678));
  nor_5  g0363(.A(pi100), .B(pi014), .Y(new_n679));
  or_6   g0364(.A(new_n679), .B(new_n678), .Y(new_n680));
  nor_5  g0365(.A(new_n680), .B(new_n677), .Y(new_n681));
  nand_5 g0366(.A(pi149), .B(pi131), .Y(new_n682));
  nand_5 g0367(.A(pi100), .B(pi014), .Y(new_n683));
  nand_5 g0368(.A(new_n683), .B(new_n682), .Y(new_n684));
  nor_5  g0369(.A(new_n684), .B(new_n681), .Y(new_n685));
  nor_5  g0370(.A(pi149), .B(pi131), .Y(new_n686));
  nor_5  g0371(.A(pi201), .B(pi156), .Y(new_n687));
  or_6   g0372(.A(new_n687), .B(new_n686), .Y(new_n688));
  nor_5  g0373(.A(new_n688), .B(new_n685), .Y(new_n689));
  nand_5 g0374(.A(pi189), .B(pi113), .Y(new_n690));
  nand_5 g0375(.A(pi201), .B(pi156), .Y(new_n691));
  nand_5 g0376(.A(new_n691), .B(new_n690), .Y(new_n692));
  nor_5  g0377(.A(new_n692), .B(new_n689), .Y(new_n693));
  nor_5  g0378(.A(pi166), .B(pi094), .Y(new_n694));
  nor_5  g0379(.A(pi189), .B(pi113), .Y(new_n695));
  or_6   g0380(.A(new_n695), .B(new_n694), .Y(new_n696));
  nor_5  g0381(.A(new_n696), .B(new_n693), .Y(new_n697));
  nand_5 g0382(.A(pi142), .B(pi138), .Y(new_n698));
  nand_5 g0383(.A(pi166), .B(pi094), .Y(new_n699));
  nand_5 g0384(.A(new_n699), .B(new_n698), .Y(new_n700));
  nor_5  g0385(.A(new_n700), .B(new_n697), .Y(new_n701));
  nor_5  g0386(.A(pi142), .B(pi138), .Y(new_n702));
  nor_5  g0387(.A(pi179), .B(pi086), .Y(new_n703));
  or_6   g0388(.A(new_n703), .B(new_n702), .Y(new_n704));
  nor_5  g0389(.A(new_n704), .B(new_n701), .Y(new_n705));
  nand_5 g0390(.A(pi146), .B(pi016), .Y(new_n706));
  nand_5 g0391(.A(pi179), .B(pi086), .Y(new_n707));
  nand_5 g0392(.A(new_n707), .B(new_n706), .Y(new_n708));
  nor_5  g0393(.A(new_n708), .B(new_n705), .Y(new_n709));
  nor_5  g0394(.A(pi139), .B(pi068), .Y(new_n710));
  nor_5  g0395(.A(pi146), .B(pi016), .Y(new_n711));
  or_6   g0396(.A(new_n711), .B(new_n710), .Y(new_n712));
  nor_5  g0397(.A(new_n712), .B(new_n709), .Y(new_n713));
  nand_5 g0398(.A(pi139), .B(pi068), .Y(new_n714));
  nand_5 g0399(.A(new_n714), .B(new_n319), .Y(new_n715));
  nor_5  g0400(.A(new_n715), .B(new_n713), .Y(new_n716));
  nand_5 g0401(.A(new_n716), .B(new_n367), .Y(new_n717));
  and_6  g0402(.A(new_n717), .B(pi104), .Y(new_n718));
  nor_5  g0403(.A(new_n716), .B(new_n369), .Y(new_n719));
  nor_5  g0404(.A(new_n719), .B(new_n718), .Y(new_n720));
  nor_5  g0405(.A(new_n720), .B(new_n647), .Y(po084));
  nand_5 g0406(.A(pi150), .B(pi082), .Y(new_n722));
  nor_5  g0407(.A(new_n722), .B(pi162), .Y(new_n723));
  not_3  g0408(.A(pi121), .Y(new_n724));
  nor_5  g0409(.A(new_n361), .B(new_n724), .Y(new_n725));
  or_6   g0410(.A(new_n725), .B(new_n723), .Y(new_n726));
  or_6   g0411(.A(new_n726), .B(po084), .Y(new_n727));
  nor_5  g0412(.A(new_n354), .B(pi174), .Y(new_n728));
  nor_5  g0413(.A(new_n360), .B(pi082), .Y(new_n729));
  or_6   g0414(.A(new_n729), .B(new_n728), .Y(new_n730));
  nand_5 g0415(.A(new_n730), .B(pi150), .Y(new_n731));
  nand_5 g0416(.A(new_n319), .B(new_n724), .Y(new_n732));
  or_6   g0417(.A(new_n732), .B(pi151), .Y(new_n733));
  and_6  g0418(.A(new_n733), .B(new_n731), .Y(new_n734));
  nand_5 g0419(.A(new_n734), .B(new_n727), .Y(new_n735));
  and_6  g0420(.A(new_n735), .B(new_n574), .Y(new_n736));
  nor_5  g0421(.A(pi088), .B(pi073), .Y(new_n737));
  nor_5  g0422(.A(pi141), .B(pi112), .Y(new_n738));
  nand_5 g0423(.A(new_n738), .B(new_n737), .Y(new_n739));
  nor_5  g0424(.A(pi065), .B(pi003), .Y(new_n740));
  or_6   g0425(.A(pi019), .B(pi010), .Y(new_n741));
  nor_5  g0426(.A(new_n741), .B(new_n554), .Y(new_n742));
  nand_5 g0427(.A(new_n742), .B(new_n740), .Y(new_n743));
  nor_5  g0428(.A(new_n743), .B(new_n739), .Y(new_n744));
  not_3  g0429(.A(pi204), .Y(new_n745));
  nor_5  g0430(.A(pi101), .B(pi085), .Y(new_n746));
  nand_5 g0431(.A(new_n746), .B(new_n745), .Y(new_n747));
  not_3  g0432(.A(pi050), .Y(new_n748));
  nand_5 g0433(.A(new_n316), .B(new_n748), .Y(new_n749));
  not_3  g0434(.A(pi018), .Y(new_n750));
  nand_5 g0435(.A(new_n536), .B(new_n750), .Y(new_n751));
  or_6   g0436(.A(new_n751), .B(new_n749), .Y(new_n752));
  or_6   g0437(.A(new_n752), .B(new_n747), .Y(new_n753));
  not_3  g0438(.A(pi101), .Y(new_n754));
  nor_5  g0439(.A(pi159), .B(new_n754), .Y(new_n755));
  nor_5  g0440(.A(new_n750), .B(pi013), .Y(new_n756));
  nor_5  g0441(.A(new_n756), .B(new_n755), .Y(new_n757));
  nor_5  g0442(.A(new_n316), .B(pi095), .Y(new_n758));
  nor_5  g0443(.A(new_n758), .B(new_n318), .Y(new_n759));
  nand_5 g0444(.A(new_n759), .B(new_n757), .Y(new_n760));
  nand_5 g0445(.A(new_n760), .B(new_n753), .Y(new_n761));
  or_6   g0446(.A(new_n748), .B(pi015), .Y(new_n762));
  nand_5 g0447(.A(new_n762), .B(pi150), .Y(new_n763));
  not_3  g0448(.A(pi085), .Y(new_n764));
  nor_5  g0449(.A(pi185), .B(new_n764), .Y(new_n765));
  nor_5  g0450(.A(pi105), .B(new_n536), .Y(new_n766));
  or_6   g0451(.A(new_n766), .B(new_n765), .Y(new_n767));
  nor_5  g0452(.A(new_n767), .B(new_n763), .Y(new_n768));
  nand_5 g0453(.A(new_n768), .B(new_n761), .Y(new_n769));
  nand_5 g0454(.A(new_n319), .B(pi141), .Y(new_n770));
  nand_5 g0455(.A(pi065), .B(pi003), .Y(new_n771));
  nor_5  g0456(.A(new_n771), .B(new_n770), .Y(new_n772));
  nand_5 g0457(.A(pi088), .B(pi019), .Y(new_n773));
  nand_5 g0458(.A(pi112), .B(pi073), .Y(new_n774));
  nor_5  g0459(.A(new_n774), .B(new_n773), .Y(new_n775));
  nand_5 g0460(.A(new_n775), .B(new_n772), .Y(new_n776));
  nand_5 g0461(.A(new_n776), .B(new_n769), .Y(new_n777));
  nor_5  g0462(.A(new_n319), .B(pi047), .Y(new_n778));
  or_6   g0463(.A(new_n778), .B(new_n564), .Y(new_n779));
  and_6  g0464(.A(new_n779), .B(new_n331), .Y(new_n780));
  not_3  g0465(.A(pi190), .Y(new_n781));
  nand_5 g0466(.A(new_n319), .B(pi010), .Y(new_n782));
  nor_5  g0467(.A(new_n782), .B(new_n781), .Y(new_n783));
  nor_5  g0468(.A(pi110), .B(new_n336), .Y(new_n784));
  nand_5 g0469(.A(new_n317), .B(pi084), .Y(new_n785));
  nor_5  g0470(.A(new_n785), .B(new_n784), .Y(new_n786));
  or_6   g0471(.A(new_n786), .B(new_n783), .Y(new_n787));
  or_6   g0472(.A(new_n787), .B(new_n780), .Y(new_n788));
  and_6  g0473(.A(new_n788), .B(new_n777), .Y(new_n789));
  or_6   g0474(.A(new_n789), .B(new_n744), .Y(new_n790));
  nor_5  g0475(.A(new_n566), .B(pi119), .Y(new_n791));
  nor_5  g0476(.A(new_n348), .B(pi006), .Y(new_n792));
  nor_5  g0477(.A(new_n792), .B(new_n791), .Y(new_n793));
  nor_5  g0478(.A(new_n793), .B(new_n569), .Y(new_n794));
  not_3  g0479(.A(pi161), .Y(new_n795));
  and_6  g0480(.A(new_n341), .B(new_n795), .Y(new_n796));
  nor_5  g0481(.A(pi177), .B(pi173), .Y(new_n797));
  nor_5  g0482(.A(pi203), .B(pi140), .Y(new_n798));
  or_6   g0483(.A(new_n798), .B(new_n797), .Y(new_n799));
  and_6  g0484(.A(new_n799), .B(new_n562), .Y(new_n800));
  or_6   g0485(.A(new_n800), .B(new_n796), .Y(new_n801));
  nor_5  g0486(.A(new_n801), .B(new_n794), .Y(new_n802));
  nand_5 g0487(.A(new_n802), .B(new_n790), .Y(new_n803));
  or_6   g0488(.A(new_n803), .B(new_n736), .Y(new_n804));
  nand_5 g0489(.A(new_n744), .B(pi190), .Y(new_n805));
  nand_5 g0490(.A(new_n331), .B(pi084), .Y(new_n806));
  nand_5 g0491(.A(pi105), .B(new_n536), .Y(new_n807));
  nand_5 g0492(.A(new_n807), .B(new_n806), .Y(new_n808));
  nand_5 g0493(.A(new_n808), .B(new_n777), .Y(new_n809));
  nand_5 g0494(.A(new_n748), .B(pi015), .Y(new_n810));
  nor_5  g0495(.A(new_n810), .B(new_n758), .Y(new_n811));
  nand_5 g0496(.A(new_n316), .B(pi095), .Y(new_n812));
  nand_5 g0497(.A(new_n812), .B(pi204), .Y(new_n813));
  nor_5  g0498(.A(new_n813), .B(new_n811), .Y(new_n814));
  nor_5  g0499(.A(new_n814), .B(new_n765), .Y(new_n815));
  nand_5 g0500(.A(pi159), .B(new_n754), .Y(new_n816));
  nand_5 g0501(.A(pi185), .B(new_n764), .Y(new_n817));
  nand_5 g0502(.A(new_n817), .B(new_n816), .Y(new_n818));
  or_6   g0503(.A(new_n818), .B(new_n815), .Y(new_n819));
  and_6  g0504(.A(new_n819), .B(new_n757), .Y(new_n820));
  nand_5 g0505(.A(new_n750), .B(pi013), .Y(new_n821));
  nand_5 g0506(.A(new_n555), .B(new_n552), .Y(new_n822));
  nand_5 g0507(.A(new_n822), .B(new_n821), .Y(new_n823));
  nor_5  g0508(.A(new_n823), .B(new_n820), .Y(new_n824));
  or_6   g0509(.A(new_n824), .B(new_n744), .Y(new_n825));
  nand_5 g0510(.A(new_n825), .B(new_n809), .Y(new_n826));
  nand_5 g0511(.A(new_n826), .B(new_n317), .Y(new_n827));
  and_6  g0512(.A(new_n827), .B(new_n805), .Y(new_n828));
  and_6  g0513(.A(new_n828), .B(new_n804), .Y(new_n829));
  or_6   g0514(.A(new_n829), .B(new_n557), .Y(new_n830));
  or_6   g0515(.A(pi078), .B(pi071), .Y(new_n831));
  not_3  g0516(.A(new_n831), .Y(new_n832));
  nand_5 g0517(.A(new_n832), .B(pi022), .Y(new_n833));
  nand_5 g0518(.A(new_n833), .B(pi124), .Y(new_n834));
  and_6  g0519(.A(new_n834), .B(new_n830), .Y(new_n835));
  nand_5 g0520(.A(pi078), .B(pi071), .Y(new_n836));
  not_3  g0521(.A(new_n836), .Y(new_n837));
  not_3  g0522(.A(pi124), .Y(new_n838));
  nand_5 g0523(.A(new_n838), .B(pi022), .Y(new_n839));
  nor_5  g0524(.A(new_n839), .B(new_n837), .Y(new_n840));
  nor_5  g0525(.A(new_n840), .B(new_n835), .Y(po008));
  xor_4  g0526(.A(new_n531), .B(new_n340), .Y(po009));
  xor_4  g0527(.A(new_n533), .B(new_n335), .Y(po011));
  or_6   g0528(.A(new_n319), .B(pi062), .Y(new_n844));
  nand_5 g0529(.A(new_n844), .B(new_n317), .Y(new_n845));
  xor_4  g0530(.A(new_n845), .B(pi101), .Y(new_n846));
  not_3  g0531(.A(pi145), .Y(new_n847));
  nand_5 g0532(.A(pi150), .B(new_n847), .Y(new_n848));
  nand_5 g0533(.A(new_n848), .B(new_n317), .Y(new_n849));
  and_6  g0534(.A(new_n849), .B(pi085), .Y(new_n850));
  xor_4  g0535(.A(new_n849), .B(pi085), .Y(new_n851));
  not_3  g0536(.A(new_n851), .Y(new_n852));
  nor_5  g0537(.A(new_n321), .B(new_n316), .Y(new_n853));
  not_3  g0538(.A(new_n322), .Y(new_n854));
  nor_5  g0539(.A(new_n543), .B(new_n854), .Y(new_n855));
  nor_5  g0540(.A(new_n855), .B(new_n853), .Y(new_n856));
  nor_5  g0541(.A(new_n856), .B(new_n745), .Y(new_n857));
  not_3  g0542(.A(pi061), .Y(new_n858));
  nand_5 g0543(.A(pi150), .B(new_n858), .Y(new_n859));
  nand_5 g0544(.A(new_n859), .B(new_n317), .Y(new_n860));
  not_3  g0545(.A(new_n860), .Y(new_n861));
  xor_4  g0546(.A(new_n856), .B(pi204), .Y(new_n862));
  nor_5  g0547(.A(new_n862), .B(new_n861), .Y(new_n863));
  nor_5  g0548(.A(new_n863), .B(new_n857), .Y(new_n864));
  nor_5  g0549(.A(new_n864), .B(new_n852), .Y(new_n865));
  nor_5  g0550(.A(new_n865), .B(new_n850), .Y(new_n866));
  xor_4  g0551(.A(new_n866), .B(new_n846), .Y(po013));
  xor_4  g0552(.A(pi132), .B(pi051), .Y(new_n868));
  xor_4  g0553(.A(pi180), .B(pi083), .Y(new_n869));
  xor_4  g0554(.A(new_n869), .B(pi092), .Y(new_n870));
  xor_4  g0555(.A(new_n870), .B(new_n868), .Y(new_n871));
  and_6  g0556(.A(new_n485), .B(new_n423), .Y(new_n872));
  or_6   g0557(.A(new_n491), .B(new_n872), .Y(new_n873));
  xor_4  g0558(.A(new_n873), .B(new_n871), .Y(new_n874));
  nor_5  g0559(.A(new_n448), .B(new_n445), .Y(new_n875));
  or_6   g0560(.A(new_n875), .B(new_n465), .Y(new_n876));
  nand_5 g0561(.A(new_n465), .B(new_n449), .Y(new_n877));
  nand_5 g0562(.A(new_n877), .B(new_n876), .Y(new_n878));
  nor_5  g0563(.A(new_n433), .B(new_n430), .Y(new_n879));
  and_6  g0564(.A(new_n879), .B(new_n439), .Y(new_n880));
  nor_5  g0565(.A(new_n439), .B(new_n434), .Y(new_n881));
  nor_5  g0566(.A(new_n881), .B(new_n880), .Y(new_n882));
  nor_5  g0567(.A(new_n882), .B(new_n474), .Y(new_n883));
  nand_5 g0568(.A(new_n476), .B(new_n434), .Y(new_n884));
  or_6   g0569(.A(new_n879), .B(new_n476), .Y(new_n885));
  nand_5 g0570(.A(new_n885), .B(new_n884), .Y(new_n886));
  and_6  g0571(.A(new_n886), .B(new_n474), .Y(new_n887));
  nor_5  g0572(.A(new_n887), .B(new_n883), .Y(new_n888));
  xor_4  g0573(.A(pi043), .B(pi035), .Y(new_n889));
  xnor_4 g0574(.A(pi169), .B(pi087), .Y(new_n890));
  xor_4  g0575(.A(pi197), .B(pi193), .Y(new_n891));
  xor_4  g0576(.A(new_n891), .B(new_n890), .Y(new_n892));
  xor_4  g0577(.A(new_n892), .B(new_n889), .Y(new_n893));
  nand_5 g0578(.A(new_n893), .B(pi150), .Y(new_n894));
  xor_4  g0579(.A(pi152), .B(pi014), .Y(new_n895));
  xnor_4 g0580(.A(pi069), .B(pi033), .Y(new_n896));
  xor_4  g0581(.A(new_n896), .B(pi007), .Y(new_n897));
  xor_4  g0582(.A(new_n897), .B(new_n895), .Y(new_n898));
  xor_4  g0583(.A(pi143), .B(pi081), .Y(new_n899));
  xor_4  g0584(.A(new_n899), .B(new_n898), .Y(new_n900));
  and_6  g0585(.A(new_n456), .B(new_n455), .Y(new_n901));
  or_6   g0586(.A(new_n901), .B(new_n457), .Y(new_n902));
  xor_4  g0587(.A(new_n902), .B(new_n900), .Y(new_n903));
  nand_5 g0588(.A(new_n903), .B(new_n319), .Y(new_n904));
  nand_5 g0589(.A(new_n904), .B(new_n894), .Y(new_n905));
  xor_4  g0590(.A(new_n905), .B(new_n888), .Y(new_n906));
  xor_4  g0591(.A(new_n906), .B(new_n878), .Y(new_n907));
  xor_4  g0592(.A(new_n907), .B(new_n874), .Y(po015));
  xnor_4 g0593(.A(new_n510), .B(new_n507), .Y(po016));
  not_3  g0594(.A(pi125), .Y(po017));
  and_6  g0595(.A(pi109), .B(pi060), .Y(po020));
  not_3  g0596(.A(new_n539), .Y(new_n912));
  xor_4  g0597(.A(new_n541), .B(new_n912), .Y(po024));
  xor_4  g0598(.A(new_n512), .B(new_n397), .Y(po025));
  or_6   g0599(.A(new_n319), .B(pi077), .Y(new_n915));
  nand_5 g0600(.A(new_n915), .B(new_n317), .Y(new_n916));
  nand_5 g0601(.A(new_n916), .B(pi181), .Y(new_n917));
  and_6  g0602(.A(new_n845), .B(pi101), .Y(new_n918));
  not_3  g0603(.A(new_n846), .Y(new_n919));
  nor_5  g0604(.A(new_n866), .B(new_n919), .Y(new_n920));
  nor_5  g0605(.A(new_n920), .B(new_n918), .Y(new_n921));
  and_6  g0606(.A(new_n921), .B(new_n750), .Y(new_n922));
  or_6   g0607(.A(pi184), .B(new_n319), .Y(new_n923));
  nand_5 g0608(.A(new_n923), .B(new_n317), .Y(new_n924));
  xor_4  g0609(.A(new_n921), .B(pi018), .Y(new_n925));
  nor_5  g0610(.A(new_n925), .B(new_n924), .Y(new_n926));
  nor_5  g0611(.A(new_n926), .B(new_n922), .Y(new_n927));
  xor_4  g0612(.A(new_n916), .B(pi181), .Y(new_n928));
  nand_5 g0613(.A(new_n928), .B(new_n927), .Y(new_n929));
  nand_5 g0614(.A(new_n929), .B(new_n917), .Y(new_n930));
  xor_4  g0615(.A(new_n930), .B(new_n838), .Y(new_n931));
  nand_5 g0616(.A(pi064), .B(pi022), .Y(new_n932));
  nor_5  g0617(.A(new_n932), .B(new_n931), .Y(new_n933));
  nand_5 g0618(.A(new_n930), .B(pi124), .Y(new_n934));
  and_6  g0619(.A(pi064), .B(pi024), .Y(new_n935));
  nor_5  g0620(.A(pi064), .B(pi024), .Y(new_n936));
  nor_5  g0621(.A(new_n936), .B(new_n935), .Y(new_n937));
  nand_5 g0622(.A(new_n937), .B(pi022), .Y(new_n938));
  nor_5  g0623(.A(new_n938), .B(new_n934), .Y(new_n939));
  nor_5  g0624(.A(new_n930), .B(pi124), .Y(new_n940));
  and_6  g0625(.A(new_n938), .B(new_n940), .Y(new_n941));
  or_6   g0626(.A(new_n941), .B(new_n939), .Y(new_n942));
  nor_5  g0627(.A(new_n942), .B(new_n933), .Y(po029));
  nor_5  g0628(.A(new_n921), .B(new_n750), .Y(new_n944));
  or_6   g0629(.A(new_n926), .B(new_n944), .Y(new_n945));
  nand_5 g0630(.A(new_n856), .B(new_n745), .Y(new_n946));
  nand_5 g0631(.A(new_n946), .B(new_n852), .Y(new_n947));
  xor_4  g0632(.A(new_n947), .B(new_n945), .Y(new_n948));
  xor_4  g0633(.A(new_n948), .B(po029), .Y(new_n949));
  xor_4  g0634(.A(pi181), .B(pi101), .Y(new_n950));
  xor_4  g0635(.A(pi184), .B(pi077), .Y(new_n951));
  xor_4  g0636(.A(new_n951), .B(pi062), .Y(new_n952));
  nand_5 g0637(.A(pi145), .B(pi061), .Y(new_n953));
  nand_5 g0638(.A(new_n847), .B(new_n858), .Y(new_n954));
  nand_5 g0639(.A(new_n954), .B(new_n764), .Y(new_n955));
  nand_5 g0640(.A(new_n955), .B(new_n953), .Y(new_n956));
  nor_5  g0641(.A(new_n956), .B(new_n952), .Y(new_n957));
  nand_5 g0642(.A(new_n956), .B(new_n952), .Y(new_n958));
  nand_5 g0643(.A(new_n317), .B(pi150), .Y(new_n959));
  not_3  g0644(.A(new_n959), .Y(new_n960));
  nand_5 g0645(.A(new_n960), .B(new_n958), .Y(new_n961));
  nor_5  g0646(.A(new_n961), .B(new_n957), .Y(new_n962));
  nand_5 g0647(.A(new_n861), .B(new_n852), .Y(new_n963));
  nand_5 g0648(.A(new_n963), .B(new_n862), .Y(new_n964));
  xor_4  g0649(.A(new_n964), .B(new_n962), .Y(new_n965));
  xor_4  g0650(.A(new_n965), .B(new_n950), .Y(new_n966));
  nand_5 g0651(.A(pi024), .B(pi022), .Y(new_n967));
  xor_4  g0652(.A(new_n967), .B(new_n931), .Y(po030));
  xor_4  g0653(.A(po030), .B(new_n966), .Y(new_n969));
  xor_4  g0654(.A(new_n969), .B(new_n949), .Y(po026));
  xnor_4 g0655(.A(new_n537), .B(new_n535), .Y(po027));
  xor_4  g0656(.A(new_n521), .B(new_n373), .Y(po038));
  xor_4  g0657(.A(new_n527), .B(new_n353), .Y(po039));
  nand_5 g0658(.A(new_n935), .B(pi022), .Y(new_n974));
  nand_5 g0659(.A(new_n974), .B(pi124), .Y(new_n975));
  and_6  g0660(.A(new_n975), .B(new_n930), .Y(new_n976));
  nor_5  g0661(.A(new_n936), .B(new_n839), .Y(new_n977));
  nor_5  g0662(.A(new_n977), .B(new_n976), .Y(po040));
  xor_4  g0663(.A(new_n459), .B(new_n455), .Y(po043));
  xnor_4 g0664(.A(new_n499), .B(new_n498), .Y(po069));
  and_6  g0665(.A(new_n505), .B(new_n399), .Y(new_n981));
  nor_5  g0666(.A(new_n511), .B(new_n981), .Y(new_n982));
  xor_4  g0667(.A(new_n982), .B(po069), .Y(new_n983));
  xor_4  g0668(.A(new_n983), .B(po005), .Y(new_n984));
  nor_5  g0669(.A(new_n517), .B(new_n386), .Y(new_n985));
  not_3  g0670(.A(new_n385), .Y(new_n986));
  and_6  g0671(.A(new_n517), .B(new_n986), .Y(new_n987));
  nor_5  g0672(.A(new_n987), .B(new_n985), .Y(new_n988));
  nand_5 g0673(.A(pi189), .B(pi139), .Y(new_n989));
  nand_5 g0674(.A(new_n401), .B(new_n375), .Y(new_n990));
  nand_5 g0675(.A(new_n990), .B(new_n989), .Y(new_n991));
  nand_5 g0676(.A(new_n991), .B(new_n402), .Y(new_n992));
  xor_4  g0677(.A(pi142), .B(pi094), .Y(new_n993));
  nor_5  g0678(.A(new_n993), .B(pi150), .Y(new_n994));
  xor_4  g0679(.A(pi187), .B(pi090), .Y(new_n995));
  not_3  g0680(.A(new_n995), .Y(new_n996));
  and_6  g0681(.A(new_n996), .B(pi032), .Y(new_n997));
  or_6   g0682(.A(new_n996), .B(pi032), .Y(new_n998));
  nand_5 g0683(.A(new_n998), .B(pi150), .Y(new_n999));
  nor_5  g0684(.A(new_n999), .B(new_n997), .Y(new_n1000));
  nor_5  g0685(.A(new_n1000), .B(new_n994), .Y(new_n1001));
  xor_4  g0686(.A(new_n1001), .B(new_n992), .Y(new_n1002));
  xor_4  g0687(.A(new_n1002), .B(new_n988), .Y(new_n1003));
  not_3  g0688(.A(new_n411), .Y(new_n1004));
  and_6  g0689(.A(new_n501), .B(new_n1004), .Y(new_n1005));
  nor_5  g0690(.A(new_n501), .B(new_n412), .Y(new_n1006));
  or_6   g0691(.A(new_n1006), .B(new_n1005), .Y(new_n1007));
  xor_4  g0692(.A(pi192), .B(pi107), .Y(new_n1008));
  xor_4  g0693(.A(new_n1008), .B(pi057), .Y(new_n1009));
  xor_4  g0694(.A(new_n1009), .B(new_n1007), .Y(new_n1010));
  xor_4  g0695(.A(new_n1010), .B(new_n1003), .Y(new_n1011));
  xor_4  g0696(.A(new_n1011), .B(po038), .Y(new_n1012));
  xor_4  g0697(.A(new_n1012), .B(new_n984), .Y(po044));
  nand_5 g0698(.A(pi126), .B(pi046), .Y(new_n1014));
  nand_5 g0699(.A(pi191), .B(pi176), .Y(new_n1015));
  or_6   g0700(.A(new_n1015), .B(new_n1014), .Y(po047));
  nor_5  g0701(.A(new_n1006), .B(new_n503), .Y(new_n1017));
  or_6   g0702(.A(new_n1017), .B(new_n1005), .Y(po048));
  xor_4  g0703(.A(new_n495), .B(new_n492), .Y(po049));
  or_6   g0704(.A(pi165), .B(pi148), .Y(po050));
  xor_4  g0705(.A(new_n468), .B(new_n465), .Y(po054));
  nand_5 g0706(.A(new_n529), .B(new_n347), .Y(new_n1022));
  nor_5  g0707(.A(new_n529), .B(new_n345), .Y(new_n1023));
  or_6   g0708(.A(new_n1023), .B(new_n531), .Y(new_n1024));
  nand_5 g0709(.A(new_n1024), .B(new_n1022), .Y(po057));
  xor_4  g0710(.A(new_n862), .B(new_n860), .Y(po058));
  xor_4  g0711(.A(pi028), .B(pi013), .Y(new_n1027));
  xor_4  g0712(.A(new_n1027), .B(pi008), .Y(new_n1028));
  xor_4  g0713(.A(pi159), .B(pi031), .Y(new_n1029));
  xor_4  g0714(.A(pi185), .B(pi168), .Y(new_n1030));
  xor_4  g0715(.A(new_n1030), .B(new_n1029), .Y(new_n1031));
  xor_4  g0716(.A(new_n1031), .B(new_n1028), .Y(new_n1032));
  or_6   g0717(.A(new_n1032), .B(new_n318), .Y(new_n1033));
  nand_5 g0718(.A(new_n1033), .B(pi150), .Y(new_n1034));
  xor_4  g0719(.A(pi084), .B(pi015), .Y(new_n1035));
  xor_4  g0720(.A(pi110), .B(pi105), .Y(new_n1036));
  xor_4  g0721(.A(new_n1036), .B(pi095), .Y(new_n1037));
  nand_5 g0722(.A(new_n1037), .B(new_n1035), .Y(new_n1038));
  nor_5  g0723(.A(new_n1037), .B(new_n1035), .Y(new_n1039));
  nor_5  g0724(.A(new_n1039), .B(new_n318), .Y(new_n1040));
  nand_5 g0725(.A(new_n1040), .B(new_n1038), .Y(new_n1041));
  xor_4  g0726(.A(pi082), .B(pi006), .Y(new_n1042));
  xor_4  g0727(.A(new_n1042), .B(pi127), .Y(new_n1043));
  xor_4  g0728(.A(pi174), .B(pi119), .Y(new_n1044));
  xor_4  g0729(.A(new_n1044), .B(new_n1043), .Y(new_n1045));
  xor_4  g0730(.A(new_n1045), .B(new_n1041), .Y(new_n1046));
  or_6   g0731(.A(new_n1046), .B(new_n1034), .Y(new_n1047));
  xnor_4 g0732(.A(pi072), .B(pi052), .Y(new_n1048));
  nor_5  g0733(.A(pi195), .B(new_n624), .Y(new_n1049));
  nand_5 g0734(.A(pi195), .B(new_n624), .Y(new_n1050));
  nand_5 g0735(.A(new_n1050), .B(pi150), .Y(new_n1051));
  nor_5  g0736(.A(new_n1051), .B(new_n1049), .Y(new_n1052));
  nor_5  g0737(.A(new_n1052), .B(new_n994), .Y(new_n1053));
  nand_5 g0738(.A(pi036), .B(pi011), .Y(new_n1054));
  nor_5  g0739(.A(pi036), .B(pi011), .Y(new_n1055));
  nor_5  g0740(.A(new_n1055), .B(new_n319), .Y(new_n1056));
  nand_5 g0741(.A(new_n1056), .B(new_n1054), .Y(new_n1057));
  nand_5 g0742(.A(new_n1057), .B(new_n991), .Y(new_n1058));
  xor_4  g0743(.A(new_n1058), .B(new_n1053), .Y(new_n1059));
  xor_4  g0744(.A(pi156), .B(pi131), .Y(new_n1060));
  or_6   g0745(.A(new_n1060), .B(pi150), .Y(new_n1061));
  xor_4  g0746(.A(pi135), .B(new_n606), .Y(new_n1062));
  nand_5 g0747(.A(new_n1062), .B(pi150), .Y(new_n1063));
  nand_5 g0748(.A(new_n1063), .B(new_n1061), .Y(new_n1064));
  xor_4  g0749(.A(new_n1064), .B(new_n1059), .Y(new_n1065));
  xor_4  g0750(.A(pi114), .B(new_n633), .Y(new_n1066));
  nand_5 g0751(.A(new_n1066), .B(pi150), .Y(new_n1067));
  xor_4  g0752(.A(pi146), .B(pi086), .Y(new_n1068));
  or_6   g0753(.A(new_n1068), .B(pi150), .Y(new_n1069));
  nand_5 g0754(.A(new_n1069), .B(new_n1067), .Y(new_n1070));
  xor_4  g0755(.A(new_n1070), .B(new_n1065), .Y(new_n1071));
  xor_4  g0756(.A(new_n1071), .B(new_n1048), .Y(new_n1072));
  or_6   g0757(.A(new_n1072), .B(new_n1047), .Y(new_n1073));
  xor_4  g0758(.A(pi136), .B(pi034), .Y(new_n1074));
  nand_5 g0759(.A(new_n1071), .B(new_n1074), .Y(new_n1075));
  xor_4  g0760(.A(pi203), .B(pi186), .Y(new_n1076));
  xor_4  g0761(.A(new_n1076), .B(pi134), .Y(new_n1077));
  xor_4  g0762(.A(pi177), .B(pi151), .Y(new_n1078));
  xor_4  g0763(.A(new_n1078), .B(new_n317), .Y(new_n1079));
  nand_5 g0764(.A(new_n1079), .B(new_n1077), .Y(new_n1080));
  nor_5  g0765(.A(new_n1079), .B(new_n1077), .Y(new_n1081));
  nor_5  g0766(.A(new_n1081), .B(pi150), .Y(new_n1082));
  nand_5 g0767(.A(new_n1082), .B(new_n1080), .Y(new_n1083));
  nor_5  g0768(.A(new_n1071), .B(new_n1074), .Y(new_n1084));
  nor_5  g0769(.A(new_n1084), .B(new_n1083), .Y(new_n1085));
  nand_5 g0770(.A(new_n1085), .B(new_n1075), .Y(new_n1086));
  nand_5 g0771(.A(new_n1086), .B(new_n1073), .Y(new_n1087));
  nor_5  g0772(.A(pi067), .B(pi038), .Y(new_n1088));
  nand_5 g0773(.A(pi067), .B(pi038), .Y(new_n1089));
  nand_5 g0774(.A(new_n1089), .B(pi150), .Y(new_n1090));
  nor_5  g0775(.A(new_n1090), .B(new_n1088), .Y(new_n1091));
  nor_5  g0776(.A(new_n431), .B(pi081), .Y(new_n1092));
  nor_5  g0777(.A(new_n487), .B(pi042), .Y(new_n1093));
  or_6   g0778(.A(new_n1093), .B(new_n1092), .Y(new_n1094));
  nor_5  g0779(.A(new_n1094), .B(new_n1091), .Y(new_n1095));
  nand_5 g0780(.A(new_n897), .B(new_n319), .Y(new_n1096));
  xor_4  g0781(.A(pi171), .B(new_n597), .Y(new_n1097));
  nand_5 g0782(.A(new_n1097), .B(pi150), .Y(new_n1098));
  nand_5 g0783(.A(new_n1098), .B(new_n1096), .Y(new_n1099));
  xor_4  g0784(.A(new_n1099), .B(new_n1095), .Y(new_n1100));
  nor_5  g0785(.A(new_n895), .B(pi150), .Y(new_n1101));
  xor_4  g0786(.A(pi206), .B(pi103), .Y(new_n1102));
  nor_5  g0787(.A(new_n1102), .B(new_n319), .Y(new_n1103));
  nor_5  g0788(.A(new_n1103), .B(new_n1101), .Y(new_n1104));
  nand_5 g0789(.A(pi055), .B(pi002), .Y(new_n1105));
  nor_5  g0790(.A(pi055), .B(pi002), .Y(new_n1106));
  nor_5  g0791(.A(new_n1106), .B(new_n319), .Y(new_n1107));
  nand_5 g0792(.A(new_n1107), .B(new_n1105), .Y(new_n1108));
  nand_5 g0793(.A(new_n1108), .B(new_n446), .Y(new_n1109));
  xor_4  g0794(.A(pi129), .B(pi089), .Y(new_n1110));
  nand_5 g0795(.A(new_n1110), .B(pi150), .Y(new_n1111));
  nand_5 g0796(.A(pi143), .B(pi040), .Y(new_n1112));
  nor_5  g0797(.A(pi143), .B(pi040), .Y(new_n1113));
  nor_5  g0798(.A(new_n1113), .B(pi150), .Y(new_n1114));
  nand_5 g0799(.A(new_n1114), .B(new_n1112), .Y(new_n1115));
  nand_5 g0800(.A(new_n1115), .B(new_n1111), .Y(new_n1116));
  xor_4  g0801(.A(new_n1116), .B(new_n1109), .Y(new_n1117));
  xor_4  g0802(.A(new_n1117), .B(new_n1104), .Y(new_n1118));
  xor_4  g0803(.A(new_n1118), .B(new_n1100), .Y(new_n1119));
  nand_5 g0804(.A(new_n1119), .B(new_n1087), .Y(po090));
  xor_4  g0805(.A(pi112), .B(pi041), .Y(new_n1121));
  nor_5  g0806(.A(new_n837), .B(pi150), .Y(new_n1122));
  nand_5 g0807(.A(new_n1122), .B(new_n831), .Y(new_n1123));
  nand_5 g0808(.A(new_n937), .B(pi150), .Y(new_n1124));
  nand_5 g0809(.A(new_n1124), .B(new_n1123), .Y(new_n1125));
  xor_4  g0810(.A(pi108), .B(pi018), .Y(new_n1126));
  nand_5 g0811(.A(new_n1126), .B(pi150), .Y(new_n1127));
  nand_5 g0812(.A(pi163), .B(pi073), .Y(new_n1128));
  nor_5  g0813(.A(pi163), .B(pi073), .Y(new_n1129));
  nor_5  g0814(.A(new_n1129), .B(pi150), .Y(new_n1130));
  nand_5 g0815(.A(new_n1130), .B(new_n1128), .Y(new_n1131));
  nand_5 g0816(.A(new_n1131), .B(new_n1127), .Y(new_n1132));
  xor_4  g0817(.A(pi204), .B(new_n764), .Y(new_n1133));
  nor_5  g0818(.A(new_n1133), .B(new_n319), .Y(new_n1134));
  nor_5  g0819(.A(pi088), .B(pi019), .Y(new_n1135));
  nand_5 g0820(.A(new_n773), .B(new_n319), .Y(new_n1136));
  nor_5  g0821(.A(new_n1136), .B(new_n1135), .Y(new_n1137));
  nor_5  g0822(.A(new_n1137), .B(new_n1134), .Y(new_n1138));
  xor_4  g0823(.A(new_n1138), .B(new_n1132), .Y(new_n1139));
  xor_4  g0824(.A(new_n1139), .B(new_n1125), .Y(new_n1140));
  not_3  g0825(.A(new_n1140), .Y(new_n1141));
  nand_5 g0826(.A(new_n1141), .B(new_n1121), .Y(new_n1142));
  xor_4  g0827(.A(pi048), .B(pi029), .Y(new_n1143));
  xor_4  g0828(.A(new_n1143), .B(pi117), .Y(new_n1144));
  xor_4  g0829(.A(pi111), .B(pi100), .Y(new_n1145));
  xor_4  g0830(.A(new_n1145), .B(new_n1144), .Y(new_n1146));
  xnor_4 g0831(.A(pi098), .B(pi096), .Y(new_n1147));
  xor_4  g0832(.A(new_n1147), .B(pi066), .Y(new_n1148));
  xor_4  g0833(.A(pi023), .B(pi021), .Y(new_n1149));
  xor_4  g0834(.A(new_n1149), .B(new_n1148), .Y(new_n1150));
  xor_4  g0835(.A(new_n1150), .B(new_n1146), .Y(new_n1151));
  nor_5  g0836(.A(new_n1151), .B(pi150), .Y(new_n1152));
  nand_5 g0837(.A(new_n1152), .B(new_n1142), .Y(new_n1153));
  xor_4  g0838(.A(pi116), .B(pi039), .Y(new_n1154));
  nand_5 g0839(.A(new_n1154), .B(pi150), .Y(new_n1155));
  nand_5 g0840(.A(pi179), .B(pi016), .Y(new_n1156));
  nor_5  g0841(.A(pi179), .B(pi016), .Y(new_n1157));
  nor_5  g0842(.A(new_n1157), .B(pi150), .Y(new_n1158));
  nand_5 g0843(.A(new_n1158), .B(new_n1156), .Y(new_n1159));
  nand_5 g0844(.A(new_n1159), .B(new_n1155), .Y(new_n1160));
  xor_4  g0845(.A(pi160), .B(pi020), .Y(new_n1161));
  nand_5 g0846(.A(new_n1161), .B(pi150), .Y(new_n1162));
  nand_5 g0847(.A(pi201), .B(pi104), .Y(new_n1163));
  nor_5  g0848(.A(pi201), .B(pi104), .Y(new_n1164));
  nor_5  g0849(.A(new_n1164), .B(pi150), .Y(new_n1165));
  nand_5 g0850(.A(new_n1165), .B(new_n1163), .Y(new_n1166));
  nand_5 g0851(.A(new_n1166), .B(new_n1162), .Y(new_n1167));
  xor_4  g0852(.A(new_n1167), .B(new_n1160), .Y(new_n1168));
  xor_4  g0853(.A(pi183), .B(pi170), .Y(new_n1169));
  nand_5 g0854(.A(new_n1169), .B(pi150), .Y(new_n1170));
  nand_5 g0855(.A(pi166), .B(pi149), .Y(new_n1171));
  nor_5  g0856(.A(pi166), .B(pi149), .Y(new_n1172));
  nor_5  g0857(.A(new_n1172), .B(pi150), .Y(new_n1173));
  nand_5 g0858(.A(new_n1173), .B(new_n1171), .Y(new_n1174));
  nand_5 g0859(.A(new_n1174), .B(new_n1170), .Y(new_n1175));
  xor_4  g0860(.A(new_n1175), .B(new_n1168), .Y(new_n1176));
  xor_4  g0861(.A(pi113), .B(pi068), .Y(new_n1177));
  xor_4  g0862(.A(pi205), .B(pi138), .Y(new_n1178));
  xor_4  g0863(.A(new_n1178), .B(new_n1177), .Y(new_n1179));
  nand_5 g0864(.A(new_n1179), .B(new_n1176), .Y(new_n1180));
  nor_5  g0865(.A(new_n1141), .B(new_n1121), .Y(new_n1181));
  nor_5  g0866(.A(new_n1179), .B(new_n1176), .Y(new_n1182));
  nor_5  g0867(.A(new_n1182), .B(new_n1181), .Y(new_n1183));
  nand_5 g0868(.A(new_n1183), .B(new_n1180), .Y(new_n1184));
  nor_5  g0869(.A(new_n1184), .B(new_n1153), .Y(new_n1185));
  xnor_4 g0870(.A(new_n1009), .B(pi118), .Y(new_n1186));
  xor_4  g0871(.A(new_n1186), .B(new_n1176), .Y(new_n1187));
  nor_5  g0872(.A(new_n1141), .B(new_n950), .Y(new_n1188));
  nand_5 g0873(.A(new_n1141), .B(new_n950), .Y(new_n1189));
  xor_4  g0874(.A(pi074), .B(new_n445), .Y(new_n1190));
  xor_4  g0875(.A(pi147), .B(pi137), .Y(new_n1191));
  xor_4  g0876(.A(new_n1191), .B(new_n1190), .Y(new_n1192));
  xor_4  g0877(.A(new_n871), .B(new_n430), .Y(new_n1193));
  nand_5 g0878(.A(new_n1193), .B(new_n1192), .Y(new_n1194));
  nand_5 g0879(.A(new_n1194), .B(new_n1189), .Y(new_n1195));
  or_6   g0880(.A(new_n1195), .B(new_n1188), .Y(new_n1196));
  or_6   g0881(.A(new_n1193), .B(new_n1192), .Y(new_n1197));
  nand_5 g0882(.A(new_n1197), .B(pi150), .Y(new_n1198));
  or_6   g0883(.A(new_n1198), .B(new_n1196), .Y(new_n1199));
  nor_5  g0884(.A(new_n1199), .B(new_n1187), .Y(new_n1200));
  nor_5  g0885(.A(new_n1200), .B(new_n1185), .Y(new_n1201));
  xor_4  g0886(.A(pi178), .B(pi162), .Y(new_n1202));
  nand_5 g0887(.A(new_n1202), .B(pi150), .Y(new_n1203));
  nand_5 g0888(.A(pi140), .B(pi121), .Y(new_n1204));
  nor_5  g0889(.A(pi140), .B(pi121), .Y(new_n1205));
  nor_5  g0890(.A(new_n1205), .B(pi150), .Y(new_n1206));
  nand_5 g0891(.A(new_n1206), .B(new_n1204), .Y(new_n1207));
  nand_5 g0892(.A(new_n1207), .B(new_n1203), .Y(new_n1208));
  xor_4  g0893(.A(pi196), .B(pi001), .Y(new_n1209));
  nand_5 g0894(.A(new_n1209), .B(pi150), .Y(new_n1210));
  nand_5 g0895(.A(pi202), .B(pi161), .Y(new_n1211));
  nor_5  g0896(.A(pi202), .B(pi161), .Y(new_n1212));
  nor_5  g0897(.A(new_n1212), .B(pi150), .Y(new_n1213));
  nand_5 g0898(.A(new_n1213), .B(new_n1211), .Y(new_n1214));
  nand_5 g0899(.A(new_n1214), .B(new_n1210), .Y(new_n1215));
  nand_5 g0900(.A(pi141), .B(pi010), .Y(new_n1216));
  nand_5 g0901(.A(new_n782), .B(new_n770), .Y(new_n1217));
  nand_5 g0902(.A(new_n1217), .B(new_n1216), .Y(new_n1218));
  nand_5 g0903(.A(pi122), .B(pi056), .Y(new_n1219));
  nor_5  g0904(.A(pi122), .B(pi056), .Y(new_n1220));
  nor_5  g0905(.A(new_n1220), .B(new_n319), .Y(new_n1221));
  nand_5 g0906(.A(new_n1221), .B(new_n1219), .Y(new_n1222));
  nand_5 g0907(.A(new_n1222), .B(new_n1218), .Y(new_n1223));
  xor_4  g0908(.A(new_n1223), .B(new_n1215), .Y(new_n1224));
  xor_4  g0909(.A(new_n1224), .B(new_n1208), .Y(new_n1225));
  nor_5  g0910(.A(new_n316), .B(new_n748), .Y(new_n1226));
  nand_5 g0911(.A(new_n749), .B(pi150), .Y(new_n1227));
  nor_5  g0912(.A(new_n1227), .B(new_n1226), .Y(new_n1228));
  nor_5  g0913(.A(new_n740), .B(pi150), .Y(new_n1229));
  and_6  g0914(.A(new_n1229), .B(new_n771), .Y(new_n1230));
  nor_5  g0915(.A(new_n1230), .B(new_n1228), .Y(new_n1231));
  xor_4  g0916(.A(pi199), .B(pi047), .Y(new_n1232));
  nor_5  g0917(.A(new_n1232), .B(new_n319), .Y(new_n1233));
  xor_4  g0918(.A(pi190), .B(pi173), .Y(new_n1234));
  nor_5  g0919(.A(new_n1234), .B(pi150), .Y(new_n1235));
  or_6   g0920(.A(new_n1235), .B(new_n1233), .Y(new_n1236));
  xor_4  g0921(.A(new_n1236), .B(new_n1231), .Y(new_n1237));
  xor_4  g0922(.A(new_n1237), .B(new_n1225), .Y(new_n1238));
  not_3  g0923(.A(new_n1238), .Y(new_n1239));
  nor_5  g0924(.A(new_n1239), .B(new_n1201), .Y(new_n1240));
  xor_4  g0925(.A(pi058), .B(pi042), .Y(new_n1241));
  xor_4  g0926(.A(new_n1241), .B(pi040), .Y(new_n1242));
  xor_4  g0927(.A(new_n1242), .B(new_n900), .Y(new_n1243));
  nor_5  g0928(.A(new_n1243), .B(new_n1083), .Y(new_n1244));
  not_3  g0929(.A(new_n952), .Y(new_n1245));
  xor_4  g0930(.A(pi102), .B(new_n858), .Y(new_n1246));
  xor_4  g0931(.A(pi200), .B(pi145), .Y(new_n1247));
  xor_4  g0932(.A(new_n1247), .B(new_n1246), .Y(new_n1248));
  not_3  g0933(.A(new_n1248), .Y(new_n1249));
  nand_5 g0934(.A(new_n1249), .B(new_n1245), .Y(new_n1250));
  nor_5  g0935(.A(new_n1249), .B(new_n1245), .Y(new_n1251));
  nor_5  g0936(.A(new_n1251), .B(new_n318), .Y(new_n1252));
  nand_5 g0937(.A(new_n1252), .B(new_n1250), .Y(new_n1253));
  and_6  g0938(.A(new_n1253), .B(pi150), .Y(new_n1254));
  xor_4  g0939(.A(pi044), .B(pi025), .Y(new_n1255));
  xor_4  g0940(.A(pi155), .B(pi120), .Y(new_n1256));
  xor_4  g0941(.A(new_n1256), .B(new_n1255), .Y(new_n1257));
  xnor_4 g0942(.A(new_n1257), .B(new_n893), .Y(new_n1258));
  nand_5 g0943(.A(new_n1258), .B(new_n1254), .Y(new_n1259));
  xor_4  g0944(.A(pi182), .B(pi009), .Y(new_n1260));
  xor_4  g0945(.A(new_n1260), .B(pi017), .Y(new_n1261));
  xor_4  g0946(.A(pi154), .B(pi115), .Y(new_n1262));
  not_3  g0947(.A(new_n1262), .Y(new_n1263));
  xor_4  g0948(.A(pi175), .B(pi026), .Y(new_n1264));
  xor_4  g0949(.A(new_n1264), .B(pi054), .Y(new_n1265));
  not_3  g0950(.A(new_n1265), .Y(new_n1266));
  nand_5 g0951(.A(new_n1266), .B(new_n1263), .Y(new_n1267));
  nor_5  g0952(.A(new_n1266), .B(new_n1263), .Y(new_n1268));
  nor_5  g0953(.A(new_n1268), .B(new_n318), .Y(new_n1269));
  nand_5 g0954(.A(new_n1269), .B(new_n1267), .Y(new_n1270));
  xor_4  g0955(.A(pi172), .B(pi080), .Y(new_n1271));
  xor_4  g0956(.A(new_n1271), .B(new_n1270), .Y(new_n1272));
  xor_4  g0957(.A(new_n1272), .B(new_n1261), .Y(new_n1273));
  nor_5  g0958(.A(new_n1273), .B(new_n1259), .Y(new_n1274));
  nor_5  g0959(.A(new_n1274), .B(new_n1244), .Y(new_n1275));
  xor_4  g0960(.A(pi194), .B(pi164), .Y(new_n1276));
  xor_4  g0961(.A(pi158), .B(pi045), .Y(new_n1277));
  xor_4  g0962(.A(pi030), .B(pi012), .Y(new_n1278));
  xor_4  g0963(.A(new_n1278), .B(new_n1277), .Y(new_n1279));
  xor_4  g0964(.A(new_n1279), .B(new_n1276), .Y(new_n1280));
  nor_5  g0965(.A(new_n1280), .B(new_n319), .Y(new_n1281));
  xor_4  g0966(.A(new_n1068), .B(new_n1060), .Y(new_n1282));
  xor_4  g0967(.A(new_n1282), .B(new_n1074), .Y(new_n1283));
  nor_5  g0968(.A(new_n1283), .B(pi150), .Y(new_n1284));
  nor_5  g0969(.A(new_n1284), .B(new_n1281), .Y(new_n1285));
  xor_4  g0970(.A(new_n1285), .B(new_n1002), .Y(new_n1286));
  not_3  g0971(.A(new_n1286), .Y(new_n1287));
  nor_5  g0972(.A(new_n1287), .B(new_n1275), .Y(new_n1288));
  not_3  g0973(.A(new_n1288), .Y(po080));
  nor_5  g0974(.A(po047), .B(po006), .Y(new_n1290));
  nand_5 g0975(.A(pi128), .B(pi079), .Y(new_n1291));
  nand_5 g0976(.A(pi157), .B(pi130), .Y(new_n1292));
  or_6   g0977(.A(new_n1292), .B(new_n1291), .Y(po100));
  nand_5 g0978(.A(pi076), .B(pi063), .Y(new_n1294));
  nand_5 g0979(.A(pi133), .B(pi099), .Y(new_n1295));
  or_6   g0980(.A(new_n1295), .B(new_n1294), .Y(po107));
  nor_5  g0981(.A(po107), .B(po100), .Y(new_n1297));
  nand_5 g0982(.A(new_n1297), .B(new_n1290), .Y(new_n1298));
  nor_5  g0983(.A(new_n1298), .B(po080), .Y(new_n1299));
  nand_5 g0984(.A(new_n1299), .B(new_n1240), .Y(new_n1300));
  or_6   g0985(.A(new_n1300), .B(po090), .Y(po059));
  xor_4  g0986(.A(new_n503), .B(new_n405), .Y(po060));
  or_6   g0987(.A(new_n928), .B(new_n927), .Y(new_n1303));
  nand_5 g0988(.A(new_n1303), .B(new_n929), .Y(po061));
  xor_4  g0989(.A(new_n481), .B(new_n480), .Y(po062));
  nand_5 g0990(.A(pi093), .B(pi053), .Y(new_n1306));
  or_6   g0991(.A(new_n1306), .B(pi165), .Y(po065));
  nor_5  g0992(.A(new_n525), .B(new_n359), .Y(new_n1308));
  not_3  g0993(.A(new_n358), .Y(new_n1309));
  and_6  g0994(.A(new_n525), .B(new_n1309), .Y(new_n1310));
  not_3  g0995(.A(new_n1310), .Y(new_n1311));
  and_6  g0996(.A(new_n1311), .B(new_n527), .Y(new_n1312));
  nor_5  g0997(.A(new_n1312), .B(new_n1308), .Y(po066));
  xor_4  g0998(.A(new_n472), .B(new_n470), .Y(po067));
  nor_5  g0999(.A(new_n985), .B(new_n519), .Y(new_n1315));
  or_6   g1000(.A(new_n1315), .B(new_n987), .Y(po068));
  nand_5 g1001(.A(new_n540), .B(new_n539), .Y(new_n1317));
  nand_5 g1002(.A(new_n912), .B(new_n325), .Y(new_n1318));
  nand_5 g1003(.A(new_n1318), .B(new_n1317), .Y(new_n1319));
  xor_4  g1004(.A(po011), .B(new_n351), .Y(new_n1320));
  nor_5  g1005(.A(new_n1310), .B(new_n1308), .Y(new_n1321));
  xor_4  g1006(.A(new_n1321), .B(new_n1320), .Y(new_n1322));
  xor_4  g1007(.A(new_n1322), .B(new_n1319), .Y(new_n1323));
  and_6  g1008(.A(new_n529), .B(new_n347), .Y(new_n1324));
  or_6   g1009(.A(new_n1023), .B(new_n1324), .Y(new_n1325));
  xor_4  g1010(.A(new_n1325), .B(new_n1232), .Y(new_n1326));
  xor_4  g1011(.A(new_n523), .B(new_n365), .Y(po095));
  xor_4  g1012(.A(po095), .B(po027), .Y(new_n1328));
  xor_4  g1013(.A(new_n1328), .B(new_n1326), .Y(new_n1329));
  nand_5 g1014(.A(new_n1264), .B(new_n960), .Y(new_n1330));
  xor_4  g1015(.A(new_n1330), .B(pi153), .Y(new_n1331));
  xor_4  g1016(.A(new_n1331), .B(new_n1329), .Y(new_n1332));
  xor_4  g1017(.A(new_n1332), .B(new_n1323), .Y(po070));
  xnor_4 g1018(.A(new_n490), .B(new_n489), .Y(po073));
  xor_4  g1019(.A(new_n864), .B(new_n851), .Y(po083));
  not_3  g1020(.A(new_n1240), .Y(po086));
  xor_4  g1021(.A(new_n925), .B(new_n924), .Y(po091));
  xor_4  g1022(.A(new_n463), .B(new_n462), .Y(po092));
  xor_4  g1023(.A(new_n483), .B(new_n429), .Y(po094));
  xor_4  g1024(.A(new_n478), .B(new_n474), .Y(po102));
  xor_4  g1025(.A(new_n519), .B(new_n379), .Y(po104));
  buf_8  g1026(.A(pi050), .Y(po001));
  buf_8  g1027(.A(pi118), .Y(po002));
  buf_8  g1028(.A(pi020), .Y(po004));
  buf_8  g1029(.A(pi196), .Y(po007));
  buf_8  g1030(.A(pi107), .Y(po010));
  buf_8  g1031(.A(pi060), .Y(po012));
  buf_8  g1032(.A(pi108), .Y(po014));
  buf_8  g1033(.A(pi057), .Y(po018));
  buf_8  g1034(.A(pi047), .Y(po019));
  buf_8  g1035(.A(pi085), .Y(po021));
  buf_8  g1036(.A(pi180), .Y(po022));
  nand_5 g1037(.A(pi167), .B(new_n545), .Y(po023));
  buf_8  g1038(.A(pi056), .Y(po028));
  nor_5  g1039(.A(new_n840), .B(new_n835), .Y(po031));
  buf_8  g1040(.A(pi001), .Y(po032));
  buf_8  g1041(.A(pi204), .Y(po033));
  buf_8  g1042(.A(pi039), .Y(po034));
  buf_8  g1043(.A(pi024), .Y(po035));
  buf_8  g1044(.A(pi101), .Y(po036));
  buf_8  g1045(.A(pi144), .Y(po037));
  nor_5  g1046(.A(new_n977), .B(new_n976), .Y(po041));
  buf_8  g1047(.A(pi160), .Y(po042));
  buf_8  g1048(.A(pi060), .Y(po045));
  buf_8  g1049(.A(pi162), .Y(po046));
  not_3  g1050(.A(pi125), .Y(po051));
  buf_8  g1051(.A(pi122), .Y(po052));
  buf_8  g1052(.A(pi027), .Y(po053));
  buf_8  g1053(.A(pi051), .Y(po055));
  buf_8  g1054(.A(pi147), .Y(po056));
  buf_8  g1055(.A(pi183), .Y(po063));
  buf_8  g1056(.A(pi192), .Y(po064));
  buf_8  g1057(.A(pi064), .Y(po071));
  nor_5  g1058(.A(new_n977), .B(new_n976), .Y(po072));
  buf_8  g1059(.A(pi132), .Y(po074));
  nor_5  g1060(.A(new_n840), .B(new_n835), .Y(po075));
  buf_8  g1061(.A(pi181), .Y(po076));
  buf_8  g1062(.A(pi083), .Y(po077));
  or_6   g1063(.A(new_n1306), .B(pi165), .Y(po078));
  buf_8  g1064(.A(pi170), .Y(po079));
  buf_8  g1065(.A(pi199), .Y(po081));
  not_3  g1066(.A(pi125), .Y(po082));
  buf_8  g1067(.A(pi153), .Y(po085));
  buf_8  g1068(.A(pi137), .Y(po087));
  xor_4  g1069(.A(new_n967), .B(new_n931), .Y(po088));
  buf_8  g1070(.A(pi060), .Y(po089));
  buf_8  g1071(.A(pi092), .Y(po093));
  buf_8  g1072(.A(pi116), .Y(po096));
  buf_8  g1073(.A(pi060), .Y(po097));
  buf_8  g1074(.A(pi074), .Y(po098));
  nor_5  g1075(.A(new_n942), .B(new_n933), .Y(po099));
  nor_5  g1076(.A(new_n977), .B(new_n976), .Y(po101));
  buf_8  g1077(.A(pi178), .Y(po103));
  buf_8  g1078(.A(pi018), .Y(po105));
  buf_8  g1079(.A(pi004), .Y(po106));
endmodule


