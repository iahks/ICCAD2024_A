 module top_810026173_843396535_809698999_829556405_809567927 (a, b, o);

      input a, b; output o; nor_8 g0(a,b,o); endmodule