// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Sun Aug 18 20:53:50 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119;
  wire new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n386, new_n387, new_n388, new_n389, new_n390, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1875, new_n1876, new_n1877, new_n1878, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1890, new_n1891, new_n1892,
    new_n1893, new_n1894, new_n1895, new_n1896, new_n1897, new_n1898,
    new_n1899, new_n1900, new_n1901, new_n1902, new_n1903, new_n1904,
    new_n1905, new_n1906, new_n1907, new_n1908, new_n1909, new_n1910,
    new_n1911, new_n1912, new_n1913, new_n1914, new_n1915, new_n1916,
    new_n1917, new_n1918, new_n1919, new_n1920, new_n1921, new_n1922,
    new_n1923, new_n1924, new_n1925, new_n1926, new_n1927, new_n1928,
    new_n1929, new_n1930, new_n1931, new_n1932, new_n1933, new_n1934,
    new_n1935, new_n1936, new_n1937, new_n1938, new_n1939, new_n1940,
    new_n1941, new_n1942, new_n1943, new_n1944, new_n1945, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019,
    new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025,
    new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031,
    new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055,
    new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061,
    new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067,
    new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896,
    new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914,
    new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944,
    new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956,
    new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962,
    new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046,
    new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052,
    new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058,
    new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064,
    new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070,
    new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076,
    new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088,
    new_n3089, new_n3090, new_n3091, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3101, new_n3102, new_n3103, new_n3104, new_n3105, new_n3106,
    new_n3107, new_n3108, new_n3109, new_n3110, new_n3111, new_n3112,
    new_n3113, new_n3114, new_n3115, new_n3116, new_n3117, new_n3118,
    new_n3119, new_n3120, new_n3121, new_n3122, new_n3123, new_n3124,
    new_n3125, new_n3126, new_n3127, new_n3128, new_n3129, new_n3130,
    new_n3131, new_n3132, new_n3133, new_n3134, new_n3135, new_n3136,
    new_n3137, new_n3138, new_n3139, new_n3140, new_n3141, new_n3142,
    new_n3143, new_n3144, new_n3145, new_n3146, new_n3147, new_n3148,
    new_n3149, new_n3150, new_n3151, new_n3152, new_n3153, new_n3154,
    new_n3155, new_n3156, new_n3157, new_n3158, new_n3159, new_n3160,
    new_n3161, new_n3162, new_n3163, new_n3164, new_n3165, new_n3166,
    new_n3167, new_n3168, new_n3169, new_n3170, new_n3171, new_n3172,
    new_n3173, new_n3174, new_n3175, new_n3176, new_n3177, new_n3178,
    new_n3179, new_n3180, new_n3181, new_n3182, new_n3183, new_n3184,
    new_n3185, new_n3186, new_n3187, new_n3188, new_n3189, new_n3190,
    new_n3191, new_n3192, new_n3193, new_n3194, new_n3195, new_n3196,
    new_n3197, new_n3198, new_n3199, new_n3200, new_n3201, new_n3202,
    new_n3203, new_n3204, new_n3205, new_n3206, new_n3207, new_n3208,
    new_n3209, new_n3210, new_n3211, new_n3213, new_n3214, new_n3215,
    new_n3216, new_n3217, new_n3218, new_n3219, new_n3220, new_n3221,
    new_n3222, new_n3223, new_n3224, new_n3225, new_n3226, new_n3227,
    new_n3228, new_n3229, new_n3230, new_n3231, new_n3232, new_n3233,
    new_n3234, new_n3235, new_n3236, new_n3237, new_n3238, new_n3239,
    new_n3240, new_n3241, new_n3242, new_n3243, new_n3244, new_n3245,
    new_n3246, new_n3247, new_n3248, new_n3249, new_n3250, new_n3251,
    new_n3252, new_n3253, new_n3254, new_n3255, new_n3256, new_n3257,
    new_n3258, new_n3259, new_n3260, new_n3261, new_n3262, new_n3263,
    new_n3264, new_n3265, new_n3266, new_n3267, new_n3268, new_n3269,
    new_n3270, new_n3271, new_n3272, new_n3273, new_n3274, new_n3275,
    new_n3276, new_n3277, new_n3278, new_n3279, new_n3280, new_n3281,
    new_n3282, new_n3283, new_n3284, new_n3285, new_n3286, new_n3287,
    new_n3288, new_n3289, new_n3290, new_n3291, new_n3292, new_n3293,
    new_n3294, new_n3295, new_n3296, new_n3297, new_n3298, new_n3299,
    new_n3300, new_n3301, new_n3302, new_n3303, new_n3304, new_n3305,
    new_n3306, new_n3307, new_n3308, new_n3309, new_n3310, new_n3311,
    new_n3312, new_n3313, new_n3314, new_n3315, new_n3316, new_n3317,
    new_n3318, new_n3319, new_n3320, new_n3321, new_n3322, new_n3323,
    new_n3324, new_n3325, new_n3326, new_n3327, new_n3328, new_n3329,
    new_n3330, new_n3331, new_n3332, new_n3333, new_n3334, new_n3335,
    new_n3336, new_n3337, new_n3338, new_n3339, new_n3340, new_n3341,
    new_n3342, new_n3343, new_n3344, new_n3345, new_n3346, new_n3347,
    new_n3348, new_n3349, new_n3350, new_n3351, new_n3352, new_n3353,
    new_n3354, new_n3355, new_n3356, new_n3357, new_n3358, new_n3359,
    new_n3360, new_n3361, new_n3362, new_n3363, new_n3364, new_n3365,
    new_n3366, new_n3367, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516,
    new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552,
    new_n3553, new_n3554, new_n3555, new_n3556, new_n3557, new_n3558,
    new_n3559, new_n3560, new_n3561, new_n3562, new_n3563, new_n3564,
    new_n3565, new_n3566, new_n3567, new_n3568, new_n3569, new_n3570,
    new_n3571, new_n3572, new_n3573, new_n3574, new_n3575, new_n3576,
    new_n3577, new_n3578, new_n3579, new_n3580, new_n3581, new_n3582,
    new_n3583, new_n3584, new_n3585, new_n3586, new_n3587, new_n3588,
    new_n3589, new_n3590, new_n3591, new_n3592, new_n3593, new_n3594,
    new_n3595, new_n3596, new_n3597, new_n3598, new_n3599, new_n3600,
    new_n3601, new_n3602, new_n3603, new_n3604, new_n3605, new_n3606,
    new_n3608, new_n3609, new_n3610, new_n3611, new_n3612, new_n3613,
    new_n3614, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4293, new_n4294,
    new_n4295, new_n4296, new_n4297, new_n4298, new_n4299, new_n4300,
    new_n4301, new_n4302, new_n4303, new_n4304, new_n4305, new_n4306,
    new_n4307, new_n4308, new_n4309, new_n4310, new_n4311, new_n4312,
    new_n4313, new_n4314, new_n4315, new_n4316, new_n4317, new_n4318,
    new_n4319, new_n4320, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577,
    new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583,
    new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589,
    new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595,
    new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601,
    new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607,
    new_n4608, new_n4609, new_n4610, new_n4611, new_n4612, new_n4613,
    new_n4614, new_n4615, new_n4616, new_n4617, new_n4618, new_n4619,
    new_n4620, new_n4621, new_n4622, new_n4623, new_n4624, new_n4625,
    new_n4626, new_n4627, new_n4628, new_n4629, new_n4630, new_n4631,
    new_n4632, new_n4633, new_n4634, new_n4635, new_n4636, new_n4637,
    new_n4638, new_n4639, new_n4640, new_n4641, new_n4642, new_n4643,
    new_n4644, new_n4645, new_n4646, new_n4647, new_n4648, new_n4649,
    new_n4650, new_n4651, new_n4652, new_n4653, new_n4654, new_n4655,
    new_n4656, new_n4657, new_n4658, new_n4659, new_n4660, new_n4661,
    new_n4662, new_n4663, new_n4664, new_n4665, new_n4666, new_n4667,
    new_n4668, new_n4669, new_n4670, new_n4671, new_n4672, new_n4673,
    new_n4674, new_n4675, new_n4676, new_n4677, new_n4678, new_n4679,
    new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685,
    new_n4686, new_n4687, new_n4688, new_n4689, new_n4690, new_n4691,
    new_n4692, new_n4693, new_n4694, new_n4695, new_n4696, new_n4697,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4927, new_n4929, new_n4930, new_n4931, new_n4932, new_n4933,
    new_n4934, new_n4935, new_n4936, new_n4937, new_n4938, new_n4939,
    new_n4940, new_n4941, new_n4942, new_n4943, new_n4944, new_n4945,
    new_n4946, new_n4947, new_n4948, new_n4949, new_n4950, new_n4951,
    new_n4952, new_n4953, new_n4954, new_n4955, new_n4956, new_n4957,
    new_n4958, new_n4959, new_n4960, new_n4961, new_n4962, new_n4963,
    new_n4964, new_n4965, new_n4966, new_n4967, new_n4968, new_n4969,
    new_n4970, new_n4971, new_n4972, new_n4973, new_n4974, new_n4975,
    new_n4976, new_n4977, new_n4978, new_n4979, new_n4980, new_n4981,
    new_n4982, new_n4983, new_n4984, new_n4985, new_n4986, new_n4987,
    new_n4988, new_n4989, new_n4990, new_n4991, new_n4992, new_n4993,
    new_n4994, new_n4995, new_n4996, new_n4997, new_n4998, new_n4999,
    new_n5000, new_n5001, new_n5002, new_n5003, new_n5004, new_n5005,
    new_n5006, new_n5007, new_n5008, new_n5009, new_n5010, new_n5011,
    new_n5012, new_n5013, new_n5014, new_n5015, new_n5016, new_n5017,
    new_n5018, new_n5019, new_n5020, new_n5021, new_n5022, new_n5023,
    new_n5024, new_n5025, new_n5026, new_n5027, new_n5028, new_n5029,
    new_n5030, new_n5031, new_n5032, new_n5033, new_n5034, new_n5035,
    new_n5036, new_n5037, new_n5038, new_n5039, new_n5040, new_n5041,
    new_n5042, new_n5043, new_n5044, new_n5045, new_n5046, new_n5047,
    new_n5048, new_n5049, new_n5050, new_n5051, new_n5052, new_n5053,
    new_n5054, new_n5055, new_n5056, new_n5057, new_n5058, new_n5059,
    new_n5060, new_n5061, new_n5062, new_n5063, new_n5064, new_n5065,
    new_n5066, new_n5067, new_n5068, new_n5069, new_n5070, new_n5071,
    new_n5072, new_n5074, new_n5075, new_n5076, new_n5077, new_n5078,
    new_n5079, new_n5080, new_n5081, new_n5082, new_n5083, new_n5084,
    new_n5085, new_n5086, new_n5087, new_n5088, new_n5089, new_n5090,
    new_n5091, new_n5092, new_n5093, new_n5094, new_n5095, new_n5096,
    new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102,
    new_n5103, new_n5104, new_n5105, new_n5106, new_n5107, new_n5108,
    new_n5109, new_n5110, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523,
    new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559,
    new_n6560, new_n6561, new_n6562, new_n6563, new_n6564, new_n6565,
    new_n6566, new_n6567, new_n6568, new_n6569, new_n6570, new_n6571,
    new_n6572, new_n6573, new_n6574, new_n6575, new_n6576, new_n6577,
    new_n6578, new_n6579, new_n6580, new_n6581, new_n6582, new_n6583,
    new_n6584, new_n6585, new_n6586, new_n6587, new_n6588, new_n6589,
    new_n6590, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595,
    new_n6596, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601,
    new_n6602, new_n6603, new_n6604, new_n6605, new_n6606, new_n6607,
    new_n6608, new_n6609, new_n6610, new_n6611, new_n6612, new_n6613,
    new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619,
    new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6625,
    new_n6626, new_n6627, new_n6628, new_n6629, new_n6630, new_n6631,
    new_n6632, new_n6633, new_n6634, new_n6635, new_n6636, new_n6637,
    new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643,
    new_n6644, new_n6645, new_n6646, new_n6647, new_n6648, new_n6649,
    new_n6653, new_n6654, new_n6655, new_n6656, new_n6657, new_n6658,
    new_n6659, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672,
    new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684,
    new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690,
    new_n6691, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6717, new_n6718, new_n6719, new_n6720,
    new_n6721, new_n6722, new_n6723, new_n6724, new_n6725, new_n6726,
    new_n6727, new_n6728, new_n6729, new_n6730, new_n6731, new_n6732,
    new_n6733, new_n6734, new_n6735, new_n6736, new_n6737, new_n6738,
    new_n6739, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229, new_n7230, new_n7231, new_n7232, new_n7233,
    new_n7234, new_n7235, new_n7236, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253, new_n7254, new_n7255, new_n7256, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7265, new_n7266, new_n7267, new_n7268, new_n7269,
    new_n7270, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275,
    new_n7276, new_n7277, new_n7278, new_n7279, new_n7280, new_n7281,
    new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287,
    new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293,
    new_n7294, new_n7295, new_n7296, new_n7297, new_n7298, new_n7299,
    new_n7300, new_n7301, new_n7302, new_n7303, new_n7304, new_n7305,
    new_n7306, new_n7307, new_n7308, new_n7309, new_n7310, new_n7311,
    new_n7312, new_n7313, new_n7314, new_n7315, new_n7316, new_n7317,
    new_n7318, new_n7319, new_n7320, new_n7321, new_n7322, new_n7323,
    new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329,
    new_n7330, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335,
    new_n7336, new_n7337, new_n7338, new_n7339, new_n7340, new_n7341,
    new_n7342, new_n7343, new_n7344, new_n7345, new_n7346, new_n7347,
    new_n7348, new_n7349, new_n7350, new_n7351, new_n7352, new_n7353,
    new_n7354, new_n7355, new_n7356, new_n7357, new_n7358, new_n7359,
    new_n7360, new_n7361, new_n7362, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052,
    new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058,
    new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064,
    new_n8065, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070,
    new_n8071, new_n8072, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819,
    new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825,
    new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528,
    new_n9529, new_n9530, new_n9531, new_n9532, new_n9533, new_n9534,
    new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540,
    new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546,
    new_n9547, new_n9548, new_n9549, new_n9550, new_n9560, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763, new_n9764, new_n9765, new_n9766, new_n9767,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865,
    new_n9866, new_n9867, new_n9868, new_n9869, new_n9870, new_n9871,
    new_n9872, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877,
    new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883,
    new_n9884, new_n9885, new_n9886, new_n9887, new_n9888, new_n9889,
    new_n9890, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895,
    new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901,
    new_n9902, new_n9903, new_n9904, new_n9905, new_n9906, new_n9907,
    new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915, new_n9916, new_n9917, new_n9918, new_n9919,
    new_n9920, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937,
    new_n9938, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997,
    new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003,
    new_n10004, new_n10005, new_n10006, new_n10007, new_n10008, new_n10009,
    new_n10010, new_n10011, new_n10012, new_n10013, new_n10014, new_n10015,
    new_n10016, new_n10017, new_n10018, new_n10019, new_n10020, new_n10021,
    new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035,
    new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041,
    new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047,
    new_n10048, new_n10049, new_n10050, new_n10051, new_n10052, new_n10053,
    new_n10054, new_n10055, new_n10056, new_n10057, new_n10058, new_n10059,
    new_n10060, new_n10061, new_n10062, new_n10063, new_n10064, new_n10065,
    new_n10066, new_n10067, new_n10068, new_n10069, new_n10070, new_n10071,
    new_n10072, new_n10073, new_n10074, new_n10075, new_n10076, new_n10077,
    new_n10078, new_n10079, new_n10080, new_n10081, new_n10082, new_n10083,
    new_n10084, new_n10085, new_n10086, new_n10087, new_n10088, new_n10089,
    new_n10090, new_n10091, new_n10092, new_n10093, new_n10094, new_n10095,
    new_n10096, new_n10097, new_n10098, new_n10099, new_n10100, new_n10101,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111, new_n10112, new_n10113,
    new_n10114, new_n10115, new_n10116, new_n10117, new_n10118, new_n10119,
    new_n10120, new_n10121, new_n10122, new_n10123, new_n10124, new_n10125,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10133, new_n10134, new_n10135, new_n10136, new_n10137,
    new_n10138, new_n10139, new_n10140, new_n10141, new_n10142, new_n10143,
    new_n10144, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158, new_n10159, new_n10160, new_n10161,
    new_n10162, new_n10163, new_n10164, new_n10165, new_n10166, new_n10167,
    new_n10168, new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174, new_n10175, new_n10176, new_n10177, new_n10178, new_n10179,
    new_n10180, new_n10181, new_n10182, new_n10183, new_n10184, new_n10185,
    new_n10186, new_n10187, new_n10188, new_n10189, new_n10190, new_n10191,
    new_n10192, new_n10193, new_n10194, new_n10195, new_n10196, new_n10197,
    new_n10198, new_n10199, new_n10200, new_n10201, new_n10202, new_n10203,
    new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209,
    new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215,
    new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236, new_n10237, new_n10238, new_n10239,
    new_n10240, new_n10241, new_n10242, new_n10243, new_n10244, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250, new_n10251,
    new_n10252, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10263,
    new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269,
    new_n10270, new_n10271, new_n10272, new_n10273, new_n10274, new_n10275,
    new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283, new_n10284, new_n10285, new_n10286, new_n10287,
    new_n10288, new_n10289, new_n10290, new_n10291, new_n10292, new_n10293,
    new_n10294, new_n10295, new_n10296, new_n10297, new_n10298, new_n10299,
    new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305,
    new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311,
    new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317,
    new_n10318, new_n10319, new_n10320, new_n10321, new_n10322, new_n10323,
    new_n10324, new_n10325, new_n10326, new_n10327, new_n10328, new_n10329,
    new_n10330, new_n10331, new_n10332, new_n10333, new_n10334, new_n10335,
    new_n10336, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377,
    new_n10378, new_n10379, new_n10380, new_n10381, new_n10382, new_n10383,
    new_n10384, new_n10385, new_n10386, new_n10387, new_n10388, new_n10389,
    new_n10390, new_n10391, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439, new_n10440, new_n10441, new_n10442, new_n10443,
    new_n10444, new_n10445, new_n10446, new_n10447, new_n10448, new_n10449,
    new_n10450, new_n10451, new_n10452, new_n10453, new_n10454, new_n10455,
    new_n10456, new_n10457, new_n10458, new_n10459, new_n10460, new_n10461,
    new_n10462, new_n10463, new_n10464, new_n10465, new_n10466, new_n10467,
    new_n10468, new_n10469, new_n10470, new_n10471, new_n10472, new_n10473,
    new_n10474, new_n10475, new_n10476, new_n10477, new_n10478, new_n10479,
    new_n10480, new_n10481, new_n10482, new_n10483, new_n10484, new_n10485,
    new_n10486, new_n10487, new_n10488, new_n10489, new_n10490, new_n10491,
    new_n10492, new_n10493, new_n10494, new_n10495, new_n10496, new_n10497,
    new_n10498, new_n10499, new_n10500, new_n10501, new_n10502, new_n10503,
    new_n10504, new_n10505, new_n10506, new_n10507, new_n10508, new_n10509,
    new_n10510, new_n10511, new_n10512, new_n10513, new_n10514, new_n10515,
    new_n10516, new_n10517, new_n10518, new_n10519, new_n10520, new_n10521,
    new_n10522, new_n10523, new_n10524, new_n10525, new_n10526, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545, new_n10546, new_n10547,
    new_n10548, new_n10549, new_n10550, new_n10551, new_n10552, new_n10553,
    new_n10554, new_n10555, new_n10556, new_n10557, new_n10558, new_n10559,
    new_n10560, new_n10561, new_n10562, new_n10563, new_n10564, new_n10565,
    new_n10566, new_n10567, new_n10568, new_n10569, new_n10570, new_n10571,
    new_n10572, new_n10573, new_n10574, new_n10575, new_n10576, new_n10577,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588, new_n10589,
    new_n10590, new_n10591, new_n10592, new_n10593, new_n10594, new_n10595,
    new_n10596, new_n10597, new_n10598, new_n10599, new_n10600, new_n10601,
    new_n10602, new_n10603, new_n10604, new_n10605, new_n10606, new_n10607,
    new_n10608, new_n10609, new_n10610, new_n10611, new_n10612, new_n10613,
    new_n10614, new_n10615, new_n10616, new_n10617, new_n10618, new_n10619,
    new_n10620, new_n10621, new_n10622, new_n10623, new_n10624, new_n10625,
    new_n10626, new_n10627, new_n10628, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647, new_n10648, new_n10649,
    new_n10650, new_n10651, new_n10652, new_n10653, new_n10654, new_n10655,
    new_n10656, new_n10657, new_n10658, new_n10659, new_n10660, new_n10661,
    new_n10662, new_n10663, new_n10664, new_n10665, new_n10666, new_n10667,
    new_n10668, new_n10669, new_n10670, new_n10671, new_n10672, new_n10673,
    new_n10674, new_n10675, new_n10676, new_n10677, new_n10678, new_n10679,
    new_n10680, new_n10681, new_n10682, new_n10683, new_n10684, new_n10685,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695, new_n10696, new_n10697,
    new_n10698, new_n10699, new_n10700, new_n10701, new_n10702, new_n10703,
    new_n10704, new_n10705, new_n10706, new_n10707, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923, new_n10924,
    new_n10925, new_n10926, new_n10927, new_n10928, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954,
    new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961, new_n10962, new_n10963, new_n10964, new_n10965, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990,
    new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996,
    new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002,
    new_n11003, new_n11004, new_n11005, new_n11006, new_n11007, new_n11008,
    new_n11009, new_n11010, new_n11011, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023, new_n11024, new_n11025, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054, new_n11055, new_n11056,
    new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062,
    new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068,
    new_n11069, new_n11070, new_n11071, new_n11072, new_n11073, new_n11074,
    new_n11075, new_n11076, new_n11077, new_n11078, new_n11079, new_n11080,
    new_n11081, new_n11082, new_n11083;
  nand     g00000 ( new_n377 , pi119 , pi131 );
  nand     g00001 ( new_n378 , pi147 , pi168 );
  nand     g00002 ( new_n379 , pi164 , pi213 );
  nand     g00003 ( new_n380 , pi027 , pi236 );
  nand g00004 ( new_n381 , new_n380 , new_n380 );
  xor      g00005 ( new_n382 , new_n379 , new_n381 );
  xor      g00006 ( new_n383 , new_n378 , new_n382 );
  nand g00007 ( new_n384 , new_n383 , new_n383 );
  xor      g00008 ( po000 , new_n377 , new_n384 );
  nand     g00009 ( new_n386 , pi072 , pi103 );
  nand     g00010 ( new_n387 , pi016 , pi119 );
  nand     g00011 ( new_n388 , pi045 , pi117 );
  nand     g00012 ( new_n389 , pi103 , pi250 );
  xor      g00013 ( new_n390 , new_n388 , new_n389 );
  xor      g00014 ( new_n391 , new_n387 , new_n390 );
  nand g00015 ( new_n392 , new_n391 , new_n391 );
  nand     g00016 ( new_n393 , pi103 , pi119 );
  nor      g00017 ( new_n394 , new_n388 , new_n393 );
  nand     g00018 ( new_n395 , new_n392 , new_n394 );
  nand     g00019 ( new_n396 , pi117 , pi250 );
  nand     g00020 ( new_n397 , pi016 , pi045 );
  nand     g00021 ( new_n398 , pi080 , pi119 );
  xor      g00022 ( new_n399 , new_n397 , new_n398 );
  xor      g00023 ( new_n400 , new_n396 , new_n399 );
  nand     g00024 ( new_n401 , pi044 , pi103 );
  nand     g00025 ( new_n402 , new_n388 , new_n389 );
  nand     g00026 ( new_n403 , new_n387 , new_n390 );
  nand     g00027 ( new_n404 , new_n402 , new_n403 );
  xor      g00028 ( new_n405 , new_n401 , new_n404 );
  xor      g00029 ( new_n406 , new_n400 , new_n405 );
  nor      g00030 ( new_n407 , new_n395 , new_n406 );
  nand g00031 ( new_n408 , new_n407 , new_n407 );
  nand     g00032 ( new_n409 , pi054 , pi103 );
  nand     g00033 ( new_n410 , pi016 , pi250 );
  nand     g00034 ( new_n411 , pi119 , pi247 );
  nand     g00035 ( new_n412 , pi045 , pi080 );
  xor      g00036 ( new_n413 , new_n411 , new_n412 );
  xor      g00037 ( new_n414 , new_n410 , new_n413 );
  nand     g00038 ( new_n415 , pi044 , pi117 );
  nand     g00039 ( new_n416 , new_n397 , new_n398 );
  nand     g00040 ( new_n417 , new_n396 , new_n399 );
  nand     g00041 ( new_n418 , new_n416 , new_n417 );
  xor      g00042 ( new_n419 , new_n415 , new_n418 );
  xor      g00043 ( new_n420 , new_n414 , new_n419 );
  xor      g00044 ( new_n421 , new_n409 , new_n420 );
  nor      g00045 ( new_n422 , new_n401 , new_n404 );
  nand g00046 ( new_n423 , new_n400 , new_n400 );
  nand     g00047 ( new_n424 , new_n423 , new_n405 );
  nand g00048 ( new_n425 , new_n424 , new_n424 );
  nor      g00049 ( new_n426 , new_n422 , new_n425 );
  xor      g00050 ( new_n427 , new_n421 , new_n426 );
  nor      g00051 ( new_n428 , new_n408 , new_n427 );
  nand g00052 ( new_n429 , new_n428 , new_n428 );
  nand     g00053 ( new_n430 , new_n386 , new_n429 );
  nor      g00054 ( new_n431 , new_n409 , new_n420 );
  nand g00055 ( new_n432 , new_n421 , new_n421 );
  nor      g00056 ( new_n433 , new_n432 , new_n426 );
  nor      g00057 ( new_n434 , new_n431 , new_n433 );
  nand     g00058 ( new_n435 , pi054 , pi117 );
  nand     g00059 ( new_n436 , pi016 , pi044 );
  and      g00060 ( new_n437 , new_n435 , new_n436 );
  nand     g00061 ( new_n438 , pi016 , pi054 );
  nor      g00062 ( new_n439 , new_n415 , new_n438 );
  or       g00063 ( new_n440 , new_n437 , new_n439 );
  nand     g00064 ( new_n441 , pi045 , pi247 );
  nand     g00065 ( new_n442 , pi119 , pi234 );
  nand     g00066 ( new_n443 , new_n441 , new_n442 );
  nand     g00067 ( new_n444 , pi045 , pi234 );
  nor      g00068 ( new_n445 , new_n411 , new_n444 );
  nand g00069 ( new_n446 , new_n445 , new_n445 );
  nand     g00070 ( new_n447 , new_n443 , new_n446 );
  nand     g00071 ( new_n448 , pi080 , pi250 );
  nand     g00072 ( new_n449 , new_n411 , new_n412 );
  nand     g00073 ( new_n450 , new_n410 , new_n413 );
  nand     g00074 ( new_n451 , new_n449 , new_n450 );
  xor      g00075 ( new_n452 , new_n448 , new_n451 );
  xor      g00076 ( new_n453 , new_n447 , new_n452 );
  xor      g00077 ( new_n454 , new_n440 , new_n453 );
  nand     g00078 ( new_n455 , new_n415 , new_n418 );
  nand     g00079 ( new_n456 , new_n414 , new_n419 );
  nand     g00080 ( new_n457 , new_n455 , new_n456 );
  xor      g00081 ( new_n458 , new_n454 , new_n457 );
  xor      g00082 ( new_n459 , new_n434 , new_n458 );
  xor      g00083 ( new_n460 , new_n386 , new_n428 );
  or       g00084 ( new_n461 , new_n459 , new_n460 );
  nand     g00085 ( new_n462 , new_n430 , new_n461 );
  or       g00086 ( new_n463 , new_n434 , new_n458 );
  nand g00087 ( new_n464 , new_n454 , new_n454 );
  nor      g00088 ( new_n465 , new_n464 , new_n457 );
  nand g00089 ( new_n466 , new_n465 , new_n465 );
  nor      g00090 ( new_n467 , new_n440 , new_n453 );
  nor      g00091 ( new_n468 , new_n439 , new_n467 );
  nand     g00092 ( new_n469 , new_n466 , new_n468 );
  nand     g00093 ( new_n470 , new_n439 , new_n465 );
  nand     g00094 ( new_n471 , new_n469 , new_n470 );
  nand     g00095 ( new_n472 , pi247 , pi250 );
  nand     g00096 ( new_n473 , pi119 , pi214 );
  xor      g00097 ( new_n474 , new_n472 , new_n473 );
  xor      g00098 ( new_n475 , new_n444 , new_n474 );
  nand     g00099 ( new_n476 , pi044 , pi080 );
  xor      g00100 ( new_n477 , new_n445 , new_n476 );
  xor      g00101 ( new_n478 , new_n475 , new_n477 );
  nand     g00102 ( new_n479 , new_n448 , new_n451 );
  nand     g00103 ( new_n480 , new_n447 , new_n452 );
  nand     g00104 ( new_n481 , new_n479 , new_n480 );
  nand     g00105 ( new_n482 , pi103 , pi248 );
  nand     g00106 ( new_n483 , pi072 , pi117 );
  xor      g00107 ( new_n484 , new_n438 , new_n483 );
  xor      g00108 ( new_n485 , new_n482 , new_n484 );
  xnor     g00109 ( new_n486 , new_n481 , new_n485 );
  xor      g00110 ( new_n487 , new_n478 , new_n486 );
  nand g00111 ( new_n488 , new_n487 , new_n487 );
  xor      g00112 ( new_n489 , new_n471 , new_n488 );
  xnor     g00113 ( new_n490 , new_n463 , new_n489 );
  xor      g00114 ( new_n491 , new_n462 , new_n490 );
  nand     g00115 ( new_n492 , pi164 , pi228 );
  nand     g00116 ( new_n493 , pi148 , pi206 );
  nand     g00117 ( new_n494 , pi032 , pi163 );
  xor      g00118 ( new_n495 , new_n493 , new_n494 );
  xnor     g00119 ( new_n496 , new_n492 , new_n495 );
  nand     g00120 ( new_n497 , pi163 , pi164 );
  or       g00121 ( new_n498 , new_n493 , new_n497 );
  nand g00122 ( new_n499 , new_n498 , new_n498 );
  nand     g00123 ( new_n500 , new_n496 , new_n499 );
  nand     g00124 ( new_n501 , pi145 , pi163 );
  nand     g00125 ( new_n502 , new_n493 , new_n494 );
  nand     g00126 ( new_n503 , new_n492 , new_n495 );
  nand     g00127 ( new_n504 , new_n502 , new_n503 );
  xor      g00128 ( new_n505 , new_n501 , new_n504 );
  nand     g00129 ( new_n506 , pi206 , pi228 );
  nand     g00130 ( new_n507 , pi032 , pi148 );
  nand     g00131 ( new_n508 , pi039 , pi164 );
  xor      g00132 ( new_n509 , new_n507 , new_n508 );
  xor      g00133 ( new_n510 , new_n506 , new_n509 );
  xor      g00134 ( new_n511 , new_n505 , new_n510 );
  nor      g00135 ( new_n512 , new_n500 , new_n511 );
  nand     g00136 ( new_n513 , pi163 , pi246 );
  nand     g00137 ( new_n514 , new_n501 , new_n504 );
  nand     g00138 ( new_n515 , new_n505 , new_n510 );
  nand     g00139 ( new_n516 , new_n514 , new_n515 );
  xor      g00140 ( new_n517 , new_n513 , new_n516 );
  nand     g00141 ( new_n518 , new_n507 , new_n508 );
  nand     g00142 ( new_n519 , new_n506 , new_n509 );
  nand     g00143 ( new_n520 , new_n518 , new_n519 );
  nand     g00144 ( new_n521 , pi145 , pi148 );
  xor      g00145 ( new_n522 , new_n520 , new_n521 );
  nand     g00146 ( new_n523 , pi116 , pi164 );
  nand     g00147 ( new_n524 , pi032 , pi228 );
  nand     g00148 ( new_n525 , pi039 , pi206 );
  xor      g00149 ( new_n526 , new_n524 , new_n525 );
  xor      g00150 ( new_n527 , new_n523 , new_n526 );
  xnor     g00151 ( new_n528 , new_n522 , new_n527 );
  xor      g00152 ( new_n529 , new_n517 , new_n528 );
  nand     g00153 ( new_n530 , new_n512 , new_n529 );
  nand     g00154 ( new_n531 , pi114 , pi163 );
  xor      g00155 ( new_n532 , new_n530 , new_n531 );
  nor      g00156 ( new_n533 , new_n513 , new_n516 );
  and      g00157 ( new_n534 , new_n517 , new_n528 );
  nor      g00158 ( new_n535 , new_n533 , new_n534 );
  nand     g00159 ( new_n536 , pi032 , pi039 );
  nand     g00160 ( new_n537 , pi116 , pi206 );
  nand     g00161 ( new_n538 , pi070 , pi164 );
  nand     g00162 ( new_n539 , new_n537 , new_n538 );
  nand     g00163 ( new_n540 , pi070 , pi206 );
  or       g00164 ( new_n541 , new_n523 , new_n540 );
  nand     g00165 ( new_n542 , new_n539 , new_n541 );
  xor      g00166 ( new_n543 , new_n536 , new_n542 );
  nand     g00167 ( new_n544 , new_n524 , new_n525 );
  nand     g00168 ( new_n545 , new_n523 , new_n526 );
  nand     g00169 ( new_n546 , new_n544 , new_n545 );
  xor      g00170 ( new_n547 , new_n543 , new_n546 );
  nand     g00171 ( new_n548 , pi145 , pi228 );
  nand     g00172 ( new_n549 , pi148 , pi246 );
  and      g00173 ( new_n550 , new_n548 , new_n549 );
  nand     g00174 ( new_n551 , pi228 , pi246 );
  nor      g00175 ( new_n552 , new_n521 , new_n551 );
  or       g00176 ( new_n553 , new_n550 , new_n552 );
  xnor     g00177 ( new_n554 , new_n547 , new_n553 );
  nand     g00178 ( new_n555 , new_n520 , new_n521 );
  nand     g00179 ( new_n556 , new_n522 , new_n527 );
  nand     g00180 ( new_n557 , new_n555 , new_n556 );
  xnor     g00181 ( new_n558 , new_n554 , new_n557 );
  xnor     g00182 ( new_n559 , new_n535 , new_n558 );
  xor      g00183 ( new_n560 , new_n532 , new_n559 );
  nand     g00184 ( new_n561 , pi026 , pi171 );
  nand     g00185 ( new_n562 , pi027 , pi049 );
  nand     g00186 ( new_n563 , pi008 , pi107 );
  nor      g00187 ( new_n564 , new_n562 , new_n563 );
  nand g00188 ( new_n565 , new_n561 , new_n561 );
  nand     g00189 ( new_n566 , pi027 , pi107 );
  and      g00190 ( new_n567 , new_n565 , new_n566 );
  and      g00191 ( new_n568 , new_n562 , new_n563 );
  nand g00192 ( new_n569 , new_n568 , new_n568 );
  nor      g00193 ( new_n570 , new_n567 , new_n569 );
  nor      g00194 ( new_n571 , new_n564 , new_n570 );
  nor      g00195 ( new_n572 , new_n561 , new_n571 );
  nand g00196 ( new_n573 , new_n572 , new_n572 );
  nand     g00197 ( new_n574 , pi027 , pi245 );
  nand     g00198 ( new_n575 , pi026 , pi049 );
  nand     g00199 ( new_n576 , pi008 , pi171 );
  xor      g00200 ( new_n577 , new_n575 , new_n576 );
  xor      g00201 ( new_n578 , new_n574 , new_n577 );
  nor      g00202 ( new_n579 , new_n565 , new_n564 );
  or       g00203 ( new_n580 , new_n568 , new_n579 );
  nand     g00204 ( new_n581 , pi056 , pi107 );
  xnor     g00205 ( new_n582 , new_n580 , new_n581 );
  xnor     g00206 ( new_n583 , new_n578 , new_n582 );
  or       g00207 ( new_n584 , new_n573 , new_n583 );
  nand     g00208 ( new_n585 , pi107 , pi136 );
  nor      g00209 ( new_n586 , new_n580 , new_n581 );
  nor      g00210 ( new_n587 , new_n578 , new_n582 );
  nor      g00211 ( new_n588 , new_n586 , new_n587 );
  xnor     g00212 ( new_n589 , new_n585 , new_n588 );
  nand     g00213 ( new_n590 , pi027 , pi201 );
  nand     g00214 ( new_n591 , pi008 , pi049 );
  nand     g00215 ( new_n592 , pi026 , pi245 );
  xor      g00216 ( new_n593 , new_n591 , new_n592 );
  xor      g00217 ( new_n594 , new_n590 , new_n593 );
  nand     g00218 ( new_n595 , new_n575 , new_n576 );
  nand     g00219 ( new_n596 , new_n574 , new_n577 );
  nand     g00220 ( new_n597 , new_n595 , new_n596 );
  nand     g00221 ( new_n598 , pi056 , pi171 );
  xor      g00222 ( new_n599 , new_n597 , new_n598 );
  xor      g00223 ( new_n600 , new_n594 , new_n599 );
  xnor     g00224 ( new_n601 , new_n589 , new_n600 );
  or       g00225 ( new_n602 , new_n584 , new_n601 );
  nand     g00226 ( new_n603 , pi096 , pi107 );
  xor      g00227 ( new_n604 , new_n602 , new_n603 );
  nor      g00228 ( new_n605 , new_n585 , new_n588 );
  nor      g00229 ( new_n606 , new_n589 , new_n600 );
  or       g00230 ( new_n607 , new_n605 , new_n606 );
  nand     g00231 ( new_n608 , new_n591 , new_n592 );
  nand     g00232 ( new_n609 , new_n590 , new_n593 );
  nand     g00233 ( new_n610 , new_n608 , new_n609 );
  nand     g00234 ( new_n611 , pi008 , pi245 );
  nand     g00235 ( new_n612 , pi027 , pi156 );
  nand     g00236 ( new_n613 , pi026 , pi201 );
  nand     g00237 ( new_n614 , new_n612 , new_n613 );
  nand     g00238 ( new_n615 , pi026 , pi156 );
  nor      g00239 ( new_n616 , new_n590 , new_n615 );
  nand g00240 ( new_n617 , new_n616 , new_n616 );
  nand     g00241 ( new_n618 , new_n614 , new_n617 );
  xor      g00242 ( new_n619 , new_n611 , new_n618 );
  xor      g00243 ( new_n620 , new_n610 , new_n619 );
  nand     g00244 ( new_n621 , new_n597 , new_n598 );
  nand     g00245 ( new_n622 , new_n594 , new_n599 );
  nand     g00246 ( new_n623 , new_n621 , new_n622 );
  nand     g00247 ( new_n624 , pi049 , pi056 );
  nand     g00248 ( new_n625 , pi136 , pi171 );
  nand     g00249 ( new_n626 , new_n624 , new_n625 );
  nand     g00250 ( new_n627 , pi049 , pi136 );
  nor      g00251 ( new_n628 , new_n598 , new_n627 );
  nand g00252 ( new_n629 , new_n628 , new_n628 );
  nand     g00253 ( new_n630 , new_n626 , new_n629 );
  xor      g00254 ( new_n631 , new_n623 , new_n630 );
  xnor     g00255 ( new_n632 , new_n620 , new_n631 );
  xnor     g00256 ( new_n633 , new_n607 , new_n632 );
  xnor     g00257 ( new_n634 , new_n604 , new_n633 );
  xor      g00258 ( new_n635 , new_n560 , new_n634 );
  xor      g00259 ( new_n636 , new_n572 , new_n583 );
  nand     g00260 ( new_n637 , pi026 , pi107 );
  nand     g00261 ( new_n638 , pi027 , pi171 );
  xnor     g00262 ( new_n639 , new_n637 , new_n638 );
  nand     g00263 ( new_n640 , pi163 , pi206 );
  nand     g00264 ( new_n641 , pi148 , pi164 );
  nand     g00265 ( new_n642 , new_n640 , new_n641 );
  nand     g00266 ( new_n643 , new_n498 , new_n642 );
  nand     g00267 ( new_n644 , new_n639 , new_n643 );
  or       g00268 ( new_n645 , new_n497 , new_n566 );
  xor      g00269 ( new_n646 , new_n639 , new_n643 );
  nand     g00270 ( new_n647 , new_n645 , new_n646 );
  nand     g00271 ( new_n648 , new_n644 , new_n647 );
  nand     g00272 ( new_n649 , new_n567 , new_n569 );
  nand     g00273 ( new_n650 , new_n571 , new_n649 );
  nand     g00274 ( new_n651 , new_n648 , new_n650 );
  xor      g00275 ( new_n652 , new_n496 , new_n498 );
  xor      g00276 ( new_n653 , new_n648 , new_n650 );
  nand     g00277 ( new_n654 , new_n652 , new_n653 );
  nand     g00278 ( new_n655 , new_n651 , new_n654 );
  and      g00279 ( new_n656 , new_n636 , new_n655 );
  and      g00280 ( new_n657 , new_n648 , new_n650 );
  and      g00281 ( new_n658 , new_n652 , new_n653 );
  nor      g00282 ( new_n659 , new_n657 , new_n658 );
  xor      g00283 ( new_n660 , new_n636 , new_n659 );
  xor      g00284 ( new_n661 , new_n500 , new_n511 );
  nor      g00285 ( new_n662 , new_n660 , new_n661 );
  nor      g00286 ( new_n663 , new_n656 , new_n662 );
  xor      g00287 ( new_n664 , new_n584 , new_n601 );
  nor      g00288 ( new_n665 , new_n663 , new_n664 );
  nand     g00289 ( new_n666 , new_n636 , new_n655 );
  xor      g00290 ( new_n667 , new_n636 , new_n655 );
  nand g00291 ( new_n668 , new_n661 , new_n661 );
  nand     g00292 ( new_n669 , new_n667 , new_n668 );
  nand     g00293 ( new_n670 , new_n666 , new_n669 );
  xor      g00294 ( new_n671 , new_n670 , new_n664 );
  xor      g00295 ( new_n672 , new_n512 , new_n529 );
  nor      g00296 ( new_n673 , new_n671 , new_n672 );
  nor      g00297 ( new_n674 , new_n665 , new_n673 );
  xor      g00298 ( new_n675 , new_n635 , new_n674 );
  nand     g00299 ( new_n676 , pi075 , pi175 );
  nand     g00300 ( new_n677 , pi134 , pi151 );
  nand     g00301 ( new_n678 , pi147 , pi240 );
  nand     g00302 ( new_n679 , pi019 , pi175 );
  or       g00303 ( new_n680 , new_n678 , new_n679 );
  nand     g00304 ( new_n681 , new_n677 , new_n680 );
  nand     g00305 ( new_n682 , new_n678 , new_n679 );
  nand     g00306 ( new_n683 , new_n681 , new_n682 );
  nand     g00307 ( new_n684 , pi097 , pi175 );
  nor      g00308 ( new_n685 , new_n683 , new_n684 );
  xnor     g00309 ( new_n686 , new_n683 , new_n684 );
  nand     g00310 ( new_n687 , pi147 , pi149 );
  nand     g00311 ( new_n688 , pi019 , pi134 );
  nand     g00312 ( new_n689 , pi151 , pi240 );
  xor      g00313 ( new_n690 , new_n688 , new_n689 );
  xor      g00314 ( new_n691 , new_n687 , new_n690 );
  nor      g00315 ( new_n692 , new_n686 , new_n691 );
  nor      g00316 ( new_n693 , new_n685 , new_n692 );
  xor      g00317 ( new_n694 , new_n676 , new_n693 );
  nand     g00318 ( new_n695 , pi019 , pi240 );
  nand     g00319 ( new_n696 , pi147 , pi167 );
  nand     g00320 ( new_n697 , pi149 , pi151 );
  xor      g00321 ( new_n698 , new_n696 , new_n697 );
  xor      g00322 ( new_n699 , new_n695 , new_n698 );
  nand     g00323 ( new_n700 , pi097 , pi134 );
  nand     g00324 ( new_n701 , new_n688 , new_n689 );
  nand     g00325 ( new_n702 , new_n687 , new_n690 );
  nand     g00326 ( new_n703 , new_n701 , new_n702 );
  xor      g00327 ( new_n704 , new_n700 , new_n703 );
  xnor     g00328 ( new_n705 , new_n699 , new_n704 );
  xor      g00329 ( new_n706 , new_n694 , new_n705 );
  nand g00330 ( new_n707 , pi147 , pi147 );
  nand g00331 ( new_n708 , pi175 , pi175 );
  nor      g00332 ( new_n709 , new_n707 , new_n708 );
  nor      g00333 ( new_n710 , new_n677 , new_n709 );
  and      g00334 ( new_n711 , new_n680 , new_n682 );
  or       g00335 ( new_n712 , new_n710 , new_n711 );
  nor      g00336 ( new_n713 , new_n677 , new_n712 );
  nand g00337 ( new_n714 , new_n713 , new_n713 );
  xnor     g00338 ( new_n715 , new_n686 , new_n691 );
  nor      g00339 ( new_n716 , new_n714 , new_n715 );
  nand     g00340 ( new_n717 , new_n706 , new_n716 );
  nand     g00341 ( new_n718 , pi093 , pi175 );
  nand     g00342 ( new_n719 , new_n700 , new_n703 );
  nand     g00343 ( new_n720 , new_n699 , new_n704 );
  nand     g00344 ( new_n721 , new_n719 , new_n720 );
  nand     g00345 ( new_n722 , pi097 , pi240 );
  nand     g00346 ( new_n723 , pi075 , pi134 );
  and      g00347 ( new_n724 , new_n722 , new_n723 );
  nand     g00348 ( new_n725 , pi075 , pi240 );
  nor      g00349 ( new_n726 , new_n700 , new_n725 );
  or       g00350 ( new_n727 , new_n724 , new_n726 );
  nand     g00351 ( new_n728 , new_n696 , new_n697 );
  nand     g00352 ( new_n729 , new_n695 , new_n698 );
  nand     g00353 ( new_n730 , new_n728 , new_n729 );
  nand     g00354 ( new_n731 , pi019 , pi149 );
  nand     g00355 ( new_n732 , pi151 , pi167 );
  nand     g00356 ( new_n733 , pi147 , pi181 );
  nand     g00357 ( new_n734 , new_n732 , new_n733 );
  nand     g00358 ( new_n735 , pi151 , pi181 );
  or       g00359 ( new_n736 , new_n696 , new_n735 );
  nand     g00360 ( new_n737 , new_n734 , new_n736 );
  xor      g00361 ( new_n738 , new_n731 , new_n737 );
  xor      g00362 ( new_n739 , new_n730 , new_n738 );
  xor      g00363 ( new_n740 , new_n727 , new_n739 );
  nand g00364 ( new_n741 , new_n740 , new_n740 );
  xor      g00365 ( new_n742 , new_n721 , new_n741 );
  nor      g00366 ( new_n743 , new_n676 , new_n693 );
  and      g00367 ( new_n744 , new_n694 , new_n705 );
  nor      g00368 ( new_n745 , new_n743 , new_n744 );
  xor      g00369 ( new_n746 , new_n742 , new_n745 );
  xnor     g00370 ( new_n747 , new_n718 , new_n746 );
  xnor     g00371 ( new_n748 , new_n717 , new_n747 );
  nor      g00372 ( new_n749 , new_n675 , new_n748 );
  xor      g00373 ( new_n750 , new_n706 , new_n716 );
  nand g00374 ( new_n751 , new_n750 , new_n750 );
  nand     g00375 ( new_n752 , new_n682 , new_n710 );
  nand     g00376 ( new_n753 , new_n712 , new_n752 );
  xor      g00377 ( new_n754 , new_n652 , new_n653 );
  or       g00378 ( new_n755 , new_n753 , new_n754 );
  nand     g00379 ( new_n756 , pi147 , pi175 );
  xnor     g00380 ( new_n757 , new_n497 , new_n566 );
  nor      g00381 ( new_n758 , new_n756 , new_n757 );
  nand     g00382 ( new_n759 , pi151 , pi175 );
  nand     g00383 ( new_n760 , pi134 , pi147 );
  xor      g00384 ( new_n761 , new_n759 , new_n760 );
  nand     g00385 ( new_n762 , new_n758 , new_n761 );
  xor      g00386 ( new_n763 , new_n645 , new_n646 );
  xnor     g00387 ( new_n764 , new_n758 , new_n761 );
  or       g00388 ( new_n765 , new_n763 , new_n764 );
  nand     g00389 ( new_n766 , new_n762 , new_n765 );
  xor      g00390 ( new_n767 , new_n753 , new_n754 );
  nand     g00391 ( new_n768 , new_n766 , new_n767 );
  and      g00392 ( new_n769 , new_n755 , new_n768 );
  xor      g00393 ( new_n770 , new_n713 , new_n715 );
  nor      g00394 ( new_n771 , new_n769 , new_n770 );
  nand     g00395 ( new_n772 , new_n755 , new_n768 );
  xor      g00396 ( new_n773 , new_n772 , new_n770 );
  xor      g00397 ( new_n774 , new_n667 , new_n668 );
  nor      g00398 ( new_n775 , new_n773 , new_n774 );
  nor      g00399 ( new_n776 , new_n771 , new_n775 );
  nor      g00400 ( new_n777 , new_n751 , new_n776 );
  xor      g00401 ( new_n778 , new_n663 , new_n664 );
  nand g00402 ( new_n779 , new_n672 , new_n672 );
  xor      g00403 ( new_n780 , new_n778 , new_n779 );
  xor      g00404 ( new_n781 , new_n750 , new_n776 );
  nor      g00405 ( new_n782 , new_n780 , new_n781 );
  nor      g00406 ( new_n783 , new_n777 , new_n782 );
  xor      g00407 ( new_n784 , new_n717 , new_n747 );
  xor      g00408 ( new_n785 , new_n675 , new_n784 );
  nor      g00409 ( new_n786 , new_n783 , new_n785 );
  or       g00410 ( new_n787 , new_n749 , new_n786 );
  nand g00411 ( new_n788 , new_n742 , new_n742 );
  nor      g00412 ( new_n789 , new_n788 , new_n745 );
  nor      g00413 ( new_n790 , new_n727 , new_n739 );
  nor      g00414 ( new_n791 , new_n721 , new_n741 );
  xor      g00415 ( new_n792 , new_n726 , new_n791 );
  nor      g00416 ( new_n793 , new_n790 , new_n792 );
  nand g00417 ( new_n794 , new_n725 , new_n725 );
  nand     g00418 ( new_n795 , pi093 , pi134 );
  and      g00419 ( new_n796 , pi166 , pi175 );
  xor      g00420 ( new_n797 , new_n795 , new_n796 );
  xor      g00421 ( new_n798 , new_n794 , new_n797 );
  nand     g00422 ( new_n799 , new_n731 , new_n737 );
  nand     g00423 ( new_n800 , new_n730 , new_n738 );
  nand     g00424 ( new_n801 , new_n799 , new_n800 );
  xor      g00425 ( new_n802 , new_n798 , new_n801 );
  nand     g00426 ( new_n803 , pi097 , pi149 );
  xor      g00427 ( new_n804 , new_n736 , new_n803 );
  nand     g00428 ( new_n805 , pi019 , pi167 );
  nand     g00429 ( new_n806 , pi147 , pi200 );
  xor      g00430 ( new_n807 , new_n805 , new_n806 );
  xor      g00431 ( new_n808 , new_n735 , new_n807 );
  xor      g00432 ( new_n809 , new_n804 , new_n808 );
  xor      g00433 ( new_n810 , new_n802 , new_n809 );
  xor      g00434 ( new_n811 , new_n793 , new_n810 );
  xor      g00435 ( new_n812 , new_n789 , new_n811 );
  nor      g00436 ( new_n813 , new_n718 , new_n746 );
  nor      g00437 ( new_n814 , new_n717 , new_n747 );
  nor      g00438 ( new_n815 , new_n813 , new_n814 );
  xor      g00439 ( new_n816 , new_n812 , new_n815 );
  nand g00440 ( new_n817 , new_n560 , new_n560 );
  and      g00441 ( new_n818 , new_n817 , new_n634 );
  or       g00442 ( new_n819 , new_n663 , new_n664 );
  nand     g00443 ( new_n820 , new_n778 , new_n779 );
  nand     g00444 ( new_n821 , new_n819 , new_n820 );
  nor      g00445 ( new_n822 , new_n635 , new_n821 );
  nor      g00446 ( new_n823 , new_n818 , new_n822 );
  nand     g00447 ( new_n824 , new_n602 , new_n603 );
  nand     g00448 ( new_n825 , new_n604 , new_n633 );
  nand     g00449 ( new_n826 , new_n824 , new_n825 );
  nand     g00450 ( new_n827 , new_n607 , new_n632 );
  nand     g00451 ( new_n828 , new_n623 , new_n630 );
  nand     g00452 ( new_n829 , new_n620 , new_n631 );
  nand     g00453 ( new_n830 , new_n828 , new_n829 );
  xor      g00454 ( new_n831 , new_n628 , new_n830 );
  nand     g00455 ( new_n832 , pi096 , pi171 );
  nand     g00456 ( new_n833 , pi107 , pi235 );
  xor      g00457 ( new_n834 , new_n832 , new_n833 );
  xor      g00458 ( new_n835 , new_n627 , new_n834 );
  nand     g00459 ( new_n836 , new_n611 , new_n618 );
  nand     g00460 ( new_n837 , new_n610 , new_n619 );
  nand     g00461 ( new_n838 , new_n836 , new_n837 );
  xnor     g00462 ( new_n839 , new_n835 , new_n838 );
  nand     g00463 ( new_n840 , pi056 , pi245 );
  xor      g00464 ( new_n841 , new_n616 , new_n840 );
  nand     g00465 ( new_n842 , pi008 , pi201 );
  nand     g00466 ( new_n843 , pi027 , pi063 );
  xor      g00467 ( new_n844 , new_n842 , new_n843 );
  xor      g00468 ( new_n845 , new_n615 , new_n844 );
  xnor     g00469 ( new_n846 , new_n841 , new_n845 );
  xor      g00470 ( new_n847 , new_n839 , new_n846 );
  xor      g00471 ( new_n848 , new_n831 , new_n847 );
  xnor     g00472 ( new_n849 , new_n827 , new_n848 );
  xnor     g00473 ( new_n850 , new_n826 , new_n849 );
  nand     g00474 ( new_n851 , new_n530 , new_n531 );
  nand     g00475 ( new_n852 , new_n532 , new_n559 );
  nand     g00476 ( new_n853 , new_n851 , new_n852 );
  nand g00477 ( new_n854 , new_n853 , new_n853 );
  nor      g00478 ( new_n855 , new_n535 , new_n558 );
  nand     g00479 ( new_n856 , pi039 , pi145 );
  xnor     g00480 ( new_n857 , new_n541 , new_n856 );
  nand     g00481 ( new_n858 , pi115 , pi164 );
  nand     g00482 ( new_n859 , pi032 , pi116 );
  xor      g00483 ( new_n860 , new_n858 , new_n859 );
  xor      g00484 ( new_n861 , new_n540 , new_n860 );
  xnor     g00485 ( new_n862 , new_n857 , new_n861 );
  nand     g00486 ( new_n863 , new_n536 , new_n542 );
  nand     g00487 ( new_n864 , new_n543 , new_n546 );
  nand     g00488 ( new_n865 , new_n863 , new_n864 );
  nand     g00489 ( new_n866 , pi114 , pi148 );
  nand     g00490 ( new_n867 , pi091 , pi163 );
  xor      g00491 ( new_n868 , new_n866 , new_n867 );
  xor      g00492 ( new_n869 , new_n551 , new_n868 );
  xor      g00493 ( new_n870 , new_n865 , new_n869 );
  xor      g00494 ( new_n871 , new_n862 , new_n870 );
  nor      g00495 ( new_n872 , new_n547 , new_n553 );
  nor      g00496 ( new_n873 , new_n554 , new_n557 );
  xor      g00497 ( new_n874 , new_n552 , new_n873 );
  nor      g00498 ( new_n875 , new_n872 , new_n874 );
  xor      g00499 ( new_n876 , new_n871 , new_n875 );
  xor      g00500 ( new_n877 , new_n855 , new_n876 );
  xor      g00501 ( new_n878 , new_n854 , new_n877 );
  xnor     g00502 ( new_n879 , new_n850 , new_n878 );
  xor      g00503 ( new_n880 , new_n823 , new_n879 );
  xnor     g00504 ( new_n881 , new_n816 , new_n880 );
  xor      g00505 ( new_n882 , new_n787 , new_n881 );
  xor      g00506 ( new_n883 , new_n491 , new_n882 );
  xor      g00507 ( new_n884 , new_n408 , new_n427 );
  xor      g00508 ( new_n885 , new_n773 , new_n774 );
  xor      g00509 ( new_n886 , new_n395 , new_n406 );
  nor      g00510 ( new_n887 , new_n885 , new_n886 );
  xor      g00511 ( new_n888 , new_n392 , new_n394 );
  xor      g00512 ( new_n889 , new_n756 , new_n757 );
  nand g00513 ( new_n890 , new_n889 , new_n889 );
  nor      g00514 ( new_n891 , new_n393 , new_n890 );
  nand g00515 ( new_n892 , new_n891 , new_n891 );
  nand     g00516 ( new_n893 , pi045 , pi103 );
  nand     g00517 ( new_n894 , pi117 , pi119 );
  and      g00518 ( new_n895 , new_n893 , new_n894 );
  or       g00519 ( new_n896 , new_n394 , new_n895 );
  nand     g00520 ( new_n897 , new_n892 , new_n896 );
  nand g00521 ( new_n898 , new_n897 , new_n897 );
  xor      g00522 ( new_n899 , new_n891 , new_n896 );
  xor      g00523 ( new_n900 , new_n763 , new_n764 );
  nor      g00524 ( new_n901 , new_n899 , new_n900 );
  or       g00525 ( new_n902 , new_n898 , new_n901 );
  nand g00526 ( new_n903 , new_n902 , new_n902 );
  nor      g00527 ( new_n904 , new_n888 , new_n903 );
  xor      g00528 ( new_n905 , new_n888 , new_n902 );
  xor      g00529 ( new_n906 , new_n766 , new_n767 );
  nor      g00530 ( new_n907 , new_n905 , new_n906 );
  nor      g00531 ( new_n908 , new_n904 , new_n907 );
  xnor     g00532 ( new_n909 , new_n885 , new_n886 );
  nor      g00533 ( new_n910 , new_n908 , new_n909 );
  nor      g00534 ( new_n911 , new_n887 , new_n910 );
  nand     g00535 ( new_n912 , new_n884 , new_n911 );
  xor      g00536 ( new_n913 , new_n780 , new_n781 );
  xor      g00537 ( new_n914 , new_n884 , new_n911 );
  nand     g00538 ( new_n915 , new_n913 , new_n914 );
  nand     g00539 ( new_n916 , new_n912 , new_n915 );
  xor      g00540 ( new_n917 , new_n459 , new_n460 );
  nand g00541 ( new_n918 , new_n917 , new_n917 );
  nor      g00542 ( new_n919 , new_n916 , new_n918 );
  xor      g00543 ( new_n920 , new_n916 , new_n917 );
  xor      g00544 ( new_n921 , new_n783 , new_n785 );
  nor      g00545 ( new_n922 , new_n920 , new_n921 );
  nor      g00546 ( new_n923 , new_n919 , new_n922 );
  xnor     g00547 ( po001 , new_n883 , new_n923 );
  nand     g00548 ( new_n925 , pi103 , pi143 );
  nand     g00549 ( new_n926 , pi162 , pi175 );
  nand     g00550 ( new_n927 , pi051 , pi107 );
  nand     g00551 ( new_n928 , pi163 , pi188 );
  xor      g00552 ( new_n929 , new_n927 , new_n928 );
  xor      g00553 ( new_n930 , new_n926 , new_n929 );
  or       g00554 ( new_n931 , new_n925 , new_n930 );
  nand     g00555 ( new_n932 , pi057 , pi117 );
  nor      g00556 ( new_n933 , new_n925 , new_n932 );
  nand     g00557 ( new_n934 , pi117 , pi143 );
  nand     g00558 ( new_n935 , pi057 , pi103 );
  and      g00559 ( new_n936 , new_n934 , new_n935 );
  or       g00560 ( new_n937 , new_n933 , new_n936 );
  nand     g00561 ( new_n938 , new_n931 , new_n937 );
  xnor     g00562 ( new_n939 , new_n931 , new_n937 );
  nor      g00563 ( new_n940 , new_n927 , new_n928 );
  nand     g00564 ( new_n941 , pi042 , pi171 );
  or       g00565 ( new_n942 , new_n927 , new_n941 );
  nand     g00566 ( new_n943 , pi051 , pi171 );
  nand     g00567 ( new_n944 , pi042 , pi107 );
  nand     g00568 ( new_n945 , new_n943 , new_n944 );
  nand     g00569 ( new_n946 , new_n942 , new_n945 );
  nand     g00570 ( new_n947 , pi148 , pi178 );
  nor      g00571 ( new_n948 , new_n928 , new_n947 );
  nand g00572 ( new_n949 , pi148 , pi148 );
  nand g00573 ( new_n950 , pi188 , pi188 );
  nor      g00574 ( new_n951 , new_n949 , new_n950 );
  nand g00575 ( new_n952 , pi163 , pi163 );
  nand g00576 ( new_n953 , pi178 , pi178 );
  nor      g00577 ( new_n954 , new_n952 , new_n953 );
  nor      g00578 ( new_n955 , new_n951 , new_n954 );
  or       g00579 ( new_n956 , new_n948 , new_n955 );
  xnor     g00580 ( new_n957 , new_n946 , new_n956 );
  xor      g00581 ( new_n958 , new_n940 , new_n957 );
  nand g00582 ( new_n959 , new_n929 , new_n929 );
  nor      g00583 ( new_n960 , new_n926 , new_n959 );
  nand     g00584 ( new_n961 , pi134 , pi162 );
  nand     g00585 ( new_n962 , pi033 , pi175 );
  xor      g00586 ( new_n963 , new_n961 , new_n962 );
  xnor     g00587 ( new_n964 , new_n960 , new_n963 );
  xor      g00588 ( new_n965 , new_n958 , new_n964 );
  or       g00589 ( new_n966 , new_n939 , new_n965 );
  nand     g00590 ( new_n967 , new_n938 , new_n966 );
  nand     g00591 ( new_n968 , pi016 , pi143 );
  nand     g00592 ( new_n969 , pi103 , pi194 );
  xor      g00593 ( new_n970 , new_n932 , new_n969 );
  xor      g00594 ( new_n971 , new_n968 , new_n970 );
  nand g00595 ( new_n972 , new_n971 , new_n971 );
  xor      g00596 ( new_n973 , new_n933 , new_n972 );
  nand g00597 ( new_n974 , new_n973 , new_n973 );
  or       g00598 ( new_n975 , new_n967 , new_n974 );
  xor      g00599 ( new_n976 , new_n967 , new_n974 );
  nand     g00600 ( new_n977 , new_n960 , new_n963 );
  or       g00601 ( new_n978 , new_n958 , new_n964 );
  nand     g00602 ( new_n979 , new_n977 , new_n978 );
  nand     g00603 ( new_n980 , pi188 , pi228 );
  nand     g00604 ( new_n981 , pi061 , pi163 );
  xor      g00605 ( new_n982 , new_n947 , new_n981 );
  xor      g00606 ( new_n983 , new_n980 , new_n982 );
  xor      g00607 ( new_n984 , new_n948 , new_n983 );
  nand     g00608 ( new_n985 , pi049 , pi051 );
  nand     g00609 ( new_n986 , pi107 , pi108 );
  xor      g00610 ( new_n987 , new_n941 , new_n986 );
  xor      g00611 ( new_n988 , new_n985 , new_n987 );
  xnor     g00612 ( new_n989 , new_n942 , new_n988 );
  xor      g00613 ( new_n990 , new_n984 , new_n989 );
  and      g00614 ( new_n991 , new_n946 , new_n956 );
  nor      g00615 ( new_n992 , new_n940 , new_n957 );
  or       g00616 ( new_n993 , new_n991 , new_n992 );
  xor      g00617 ( new_n994 , new_n990 , new_n993 );
  nand     g00618 ( new_n995 , pi162 , pi240 );
  nand     g00619 ( new_n996 , pi175 , pi179 );
  nor      g00620 ( new_n997 , new_n995 , new_n996 );
  nand     g00621 ( new_n998 , new_n995 , new_n996 );
  nand     g00622 ( new_n999 , pi033 , pi134 );
  nand g00623 ( new_n1000 , new_n999 , new_n999 );
  and      g00624 ( new_n1001 , new_n926 , new_n1000 );
  nor      g00625 ( new_n1002 , new_n998 , new_n1001 );
  nor      g00626 ( new_n1003 , new_n997 , new_n1002 );
  nand     g00627 ( new_n1004 , new_n998 , new_n1001 );
  nand     g00628 ( new_n1005 , new_n1003 , new_n1004 );
  and      g00629 ( new_n1006 , new_n994 , new_n1005 );
  nor      g00630 ( new_n1007 , new_n994 , new_n1005 );
  nor      g00631 ( new_n1008 , new_n1006 , new_n1007 );
  xor      g00632 ( new_n1009 , new_n979 , new_n1008 );
  nand     g00633 ( new_n1010 , new_n976 , new_n1009 );
  nand     g00634 ( new_n1011 , new_n975 , new_n1010 );
  nand     g00635 ( new_n1012 , new_n933 , new_n972 );
  nand     g00636 ( new_n1013 , pi085 , pi103 );
  nand     g00637 ( new_n1014 , new_n932 , new_n969 );
  nand     g00638 ( new_n1015 , new_n968 , new_n970 );
  nand     g00639 ( new_n1016 , new_n1014 , new_n1015 );
  xor      g00640 ( new_n1017 , new_n1013 , new_n1016 );
  nand     g00641 ( new_n1018 , pi080 , pi143 );
  nand     g00642 ( new_n1019 , pi117 , pi194 );
  nand     g00643 ( new_n1020 , pi016 , pi057 );
  xor      g00644 ( new_n1021 , new_n1019 , new_n1020 );
  xor      g00645 ( new_n1022 , new_n1018 , new_n1021 );
  xor      g00646 ( new_n1023 , new_n1017 , new_n1022 );
  xnor     g00647 ( new_n1024 , new_n1012 , new_n1023 );
  xor      g00648 ( new_n1025 , new_n1011 , new_n1024 );
  nor      g00649 ( new_n1026 , new_n984 , new_n989 );
  nand g00650 ( new_n1027 , new_n990 , new_n990 );
  nor      g00651 ( new_n1028 , new_n1027 , new_n993 );
  or       g00652 ( new_n1029 , new_n1026 , new_n1028 );
  or       g00653 ( new_n1030 , new_n942 , new_n988 );
  nand     g00654 ( new_n1031 , pi108 , pi171 );
  nand     g00655 ( new_n1032 , pi051 , pi245 );
  nand     g00656 ( new_n1033 , pi042 , pi049 );
  xor      g00657 ( new_n1034 , new_n1032 , new_n1033 );
  xor      g00658 ( new_n1035 , new_n1031 , new_n1034 );
  nand     g00659 ( new_n1036 , pi007 , pi107 );
  nand     g00660 ( new_n1037 , new_n941 , new_n986 );
  nand     g00661 ( new_n1038 , new_n985 , new_n987 );
  nand     g00662 ( new_n1039 , new_n1037 , new_n1038 );
  xnor     g00663 ( new_n1040 , new_n1036 , new_n1039 );
  xnor     g00664 ( new_n1041 , new_n1035 , new_n1040 );
  xor      g00665 ( new_n1042 , new_n1030 , new_n1041 );
  nand g00666 ( new_n1043 , new_n983 , new_n983 );
  nand     g00667 ( new_n1044 , new_n948 , new_n1043 );
  nand     g00668 ( new_n1045 , pi012 , pi163 );
  nand     g00669 ( new_n1046 , new_n947 , new_n981 );
  nand     g00670 ( new_n1047 , new_n980 , new_n982 );
  nand     g00671 ( new_n1048 , new_n1046 , new_n1047 );
  xor      g00672 ( new_n1049 , new_n1045 , new_n1048 );
  nand     g00673 ( new_n1050 , pi061 , pi148 );
  nand     g00674 ( new_n1051 , pi039 , pi188 );
  nand     g00675 ( new_n1052 , pi178 , pi228 );
  xor      g00676 ( new_n1053 , new_n1051 , new_n1052 );
  xor      g00677 ( new_n1054 , new_n1050 , new_n1053 );
  xor      g00678 ( new_n1055 , new_n1049 , new_n1054 );
  xor      g00679 ( new_n1056 , new_n1044 , new_n1055 );
  xor      g00680 ( new_n1057 , new_n1042 , new_n1056 );
  xor      g00681 ( new_n1058 , new_n1029 , new_n1057 );
  nor      g00682 ( new_n1059 , new_n979 , new_n1007 );
  or       g00683 ( new_n1060 , new_n1006 , new_n1059 );
  nor      g00684 ( new_n1061 , new_n999 , new_n1003 );
  or       g00685 ( new_n1062 , new_n997 , new_n1000 );
  nand     g00686 ( new_n1063 , new_n998 , new_n1062 );
  nand     g00687 ( new_n1064 , pi048 , pi175 );
  xor      g00688 ( new_n1065 , new_n1063 , new_n1064 );
  nand     g00689 ( new_n1066 , pi134 , pi179 );
  nand     g00690 ( new_n1067 , pi149 , pi162 );
  nand     g00691 ( new_n1068 , pi033 , pi240 );
  xor      g00692 ( new_n1069 , new_n1067 , new_n1068 );
  xor      g00693 ( new_n1070 , new_n1066 , new_n1069 );
  xor      g00694 ( new_n1071 , new_n1065 , new_n1070 );
  xor      g00695 ( new_n1072 , new_n1061 , new_n1071 );
  xnor     g00696 ( new_n1073 , new_n1060 , new_n1072 );
  xor      g00697 ( new_n1074 , new_n1058 , new_n1073 );
  xor      g00698 ( po002 , new_n1025 , new_n1074 );
  nand     g00699 ( new_n1076 , pi119 , pi160 );
  nand g00700 ( new_n1077 , new_n1076 , new_n1076 );
  nand     g00701 ( new_n1078 , pi138 , pi147 );
  nand     g00702 ( new_n1079 , pi027 , pi087 );
  nand     g00703 ( new_n1080 , pi142 , pi164 );
  xnor     g00704 ( new_n1081 , new_n1079 , new_n1080 );
  xor      g00705 ( new_n1082 , new_n1078 , new_n1081 );
  xor      g00706 ( po003 , new_n1077 , new_n1082 );
  nand     g00707 ( new_n1084 , pi131 , pi217 );
  nand g00708 ( new_n1085 , new_n1084 , new_n1084 );
  nand     g00709 ( new_n1086 , pi168 , pi249 );
  nand     g00710 ( new_n1087 , pi236 , pi242 );
  nand     g00711 ( new_n1088 , pi210 , pi213 );
  nand g00712 ( new_n1089 , new_n1088 , new_n1088 );
  xor      g00713 ( new_n1090 , new_n1087 , new_n1089 );
  xor      g00714 ( new_n1091 , new_n1086 , new_n1090 );
  nand     g00715 ( new_n1092 , new_n1085 , new_n1091 );
  nand g00716 ( new_n1093 , new_n1092 , new_n1092 );
  nand     g00717 ( new_n1094 , pi100 , pi131 );
  nand     g00718 ( new_n1095 , pi052 , pi217 );
  xor      g00719 ( new_n1096 , new_n1094 , new_n1095 );
  nor      g00720 ( new_n1097 , new_n1093 , new_n1096 );
  or       g00721 ( new_n1098 , new_n1086 , new_n1090 );
  nand     g00722 ( new_n1099 , pi208 , pi222 );
  nor      g00723 ( new_n1100 , new_n1086 , new_n1099 );
  nand g00724 ( new_n1101 , new_n1100 , new_n1100 );
  nand     g00725 ( new_n1102 , pi168 , pi222 );
  nand     g00726 ( new_n1103 , pi208 , pi249 );
  nand     g00727 ( new_n1104 , new_n1102 , new_n1103 );
  nand     g00728 ( new_n1105 , new_n1101 , new_n1104 );
  xor      g00729 ( new_n1106 , new_n1098 , new_n1105 );
  nor      g00730 ( new_n1107 , new_n1087 , new_n1088 );
  nand     g00731 ( new_n1108 , pi210 , pi212 );
  nand     g00732 ( new_n1109 , pi111 , pi213 );
  xor      g00733 ( new_n1110 , new_n1108 , new_n1109 );
  nand     g00734 ( new_n1111 , pi241 , pi242 );
  nand     g00735 ( new_n1112 , pi140 , pi236 );
  xor      g00736 ( new_n1113 , new_n1111 , new_n1112 );
  xor      g00737 ( new_n1114 , new_n1110 , new_n1113 );
  xor      g00738 ( new_n1115 , new_n1107 , new_n1114 );
  xor      g00739 ( new_n1116 , new_n1106 , new_n1115 );
  xor      g00740 ( new_n1117 , new_n1092 , new_n1096 );
  nor      g00741 ( new_n1118 , new_n1116 , new_n1117 );
  nor      g00742 ( new_n1119 , new_n1097 , new_n1118 );
  nand g00743 ( new_n1120 , new_n1119 , new_n1119 );
  nand     g00744 ( new_n1121 , pi077 , pi217 );
  nand     g00745 ( new_n1122 , pi131 , pi227 );
  nor      g00746 ( new_n1123 , new_n1121 , new_n1122 );
  nand     g00747 ( new_n1124 , new_n1121 , new_n1122 );
  nand     g00748 ( new_n1125 , pi052 , pi100 );
  nor      g00749 ( new_n1126 , new_n1085 , new_n1125 );
  nor      g00750 ( new_n1127 , new_n1124 , new_n1126 );
  nor      g00751 ( new_n1128 , new_n1123 , new_n1127 );
  nand     g00752 ( new_n1129 , new_n1124 , new_n1126 );
  nand     g00753 ( new_n1130 , new_n1128 , new_n1129 );
  nand     g00754 ( new_n1131 , new_n1120 , new_n1130 );
  xor      g00755 ( new_n1132 , new_n1119 , new_n1130 );
  nor      g00756 ( new_n1133 , new_n1098 , new_n1105 );
  nand g00757 ( new_n1134 , new_n1133 , new_n1133 );
  nand     g00758 ( new_n1135 , new_n1106 , new_n1115 );
  nand     g00759 ( new_n1136 , new_n1134 , new_n1135 );
  nand     g00760 ( new_n1137 , pi139 , pi249 );
  nand     g00761 ( new_n1138 , pi125 , pi168 );
  xor      g00762 ( new_n1139 , new_n1099 , new_n1138 );
  xor      g00763 ( new_n1140 , new_n1137 , new_n1139 );
  xor      g00764 ( new_n1141 , new_n1101 , new_n1140 );
  nor      g00765 ( new_n1142 , new_n1110 , new_n1113 );
  nand g00766 ( new_n1143 , new_n1107 , new_n1107 );
  and      g00767 ( new_n1144 , new_n1143 , new_n1114 );
  nor      g00768 ( new_n1145 , new_n1142 , new_n1144 );
  nand     g00769 ( new_n1146 , pi140 , pi241 );
  nand g00770 ( new_n1147 , new_n1146 , new_n1146 );
  and      g00771 ( new_n1148 , new_n1087 , new_n1147 );
  nand     g00772 ( new_n1149 , pi161 , pi242 );
  nand     g00773 ( new_n1150 , pi236 , pi252 );
  nor      g00774 ( new_n1151 , new_n1149 , new_n1150 );
  nand     g00775 ( new_n1152 , new_n1149 , new_n1150 );
  nand g00776 ( new_n1153 , new_n1152 , new_n1152 );
  nor      g00777 ( new_n1154 , new_n1151 , new_n1153 );
  nor      g00778 ( new_n1155 , new_n1148 , new_n1154 );
  and      g00779 ( new_n1156 , new_n1152 , new_n1148 );
  nor      g00780 ( new_n1157 , new_n1155 , new_n1156 );
  nand     g00781 ( new_n1158 , pi104 , pi210 );
  nand     g00782 ( new_n1159 , pi024 , pi213 );
  or       g00783 ( new_n1160 , new_n1158 , new_n1159 );
  nand     g00784 ( new_n1161 , pi111 , pi212 );
  nor      g00785 ( new_n1162 , new_n1089 , new_n1161 );
  nand     g00786 ( new_n1163 , new_n1158 , new_n1159 );
  or       g00787 ( new_n1164 , new_n1162 , new_n1163 );
  nand     g00788 ( new_n1165 , new_n1160 , new_n1164 );
  and      g00789 ( new_n1166 , new_n1162 , new_n1163 );
  nor      g00790 ( new_n1167 , new_n1165 , new_n1166 );
  xnor     g00791 ( new_n1168 , new_n1157 , new_n1167 );
  xnor     g00792 ( new_n1169 , new_n1145 , new_n1168 );
  xor      g00793 ( new_n1170 , new_n1141 , new_n1169 );
  xor      g00794 ( new_n1171 , new_n1136 , new_n1170 );
  or       g00795 ( new_n1172 , new_n1132 , new_n1171 );
  nand     g00796 ( new_n1173 , new_n1131 , new_n1172 );
  nand g00797 ( new_n1174 , new_n1125 , new_n1125 );
  or       g00798 ( new_n1175 , new_n1123 , new_n1174 );
  nand     g00799 ( new_n1176 , new_n1124 , new_n1175 );
  nand     g00800 ( new_n1177 , pi081 , pi131 );
  xor      g00801 ( new_n1178 , new_n1176 , new_n1177 );
  nand     g00802 ( new_n1179 , pi077 , pi100 );
  nand     g00803 ( new_n1180 , pi133 , pi217 );
  nand     g00804 ( new_n1181 , pi052 , pi227 );
  xor      g00805 ( new_n1182 , new_n1180 , new_n1181 );
  xor      g00806 ( new_n1183 , new_n1179 , new_n1182 );
  xor      g00807 ( new_n1184 , new_n1178 , new_n1183 );
  nor      g00808 ( new_n1185 , new_n1125 , new_n1128 );
  xor      g00809 ( new_n1186 , new_n1184 , new_n1185 );
  xor      g00810 ( new_n1187 , new_n1173 , new_n1186 );
  nand     g00811 ( new_n1188 , new_n1141 , new_n1169 );
  nand     g00812 ( new_n1189 , new_n1136 , new_n1170 );
  nand     g00813 ( new_n1190 , new_n1188 , new_n1189 );
  and      g00814 ( new_n1191 , new_n1147 , new_n1155 );
  nand     g00815 ( new_n1192 , pi140 , pi161 );
  nand     g00816 ( new_n1193 , pi141 , pi242 );
  nand     g00817 ( new_n1194 , pi241 , pi252 );
  xor      g00818 ( new_n1195 , new_n1193 , new_n1194 );
  xor      g00819 ( new_n1196 , new_n1192 , new_n1195 );
  nor      g00820 ( new_n1197 , new_n1151 , new_n1147 );
  or       g00821 ( new_n1198 , new_n1153 , new_n1197 );
  nand     g00822 ( new_n1199 , pi121 , pi236 );
  xnor     g00823 ( new_n1200 , new_n1198 , new_n1199 );
  xor      g00824 ( new_n1201 , new_n1196 , new_n1200 );
  xnor     g00825 ( new_n1202 , new_n1191 , new_n1201 );
  nand g00826 ( new_n1203 , new_n1161 , new_n1161 );
  and      g00827 ( new_n1204 , new_n1203 , new_n1165 );
  nand     g00828 ( new_n1205 , pi104 , pi111 );
  nand     g00829 ( new_n1206 , pi013 , pi210 );
  nand     g00830 ( new_n1207 , pi024 , pi212 );
  xor      g00831 ( new_n1208 , new_n1206 , new_n1207 );
  xor      g00832 ( new_n1209 , new_n1205 , new_n1208 );
  nand     g00833 ( new_n1210 , new_n1160 , new_n1161 );
  nand     g00834 ( new_n1211 , new_n1163 , new_n1210 );
  nand     g00835 ( new_n1212 , pi213 , pi224 );
  xor      g00836 ( new_n1213 , new_n1211 , new_n1212 );
  xor      g00837 ( new_n1214 , new_n1209 , new_n1213 );
  xor      g00838 ( new_n1215 , new_n1204 , new_n1214 );
  xor      g00839 ( new_n1216 , new_n1202 , new_n1215 );
  nor      g00840 ( new_n1217 , new_n1157 , new_n1167 );
  nor      g00841 ( new_n1218 , new_n1145 , new_n1168 );
  nor      g00842 ( new_n1219 , new_n1217 , new_n1218 );
  xor      g00843 ( new_n1220 , new_n1216 , new_n1219 );
  nor      g00844 ( new_n1221 , new_n1101 , new_n1140 );
  nand     g00845 ( new_n1222 , pi125 , pi208 );
  nand     g00846 ( new_n1223 , pi035 , pi249 );
  nand     g00847 ( new_n1224 , pi139 , pi222 );
  xor      g00848 ( new_n1225 , new_n1223 , new_n1224 );
  xor      g00849 ( new_n1226 , new_n1222 , new_n1225 );
  nand     g00850 ( new_n1227 , pi168 , pi176 );
  nand     g00851 ( new_n1228 , new_n1099 , new_n1138 );
  nand     g00852 ( new_n1229 , new_n1137 , new_n1139 );
  nand     g00853 ( new_n1230 , new_n1228 , new_n1229 );
  xor      g00854 ( new_n1231 , new_n1227 , new_n1230 );
  xnor     g00855 ( new_n1232 , new_n1226 , new_n1231 );
  xor      g00856 ( new_n1233 , new_n1221 , new_n1232 );
  xor      g00857 ( new_n1234 , new_n1220 , new_n1233 );
  xor      g00858 ( new_n1235 , new_n1190 , new_n1234 );
  xor      g00859 ( po004 , new_n1187 , new_n1235 );
  nand     g00860 ( new_n1237 , pi071 , pi114 );
  nand     g00861 ( new_n1238 , pi091 , pi142 );
  nand     g00862 ( new_n1239 , new_n1237 , new_n1238 );
  nand     g00863 ( new_n1240 , pi169 , pi246 );
  xor      g00864 ( new_n1241 , new_n1237 , new_n1238 );
  nand     g00865 ( new_n1242 , new_n1240 , new_n1241 );
  nand     g00866 ( new_n1243 , new_n1239 , new_n1242 );
  nand     g00867 ( new_n1244 , pi101 , pi119 );
  nand g00868 ( new_n1245 , new_n1244 , new_n1244 );
  nand     g00869 ( new_n1246 , pi045 , pi225 );
  nand g00870 ( new_n1247 , new_n1246 , new_n1246 );
  nand     g00871 ( new_n1248 , new_n1245 , new_n1247 );
  nand     g00872 ( new_n1249 , pi044 , pi223 );
  nor      g00873 ( new_n1250 , new_n1248 , new_n1249 );
  xnor     g00874 ( new_n1251 , new_n1248 , new_n1249 );
  nand     g00875 ( new_n1252 , pi101 , pi250 );
  nand     g00876 ( new_n1253 , pi119 , pi177 );
  xor      g00877 ( new_n1254 , new_n1247 , new_n1253 );
  xor      g00878 ( new_n1255 , new_n1252 , new_n1254 );
  nand g00879 ( new_n1256 , new_n1255 , new_n1255 );
  nor      g00880 ( new_n1257 , new_n1251 , new_n1256 );
  nor      g00881 ( new_n1258 , new_n1250 , new_n1257 );
  nand     g00882 ( new_n1259 , new_n1246 , new_n1253 );
  nand g00883 ( new_n1260 , new_n1254 , new_n1254 );
  nand     g00884 ( new_n1261 , new_n1252 , new_n1260 );
  nand     g00885 ( new_n1262 , new_n1259 , new_n1261 );
  xor      g00886 ( new_n1263 , new_n1258 , new_n1262 );
  xor      g00887 ( new_n1264 , new_n1243 , new_n1263 );
  nand     g00888 ( new_n1265 , pi001 , pi136 );
  nand     g00889 ( new_n1266 , pi147 , pi192 );
  nand     g00890 ( new_n1267 , pi225 , pi250 );
  xor      g00891 ( new_n1268 , new_n1266 , new_n1267 );
  xor      g00892 ( new_n1269 , new_n1265 , new_n1268 );
  xor      g00893 ( new_n1270 , new_n1264 , new_n1269 );
  nand     g00894 ( new_n1271 , pi056 , pi219 );
  nand     g00895 ( new_n1272 , pi102 , pi136 );
  nor      g00896 ( new_n1273 , new_n1271 , new_n1272 );
  nand     g00897 ( new_n1274 , pi001 , pi027 );
  nand     g00898 ( new_n1275 , pi026 , pi102 );
  nand     g00899 ( new_n1276 , new_n1274 , new_n1275 );
  nand     g00900 ( new_n1277 , pi008 , pi219 );
  xor      g00901 ( new_n1278 , new_n1274 , new_n1275 );
  nand     g00902 ( new_n1279 , new_n1277 , new_n1278 );
  nand     g00903 ( new_n1280 , new_n1276 , new_n1279 );
  nand     g00904 ( new_n1281 , new_n1271 , new_n1280 );
  nand     g00905 ( new_n1282 , pi008 , pi102 );
  nand     g00906 ( new_n1283 , pi027 , pi122 );
  nand     g00907 ( new_n1284 , pi001 , pi026 );
  xor      g00908 ( new_n1285 , new_n1283 , new_n1284 );
  xor      g00909 ( new_n1286 , new_n1282 , new_n1285 );
  xor      g00910 ( new_n1287 , new_n1271 , new_n1280 );
  nand     g00911 ( new_n1288 , new_n1286 , new_n1287 );
  nand     g00912 ( new_n1289 , new_n1281 , new_n1288 );
  nand     g00913 ( new_n1290 , pi136 , pi219 );
  nand     g00914 ( new_n1291 , pi056 , pi102 );
  and      g00915 ( new_n1292 , new_n1290 , new_n1291 );
  nor      g00916 ( new_n1293 , new_n1273 , new_n1292 );
  nand     g00917 ( new_n1294 , new_n1283 , new_n1284 );
  nand     g00918 ( new_n1295 , new_n1282 , new_n1285 );
  nand     g00919 ( new_n1296 , new_n1294 , new_n1295 );
  nand     g00920 ( new_n1297 , pi001 , pi008 );
  nand     g00921 ( new_n1298 , pi027 , pi135 );
  nand     g00922 ( new_n1299 , pi026 , pi122 );
  nand     g00923 ( new_n1300 , new_n1298 , new_n1299 );
  nand     g00924 ( new_n1301 , pi026 , pi135 );
  nor      g00925 ( new_n1302 , new_n1283 , new_n1301 );
  nand g00926 ( new_n1303 , new_n1302 , new_n1302 );
  nand     g00927 ( new_n1304 , new_n1300 , new_n1303 );
  xor      g00928 ( new_n1305 , new_n1297 , new_n1304 );
  xor      g00929 ( new_n1306 , new_n1296 , new_n1305 );
  xor      g00930 ( new_n1307 , new_n1293 , new_n1306 );
  nor      g00931 ( new_n1308 , new_n1289 , new_n1307 );
  nand     g00932 ( new_n1309 , new_n1273 , new_n1308 );
  nand g00933 ( new_n1310 , new_n1306 , new_n1306 );
  nand     g00934 ( new_n1311 , new_n1293 , new_n1310 );
  nand g00935 ( new_n1312 , new_n1311 , new_n1311 );
  xor      g00936 ( new_n1313 , new_n1273 , new_n1308 );
  nor      g00937 ( new_n1314 , new_n1312 , new_n1313 );
  nand g00938 ( new_n1315 , new_n1314 , new_n1314 );
  nand     g00939 ( new_n1316 , pi008 , pi122 );
  nand     g00940 ( new_n1317 , pi027 , pi059 );
  xor      g00941 ( new_n1318 , new_n1316 , new_n1317 );
  xor      g00942 ( new_n1319 , new_n1301 , new_n1318 );
  nand     g00943 ( new_n1320 , pi001 , pi056 );
  xor      g00944 ( new_n1321 , new_n1302 , new_n1320 );
  xor      g00945 ( new_n1322 , new_n1319 , new_n1321 );
  nand     g00946 ( new_n1323 , new_n1297 , new_n1304 );
  nand     g00947 ( new_n1324 , new_n1296 , new_n1305 );
  nand     g00948 ( new_n1325 , new_n1323 , new_n1324 );
  nand     g00949 ( new_n1326 , pi087 , pi235 );
  nand     g00950 ( new_n1327 , pi096 , pi219 );
  xor      g00951 ( new_n1328 , new_n1272 , new_n1327 );
  xnor     g00952 ( new_n1329 , new_n1326 , new_n1328 );
  xor      g00953 ( new_n1330 , new_n1325 , new_n1329 );
  xnor     g00954 ( new_n1331 , new_n1322 , new_n1330 );
  nand     g00955 ( new_n1332 , new_n1315 , new_n1331 );
  nand     g00956 ( new_n1333 , new_n1309 , new_n1332 );
  nand     g00957 ( new_n1334 , pi114 , pi169 );
  xor      g00958 ( new_n1335 , new_n1333 , new_n1334 );
  xor      g00959 ( new_n1336 , new_n1270 , new_n1335 );
  nand     g00960 ( new_n1337 , pi027 , pi094 );
  nand     g00961 ( new_n1338 , new_n1316 , new_n1317 );
  nand     g00962 ( new_n1339 , new_n1301 , new_n1318 );
  nand     g00963 ( new_n1340 , new_n1338 , new_n1339 );
  xor      g00964 ( new_n1341 , new_n1337 , new_n1340 );
  xor      g00965 ( new_n1342 , new_n1336 , new_n1341 );
  nand     g00966 ( new_n1343 , pi075 , pi216 );
  nand     g00967 ( new_n1344 , pi151 , pi251 );
  nand     g00968 ( new_n1345 , pi142 , pi246 );
  nand     g00969 ( new_n1346 , pi164 , pi169 );
  nand     g00970 ( new_n1347 , pi032 , pi142 );
  and      g00971 ( new_n1348 , new_n1346 , new_n1347 );
  nand g00972 ( new_n1349 , new_n1348 , new_n1348 );
  nand     g00973 ( new_n1350 , pi071 , pi206 );
  or       g00974 ( new_n1351 , new_n1346 , new_n1347 );
  nand     g00975 ( new_n1352 , new_n1350 , new_n1351 );
  nand     g00976 ( new_n1353 , new_n1349 , new_n1352 );
  nand     g00977 ( new_n1354 , pi142 , pi145 );
  nand     g00978 ( new_n1355 , new_n1353 , new_n1354 );
  nand     g00979 ( new_n1356 , pi032 , pi071 );
  nand     g00980 ( new_n1357 , pi123 , pi164 );
  nand     g00981 ( new_n1358 , pi169 , pi206 );
  xor      g00982 ( new_n1359 , new_n1357 , new_n1358 );
  xor      g00983 ( new_n1360 , new_n1356 , new_n1359 );
  xor      g00984 ( new_n1361 , new_n1353 , new_n1354 );
  nand     g00985 ( new_n1362 , new_n1360 , new_n1361 );
  nand     g00986 ( new_n1363 , new_n1355 , new_n1362 );
  nor      g00987 ( new_n1364 , new_n1345 , new_n1363 );
  xor      g00988 ( new_n1365 , new_n1345 , new_n1363 );
  nand     g00989 ( new_n1366 , pi032 , pi169 );
  nand     g00990 ( new_n1367 , pi099 , pi164 );
  nand     g00991 ( new_n1368 , pi123 , pi206 );
  xor      g00992 ( new_n1369 , new_n1367 , new_n1368 );
  xor      g00993 ( new_n1370 , new_n1366 , new_n1369 );
  nand     g00994 ( new_n1371 , pi071 , pi145 );
  nand     g00995 ( new_n1372 , new_n1357 , new_n1358 );
  nand     g00996 ( new_n1373 , new_n1356 , new_n1359 );
  nand     g00997 ( new_n1374 , new_n1372 , new_n1373 );
  xor      g00998 ( new_n1375 , new_n1371 , new_n1374 );
  xnor     g00999 ( new_n1376 , new_n1370 , new_n1375 );
  nand     g01000 ( new_n1377 , new_n1365 , new_n1376 );
  nand g01001 ( new_n1378 , new_n1377 , new_n1377 );
  nor      g01002 ( new_n1379 , new_n1364 , new_n1378 );
  nand g01003 ( new_n1380 , new_n1379 , new_n1379 );
  nand     g01004 ( new_n1381 , new_n1371 , new_n1374 );
  nand     g01005 ( new_n1382 , new_n1370 , new_n1375 );
  nand     g01006 ( new_n1383 , new_n1381 , new_n1382 );
  nand     g01007 ( new_n1384 , pi071 , pi246 );
  nand     g01008 ( new_n1385 , pi145 , pi169 );
  nand     g01009 ( new_n1386 , new_n1384 , new_n1385 );
  nor      g01010 ( new_n1387 , new_n1240 , new_n1371 );
  nand g01011 ( new_n1388 , new_n1387 , new_n1387 );
  nand     g01012 ( new_n1389 , new_n1386 , new_n1388 );
  nand     g01013 ( new_n1390 , pi099 , pi206 );
  nand     g01014 ( new_n1391 , pi023 , pi164 );
  nand     g01015 ( new_n1392 , new_n1390 , new_n1391 );
  nand     g01016 ( new_n1393 , pi023 , pi206 );
  or       g01017 ( new_n1394 , new_n1367 , new_n1393 );
  nand     g01018 ( new_n1395 , new_n1392 , new_n1394 );
  nand     g01019 ( new_n1396 , pi032 , pi123 );
  nand     g01020 ( new_n1397 , new_n1367 , new_n1368 );
  nand     g01021 ( new_n1398 , new_n1366 , new_n1369 );
  nand     g01022 ( new_n1399 , new_n1397 , new_n1398 );
  xor      g01023 ( new_n1400 , new_n1396 , new_n1399 );
  xor      g01024 ( new_n1401 , new_n1395 , new_n1400 );
  xor      g01025 ( new_n1402 , new_n1389 , new_n1401 );
  xnor     g01026 ( new_n1403 , new_n1383 , new_n1402 );
  nand     g01027 ( new_n1404 , new_n1380 , new_n1403 );
  nand     g01028 ( new_n1405 , pi123 , pi145 );
  xnor     g01029 ( new_n1406 , new_n1394 , new_n1405 );
  nand     g01030 ( new_n1407 , pi032 , pi099 );
  nand     g01031 ( new_n1408 , pi155 , pi164 );
  xor      g01032 ( new_n1409 , new_n1393 , new_n1408 );
  xor      g01033 ( new_n1410 , new_n1407 , new_n1409 );
  xor      g01034 ( new_n1411 , new_n1406 , new_n1410 );
  nand     g01035 ( new_n1412 , new_n1396 , new_n1399 );
  nand     g01036 ( new_n1413 , new_n1395 , new_n1400 );
  nand     g01037 ( new_n1414 , new_n1412 , new_n1413 );
  xnor     g01038 ( new_n1415 , new_n1240 , new_n1241 );
  xor      g01039 ( new_n1416 , new_n1414 , new_n1415 );
  xor      g01040 ( new_n1417 , new_n1411 , new_n1416 );
  nand     g01041 ( new_n1418 , new_n1389 , new_n1401 );
  nand     g01042 ( new_n1419 , new_n1383 , new_n1402 );
  nand     g01043 ( new_n1420 , new_n1418 , new_n1419 );
  xor      g01044 ( new_n1421 , new_n1388 , new_n1420 );
  xor      g01045 ( new_n1422 , new_n1417 , new_n1421 );
  nor      g01046 ( new_n1423 , new_n1404 , new_n1422 );
  and      g01047 ( new_n1424 , pi142 , pi164 );
  nor      g01048 ( new_n1425 , new_n1424 , new_n1350 );
  and      g01049 ( new_n1426 , new_n1349 , new_n1351 );
  nor      g01050 ( new_n1427 , new_n1425 , new_n1426 );
  nand g01051 ( new_n1428 , new_n1427 , new_n1427 );
  nor      g01052 ( new_n1429 , new_n1350 , new_n1428 );
  xor      g01053 ( new_n1430 , new_n1360 , new_n1361 );
  nand g01054 ( new_n1431 , new_n1430 , new_n1430 );
  nand     g01055 ( new_n1432 , new_n1429 , new_n1431 );
  nand g01056 ( new_n1433 , new_n1432 , new_n1432 );
  xor      g01057 ( new_n1434 , new_n1365 , new_n1376 );
  nand     g01058 ( new_n1435 , new_n1433 , new_n1434 );
  nand     g01059 ( new_n1436 , pi114 , pi142 );
  nand     g01060 ( new_n1437 , new_n1435 , new_n1436 );
  xor      g01061 ( new_n1438 , new_n1435 , new_n1436 );
  xor      g01062 ( new_n1439 , new_n1379 , new_n1403 );
  nand     g01063 ( new_n1440 , new_n1438 , new_n1439 );
  nand     g01064 ( new_n1441 , new_n1437 , new_n1440 );
  xor      g01065 ( new_n1442 , new_n1404 , new_n1422 );
  nand g01066 ( new_n1443 , new_n1442 , new_n1442 );
  nor      g01067 ( new_n1444 , new_n1441 , new_n1443 );
  or       g01068 ( new_n1445 , new_n1423 , new_n1444 );
  xor      g01069 ( new_n1446 , new_n1344 , new_n1445 );
  xor      g01070 ( new_n1447 , new_n1343 , new_n1446 );
  nand     g01071 ( new_n1448 , pi060 , pi250 );
  nand     g01072 ( new_n1449 , new_n1244 , new_n1448 );
  nand     g01073 ( new_n1450 , pi045 , pi223 );
  xor      g01074 ( new_n1451 , new_n1245 , new_n1448 );
  nand g01075 ( new_n1452 , new_n1451 , new_n1451 );
  nand     g01076 ( new_n1453 , new_n1450 , new_n1452 );
  nand     g01077 ( new_n1454 , new_n1449 , new_n1453 );
  nand     g01078 ( new_n1455 , pi119 , pi225 );
  nand     g01079 ( new_n1456 , pi045 , pi101 );
  nand     g01080 ( new_n1457 , new_n1455 , new_n1456 );
  nand     g01081 ( new_n1458 , new_n1248 , new_n1457 );
  nand     g01082 ( new_n1459 , new_n1454 , new_n1458 );
  nand     g01083 ( new_n1460 , pi223 , pi250 );
  xor      g01084 ( new_n1461 , new_n1454 , new_n1458 );
  nand     g01085 ( new_n1462 , new_n1460 , new_n1461 );
  nand     g01086 ( new_n1463 , new_n1459 , new_n1462 );
  nand     g01087 ( new_n1464 , pi054 , pi060 );
  nand     g01088 ( new_n1465 , pi160 , pi248 );
  nand     g01089 ( new_n1466 , pi020 , pi072 );
  xor      g01090 ( new_n1467 , new_n1465 , new_n1466 );
  xor      g01091 ( new_n1468 , new_n1464 , new_n1467 );
  nor      g01092 ( new_n1469 , new_n1463 , new_n1468 );
  xor      g01093 ( new_n1470 , new_n1251 , new_n1255 );
  xnor     g01094 ( new_n1471 , new_n1463 , new_n1468 );
  nor      g01095 ( new_n1472 , new_n1470 , new_n1471 );
  nor      g01096 ( new_n1473 , new_n1469 , new_n1472 );
  nand     g01097 ( new_n1474 , pi011 , pi138 );
  xor      g01098 ( new_n1475 , new_n1473 , new_n1474 );
  xor      g01099 ( new_n1476 , new_n1447 , new_n1475 );
  nand     g01100 ( new_n1477 , pi087 , pi096 );
  nand     g01101 ( new_n1478 , pi056 , pi087 );
  nand     g01102 ( new_n1479 , pi008 , pi087 );
  nand     g01103 ( new_n1480 , pi026 , pi219 );
  nand     g01104 ( new_n1481 , new_n1479 , new_n1480 );
  nand     g01105 ( new_n1482 , pi027 , pi102 );
  xor      g01106 ( new_n1483 , new_n1479 , new_n1480 );
  nand     g01107 ( new_n1484 , new_n1482 , new_n1483 );
  nand     g01108 ( new_n1485 , new_n1481 , new_n1484 );
  nor      g01109 ( new_n1486 , new_n1478 , new_n1485 );
  xor      g01110 ( new_n1487 , new_n1478 , new_n1485 );
  nand g01111 ( new_n1488 , new_n1487 , new_n1487 );
  xor      g01112 ( new_n1489 , new_n1277 , new_n1278 );
  nor      g01113 ( new_n1490 , new_n1488 , new_n1489 );
  nor      g01114 ( new_n1491 , new_n1486 , new_n1490 );
  nand     g01115 ( new_n1492 , pi087 , pi136 );
  xor      g01116 ( new_n1493 , new_n1286 , new_n1287 );
  xor      g01117 ( new_n1494 , new_n1492 , new_n1493 );
  nand g01118 ( new_n1495 , new_n1494 , new_n1494 );
  xor      g01119 ( new_n1496 , new_n1491 , new_n1495 );
  xor      g01120 ( new_n1497 , new_n1482 , new_n1483 );
  nand g01121 ( new_n1498 , new_n1497 , new_n1497 );
  nor      g01122 ( new_n1499 , new_n1079 , new_n1480 );
  nand     g01123 ( new_n1500 , new_n1498 , new_n1499 );
  xor      g01124 ( new_n1501 , new_n1487 , new_n1489 );
  nor      g01125 ( new_n1502 , new_n1500 , new_n1501 );
  nand     g01126 ( new_n1503 , new_n1496 , new_n1502 );
  xor      g01127 ( new_n1504 , new_n1477 , new_n1503 );
  nand g01128 ( new_n1505 , new_n1504 , new_n1504 );
  nor      g01129 ( new_n1506 , new_n1492 , new_n1493 );
  nor      g01130 ( new_n1507 , new_n1491 , new_n1495 );
  nor      g01131 ( new_n1508 , new_n1506 , new_n1507 );
  xnor     g01132 ( new_n1509 , new_n1289 , new_n1307 );
  xor      g01133 ( new_n1510 , new_n1508 , new_n1509 );
  xor      g01134 ( new_n1511 , new_n1505 , new_n1510 );
  nand g01135 ( new_n1512 , new_n1511 , new_n1511 );
  xor      g01136 ( new_n1513 , new_n1432 , new_n1434 );
  nand g01137 ( new_n1514 , new_n1513 , new_n1513 );
  xnor     g01138 ( new_n1515 , new_n1500 , new_n1501 );
  nand g01139 ( new_n1516 , new_n1515 , new_n1515 );
  nand     g01140 ( new_n1517 , pi026 , pi087 );
  nand     g01141 ( new_n1518 , pi027 , pi219 );
  and      g01142 ( new_n1519 , new_n1517 , new_n1518 );
  or       g01143 ( new_n1520 , new_n1499 , new_n1519 );
  nand     g01144 ( new_n1521 , pi071 , pi164 );
  nand     g01145 ( new_n1522 , pi142 , pi206 );
  xnor     g01146 ( new_n1523 , new_n1521 , new_n1522 );
  nand     g01147 ( new_n1524 , new_n1520 , new_n1523 );
  nor      g01148 ( new_n1525 , new_n1079 , new_n1080 );
  xnor     g01149 ( new_n1526 , new_n1520 , new_n1523 );
  or       g01150 ( new_n1527 , new_n1525 , new_n1526 );
  nand     g01151 ( new_n1528 , new_n1524 , new_n1527 );
  nand     g01152 ( new_n1529 , new_n1349 , new_n1425 );
  nand     g01153 ( new_n1530 , new_n1428 , new_n1529 );
  and      g01154 ( new_n1531 , new_n1528 , new_n1530 );
  xnor     g01155 ( new_n1532 , new_n1528 , new_n1530 );
  xor      g01156 ( new_n1533 , new_n1497 , new_n1499 );
  nand g01157 ( new_n1534 , new_n1533 , new_n1533 );
  nor      g01158 ( new_n1535 , new_n1532 , new_n1534 );
  nor      g01159 ( new_n1536 , new_n1531 , new_n1535 );
  nor      g01160 ( new_n1537 , new_n1516 , new_n1536 );
  xor      g01161 ( new_n1538 , new_n1429 , new_n1431 );
  xor      g01162 ( new_n1539 , new_n1515 , new_n1536 );
  nor      g01163 ( new_n1540 , new_n1538 , new_n1539 );
  nor      g01164 ( new_n1541 , new_n1537 , new_n1540 );
  nor      g01165 ( new_n1542 , new_n1514 , new_n1541 );
  xor      g01166 ( new_n1543 , new_n1496 , new_n1502 );
  xor      g01167 ( new_n1544 , new_n1513 , new_n1541 );
  nor      g01168 ( new_n1545 , new_n1543 , new_n1544 );
  nor      g01169 ( new_n1546 , new_n1542 , new_n1545 );
  nor      g01170 ( new_n1547 , new_n1512 , new_n1546 );
  xor      g01171 ( new_n1548 , new_n1438 , new_n1439 );
  nand g01172 ( new_n1549 , new_n1548 , new_n1548 );
  xor      g01173 ( new_n1550 , new_n1511 , new_n1546 );
  nor      g01174 ( new_n1551 , new_n1549 , new_n1550 );
  nor      g01175 ( new_n1552 , new_n1547 , new_n1551 );
  nand     g01176 ( new_n1553 , new_n1477 , new_n1503 );
  or       g01177 ( new_n1554 , new_n1505 , new_n1510 );
  nand     g01178 ( new_n1555 , new_n1553 , new_n1554 );
  nor      g01179 ( new_n1556 , new_n1508 , new_n1509 );
  xor      g01180 ( new_n1557 , new_n1314 , new_n1331 );
  xor      g01181 ( new_n1558 , new_n1556 , new_n1557 );
  xor      g01182 ( new_n1559 , new_n1555 , new_n1558 );
  nand     g01183 ( new_n1560 , new_n1552 , new_n1559 );
  xor      g01184 ( new_n1561 , new_n1552 , new_n1559 );
  xor      g01185 ( new_n1562 , new_n1441 , new_n1443 );
  nand     g01186 ( new_n1563 , new_n1561 , new_n1562 );
  nand     g01187 ( new_n1564 , new_n1560 , new_n1563 );
  nand     g01188 ( new_n1565 , new_n1465 , new_n1466 );
  nand     g01189 ( new_n1566 , new_n1464 , new_n1467 );
  nand     g01190 ( new_n1567 , new_n1565 , new_n1566 );
  nand     g01191 ( new_n1568 , pi086 , pi164 );
  xnor     g01192 ( new_n1569 , new_n1567 , new_n1568 );
  xor      g01193 ( new_n1570 , new_n1564 , new_n1569 );
  xor      g01194 ( new_n1571 , new_n1476 , new_n1570 );
  xor      g01195 ( new_n1572 , new_n1342 , new_n1571 );
  nand     g01196 ( new_n1573 , pi020 , pi248 );
  nand g01197 ( new_n1574 , new_n1556 , new_n1556 );
  nand     g01198 ( new_n1575 , new_n1574 , new_n1557 );
  nand g01199 ( new_n1576 , new_n1558 , new_n1558 );
  nand     g01200 ( new_n1577 , new_n1555 , new_n1576 );
  nand     g01201 ( new_n1578 , new_n1575 , new_n1577 );
  nor      g01202 ( new_n1579 , new_n1303 , new_n1320 );
  nor      g01203 ( new_n1580 , new_n1319 , new_n1321 );
  nor      g01204 ( new_n1581 , new_n1579 , new_n1580 );
  nand     g01205 ( new_n1582 , pi138 , pi166 );
  nand     g01206 ( new_n1583 , pi093 , pi182 );
  nand     g01207 ( new_n1584 , new_n1582 , new_n1583 );
  nand     g01208 ( new_n1585 , pi041 , pi075 );
  xor      g01209 ( new_n1586 , new_n1582 , new_n1583 );
  nand     g01210 ( new_n1587 , new_n1585 , new_n1586 );
  nand     g01211 ( new_n1588 , new_n1584 , new_n1587 );
  nand     g01212 ( new_n1589 , pi026 , pi059 );
  nand     g01213 ( new_n1590 , pi009 , pi160 );
  xor      g01214 ( new_n1591 , new_n1589 , new_n1590 );
  xor      g01215 ( new_n1592 , new_n1588 , new_n1591 );
  xor      g01216 ( new_n1593 , new_n1581 , new_n1592 );
  nand     g01217 ( new_n1594 , new_n1272 , new_n1327 );
  nand     g01218 ( new_n1595 , new_n1326 , new_n1328 );
  nand     g01219 ( new_n1596 , new_n1594 , new_n1595 );
  nand     g01220 ( new_n1597 , pi087 , pi110 );
  nand     g01221 ( new_n1598 , pi008 , pi135 );
  xor      g01222 ( new_n1599 , new_n1597 , new_n1598 );
  xor      g01223 ( new_n1600 , new_n1596 , new_n1599 );
  xor      g01224 ( new_n1601 , new_n1593 , new_n1600 );
  xor      g01225 ( new_n1602 , new_n1578 , new_n1601 );
  xor      g01226 ( new_n1603 , new_n1573 , new_n1602 );
  nand     g01227 ( new_n1604 , pi020 , pi044 );
  nor      g01228 ( new_n1605 , new_n1464 , new_n1604 );
  nand     g01229 ( new_n1606 , pi045 , pi060 );
  nand     g01230 ( new_n1607 , pi119 , pi223 );
  nand     g01231 ( new_n1608 , new_n1606 , new_n1607 );
  nand     g01232 ( new_n1609 , pi020 , pi250 );
  xor      g01233 ( new_n1610 , new_n1606 , new_n1607 );
  nand     g01234 ( new_n1611 , new_n1609 , new_n1610 );
  nand     g01235 ( new_n1612 , new_n1608 , new_n1611 );
  nand     g01236 ( new_n1613 , new_n1604 , new_n1612 );
  xor      g01237 ( new_n1614 , new_n1450 , new_n1451 );
  nand g01238 ( new_n1615 , new_n1614 , new_n1614 );
  xor      g01239 ( new_n1616 , new_n1604 , new_n1612 );
  nand     g01240 ( new_n1617 , new_n1615 , new_n1616 );
  nand     g01241 ( new_n1618 , new_n1613 , new_n1617 );
  nand     g01242 ( new_n1619 , pi044 , pi060 );
  nand     g01243 ( new_n1620 , pi020 , pi054 );
  nand     g01244 ( new_n1621 , new_n1619 , new_n1620 );
  nand g01245 ( new_n1622 , new_n1621 , new_n1621 );
  nor      g01246 ( new_n1623 , new_n1605 , new_n1622 );
  nand g01247 ( new_n1624 , new_n1623 , new_n1623 );
  nand     g01248 ( new_n1625 , new_n1618 , new_n1624 );
  xor      g01249 ( new_n1626 , new_n1460 , new_n1461 );
  xor      g01250 ( new_n1627 , new_n1618 , new_n1624 );
  nand     g01251 ( new_n1628 , new_n1626 , new_n1627 );
  nand     g01252 ( new_n1629 , new_n1625 , new_n1628 );
  xor      g01253 ( new_n1630 , new_n1605 , new_n1629 );
  xor      g01254 ( new_n1631 , new_n1470 , new_n1471 );
  xor      g01255 ( new_n1632 , new_n1630 , new_n1631 );
  nand     g01256 ( new_n1633 , pi054 , pi160 );
  xor      g01257 ( new_n1634 , new_n1614 , new_n1616 );
  nand g01258 ( new_n1635 , new_n1634 , new_n1634 );
  nor      g01259 ( new_n1636 , new_n1633 , new_n1635 );
  nand     g01260 ( new_n1637 , pi020 , pi045 );
  nand g01261 ( new_n1638 , new_n1637 , new_n1637 );
  nand     g01262 ( new_n1639 , pi060 , pi119 );
  nand     g01263 ( new_n1640 , pi160 , pi250 );
  nor      g01264 ( new_n1641 , new_n1639 , new_n1640 );
  or       g01265 ( new_n1642 , new_n1638 , new_n1641 );
  nand     g01266 ( new_n1643 , new_n1639 , new_n1640 );
  nand     g01267 ( new_n1644 , new_n1642 , new_n1643 );
  nand     g01268 ( new_n1645 , pi044 , pi160 );
  nor      g01269 ( new_n1646 , new_n1644 , new_n1645 );
  xor      g01270 ( new_n1647 , new_n1609 , new_n1610 );
  xor      g01271 ( new_n1648 , new_n1644 , new_n1645 );
  nand g01272 ( new_n1649 , new_n1648 , new_n1648 );
  nor      g01273 ( new_n1650 , new_n1647 , new_n1649 );
  nor      g01274 ( new_n1651 , new_n1646 , new_n1650 );
  xor      g01275 ( new_n1652 , new_n1633 , new_n1634 );
  nor      g01276 ( new_n1653 , new_n1651 , new_n1652 );
  nor      g01277 ( new_n1654 , new_n1636 , new_n1653 );
  xor      g01278 ( new_n1655 , new_n1626 , new_n1627 );
  nor      g01279 ( new_n1656 , new_n1654 , new_n1655 );
  nand g01280 ( new_n1657 , new_n1656 , new_n1656 );
  nor      g01281 ( new_n1658 , new_n1632 , new_n1657 );
  xor      g01282 ( new_n1659 , new_n1632 , new_n1656 );
  nand     g01283 ( new_n1660 , pi072 , pi160 );
  xor      g01284 ( new_n1661 , new_n1651 , new_n1652 );
  nor      g01285 ( new_n1662 , new_n1077 , new_n1637 );
  nor      g01286 ( new_n1663 , new_n1643 , new_n1662 );
  nor      g01287 ( new_n1664 , new_n1641 , new_n1663 );
  nor      g01288 ( new_n1665 , new_n1637 , new_n1664 );
  xor      g01289 ( new_n1666 , new_n1647 , new_n1648 );
  nand g01290 ( new_n1667 , new_n1666 , new_n1666 );
  nand     g01291 ( new_n1668 , new_n1665 , new_n1667 );
  nand g01292 ( new_n1669 , new_n1668 , new_n1668 );
  nand     g01293 ( new_n1670 , new_n1661 , new_n1669 );
  nand     g01294 ( new_n1671 , new_n1660 , new_n1670 );
  xor      g01295 ( new_n1672 , new_n1660 , new_n1670 );
  xnor     g01296 ( new_n1673 , new_n1654 , new_n1655 );
  nand     g01297 ( new_n1674 , new_n1672 , new_n1673 );
  nand     g01298 ( new_n1675 , new_n1671 , new_n1674 );
  nor      g01299 ( new_n1676 , new_n1659 , new_n1675 );
  nor      g01300 ( new_n1677 , new_n1658 , new_n1676 );
  nand g01301 ( new_n1678 , new_n1325 , new_n1325 );
  nor      g01302 ( new_n1679 , new_n1678 , new_n1329 );
  nor      g01303 ( new_n1680 , new_n1322 , new_n1330 );
  nor      g01304 ( new_n1681 , new_n1679 , new_n1680 );
  nand g01305 ( new_n1682 , new_n1414 , new_n1414 );
  nor      g01306 ( new_n1683 , new_n1682 , new_n1415 );
  nor      g01307 ( new_n1684 , new_n1411 , new_n1416 );
  nor      g01308 ( new_n1685 , new_n1683 , new_n1684 );
  xor      g01309 ( new_n1686 , new_n1681 , new_n1685 );
  xor      g01310 ( new_n1687 , new_n1677 , new_n1686 );
  nand     g01311 ( new_n1688 , pi166 , pi182 );
  nand     g01312 ( new_n1689 , pi041 , pi093 );
  xor      g01313 ( new_n1690 , new_n1688 , new_n1689 );
  nand g01314 ( new_n1691 , new_n1629 , new_n1629 );
  nand     g01315 ( new_n1692 , new_n1605 , new_n1691 );
  nand g01316 ( new_n1693 , new_n1630 , new_n1630 );
  nand     g01317 ( new_n1694 , new_n1693 , new_n1631 );
  nand     g01318 ( new_n1695 , new_n1692 , new_n1694 );
  nand     g01319 ( new_n1696 , pi096 , pi102 );
  nand     g01320 ( new_n1697 , pi219 , pi235 );
  xor      g01321 ( new_n1698 , new_n1696 , new_n1697 );
  xor      g01322 ( new_n1699 , new_n1695 , new_n1698 );
  xor      g01323 ( new_n1700 , new_n1690 , new_n1699 );
  xor      g01324 ( new_n1701 , new_n1687 , new_n1700 );
  nand     g01325 ( new_n1702 , pi071 , pi091 );
  nand     g01326 ( new_n1703 , pi123 , pi246 );
  nor      g01327 ( new_n1704 , new_n1394 , new_n1405 );
  nor      g01328 ( new_n1705 , new_n1406 , new_n1410 );
  or       g01329 ( new_n1706 , new_n1704 , new_n1705 );
  xor      g01330 ( new_n1707 , new_n1703 , new_n1706 );
  nand     g01331 ( new_n1708 , pi054 , pi223 );
  nand     g01332 ( new_n1709 , pi076 , pi147 );
  nand     g01333 ( new_n1710 , pi079 , pi151 );
  nor      g01334 ( new_n1711 , new_n1709 , new_n1710 );
  nand g01335 ( new_n1712 , new_n1711 , new_n1711 );
  nand     g01336 ( new_n1713 , pi097 , pi216 );
  nor      g01337 ( new_n1714 , new_n1712 , new_n1713 );
  nand     g01338 ( new_n1715 , pi019 , pi076 );
  nand     g01339 ( new_n1716 , pi147 , pi251 );
  xor      g01340 ( new_n1717 , new_n1715 , new_n1716 );
  xor      g01341 ( new_n1718 , new_n1710 , new_n1717 );
  xor      g01342 ( new_n1719 , new_n1711 , new_n1713 );
  nor      g01343 ( new_n1720 , new_n1718 , new_n1719 );
  nor      g01344 ( new_n1721 , new_n1714 , new_n1720 );
  xor      g01345 ( new_n1722 , new_n1708 , new_n1721 );
  nand     g01346 ( new_n1723 , pi056 , pi122 );
  nand     g01347 ( new_n1724 , pi099 , pi145 );
  xor      g01348 ( new_n1725 , new_n1723 , new_n1724 );
  xor      g01349 ( new_n1726 , new_n1722 , new_n1725 );
  xor      g01350 ( new_n1727 , new_n1707 , new_n1726 );
  xnor     g01351 ( new_n1728 , new_n1702 , new_n1727 );
  nand     g01352 ( new_n1729 , new_n1393 , new_n1408 );
  nand     g01353 ( new_n1730 , new_n1407 , new_n1409 );
  nand     g01354 ( new_n1731 , new_n1729 , new_n1730 );
  nand     g01355 ( new_n1732 , pi075 , pi138 );
  nand     g01356 ( new_n1733 , pi097 , pi138 );
  nand     g01357 ( new_n1734 , pi019 , pi138 );
  nand     g01358 ( new_n1735 , pi151 , pi182 );
  nand     g01359 ( new_n1736 , new_n1734 , new_n1735 );
  xor      g01360 ( new_n1737 , new_n1734 , new_n1735 );
  nand     g01361 ( new_n1738 , pi041 , pi147 );
  nand     g01362 ( new_n1739 , new_n1737 , new_n1738 );
  nand     g01363 ( new_n1740 , new_n1736 , new_n1739 );
  nor      g01364 ( new_n1741 , new_n1733 , new_n1740 );
  nand     g01365 ( new_n1742 , pi019 , pi182 );
  nand     g01366 ( new_n1743 , pi147 , pi216 );
  nand     g01367 ( new_n1744 , pi041 , pi151 );
  xor      g01368 ( new_n1745 , new_n1743 , new_n1744 );
  xor      g01369 ( new_n1746 , new_n1742 , new_n1745 );
  nand g01370 ( new_n1747 , new_n1746 , new_n1746 );
  xor      g01371 ( new_n1748 , new_n1733 , new_n1740 );
  and      g01372 ( new_n1749 , new_n1747 , new_n1748 );
  nor      g01373 ( new_n1750 , new_n1741 , new_n1749 );
  nor      g01374 ( new_n1751 , new_n1732 , new_n1750 );
  nand g01375 ( new_n1752 , new_n1751 , new_n1751 );
  xor      g01376 ( new_n1753 , new_n1732 , new_n1750 );
  nand     g01377 ( new_n1754 , pi151 , pi216 );
  nand     g01378 ( new_n1755 , pi019 , pi041 );
  xor      g01379 ( new_n1756 , new_n1709 , new_n1755 );
  xor      g01380 ( new_n1757 , new_n1754 , new_n1756 );
  nand     g01381 ( new_n1758 , pi097 , pi182 );
  nand     g01382 ( new_n1759 , new_n1743 , new_n1744 );
  nand     g01383 ( new_n1760 , new_n1742 , new_n1745 );
  nand     g01384 ( new_n1761 , new_n1759 , new_n1760 );
  xor      g01385 ( new_n1762 , new_n1758 , new_n1761 );
  xnor     g01386 ( new_n1763 , new_n1757 , new_n1762 );
  nand     g01387 ( new_n1764 , new_n1753 , new_n1763 );
  nand     g01388 ( new_n1765 , new_n1752 , new_n1764 );
  nand     g01389 ( new_n1766 , new_n1758 , new_n1761 );
  nand     g01390 ( new_n1767 , new_n1757 , new_n1762 );
  nand     g01391 ( new_n1768 , new_n1766 , new_n1767 );
  nor      g01392 ( new_n1769 , new_n1758 , new_n1585 );
  nand     g01393 ( new_n1770 , pi041 , pi097 );
  nand     g01394 ( new_n1771 , pi075 , pi182 );
  and      g01395 ( new_n1772 , new_n1770 , new_n1771 );
  nor      g01396 ( new_n1773 , new_n1769 , new_n1772 );
  nand     g01397 ( new_n1774 , pi019 , pi216 );
  nand     g01398 ( new_n1775 , new_n1709 , new_n1755 );
  nand     g01399 ( new_n1776 , new_n1754 , new_n1756 );
  nand     g01400 ( new_n1777 , new_n1775 , new_n1776 );
  nand     g01401 ( new_n1778 , pi079 , pi147 );
  nand     g01402 ( new_n1779 , pi076 , pi151 );
  nand     g01403 ( new_n1780 , new_n1778 , new_n1779 );
  nand     g01404 ( new_n1781 , new_n1712 , new_n1780 );
  xor      g01405 ( new_n1782 , new_n1777 , new_n1781 );
  xor      g01406 ( new_n1783 , new_n1774 , new_n1782 );
  xor      g01407 ( new_n1784 , new_n1773 , new_n1783 );
  xor      g01408 ( new_n1785 , new_n1768 , new_n1784 );
  and      g01409 ( new_n1786 , new_n1765 , new_n1785 );
  nand g01410 ( new_n1787 , new_n1786 , new_n1786 );
  nor      g01411 ( new_n1788 , new_n1768 , new_n1784 );
  nand g01412 ( new_n1789 , new_n1788 , new_n1788 );
  nand g01413 ( new_n1790 , new_n1773 , new_n1773 );
  nor      g01414 ( new_n1791 , new_n1790 , new_n1783 );
  nor      g01415 ( new_n1792 , new_n1769 , new_n1791 );
  nand     g01416 ( new_n1793 , new_n1789 , new_n1792 );
  nand     g01417 ( new_n1794 , new_n1769 , new_n1788 );
  nand     g01418 ( new_n1795 , new_n1793 , new_n1794 );
  xor      g01419 ( new_n1796 , new_n1718 , new_n1719 );
  nand     g01420 ( new_n1797 , new_n1777 , new_n1781 );
  nand     g01421 ( new_n1798 , new_n1774 , new_n1782 );
  nand     g01422 ( new_n1799 , new_n1797 , new_n1798 );
  xnor     g01423 ( new_n1800 , new_n1585 , new_n1586 );
  xor      g01424 ( new_n1801 , new_n1799 , new_n1800 );
  xnor     g01425 ( new_n1802 , new_n1796 , new_n1801 );
  xor      g01426 ( new_n1803 , new_n1795 , new_n1802 );
  nor      g01427 ( new_n1804 , new_n1787 , new_n1803 );
  nand     g01428 ( new_n1805 , pi093 , pi138 );
  xor      g01429 ( new_n1806 , new_n1753 , new_n1763 );
  xor      g01430 ( new_n1807 , new_n1746 , new_n1748 );
  xor      g01431 ( new_n1808 , new_n1737 , new_n1738 );
  nor      g01432 ( new_n1809 , new_n1078 , new_n1735 );
  nand g01433 ( new_n1810 , new_n1809 , new_n1809 );
  nor      g01434 ( new_n1811 , new_n1808 , new_n1810 );
  nand g01435 ( new_n1812 , new_n1811 , new_n1811 );
  nor      g01436 ( new_n1813 , new_n1807 , new_n1812 );
  nand     g01437 ( new_n1814 , new_n1806 , new_n1813 );
  nand     g01438 ( new_n1815 , new_n1805 , new_n1814 );
  xor      g01439 ( new_n1816 , new_n1805 , new_n1814 );
  xnor     g01440 ( new_n1817 , new_n1765 , new_n1785 );
  nand     g01441 ( new_n1818 , new_n1816 , new_n1817 );
  nand     g01442 ( new_n1819 , new_n1815 , new_n1818 );
  xor      g01443 ( new_n1820 , new_n1786 , new_n1803 );
  nor      g01444 ( new_n1821 , new_n1819 , new_n1820 );
  nor      g01445 ( new_n1822 , new_n1804 , new_n1821 );
  nand     g01446 ( new_n1823 , pi119 , pi137 );
  xor      g01447 ( new_n1824 , new_n1822 , new_n1823 );
  xor      g01448 ( new_n1825 , new_n1731 , new_n1824 );
  xor      g01449 ( new_n1826 , new_n1728 , new_n1825 );
  xor      g01450 ( new_n1827 , new_n1701 , new_n1826 );
  xor      g01451 ( new_n1828 , new_n1603 , new_n1827 );
  xor      g01452 ( new_n1829 , new_n1665 , new_n1667 );
  or       g01453 ( new_n1830 , new_n1078 , new_n1081 );
  nand     g01454 ( new_n1831 , pi138 , pi151 );
  nand     g01455 ( new_n1832 , pi147 , pi182 );
  and      g01456 ( new_n1833 , new_n1831 , new_n1832 );
  or       g01457 ( new_n1834 , new_n1809 , new_n1833 );
  or       g01458 ( new_n1835 , new_n1830 , new_n1834 );
  xor      g01459 ( new_n1836 , new_n1525 , new_n1526 );
  xnor     g01460 ( new_n1837 , new_n1830 , new_n1834 );
  or       g01461 ( new_n1838 , new_n1836 , new_n1837 );
  and      g01462 ( new_n1839 , new_n1835 , new_n1838 );
  xor      g01463 ( new_n1840 , new_n1808 , new_n1809 );
  xor      g01464 ( new_n1841 , new_n1839 , new_n1840 );
  xor      g01465 ( new_n1842 , new_n1532 , new_n1533 );
  xnor     g01466 ( new_n1843 , new_n1841 , new_n1842 );
  nand     g01467 ( new_n1844 , new_n1077 , new_n1082 );
  nand g01468 ( new_n1845 , new_n1844 , new_n1844 );
  nand     g01469 ( new_n1846 , pi045 , pi160 );
  nand     g01470 ( new_n1847 , pi020 , pi119 );
  xor      g01471 ( new_n1848 , new_n1846 , new_n1847 );
  nor      g01472 ( new_n1849 , new_n1845 , new_n1848 );
  xor      g01473 ( new_n1850 , new_n1844 , new_n1848 );
  xor      g01474 ( new_n1851 , new_n1836 , new_n1837 );
  nor      g01475 ( new_n1852 , new_n1850 , new_n1851 );
  or       g01476 ( new_n1853 , new_n1849 , new_n1852 );
  nor      g01477 ( new_n1854 , new_n1843 , new_n1853 );
  xnor     g01478 ( new_n1855 , new_n1843 , new_n1853 );
  nand     g01479 ( new_n1856 , new_n1643 , new_n1662 );
  nand     g01480 ( new_n1857 , new_n1664 , new_n1856 );
  nor      g01481 ( new_n1858 , new_n1855 , new_n1857 );
  or       g01482 ( new_n1859 , new_n1854 , new_n1858 );
  nor      g01483 ( new_n1860 , new_n1829 , new_n1859 );
  xnor     g01484 ( new_n1861 , new_n1829 , new_n1859 );
  nor      g01485 ( new_n1862 , new_n1839 , new_n1840 );
  and      g01486 ( new_n1863 , new_n1841 , new_n1842 );
  nor      g01487 ( new_n1864 , new_n1862 , new_n1863 );
  xor      g01488 ( new_n1865 , new_n1807 , new_n1811 );
  xor      g01489 ( new_n1866 , new_n1864 , new_n1865 );
  xnor     g01490 ( new_n1867 , new_n1538 , new_n1539 );
  xor      g01491 ( new_n1868 , new_n1866 , new_n1867 );
  nor      g01492 ( new_n1869 , new_n1861 , new_n1868 );
  or       g01493 ( new_n1870 , new_n1860 , new_n1869 );
  xor      g01494 ( new_n1871 , new_n1661 , new_n1668 );
  nor      g01495 ( new_n1872 , new_n1870 , new_n1871 );
  nor      g01496 ( new_n1873 , new_n1864 , new_n1865 );
  nand g01497 ( new_n1874 , new_n1873 , new_n1873 );
  nand     g01498 ( new_n1875 , new_n1866 , new_n1867 );
  nand     g01499 ( new_n1876 , new_n1874 , new_n1875 );
  xnor     g01500 ( new_n1877 , new_n1543 , new_n1544 );
  xor      g01501 ( new_n1878 , new_n1806 , new_n1813 );
  xnor     g01502 ( new_n1879 , new_n1877 , new_n1878 );
  xor      g01503 ( new_n1880 , new_n1876 , new_n1879 );
  xnor     g01504 ( new_n1881 , new_n1870 , new_n1871 );
  nor      g01505 ( new_n1882 , new_n1880 , new_n1881 );
  or       g01506 ( new_n1883 , new_n1872 , new_n1882 );
  xnor     g01507 ( new_n1884 , new_n1672 , new_n1673 );
  nor      g01508 ( new_n1885 , new_n1883 , new_n1884 );
  xnor     g01509 ( new_n1886 , new_n1883 , new_n1884 );
  nor      g01510 ( new_n1887 , new_n1877 , new_n1878 );
  nor      g01511 ( new_n1888 , new_n1876 , new_n1879 );
  or       g01512 ( new_n1889 , new_n1887 , new_n1888 );
  xor      g01513 ( new_n1890 , new_n1549 , new_n1550 );
  xor      g01514 ( new_n1891 , new_n1816 , new_n1817 );
  xnor     g01515 ( new_n1892 , new_n1890 , new_n1891 );
  xor      g01516 ( new_n1893 , new_n1889 , new_n1892 );
  nor      g01517 ( new_n1894 , new_n1886 , new_n1893 );
  nor      g01518 ( new_n1895 , new_n1885 , new_n1894 );
  xor      g01519 ( new_n1896 , new_n1659 , new_n1675 );
  nand     g01520 ( new_n1897 , new_n1895 , new_n1896 );
  xor      g01521 ( new_n1898 , new_n1895 , new_n1896 );
  nor      g01522 ( new_n1899 , new_n1890 , new_n1891 );
  nor      g01523 ( new_n1900 , new_n1889 , new_n1892 );
  or       g01524 ( new_n1901 , new_n1899 , new_n1900 );
  xor      g01525 ( new_n1902 , new_n1819 , new_n1820 );
  xnor     g01526 ( new_n1903 , new_n1901 , new_n1902 );
  xor      g01527 ( new_n1904 , new_n1561 , new_n1562 );
  xnor     g01528 ( new_n1905 , new_n1903 , new_n1904 );
  nand     g01529 ( new_n1906 , new_n1898 , new_n1905 );
  nand     g01530 ( new_n1907 , new_n1897 , new_n1906 );
  nor      g01531 ( new_n1908 , new_n1901 , new_n1902 );
  nor      g01532 ( new_n1909 , new_n1903 , new_n1904 );
  nor      g01533 ( new_n1910 , new_n1908 , new_n1909 );
  nand     g01534 ( new_n1911 , pi045 , pi177 );
  nor      g01535 ( new_n1912 , new_n1388 , new_n1420 );
  nand g01536 ( new_n1913 , new_n1421 , new_n1421 );
  nor      g01537 ( new_n1914 , new_n1417 , new_n1913 );
  nor      g01538 ( new_n1915 , new_n1912 , new_n1914 );
  xor      g01539 ( new_n1916 , new_n1911 , new_n1915 );
  nand     g01540 ( new_n1917 , pi031 , pi142 );
  xor      g01541 ( new_n1918 , new_n1916 , new_n1917 );
  nand     g01542 ( new_n1919 , pi044 , pi101 );
  nand     g01543 ( new_n1920 , pi155 , pi206 );
  nand     g01544 ( new_n1921 , pi060 , pi072 );
  xor      g01545 ( new_n1922 , new_n1920 , new_n1921 );
  xor      g01546 ( new_n1923 , new_n1919 , new_n1922 );
  nand     g01547 ( new_n1924 , pi019 , pi079 );
  nand     g01548 ( new_n1925 , new_n1715 , new_n1716 );
  nand     g01549 ( new_n1926 , new_n1710 , new_n1717 );
  nand     g01550 ( new_n1927 , new_n1925 , new_n1926 );
  xor      g01551 ( new_n1928 , new_n1924 , new_n1927 );
  xor      g01552 ( new_n1929 , new_n1923 , new_n1928 );
  xor      g01553 ( new_n1930 , new_n1918 , new_n1929 );
  xor      g01554 ( new_n1931 , new_n1910 , new_n1930 );
  nand     g01555 ( new_n1932 , pi076 , pi097 );
  or       g01556 ( new_n1933 , new_n1795 , new_n1802 );
  nand     g01557 ( new_n1934 , new_n1793 , new_n1933 );
  nand     g01558 ( new_n1935 , pi023 , pi032 );
  nand g01559 ( new_n1936 , new_n1799 , new_n1799 );
  nor      g01560 ( new_n1937 , new_n1936 , new_n1800 );
  nor      g01561 ( new_n1938 , new_n1796 , new_n1801 );
  nor      g01562 ( new_n1939 , new_n1937 , new_n1938 );
  xnor     g01563 ( new_n1940 , new_n1935 , new_n1939 );
  xor      g01564 ( new_n1941 , new_n1934 , new_n1940 );
  xor      g01565 ( new_n1942 , new_n1932 , new_n1941 );
  xor      g01566 ( new_n1943 , new_n1931 , new_n1942 );
  xor      g01567 ( new_n1944 , new_n1907 , new_n1943 );
  xor      g01568 ( new_n1945 , new_n1828 , new_n1944 );
  xor      g01569 ( po005 , new_n1572 , new_n1945 );
  nand     g01570 ( new_n1947 , pi070 , pi073 );
  nand     g01571 ( new_n1948 , pi030 , pi117 );
  xor      g01572 ( new_n1949 , new_n1947 , new_n1948 );
  nand     g01573 ( new_n1950 , pi000 , pi170 );
  nand     g01574 ( new_n1951 , pi065 , pi203 );
  nand     g01575 ( new_n1952 , pi022 , pi163 );
  xor      g01576 ( new_n1953 , new_n1951 , new_n1952 );
  xor      g01577 ( new_n1954 , new_n1950 , new_n1953 );
  xor      g01578 ( new_n1955 , new_n1949 , new_n1954 );
  nand     g01579 ( new_n1956 , pi065 , pi167 );
  nand     g01580 ( new_n1957 , pi120 , pi240 );
  nand     g01581 ( new_n1958 , pi062 , pi149 );
  xor      g01582 ( new_n1959 , new_n1957 , new_n1958 );
  xor      g01583 ( new_n1960 , new_n1956 , new_n1959 );
  nand     g01584 ( new_n1961 , pi062 , pi240 );
  nand     g01585 ( new_n1962 , pi065 , pi149 );
  nand     g01586 ( new_n1963 , new_n1961 , new_n1962 );
  nand     g01587 ( new_n1964 , pi120 , pi134 );
  xor      g01588 ( new_n1965 , new_n1961 , new_n1962 );
  nand     g01589 ( new_n1966 , new_n1964 , new_n1965 );
  nand     g01590 ( new_n1967 , new_n1963 , new_n1966 );
  nand     g01591 ( new_n1968 , pi134 , pi172 );
  xor      g01592 ( new_n1969 , new_n1967 , new_n1968 );
  xor      g01593 ( new_n1970 , new_n1960 , new_n1969 );
  nand     g01594 ( new_n1971 , pi175 , pi198 );
  nor      g01595 ( new_n1972 , new_n1970 , new_n1971 );
  xor      g01596 ( new_n1973 , new_n1970 , new_n1971 );
  nand g01597 ( new_n1974 , new_n1973 , new_n1973 );
  nand     g01598 ( new_n1975 , pi062 , pi134 );
  nand g01599 ( new_n1976 , new_n1975 , new_n1975 );
  nand     g01600 ( new_n1977 , pi065 , pi240 );
  nand     g01601 ( new_n1978 , pi120 , pi175 );
  nor      g01602 ( new_n1979 , new_n1977 , new_n1978 );
  or       g01603 ( new_n1980 , new_n1976 , new_n1979 );
  nand     g01604 ( new_n1981 , new_n1977 , new_n1978 );
  nand     g01605 ( new_n1982 , new_n1980 , new_n1981 );
  nand     g01606 ( new_n1983 , pi172 , pi175 );
  nor      g01607 ( new_n1984 , new_n1982 , new_n1983 );
  xor      g01608 ( new_n1985 , new_n1964 , new_n1965 );
  xor      g01609 ( new_n1986 , new_n1982 , new_n1983 );
  nand g01610 ( new_n1987 , new_n1986 , new_n1986 );
  nor      g01611 ( new_n1988 , new_n1985 , new_n1987 );
  nor      g01612 ( new_n1989 , new_n1984 , new_n1988 );
  nor      g01613 ( new_n1990 , new_n1974 , new_n1989 );
  nor      g01614 ( new_n1991 , new_n1972 , new_n1990 );
  nand     g01615 ( new_n1992 , pi172 , pi240 );
  nand     g01616 ( new_n1993 , pi134 , pi198 );
  nand     g01617 ( new_n1994 , new_n1992 , new_n1993 );
  nand     g01618 ( new_n1995 , pi198 , pi240 );
  nor      g01619 ( new_n1996 , new_n1968 , new_n1995 );
  nand g01620 ( new_n1997 , new_n1996 , new_n1996 );
  nand     g01621 ( new_n1998 , new_n1994 , new_n1997 );
  nand     g01622 ( new_n1999 , new_n1957 , new_n1958 );
  nand     g01623 ( new_n2000 , new_n1956 , new_n1959 );
  nand     g01624 ( new_n2001 , new_n1999 , new_n2000 );
  nand     g01625 ( new_n2002 , pi120 , pi149 );
  nand     g01626 ( new_n2003 , pi062 , pi167 );
  nand     g01627 ( new_n2004 , pi065 , pi181 );
  nand     g01628 ( new_n2005 , new_n2003 , new_n2004 );
  nand     g01629 ( new_n2006 , pi062 , pi181 );
  or       g01630 ( new_n2007 , new_n2006 , new_n1956 );
  nand     g01631 ( new_n2008 , new_n2005 , new_n2007 );
  xor      g01632 ( new_n2009 , new_n2002 , new_n2008 );
  xor      g01633 ( new_n2010 , new_n2001 , new_n2009 );
  xor      g01634 ( new_n2011 , new_n1998 , new_n2010 );
  nand     g01635 ( new_n2012 , new_n1967 , new_n1968 );
  nand     g01636 ( new_n2013 , new_n1960 , new_n1969 );
  nand     g01637 ( new_n2014 , new_n2012 , new_n2013 );
  xor      g01638 ( new_n2015 , new_n2011 , new_n2014 );
  nor      g01639 ( new_n2016 , new_n1991 , new_n2015 );
  nand     g01640 ( new_n2017 , pi134 , pi165 );
  nand     g01641 ( new_n2018 , pi175 , pi197 );
  xor      g01642 ( new_n2019 , new_n2017 , new_n2018 );
  xor      g01643 ( new_n2020 , new_n1995 , new_n2019 );
  nand     g01644 ( new_n2021 , new_n2002 , new_n2008 );
  nand     g01645 ( new_n2022 , new_n2001 , new_n2009 );
  nand     g01646 ( new_n2023 , new_n2021 , new_n2022 );
  xor      g01647 ( new_n2024 , new_n2020 , new_n2023 );
  nand     g01648 ( new_n2025 , pi149 , pi172 );
  xor      g01649 ( new_n2026 , new_n2007 , new_n2025 );
  nand     g01650 ( new_n2027 , pi065 , pi200 );
  and      g01651 ( new_n2028 , pi120 , pi167 );
  xor      g01652 ( new_n2029 , new_n2027 , new_n2028 );
  xor      g01653 ( new_n2030 , new_n2006 , new_n2029 );
  xnor     g01654 ( new_n2031 , new_n2026 , new_n2030 );
  xor      g01655 ( new_n2032 , new_n2024 , new_n2031 );
  nand     g01656 ( new_n2033 , new_n1998 , new_n2010 );
  nand     g01657 ( new_n2034 , new_n2011 , new_n2014 );
  nand     g01658 ( new_n2035 , new_n2033 , new_n2034 );
  xor      g01659 ( new_n2036 , new_n1996 , new_n2035 );
  xor      g01660 ( new_n2037 , new_n2032 , new_n2036 );
  or       g01661 ( new_n2038 , new_n2016 , new_n2037 );
  xor      g01662 ( new_n2039 , new_n2016 , new_n2037 );
  nand     g01663 ( new_n2040 , pi165 , pi175 );
  xor      g01664 ( new_n2041 , new_n1985 , new_n1987 );
  nand     g01665 ( new_n2042 , pi065 , pi175 );
  nand g01666 ( new_n2043 , new_n2042 , new_n2042 );
  nor      g01667 ( new_n2044 , new_n1975 , new_n2043 );
  nor      g01668 ( new_n2045 , new_n1981 , new_n2044 );
  nor      g01669 ( new_n2046 , new_n1979 , new_n2045 );
  nor      g01670 ( new_n2047 , new_n1975 , new_n2046 );
  nand     g01671 ( new_n2048 , new_n2041 , new_n2047 );
  xor      g01672 ( new_n2049 , new_n1973 , new_n1989 );
  nor      g01673 ( new_n2050 , new_n2048 , new_n2049 );
  nand g01674 ( new_n2051 , new_n2050 , new_n2050 );
  nand     g01675 ( new_n2052 , new_n2040 , new_n2051 );
  nand g01676 ( new_n2053 , new_n2052 , new_n2052 );
  xor      g01677 ( new_n2054 , new_n1991 , new_n2015 );
  xor      g01678 ( new_n2055 , new_n2040 , new_n2050 );
  nor      g01679 ( new_n2056 , new_n2054 , new_n2055 );
  nor      g01680 ( new_n2057 , new_n2053 , new_n2056 );
  nand g01681 ( new_n2058 , new_n2057 , new_n2057 );
  nand     g01682 ( new_n2059 , new_n2039 , new_n2058 );
  nand     g01683 ( new_n2060 , new_n2038 , new_n2059 );
  nand     g01684 ( new_n2061 , pi190 , pi214 );
  nand     g01685 ( new_n2062 , pi229 , pi247 );
  nand     g01686 ( new_n2063 , new_n2061 , new_n2062 );
  nand     g01687 ( new_n2064 , pi092 , pi234 );
  xor      g01688 ( new_n2065 , new_n2061 , new_n2062 );
  nand     g01689 ( new_n2066 , new_n2064 , new_n2065 );
  nand     g01690 ( new_n2067 , new_n2063 , new_n2066 );
  xor      g01691 ( new_n2068 , new_n2060 , new_n2067 );
  nand g01692 ( new_n2069 , pi004 , pi004 );
  nor      g01693 ( new_n2070 , new_n2069 , new_n949 );
  nand g01694 ( new_n2071 , new_n2070 , new_n2070 );
  nand     g01695 ( new_n2072 , pi073 , pi163 );
  nand     g01696 ( new_n2073 , pi170 , pi228 );
  nor      g01697 ( new_n2074 , new_n2072 , new_n2073 );
  nand     g01698 ( new_n2075 , pi163 , pi170 );
  and      g01699 ( new_n2076 , new_n2070 , new_n2075 );
  nand     g01700 ( new_n2077 , new_n2072 , new_n2073 );
  nor      g01701 ( new_n2078 , new_n2076 , new_n2077 );
  nor      g01702 ( new_n2079 , new_n2074 , new_n2078 );
  nor      g01703 ( new_n2080 , new_n2071 , new_n2079 );
  nand     g01704 ( new_n2081 , pi039 , pi170 );
  nand     g01705 ( new_n2082 , pi004 , pi228 );
  nand     g01706 ( new_n2083 , pi073 , pi148 );
  xor      g01707 ( new_n2084 , new_n2082 , new_n2083 );
  xor      g01708 ( new_n2085 , new_n2081 , new_n2084 );
  or       g01709 ( new_n2086 , new_n2070 , new_n2074 );
  nand     g01710 ( new_n2087 , new_n2077 , new_n2086 );
  nand     g01711 ( new_n2088 , pi003 , pi163 );
  xor      g01712 ( new_n2089 , new_n2087 , new_n2088 );
  xnor     g01713 ( new_n2090 , new_n2085 , new_n2089 );
  nand     g01714 ( new_n2091 , new_n2080 , new_n2090 );
  nand     g01715 ( new_n2092 , pi130 , pi163 );
  nand     g01716 ( new_n2093 , new_n2087 , new_n2088 );
  nand     g01717 ( new_n2094 , new_n2085 , new_n2089 );
  nand     g01718 ( new_n2095 , new_n2093 , new_n2094 );
  xnor     g01719 ( new_n2096 , new_n2092 , new_n2095 );
  nand     g01720 ( new_n2097 , pi004 , pi039 );
  nand     g01721 ( new_n2098 , pi073 , pi228 );
  nand     g01722 ( new_n2099 , pi116 , pi170 );
  xor      g01723 ( new_n2100 , new_n2098 , new_n2099 );
  xor      g01724 ( new_n2101 , new_n2097 , new_n2100 );
  nand     g01725 ( new_n2102 , pi003 , pi148 );
  nand     g01726 ( new_n2103 , new_n2082 , new_n2083 );
  nand     g01727 ( new_n2104 , new_n2081 , new_n2084 );
  nand     g01728 ( new_n2105 , new_n2103 , new_n2104 );
  xor      g01729 ( new_n2106 , new_n2102 , new_n2105 );
  xor      g01730 ( new_n2107 , new_n2101 , new_n2106 );
  xnor     g01731 ( new_n2108 , new_n2096 , new_n2107 );
  nor      g01732 ( new_n2109 , new_n2091 , new_n2108 );
  nand g01733 ( new_n2110 , new_n2109 , new_n2109 );
  nor      g01734 ( new_n2111 , new_n2092 , new_n2095 );
  nor      g01735 ( new_n2112 , new_n2096 , new_n2107 );
  nor      g01736 ( new_n2113 , new_n2111 , new_n2112 );
  nand     g01737 ( new_n2114 , pi130 , pi148 );
  nand     g01738 ( new_n2115 , pi003 , pi228 );
  and      g01739 ( new_n2116 , new_n2114 , new_n2115 );
  nand     g01740 ( new_n2117 , pi130 , pi228 );
  nor      g01741 ( new_n2118 , new_n2117 , new_n2102 );
  or       g01742 ( new_n2119 , new_n2116 , new_n2118 );
  nand     g01743 ( new_n2120 , pi070 , pi170 );
  nand     g01744 ( new_n2121 , pi004 , pi116 );
  nand     g01745 ( new_n2122 , new_n2120 , new_n2121 );
  nand     g01746 ( new_n2123 , pi004 , pi070 );
  nor      g01747 ( new_n2124 , new_n2099 , new_n2123 );
  nand g01748 ( new_n2125 , new_n2124 , new_n2124 );
  nand     g01749 ( new_n2126 , new_n2122 , new_n2125 );
  nand     g01750 ( new_n2127 , pi039 , pi073 );
  nand     g01751 ( new_n2128 , new_n2098 , new_n2099 );
  nand     g01752 ( new_n2129 , new_n2097 , new_n2100 );
  nand     g01753 ( new_n2130 , new_n2128 , new_n2129 );
  xor      g01754 ( new_n2131 , new_n2127 , new_n2130 );
  xor      g01755 ( new_n2132 , new_n2126 , new_n2131 );
  xor      g01756 ( new_n2133 , new_n2119 , new_n2132 );
  nand     g01757 ( new_n2134 , new_n2102 , new_n2105 );
  nand     g01758 ( new_n2135 , new_n2101 , new_n2106 );
  nand     g01759 ( new_n2136 , new_n2134 , new_n2135 );
  xor      g01760 ( new_n2137 , new_n2133 , new_n2136 );
  xor      g01761 ( new_n2138 , new_n2113 , new_n2137 );
  nand     g01762 ( new_n2139 , pi124 , pi163 );
  xor      g01763 ( new_n2140 , new_n2138 , new_n2139 );
  xor      g01764 ( new_n2141 , new_n2110 , new_n2140 );
  nand     g01765 ( new_n2142 , pi095 , pi107 );
  nand     g01766 ( new_n2143 , pi158 , pi171 );
  nand     g01767 ( new_n2144 , pi049 , pi254 );
  nand     g01768 ( new_n2145 , pi089 , pi107 );
  or       g01769 ( new_n2146 , new_n2144 , new_n2145 );
  nand     g01770 ( new_n2147 , new_n2143 , new_n2146 );
  nand     g01771 ( new_n2148 , new_n2144 , new_n2145 );
  nand     g01772 ( new_n2149 , new_n2147 , new_n2148 );
  nand     g01773 ( new_n2150 , pi107 , pi154 );
  nor      g01774 ( new_n2151 , new_n2149 , new_n2150 );
  xor      g01775 ( new_n2152 , new_n2149 , new_n2150 );
  nand     g01776 ( new_n2153 , pi049 , pi158 );
  nand     g01777 ( new_n2154 , pi245 , pi254 );
  nand g01778 ( new_n2155 , pi089 , pi089 );
  nand g01779 ( new_n2156 , pi171 , pi171 );
  nor      g01780 ( new_n2157 , new_n2155 , new_n2156 );
  xor      g01781 ( new_n2158 , new_n2154 , new_n2157 );
  xor      g01782 ( new_n2159 , new_n2153 , new_n2158 );
  and      g01783 ( new_n2160 , new_n2152 , new_n2159 );
  nor      g01784 ( new_n2161 , new_n2151 , new_n2160 );
  nor      g01785 ( new_n2162 , new_n2142 , new_n2161 );
  xor      g01786 ( new_n2163 , new_n2142 , new_n2161 );
  nand     g01787 ( new_n2164 , pi049 , pi089 );
  nand     g01788 ( new_n2165 , pi201 , pi254 );
  nand g01789 ( new_n2166 , new_n2165 , new_n2165 );
  nand     g01790 ( new_n2167 , pi158 , pi245 );
  xor      g01791 ( new_n2168 , new_n2166 , new_n2167 );
  xor      g01792 ( new_n2169 , new_n2164 , new_n2168 );
  nand g01793 ( new_n2170 , new_n2154 , new_n2154 );
  nor      g01794 ( new_n2171 , new_n2170 , new_n2157 );
  nand g01795 ( new_n2172 , new_n2153 , new_n2153 );
  nor      g01796 ( new_n2173 , new_n2172 , new_n2158 );
  nor      g01797 ( new_n2174 , new_n2171 , new_n2173 );
  nand     g01798 ( new_n2175 , pi154 , pi171 );
  xor      g01799 ( new_n2176 , new_n2174 , new_n2175 );
  xnor     g01800 ( new_n2177 , new_n2169 , new_n2176 );
  and      g01801 ( new_n2178 , new_n2163 , new_n2177 );
  nor      g01802 ( new_n2179 , new_n2162 , new_n2178 );
  nand g01803 ( new_n2180 , new_n2175 , new_n2175 );
  nor      g01804 ( new_n2181 , new_n2174 , new_n2180 );
  nor      g01805 ( new_n2182 , new_n2169 , new_n2176 );
  nor      g01806 ( new_n2183 , new_n2181 , new_n2182 );
  nand     g01807 ( new_n2184 , pi049 , pi154 );
  nand     g01808 ( new_n2185 , pi095 , pi171 );
  and      g01809 ( new_n2186 , new_n2184 , new_n2185 );
  nand     g01810 ( new_n2187 , pi049 , pi095 );
  nor      g01811 ( new_n2188 , new_n2187 , new_n2175 );
  nor      g01812 ( new_n2189 , new_n2186 , new_n2188 );
  nand     g01813 ( new_n2190 , new_n2165 , new_n2167 );
  nand g01814 ( new_n2191 , new_n2168 , new_n2168 );
  nand     g01815 ( new_n2192 , new_n2164 , new_n2191 );
  nand     g01816 ( new_n2193 , new_n2190 , new_n2192 );
  nand     g01817 ( new_n2194 , pi089 , pi245 );
  nand     g01818 ( new_n2195 , pi156 , pi158 );
  nand g01819 ( new_n2196 , new_n2195 , new_n2195 );
  nand     g01820 ( new_n2197 , new_n2196 , new_n2166 );
  nand     g01821 ( new_n2198 , pi158 , pi201 );
  nand     g01822 ( new_n2199 , pi156 , pi254 );
  nand     g01823 ( new_n2200 , new_n2198 , new_n2199 );
  nand     g01824 ( new_n2201 , new_n2197 , new_n2200 );
  xor      g01825 ( new_n2202 , new_n2194 , new_n2201 );
  xnor     g01826 ( new_n2203 , new_n2193 , new_n2202 );
  xnor     g01827 ( new_n2204 , new_n2189 , new_n2203 );
  xor      g01828 ( new_n2205 , new_n2183 , new_n2204 );
  xnor     g01829 ( new_n2206 , new_n2179 , new_n2205 );
  nand     g01830 ( new_n2207 , pi006 , pi107 );
  xor      g01831 ( new_n2208 , new_n2163 , new_n2177 );
  xor      g01832 ( new_n2209 , new_n2152 , new_n2159 );
  nand     g01833 ( new_n2210 , pi107 , pi254 );
  nand g01834 ( new_n2211 , new_n2210 , new_n2210 );
  nor      g01835 ( new_n2212 , new_n2143 , new_n2211 );
  and      g01836 ( new_n2213 , new_n2146 , new_n2148 );
  or       g01837 ( new_n2214 , new_n2212 , new_n2213 );
  nor      g01838 ( new_n2215 , new_n2143 , new_n2214 );
  and      g01839 ( new_n2216 , new_n2209 , new_n2215 );
  nand     g01840 ( new_n2217 , new_n2208 , new_n2216 );
  xor      g01841 ( new_n2218 , new_n2207 , new_n2217 );
  xnor     g01842 ( new_n2219 , new_n2206 , new_n2218 );
  nand     g01843 ( new_n2220 , new_n2141 , new_n2219 );
  xor      g01844 ( new_n2221 , new_n2141 , new_n2219 );
  xor      g01845 ( new_n2222 , new_n2208 , new_n2216 );
  xor      g01846 ( new_n2223 , new_n2209 , new_n2215 );
  nand     g01847 ( new_n2224 , new_n2148 , new_n2212 );
  nand     g01848 ( new_n2225 , new_n2214 , new_n2224 );
  nand     g01849 ( new_n2226 , new_n2076 , new_n2077 );
  nand     g01850 ( new_n2227 , new_n2079 , new_n2226 );
  nor      g01851 ( new_n2228 , new_n2225 , new_n2227 );
  and      g01852 ( new_n2229 , new_n2225 , new_n2227 );
  nand     g01853 ( new_n2230 , pi171 , pi254 );
  nand     g01854 ( new_n2231 , pi107 , pi158 );
  xor      g01855 ( new_n2232 , new_n2230 , new_n2231 );
  nor      g01856 ( new_n2233 , new_n2075 , new_n2210 );
  nand     g01857 ( new_n2234 , new_n2232 , new_n2233 );
  xor      g01858 ( new_n2235 , new_n2232 , new_n2233 );
  nand     g01859 ( new_n2236 , pi004 , pi163 );
  nand     g01860 ( new_n2237 , pi148 , pi170 );
  xor      g01861 ( new_n2238 , new_n2236 , new_n2237 );
  nand     g01862 ( new_n2239 , new_n2235 , new_n2238 );
  and      g01863 ( new_n2240 , new_n2234 , new_n2239 );
  nor      g01864 ( new_n2241 , new_n2229 , new_n2240 );
  or       g01865 ( new_n2242 , new_n2228 , new_n2241 );
  nor      g01866 ( new_n2243 , new_n2223 , new_n2242 );
  xor      g01867 ( new_n2244 , new_n2080 , new_n2090 );
  nor      g01868 ( new_n2245 , new_n2228 , new_n2241 );
  xor      g01869 ( new_n2246 , new_n2223 , new_n2245 );
  nor      g01870 ( new_n2247 , new_n2244 , new_n2246 );
  nor      g01871 ( new_n2248 , new_n2243 , new_n2247 );
  nor      g01872 ( new_n2249 , new_n2222 , new_n2248 );
  nand g01873 ( new_n2250 , new_n2222 , new_n2222 );
  xor      g01874 ( new_n2251 , new_n2250 , new_n2248 );
  xor      g01875 ( new_n2252 , new_n2091 , new_n2108 );
  nor      g01876 ( new_n2253 , new_n2251 , new_n2252 );
  nor      g01877 ( new_n2254 , new_n2249 , new_n2253 );
  nand     g01878 ( new_n2255 , new_n2221 , new_n2254 );
  and      g01879 ( new_n2256 , new_n2220 , new_n2255 );
  nand     g01880 ( new_n2257 , new_n2207 , new_n2217 );
  nand     g01881 ( new_n2258 , new_n2206 , new_n2218 );
  nand     g01882 ( new_n2259 , new_n2257 , new_n2258 );
  or       g01883 ( new_n2260 , new_n2179 , new_n2205 );
  nand     g01884 ( new_n2261 , pi006 , pi171 );
  nand     g01885 ( new_n2262 , pi107 , pi209 );
  xor      g01886 ( new_n2263 , new_n2261 , new_n2262 );
  xnor     g01887 ( new_n2264 , new_n2187 , new_n2263 );
  nand     g01888 ( new_n2265 , new_n2194 , new_n2201 );
  nand     g01889 ( new_n2266 , new_n2193 , new_n2202 );
  nand     g01890 ( new_n2267 , new_n2265 , new_n2266 );
  nand g01891 ( new_n2268 , new_n2267 , new_n2267 );
  xor      g01892 ( new_n2269 , new_n2264 , new_n2268 );
  nand     g01893 ( new_n2270 , pi089 , pi201 );
  and      g01894 ( new_n2271 , pi063 , pi254 );
  xor      g01895 ( new_n2272 , new_n2270 , new_n2271 );
  xor      g01896 ( new_n2273 , new_n2196 , new_n2272 );
  nand     g01897 ( new_n2274 , pi154 , pi245 );
  xnor     g01898 ( new_n2275 , new_n2197 , new_n2274 );
  xor      g01899 ( new_n2276 , new_n2273 , new_n2275 );
  nand g01900 ( new_n2277 , new_n2276 , new_n2276 );
  xor      g01901 ( new_n2278 , new_n2269 , new_n2277 );
  nor      g01902 ( new_n2279 , new_n2189 , new_n2203 );
  nor      g01903 ( new_n2280 , new_n2183 , new_n2204 );
  nor      g01904 ( new_n2281 , new_n2279 , new_n2280 );
  xor      g01905 ( new_n2282 , new_n2188 , new_n2281 );
  xor      g01906 ( new_n2283 , new_n2278 , new_n2282 );
  xor      g01907 ( new_n2284 , new_n2260 , new_n2283 );
  xnor     g01908 ( new_n2285 , new_n2259 , new_n2284 );
  nand g01909 ( new_n2286 , new_n2139 , new_n2139 );
  nand     g01910 ( new_n2287 , new_n2138 , new_n2286 );
  or       g01911 ( new_n2288 , new_n2110 , new_n2140 );
  nand     g01912 ( new_n2289 , new_n2287 , new_n2288 );
  nor      g01913 ( new_n2290 , new_n2113 , new_n2137 );
  nand g01914 ( new_n2291 , new_n2133 , new_n2133 );
  nor      g01915 ( new_n2292 , new_n2291 , new_n2136 );
  nand     g01916 ( new_n2293 , new_n2118 , new_n2292 );
  nor      g01917 ( new_n2294 , new_n2119 , new_n2132 );
  nor      g01918 ( new_n2295 , new_n2118 , new_n2294 );
  nand g01919 ( new_n2296 , new_n2295 , new_n2295 );
  or       g01920 ( new_n2297 , new_n2292 , new_n2296 );
  nand     g01921 ( new_n2298 , new_n2293 , new_n2297 );
  nand     g01922 ( new_n2299 , pi003 , pi039 );
  xor      g01923 ( new_n2300 , new_n2124 , new_n2299 );
  nand     g01924 ( new_n2301 , pi073 , pi116 );
  nand     g01925 ( new_n2302 , pi115 , pi170 );
  xor      g01926 ( new_n2303 , new_n2301 , new_n2302 );
  xor      g01927 ( new_n2304 , new_n2123 , new_n2303 );
  xor      g01928 ( new_n2305 , new_n2300 , new_n2304 );
  nand     g01929 ( new_n2306 , new_n2127 , new_n2130 );
  nand     g01930 ( new_n2307 , new_n2126 , new_n2131 );
  nand     g01931 ( new_n2308 , new_n2306 , new_n2307 );
  nand     g01932 ( new_n2309 , pi124 , pi148 );
  nand     g01933 ( new_n2310 , pi163 , pi215 );
  xor      g01934 ( new_n2311 , new_n2117 , new_n2310 );
  xor      g01935 ( new_n2312 , new_n2309 , new_n2311 );
  xor      g01936 ( new_n2313 , new_n2308 , new_n2312 );
  xor      g01937 ( new_n2314 , new_n2305 , new_n2313 );
  xor      g01938 ( new_n2315 , new_n2298 , new_n2314 );
  xor      g01939 ( new_n2316 , new_n2290 , new_n2315 );
  xor      g01940 ( new_n2317 , new_n2289 , new_n2316 );
  xor      g01941 ( new_n2318 , new_n2285 , new_n2317 );
  xor      g01942 ( new_n2319 , new_n2256 , new_n2318 );
  xor      g01943 ( new_n2320 , new_n2251 , new_n2252 );
  xnor     g01944 ( new_n2321 , new_n2048 , new_n2049 );
  or       g01945 ( new_n2322 , new_n2320 , new_n2321 );
  xor      g01946 ( new_n2323 , new_n2041 , new_n2047 );
  nand g01947 ( new_n2324 , new_n2323 , new_n2323 );
  xor      g01948 ( new_n2325 , new_n2244 , new_n2246 );
  nand     g01949 ( new_n2326 , new_n2324 , new_n2325 );
  xor      g01950 ( new_n2327 , new_n2324 , new_n2325 );
  nor      g01951 ( new_n2328 , new_n2228 , new_n2229 );
  xor      g01952 ( new_n2329 , new_n2240 , new_n2328 );
  nand     g01953 ( new_n2330 , new_n1981 , new_n2044 );
  nand     g01954 ( new_n2331 , new_n2046 , new_n2330 );
  nor      g01955 ( new_n2332 , new_n2329 , new_n2331 );
  xor      g01956 ( new_n2333 , new_n2075 , new_n2210 );
  nand     g01957 ( new_n2334 , new_n2043 , new_n2333 );
  nand g01958 ( new_n2335 , new_n2334 , new_n2334 );
  nand     g01959 ( new_n2336 , pi062 , pi175 );
  nand     g01960 ( new_n2337 , pi065 , pi134 );
  xor      g01961 ( new_n2338 , new_n2336 , new_n2337 );
  nor      g01962 ( new_n2339 , new_n2335 , new_n2338 );
  xor      g01963 ( new_n2340 , new_n2235 , new_n2238 );
  xor      g01964 ( new_n2341 , new_n2334 , new_n2338 );
  nor      g01965 ( new_n2342 , new_n2340 , new_n2341 );
  nor      g01966 ( new_n2343 , new_n2339 , new_n2342 );
  nand g01967 ( new_n2344 , new_n2343 , new_n2343 );
  xnor     g01968 ( new_n2345 , new_n2329 , new_n2331 );
  nor      g01969 ( new_n2346 , new_n2344 , new_n2345 );
  nor      g01970 ( new_n2347 , new_n2332 , new_n2346 );
  nand     g01971 ( new_n2348 , new_n2327 , new_n2347 );
  and      g01972 ( new_n2349 , new_n2326 , new_n2348 );
  xor      g01973 ( new_n2350 , new_n2320 , new_n2321 );
  nand     g01974 ( new_n2351 , new_n2349 , new_n2350 );
  nand     g01975 ( new_n2352 , new_n2322 , new_n2351 );
  xnor     g01976 ( new_n2353 , new_n2054 , new_n2055 );
  nor      g01977 ( new_n2354 , new_n2352 , new_n2353 );
  xnor     g01978 ( new_n2355 , new_n2352 , new_n2353 );
  xor      g01979 ( new_n2356 , new_n2221 , new_n2254 );
  nor      g01980 ( new_n2357 , new_n2355 , new_n2356 );
  nor      g01981 ( new_n2358 , new_n2354 , new_n2357 );
  nor      g01982 ( new_n2359 , new_n2319 , new_n2358 );
  xnor     g01983 ( new_n2360 , new_n2319 , new_n2358 );
  xor      g01984 ( new_n2361 , new_n2039 , new_n2057 );
  nor      g01985 ( new_n2362 , new_n2360 , new_n2361 );
  nor      g01986 ( new_n2363 , new_n2359 , new_n2362 );
  nand     g01987 ( new_n2364 , pi067 , pi247 );
  nand     g01988 ( new_n2365 , pi092 , pi214 );
  xor      g01989 ( new_n2366 , new_n2364 , new_n2365 );
  xor      g01990 ( new_n2367 , new_n2363 , new_n2366 );
  xor      g01991 ( new_n2368 , new_n2068 , new_n2367 );
  nand     g01992 ( new_n2369 , pi006 , pi049 );
  nand     g01993 ( new_n2370 , pi067 , pi117 );
  nand     g01994 ( new_n2371 , pi080 , pi190 );
  nand     g01995 ( new_n2372 , pi016 , pi092 );
  nand     g01996 ( new_n2373 , new_n2371 , new_n2372 );
  nand     g01997 ( new_n2374 , pi117 , pi229 );
  xor      g01998 ( new_n2375 , new_n2371 , new_n2372 );
  nand     g01999 ( new_n2376 , new_n2374 , new_n2375 );
  nand     g02000 ( new_n2377 , new_n2373 , new_n2376 );
  nand     g02001 ( new_n2378 , new_n2370 , new_n2377 );
  nand     g02002 ( new_n2379 , pi190 , pi247 );
  nand     g02003 ( new_n2380 , pi080 , pi092 );
  nand     g02004 ( new_n2381 , pi016 , pi229 );
  xor      g02005 ( new_n2382 , new_n2380 , new_n2381 );
  xor      g02006 ( new_n2383 , new_n2379 , new_n2382 );
  xor      g02007 ( new_n2384 , new_n2370 , new_n2377 );
  nand     g02008 ( new_n2385 , new_n2383 , new_n2384 );
  nand     g02009 ( new_n2386 , new_n2378 , new_n2385 );
  nand     g02010 ( new_n2387 , pi016 , pi067 );
  nand     g02011 ( new_n2388 , pi053 , pi117 );
  nand     g02012 ( new_n2389 , new_n2387 , new_n2388 );
  nand     g02013 ( new_n2390 , pi016 , pi053 );
  nor      g02014 ( new_n2391 , new_n2370 , new_n2390 );
  nand g02015 ( new_n2392 , new_n2391 , new_n2391 );
  nand     g02016 ( new_n2393 , new_n2389 , new_n2392 );
  nand     g02017 ( new_n2394 , pi190 , pi234 );
  nand     g02018 ( new_n2395 , pi092 , pi247 );
  nand     g02019 ( new_n2396 , new_n2394 , new_n2395 );
  or       g02020 ( new_n2397 , new_n2379 , new_n2064 );
  nand     g02021 ( new_n2398 , new_n2396 , new_n2397 );
  nand     g02022 ( new_n2399 , pi080 , pi229 );
  nand     g02023 ( new_n2400 , new_n2380 , new_n2381 );
  nand     g02024 ( new_n2401 , new_n2379 , new_n2382 );
  nand     g02025 ( new_n2402 , new_n2400 , new_n2401 );
  xor      g02026 ( new_n2403 , new_n2399 , new_n2402 );
  xor      g02027 ( new_n2404 , new_n2398 , new_n2403 );
  xnor     g02028 ( new_n2405 , new_n2393 , new_n2404 );
  xor      g02029 ( new_n2406 , new_n2386 , new_n2405 );
  nand     g02030 ( new_n2407 , pi053 , pi103 );
  xor      g02031 ( new_n2408 , new_n2383 , new_n2384 );
  nor      g02032 ( new_n2409 , new_n2407 , new_n2408 );
  xor      g02033 ( new_n2410 , new_n2407 , new_n2408 );
  nand g02034 ( new_n2411 , new_n2410 , new_n2410 );
  nand     g02035 ( new_n2412 , pi067 , pi103 );
  nand     g02036 ( new_n2413 , pi092 , pi117 );
  nand     g02037 ( new_n2414 , pi103 , pi229 );
  nand     g02038 ( new_n2415 , new_n2413 , new_n2414 );
  nand     g02039 ( new_n2416 , pi016 , pi190 );
  xor      g02040 ( new_n2417 , new_n2413 , new_n2414 );
  nand     g02041 ( new_n2418 , new_n2416 , new_n2417 );
  nand     g02042 ( new_n2419 , new_n2415 , new_n2418 );
  nor      g02043 ( new_n2420 , new_n2412 , new_n2419 );
  xor      g02044 ( new_n2421 , new_n2374 , new_n2375 );
  xnor     g02045 ( new_n2422 , new_n2412 , new_n2419 );
  nor      g02046 ( new_n2423 , new_n2421 , new_n2422 );
  nor      g02047 ( new_n2424 , new_n2420 , new_n2423 );
  nor      g02048 ( new_n2425 , new_n2411 , new_n2424 );
  nor      g02049 ( new_n2426 , new_n2409 , new_n2425 );
  nand g02050 ( new_n2427 , new_n2426 , new_n2426 );
  nand     g02051 ( new_n2428 , new_n2406 , new_n2427 );
  nor      g02052 ( new_n2429 , new_n2393 , new_n2404 );
  nor      g02053 ( new_n2430 , new_n2386 , new_n2405 );
  xor      g02054 ( new_n2431 , new_n2392 , new_n2430 );
  nand g02055 ( new_n2432 , new_n2431 , new_n2431 );
  nor      g02056 ( new_n2433 , new_n2429 , new_n2432 );
  nand     g02057 ( new_n2434 , pi067 , pi080 );
  xnor     g02058 ( new_n2435 , new_n2397 , new_n2434 );
  xor      g02059 ( new_n2436 , new_n2064 , new_n2065 );
  xnor     g02060 ( new_n2437 , new_n2435 , new_n2436 );
  nand     g02061 ( new_n2438 , new_n2399 , new_n2402 );
  nand     g02062 ( new_n2439 , new_n2398 , new_n2403 );
  nand     g02063 ( new_n2440 , new_n2438 , new_n2439 );
  nand     g02064 ( new_n2441 , pi030 , pi103 );
  nand     g02065 ( new_n2442 , pi117 , pi185 );
  xor      g02066 ( new_n2443 , new_n2441 , new_n2442 );
  xor      g02067 ( new_n2444 , new_n2390 , new_n2443 );
  xor      g02068 ( new_n2445 , new_n2440 , new_n2444 );
  xnor     g02069 ( new_n2446 , new_n2437 , new_n2445 );
  xor      g02070 ( new_n2447 , new_n2433 , new_n2446 );
  nand     g02071 ( new_n2448 , new_n2428 , new_n2447 );
  xor      g02072 ( new_n2449 , new_n2428 , new_n2447 );
  nand     g02073 ( new_n2450 , pi103 , pi185 );
  xor      g02074 ( new_n2451 , new_n2411 , new_n2424 );
  xor      g02075 ( new_n2452 , new_n2416 , new_n2417 );
  nand g02076 ( new_n2453 , new_n2452 , new_n2452 );
  nand     g02077 ( new_n2454 , pi103 , pi190 );
  nor      g02078 ( new_n2455 , new_n2413 , new_n2454 );
  nand     g02079 ( new_n2456 , new_n2453 , new_n2455 );
  xnor     g02080 ( new_n2457 , new_n2421 , new_n2422 );
  nor      g02081 ( new_n2458 , new_n2456 , new_n2457 );
  nand     g02082 ( new_n2459 , new_n2451 , new_n2458 );
  nand     g02083 ( new_n2460 , new_n2450 , new_n2459 );
  xor      g02084 ( new_n2461 , new_n2450 , new_n2459 );
  xor      g02085 ( new_n2462 , new_n2406 , new_n2426 );
  nand     g02086 ( new_n2463 , new_n2461 , new_n2462 );
  nand     g02087 ( new_n2464 , new_n2460 , new_n2463 );
  nand     g02088 ( new_n2465 , new_n2449 , new_n2464 );
  nand     g02089 ( new_n2466 , new_n2448 , new_n2465 );
  nand     g02090 ( new_n2467 , pi171 , pi209 );
  xor      g02091 ( new_n2468 , new_n2466 , new_n2467 );
  xor      g02092 ( new_n2469 , new_n2369 , new_n2468 );
  nand     g02093 ( new_n2470 , new_n2261 , new_n2262 );
  nand     g02094 ( new_n2471 , new_n2187 , new_n2263 );
  nand     g02095 ( new_n2472 , new_n2470 , new_n2471 );
  nand g02096 ( new_n2473 , new_n2270 , new_n2270 );
  nor      g02097 ( new_n2474 , new_n2473 , new_n2271 );
  nor      g02098 ( new_n2475 , new_n2196 , new_n2272 );
  nor      g02099 ( new_n2476 , new_n2474 , new_n2475 );
  xor      g02100 ( new_n2477 , new_n2472 , new_n2476 );
  xor      g02101 ( new_n2478 , new_n2469 , new_n2477 );
  nand     g02102 ( new_n2479 , pi078 , pi175 );
  nand     g02103 ( new_n2480 , new_n2441 , new_n2442 );
  nand     g02104 ( new_n2481 , new_n2390 , new_n2443 );
  nand     g02105 ( new_n2482 , new_n2480 , new_n2481 );
  xor      g02106 ( new_n2483 , new_n2479 , new_n2482 );
  nand     g02107 ( new_n2484 , new_n2308 , new_n2312 );
  nand g02108 ( new_n2485 , new_n2305 , new_n2305 );
  nand     g02109 ( new_n2486 , new_n2485 , new_n2313 );
  nand     g02110 ( new_n2487 , new_n2484 , new_n2486 );
  nand     g02111 ( new_n2488 , pi190 , pi202 );
  xor      g02112 ( new_n2489 , new_n2487 , new_n2488 );
  nand     g02113 ( new_n2490 , pi124 , pi228 );
  nand     g02114 ( new_n2491 , pi103 , pi220 );
  xor      g02115 ( new_n2492 , new_n2490 , new_n2491 );
  nor      g02116 ( new_n2493 , new_n2197 , new_n2274 );
  nor      g02117 ( new_n2494 , new_n2273 , new_n2275 );
  nor      g02118 ( new_n2495 , new_n2493 , new_n2494 );
  xor      g02119 ( new_n2496 , new_n2492 , new_n2495 );
  xor      g02120 ( new_n2497 , new_n2489 , new_n2496 );
  xor      g02121 ( new_n2498 , new_n2483 , new_n2497 );
  xor      g02122 ( new_n2499 , new_n2478 , new_n2498 );
  nand     g02123 ( new_n2500 , pi134 , pi197 );
  nand g02124 ( new_n2501 , new_n2027 , new_n2027 );
  nor      g02125 ( new_n2502 , new_n2501 , new_n2028 );
  nand g02126 ( new_n2503 , new_n2006 , new_n2006 );
  nor      g02127 ( new_n2504 , new_n2503 , new_n2029 );
  nor      g02128 ( new_n2505 , new_n2502 , new_n2504 );
  nand     g02129 ( new_n2506 , pi229 , pi234 );
  xor      g02130 ( new_n2507 , new_n2505 , new_n2506 );
  xor      g02131 ( new_n2508 , new_n2500 , new_n2507 );
  xor      g02132 ( new_n2509 , new_n2499 , new_n2508 );
  xor      g02133 ( new_n2510 , new_n2368 , new_n2509 );
  xor      g02134 ( new_n2511 , new_n1955 , new_n2510 );
  nand     g02135 ( new_n2512 , pi120 , pi181 );
  nand     g02136 ( new_n2513 , pi149 , pi198 );
  or       g02137 ( new_n2514 , new_n2298 , new_n2314 );
  nand     g02138 ( new_n2515 , new_n2297 , new_n2514 );
  xor      g02139 ( new_n2516 , new_n2513 , new_n2515 );
  nand     g02140 ( new_n2517 , new_n2017 , new_n2018 );
  nand     g02141 ( new_n2518 , new_n1995 , new_n2019 );
  nand     g02142 ( new_n2519 , new_n2517 , new_n2518 );
  nand g02143 ( new_n2520 , new_n2285 , new_n2285 );
  nor      g02144 ( new_n2521 , new_n2520 , new_n2317 );
  nor      g02145 ( new_n2522 , new_n2256 , new_n2318 );
  nor      g02146 ( new_n2523 , new_n2521 , new_n2522 );
  xor      g02147 ( new_n2524 , new_n2519 , new_n2523 );
  or       g02148 ( new_n2525 , new_n2007 , new_n2025 );
  nand     g02149 ( new_n2526 , new_n2026 , new_n2030 );
  nand     g02150 ( new_n2527 , new_n2525 , new_n2526 );
  nand     g02151 ( new_n2528 , pi039 , pi130 );
  nand     g02152 ( new_n2529 , pi167 , pi172 );
  nand     g02153 ( new_n2530 , pi063 , pi158 );
  xor      g02154 ( new_n2531 , new_n2529 , new_n2530 );
  xor      g02155 ( new_n2532 , new_n2528 , new_n2531 );
  xor      g02156 ( new_n2533 , new_n2527 , new_n2532 );
  xor      g02157 ( new_n2534 , new_n2524 , new_n2533 );
  nand     g02158 ( new_n2535 , pi095 , pi245 );
  xor      g02159 ( new_n2536 , new_n2534 , new_n2535 );
  xor      g02160 ( new_n2537 , new_n2516 , new_n2536 );
  xor      g02161 ( new_n2538 , new_n2512 , new_n2537 );
  xor      g02162 ( new_n2539 , new_n2511 , new_n2538 );
  nand     g02163 ( new_n2540 , pi165 , pi240 );
  nand     g02164 ( new_n2541 , pi016 , pi185 );
  xor      g02165 ( new_n2542 , new_n2540 , new_n2541 );
  nor      g02166 ( new_n2543 , new_n2397 , new_n2434 );
  nor      g02167 ( new_n2544 , new_n2435 , new_n2436 );
  nor      g02168 ( new_n2545 , new_n2543 , new_n2544 );
  nor      g02169 ( new_n2546 , new_n1997 , new_n2035 );
  nor      g02170 ( new_n2547 , new_n2032 , new_n2036 );
  nor      g02171 ( new_n2548 , new_n2546 , new_n2547 );
  nand     g02172 ( new_n2549 , pi004 , pi115 );
  nand     g02173 ( new_n2550 , pi053 , pi080 );
  xor      g02174 ( new_n2551 , new_n2549 , new_n2550 );
  xor      g02175 ( new_n2552 , new_n2548 , new_n2551 );
  xor      g02176 ( new_n2553 , new_n2545 , new_n2552 );
  xor      g02177 ( new_n2554 , new_n2542 , new_n2553 );
  nand     g02178 ( new_n2555 , pi062 , pi200 );
  nand     g02179 ( new_n2556 , new_n2440 , new_n2444 );
  nand     g02180 ( new_n2557 , new_n2437 , new_n2445 );
  nand     g02181 ( new_n2558 , new_n2556 , new_n2557 );
  nand     g02182 ( new_n2559 , new_n2020 , new_n2023 );
  nand     g02183 ( new_n2560 , new_n2024 , new_n2031 );
  nand     g02184 ( new_n2561 , new_n2559 , new_n2560 );
  xor      g02185 ( new_n2562 , new_n2558 , new_n2561 );
  xor      g02186 ( new_n2563 , new_n2449 , new_n2464 );
  xor      g02187 ( new_n2564 , new_n2360 , new_n2361 );
  nor      g02188 ( new_n2565 , new_n2563 , new_n2564 );
  xnor     g02189 ( new_n2566 , new_n2563 , new_n2564 );
  xor      g02190 ( new_n2567 , new_n2355 , new_n2356 );
  xor      g02191 ( new_n2568 , new_n2461 , new_n2462 );
  nor      g02192 ( new_n2569 , new_n2567 , new_n2568 );
  xor      g02193 ( new_n2570 , new_n2456 , new_n2457 );
  xnor     g02194 ( new_n2571 , new_n2327 , new_n2347 );
  or       g02195 ( new_n2572 , new_n2570 , new_n2571 );
  xor      g02196 ( new_n2573 , new_n2570 , new_n2571 );
  xor      g02197 ( new_n2574 , new_n2042 , new_n2333 );
  nor      g02198 ( new_n2575 , new_n2454 , new_n2574 );
  nand     g02199 ( new_n2576 , pi092 , pi103 );
  nand     g02200 ( new_n2577 , pi117 , pi190 );
  and      g02201 ( new_n2578 , new_n2576 , new_n2577 );
  nor      g02202 ( new_n2579 , new_n2455 , new_n2578 );
  nand     g02203 ( new_n2580 , new_n2575 , new_n2579 );
  nand g02204 ( new_n2581 , new_n2580 , new_n2580 );
  xor      g02205 ( new_n2582 , new_n2340 , new_n2341 );
  xor      g02206 ( new_n2583 , new_n2575 , new_n2579 );
  nand g02207 ( new_n2584 , new_n2583 , new_n2583 );
  nor      g02208 ( new_n2585 , new_n2582 , new_n2584 );
  nor      g02209 ( new_n2586 , new_n2581 , new_n2585 );
  xor      g02210 ( new_n2587 , new_n2452 , new_n2455 );
  nor      g02211 ( new_n2588 , new_n2586 , new_n2587 );
  xor      g02212 ( new_n2589 , new_n2343 , new_n2345 );
  xor      g02213 ( new_n2590 , new_n2586 , new_n2587 );
  nand g02214 ( new_n2591 , new_n2590 , new_n2590 );
  nor      g02215 ( new_n2592 , new_n2589 , new_n2591 );
  nor      g02216 ( new_n2593 , new_n2588 , new_n2592 );
  nand     g02217 ( new_n2594 , new_n2573 , new_n2593 );
  nand     g02218 ( new_n2595 , new_n2572 , new_n2594 );
  xnor     g02219 ( new_n2596 , new_n2349 , new_n2350 );
  xnor     g02220 ( new_n2597 , new_n2451 , new_n2458 );
  or       g02221 ( new_n2598 , new_n2596 , new_n2597 );
  nand     g02222 ( new_n2599 , new_n2595 , new_n2598 );
  nand     g02223 ( new_n2600 , new_n2596 , new_n2597 );
  nand     g02224 ( new_n2601 , new_n2599 , new_n2600 );
  xnor     g02225 ( new_n2602 , new_n2567 , new_n2568 );
  nor      g02226 ( new_n2603 , new_n2601 , new_n2602 );
  nor      g02227 ( new_n2604 , new_n2569 , new_n2603 );
  nor      g02228 ( new_n2605 , new_n2566 , new_n2604 );
  nor      g02229 ( new_n2606 , new_n2565 , new_n2605 );
  xor      g02230 ( new_n2607 , new_n2562 , new_n2606 );
  xor      g02231 ( new_n2608 , new_n2555 , new_n2607 );
  nand     g02232 ( new_n2609 , pi148 , pi215 );
  nand     g02233 ( new_n2610 , pi154 , pi201 );
  nand     g02234 ( new_n2611 , new_n2260 , new_n2283 );
  nand     g02235 ( new_n2612 , new_n2259 , new_n2284 );
  nand     g02236 ( new_n2613 , new_n2611 , new_n2612 );
  nand     g02237 ( new_n2614 , new_n2391 , new_n2430 );
  nand g02238 ( new_n2615 , new_n2433 , new_n2433 );
  nand     g02239 ( new_n2616 , new_n2615 , new_n2446 );
  nand     g02240 ( new_n2617 , new_n2614 , new_n2616 );
  xor      g02241 ( new_n2618 , new_n2613 , new_n2617 );
  nand     g02242 ( new_n2619 , new_n2117 , new_n2310 );
  nand     g02243 ( new_n2620 , new_n2309 , new_n2311 );
  nand     g02244 ( new_n2621 , new_n2619 , new_n2620 );
  nand g02245 ( new_n2622 , new_n2290 , new_n2290 );
  nor      g02246 ( new_n2623 , new_n2622 , new_n2315 );
  nand g02247 ( new_n2624 , new_n2289 , new_n2289 );
  nor      g02248 ( new_n2625 , new_n2624 , new_n2316 );
  nor      g02249 ( new_n2626 , new_n2623 , new_n2625 );
  xor      g02250 ( new_n2627 , new_n2621 , new_n2626 );
  xor      g02251 ( new_n2628 , new_n2618 , new_n2627 );
  xor      g02252 ( new_n2629 , new_n2610 , new_n2628 );
  nand     g02253 ( new_n2630 , pi107 , pi153 );
  nand     g02254 ( new_n2631 , pi089 , pi156 );
  nand     g02255 ( new_n2632 , pi083 , pi254 );
  xor      g02256 ( new_n2633 , new_n2631 , new_n2632 );
  xor      g02257 ( new_n2634 , new_n2630 , new_n2633 );
  or       g02258 ( new_n2635 , new_n2264 , new_n2268 );
  nand     g02259 ( new_n2636 , new_n2269 , new_n2277 );
  nand     g02260 ( new_n2637 , new_n2635 , new_n2636 );
  nand     g02261 ( new_n2638 , new_n2301 , new_n2302 );
  nand     g02262 ( new_n2639 , new_n2123 , new_n2303 );
  nand     g02263 ( new_n2640 , new_n2638 , new_n2639 );
  nand     g02264 ( new_n2641 , pi003 , pi116 );
  xnor     g02265 ( new_n2642 , new_n2640 , new_n2641 );
  xor      g02266 ( new_n2643 , new_n2637 , new_n2642 );
  xor      g02267 ( new_n2644 , new_n2634 , new_n2643 );
  nand     g02268 ( new_n2645 , new_n2188 , new_n2281 );
  nand g02269 ( new_n2646 , new_n2278 , new_n2278 );
  nand     g02270 ( new_n2647 , new_n2646 , new_n2282 );
  nand     g02271 ( new_n2648 , new_n2645 , new_n2647 );
  nor      g02272 ( new_n2649 , new_n2125 , new_n2299 );
  nor      g02273 ( new_n2650 , new_n2300 , new_n2304 );
  nor      g02274 ( new_n2651 , new_n2649 , new_n2650 );
  xor      g02275 ( new_n2652 , new_n2648 , new_n2651 );
  xor      g02276 ( new_n2653 , new_n2644 , new_n2652 );
  xor      g02277 ( new_n2654 , new_n2629 , new_n2653 );
  xor      g02278 ( new_n2655 , new_n2609 , new_n2654 );
  xor      g02279 ( new_n2656 , new_n2608 , new_n2655 );
  xor      g02280 ( new_n2657 , new_n2554 , new_n2656 );
  xor      g02281 ( po006 , new_n2539 , new_n2657 );
  nand     g02282 ( new_n2659 , pi158 , pi219 );
  nand g02283 ( new_n2660 , pi087 , pi087 );
  nand g02284 ( new_n2661 , pi254 , pi254 );
  nor      g02285 ( new_n2662 , new_n2660 , new_n2661 );
  nor      g02286 ( new_n2663 , new_n2659 , new_n2662 );
  nand     g02287 ( new_n2664 , pi102 , pi254 );
  nand     g02288 ( new_n2665 , pi087 , pi089 );
  or       g02289 ( new_n2666 , new_n2664 , new_n2665 );
  nand     g02290 ( new_n2667 , new_n2664 , new_n2665 );
  and      g02291 ( new_n2668 , new_n2666 , new_n2667 );
  or       g02292 ( new_n2669 , new_n2663 , new_n2668 );
  nor      g02293 ( new_n2670 , new_n2659 , new_n2669 );
  nand g02294 ( new_n2671 , new_n2670 , new_n2670 );
  nand     g02295 ( new_n2672 , new_n2659 , new_n2666 );
  nand     g02296 ( new_n2673 , new_n2667 , new_n2672 );
  nand     g02297 ( new_n2674 , pi087 , pi154 );
  xor      g02298 ( new_n2675 , new_n2673 , new_n2674 );
  nand     g02299 ( new_n2676 , pi001 , pi254 );
  nand     g02300 ( new_n2677 , pi102 , pi158 );
  nand     g02301 ( new_n2678 , pi089 , pi219 );
  xor      g02302 ( new_n2679 , new_n2677 , new_n2678 );
  xor      g02303 ( new_n2680 , new_n2676 , new_n2679 );
  xor      g02304 ( new_n2681 , new_n2675 , new_n2680 );
  nor      g02305 ( new_n2682 , new_n2671 , new_n2681 );
  nor      g02306 ( new_n2683 , new_n2673 , new_n2674 );
  nand g02307 ( new_n2684 , new_n2675 , new_n2675 );
  nor      g02308 ( new_n2685 , new_n2684 , new_n2680 );
  nor      g02309 ( new_n2686 , new_n2683 , new_n2685 );
  nand     g02310 ( new_n2687 , pi087 , pi095 );
  nand     g02311 ( new_n2688 , pi089 , pi102 );
  nand     g02312 ( new_n2689 , pi001 , pi158 );
  nand     g02313 ( new_n2690 , pi122 , pi254 );
  xor      g02314 ( new_n2691 , new_n2689 , new_n2690 );
  xor      g02315 ( new_n2692 , new_n2688 , new_n2691 );
  nand     g02316 ( new_n2693 , pi154 , pi219 );
  nand     g02317 ( new_n2694 , new_n2677 , new_n2678 );
  nand     g02318 ( new_n2695 , new_n2676 , new_n2679 );
  nand     g02319 ( new_n2696 , new_n2694 , new_n2695 );
  xor      g02320 ( new_n2697 , new_n2693 , new_n2696 );
  xor      g02321 ( new_n2698 , new_n2692 , new_n2697 );
  xor      g02322 ( new_n2699 , new_n2687 , new_n2698 );
  nand g02323 ( new_n2700 , new_n2699 , new_n2699 );
  xor      g02324 ( new_n2701 , new_n2686 , new_n2700 );
  xor      g02325 ( new_n2702 , new_n2682 , new_n2701 );
  nand     g02326 ( new_n2703 , pi004 , pi071 );
  nand     g02327 ( new_n2704 , pi142 , pi170 );
  nand g02328 ( new_n2705 , new_n2704 , new_n2704 );
  nor      g02329 ( new_n2706 , new_n2703 , new_n2705 );
  nand     g02330 ( new_n2707 , pi169 , pi170 );
  nand     g02331 ( new_n2708 , pi073 , pi142 );
  or       g02332 ( new_n2709 , new_n2707 , new_n2708 );
  nand     g02333 ( new_n2710 , new_n2707 , new_n2708 );
  and      g02334 ( new_n2711 , new_n2709 , new_n2710 );
  or       g02335 ( new_n2712 , new_n2706 , new_n2711 );
  nor      g02336 ( new_n2713 , new_n2703 , new_n2712 );
  nand     g02337 ( new_n2714 , new_n2703 , new_n2709 );
  nand     g02338 ( new_n2715 , new_n2710 , new_n2714 );
  nand     g02339 ( new_n2716 , pi003 , pi142 );
  xor      g02340 ( new_n2717 , new_n2715 , new_n2716 );
  nand     g02341 ( new_n2718 , pi123 , pi170 );
  nand     g02342 ( new_n2719 , pi004 , pi169 );
  nand     g02343 ( new_n2720 , pi071 , pi073 );
  xor      g02344 ( new_n2721 , new_n2719 , new_n2720 );
  xor      g02345 ( new_n2722 , new_n2718 , new_n2721 );
  xor      g02346 ( new_n2723 , new_n2717 , new_n2722 );
  nand g02347 ( new_n2724 , new_n2723 , new_n2723 );
  nand     g02348 ( new_n2725 , new_n2713 , new_n2724 );
  nand     g02349 ( new_n2726 , pi130 , pi142 );
  nand     g02350 ( new_n2727 , pi099 , pi170 );
  nand     g02351 ( new_n2728 , pi073 , pi169 );
  nand     g02352 ( new_n2729 , pi004 , pi123 );
  xor      g02353 ( new_n2730 , new_n2728 , new_n2729 );
  xor      g02354 ( new_n2731 , new_n2727 , new_n2730 );
  nand     g02355 ( new_n2732 , pi003 , pi071 );
  nand     g02356 ( new_n2733 , new_n2719 , new_n2720 );
  nand     g02357 ( new_n2734 , new_n2718 , new_n2721 );
  nand     g02358 ( new_n2735 , new_n2733 , new_n2734 );
  xor      g02359 ( new_n2736 , new_n2732 , new_n2735 );
  xor      g02360 ( new_n2737 , new_n2731 , new_n2736 );
  xor      g02361 ( new_n2738 , new_n2726 , new_n2737 );
  nor      g02362 ( new_n2739 , new_n2715 , new_n2716 );
  nand g02363 ( new_n2740 , new_n2717 , new_n2717 );
  nor      g02364 ( new_n2741 , new_n2740 , new_n2722 );
  nor      g02365 ( new_n2742 , new_n2739 , new_n2741 );
  xor      g02366 ( new_n2743 , new_n2738 , new_n2742 );
  xor      g02367 ( new_n2744 , new_n2725 , new_n2743 );
  nand     g02368 ( new_n2745 , new_n2702 , new_n2744 );
  nand g02369 ( new_n2746 , new_n2745 , new_n2745 );
  xor      g02370 ( new_n2747 , new_n2670 , new_n2681 );
  nand g02371 ( new_n2748 , new_n2747 , new_n2747 );
  nand     g02372 ( new_n2749 , new_n2710 , new_n2706 );
  nand     g02373 ( new_n2750 , new_n2712 , new_n2749 );
  nand     g02374 ( new_n2751 , new_n2663 , new_n2667 );
  nand     g02375 ( new_n2752 , new_n2669 , new_n2751 );
  or       g02376 ( new_n2753 , new_n2750 , new_n2752 );
  nand     g02377 ( new_n2754 , new_n2750 , new_n2752 );
  nand     g02378 ( new_n2755 , pi087 , pi254 );
  nor      g02379 ( new_n2756 , new_n2755 , new_n2704 );
  nand     g02380 ( new_n2757 , pi087 , pi158 );
  nand     g02381 ( new_n2758 , pi219 , pi254 );
  xor      g02382 ( new_n2759 , new_n2757 , new_n2758 );
  nand     g02383 ( new_n2760 , new_n2756 , new_n2759 );
  nand     g02384 ( new_n2761 , pi004 , pi142 );
  nand     g02385 ( new_n2762 , pi071 , pi170 );
  xor      g02386 ( new_n2763 , new_n2761 , new_n2762 );
  xor      g02387 ( new_n2764 , new_n2756 , new_n2759 );
  nand     g02388 ( new_n2765 , new_n2763 , new_n2764 );
  nand     g02389 ( new_n2766 , new_n2760 , new_n2765 );
  nand     g02390 ( new_n2767 , new_n2754 , new_n2766 );
  nand     g02391 ( new_n2768 , new_n2753 , new_n2767 );
  nor      g02392 ( new_n2769 , new_n2748 , new_n2768 );
  nand g02393 ( new_n2770 , new_n2769 , new_n2769 );
  xor      g02394 ( new_n2771 , new_n2713 , new_n2724 );
  nand g02395 ( new_n2772 , new_n2771 , new_n2771 );
  xor      g02396 ( new_n2773 , new_n2748 , new_n2768 );
  nand     g02397 ( new_n2774 , new_n2772 , new_n2773 );
  nand     g02398 ( new_n2775 , new_n2770 , new_n2774 );
  xnor     g02399 ( new_n2776 , new_n2702 , new_n2744 );
  nor      g02400 ( new_n2777 , new_n2775 , new_n2776 );
  nor      g02401 ( new_n2778 , new_n2746 , new_n2777 );
  nand     g02402 ( new_n2779 , new_n2682 , new_n2701 );
  nand     g02403 ( new_n2780 , pi006 , pi087 );
  xor      g02404 ( new_n2781 , new_n2779 , new_n2780 );
  nand     g02405 ( new_n2782 , pi095 , pi219 );
  nand     g02406 ( new_n2783 , pi102 , pi154 );
  nand     g02407 ( new_n2784 , new_n2782 , new_n2783 );
  nand     g02408 ( new_n2785 , pi095 , pi102 );
  nor      g02409 ( new_n2786 , new_n2693 , new_n2785 );
  nand g02410 ( new_n2787 , new_n2786 , new_n2786 );
  nand     g02411 ( new_n2788 , new_n2784 , new_n2787 );
  nand     g02412 ( new_n2789 , pi122 , pi158 );
  nand     g02413 ( new_n2790 , pi135 , pi254 );
  nand     g02414 ( new_n2791 , new_n2789 , new_n2790 );
  nand     g02415 ( new_n2792 , pi135 , pi158 );
  nor      g02416 ( new_n2793 , new_n2690 , new_n2792 );
  nand g02417 ( new_n2794 , new_n2793 , new_n2793 );
  nand     g02418 ( new_n2795 , new_n2791 , new_n2794 );
  nand     g02419 ( new_n2796 , pi001 , pi089 );
  nand     g02420 ( new_n2797 , new_n2689 , new_n2690 );
  nand     g02421 ( new_n2798 , new_n2688 , new_n2691 );
  nand     g02422 ( new_n2799 , new_n2797 , new_n2798 );
  xor      g02423 ( new_n2800 , new_n2796 , new_n2799 );
  xor      g02424 ( new_n2801 , new_n2795 , new_n2800 );
  xor      g02425 ( new_n2802 , new_n2788 , new_n2801 );
  nand g02426 ( new_n2803 , new_n2802 , new_n2802 );
  nand     g02427 ( new_n2804 , new_n2693 , new_n2696 );
  nand     g02428 ( new_n2805 , new_n2692 , new_n2697 );
  nand     g02429 ( new_n2806 , new_n2804 , new_n2805 );
  xor      g02430 ( new_n2807 , new_n2803 , new_n2806 );
  nor      g02431 ( new_n2808 , new_n2687 , new_n2698 );
  nor      g02432 ( new_n2809 , new_n2686 , new_n2700 );
  nor      g02433 ( new_n2810 , new_n2808 , new_n2809 );
  xor      g02434 ( new_n2811 , new_n2807 , new_n2810 );
  xor      g02435 ( new_n2812 , new_n2781 , new_n2811 );
  nor      g02436 ( new_n2813 , new_n2726 , new_n2737 );
  nand g02437 ( new_n2814 , new_n2738 , new_n2738 );
  nor      g02438 ( new_n2815 , new_n2814 , new_n2742 );
  nor      g02439 ( new_n2816 , new_n2813 , new_n2815 );
  nand     g02440 ( new_n2817 , new_n2732 , new_n2735 );
  nand     g02441 ( new_n2818 , new_n2731 , new_n2736 );
  nand     g02442 ( new_n2819 , new_n2817 , new_n2818 );
  nand     g02443 ( new_n2820 , pi071 , pi130 );
  nand     g02444 ( new_n2821 , pi003 , pi169 );
  nand     g02445 ( new_n2822 , new_n2820 , new_n2821 );
  nand     g02446 ( new_n2823 , pi130 , pi169 );
  nor      g02447 ( new_n2824 , new_n2732 , new_n2823 );
  nand g02448 ( new_n2825 , new_n2824 , new_n2824 );
  nand     g02449 ( new_n2826 , new_n2822 , new_n2825 );
  nand     g02450 ( new_n2827 , pi004 , pi099 );
  nand     g02451 ( new_n2828 , pi023 , pi170 );
  nand     g02452 ( new_n2829 , new_n2827 , new_n2828 );
  nand     g02453 ( new_n2830 , pi004 , pi023 );
  nor      g02454 ( new_n2831 , new_n2727 , new_n2830 );
  nand g02455 ( new_n2832 , new_n2831 , new_n2831 );
  nand     g02456 ( new_n2833 , new_n2829 , new_n2832 );
  nand     g02457 ( new_n2834 , pi073 , pi123 );
  nand     g02458 ( new_n2835 , new_n2728 , new_n2729 );
  nand     g02459 ( new_n2836 , new_n2727 , new_n2730 );
  nand     g02460 ( new_n2837 , new_n2835 , new_n2836 );
  xor      g02461 ( new_n2838 , new_n2834 , new_n2837 );
  xor      g02462 ( new_n2839 , new_n2833 , new_n2838 );
  xor      g02463 ( new_n2840 , new_n2826 , new_n2839 );
  xor      g02464 ( new_n2841 , new_n2819 , new_n2840 );
  xnor     g02465 ( new_n2842 , new_n2816 , new_n2841 );
  nor      g02466 ( new_n2843 , new_n2725 , new_n2743 );
  nand     g02467 ( new_n2844 , pi124 , pi142 );
  xor      g02468 ( new_n2845 , new_n2843 , new_n2844 );
  xor      g02469 ( new_n2846 , new_n2842 , new_n2845 );
  xor      g02470 ( new_n2847 , new_n2812 , new_n2846 );
  xnor     g02471 ( new_n2848 , new_n2778 , new_n2847 );
  nand     g02472 ( new_n2849 , pi138 , pi198 );
  nand     g02473 ( new_n2850 , pi062 , pi216 );
  nand     g02474 ( new_n2851 , pi065 , pi076 );
  nand     g02475 ( new_n2852 , pi041 , pi120 );
  xor      g02476 ( new_n2853 , new_n2851 , new_n2852 );
  xor      g02477 ( new_n2854 , new_n2850 , new_n2853 );
  nand     g02478 ( new_n2855 , pi172 , pi182 );
  nand     g02479 ( new_n2856 , pi041 , pi062 );
  nand     g02480 ( new_n2857 , pi065 , pi216 );
  nand     g02481 ( new_n2858 , new_n2856 , new_n2857 );
  nand     g02482 ( new_n2859 , pi120 , pi182 );
  xor      g02483 ( new_n2860 , new_n2856 , new_n2857 );
  nand     g02484 ( new_n2861 , new_n2859 , new_n2860 );
  nand     g02485 ( new_n2862 , new_n2858 , new_n2861 );
  xor      g02486 ( new_n2863 , new_n2855 , new_n2862 );
  xor      g02487 ( new_n2864 , new_n2854 , new_n2863 );
  nor      g02488 ( new_n2865 , new_n2849 , new_n2864 );
  nand     g02489 ( new_n2866 , pi138 , pi172 );
  nand     g02490 ( new_n2867 , pi120 , pi138 );
  nand     g02491 ( new_n2868 , pi062 , pi182 );
  nand     g02492 ( new_n2869 , new_n2867 , new_n2868 );
  nand     g02493 ( new_n2870 , pi041 , pi065 );
  xor      g02494 ( new_n2871 , new_n2867 , new_n2868 );
  nand     g02495 ( new_n2872 , new_n2870 , new_n2871 );
  nand     g02496 ( new_n2873 , new_n2869 , new_n2872 );
  nor      g02497 ( new_n2874 , new_n2866 , new_n2873 );
  xor      g02498 ( new_n2875 , new_n2859 , new_n2860 );
  nand g02499 ( new_n2876 , new_n2875 , new_n2875 );
  xor      g02500 ( new_n2877 , new_n2866 , new_n2873 );
  nand     g02501 ( new_n2878 , new_n2876 , new_n2877 );
  nand g02502 ( new_n2879 , new_n2878 , new_n2878 );
  nor      g02503 ( new_n2880 , new_n2874 , new_n2879 );
  nand g02504 ( new_n2881 , new_n2880 , new_n2880 );
  xor      g02505 ( new_n2882 , new_n2849 , new_n2864 );
  nand     g02506 ( new_n2883 , new_n2881 , new_n2882 );
  nand g02507 ( new_n2884 , new_n2883 , new_n2883 );
  or       g02508 ( new_n2885 , new_n2865 , new_n2884 );
  nand     g02509 ( new_n2886 , pi041 , pi172 );
  nand     g02510 ( new_n2887 , pi182 , pi198 );
  and      g02511 ( new_n2888 , new_n2886 , new_n2887 );
  nand     g02512 ( new_n2889 , pi041 , pi198 );
  nor      g02513 ( new_n2890 , new_n2855 , new_n2889 );
  or       g02514 ( new_n2891 , new_n2888 , new_n2890 );
  nand     g02515 ( new_n2892 , new_n2851 , new_n2852 );
  nand     g02516 ( new_n2893 , new_n2850 , new_n2853 );
  nand     g02517 ( new_n2894 , new_n2892 , new_n2893 );
  nand     g02518 ( new_n2895 , pi120 , pi216 );
  nand     g02519 ( new_n2896 , pi062 , pi076 );
  nand     g02520 ( new_n2897 , pi065 , pi079 );
  nand     g02521 ( new_n2898 , new_n2896 , new_n2897 );
  nand     g02522 ( new_n2899 , pi062 , pi079 );
  nor      g02523 ( new_n2900 , new_n2851 , new_n2899 );
  nand g02524 ( new_n2901 , new_n2900 , new_n2900 );
  nand     g02525 ( new_n2902 , new_n2898 , new_n2901 );
  xor      g02526 ( new_n2903 , new_n2895 , new_n2902 );
  xor      g02527 ( new_n2904 , new_n2894 , new_n2903 );
  xor      g02528 ( new_n2905 , new_n2891 , new_n2904 );
  nand     g02529 ( new_n2906 , new_n2855 , new_n2862 );
  nand     g02530 ( new_n2907 , new_n2854 , new_n2863 );
  nand     g02531 ( new_n2908 , new_n2906 , new_n2907 );
  xor      g02532 ( new_n2909 , new_n2905 , new_n2908 );
  xor      g02533 ( new_n2910 , new_n2885 , new_n2909 );
  xor      g02534 ( new_n2911 , new_n2870 , new_n2871 );
  nand g02535 ( new_n2912 , new_n2911 , new_n2911 );
  nand     g02536 ( new_n2913 , pi065 , pi138 );
  nor      g02537 ( new_n2914 , new_n2868 , new_n2913 );
  nand     g02538 ( new_n2915 , new_n2912 , new_n2914 );
  xor      g02539 ( new_n2916 , new_n2875 , new_n2877 );
  or       g02540 ( new_n2917 , new_n2915 , new_n2916 );
  xor      g02541 ( new_n2918 , new_n2880 , new_n2882 );
  nor      g02542 ( new_n2919 , new_n2917 , new_n2918 );
  nand     g02543 ( new_n2920 , pi138 , pi165 );
  xor      g02544 ( new_n2921 , new_n2919 , new_n2920 );
  xor      g02545 ( new_n2922 , new_n2910 , new_n2921 );
  nand g02546 ( new_n2923 , new_n2922 , new_n2922 );
  nor      g02547 ( new_n2924 , new_n2848 , new_n2923 );
  xor      g02548 ( new_n2925 , new_n2917 , new_n2918 );
  xor      g02549 ( new_n2926 , new_n2915 , new_n2916 );
  xor      g02550 ( new_n2927 , new_n2771 , new_n2773 );
  nor      g02551 ( new_n2928 , new_n2926 , new_n2927 );
  xor      g02552 ( new_n2929 , new_n2755 , new_n2704 );
  nand g02553 ( new_n2930 , new_n2929 , new_n2929 );
  nor      g02554 ( new_n2931 , new_n2913 , new_n2930 );
  nand g02555 ( new_n2932 , new_n2931 , new_n2931 );
  nand     g02556 ( new_n2933 , pi062 , pi138 );
  nand     g02557 ( new_n2934 , pi065 , pi182 );
  and      g02558 ( new_n2935 , new_n2933 , new_n2934 );
  or       g02559 ( new_n2936 , new_n2914 , new_n2935 );
  nand     g02560 ( new_n2937 , new_n2932 , new_n2936 );
  xor      g02561 ( new_n2938 , new_n2932 , new_n2936 );
  xnor     g02562 ( new_n2939 , new_n2763 , new_n2764 );
  nand     g02563 ( new_n2940 , new_n2938 , new_n2939 );
  nand     g02564 ( new_n2941 , new_n2937 , new_n2940 );
  xor      g02565 ( new_n2942 , new_n2912 , new_n2914 );
  nand g02566 ( new_n2943 , new_n2942 , new_n2942 );
  nor      g02567 ( new_n2944 , new_n2941 , new_n2943 );
  nand g02568 ( new_n2945 , new_n2944 , new_n2944 );
  xor      g02569 ( new_n2946 , new_n2941 , new_n2943 );
  xor      g02570 ( new_n2947 , new_n2750 , new_n2752 );
  xor      g02571 ( new_n2948 , new_n2766 , new_n2947 );
  nand     g02572 ( new_n2949 , new_n2946 , new_n2948 );
  nand     g02573 ( new_n2950 , new_n2945 , new_n2949 );
  xnor     g02574 ( new_n2951 , new_n2926 , new_n2927 );
  nor      g02575 ( new_n2952 , new_n2950 , new_n2951 );
  nor      g02576 ( new_n2953 , new_n2928 , new_n2952 );
  nor      g02577 ( new_n2954 , new_n2925 , new_n2953 );
  xnor     g02578 ( new_n2955 , new_n2775 , new_n2776 );
  xor      g02579 ( new_n2956 , new_n2925 , new_n2953 );
  and      g02580 ( new_n2957 , new_n2955 , new_n2956 );
  or       g02581 ( new_n2958 , new_n2954 , new_n2957 );
  xor      g02582 ( new_n2959 , new_n2848 , new_n2922 );
  nor      g02583 ( new_n2960 , new_n2958 , new_n2959 );
  nor      g02584 ( new_n2961 , new_n2924 , new_n2960 );
  nand g02585 ( new_n2962 , new_n2919 , new_n2919 );
  nand     g02586 ( new_n2963 , new_n2962 , new_n2920 );
  nand g02587 ( new_n2964 , new_n2921 , new_n2921 );
  nand     g02588 ( new_n2965 , new_n2910 , new_n2964 );
  nand     g02589 ( new_n2966 , new_n2963 , new_n2965 );
  nand g02590 ( new_n2967 , new_n2885 , new_n2885 );
  or       g02591 ( new_n2968 , new_n2967 , new_n2909 );
  nand g02592 ( new_n2969 , new_n2905 , new_n2905 );
  nor      g02593 ( new_n2970 , new_n2969 , new_n2908 );
  and      g02594 ( new_n2971 , new_n2890 , new_n2970 );
  nor      g02595 ( new_n2972 , new_n2891 , new_n2904 );
  nor      g02596 ( new_n2973 , new_n2890 , new_n2972 );
  nand g02597 ( new_n2974 , new_n2973 , new_n2973 );
  nor      g02598 ( new_n2975 , new_n2970 , new_n2974 );
  or       g02599 ( new_n2976 , new_n2971 , new_n2975 );
  nand     g02600 ( new_n2977 , pi172 , pi216 );
  xor      g02601 ( new_n2978 , new_n2900 , new_n2977 );
  nand     g02602 ( new_n2979 , pi076 , pi120 );
  nand     g02603 ( new_n2980 , pi065 , pi251 );
  xor      g02604 ( new_n2981 , new_n2979 , new_n2980 );
  xor      g02605 ( new_n2982 , new_n2899 , new_n2981 );
  xor      g02606 ( new_n2983 , new_n2978 , new_n2982 );
  nand     g02607 ( new_n2984 , new_n2895 , new_n2902 );
  nand     g02608 ( new_n2985 , new_n2894 , new_n2903 );
  nand     g02609 ( new_n2986 , new_n2984 , new_n2985 );
  nand     g02610 ( new_n2987 , pi138 , pi197 );
  nand     g02611 ( new_n2988 , pi165 , pi182 );
  xor      g02612 ( new_n2989 , new_n2987 , new_n2988 );
  xor      g02613 ( new_n2990 , new_n2889 , new_n2989 );
  xor      g02614 ( new_n2991 , new_n2986 , new_n2990 );
  xor      g02615 ( new_n2992 , new_n2983 , new_n2991 );
  xor      g02616 ( new_n2993 , new_n2976 , new_n2992 );
  xnor     g02617 ( new_n2994 , new_n2968 , new_n2993 );
  xnor     g02618 ( new_n2995 , new_n2966 , new_n2994 );
  nand g02619 ( new_n2996 , new_n2846 , new_n2846 );
  nor      g02620 ( new_n2997 , new_n2812 , new_n2996 );
  nor      g02621 ( new_n2998 , new_n2778 , new_n2847 );
  nor      g02622 ( new_n2999 , new_n2997 , new_n2998 );
  nand     g02623 ( new_n3000 , new_n2779 , new_n2780 );
  nand     g02624 ( new_n3001 , new_n2781 , new_n2811 );
  nand     g02625 ( new_n3002 , new_n3000 , new_n3001 );
  nand g02626 ( new_n3003 , new_n2807 , new_n2807 );
  nor      g02627 ( new_n3004 , new_n3003 , new_n2810 );
  nand g02628 ( new_n3005 , new_n3004 , new_n3004 );
  nand     g02629 ( new_n3006 , pi001 , pi154 );
  xor      g02630 ( new_n3007 , new_n2793 , new_n3006 );
  nand     g02631 ( new_n3008 , pi089 , pi122 );
  nand     g02632 ( new_n3009 , pi059 , pi254 );
  xor      g02633 ( new_n3010 , new_n3008 , new_n3009 );
  xor      g02634 ( new_n3011 , new_n2792 , new_n3010 );
  xnor     g02635 ( new_n3012 , new_n3007 , new_n3011 );
  nand     g02636 ( new_n3013 , new_n2796 , new_n2799 );
  nand     g02637 ( new_n3014 , new_n2795 , new_n2800 );
  nand     g02638 ( new_n3015 , new_n3013 , new_n3014 );
  nand     g02639 ( new_n3016 , pi087 , pi209 );
  nand     g02640 ( new_n3017 , pi006 , pi219 );
  xor      g02641 ( new_n3018 , new_n2785 , new_n3017 );
  xor      g02642 ( new_n3019 , new_n3016 , new_n3018 );
  xnor     g02643 ( new_n3020 , new_n3015 , new_n3019 );
  xor      g02644 ( new_n3021 , new_n3012 , new_n3020 );
  nor      g02645 ( new_n3022 , new_n2803 , new_n2806 );
  nand     g02646 ( new_n3023 , new_n2786 , new_n3022 );
  or       g02647 ( new_n3024 , new_n2788 , new_n2801 );
  nand     g02648 ( new_n3025 , new_n2787 , new_n3024 );
  or       g02649 ( new_n3026 , new_n3022 , new_n3025 );
  nand     g02650 ( new_n3027 , new_n3023 , new_n3026 );
  xor      g02651 ( new_n3028 , new_n3021 , new_n3027 );
  xor      g02652 ( new_n3029 , new_n3005 , new_n3028 );
  xor      g02653 ( new_n3030 , new_n3002 , new_n3029 );
  nand g02654 ( new_n3031 , new_n2843 , new_n2843 );
  nand     g02655 ( new_n3032 , new_n3031 , new_n2844 );
  nand g02656 ( new_n3033 , new_n2845 , new_n2845 );
  nand     g02657 ( new_n3034 , new_n2842 , new_n3033 );
  nand     g02658 ( new_n3035 , new_n3032 , new_n3034 );
  nor      g02659 ( new_n3036 , new_n2816 , new_n2841 );
  nand     g02660 ( new_n3037 , new_n2826 , new_n2839 );
  nand     g02661 ( new_n3038 , new_n2819 , new_n2840 );
  nand     g02662 ( new_n3039 , new_n3037 , new_n3038 );
  xor      g02663 ( new_n3040 , new_n2825 , new_n3039 );
  nand     g02664 ( new_n3041 , new_n2834 , new_n2837 );
  nand     g02665 ( new_n3042 , new_n2833 , new_n2838 );
  nand     g02666 ( new_n3043 , new_n3041 , new_n3042 );
  nand     g02667 ( new_n3044 , pi142 , pi215 );
  nand     g02668 ( new_n3045 , pi071 , pi124 );
  xor      g02669 ( new_n3046 , new_n3044 , new_n3045 );
  xor      g02670 ( new_n3047 , new_n2823 , new_n3046 );
  xnor     g02671 ( new_n3048 , new_n3043 , new_n3047 );
  nand     g02672 ( new_n3049 , pi003 , pi123 );
  xor      g02673 ( new_n3050 , new_n2831 , new_n3049 );
  nand     g02674 ( new_n3051 , pi073 , pi099 );
  nand     g02675 ( new_n3052 , pi155 , pi170 );
  xor      g02676 ( new_n3053 , new_n3051 , new_n3052 );
  xor      g02677 ( new_n3054 , new_n2830 , new_n3053 );
  xnor     g02678 ( new_n3055 , new_n3050 , new_n3054 );
  xor      g02679 ( new_n3056 , new_n3048 , new_n3055 );
  nand g02680 ( new_n3057 , new_n3056 , new_n3056 );
  xor      g02681 ( new_n3058 , new_n3040 , new_n3057 );
  xor      g02682 ( new_n3059 , new_n3036 , new_n3058 );
  xnor     g02683 ( new_n3060 , new_n3035 , new_n3059 );
  xnor     g02684 ( new_n3061 , new_n3030 , new_n3060 );
  xnor     g02685 ( new_n3062 , new_n2999 , new_n3061 );
  xor      g02686 ( new_n3063 , new_n2995 , new_n3062 );
  xor      g02687 ( new_n3064 , new_n2961 , new_n3063 );
  nand     g02688 ( new_n3065 , pi101 , pi190 );
  nand     g02689 ( new_n3066 , pi092 , pi225 );
  nor      g02690 ( new_n3067 , new_n3065 , new_n3066 );
  nand     g02691 ( new_n3068 , pi067 , pi223 );
  xor      g02692 ( new_n3069 , new_n3067 , new_n3068 );
  nand     g02693 ( new_n3070 , pi177 , pi190 );
  nand     g02694 ( new_n3071 , pi101 , pi229 );
  xor      g02695 ( new_n3072 , new_n3070 , new_n3071 );
  xor      g02696 ( new_n3073 , new_n3066 , new_n3072 );
  xnor     g02697 ( new_n3074 , new_n3069 , new_n3073 );
  nand     g02698 ( new_n3075 , pi053 , pi060 );
  nand     g02699 ( new_n3076 , pi030 , pi160 );
  nand     g02700 ( new_n3077 , pi020 , pi185 );
  xor      g02701 ( new_n3078 , new_n3076 , new_n3077 );
  xor      g02702 ( new_n3079 , new_n3075 , new_n3078 );
  nand     g02703 ( new_n3080 , pi060 , pi229 );
  nand     g02704 ( new_n3081 , pi092 , pi223 );
  nand     g02705 ( new_n3082 , new_n3080 , new_n3081 );
  xor      g02706 ( new_n3083 , new_n3080 , new_n3081 );
  nand     g02707 ( new_n3084 , new_n3065 , new_n3083 );
  nand     g02708 ( new_n3085 , new_n3082 , new_n3084 );
  nand g02709 ( new_n3086 , new_n3067 , new_n3067 );
  nand     g02710 ( new_n3087 , pi190 , pi225 );
  nand     g02711 ( new_n3088 , pi092 , pi101 );
  nand     g02712 ( new_n3089 , new_n3087 , new_n3088 );
  nand     g02713 ( new_n3090 , new_n3086 , new_n3089 );
  nor      g02714 ( new_n3091 , new_n3085 , new_n3090 );
  nand     g02715 ( new_n3092 , pi223 , pi229 );
  xor      g02716 ( new_n3093 , new_n3085 , new_n3090 );
  nand g02717 ( new_n3094 , new_n3093 , new_n3093 );
  nor      g02718 ( new_n3095 , new_n3092 , new_n3094 );
  nor      g02719 ( new_n3096 , new_n3091 , new_n3095 );
  xor      g02720 ( new_n3097 , new_n3079 , new_n3096 );
  xnor     g02721 ( new_n3098 , new_n3074 , new_n3097 );
  nand     g02722 ( new_n3099 , pi020 , pi067 );
  nor      g02723 ( new_n3100 , new_n3075 , new_n3099 );
  nand g02724 ( new_n3101 , new_n3100 , new_n3100 );
  nand     g02725 ( new_n3102 , pi060 , pi092 );
  nand     g02726 ( new_n3103 , pi020 , pi229 );
  nand     g02727 ( new_n3104 , new_n3102 , new_n3103 );
  nand     g02728 ( new_n3105 , pi190 , pi223 );
  xor      g02729 ( new_n3106 , new_n3102 , new_n3103 );
  nand     g02730 ( new_n3107 , new_n3105 , new_n3106 );
  nand     g02731 ( new_n3108 , new_n3104 , new_n3107 );
  nand     g02732 ( new_n3109 , new_n3099 , new_n3108 );
  xor      g02733 ( new_n3110 , new_n3065 , new_n3083 );
  xor      g02734 ( new_n3111 , new_n3099 , new_n3108 );
  nand     g02735 ( new_n3112 , new_n3110 , new_n3111 );
  nand     g02736 ( new_n3113 , new_n3109 , new_n3112 );
  xor      g02737 ( new_n3114 , new_n3092 , new_n3093 );
  nand     g02738 ( new_n3115 , new_n3113 , new_n3114 );
  nand     g02739 ( new_n3116 , pi060 , pi067 );
  nand     g02740 ( new_n3117 , pi020 , pi053 );
  nand     g02741 ( new_n3118 , new_n3116 , new_n3117 );
  nand     g02742 ( new_n3119 , new_n3101 , new_n3118 );
  xor      g02743 ( new_n3120 , new_n3113 , new_n3114 );
  nand     g02744 ( new_n3121 , new_n3119 , new_n3120 );
  nand     g02745 ( new_n3122 , new_n3115 , new_n3121 );
  nand     g02746 ( new_n3123 , new_n3101 , new_n3122 );
  nor      g02747 ( new_n3124 , new_n3113 , new_n3114 );
  nand     g02748 ( new_n3125 , new_n3100 , new_n3124 );
  nand     g02749 ( new_n3126 , new_n3123 , new_n3125 );
  xor      g02750 ( new_n3127 , new_n3098 , new_n3126 );
  xor      g02751 ( new_n3128 , new_n3119 , new_n3120 );
  nand     g02752 ( new_n3129 , pi053 , pi160 );
  xor      g02753 ( new_n3130 , new_n3110 , new_n3111 );
  nor      g02754 ( new_n3131 , new_n3129 , new_n3130 );
  xor      g02755 ( new_n3132 , new_n3129 , new_n3130 );
  nand g02756 ( new_n3133 , new_n3132 , new_n3132 );
  nand     g02757 ( new_n3134 , pi020 , pi092 );
  nand     g02758 ( new_n3135 , pi060 , pi190 );
  nand     g02759 ( new_n3136 , pi160 , pi229 );
  or       g02760 ( new_n3137 , new_n3135 , new_n3136 );
  nand     g02761 ( new_n3138 , new_n3134 , new_n3137 );
  nand     g02762 ( new_n3139 , new_n3135 , new_n3136 );
  nand     g02763 ( new_n3140 , new_n3138 , new_n3139 );
  nand     g02764 ( new_n3141 , pi067 , pi160 );
  nor      g02765 ( new_n3142 , new_n3140 , new_n3141 );
  xor      g02766 ( new_n3143 , new_n3140 , new_n3141 );
  nand g02767 ( new_n3144 , new_n3143 , new_n3143 );
  xor      g02768 ( new_n3145 , new_n3105 , new_n3106 );
  nor      g02769 ( new_n3146 , new_n3144 , new_n3145 );
  nor      g02770 ( new_n3147 , new_n3142 , new_n3146 );
  nor      g02771 ( new_n3148 , new_n3133 , new_n3147 );
  nor      g02772 ( new_n3149 , new_n3131 , new_n3148 );
  nor      g02773 ( new_n3150 , new_n3128 , new_n3149 );
  xor      g02774 ( new_n3151 , new_n3127 , new_n3150 );
  nand     g02775 ( new_n3152 , pi160 , pi185 );
  xor      g02776 ( new_n3153 , new_n3133 , new_n3147 );
  nand     g02777 ( new_n3154 , pi160 , pi190 );
  nand g02778 ( new_n3155 , new_n3154 , new_n3154 );
  nor      g02779 ( new_n3156 , new_n3134 , new_n3155 );
  or       g02780 ( new_n3157 , new_n3139 , new_n3156 );
  nand     g02781 ( new_n3158 , new_n3137 , new_n3157 );
  nand g02782 ( new_n3159 , new_n3158 , new_n3158 );
  nor      g02783 ( new_n3160 , new_n3134 , new_n3159 );
  xor      g02784 ( new_n3161 , new_n3143 , new_n3145 );
  nand g02785 ( new_n3162 , new_n3161 , new_n3161 );
  nand     g02786 ( new_n3163 , new_n3160 , new_n3162 );
  nand g02787 ( new_n3164 , new_n3163 , new_n3163 );
  nand     g02788 ( new_n3165 , new_n3153 , new_n3164 );
  nand     g02789 ( new_n3166 , new_n3152 , new_n3165 );
  xor      g02790 ( new_n3167 , new_n3152 , new_n3165 );
  nand g02791 ( new_n3168 , new_n3167 , new_n3167 );
  xor      g02792 ( new_n3169 , new_n3128 , new_n3149 );
  or       g02793 ( new_n3170 , new_n3168 , new_n3169 );
  nand     g02794 ( new_n3171 , new_n3166 , new_n3170 );
  xnor     g02795 ( new_n3172 , new_n3151 , new_n3171 );
  xor      g02796 ( new_n3173 , new_n3064 , new_n3172 );
  xor      g02797 ( new_n3174 , new_n3168 , new_n3169 );
  xnor     g02798 ( new_n3175 , new_n2958 , new_n2959 );
  nor      g02799 ( new_n3176 , new_n3174 , new_n3175 );
  xor      g02800 ( new_n3177 , new_n3160 , new_n3162 );
  xor      g02801 ( new_n3178 , new_n2913 , new_n2929 );
  nor      g02802 ( new_n3179 , new_n3154 , new_n3178 );
  nand     g02803 ( new_n3180 , pi092 , pi160 );
  nand     g02804 ( new_n3181 , pi020 , pi190 );
  xor      g02805 ( new_n3182 , new_n3180 , new_n3181 );
  nand     g02806 ( new_n3183 , new_n3179 , new_n3182 );
  xor      g02807 ( new_n3184 , new_n3179 , new_n3182 );
  xnor     g02808 ( new_n3185 , new_n2938 , new_n2939 );
  nand     g02809 ( new_n3186 , new_n3184 , new_n3185 );
  nand     g02810 ( new_n3187 , new_n3183 , new_n3186 );
  nand     g02811 ( new_n3188 , new_n3139 , new_n3156 );
  nand     g02812 ( new_n3189 , new_n3159 , new_n3188 );
  nand g02813 ( new_n3190 , new_n3189 , new_n3189 );
  nor      g02814 ( new_n3191 , new_n3187 , new_n3190 );
  xor      g02815 ( new_n3192 , new_n3187 , new_n3189 );
  xor      g02816 ( new_n3193 , new_n2946 , new_n2948 );
  nor      g02817 ( new_n3194 , new_n3192 , new_n3193 );
  nor      g02818 ( new_n3195 , new_n3191 , new_n3194 );
  nand     g02819 ( new_n3196 , new_n3177 , new_n3195 );
  xor      g02820 ( new_n3197 , new_n3177 , new_n3195 );
  xor      g02821 ( new_n3198 , new_n2950 , new_n2951 );
  nand g02822 ( new_n3199 , new_n3198 , new_n3198 );
  nand     g02823 ( new_n3200 , new_n3197 , new_n3199 );
  nand     g02824 ( new_n3201 , new_n3196 , new_n3200 );
  nand g02825 ( new_n3202 , new_n3201 , new_n3201 );
  xor      g02826 ( new_n3203 , new_n3153 , new_n3163 );
  nor      g02827 ( new_n3204 , new_n3202 , new_n3203 );
  xor      g02828 ( new_n3205 , new_n2955 , new_n2956 );
  xor      g02829 ( new_n3206 , new_n3201 , new_n3203 );
  nor      g02830 ( new_n3207 , new_n3205 , new_n3206 );
  nor      g02831 ( new_n3208 , new_n3204 , new_n3207 );
  xnor     g02832 ( new_n3209 , new_n3174 , new_n3175 );
  nor      g02833 ( new_n3210 , new_n3208 , new_n3209 );
  nor      g02834 ( new_n3211 , new_n3176 , new_n3210 );
  xnor     g02835 ( po007 , new_n3173 , new_n3211 );
  nand     g02836 ( new_n3213 , pi029 , pi131 );
  nand     g02837 ( new_n3214 , pi132 , pi168 );
  nand     g02838 ( new_n3215 , pi213 , pi226 );
  nand     g02839 ( new_n3216 , pi109 , pi236 );
  xor      g02840 ( new_n3217 , new_n3215 , new_n3216 );
  xor      g02841 ( new_n3218 , new_n3214 , new_n3217 );
  nor      g02842 ( new_n3219 , new_n3213 , new_n3218 );
  nand g02843 ( new_n3220 , new_n3219 , new_n3219 );
  nand     g02844 ( new_n3221 , pi052 , pi069 );
  nor      g02845 ( new_n3222 , new_n3213 , new_n3221 );
  nand     g02846 ( new_n3223 , pi029 , pi052 );
  nand     g02847 ( new_n3224 , pi069 , pi131 );
  and      g02848 ( new_n3225 , new_n3223 , new_n3224 );
  or       g02849 ( new_n3226 , new_n3222 , new_n3225 );
  nand     g02850 ( new_n3227 , new_n3220 , new_n3226 );
  nand g02851 ( new_n3228 , new_n3214 , new_n3214 );
  nand     g02852 ( new_n3229 , new_n3228 , new_n3217 );
  nand     g02853 ( new_n3230 , pi186 , pi208 );
  nor      g02854 ( new_n3231 , new_n3214 , new_n3230 );
  nand     g02855 ( new_n3232 , pi168 , pi186 );
  nand     g02856 ( new_n3233 , pi132 , pi208 );
  and      g02857 ( new_n3234 , new_n3232 , new_n3233 );
  or       g02858 ( new_n3235 , new_n3231 , new_n3234 );
  xor      g02859 ( new_n3236 , new_n3229 , new_n3235 );
  nor      g02860 ( new_n3237 , new_n3215 , new_n3216 );
  nand     g02861 ( new_n3238 , pi207 , pi212 );
  nor      g02862 ( new_n3239 , new_n3215 , new_n3238 );
  nand     g02863 ( new_n3240 , pi207 , pi213 );
  nand     g02864 ( new_n3241 , pi212 , pi226 );
  and      g02865 ( new_n3242 , new_n3240 , new_n3241 );
  or       g02866 ( new_n3243 , new_n3239 , new_n3242 );
  nand     g02867 ( new_n3244 , pi014 , pi241 );
  or       g02868 ( new_n3245 , new_n3216 , new_n3244 );
  nand     g02869 ( new_n3246 , pi109 , pi241 );
  nand     g02870 ( new_n3247 , pi014 , pi236 );
  nand     g02871 ( new_n3248 , new_n3246 , new_n3247 );
  nand     g02872 ( new_n3249 , new_n3245 , new_n3248 );
  xor      g02873 ( new_n3250 , new_n3243 , new_n3249 );
  xor      g02874 ( new_n3251 , new_n3237 , new_n3250 );
  xnor     g02875 ( new_n3252 , new_n3236 , new_n3251 );
  xor      g02876 ( new_n3253 , new_n3219 , new_n3226 );
  nand g02877 ( new_n3254 , new_n3253 , new_n3253 );
  nand     g02878 ( new_n3255 , new_n3252 , new_n3254 );
  nand     g02879 ( new_n3256 , new_n3227 , new_n3255 );
  nand     g02880 ( new_n3257 , pi029 , pi077 );
  nand     g02881 ( new_n3258 , pi131 , pi244 );
  xor      g02882 ( new_n3259 , new_n3221 , new_n3258 );
  xor      g02883 ( new_n3260 , new_n3257 , new_n3259 );
  xor      g02884 ( new_n3261 , new_n3222 , new_n3260 );
  and      g02885 ( new_n3262 , new_n3256 , new_n3261 );
  xnor     g02886 ( new_n3263 , new_n3256 , new_n3261 );
  nand     g02887 ( new_n3264 , pi104 , pi226 );
  nand     g02888 ( new_n3265 , pi066 , pi213 );
  xor      g02889 ( new_n3266 , new_n3238 , new_n3265 );
  xor      g02890 ( new_n3267 , new_n3264 , new_n3266 );
  xor      g02891 ( new_n3268 , new_n3239 , new_n3267 );
  nand     g02892 ( new_n3269 , new_n3243 , new_n3249 );
  nand g02893 ( new_n3270 , new_n3237 , new_n3237 );
  nand     g02894 ( new_n3271 , new_n3270 , new_n3250 );
  nand     g02895 ( new_n3272 , new_n3269 , new_n3271 );
  xor      g02896 ( new_n3273 , new_n3268 , new_n3272 );
  nand     g02897 ( new_n3274 , pi173 , pi236 );
  nand     g02898 ( new_n3275 , pi109 , pi161 );
  xor      g02899 ( new_n3276 , new_n3274 , new_n3275 );
  nor      g02900 ( new_n3277 , new_n3245 , new_n3276 );
  nor      g02901 ( new_n3278 , new_n3244 , new_n3276 );
  nand     g02902 ( new_n3279 , new_n3244 , new_n3276 );
  nand     g02903 ( new_n3280 , new_n3245 , new_n3279 );
  nor      g02904 ( new_n3281 , new_n3278 , new_n3280 );
  nor      g02905 ( new_n3282 , new_n3277 , new_n3281 );
  nand g02906 ( new_n3283 , new_n3282 , new_n3282 );
  xor      g02907 ( new_n3284 , new_n3273 , new_n3283 );
  nor      g02908 ( new_n3285 , new_n3229 , new_n3235 );
  and      g02909 ( new_n3286 , new_n3236 , new_n3251 );
  nor      g02910 ( new_n3287 , new_n3285 , new_n3286 );
  nand     g02911 ( new_n3288 , pi132 , pi139 );
  nand     g02912 ( new_n3289 , pi058 , pi168 );
  xor      g02913 ( new_n3290 , new_n3230 , new_n3289 );
  xor      g02914 ( new_n3291 , new_n3288 , new_n3290 );
  xor      g02915 ( new_n3292 , new_n3231 , new_n3291 );
  xnor     g02916 ( new_n3293 , new_n3287 , new_n3292 );
  xor      g02917 ( new_n3294 , new_n3284 , new_n3293 );
  nor      g02918 ( new_n3295 , new_n3263 , new_n3294 );
  or       g02919 ( new_n3296 , new_n3262 , new_n3295 );
  nand g02920 ( new_n3297 , new_n3260 , new_n3260 );
  nand     g02921 ( new_n3298 , new_n3222 , new_n3297 );
  nand     g02922 ( new_n3299 , pi029 , pi133 );
  nand     g02923 ( new_n3300 , pi052 , pi244 );
  nand     g02924 ( new_n3301 , pi069 , pi077 );
  xor      g02925 ( new_n3302 , new_n3300 , new_n3301 );
  xor      g02926 ( new_n3303 , new_n3299 , new_n3302 );
  nand     g02927 ( new_n3304 , pi131 , pi150 );
  nand     g02928 ( new_n3305 , new_n3221 , new_n3258 );
  nand     g02929 ( new_n3306 , new_n3257 , new_n3259 );
  nand     g02930 ( new_n3307 , new_n3305 , new_n3306 );
  xor      g02931 ( new_n3308 , new_n3304 , new_n3307 );
  xor      g02932 ( new_n3309 , new_n3303 , new_n3308 );
  xnor     g02933 ( new_n3310 , new_n3298 , new_n3309 );
  xor      g02934 ( new_n3311 , new_n3296 , new_n3310 );
  nor      g02935 ( new_n3312 , new_n3287 , new_n3292 );
  nor      g02936 ( new_n3313 , new_n3284 , new_n3293 );
  nor      g02937 ( new_n3314 , new_n3312 , new_n3313 );
  nand g02938 ( new_n3315 , new_n3291 , new_n3291 );
  nand     g02939 ( new_n3316 , new_n3231 , new_n3315 );
  nand     g02940 ( new_n3317 , pi035 , pi132 );
  nand     g02941 ( new_n3318 , pi058 , pi208 );
  nand     g02942 ( new_n3319 , pi139 , pi186 );
  xor      g02943 ( new_n3320 , new_n3318 , new_n3319 );
  xor      g02944 ( new_n3321 , new_n3317 , new_n3320 );
  nand     g02945 ( new_n3322 , pi168 , pi211 );
  nand     g02946 ( new_n3323 , new_n3230 , new_n3289 );
  nand     g02947 ( new_n3324 , new_n3288 , new_n3290 );
  nand     g02948 ( new_n3325 , new_n3323 , new_n3324 );
  xor      g02949 ( new_n3326 , new_n3322 , new_n3325 );
  nand g02950 ( new_n3327 , new_n3326 , new_n3326 );
  xor      g02951 ( new_n3328 , new_n3321 , new_n3327 );
  xor      g02952 ( new_n3329 , new_n3316 , new_n3328 );
  xor      g02953 ( new_n3330 , new_n3314 , new_n3329 );
  nand     g02954 ( new_n3331 , new_n3268 , new_n3272 );
  nand g02955 ( new_n3332 , new_n3331 , new_n3331 );
  and      g02956 ( new_n3333 , new_n3273 , new_n3283 );
  nor      g02957 ( new_n3334 , new_n3332 , new_n3333 );
  nand     g02958 ( new_n3335 , pi230 , pi236 );
  nand     g02959 ( new_n3336 , new_n3274 , new_n3275 );
  nand     g02960 ( new_n3337 , new_n3336 , new_n3279 );
  xor      g02961 ( new_n3338 , new_n3335 , new_n3337 );
  nand     g02962 ( new_n3339 , pi014 , pi161 );
  nand     g02963 ( new_n3340 , pi109 , pi141 );
  nand     g02964 ( new_n3341 , pi173 , pi241 );
  xor      g02965 ( new_n3342 , new_n3340 , new_n3341 );
  xor      g02966 ( new_n3343 , new_n3339 , new_n3342 );
  nand g02967 ( new_n3344 , new_n3343 , new_n3343 );
  xor      g02968 ( new_n3345 , new_n3338 , new_n3344 );
  xor      g02969 ( new_n3346 , new_n3277 , new_n3345 );
  nand g02970 ( new_n3347 , new_n3346 , new_n3346 );
  nand g02971 ( new_n3348 , new_n3267 , new_n3267 );
  nand     g02972 ( new_n3349 , new_n3239 , new_n3348 );
  nand     g02973 ( new_n3350 , pi066 , pi212 );
  nand     g02974 ( new_n3351 , pi104 , pi207 );
  nand     g02975 ( new_n3352 , pi013 , pi226 );
  xor      g02976 ( new_n3353 , new_n3351 , new_n3352 );
  xor      g02977 ( new_n3354 , new_n3350 , new_n3353 );
  nand     g02978 ( new_n3355 , pi055 , pi213 );
  nand     g02979 ( new_n3356 , new_n3238 , new_n3265 );
  nand     g02980 ( new_n3357 , new_n3264 , new_n3266 );
  nand     g02981 ( new_n3358 , new_n3356 , new_n3357 );
  xor      g02982 ( new_n3359 , new_n3355 , new_n3358 );
  xor      g02983 ( new_n3360 , new_n3354 , new_n3359 );
  xnor     g02984 ( new_n3361 , new_n3349 , new_n3360 );
  nand     g02985 ( new_n3362 , new_n3347 , new_n3361 );
  nand g02986 ( new_n3363 , new_n3362 , new_n3362 );
  nor      g02987 ( new_n3364 , new_n3347 , new_n3361 );
  nor      g02988 ( new_n3365 , new_n3363 , new_n3364 );
  xnor     g02989 ( new_n3366 , new_n3334 , new_n3365 );
  xnor     g02990 ( new_n3367 , new_n3330 , new_n3366 );
  xor      g02991 ( po008 , new_n3311 , new_n3367 );
  nand     g02992 ( new_n3369 , pi065 , pi139 );
  nand     g02993 ( new_n3370 , pi062 , pi208 );
  nand     g02994 ( new_n3371 , pi120 , pi168 );
  xnor     g02995 ( new_n3372 , new_n3370 , new_n3371 );
  xor      g02996 ( new_n3373 , new_n3369 , new_n3372 );
  nand     g02997 ( new_n3374 , pi065 , pi168 );
  nor      g02998 ( new_n3375 , new_n3370 , new_n3374 );
  nand     g02999 ( new_n3376 , new_n3373 , new_n3375 );
  nand     g03000 ( new_n3377 , pi120 , pi208 );
  nand     g03001 ( new_n3378 , pi035 , pi065 );
  nand     g03002 ( new_n3379 , pi062 , pi139 );
  xor      g03003 ( new_n3380 , new_n3378 , new_n3379 );
  xor      g03004 ( new_n3381 , new_n3377 , new_n3380 );
  nand     g03005 ( new_n3382 , pi168 , pi172 );
  nand     g03006 ( new_n3383 , new_n3370 , new_n3371 );
  nand g03007 ( new_n3384 , new_n3372 , new_n3372 );
  nand     g03008 ( new_n3385 , new_n3369 , new_n3384 );
  nand     g03009 ( new_n3386 , new_n3383 , new_n3385 );
  xnor     g03010 ( new_n3387 , new_n3382 , new_n3386 );
  xnor     g03011 ( new_n3388 , new_n3381 , new_n3387 );
  xor      g03012 ( new_n3389 , new_n3376 , new_n3388 );
  nand     g03013 ( new_n3390 , pi104 , pi170 );
  nand     g03014 ( new_n3391 , pi073 , pi213 );
  nor      g03015 ( new_n3392 , new_n3390 , new_n3391 );
  nand     g03016 ( new_n3393 , new_n3390 , new_n3391 );
  nand     g03017 ( new_n3394 , pi004 , pi212 );
  nand g03018 ( new_n3395 , new_n3394 , new_n3394 );
  nand     g03019 ( new_n3396 , pi170 , pi213 );
  and      g03020 ( new_n3397 , new_n3395 , new_n3396 );
  nor      g03021 ( new_n3398 , new_n3393 , new_n3397 );
  nor      g03022 ( new_n3399 , new_n3392 , new_n3398 );
  nand     g03023 ( new_n3400 , new_n3393 , new_n3397 );
  nand     g03024 ( new_n3401 , new_n3399 , new_n3400 );
  nand     g03025 ( new_n3402 , pi161 , pi254 );
  nand     g03026 ( new_n3403 , pi158 , pi241 );
  nand     g03027 ( new_n3404 , pi089 , pi236 );
  xor      g03028 ( new_n3405 , new_n3403 , new_n3404 );
  xor      g03029 ( new_n3406 , new_n3402 , new_n3405 );
  nand     g03030 ( new_n3407 , pi236 , pi254 );
  nor      g03031 ( new_n3408 , new_n3403 , new_n3407 );
  xor      g03032 ( new_n3409 , new_n3406 , new_n3408 );
  or       g03033 ( new_n3410 , new_n3401 , new_n3409 );
  xor      g03034 ( new_n3411 , new_n3401 , new_n3409 );
  nand     g03035 ( new_n3412 , pi158 , pi236 );
  nand     g03036 ( new_n3413 , pi241 , pi254 );
  and      g03037 ( new_n3414 , new_n3412 , new_n3413 );
  nor      g03038 ( new_n3415 , new_n3408 , new_n3414 );
  nand     g03039 ( new_n3416 , pi004 , pi213 );
  nand     g03040 ( new_n3417 , pi170 , pi212 );
  xor      g03041 ( new_n3418 , new_n3416 , new_n3417 );
  nor      g03042 ( new_n3419 , new_n3415 , new_n3418 );
  nor      g03043 ( new_n3420 , new_n3396 , new_n3407 );
  xnor     g03044 ( new_n3421 , new_n3415 , new_n3418 );
  nor      g03045 ( new_n3422 , new_n3420 , new_n3421 );
  nor      g03046 ( new_n3423 , new_n3419 , new_n3422 );
  nand     g03047 ( new_n3424 , new_n3411 , new_n3423 );
  nand     g03048 ( new_n3425 , new_n3410 , new_n3424 );
  nand g03049 ( new_n3426 , new_n3408 , new_n3408 );
  or       g03050 ( new_n3427 , new_n3406 , new_n3426 );
  nand     g03051 ( new_n3428 , pi158 , pi161 );
  nand     g03052 ( new_n3429 , pi089 , pi241 );
  nand     g03053 ( new_n3430 , pi141 , pi254 );
  xor      g03054 ( new_n3431 , new_n3429 , new_n3430 );
  xor      g03055 ( new_n3432 , new_n3428 , new_n3431 );
  nand     g03056 ( new_n3433 , pi154 , pi236 );
  nand     g03057 ( new_n3434 , new_n3403 , new_n3404 );
  nand     g03058 ( new_n3435 , new_n3402 , new_n3405 );
  nand     g03059 ( new_n3436 , new_n3434 , new_n3435 );
  xnor     g03060 ( new_n3437 , new_n3433 , new_n3436 );
  xnor     g03061 ( new_n3438 , new_n3432 , new_n3437 );
  xor      g03062 ( new_n3439 , new_n3427 , new_n3438 );
  nand     g03063 ( new_n3440 , pi013 , pi170 );
  nand     g03064 ( new_n3441 , pi073 , pi212 );
  nand     g03065 ( new_n3442 , pi004 , pi104 );
  xor      g03066 ( new_n3443 , new_n3441 , new_n3442 );
  xor      g03067 ( new_n3444 , new_n3440 , new_n3443 );
  nand     g03068 ( new_n3445 , pi003 , pi213 );
  or       g03069 ( new_n3446 , new_n3392 , new_n3395 );
  nand     g03070 ( new_n3447 , new_n3393 , new_n3446 );
  xnor     g03071 ( new_n3448 , new_n3445 , new_n3447 );
  xor      g03072 ( new_n3449 , new_n3444 , new_n3448 );
  nor      g03073 ( new_n3450 , new_n3394 , new_n3399 );
  xor      g03074 ( new_n3451 , new_n3449 , new_n3450 );
  xor      g03075 ( new_n3452 , new_n3439 , new_n3451 );
  xor      g03076 ( new_n3453 , new_n3425 , new_n3452 );
  xnor     g03077 ( new_n3454 , new_n3389 , new_n3453 );
  xor      g03078 ( new_n3455 , new_n3373 , new_n3375 );
  xor      g03079 ( new_n3456 , new_n3411 , new_n3423 );
  nor      g03080 ( new_n3457 , new_n3455 , new_n3456 );
  nand     g03081 ( new_n3458 , pi062 , pi168 );
  nand     g03082 ( new_n3459 , pi065 , pi208 );
  and      g03083 ( new_n3460 , new_n3458 , new_n3459 );
  or       g03084 ( new_n3461 , new_n3375 , new_n3460 );
  nand g03085 ( new_n3462 , new_n3374 , new_n3374 );
  xor      g03086 ( new_n3463 , new_n3396 , new_n3407 );
  nand     g03087 ( new_n3464 , new_n3462 , new_n3463 );
  nor      g03088 ( new_n3465 , new_n3461 , new_n3464 );
  xnor     g03089 ( new_n3466 , new_n3461 , new_n3464 );
  xor      g03090 ( new_n3467 , new_n3420 , new_n3421 );
  nor      g03091 ( new_n3468 , new_n3466 , new_n3467 );
  or       g03092 ( new_n3469 , new_n3465 , new_n3468 );
  xnor     g03093 ( new_n3470 , new_n3455 , new_n3456 );
  nor      g03094 ( new_n3471 , new_n3469 , new_n3470 );
  nor      g03095 ( new_n3472 , new_n3457 , new_n3471 );
  xor      g03096 ( new_n3473 , new_n3454 , new_n3472 );
  nand     g03097 ( new_n3474 , pi052 , pi229 );
  nand     g03098 ( new_n3475 , pi133 , pi190 );
  nand     g03099 ( new_n3476 , pi077 , pi092 );
  xor      g03100 ( new_n3477 , new_n3475 , new_n3476 );
  xor      g03101 ( new_n3478 , new_n3474 , new_n3477 );
  nand     g03102 ( new_n3479 , pi067 , pi131 );
  nand     g03103 ( new_n3480 , pi131 , pi229 );
  nand     g03104 ( new_n3481 , pi052 , pi092 );
  nand     g03105 ( new_n3482 , new_n3480 , new_n3481 );
  nand     g03106 ( new_n3483 , pi077 , pi190 );
  xor      g03107 ( new_n3484 , new_n3480 , new_n3481 );
  nand     g03108 ( new_n3485 , new_n3483 , new_n3484 );
  nand     g03109 ( new_n3486 , new_n3482 , new_n3485 );
  xor      g03110 ( new_n3487 , new_n3479 , new_n3486 );
  nand g03111 ( new_n3488 , new_n3487 , new_n3487 );
  xor      g03112 ( new_n3489 , new_n3478 , new_n3488 );
  xor      g03113 ( new_n3490 , new_n3483 , new_n3484 );
  nand g03114 ( new_n3491 , new_n3490 , new_n3490 );
  nand     g03115 ( new_n3492 , pi131 , pi190 );
  nor      g03116 ( new_n3493 , new_n3481 , new_n3492 );
  nand     g03117 ( new_n3494 , new_n3491 , new_n3493 );
  xor      g03118 ( new_n3495 , new_n3489 , new_n3494 );
  nand     g03119 ( new_n3496 , new_n3473 , new_n3495 );
  xor      g03120 ( new_n3497 , new_n3374 , new_n3463 );
  nor      g03121 ( new_n3498 , new_n3492 , new_n3497 );
  nand     g03122 ( new_n3499 , pi092 , pi131 );
  nand     g03123 ( new_n3500 , pi052 , pi190 );
  and      g03124 ( new_n3501 , new_n3499 , new_n3500 );
  nor      g03125 ( new_n3502 , new_n3493 , new_n3501 );
  or       g03126 ( new_n3503 , new_n3498 , new_n3502 );
  xnor     g03127 ( new_n3504 , new_n3466 , new_n3467 );
  xor      g03128 ( new_n3505 , new_n3498 , new_n3502 );
  nand     g03129 ( new_n3506 , new_n3504 , new_n3505 );
  nand     g03130 ( new_n3507 , new_n3503 , new_n3506 );
  xor      g03131 ( new_n3508 , new_n3490 , new_n3493 );
  or       g03132 ( new_n3509 , new_n3507 , new_n3508 );
  xor      g03133 ( new_n3510 , new_n3507 , new_n3508 );
  xnor     g03134 ( new_n3511 , new_n3469 , new_n3470 );
  nand     g03135 ( new_n3512 , new_n3510 , new_n3511 );
  nand     g03136 ( new_n3513 , new_n3509 , new_n3512 );
  xnor     g03137 ( new_n3514 , new_n3473 , new_n3495 );
  or       g03138 ( new_n3515 , new_n3513 , new_n3514 );
  nand     g03139 ( new_n3516 , new_n3496 , new_n3515 );
  nand g03140 ( new_n3517 , new_n3494 , new_n3494 );
  nand     g03141 ( new_n3518 , new_n3489 , new_n3517 );
  nand     g03142 ( new_n3519 , pi077 , pi229 );
  nand     g03143 ( new_n3520 , pi189 , pi190 );
  nand     g03144 ( new_n3521 , pi092 , pi133 );
  xor      g03145 ( new_n3522 , new_n3520 , new_n3521 );
  xor      g03146 ( new_n3523 , new_n3519 , new_n3522 );
  nand     g03147 ( new_n3524 , new_n3475 , new_n3476 );
  nand     g03148 ( new_n3525 , new_n3474 , new_n3477 );
  nand     g03149 ( new_n3526 , new_n3524 , new_n3525 );
  nand     g03150 ( new_n3527 , pi052 , pi067 );
  xor      g03151 ( new_n3528 , new_n3526 , new_n3527 );
  xor      g03152 ( new_n3529 , new_n3523 , new_n3528 );
  nand     g03153 ( new_n3530 , pi053 , pi131 );
  nor      g03154 ( new_n3531 , new_n3479 , new_n3486 );
  nor      g03155 ( new_n3532 , new_n3478 , new_n3488 );
  nor      g03156 ( new_n3533 , new_n3531 , new_n3532 );
  xnor     g03157 ( new_n3534 , new_n3530 , new_n3533 );
  xor      g03158 ( new_n3535 , new_n3529 , new_n3534 );
  xor      g03159 ( new_n3536 , new_n3518 , new_n3535 );
  xnor     g03160 ( new_n3537 , new_n3516 , new_n3536 );
  nor      g03161 ( new_n3538 , new_n3376 , new_n3388 );
  nand g03162 ( new_n3539 , new_n3538 , new_n3538 );
  nand     g03163 ( new_n3540 , pi168 , pi198 );
  nor      g03164 ( new_n3541 , new_n3382 , new_n3386 );
  nor      g03165 ( new_n3542 , new_n3381 , new_n3387 );
  nor      g03166 ( new_n3543 , new_n3541 , new_n3542 );
  xnor     g03167 ( new_n3544 , new_n3540 , new_n3543 );
  nand     g03168 ( new_n3545 , pi120 , pi139 );
  nand     g03169 ( new_n3546 , pi035 , pi062 );
  nand     g03170 ( new_n3547 , pi015 , pi065 );
  xor      g03171 ( new_n3548 , new_n3546 , new_n3547 );
  xor      g03172 ( new_n3549 , new_n3545 , new_n3548 );
  nand     g03173 ( new_n3550 , new_n3378 , new_n3379 );
  nand     g03174 ( new_n3551 , new_n3377 , new_n3380 );
  nand     g03175 ( new_n3552 , new_n3550 , new_n3551 );
  nand     g03176 ( new_n3553 , pi172 , pi208 );
  xor      g03177 ( new_n3554 , new_n3552 , new_n3553 );
  xor      g03178 ( new_n3555 , new_n3549 , new_n3554 );
  xnor     g03179 ( new_n3556 , new_n3544 , new_n3555 );
  xor      g03180 ( new_n3557 , new_n3539 , new_n3556 );
  nor      g03181 ( new_n3558 , new_n3389 , new_n3453 );
  nor      g03182 ( new_n3559 , new_n3454 , new_n3472 );
  nor      g03183 ( new_n3560 , new_n3558 , new_n3559 );
  xor      g03184 ( new_n3561 , new_n3557 , new_n3560 );
  nand     g03185 ( new_n3562 , new_n3449 , new_n3450 );
  nand g03186 ( new_n3563 , new_n3562 , new_n3562 );
  nand     g03187 ( new_n3564 , pi073 , pi104 );
  nand     g03188 ( new_n3565 , pi112 , pi170 );
  nand     g03189 ( new_n3566 , pi004 , pi013 );
  xor      g03190 ( new_n3567 , new_n3565 , new_n3566 );
  xor      g03191 ( new_n3568 , new_n3564 , new_n3567 );
  nand     g03192 ( new_n3569 , pi003 , pi212 );
  nand     g03193 ( new_n3570 , new_n3441 , new_n3442 );
  nand     g03194 ( new_n3571 , new_n3440 , new_n3443 );
  nand     g03195 ( new_n3572 , new_n3570 , new_n3571 );
  xor      g03196 ( new_n3573 , new_n3569 , new_n3572 );
  xor      g03197 ( new_n3574 , new_n3568 , new_n3573 );
  nand     g03198 ( new_n3575 , pi130 , pi213 );
  nor      g03199 ( new_n3576 , new_n3445 , new_n3447 );
  nor      g03200 ( new_n3577 , new_n3444 , new_n3448 );
  nor      g03201 ( new_n3578 , new_n3576 , new_n3577 );
  xor      g03202 ( new_n3579 , new_n3575 , new_n3578 );
  xnor     g03203 ( new_n3580 , new_n3574 , new_n3579 );
  xor      g03204 ( new_n3581 , new_n3563 , new_n3580 );
  nand     g03205 ( new_n3582 , new_n3439 , new_n3451 );
  nand     g03206 ( new_n3583 , new_n3425 , new_n3452 );
  nand     g03207 ( new_n3584 , new_n3582 , new_n3583 );
  nor      g03208 ( new_n3585 , new_n3427 , new_n3438 );
  nand     g03209 ( new_n3586 , pi095 , pi236 );
  nor      g03210 ( new_n3587 , new_n3433 , new_n3436 );
  nor      g03211 ( new_n3588 , new_n3432 , new_n3437 );
  nor      g03212 ( new_n3589 , new_n3587 , new_n3588 );
  xor      g03213 ( new_n3590 , new_n3586 , new_n3589 );
  nand     g03214 ( new_n3591 , pi141 , pi158 );
  nand     g03215 ( new_n3592 , pi089 , pi161 );
  nand     g03216 ( new_n3593 , pi090 , pi254 );
  xor      g03217 ( new_n3594 , new_n3592 , new_n3593 );
  xnor     g03218 ( new_n3595 , new_n3591 , new_n3594 );
  and      g03219 ( new_n3596 , new_n3429 , new_n3430 );
  and      g03220 ( new_n3597 , new_n3428 , new_n3431 );
  or       g03221 ( new_n3598 , new_n3596 , new_n3597 );
  nand     g03222 ( new_n3599 , pi154 , pi241 );
  xnor     g03223 ( new_n3600 , new_n3598 , new_n3599 );
  xnor     g03224 ( new_n3601 , new_n3595 , new_n3600 );
  xor      g03225 ( new_n3602 , new_n3590 , new_n3601 );
  xor      g03226 ( new_n3603 , new_n3585 , new_n3602 );
  xnor     g03227 ( new_n3604 , new_n3584 , new_n3603 );
  xnor     g03228 ( new_n3605 , new_n3581 , new_n3604 );
  xor      g03229 ( new_n3606 , new_n3561 , new_n3605 );
  xnor     g03230 ( po009 , new_n3537 , new_n3606 );
  nand     g03231 ( new_n3608 , pi162 , pi168 );
  nand     g03232 ( new_n3609 , pi051 , pi236 );
  nand     g03233 ( new_n3610 , pi188 , pi213 );
  xnor     g03234 ( new_n3611 , new_n3609 , new_n3610 );
  xor      g03235 ( new_n3612 , new_n3608 , new_n3611 );
  nand g03236 ( new_n3613 , new_n3612 , new_n3612 );
  nand     g03237 ( new_n3614 , pi131 , pi143 );
  xor      g03238 ( po010 , new_n3613 , new_n3614 );
  xnor     g03239 ( po011 , new_n1886 , new_n1893 );
  xnor     g03240 ( po012 , new_n3513 , new_n3514 );
  nand     g03241 ( new_n3618 , pi155 , pi207 );
  nand     g03242 ( new_n3619 , pi132 , pi192 );
  xor      g03243 ( new_n3620 , new_n3618 , new_n3619 );
  nand     g03244 ( new_n3621 , pi029 , pi137 );
  nand     g03245 ( new_n3622 , pi087 , pi205 );
  nand     g03246 ( new_n3623 , pi001 , pi050 );
  xor      g03247 ( new_n3624 , new_n3622 , new_n3623 );
  nand     g03248 ( new_n3625 , pi025 , pi169 );
  nand     g03249 ( new_n3626 , pi074 , pi087 );
  nand     g03250 ( new_n3627 , pi219 , pi253 );
  nand     g03251 ( new_n3628 , new_n3626 , new_n3627 );
  nand     g03252 ( new_n3629 , pi050 , pi102 );
  xor      g03253 ( new_n3630 , new_n3626 , new_n3627 );
  nand     g03254 ( new_n3631 , new_n3629 , new_n3630 );
  nand     g03255 ( new_n3632 , new_n3628 , new_n3631 );
  nand     g03256 ( new_n3633 , pi066 , pi123 );
  nand     g03257 ( new_n3634 , pi023 , pi226 );
  nand     g03258 ( new_n3635 , pi099 , pi207 );
  nand     g03259 ( new_n3636 , new_n3634 , new_n3635 );
  nand     g03260 ( new_n3637 , pi099 , pi226 );
  nand     g03261 ( new_n3638 , pi023 , pi207 );
  nor      g03262 ( new_n3639 , new_n3637 , new_n3638 );
  nand g03263 ( new_n3640 , new_n3639 , new_n3639 );
  nand     g03264 ( new_n3641 , new_n3636 , new_n3640 );
  nand     g03265 ( new_n3642 , new_n3633 , new_n3641 );
  nand     g03266 ( new_n3643 , pi066 , pi169 );
  nand     g03267 ( new_n3644 , new_n3637 , new_n3643 );
  nand     g03268 ( new_n3645 , pi123 , pi207 );
  xor      g03269 ( new_n3646 , new_n3637 , new_n3643 );
  nand     g03270 ( new_n3647 , new_n3645 , new_n3646 );
  nand     g03271 ( new_n3648 , new_n3644 , new_n3647 );
  xor      g03272 ( new_n3649 , new_n3633 , new_n3641 );
  nand     g03273 ( new_n3650 , new_n3648 , new_n3649 );
  nand     g03274 ( new_n3651 , new_n3642 , new_n3650 );
  nand     g03275 ( new_n3652 , pi025 , pi071 );
  nand     g03276 ( new_n3653 , pi142 , pi239 );
  xor      g03277 ( new_n3654 , new_n3652 , new_n3653 );
  nand     g03278 ( new_n3655 , pi002 , pi169 );
  xor      g03279 ( new_n3656 , new_n3654 , new_n3655 );
  nand     g03280 ( new_n3657 , new_n3651 , new_n3656 );
  nand     g03281 ( new_n3658 , pi055 , pi123 );
  xor      g03282 ( new_n3659 , new_n3639 , new_n3658 );
  nand     g03283 ( new_n3660 , pi066 , pi099 );
  nand     g03284 ( new_n3661 , pi155 , pi226 );
  xor      g03285 ( new_n3662 , new_n3638 , new_n3661 );
  xor      g03286 ( new_n3663 , new_n3660 , new_n3662 );
  xnor     g03287 ( new_n3664 , new_n3659 , new_n3663 );
  xnor     g03288 ( new_n3665 , new_n3651 , new_n3656 );
  nand g03289 ( new_n3666 , new_n3665 , new_n3665 );
  nand     g03290 ( new_n3667 , new_n3664 , new_n3666 );
  nand     g03291 ( new_n3668 , new_n3657 , new_n3667 );
  xor      g03292 ( new_n3669 , new_n3632 , new_n3668 );
  xor      g03293 ( new_n3670 , new_n3625 , new_n3669 );
  xor      g03294 ( new_n3671 , new_n3624 , new_n3670 );
  xor      g03295 ( new_n3672 , new_n3621 , new_n3671 );
  xor      g03296 ( new_n3673 , new_n3620 , new_n3672 );
  nand     g03297 ( new_n3674 , pi041 , pi195 );
  nand     g03298 ( new_n3675 , pi060 , pi221 );
  nand     g03299 ( new_n3676 , pi020 , pi196 );
  nand     g03300 ( new_n3677 , pi160 , pi184 );
  xor      g03301 ( new_n3678 , new_n3676 , new_n3677 );
  xor      g03302 ( new_n3679 , new_n3675 , new_n3678 );
  nand     g03303 ( new_n3680 , pi223 , pi244 );
  nand     g03304 ( new_n3681 , pi069 , pi101 );
  nand     g03305 ( new_n3682 , pi029 , pi225 );
  nand     g03306 ( new_n3683 , new_n3681 , new_n3682 );
  nand     g03307 ( new_n3684 , pi029 , pi101 );
  nand g03308 ( new_n3685 , new_n3684 , new_n3684 );
  nand     g03309 ( new_n3686 , pi069 , pi225 );
  nand g03310 ( new_n3687 , new_n3686 , new_n3686 );
  nand     g03311 ( new_n3688 , new_n3685 , new_n3687 );
  nand     g03312 ( new_n3689 , new_n3683 , new_n3688 );
  nand     g03313 ( new_n3690 , new_n3680 , new_n3689 );
  nand     g03314 ( new_n3691 , pi069 , pi223 );
  nand     g03315 ( new_n3692 , new_n3684 , new_n3691 );
  nand     g03316 ( new_n3693 , pi060 , pi244 );
  xor      g03317 ( new_n3694 , new_n3685 , new_n3691 );
  nand g03318 ( new_n3695 , new_n3694 , new_n3694 );
  nand     g03319 ( new_n3696 , new_n3693 , new_n3695 );
  nand     g03320 ( new_n3697 , new_n3692 , new_n3696 );
  xor      g03321 ( new_n3698 , new_n3680 , new_n3689 );
  nand     g03322 ( new_n3699 , new_n3697 , new_n3698 );
  nand     g03323 ( new_n3700 , new_n3690 , new_n3699 );
  nand     g03324 ( new_n3701 , new_n3679 , new_n3700 );
  xor      g03325 ( new_n3702 , new_n3679 , new_n3700 );
  nand     g03326 ( new_n3703 , pi150 , pi223 );
  xor      g03327 ( new_n3704 , new_n3688 , new_n3703 );
  nand     g03328 ( new_n3705 , pi029 , pi177 );
  and      g03329 ( new_n3706 , pi101 , pi244 );
  xor      g03330 ( new_n3707 , new_n3705 , new_n3706 );
  xor      g03331 ( new_n3708 , new_n3686 , new_n3707 );
  xnor     g03332 ( new_n3709 , new_n3704 , new_n3708 );
  nand     g03333 ( new_n3710 , new_n3702 , new_n3709 );
  nand     g03334 ( new_n3711 , new_n3701 , new_n3710 );
  xor      g03335 ( new_n3712 , new_n3674 , new_n3711 );
  nand     g03336 ( new_n3713 , pi058 , pi216 );
  nand     g03337 ( new_n3714 , pi076 , pi132 );
  nand g03338 ( new_n3715 , new_n3714 , new_n3714 );
  nand     g03339 ( new_n3716 , pi079 , pi186 );
  nand g03340 ( new_n3717 , new_n3716 , new_n3716 );
  nand     g03341 ( new_n3718 , new_n3715 , new_n3717 );
  nand     g03342 ( new_n3719 , pi079 , pi132 );
  nand     g03343 ( new_n3720 , pi076 , pi186 );
  nand     g03344 ( new_n3721 , new_n3719 , new_n3720 );
  nand     g03345 ( new_n3722 , new_n3718 , new_n3721 );
  nand     g03346 ( new_n3723 , new_n3713 , new_n3722 );
  nand     g03347 ( new_n3724 , pi186 , pi216 );
  nand     g03348 ( new_n3725 , pi041 , pi058 );
  nand     g03349 ( new_n3726 , new_n3724 , new_n3725 );
  xor      g03350 ( new_n3727 , new_n3724 , new_n3725 );
  nand     g03351 ( new_n3728 , new_n3714 , new_n3727 );
  nand     g03352 ( new_n3729 , new_n3726 , new_n3728 );
  xor      g03353 ( new_n3730 , new_n3713 , new_n3722 );
  nand     g03354 ( new_n3731 , new_n3729 , new_n3730 );
  nand     g03355 ( new_n3732 , new_n3723 , new_n3731 );
  nand     g03356 ( new_n3733 , pi041 , pi199 );
  nand     g03357 ( new_n3734 , pi138 , pi218 );
  nand     g03358 ( new_n3735 , pi182 , pi195 );
  xor      g03359 ( new_n3736 , new_n3734 , new_n3735 );
  xor      g03360 ( new_n3737 , new_n3733 , new_n3736 );
  or       g03361 ( new_n3738 , new_n3732 , new_n3737 );
  nand     g03362 ( new_n3739 , pi211 , pi216 );
  xor      g03363 ( new_n3740 , new_n3718 , new_n3739 );
  nand     g03364 ( new_n3741 , pi132 , pi251 );
  nand     g03365 ( new_n3742 , pi058 , pi076 );
  xor      g03366 ( new_n3743 , new_n3717 , new_n3742 );
  xor      g03367 ( new_n3744 , new_n3741 , new_n3743 );
  xor      g03368 ( new_n3745 , new_n3740 , new_n3744 );
  xor      g03369 ( new_n3746 , new_n3732 , new_n3737 );
  nand     g03370 ( new_n3747 , new_n3745 , new_n3746 );
  nand     g03371 ( new_n3748 , new_n3738 , new_n3747 );
  xor      g03372 ( new_n3749 , new_n3712 , new_n3748 );
  nand     g03373 ( new_n3750 , pi225 , pi244 );
  nand     g03374 ( new_n3751 , pi086 , pi226 );
  xor      g03375 ( new_n3752 , new_n3750 , new_n3751 );
  nand     g03376 ( new_n3753 , pi102 , pi253 );
  nand     g03377 ( new_n3754 , pi002 , pi142 );
  nand     g03378 ( new_n3755 , pi055 , pi142 );
  nand     g03379 ( new_n3756 , pi071 , pi207 );
  nand     g03380 ( new_n3757 , pi066 , pi142 );
  nand     g03381 ( new_n3758 , new_n3756 , new_n3757 );
  nand     g03382 ( new_n3759 , pi169 , pi226 );
  xor      g03383 ( new_n3760 , new_n3756 , new_n3757 );
  nand     g03384 ( new_n3761 , new_n3759 , new_n3760 );
  nand     g03385 ( new_n3762 , new_n3758 , new_n3761 );
  nor      g03386 ( new_n3763 , new_n3755 , new_n3762 );
  nand     g03387 ( new_n3764 , pi066 , pi071 );
  nand     g03388 ( new_n3765 , pi123 , pi226 );
  xor      g03389 ( new_n3766 , new_n3764 , new_n3765 );
  nand     g03390 ( new_n3767 , pi169 , pi207 );
  xor      g03391 ( new_n3768 , new_n3766 , new_n3767 );
  xnor     g03392 ( new_n3769 , new_n3755 , new_n3762 );
  nor      g03393 ( new_n3770 , new_n3768 , new_n3769 );
  nor      g03394 ( new_n3771 , new_n3763 , new_n3770 );
  nor      g03395 ( new_n3772 , new_n3754 , new_n3771 );
  xor      g03396 ( new_n3773 , new_n3754 , new_n3771 );
  xor      g03397 ( new_n3774 , new_n3645 , new_n3646 );
  nand     g03398 ( new_n3775 , new_n3764 , new_n3765 );
  nand     g03399 ( new_n3776 , new_n3766 , new_n3767 );
  nand     g03400 ( new_n3777 , new_n3775 , new_n3776 );
  nand     g03401 ( new_n3778 , pi055 , pi071 );
  xor      g03402 ( new_n3779 , new_n3777 , new_n3778 );
  xnor     g03403 ( new_n3780 , new_n3774 , new_n3779 );
  and      g03404 ( new_n3781 , new_n3773 , new_n3780 );
  nor      g03405 ( new_n3782 , new_n3772 , new_n3781 );
  xor      g03406 ( new_n3783 , new_n3648 , new_n3649 );
  nand g03407 ( new_n3784 , new_n3783 , new_n3783 );
  nand     g03408 ( new_n3785 , new_n3777 , new_n3778 );
  nand     g03409 ( new_n3786 , new_n3774 , new_n3779 );
  nand     g03410 ( new_n3787 , new_n3785 , new_n3786 );
  nand     g03411 ( new_n3788 , pi002 , pi071 );
  nand     g03412 ( new_n3789 , pi055 , pi169 );
  and      g03413 ( new_n3790 , new_n3788 , new_n3789 );
  nor      g03414 ( new_n3791 , new_n3655 , new_n3778 );
  nor      g03415 ( new_n3792 , new_n3790 , new_n3791 );
  xor      g03416 ( new_n3793 , new_n3787 , new_n3792 );
  xor      g03417 ( new_n3794 , new_n3784 , new_n3793 );
  or       g03418 ( new_n3795 , new_n3782 , new_n3794 );
  xor      g03419 ( new_n3796 , new_n3664 , new_n3665 );
  nand g03420 ( new_n3797 , new_n3792 , new_n3792 );
  nand     g03421 ( new_n3798 , new_n3787 , new_n3797 );
  or       g03422 ( new_n3799 , new_n3784 , new_n3793 );
  nand     g03423 ( new_n3800 , new_n3798 , new_n3799 );
  xor      g03424 ( new_n3801 , new_n3791 , new_n3800 );
  xor      g03425 ( new_n3802 , new_n3796 , new_n3801 );
  or       g03426 ( new_n3803 , new_n3795 , new_n3802 );
  nand     g03427 ( new_n3804 , pi025 , pi142 );
  xnor     g03428 ( new_n3805 , new_n3782 , new_n3794 );
  or       g03429 ( new_n3806 , new_n3804 , new_n3805 );
  xnor     g03430 ( new_n3807 , new_n3759 , new_n3760 );
  nand     g03431 ( new_n3808 , pi142 , pi207 );
  nand     g03432 ( new_n3809 , pi071 , pi226 );
  nor      g03433 ( new_n3810 , new_n3808 , new_n3809 );
  and      g03434 ( new_n3811 , new_n3807 , new_n3810 );
  nand g03435 ( new_n3812 , new_n3811 , new_n3811 );
  xnor     g03436 ( new_n3813 , new_n3768 , new_n3769 );
  nor      g03437 ( new_n3814 , new_n3812 , new_n3813 );
  xor      g03438 ( new_n3815 , new_n3773 , new_n3780 );
  and      g03439 ( new_n3816 , new_n3814 , new_n3815 );
  xor      g03440 ( new_n3817 , new_n3804 , new_n3805 );
  nand     g03441 ( new_n3818 , new_n3816 , new_n3817 );
  nand     g03442 ( new_n3819 , new_n3806 , new_n3818 );
  xor      g03443 ( new_n3820 , new_n3795 , new_n3802 );
  nand     g03444 ( new_n3821 , new_n3819 , new_n3820 );
  nand     g03445 ( new_n3822 , new_n3803 , new_n3821 );
  nand     g03446 ( new_n3823 , pi023 , pi066 );
  xor      g03447 ( new_n3824 , new_n3822 , new_n3823 );
  xor      g03448 ( new_n3825 , new_n3753 , new_n3824 );
  nand     g03449 ( new_n3826 , new_n3716 , new_n3742 );
  nand g03450 ( new_n3827 , new_n3743 , new_n3743 );
  nand     g03451 ( new_n3828 , new_n3741 , new_n3827 );
  nand     g03452 ( new_n3829 , new_n3826 , new_n3828 );
  nand     g03453 ( new_n3830 , pi094 , pi109 );
  xor      g03454 ( new_n3831 , new_n3829 , new_n3830 );
  nand     g03455 ( new_n3832 , pi138 , pi199 );
  nand     g03456 ( new_n3833 , pi138 , pi211 );
  nand     g03457 ( new_n3834 , pi058 , pi138 );
  nand     g03458 ( new_n3835 , pi182 , pi186 );
  nand     g03459 ( new_n3836 , new_n3834 , new_n3835 );
  nand     g03460 ( new_n3837 , pi041 , pi132 );
  xor      g03461 ( new_n3838 , new_n3834 , new_n3835 );
  nand     g03462 ( new_n3839 , new_n3837 , new_n3838 );
  nand     g03463 ( new_n3840 , new_n3836 , new_n3839 );
  nor      g03464 ( new_n3841 , new_n3833 , new_n3840 );
  xnor     g03465 ( new_n3842 , new_n3833 , new_n3840 );
  nand     g03466 ( new_n3843 , pi058 , pi182 );
  nand     g03467 ( new_n3844 , pi041 , pi186 );
  nand     g03468 ( new_n3845 , pi132 , pi216 );
  xor      g03469 ( new_n3846 , new_n3844 , new_n3845 );
  xor      g03470 ( new_n3847 , new_n3843 , new_n3846 );
  nor      g03471 ( new_n3848 , new_n3842 , new_n3847 );
  nor      g03472 ( new_n3849 , new_n3841 , new_n3848 );
  nor      g03473 ( new_n3850 , new_n3832 , new_n3849 );
  xor      g03474 ( new_n3851 , new_n3832 , new_n3849 );
  xor      g03475 ( new_n3852 , new_n3715 , new_n3727 );
  nand     g03476 ( new_n3853 , pi182 , pi211 );
  nand     g03477 ( new_n3854 , new_n3844 , new_n3845 );
  nand     g03478 ( new_n3855 , new_n3843 , new_n3846 );
  nand     g03479 ( new_n3856 , new_n3854 , new_n3855 );
  xnor     g03480 ( new_n3857 , new_n3853 , new_n3856 );
  xnor     g03481 ( new_n3858 , new_n3852 , new_n3857 );
  and      g03482 ( new_n3859 , new_n3851 , new_n3858 );
  nor      g03483 ( new_n3860 , new_n3850 , new_n3859 );
  nand     g03484 ( new_n3861 , new_n3853 , new_n3856 );
  or       g03485 ( new_n3862 , new_n3852 , new_n3857 );
  nand     g03486 ( new_n3863 , new_n3861 , new_n3862 );
  nand     g03487 ( new_n3864 , pi041 , pi211 );
  nand     g03488 ( new_n3865 , pi182 , pi199 );
  nand     g03489 ( new_n3866 , new_n3864 , new_n3865 );
  nor      g03490 ( new_n3867 , new_n3733 , new_n3853 );
  nand g03491 ( new_n3868 , new_n3867 , new_n3867 );
  nand     g03492 ( new_n3869 , new_n3866 , new_n3868 );
  xor      g03493 ( new_n3870 , new_n3729 , new_n3730 );
  xnor     g03494 ( new_n3871 , new_n3869 , new_n3870 );
  xor      g03495 ( new_n3872 , new_n3863 , new_n3871 );
  nand g03496 ( new_n3873 , new_n3872 , new_n3872 );
  or       g03497 ( new_n3874 , new_n3860 , new_n3873 );
  nor      g03498 ( new_n3875 , new_n3863 , new_n3871 );
  nand     g03499 ( new_n3876 , new_n3867 , new_n3875 );
  or       g03500 ( new_n3877 , new_n3863 , new_n3871 );
  nor      g03501 ( new_n3878 , new_n3869 , new_n3870 );
  nor      g03502 ( new_n3879 , new_n3867 , new_n3878 );
  nand     g03503 ( new_n3880 , new_n3877 , new_n3879 );
  nand     g03504 ( new_n3881 , new_n3876 , new_n3880 );
  xor      g03505 ( new_n3882 , new_n3745 , new_n3746 );
  xor      g03506 ( new_n3883 , new_n3881 , new_n3882 );
  nor      g03507 ( new_n3884 , new_n3874 , new_n3883 );
  xnor     g03508 ( new_n3885 , new_n3874 , new_n3883 );
  nand     g03509 ( new_n3886 , pi138 , pi195 );
  xor      g03510 ( new_n3887 , new_n3860 , new_n3872 );
  nor      g03511 ( new_n3888 , new_n3886 , new_n3887 );
  xor      g03512 ( new_n3889 , new_n3837 , new_n3838 );
  nand     g03513 ( new_n3890 , pi132 , pi138 );
  or       g03514 ( new_n3891 , new_n3835 , new_n3890 );
  or       g03515 ( new_n3892 , new_n3889 , new_n3891 );
  xnor     g03516 ( new_n3893 , new_n3842 , new_n3847 );
  nor      g03517 ( new_n3894 , new_n3892 , new_n3893 );
  xor      g03518 ( new_n3895 , new_n3851 , new_n3858 );
  nand     g03519 ( new_n3896 , new_n3894 , new_n3895 );
  xnor     g03520 ( new_n3897 , new_n3886 , new_n3887 );
  nor      g03521 ( new_n3898 , new_n3896 , new_n3897 );
  nor      g03522 ( new_n3899 , new_n3888 , new_n3898 );
  nor      g03523 ( new_n3900 , new_n3885 , new_n3899 );
  nor      g03524 ( new_n3901 , new_n3884 , new_n3900 );
  nand     g03525 ( new_n3902 , pi199 , pi216 );
  nand     g03526 ( new_n3903 , pi142 , pi243 );
  xor      g03527 ( new_n3904 , new_n3902 , new_n3903 );
  nand g03528 ( new_n3905 , new_n3705 , new_n3705 );
  nor      g03529 ( new_n3906 , new_n3905 , new_n3706 );
  nor      g03530 ( new_n3907 , new_n3687 , new_n3707 );
  nor      g03531 ( new_n3908 , new_n3906 , new_n3907 );
  xor      g03532 ( new_n3909 , new_n3904 , new_n3908 );
  xor      g03533 ( new_n3910 , new_n3901 , new_n3909 );
  xor      g03534 ( new_n3911 , new_n3831 , new_n3910 );
  xor      g03535 ( new_n3912 , new_n3825 , new_n3911 );
  xor      g03536 ( new_n3913 , new_n3752 , new_n3912 );
  xor      g03537 ( new_n3914 , new_n3749 , new_n3913 );
  nand     g03538 ( new_n3915 , pi058 , pi079 );
  nand g03539 ( new_n3916 , pi014 , pi014 );
  nand g03540 ( new_n3917 , pi059 , pi059 );
  nor      g03541 ( new_n3918 , new_n3916 , new_n3917 );
  xor      g03542 ( new_n3919 , new_n3915 , new_n3918 );
  nand     g03543 ( new_n3920 , pi076 , pi211 );
  xor      g03544 ( new_n3921 , new_n3919 , new_n3920 );
  nand     g03545 ( new_n3922 , pi069 , pi177 );
  or       g03546 ( new_n3923 , new_n3688 , new_n3703 );
  nand     g03547 ( new_n3924 , new_n3704 , new_n3708 );
  nand     g03548 ( new_n3925 , new_n3923 , new_n3924 );
  xor      g03549 ( new_n3926 , new_n3922 , new_n3925 );
  xor      g03550 ( new_n3927 , new_n3921 , new_n3926 );
  xor      g03551 ( new_n3928 , new_n3914 , new_n3927 );
  nand     g03552 ( new_n3929 , pi182 , pi218 );
  nand g03553 ( new_n3930 , new_n3800 , new_n3800 );
  nor      g03554 ( new_n3931 , new_n3791 , new_n3930 );
  nor      g03555 ( new_n3932 , new_n3796 , new_n3801 );
  nor      g03556 ( new_n3933 , new_n3931 , new_n3932 );
  xor      g03557 ( new_n3934 , new_n3929 , new_n3933 );
  nand     g03558 ( new_n3935 , pi060 , pi196 );
  nand     g03559 ( new_n3936 , new_n3734 , new_n3735 );
  nand     g03560 ( new_n3937 , new_n3733 , new_n3736 );
  nand     g03561 ( new_n3938 , new_n3936 , new_n3937 );
  nand     g03562 ( new_n3939 , pi101 , pi150 );
  nor      g03563 ( new_n3940 , new_n3718 , new_n3739 );
  and      g03564 ( new_n3941 , new_n3740 , new_n3744 );
  nor      g03565 ( new_n3942 , new_n3940 , new_n3941 );
  xnor     g03566 ( new_n3943 , new_n3939 , new_n3942 );
  xor      g03567 ( new_n3944 , new_n3938 , new_n3943 );
  xor      g03568 ( new_n3945 , new_n3935 , new_n3944 );
  nand     g03569 ( new_n3946 , pi037 , pi138 );
  nand     g03570 ( new_n3947 , pi087 , pi253 );
  nand     g03571 ( new_n3948 , pi014 , pi219 );
  nand g03572 ( new_n3949 , new_n3948 , new_n3948 );
  nand     g03573 ( new_n3950 , pi087 , pi109 );
  nand     g03574 ( new_n3951 , new_n3949 , new_n3950 );
  nand g03575 ( new_n3952 , new_n3951 , new_n3951 );
  nand     g03576 ( new_n3953 , pi087 , pi173 );
  nand     g03577 ( new_n3954 , pi102 , pi109 );
  nor      g03578 ( new_n3955 , new_n3953 , new_n3954 );
  and      g03579 ( new_n3956 , new_n3953 , new_n3954 );
  nor      g03580 ( new_n3957 , new_n3955 , new_n3956 );
  nor      g03581 ( new_n3958 , new_n3952 , new_n3957 );
  and      g03582 ( new_n3959 , new_n3949 , new_n3958 );
  nand     g03583 ( new_n3960 , pi001 , pi109 );
  nand     g03584 ( new_n3961 , pi173 , pi219 );
  nand     g03585 ( new_n3962 , pi014 , pi102 );
  xor      g03586 ( new_n3963 , new_n3961 , new_n3962 );
  xor      g03587 ( new_n3964 , new_n3960 , new_n3963 );
  nor      g03588 ( new_n3965 , new_n3949 , new_n3955 );
  or       g03589 ( new_n3966 , new_n3956 , new_n3965 );
  nand     g03590 ( new_n3967 , pi087 , pi230 );
  xnor     g03591 ( new_n3968 , new_n3966 , new_n3967 );
  xor      g03592 ( new_n3969 , new_n3964 , new_n3968 );
  nand     g03593 ( new_n3970 , new_n3959 , new_n3969 );
  nand     g03594 ( new_n3971 , pi050 , pi087 );
  nor      g03595 ( new_n3972 , new_n3966 , new_n3967 );
  nor      g03596 ( new_n3973 , new_n3964 , new_n3968 );
  nor      g03597 ( new_n3974 , new_n3972 , new_n3973 );
  xor      g03598 ( new_n3975 , new_n3971 , new_n3974 );
  nand     g03599 ( new_n3976 , pi102 , pi173 );
  nand     g03600 ( new_n3977 , pi109 , pi122 );
  nand     g03601 ( new_n3978 , pi001 , pi014 );
  xor      g03602 ( new_n3979 , new_n3977 , new_n3978 );
  xor      g03603 ( new_n3980 , new_n3976 , new_n3979 );
  nand     g03604 ( new_n3981 , new_n3961 , new_n3962 );
  nand     g03605 ( new_n3982 , new_n3960 , new_n3963 );
  nand     g03606 ( new_n3983 , new_n3981 , new_n3982 );
  nand     g03607 ( new_n3984 , pi219 , pi230 );
  xnor     g03608 ( new_n3985 , new_n3983 , new_n3984 );
  xor      g03609 ( new_n3986 , new_n3980 , new_n3985 );
  xnor     g03610 ( new_n3987 , new_n3975 , new_n3986 );
  or       g03611 ( new_n3988 , new_n3970 , new_n3987 );
  nand     g03612 ( new_n3989 , new_n3947 , new_n3988 );
  xor      g03613 ( new_n3990 , new_n3947 , new_n3988 );
  or       g03614 ( new_n3991 , new_n3971 , new_n3974 );
  nand     g03615 ( new_n3992 , new_n3975 , new_n3986 );
  and      g03616 ( new_n3993 , new_n3991 , new_n3992 );
  nand     g03617 ( new_n3994 , new_n3983 , new_n3984 );
  nand g03618 ( new_n3995 , new_n3980 , new_n3980 );
  or       g03619 ( new_n3996 , new_n3995 , new_n3985 );
  nand     g03620 ( new_n3997 , new_n3994 , new_n3996 );
  nand     g03621 ( new_n3998 , pi102 , pi230 );
  nand     g03622 ( new_n3999 , pi050 , pi219 );
  and      g03623 ( new_n4000 , new_n3998 , new_n3999 );
  nor      g03624 ( new_n4001 , new_n3629 , new_n3984 );
  or       g03625 ( new_n4002 , new_n4000 , new_n4001 );
  nand g03626 ( new_n4003 , new_n3977 , new_n3977 );
  nand     g03627 ( new_n4004 , pi014 , pi135 );
  nand g03628 ( new_n4005 , new_n4004 , new_n4004 );
  nand     g03629 ( new_n4006 , new_n4003 , new_n4005 );
  nand     g03630 ( new_n4007 , pi014 , pi122 );
  nand     g03631 ( new_n4008 , pi109 , pi135 );
  nand     g03632 ( new_n4009 , new_n4007 , new_n4008 );
  nand     g03633 ( new_n4010 , new_n4006 , new_n4009 );
  nand     g03634 ( new_n4011 , pi001 , pi173 );
  nand     g03635 ( new_n4012 , new_n3977 , new_n3978 );
  nand     g03636 ( new_n4013 , new_n3976 , new_n3979 );
  nand     g03637 ( new_n4014 , new_n4012 , new_n4013 );
  xor      g03638 ( new_n4015 , new_n4011 , new_n4014 );
  xor      g03639 ( new_n4016 , new_n4010 , new_n4015 );
  xnor     g03640 ( new_n4017 , new_n4002 , new_n4016 );
  xnor     g03641 ( new_n4018 , new_n3997 , new_n4017 );
  xnor     g03642 ( new_n4019 , new_n3993 , new_n4018 );
  nand     g03643 ( new_n4020 , new_n3990 , new_n4019 );
  nand     g03644 ( new_n4021 , new_n3989 , new_n4020 );
  nor      g03645 ( new_n4022 , new_n3993 , new_n4018 );
  nor      g03646 ( new_n4023 , new_n4002 , new_n4016 );
  nor      g03647 ( new_n4024 , new_n3997 , new_n4017 );
  xor      g03648 ( new_n4025 , new_n4001 , new_n4024 );
  nor      g03649 ( new_n4026 , new_n4023 , new_n4025 );
  nand     g03650 ( new_n4027 , new_n4011 , new_n4014 );
  nand     g03651 ( new_n4028 , new_n4010 , new_n4015 );
  nand     g03652 ( new_n4029 , new_n4027 , new_n4028 );
  xor      g03653 ( new_n4030 , new_n3629 , new_n3630 );
  xor      g03654 ( new_n4031 , new_n4029 , new_n4030 );
  nand     g03655 ( new_n4032 , pi122 , pi173 );
  nand g03656 ( new_n4033 , pi109 , pi109 );
  nor      g03657 ( new_n4034 , new_n3917 , new_n4033 );
  xor      g03658 ( new_n4035 , new_n4032 , new_n4034 );
  xor      g03659 ( new_n4036 , new_n4005 , new_n4035 );
  nand     g03660 ( new_n4037 , pi001 , pi230 );
  xnor     g03661 ( new_n4038 , new_n4006 , new_n4037 );
  xor      g03662 ( new_n4039 , new_n4036 , new_n4038 );
  xnor     g03663 ( new_n4040 , new_n4031 , new_n4039 );
  xor      g03664 ( new_n4041 , new_n4026 , new_n4040 );
  xnor     g03665 ( new_n4042 , new_n4022 , new_n4041 );
  xnor     g03666 ( new_n4043 , new_n4021 , new_n4042 );
  xnor     g03667 ( new_n4044 , new_n3819 , new_n3820 );
  nor      g03668 ( new_n4045 , new_n4043 , new_n4044 );
  xnor     g03669 ( new_n4046 , new_n3816 , new_n3817 );
  nand g03670 ( new_n4047 , new_n4046 , new_n4046 );
  xnor     g03671 ( new_n4048 , new_n3990 , new_n4019 );
  and      g03672 ( new_n4049 , new_n4047 , new_n4048 );
  nand     g03673 ( new_n4050 , pi142 , pi226 );
  nor      g03674 ( new_n4051 , new_n3950 , new_n4050 );
  xor      g03675 ( new_n4052 , new_n3808 , new_n3809 );
  nor      g03676 ( new_n4053 , new_n4051 , new_n4052 );
  xnor     g03677 ( new_n4054 , new_n4051 , new_n4052 );
  nand     g03678 ( new_n4055 , pi109 , pi219 );
  nand     g03679 ( new_n4056 , pi014 , pi087 );
  xor      g03680 ( new_n4057 , new_n4055 , new_n4056 );
  nor      g03681 ( new_n4058 , new_n4054 , new_n4057 );
  nor      g03682 ( new_n4059 , new_n4053 , new_n4058 );
  nor      g03683 ( new_n4060 , new_n3951 , new_n3956 );
  nor      g03684 ( new_n4061 , new_n3958 , new_n4060 );
  nor      g03685 ( new_n4062 , new_n4059 , new_n4061 );
  xor      g03686 ( new_n4063 , new_n3807 , new_n3810 );
  xnor     g03687 ( new_n4064 , new_n4059 , new_n4061 );
  nor      g03688 ( new_n4065 , new_n4063 , new_n4064 );
  or       g03689 ( new_n4066 , new_n4062 , new_n4065 );
  xor      g03690 ( new_n4067 , new_n3811 , new_n3813 );
  nand     g03691 ( new_n4068 , new_n4066 , new_n4067 );
  xnor     g03692 ( new_n4069 , new_n3959 , new_n3969 );
  nand g03693 ( new_n4070 , new_n4069 , new_n4069 );
  xnor     g03694 ( new_n4071 , new_n4066 , new_n4067 );
  or       g03695 ( new_n4072 , new_n4070 , new_n4071 );
  nand     g03696 ( new_n4073 , new_n4068 , new_n4072 );
  xnor     g03697 ( new_n4074 , new_n3970 , new_n3987 );
  nand     g03698 ( new_n4075 , new_n4073 , new_n4074 );
  xor      g03699 ( new_n4076 , new_n4073 , new_n4074 );
  xnor     g03700 ( new_n4077 , new_n3814 , new_n3815 );
  nand     g03701 ( new_n4078 , new_n4076 , new_n4077 );
  nand     g03702 ( new_n4079 , new_n4075 , new_n4078 );
  xor      g03703 ( new_n4080 , new_n4046 , new_n4048 );
  nor      g03704 ( new_n4081 , new_n4079 , new_n4080 );
  nor      g03705 ( new_n4082 , new_n4049 , new_n4081 );
  xnor     g03706 ( new_n4083 , new_n4043 , new_n4044 );
  nor      g03707 ( new_n4084 , new_n4082 , new_n4083 );
  nor      g03708 ( new_n4085 , new_n4045 , new_n4084 );
  nand     g03709 ( new_n4086 , pi020 , pi184 );
  xor      g03710 ( new_n4087 , new_n4085 , new_n4086 );
  xor      g03711 ( new_n4088 , new_n3946 , new_n4087 );
  xor      g03712 ( new_n4089 , new_n3945 , new_n4088 );
  xor      g03713 ( new_n4090 , new_n3934 , new_n4089 );
  xor      g03714 ( new_n4091 , new_n3928 , new_n4090 );
  nand     g03715 ( new_n4092 , pi002 , pi123 );
  nand     g03716 ( new_n4093 , pi055 , pi099 );
  xor      g03717 ( new_n4094 , new_n4092 , new_n4093 );
  nand     g03718 ( new_n4095 , pi122 , pi230 );
  or       g03719 ( new_n4096 , new_n4029 , new_n4030 );
  nand     g03720 ( new_n4097 , new_n4031 , new_n4039 );
  nand     g03721 ( new_n4098 , new_n4096 , new_n4097 );
  xor      g03722 ( new_n4099 , new_n4095 , new_n4098 );
  nor      g03723 ( new_n4100 , new_n3640 , new_n3658 );
  nor      g03724 ( new_n4101 , new_n3659 , new_n3663 );
  nor      g03725 ( new_n4102 , new_n4100 , new_n4101 );
  nor      g03726 ( new_n4103 , new_n4006 , new_n4037 );
  nor      g03727 ( new_n4104 , new_n4036 , new_n4038 );
  nor      g03728 ( new_n4105 , new_n4103 , new_n4104 );
  xor      g03729 ( new_n4106 , new_n4102 , new_n4105 );
  xor      g03730 ( new_n4107 , new_n4099 , new_n4106 );
  xor      g03731 ( new_n4108 , new_n4094 , new_n4107 );
  nand     g03732 ( new_n4109 , pi071 , pi239 );
  nand     g03733 ( new_n4110 , new_n3638 , new_n3661 );
  nand     g03734 ( new_n4111 , new_n3660 , new_n3662 );
  nand     g03735 ( new_n4112 , new_n4110 , new_n4111 );
  nand     g03736 ( new_n4113 , new_n3652 , new_n3653 );
  nand     g03737 ( new_n4114 , new_n3654 , new_n3655 );
  nand     g03738 ( new_n4115 , new_n4113 , new_n4114 );
  xor      g03739 ( new_n4116 , new_n4112 , new_n4115 );
  xor      g03740 ( new_n4117 , new_n4109 , new_n4116 );
  xor      g03741 ( new_n4118 , new_n4108 , new_n4117 );
  xor      g03742 ( new_n4119 , new_n4091 , new_n4118 );
  xor      g03743 ( new_n4120 , new_n3673 , new_n4119 );
  nand     g03744 ( new_n4121 , pi020 , pi150 );
  nand     g03745 ( new_n4122 , pi029 , pi223 );
  nand     g03746 ( new_n4123 , pi020 , pi244 );
  nand     g03747 ( new_n4124 , new_n4122 , new_n4123 );
  nand     g03748 ( new_n4125 , pi060 , pi069 );
  xor      g03749 ( new_n4126 , new_n4122 , new_n4123 );
  nand     g03750 ( new_n4127 , new_n4125 , new_n4126 );
  nand     g03751 ( new_n4128 , new_n4124 , new_n4127 );
  nand     g03752 ( new_n4129 , new_n4121 , new_n4128 );
  xor      g03753 ( new_n4130 , new_n3693 , new_n3694 );
  nand g03754 ( new_n4131 , new_n4130 , new_n4130 );
  xor      g03755 ( new_n4132 , new_n4121 , new_n4128 );
  nand     g03756 ( new_n4133 , new_n4131 , new_n4132 );
  nand     g03757 ( new_n4134 , new_n4129 , new_n4133 );
  nand     g03758 ( new_n4135 , pi060 , pi150 );
  nand     g03759 ( new_n4136 , pi020 , pi221 );
  and      g03760 ( new_n4137 , new_n4135 , new_n4136 );
  nor      g03761 ( new_n4138 , new_n3675 , new_n4121 );
  nor      g03762 ( new_n4139 , new_n4137 , new_n4138 );
  xor      g03763 ( new_n4140 , new_n3697 , new_n3698 );
  xor      g03764 ( new_n4141 , new_n4139 , new_n4140 );
  nor      g03765 ( new_n4142 , new_n4134 , new_n4141 );
  nand g03766 ( new_n4143 , new_n4140 , new_n4140 );
  nand     g03767 ( new_n4144 , new_n4139 , new_n4143 );
  nand g03768 ( new_n4145 , new_n4144 , new_n4144 );
  nor      g03769 ( new_n4146 , new_n4138 , new_n4145 );
  nand g03770 ( new_n4147 , new_n4146 , new_n4146 );
  nor      g03771 ( new_n4148 , new_n4142 , new_n4147 );
  and      g03772 ( new_n4149 , new_n4138 , new_n4142 );
  or       g03773 ( new_n4150 , new_n4148 , new_n4149 );
  xor      g03774 ( new_n4151 , new_n3702 , new_n3709 );
  nand g03775 ( new_n4152 , new_n4151 , new_n4151 );
  nor      g03776 ( new_n4153 , new_n4150 , new_n4152 );
  nor      g03777 ( new_n4154 , new_n4148 , new_n4153 );
  nand     g03778 ( new_n4155 , pi074 , pi219 );
  nand     g03779 ( new_n4156 , pi010 , pi160 );
  xor      g03780 ( new_n4157 , new_n4155 , new_n4156 );
  xor      g03781 ( new_n4158 , new_n4154 , new_n4157 );
  nand     g03782 ( new_n4159 , pi186 , pi251 );
  nand     g03783 ( new_n4160 , pi160 , pi196 );
  nand     g03784 ( new_n4161 , pi150 , pi160 );
  nand     g03785 ( new_n4162 , pi160 , pi244 );
  nand     g03786 ( new_n4163 , pi020 , pi069 );
  nand     g03787 ( new_n4164 , new_n4162 , new_n4163 );
  nand     g03788 ( new_n4165 , pi029 , pi060 );
  xor      g03789 ( new_n4166 , new_n4162 , new_n4163 );
  nand     g03790 ( new_n4167 , new_n4165 , new_n4166 );
  nand     g03791 ( new_n4168 , new_n4164 , new_n4167 );
  nand     g03792 ( new_n4169 , new_n4161 , new_n4168 );
  xor      g03793 ( new_n4170 , new_n4125 , new_n4126 );
  xor      g03794 ( new_n4171 , new_n4161 , new_n4168 );
  nand     g03795 ( new_n4172 , new_n4170 , new_n4171 );
  nand     g03796 ( new_n4173 , new_n4169 , new_n4172 );
  nand     g03797 ( new_n4174 , pi160 , pi221 );
  xor      g03798 ( new_n4175 , new_n4130 , new_n4132 );
  xor      g03799 ( new_n4176 , new_n4174 , new_n4175 );
  xor      g03800 ( new_n4177 , new_n4173 , new_n4176 );
  xor      g03801 ( new_n4178 , new_n4165 , new_n4166 );
  nand g03802 ( new_n4179 , new_n4178 , new_n4178 );
  nand     g03803 ( new_n4180 , pi029 , pi160 );
  nor      g03804 ( new_n4181 , new_n4163 , new_n4180 );
  nand     g03805 ( new_n4182 , new_n4179 , new_n4181 );
  nand g03806 ( new_n4183 , new_n4182 , new_n4182 );
  xnor     g03807 ( new_n4184 , new_n4170 , new_n4171 );
  and      g03808 ( new_n4185 , new_n4183 , new_n4184 );
  nand     g03809 ( new_n4186 , new_n4177 , new_n4185 );
  nand     g03810 ( new_n4187 , new_n4160 , new_n4186 );
  xor      g03811 ( new_n4188 , new_n4160 , new_n4186 );
  nand g03812 ( new_n4189 , new_n4188 , new_n4188 );
  nand g03813 ( new_n4190 , new_n4175 , new_n4175 );
  nor      g03814 ( new_n4191 , new_n4174 , new_n4190 );
  nor      g03815 ( new_n4192 , new_n4173 , new_n4176 );
  nor      g03816 ( new_n4193 , new_n4191 , new_n4192 );
  xor      g03817 ( new_n4194 , new_n4134 , new_n4141 );
  nand g03818 ( new_n4195 , new_n4194 , new_n4194 );
  xor      g03819 ( new_n4196 , new_n4193 , new_n4195 );
  or       g03820 ( new_n4197 , new_n4189 , new_n4196 );
  nand     g03821 ( new_n4198 , new_n4187 , new_n4197 );
  or       g03822 ( new_n4199 , new_n4193 , new_n4195 );
  xor      g03823 ( new_n4200 , new_n4150 , new_n4151 );
  xor      g03824 ( new_n4201 , new_n4199 , new_n4200 );
  xnor     g03825 ( new_n4202 , new_n4198 , new_n4201 );
  xor      g03826 ( new_n4203 , new_n4189 , new_n4196 );
  xor      g03827 ( new_n4204 , new_n4177 , new_n4185 );
  xor      g03828 ( new_n4205 , new_n4182 , new_n4184 );
  xor      g03829 ( new_n4206 , new_n4178 , new_n4181 );
  xnor     g03830 ( new_n4207 , new_n4063 , new_n4064 );
  xnor     g03831 ( new_n4208 , new_n3950 , new_n4050 );
  or       g03832 ( new_n4209 , new_n3890 , new_n4208 );
  nand     g03833 ( new_n4210 , pi138 , pi186 );
  nand     g03834 ( new_n4211 , pi132 , pi182 );
  nand     g03835 ( new_n4212 , new_n4210 , new_n4211 );
  nand     g03836 ( new_n4213 , new_n3891 , new_n4212 );
  nor      g03837 ( new_n4214 , new_n4209 , new_n4213 );
  xnor     g03838 ( new_n4215 , new_n4209 , new_n4213 );
  xor      g03839 ( new_n4216 , new_n4054 , new_n4057 );
  nor      g03840 ( new_n4217 , new_n4215 , new_n4216 );
  nor      g03841 ( new_n4218 , new_n4214 , new_n4217 );
  xor      g03842 ( new_n4219 , new_n3889 , new_n3891 );
  xor      g03843 ( new_n4220 , new_n4218 , new_n4219 );
  xor      g03844 ( new_n4221 , new_n4207 , new_n4220 );
  and      g03845 ( new_n4222 , new_n4206 , new_n4221 );
  xnor     g03846 ( new_n4223 , new_n4206 , new_n4221 );
  xor      g03847 ( new_n4224 , new_n3890 , new_n4208 );
  nand g03848 ( new_n4225 , new_n4224 , new_n4224 );
  nor      g03849 ( new_n4226 , new_n4180 , new_n4225 );
  nand     g03850 ( new_n4227 , pi020 , pi029 );
  nand     g03851 ( new_n4228 , pi069 , pi160 );
  and      g03852 ( new_n4229 , new_n4227 , new_n4228 );
  nor      g03853 ( new_n4230 , new_n4181 , new_n4229 );
  nor      g03854 ( new_n4231 , new_n4226 , new_n4230 );
  xnor     g03855 ( new_n4232 , new_n4226 , new_n4230 );
  xor      g03856 ( new_n4233 , new_n4215 , new_n4216 );
  nor      g03857 ( new_n4234 , new_n4232 , new_n4233 );
  nor      g03858 ( new_n4235 , new_n4231 , new_n4234 );
  nor      g03859 ( new_n4236 , new_n4223 , new_n4235 );
  or       g03860 ( new_n4237 , new_n4222 , new_n4236 );
  nor      g03861 ( new_n4238 , new_n4205 , new_n4237 );
  nand g03862 ( new_n4239 , new_n4218 , new_n4218 );
  nand     g03863 ( new_n4240 , new_n4239 , new_n4219 );
  nand g03864 ( new_n4241 , new_n4220 , new_n4220 );
  nand     g03865 ( new_n4242 , new_n4207 , new_n4241 );
  nand     g03866 ( new_n4243 , new_n4240 , new_n4242 );
  xor      g03867 ( new_n4244 , new_n3892 , new_n3893 );
  xor      g03868 ( new_n4245 , new_n4069 , new_n4071 );
  xnor     g03869 ( new_n4246 , new_n4244 , new_n4245 );
  xor      g03870 ( new_n4247 , new_n4243 , new_n4246 );
  xnor     g03871 ( new_n4248 , new_n4205 , new_n4237 );
  nor      g03872 ( new_n4249 , new_n4247 , new_n4248 );
  or       g03873 ( new_n4250 , new_n4238 , new_n4249 );
  nor      g03874 ( new_n4251 , new_n4204 , new_n4250 );
  xnor     g03875 ( new_n4252 , new_n4204 , new_n4250 );
  xor      g03876 ( new_n4253 , new_n4076 , new_n4077 );
  nor      g03877 ( new_n4254 , new_n4244 , new_n4245 );
  nor      g03878 ( new_n4255 , new_n4243 , new_n4246 );
  or       g03879 ( new_n4256 , new_n4254 , new_n4255 );
  xnor     g03880 ( new_n4257 , new_n3894 , new_n3895 );
  xnor     g03881 ( new_n4258 , new_n4256 , new_n4257 );
  xor      g03882 ( new_n4259 , new_n4253 , new_n4258 );
  nor      g03883 ( new_n4260 , new_n4252 , new_n4259 );
  or       g03884 ( new_n4261 , new_n4251 , new_n4260 );
  nor      g03885 ( new_n4262 , new_n4203 , new_n4261 );
  xor      g03886 ( new_n4263 , new_n4079 , new_n4080 );
  nor      g03887 ( new_n4264 , new_n4256 , new_n4257 );
  nor      g03888 ( new_n4265 , new_n4253 , new_n4258 );
  nor      g03889 ( new_n4266 , new_n4264 , new_n4265 );
  xor      g03890 ( new_n4267 , new_n3896 , new_n3897 );
  xor      g03891 ( new_n4268 , new_n4266 , new_n4267 );
  xor      g03892 ( new_n4269 , new_n4263 , new_n4268 );
  xnor     g03893 ( new_n4270 , new_n4203 , new_n4261 );
  nor      g03894 ( new_n4271 , new_n4269 , new_n4270 );
  nor      g03895 ( new_n4272 , new_n4262 , new_n4271 );
  nor      g03896 ( new_n4273 , new_n4202 , new_n4272 );
  xnor     g03897 ( new_n4274 , new_n4202 , new_n4272 );
  nand g03898 ( new_n4275 , new_n4267 , new_n4267 );
  nor      g03899 ( new_n4276 , new_n4266 , new_n4275 );
  nand g03900 ( new_n4277 , new_n4263 , new_n4263 );
  nor      g03901 ( new_n4278 , new_n4277 , new_n4268 );
  nor      g03902 ( new_n4279 , new_n4276 , new_n4278 );
  xnor     g03903 ( new_n4280 , new_n3885 , new_n3899 );
  xor      g03904 ( new_n4281 , new_n4279 , new_n4280 );
  xnor     g03905 ( new_n4282 , new_n4082 , new_n4083 );
  xor      g03906 ( new_n4283 , new_n4281 , new_n4282 );
  nor      g03907 ( new_n4284 , new_n4274 , new_n4283 );
  nor      g03908 ( new_n4285 , new_n4273 , new_n4284 );
  xor      g03909 ( new_n4286 , new_n4159 , new_n4285 );
  xor      g03910 ( new_n4287 , new_n4158 , new_n4286 );
  xor      g03911 ( new_n4288 , new_n4120 , new_n4287 );
  nand     g03912 ( new_n4289 , pi221 , pi223 );
  or       g03913 ( new_n4290 , new_n3881 , new_n3882 );
  nand     g03914 ( new_n4291 , new_n3880 , new_n4290 );
  xor      g03915 ( new_n4292 , new_n4289 , new_n4291 );
  nand     g03916 ( new_n4293 , new_n3676 , new_n3677 );
  nand     g03917 ( new_n4294 , new_n3675 , new_n3678 );
  nand     g03918 ( new_n4295 , new_n4293 , new_n4294 );
  and      g03919 ( new_n4296 , new_n4022 , new_n4041 );
  nor      g03920 ( new_n4297 , new_n4021 , new_n4042 );
  nor      g03921 ( new_n4298 , new_n4296 , new_n4297 );
  xor      g03922 ( new_n4299 , new_n4295 , new_n4298 );
  xor      g03923 ( new_n4300 , new_n4292 , new_n4299 );
  nand     g03924 ( new_n4301 , new_n4279 , new_n4280 );
  nand     g03925 ( new_n4302 , new_n4281 , new_n4282 );
  nand     g03926 ( new_n4303 , new_n4301 , new_n4302 );
  nand     g03927 ( new_n4304 , new_n4001 , new_n4024 );
  or       g03928 ( new_n4305 , new_n4026 , new_n4040 );
  nand     g03929 ( new_n4306 , new_n4304 , new_n4305 );
  nand g03930 ( new_n4307 , new_n4200 , new_n4200 );
  nor      g03931 ( new_n4308 , new_n4199 , new_n4307 );
  nor      g03932 ( new_n4309 , new_n4198 , new_n4201 );
  nor      g03933 ( new_n4310 , new_n4308 , new_n4309 );
  xor      g03934 ( new_n4311 , new_n4306 , new_n4310 );
  xor      g03935 ( new_n4312 , new_n4303 , new_n4311 );
  nand     g03936 ( new_n4313 , pi135 , pi173 );
  nand g03937 ( new_n4314 , new_n4032 , new_n4032 );
  nor      g03938 ( new_n4315 , new_n4314 , new_n4034 );
  nor      g03939 ( new_n4316 , new_n4005 , new_n4035 );
  nor      g03940 ( new_n4317 , new_n4315 , new_n4316 );
  xor      g03941 ( new_n4318 , new_n4313 , new_n4317 );
  xor      g03942 ( new_n4319 , new_n4312 , new_n4318 );
  xor      g03943 ( new_n4320 , new_n4300 , new_n4319 );
  xor      g03944 ( po013 , new_n4288 , new_n4320 );
  nand     g03945 ( new_n4322 , pi036 , pi103 );
  nor      g03946 ( new_n4323 , new_n1012 , new_n1023 );
  nand     g03947 ( new_n4324 , pi016 , pi194 );
  nand     g03948 ( new_n4325 , pi143 , pi247 );
  nand     g03949 ( new_n4326 , pi057 , pi080 );
  xor      g03950 ( new_n4327 , new_n4325 , new_n4326 );
  xor      g03951 ( new_n4328 , new_n4324 , new_n4327 );
  nand     g03952 ( new_n4329 , pi085 , pi117 );
  nand     g03953 ( new_n4330 , new_n1019 , new_n1020 );
  nand     g03954 ( new_n4331 , new_n1018 , new_n1021 );
  nand     g03955 ( new_n4332 , new_n4330 , new_n4331 );
  xor      g03956 ( new_n4333 , new_n4329 , new_n4332 );
  xor      g03957 ( new_n4334 , new_n4328 , new_n4333 );
  nand     g03958 ( new_n4335 , pi103 , pi180 );
  nand     g03959 ( new_n4336 , new_n1013 , new_n1016 );
  nand     g03960 ( new_n4337 , new_n1017 , new_n1022 );
  nand     g03961 ( new_n4338 , new_n4336 , new_n4337 );
  xnor     g03962 ( new_n4339 , new_n4335 , new_n4338 );
  xor      g03963 ( new_n4340 , new_n4334 , new_n4339 );
  nand     g03964 ( new_n4341 , new_n4323 , new_n4340 );
  nand     g03965 ( new_n4342 , new_n4322 , new_n4341 );
  nand     g03966 ( new_n4343 , pi016 , pi180 );
  nor      g03967 ( new_n4344 , new_n4329 , new_n4343 );
  nand g03968 ( new_n4345 , new_n4344 , new_n4344 );
  nand     g03969 ( new_n4346 , pi016 , pi085 );
  nand     g03970 ( new_n4347 , pi117 , pi180 );
  nand     g03971 ( new_n4348 , new_n4346 , new_n4347 );
  nand     g03972 ( new_n4349 , new_n4345 , new_n4348 );
  nand     g03973 ( new_n4350 , pi080 , pi194 );
  nand     g03974 ( new_n4351 , new_n4325 , new_n4326 );
  nand     g03975 ( new_n4352 , new_n4324 , new_n4327 );
  nand     g03976 ( new_n4353 , new_n4351 , new_n4352 );
  xor      g03977 ( new_n4354 , new_n4350 , new_n4353 );
  nand     g03978 ( new_n4355 , pi057 , pi247 );
  nand     g03979 ( new_n4356 , pi143 , pi234 );
  nand     g03980 ( new_n4357 , new_n4355 , new_n4356 );
  nand     g03981 ( new_n4358 , pi057 , pi234 );
  nor      g03982 ( new_n4359 , new_n4325 , new_n4358 );
  nand g03983 ( new_n4360 , new_n4359 , new_n4359 );
  nand     g03984 ( new_n4361 , new_n4357 , new_n4360 );
  xor      g03985 ( new_n4362 , new_n4354 , new_n4361 );
  xnor     g03986 ( new_n4363 , new_n4349 , new_n4362 );
  nand     g03987 ( new_n4364 , new_n4329 , new_n4332 );
  nand     g03988 ( new_n4365 , new_n4328 , new_n4333 );
  nand     g03989 ( new_n4366 , new_n4364 , new_n4365 );
  xor      g03990 ( new_n4367 , new_n4363 , new_n4366 );
  nand g03991 ( new_n4368 , new_n4367 , new_n4367 );
  nor      g03992 ( new_n4369 , new_n4335 , new_n4338 );
  nor      g03993 ( new_n4370 , new_n4334 , new_n4339 );
  nor      g03994 ( new_n4371 , new_n4369 , new_n4370 );
  xor      g03995 ( new_n4372 , new_n4368 , new_n4371 );
  nand g03996 ( new_n4373 , new_n4372 , new_n4372 );
  xor      g03997 ( new_n4374 , new_n4322 , new_n4341 );
  nand     g03998 ( new_n4375 , new_n4373 , new_n4374 );
  nand     g03999 ( new_n4376 , new_n4342 , new_n4375 );
  nor      g04000 ( new_n4377 , new_n4368 , new_n4371 );
  nor      g04001 ( new_n4378 , new_n4349 , new_n4362 );
  nor      g04002 ( new_n4379 , new_n4363 , new_n4366 );
  xor      g04003 ( new_n4380 , new_n4345 , new_n4379 );
  nand g04004 ( new_n4381 , new_n4380 , new_n4380 );
  nor      g04005 ( new_n4382 , new_n4378 , new_n4381 );
  nand     g04006 ( new_n4383 , pi080 , pi085 );
  xor      g04007 ( new_n4384 , new_n4359 , new_n4383 );
  nand     g04008 ( new_n4385 , pi143 , pi214 );
  nand     g04009 ( new_n4386 , pi194 , pi247 );
  xor      g04010 ( new_n4387 , new_n4385 , new_n4386 );
  xor      g04011 ( new_n4388 , new_n4358 , new_n4387 );
  xor      g04012 ( new_n4389 , new_n4384 , new_n4388 );
  nand     g04013 ( new_n4390 , pi036 , pi117 );
  nand     g04014 ( new_n4391 , pi068 , pi103 );
  xor      g04015 ( new_n4392 , new_n4390 , new_n4391 );
  xor      g04016 ( new_n4393 , new_n4343 , new_n4392 );
  nor      g04017 ( new_n4394 , new_n4350 , new_n4353 );
  nand g04018 ( new_n4395 , new_n4354 , new_n4354 );
  nor      g04019 ( new_n4396 , new_n4395 , new_n4361 );
  nor      g04020 ( new_n4397 , new_n4394 , new_n4396 );
  xor      g04021 ( new_n4398 , new_n4393 , new_n4397 );
  xor      g04022 ( new_n4399 , new_n4389 , new_n4398 );
  xor      g04023 ( new_n4400 , new_n4382 , new_n4399 );
  xor      g04024 ( new_n4401 , new_n4377 , new_n4400 );
  xor      g04025 ( new_n4402 , new_n4376 , new_n4401 );
  and      g04026 ( new_n4403 , new_n975 , new_n1010 );
  nor      g04027 ( new_n4404 , new_n4403 , new_n1024 );
  nor      g04028 ( new_n4405 , new_n1025 , new_n1074 );
  nor      g04029 ( new_n4406 , new_n4404 , new_n4405 );
  xnor     g04030 ( new_n4407 , new_n4323 , new_n4340 );
  nand     g04031 ( new_n4408 , new_n4406 , new_n4407 );
  xor      g04032 ( new_n4409 , new_n4406 , new_n4407 );
  nor      g04033 ( new_n4410 , new_n1044 , new_n1055 );
  nand     g04034 ( new_n4411 , pi144 , pi163 );
  nand     g04035 ( new_n4412 , new_n1051 , new_n1052 );
  nand     g04036 ( new_n4413 , new_n1050 , new_n1053 );
  nand     g04037 ( new_n4414 , new_n4412 , new_n4413 );
  nand     g04038 ( new_n4415 , pi012 , pi148 );
  xor      g04039 ( new_n4416 , new_n4414 , new_n4415 );
  nand     g04040 ( new_n4417 , pi061 , pi228 );
  nand     g04041 ( new_n4418 , pi116 , pi188 );
  nand     g04042 ( new_n4419 , pi039 , pi178 );
  xor      g04043 ( new_n4420 , new_n4418 , new_n4419 );
  xor      g04044 ( new_n4421 , new_n4417 , new_n4420 );
  xor      g04045 ( new_n4422 , new_n4416 , new_n4421 );
  xnor     g04046 ( new_n4423 , new_n4411 , new_n4422 );
  nand     g04047 ( new_n4424 , new_n1045 , new_n1048 );
  nand     g04048 ( new_n4425 , new_n1049 , new_n1054 );
  nand     g04049 ( new_n4426 , new_n4424 , new_n4425 );
  xor      g04050 ( new_n4427 , new_n4423 , new_n4426 );
  xor      g04051 ( new_n4428 , new_n4410 , new_n4427 );
  nand     g04052 ( new_n4429 , new_n1042 , new_n1056 );
  nand     g04053 ( new_n4430 , new_n1029 , new_n1057 );
  nand     g04054 ( new_n4431 , new_n4429 , new_n4430 );
  nor      g04055 ( new_n4432 , new_n1030 , new_n1041 );
  nand     g04056 ( new_n4433 , pi107 , pi118 );
  nor      g04057 ( new_n4434 , new_n1036 , new_n1039 );
  nor      g04058 ( new_n4435 , new_n1035 , new_n1040 );
  nor      g04059 ( new_n4436 , new_n4434 , new_n4435 );
  xor      g04060 ( new_n4437 , new_n4433 , new_n4436 );
  nand     g04061 ( new_n4438 , pi049 , pi108 );
  nand     g04062 ( new_n4439 , pi042 , pi245 );
  nand     g04063 ( new_n4440 , pi051 , pi201 );
  xor      g04064 ( new_n4441 , new_n4439 , new_n4440 );
  xor      g04065 ( new_n4442 , new_n4438 , new_n4441 );
  nand     g04066 ( new_n4443 , pi007 , pi171 );
  nand     g04067 ( new_n4444 , new_n1032 , new_n1033 );
  nand     g04068 ( new_n4445 , new_n1031 , new_n1034 );
  nand     g04069 ( new_n4446 , new_n4444 , new_n4445 );
  xor      g04070 ( new_n4447 , new_n4443 , new_n4446 );
  xnor     g04071 ( new_n4448 , new_n4442 , new_n4447 );
  xor      g04072 ( new_n4449 , new_n4437 , new_n4448 );
  xor      g04073 ( new_n4450 , new_n4432 , new_n4449 );
  xnor     g04074 ( new_n4451 , new_n4431 , new_n4450 );
  xor      g04075 ( new_n4452 , new_n4428 , new_n4451 );
  nand g04076 ( new_n4453 , new_n1071 , new_n1071 );
  nand     g04077 ( new_n4454 , new_n1061 , new_n4453 );
  nand g04078 ( new_n4455 , new_n4454 , new_n4454 );
  nand     g04079 ( new_n4456 , pi162 , pi167 );
  nand     g04080 ( new_n4457 , pi179 , pi240 );
  nand     g04081 ( new_n4458 , pi033 , pi149 );
  xor      g04082 ( new_n4459 , new_n4457 , new_n4458 );
  xor      g04083 ( new_n4460 , new_n4456 , new_n4459 );
  nand     g04084 ( new_n4461 , new_n1067 , new_n1068 );
  nand     g04085 ( new_n4462 , new_n1066 , new_n1069 );
  nand     g04086 ( new_n4463 , new_n4461 , new_n4462 );
  nand     g04087 ( new_n4464 , pi048 , pi134 );
  xor      g04088 ( new_n4465 , new_n4463 , new_n4464 );
  xor      g04089 ( new_n4466 , new_n4460 , new_n4465 );
  nand     g04090 ( new_n4467 , pi175 , pi237 );
  nor      g04091 ( new_n4468 , new_n1063 , new_n1064 );
  nand g04092 ( new_n4469 , new_n1070 , new_n1070 );
  nand     g04093 ( new_n4470 , new_n1065 , new_n4469 );
  nand g04094 ( new_n4471 , new_n4470 , new_n4470 );
  or       g04095 ( new_n4472 , new_n4468 , new_n4471 );
  xor      g04096 ( new_n4473 , new_n4467 , new_n4472 );
  xor      g04097 ( new_n4474 , new_n4466 , new_n4473 );
  xor      g04098 ( new_n4475 , new_n4455 , new_n4474 );
  and      g04099 ( new_n4476 , new_n1060 , new_n1072 );
  nor      g04100 ( new_n4477 , new_n1058 , new_n1073 );
  nor      g04101 ( new_n4478 , new_n4476 , new_n4477 );
  xnor     g04102 ( new_n4479 , new_n4475 , new_n4478 );
  xnor     g04103 ( new_n4480 , new_n4452 , new_n4479 );
  nand     g04104 ( new_n4481 , new_n4409 , new_n4480 );
  and      g04105 ( new_n4482 , new_n4408 , new_n4481 );
  xor      g04106 ( new_n4483 , new_n4372 , new_n4374 );
  nor      g04107 ( new_n4484 , new_n4482 , new_n4483 );
  xnor     g04108 ( new_n4485 , new_n4482 , new_n4483 );
  nor      g04109 ( new_n4486 , new_n4431 , new_n4450 );
  nor      g04110 ( new_n4487 , new_n4428 , new_n4451 );
  or       g04111 ( new_n4488 , new_n4486 , new_n4487 );
  nand     g04112 ( new_n4489 , new_n4432 , new_n4449 );
  nand     g04113 ( new_n4490 , pi107 , pi113 );
  xor      g04114 ( new_n4491 , new_n4489 , new_n4490 );
  nand     g04115 ( new_n4492 , new_n4443 , new_n4446 );
  nand     g04116 ( new_n4493 , new_n4442 , new_n4447 );
  nand     g04117 ( new_n4494 , new_n4492 , new_n4493 );
  nand     g04118 ( new_n4495 , pi007 , pi049 );
  nand     g04119 ( new_n4496 , pi118 , pi171 );
  and      g04120 ( new_n4497 , new_n4495 , new_n4496 );
  nand     g04121 ( new_n4498 , pi049 , pi118 );
  nor      g04122 ( new_n4499 , new_n4443 , new_n4498 );
  or       g04123 ( new_n4500 , new_n4497 , new_n4499 );
  nand     g04124 ( new_n4501 , new_n4439 , new_n4440 );
  nand     g04125 ( new_n4502 , new_n4438 , new_n4441 );
  nand     g04126 ( new_n4503 , new_n4501 , new_n4502 );
  nand     g04127 ( new_n4504 , pi108 , pi245 );
  nand     g04128 ( new_n4505 , pi042 , pi201 );
  nand     g04129 ( new_n4506 , pi051 , pi156 );
  nand     g04130 ( new_n4507 , new_n4505 , new_n4506 );
  nand     g04131 ( new_n4508 , pi042 , pi156 );
  nor      g04132 ( new_n4509 , new_n4440 , new_n4508 );
  nand g04133 ( new_n4510 , new_n4509 , new_n4509 );
  nand     g04134 ( new_n4511 , new_n4507 , new_n4510 );
  xor      g04135 ( new_n4512 , new_n4504 , new_n4511 );
  xor      g04136 ( new_n4513 , new_n4503 , new_n4512 );
  xor      g04137 ( new_n4514 , new_n4500 , new_n4513 );
  nand g04138 ( new_n4515 , new_n4514 , new_n4514 );
  xor      g04139 ( new_n4516 , new_n4494 , new_n4515 );
  nand g04140 ( new_n4517 , new_n4516 , new_n4516 );
  nor      g04141 ( new_n4518 , new_n4433 , new_n4436 );
  and      g04142 ( new_n4519 , new_n4437 , new_n4448 );
  nor      g04143 ( new_n4520 , new_n4518 , new_n4519 );
  xor      g04144 ( new_n4521 , new_n4517 , new_n4520 );
  xor      g04145 ( new_n4522 , new_n4491 , new_n4521 );
  nand     g04146 ( new_n4523 , new_n4410 , new_n4427 );
  nand     g04147 ( new_n4524 , pi098 , pi163 );
  nor      g04148 ( new_n4525 , new_n4411 , new_n4422 );
  nor      g04149 ( new_n4526 , new_n4423 , new_n4426 );
  nor      g04150 ( new_n4527 , new_n4525 , new_n4526 );
  nand     g04151 ( new_n4528 , new_n4414 , new_n4415 );
  nand     g04152 ( new_n4529 , new_n4416 , new_n4421 );
  nand     g04153 ( new_n4530 , new_n4528 , new_n4529 );
  nand     g04154 ( new_n4531 , pi012 , pi228 );
  nand     g04155 ( new_n4532 , pi144 , pi148 );
  and      g04156 ( new_n4533 , new_n4531 , new_n4532 );
  nand     g04157 ( new_n4534 , pi144 , pi228 );
  nor      g04158 ( new_n4535 , new_n4415 , new_n4534 );
  or       g04159 ( new_n4536 , new_n4533 , new_n4535 );
  nand     g04160 ( new_n4537 , new_n4418 , new_n4419 );
  nand     g04161 ( new_n4538 , new_n4417 , new_n4420 );
  nand     g04162 ( new_n4539 , new_n4537 , new_n4538 );
  nand     g04163 ( new_n4540 , pi039 , pi061 );
  nand     g04164 ( new_n4541 , pi070 , pi178 );
  or       g04165 ( new_n4542 , new_n4418 , new_n4541 );
  nand     g04166 ( new_n4543 , pi116 , pi178 );
  nand     g04167 ( new_n4544 , pi070 , pi188 );
  nand     g04168 ( new_n4545 , new_n4543 , new_n4544 );
  nand     g04169 ( new_n4546 , new_n4542 , new_n4545 );
  xor      g04170 ( new_n4547 , new_n4540 , new_n4546 );
  xor      g04171 ( new_n4548 , new_n4539 , new_n4547 );
  xor      g04172 ( new_n4549 , new_n4536 , new_n4548 );
  nand g04173 ( new_n4550 , new_n4549 , new_n4549 );
  xor      g04174 ( new_n4551 , new_n4530 , new_n4550 );
  xor      g04175 ( new_n4552 , new_n4527 , new_n4551 );
  xor      g04176 ( new_n4553 , new_n4524 , new_n4552 );
  xor      g04177 ( new_n4554 , new_n4523 , new_n4553 );
  xor      g04178 ( new_n4555 , new_n4522 , new_n4554 );
  xor      g04179 ( new_n4556 , new_n4488 , new_n4555 );
  nand     g04180 ( new_n4557 , new_n4475 , new_n4478 );
  or       g04181 ( new_n4558 , new_n4452 , new_n4479 );
  nand     g04182 ( new_n4559 , new_n4557 , new_n4558 );
  nand     g04183 ( new_n4560 , new_n4463 , new_n4464 );
  nand     g04184 ( new_n4561 , new_n4460 , new_n4465 );
  nand     g04185 ( new_n4562 , new_n4560 , new_n4561 );
  nand     g04186 ( new_n4563 , pi033 , pi181 );
  nor      g04187 ( new_n4564 , new_n4456 , new_n4563 );
  nand g04188 ( new_n4565 , new_n4564 , new_n4564 );
  nand     g04189 ( new_n4566 , pi033 , pi167 );
  nand     g04190 ( new_n4567 , pi162 , pi181 );
  nand     g04191 ( new_n4568 , new_n4566 , new_n4567 );
  nand     g04192 ( new_n4569 , new_n4565 , new_n4568 );
  nand     g04193 ( new_n4570 , pi149 , pi179 );
  nand     g04194 ( new_n4571 , new_n4457 , new_n4458 );
  nand     g04195 ( new_n4572 , new_n4456 , new_n4459 );
  nand     g04196 ( new_n4573 , new_n4571 , new_n4572 );
  xnor     g04197 ( new_n4574 , new_n4570 , new_n4573 );
  xor      g04198 ( new_n4575 , new_n4569 , new_n4574 );
  nand     g04199 ( new_n4576 , pi048 , pi240 );
  nand     g04200 ( new_n4577 , pi134 , pi237 );
  and      g04201 ( new_n4578 , new_n4576 , new_n4577 );
  nand     g04202 ( new_n4579 , pi237 , pi240 );
  nor      g04203 ( new_n4580 , new_n4464 , new_n4579 );
  or       g04204 ( new_n4581 , new_n4578 , new_n4580 );
  xor      g04205 ( new_n4582 , new_n4575 , new_n4581 );
  xor      g04206 ( new_n4583 , new_n4562 , new_n4582 );
  nand g04207 ( new_n4584 , new_n4583 , new_n4583 );
  nand g04208 ( new_n4585 , new_n4472 , new_n4472 );
  nor      g04209 ( new_n4586 , new_n4467 , new_n4585 );
  nor      g04210 ( new_n4587 , new_n4466 , new_n4473 );
  nor      g04211 ( new_n4588 , new_n4586 , new_n4587 );
  xor      g04212 ( new_n4589 , new_n4584 , new_n4588 );
  nand     g04213 ( new_n4590 , new_n4455 , new_n4474 );
  nand     g04214 ( new_n4591 , pi175 , pi238 );
  xor      g04215 ( new_n4592 , new_n4590 , new_n4591 );
  xor      g04216 ( new_n4593 , new_n4589 , new_n4592 );
  xor      g04217 ( new_n4594 , new_n4559 , new_n4593 );
  xor      g04218 ( new_n4595 , new_n4556 , new_n4594 );
  nor      g04219 ( new_n4596 , new_n4485 , new_n4595 );
  nor      g04220 ( new_n4597 , new_n4484 , new_n4596 );
  xnor     g04221 ( new_n4598 , new_n4402 , new_n4597 );
  nand     g04222 ( new_n4599 , new_n4524 , new_n4552 );
  nand     g04223 ( new_n4600 , new_n4523 , new_n4553 );
  nand     g04224 ( new_n4601 , new_n4599 , new_n4600 );
  nand g04225 ( new_n4602 , new_n4551 , new_n4551 );
  nor      g04226 ( new_n4603 , new_n4527 , new_n4602 );
  nor      g04227 ( new_n4604 , new_n4536 , new_n4548 );
  nor      g04228 ( new_n4605 , new_n4530 , new_n4550 );
  xor      g04229 ( new_n4606 , new_n4535 , new_n4605 );
  nor      g04230 ( new_n4607 , new_n4604 , new_n4606 );
  nand     g04231 ( new_n4608 , pi098 , pi148 );
  nand     g04232 ( new_n4609 , pi043 , pi163 );
  xor      g04233 ( new_n4610 , new_n4608 , new_n4609 );
  xnor     g04234 ( new_n4611 , new_n4534 , new_n4610 );
  nand     g04235 ( new_n4612 , new_n4540 , new_n4546 );
  nand     g04236 ( new_n4613 , new_n4539 , new_n4547 );
  nand     g04237 ( new_n4614 , new_n4612 , new_n4613 );
  nand g04238 ( new_n4615 , new_n4614 , new_n4614 );
  xor      g04239 ( new_n4616 , new_n4611 , new_n4615 );
  nand     g04240 ( new_n4617 , pi012 , pi039 );
  xor      g04241 ( new_n4618 , new_n4542 , new_n4617 );
  nand     g04242 ( new_n4619 , pi115 , pi188 );
  nand     g04243 ( new_n4620 , pi061 , pi116 );
  xor      g04244 ( new_n4621 , new_n4619 , new_n4620 );
  xor      g04245 ( new_n4622 , new_n4541 , new_n4621 );
  xor      g04246 ( new_n4623 , new_n4618 , new_n4622 );
  xor      g04247 ( new_n4624 , new_n4616 , new_n4623 );
  xor      g04248 ( new_n4625 , new_n4607 , new_n4624 );
  xor      g04249 ( new_n4626 , new_n4603 , new_n4625 );
  xor      g04250 ( new_n4627 , new_n4601 , new_n4626 );
  nor      g04251 ( new_n4628 , new_n4517 , new_n4520 );
  nor      g04252 ( new_n4629 , new_n4500 , new_n4513 );
  nor      g04253 ( new_n4630 , new_n4494 , new_n4515 );
  xor      g04254 ( new_n4631 , new_n4499 , new_n4630 );
  nor      g04255 ( new_n4632 , new_n4629 , new_n4631 );
  nand     g04256 ( new_n4633 , pi007 , pi245 );
  xor      g04257 ( new_n4634 , new_n4509 , new_n4633 );
  nand     g04258 ( new_n4635 , pi051 , pi063 );
  nand     g04259 ( new_n4636 , pi108 , pi201 );
  xor      g04260 ( new_n4637 , new_n4635 , new_n4636 );
  xor      g04261 ( new_n4638 , new_n4508 , new_n4637 );
  xnor     g04262 ( new_n4639 , new_n4634 , new_n4638 );
  nand     g04263 ( new_n4640 , new_n4504 , new_n4511 );
  nand     g04264 ( new_n4641 , new_n4503 , new_n4512 );
  nand     g04265 ( new_n4642 , new_n4640 , new_n4641 );
  nand     g04266 ( new_n4643 , pi038 , pi107 );
  nand     g04267 ( new_n4644 , pi113 , pi171 );
  xor      g04268 ( new_n4645 , new_n4643 , new_n4644 );
  xor      g04269 ( new_n4646 , new_n4498 , new_n4645 );
  xor      g04270 ( new_n4647 , new_n4642 , new_n4646 );
  xor      g04271 ( new_n4648 , new_n4639 , new_n4647 );
  xor      g04272 ( new_n4649 , new_n4632 , new_n4648 );
  xor      g04273 ( new_n4650 , new_n4628 , new_n4649 );
  nand     g04274 ( new_n4651 , new_n4489 , new_n4490 );
  nand g04275 ( new_n4652 , new_n4521 , new_n4521 );
  nand     g04276 ( new_n4653 , new_n4491 , new_n4652 );
  nand     g04277 ( new_n4654 , new_n4651 , new_n4653 );
  xor      g04278 ( new_n4655 , new_n4650 , new_n4654 );
  xor      g04279 ( new_n4656 , new_n4627 , new_n4655 );
  nand g04280 ( new_n4657 , new_n4522 , new_n4522 );
  nor      g04281 ( new_n4658 , new_n4657 , new_n4554 );
  nor      g04282 ( new_n4659 , new_n4488 , new_n4555 );
  nor      g04283 ( new_n4660 , new_n4658 , new_n4659 );
  xor      g04284 ( new_n4661 , new_n4656 , new_n4660 );
  nor      g04285 ( new_n4662 , new_n4584 , new_n4588 );
  nor      g04286 ( new_n4663 , new_n4570 , new_n4573 );
  nor      g04287 ( new_n4664 , new_n4569 , new_n4574 );
  nor      g04288 ( new_n4665 , new_n4663 , new_n4664 );
  nand     g04289 ( new_n4666 , pi134 , pi238 );
  nand     g04290 ( new_n4667 , pi175 , pi193 );
  xor      g04291 ( new_n4668 , new_n4666 , new_n4667 );
  xor      g04292 ( new_n4669 , new_n4579 , new_n4668 );
  xor      g04293 ( new_n4670 , new_n4665 , new_n4669 );
  nand     g04294 ( new_n4671 , pi162 , pi200 );
  nand     g04295 ( new_n4672 , pi167 , pi179 );
  xor      g04296 ( new_n4673 , new_n4671 , new_n4672 );
  xor      g04297 ( new_n4674 , new_n4563 , new_n4673 );
  nand     g04298 ( new_n4675 , pi048 , pi149 );
  xor      g04299 ( new_n4676 , new_n4564 , new_n4675 );
  xnor     g04300 ( new_n4677 , new_n4674 , new_n4676 );
  xor      g04301 ( new_n4678 , new_n4670 , new_n4677 );
  nand g04302 ( new_n4679 , new_n4575 , new_n4575 );
  nor      g04303 ( new_n4680 , new_n4679 , new_n4581 );
  nor      g04304 ( new_n4681 , new_n4562 , new_n4582 );
  xor      g04305 ( new_n4682 , new_n4580 , new_n4681 );
  nor      g04306 ( new_n4683 , new_n4680 , new_n4682 );
  xor      g04307 ( new_n4684 , new_n4678 , new_n4683 );
  nand     g04308 ( new_n4685 , new_n4662 , new_n4684 );
  or       g04309 ( new_n4686 , new_n4662 , new_n4684 );
  nand     g04310 ( new_n4687 , new_n4685 , new_n4686 );
  nand     g04311 ( new_n4688 , new_n4590 , new_n4591 );
  nand g04312 ( new_n4689 , new_n4589 , new_n4589 );
  nand     g04313 ( new_n4690 , new_n4689 , new_n4592 );
  nand     g04314 ( new_n4691 , new_n4688 , new_n4690 );
  xnor     g04315 ( new_n4692 , new_n4687 , new_n4691 );
  xnor     g04316 ( new_n4693 , new_n4661 , new_n4692 );
  nand     g04317 ( new_n4694 , new_n4559 , new_n4593 );
  nand     g04318 ( new_n4695 , new_n4556 , new_n4594 );
  and      g04319 ( new_n4696 , new_n4694 , new_n4695 );
  xor      g04320 ( new_n4697 , new_n4693 , new_n4696 );
  xnor     g04321 ( po014 , new_n4598 , new_n4697 );
  nand     g04322 ( new_n4699 , pi085 , pi131 );
  nand     g04323 ( new_n4700 , pi052 , pi057 );
  nand     g04324 ( new_n4701 , pi131 , pi194 );
  nand     g04325 ( new_n4702 , new_n4700 , new_n4701 );
  nand     g04326 ( new_n4703 , pi077 , pi143 );
  xor      g04327 ( new_n4704 , new_n4700 , new_n4701 );
  nand     g04328 ( new_n4705 , new_n4703 , new_n4704 );
  nand     g04329 ( new_n4706 , new_n4702 , new_n4705 );
  nor      g04330 ( new_n4707 , new_n4699 , new_n4706 );
  nand     g04331 ( new_n4708 , pi057 , pi077 );
  nand     g04332 ( new_n4709 , pi052 , pi194 );
  nand     g04333 ( new_n4710 , pi133 , pi143 );
  xor      g04334 ( new_n4711 , new_n4709 , new_n4710 );
  xor      g04335 ( new_n4712 , new_n4708 , new_n4711 );
  xnor     g04336 ( new_n4713 , new_n4699 , new_n4706 );
  nor      g04337 ( new_n4714 , new_n4712 , new_n4713 );
  nor      g04338 ( new_n4715 , new_n4707 , new_n4714 );
  nand     g04339 ( new_n4716 , pi131 , pi180 );
  nand     g04340 ( new_n4717 , pi057 , pi133 );
  nand     g04341 ( new_n4718 , pi143 , pi189 );
  nand     g04342 ( new_n4719 , pi077 , pi194 );
  xor      g04343 ( new_n4720 , new_n4718 , new_n4719 );
  xor      g04344 ( new_n4721 , new_n4717 , new_n4720 );
  nand     g04345 ( new_n4722 , pi052 , pi085 );
  nand     g04346 ( new_n4723 , new_n4709 , new_n4710 );
  nand     g04347 ( new_n4724 , new_n4708 , new_n4711 );
  nand     g04348 ( new_n4725 , new_n4723 , new_n4724 );
  xor      g04349 ( new_n4726 , new_n4722 , new_n4725 );
  xor      g04350 ( new_n4727 , new_n4721 , new_n4726 );
  xor      g04351 ( new_n4728 , new_n4716 , new_n4727 );
  nand g04352 ( new_n4729 , new_n4728 , new_n4728 );
  xor      g04353 ( new_n4730 , new_n4715 , new_n4729 );
  xor      g04354 ( new_n4731 , new_n4703 , new_n4704 );
  nand g04355 ( new_n4732 , new_n4731 , new_n4731 );
  nand     g04356 ( new_n4733 , pi057 , pi131 );
  nand     g04357 ( new_n4734 , pi052 , pi143 );
  nor      g04358 ( new_n4735 , new_n4733 , new_n4734 );
  nand     g04359 ( new_n4736 , new_n4732 , new_n4735 );
  xnor     g04360 ( new_n4737 , new_n4712 , new_n4713 );
  nor      g04361 ( new_n4738 , new_n4736 , new_n4737 );
  xor      g04362 ( new_n4739 , new_n4730 , new_n4738 );
  nand     g04363 ( new_n4740 , pi051 , pi141 );
  nand     g04364 ( new_n4741 , pi042 , pi161 );
  nand     g04365 ( new_n4742 , pi108 , pi241 );
  xor      g04366 ( new_n4743 , new_n4741 , new_n4742 );
  xor      g04367 ( new_n4744 , new_n4740 , new_n4743 );
  nand     g04368 ( new_n4745 , pi007 , pi236 );
  nand     g04369 ( new_n4746 , pi042 , pi241 );
  nand     g04370 ( new_n4747 , pi108 , pi236 );
  nand     g04371 ( new_n4748 , new_n4746 , new_n4747 );
  nand     g04372 ( new_n4749 , pi051 , pi161 );
  xor      g04373 ( new_n4750 , new_n4746 , new_n4747 );
  nand     g04374 ( new_n4751 , new_n4749 , new_n4750 );
  nand     g04375 ( new_n4752 , new_n4748 , new_n4751 );
  xnor     g04376 ( new_n4753 , new_n4745 , new_n4752 );
  xnor     g04377 ( new_n4754 , new_n4744 , new_n4753 );
  xnor     g04378 ( new_n4755 , new_n4749 , new_n4750 );
  or       g04379 ( new_n4756 , new_n3609 , new_n4746 );
  nand g04380 ( new_n4757 , new_n4756 , new_n4756 );
  nand     g04381 ( new_n4758 , new_n4755 , new_n4757 );
  xor      g04382 ( new_n4759 , new_n4754 , new_n4758 );
  nand     g04383 ( new_n4760 , pi013 , pi188 );
  nand     g04384 ( new_n4761 , pi104 , pi178 );
  nand     g04385 ( new_n4762 , pi061 , pi212 );
  xor      g04386 ( new_n4763 , new_n4761 , new_n4762 );
  xor      g04387 ( new_n4764 , new_n4760 , new_n4763 );
  nand     g04388 ( new_n4765 , pi012 , pi213 );
  nand     g04389 ( new_n4766 , pi178 , pi212 );
  nand     g04390 ( new_n4767 , pi061 , pi213 );
  nand     g04391 ( new_n4768 , new_n4766 , new_n4767 );
  and      g04392 ( new_n4769 , pi104 , pi188 );
  xnor     g04393 ( new_n4770 , new_n4766 , new_n4767 );
  or       g04394 ( new_n4771 , new_n4769 , new_n4770 );
  nand     g04395 ( new_n4772 , new_n4768 , new_n4771 );
  xor      g04396 ( new_n4773 , new_n4765 , new_n4772 );
  xor      g04397 ( new_n4774 , new_n4764 , new_n4773 );
  xnor     g04398 ( new_n4775 , new_n4769 , new_n4770 );
  nor      g04399 ( new_n4776 , new_n3610 , new_n4766 );
  nand     g04400 ( new_n4777 , new_n4775 , new_n4776 );
  xor      g04401 ( new_n4778 , new_n4774 , new_n4777 );
  nand     g04402 ( new_n4779 , new_n4759 , new_n4778 );
  xor      g04403 ( new_n4780 , new_n4759 , new_n4778 );
  or       g04404 ( new_n4781 , new_n3609 , new_n3610 );
  nand     g04405 ( new_n4782 , pi042 , pi236 );
  nand     g04406 ( new_n4783 , pi051 , pi241 );
  nand     g04407 ( new_n4784 , new_n4782 , new_n4783 );
  nand     g04408 ( new_n4785 , new_n4756 , new_n4784 );
  nor      g04409 ( new_n4786 , new_n4781 , new_n4785 );
  xnor     g04410 ( new_n4787 , new_n4781 , new_n4785 );
  nand     g04411 ( new_n4788 , pi178 , pi213 );
  nand     g04412 ( new_n4789 , pi188 , pi212 );
  and      g04413 ( new_n4790 , new_n4788 , new_n4789 );
  or       g04414 ( new_n4791 , new_n4776 , new_n4790 );
  nor      g04415 ( new_n4792 , new_n4787 , new_n4791 );
  or       g04416 ( new_n4793 , new_n4786 , new_n4792 );
  xor      g04417 ( new_n4794 , new_n4775 , new_n4776 );
  nor      g04418 ( new_n4795 , new_n4793 , new_n4794 );
  xor      g04419 ( new_n4796 , new_n4755 , new_n4757 );
  xnor     g04420 ( new_n4797 , new_n4793 , new_n4794 );
  nor      g04421 ( new_n4798 , new_n4796 , new_n4797 );
  nor      g04422 ( new_n4799 , new_n4795 , new_n4798 );
  nand     g04423 ( new_n4800 , new_n4780 , new_n4799 );
  and      g04424 ( new_n4801 , new_n4779 , new_n4800 );
  nor      g04425 ( new_n4802 , new_n4754 , new_n4758 );
  nand     g04426 ( new_n4803 , pi118 , pi236 );
  nor      g04427 ( new_n4804 , new_n4745 , new_n4752 );
  nor      g04428 ( new_n4805 , new_n4744 , new_n4753 );
  nor      g04429 ( new_n4806 , new_n4804 , new_n4805 );
  xor      g04430 ( new_n4807 , new_n4803 , new_n4806 );
  nand     g04431 ( new_n4808 , pi108 , pi161 );
  nand     g04432 ( new_n4809 , pi042 , pi141 );
  nand     g04433 ( new_n4810 , pi051 , pi090 );
  xor      g04434 ( new_n4811 , new_n4809 , new_n4810 );
  xor      g04435 ( new_n4812 , new_n4808 , new_n4811 );
  nand     g04436 ( new_n4813 , pi007 , pi241 );
  nand     g04437 ( new_n4814 , new_n4741 , new_n4742 );
  nand     g04438 ( new_n4815 , new_n4740 , new_n4743 );
  nand     g04439 ( new_n4816 , new_n4814 , new_n4815 );
  xor      g04440 ( new_n4817 , new_n4813 , new_n4816 );
  xnor     g04441 ( new_n4818 , new_n4812 , new_n4817 );
  xor      g04442 ( new_n4819 , new_n4807 , new_n4818 );
  xnor     g04443 ( new_n4820 , new_n4802 , new_n4819 );
  nor      g04444 ( new_n4821 , new_n4774 , new_n4777 );
  nand     g04445 ( new_n4822 , pi144 , pi213 );
  nand     g04446 ( new_n4823 , new_n4765 , new_n4772 );
  nand     g04447 ( new_n4824 , new_n4764 , new_n4773 );
  nand     g04448 ( new_n4825 , new_n4823 , new_n4824 );
  xor      g04449 ( new_n4826 , new_n4822 , new_n4825 );
  nand     g04450 ( new_n4827 , pi112 , pi188 );
  nand     g04451 ( new_n4828 , pi061 , pi104 );
  nand     g04452 ( new_n4829 , pi013 , pi178 );
  xor      g04453 ( new_n4830 , new_n4828 , new_n4829 );
  xor      g04454 ( new_n4831 , new_n4827 , new_n4830 );
  nand     g04455 ( new_n4832 , pi012 , pi212 );
  nand     g04456 ( new_n4833 , new_n4761 , new_n4762 );
  nand     g04457 ( new_n4834 , new_n4760 , new_n4763 );
  nand     g04458 ( new_n4835 , new_n4833 , new_n4834 );
  xor      g04459 ( new_n4836 , new_n4832 , new_n4835 );
  xnor     g04460 ( new_n4837 , new_n4831 , new_n4836 );
  xor      g04461 ( new_n4838 , new_n4826 , new_n4837 );
  xor      g04462 ( new_n4839 , new_n4821 , new_n4838 );
  xor      g04463 ( new_n4840 , new_n4820 , new_n4839 );
  xor      g04464 ( new_n4841 , new_n4801 , new_n4840 );
  nand     g04465 ( new_n4842 , pi139 , pi162 );
  nand     g04466 ( new_n4843 , pi033 , pi208 );
  nand     g04467 ( new_n4844 , pi168 , pi179 );
  xor      g04468 ( new_n4845 , new_n4843 , new_n4844 );
  xor      g04469 ( new_n4846 , new_n4842 , new_n4845 );
  nand g04470 ( new_n4847 , new_n4846 , new_n4846 );
  nor      g04471 ( new_n4848 , new_n3608 , new_n4843 );
  nand     g04472 ( new_n4849 , new_n4847 , new_n4848 );
  nand     g04473 ( new_n4850 , pi179 , pi208 );
  nand     g04474 ( new_n4851 , pi035 , pi162 );
  nand     g04475 ( new_n4852 , pi033 , pi139 );
  xor      g04476 ( new_n4853 , new_n4851 , new_n4852 );
  xor      g04477 ( new_n4854 , new_n4850 , new_n4853 );
  nand     g04478 ( new_n4855 , pi048 , pi168 );
  nand     g04479 ( new_n4856 , new_n4843 , new_n4844 );
  nand     g04480 ( new_n4857 , new_n4842 , new_n4845 );
  nand     g04481 ( new_n4858 , new_n4856 , new_n4857 );
  xor      g04482 ( new_n4859 , new_n4855 , new_n4858 );
  xor      g04483 ( new_n4860 , new_n4854 , new_n4859 );
  nor      g04484 ( new_n4861 , new_n4849 , new_n4860 );
  nand     g04485 ( new_n4862 , pi139 , pi179 );
  nand     g04486 ( new_n4863 , pi033 , pi035 );
  nand     g04487 ( new_n4864 , pi015 , pi162 );
  xor      g04488 ( new_n4865 , new_n4863 , new_n4864 );
  xor      g04489 ( new_n4866 , new_n4862 , new_n4865 );
  nand     g04490 ( new_n4867 , pi048 , pi208 );
  nand     g04491 ( new_n4868 , new_n4851 , new_n4852 );
  nand     g04492 ( new_n4869 , new_n4850 , new_n4853 );
  nand     g04493 ( new_n4870 , new_n4868 , new_n4869 );
  xor      g04494 ( new_n4871 , new_n4867 , new_n4870 );
  xor      g04495 ( new_n4872 , new_n4866 , new_n4871 );
  nand     g04496 ( new_n4873 , pi168 , pi237 );
  nor      g04497 ( new_n4874 , new_n4855 , new_n4858 );
  nand g04498 ( new_n4875 , new_n4854 , new_n4854 );
  nand     g04499 ( new_n4876 , new_n4875 , new_n4859 );
  nand g04500 ( new_n4877 , new_n4876 , new_n4876 );
  nor      g04501 ( new_n4878 , new_n4874 , new_n4877 );
  xnor     g04502 ( new_n4879 , new_n4873 , new_n4878 );
  xnor     g04503 ( new_n4880 , new_n4872 , new_n4879 );
  xor      g04504 ( new_n4881 , new_n4861 , new_n4880 );
  xor      g04505 ( new_n4882 , new_n4780 , new_n4799 );
  xor      g04506 ( new_n4883 , new_n4849 , new_n4860 );
  and      g04507 ( new_n4884 , new_n4882 , new_n4883 );
  nor      g04508 ( new_n4885 , new_n4882 , new_n4883 );
  or       g04509 ( new_n4886 , new_n3608 , new_n3611 );
  nand     g04510 ( new_n4887 , pi033 , pi168 );
  nand     g04511 ( new_n4888 , pi162 , pi208 );
  and      g04512 ( new_n4889 , new_n4887 , new_n4888 );
  or       g04513 ( new_n4890 , new_n4848 , new_n4889 );
  nand     g04514 ( new_n4891 , new_n4886 , new_n4890 );
  xor      g04515 ( new_n4892 , new_n4787 , new_n4791 );
  xnor     g04516 ( new_n4893 , new_n4886 , new_n4890 );
  or       g04517 ( new_n4894 , new_n4892 , new_n4893 );
  nand     g04518 ( new_n4895 , new_n4891 , new_n4894 );
  xor      g04519 ( new_n4896 , new_n4846 , new_n4848 );
  nor      g04520 ( new_n4897 , new_n4895 , new_n4896 );
  xor      g04521 ( new_n4898 , new_n4895 , new_n4896 );
  xnor     g04522 ( new_n4899 , new_n4796 , new_n4797 );
  and      g04523 ( new_n4900 , new_n4898 , new_n4899 );
  nor      g04524 ( new_n4901 , new_n4897 , new_n4900 );
  nor      g04525 ( new_n4902 , new_n4885 , new_n4901 );
  nor      g04526 ( new_n4903 , new_n4884 , new_n4902 );
  xnor     g04527 ( new_n4904 , new_n4881 , new_n4903 );
  xnor     g04528 ( new_n4905 , new_n4841 , new_n4904 );
  xor      g04529 ( new_n4906 , new_n4739 , new_n4905 );
  or       g04530 ( new_n4907 , new_n4884 , new_n4885 );
  xor      g04531 ( new_n4908 , new_n4901 , new_n4907 );
  xor      g04532 ( new_n4909 , new_n4736 , new_n4737 );
  nor      g04533 ( new_n4910 , new_n4908 , new_n4909 );
  xor      g04534 ( new_n4911 , new_n4898 , new_n4899 );
  xor      g04535 ( new_n4912 , new_n4732 , new_n4735 );
  nand     g04536 ( new_n4913 , new_n4911 , new_n4912 );
  xor      g04537 ( new_n4914 , new_n4911 , new_n4912 );
  nor      g04538 ( new_n4915 , new_n3613 , new_n3614 );
  xor      g04539 ( new_n4916 , new_n4733 , new_n4734 );
  nor      g04540 ( new_n4917 , new_n4915 , new_n4916 );
  xor      g04541 ( new_n4918 , new_n4915 , new_n4916 );
  xor      g04542 ( new_n4919 , new_n4892 , new_n4893 );
  nand     g04543 ( new_n4920 , new_n4918 , new_n4919 );
  nand g04544 ( new_n4921 , new_n4920 , new_n4920 );
  nor      g04545 ( new_n4922 , new_n4917 , new_n4921 );
  nand     g04546 ( new_n4923 , new_n4914 , new_n4922 );
  nand     g04547 ( new_n4924 , new_n4913 , new_n4923 );
  xnor     g04548 ( new_n4925 , new_n4908 , new_n4909 );
  nor      g04549 ( new_n4926 , new_n4924 , new_n4925 );
  nor      g04550 ( new_n4927 , new_n4910 , new_n4926 );
  xor      g04551 ( po015 , new_n4906 , new_n4927 );
  nand     g04552 ( new_n4929 , pi060 , pi143 );
  nand     g04553 ( new_n4930 , pi020 , pi057 );
  nand     g04554 ( new_n4931 , pi160 , pi194 );
  xor      g04555 ( new_n4932 , new_n4930 , new_n4931 );
  xor      g04556 ( new_n4933 , new_n4929 , new_n4932 );
  nand     g04557 ( new_n4934 , pi143 , pi160 );
  or       g04558 ( new_n4935 , new_n4930 , new_n4934 );
  xor      g04559 ( new_n4936 , new_n4933 , new_n4935 );
  nand g04560 ( new_n4937 , new_n4936 , new_n4936 );
  nand     g04561 ( new_n4938 , pi142 , pi188 );
  nand     g04562 ( new_n4939 , pi051 , pi087 );
  xnor     g04563 ( new_n4940 , new_n4938 , new_n4939 );
  nand     g04564 ( new_n4941 , pi138 , pi162 );
  xor      g04565 ( new_n4942 , new_n4940 , new_n4941 );
  nand g04566 ( new_n4943 , new_n4942 , new_n4942 );
  or       g04567 ( new_n4944 , new_n4934 , new_n4943 );
  nand     g04568 ( new_n4945 , pi057 , pi160 );
  nand     g04569 ( new_n4946 , pi020 , pi143 );
  nand     g04570 ( new_n4947 , new_n4945 , new_n4946 );
  nand     g04571 ( new_n4948 , new_n4935 , new_n4947 );
  nor      g04572 ( new_n4949 , new_n4944 , new_n4948 );
  xnor     g04573 ( new_n4950 , new_n4944 , new_n4948 );
  nor      g04574 ( new_n4951 , new_n4938 , new_n4939 );
  nand     g04575 ( new_n4952 , pi142 , pi178 );
  nand     g04576 ( new_n4953 , pi071 , pi188 );
  xor      g04577 ( new_n4954 , new_n4952 , new_n4953 );
  nand     g04578 ( new_n4955 , pi042 , pi087 );
  nand     g04579 ( new_n4956 , pi051 , pi219 );
  xor      g04580 ( new_n4957 , new_n4955 , new_n4956 );
  xnor     g04581 ( new_n4958 , new_n4954 , new_n4957 );
  xnor     g04582 ( new_n4959 , new_n4951 , new_n4958 );
  nor      g04583 ( new_n4960 , new_n4940 , new_n4941 );
  nand     g04584 ( new_n4961 , pi162 , pi182 );
  nand     g04585 ( new_n4962 , pi033 , pi138 );
  xor      g04586 ( new_n4963 , new_n4961 , new_n4962 );
  xnor     g04587 ( new_n4964 , new_n4960 , new_n4963 );
  xor      g04588 ( new_n4965 , new_n4959 , new_n4964 );
  nor      g04589 ( new_n4966 , new_n4950 , new_n4965 );
  nor      g04590 ( new_n4967 , new_n4949 , new_n4966 );
  nand     g04591 ( new_n4968 , new_n4937 , new_n4967 );
  xor      g04592 ( new_n4969 , new_n4937 , new_n4967 );
  nor      g04593 ( new_n4970 , new_n4961 , new_n4962 );
  nand     g04594 ( new_n4971 , pi041 , pi162 );
  nand     g04595 ( new_n4972 , pi033 , pi182 );
  nand     g04596 ( new_n4973 , pi138 , pi179 );
  xor      g04597 ( new_n4974 , new_n4972 , new_n4973 );
  xnor     g04598 ( new_n4975 , new_n4971 , new_n4974 );
  xor      g04599 ( new_n4976 , new_n4970 , new_n4975 );
  and      g04600 ( new_n4977 , pi042 , pi219 );
  and      g04601 ( new_n4978 , new_n4939 , new_n4977 );
  nand     g04602 ( new_n4979 , pi087 , pi108 );
  nand     g04603 ( new_n4980 , pi051 , pi102 );
  nor      g04604 ( new_n4981 , new_n4979 , new_n4980 );
  nand     g04605 ( new_n4982 , new_n4979 , new_n4980 );
  nand g04606 ( new_n4983 , new_n4982 , new_n4982 );
  nor      g04607 ( new_n4984 , new_n4981 , new_n4983 );
  nor      g04608 ( new_n4985 , new_n4978 , new_n4984 );
  and      g04609 ( new_n4986 , new_n4982 , new_n4978 );
  nor      g04610 ( new_n4987 , new_n4985 , new_n4986 );
  nor      g04611 ( new_n4988 , new_n4954 , new_n4957 );
  nor      g04612 ( new_n4989 , new_n4951 , new_n4958 );
  nor      g04613 ( new_n4990 , new_n4988 , new_n4989 );
  nand g04614 ( new_n4991 , pi071 , pi071 );
  nor      g04615 ( new_n4992 , new_n4991 , new_n953 );
  nand     g04616 ( new_n4993 , new_n4938 , new_n4992 );
  nand     g04617 ( new_n4994 , pi169 , pi188 );
  nand     g04618 ( new_n4995 , pi061 , pi142 );
  nor      g04619 ( new_n4996 , new_n4994 , new_n4995 );
  and      g04620 ( new_n4997 , new_n4994 , new_n4995 );
  or       g04621 ( new_n4998 , new_n4996 , new_n4997 );
  and      g04622 ( new_n4999 , new_n4993 , new_n4998 );
  nor      g04623 ( new_n5000 , new_n4997 , new_n4993 );
  nor      g04624 ( new_n5001 , new_n4999 , new_n5000 );
  xor      g04625 ( new_n5002 , new_n4990 , new_n5001 );
  xor      g04626 ( new_n5003 , new_n4987 , new_n5002 );
  xor      g04627 ( new_n5004 , new_n4976 , new_n5003 );
  nor      g04628 ( new_n5005 , new_n4960 , new_n4963 );
  nor      g04629 ( new_n5006 , new_n4959 , new_n4964 );
  nor      g04630 ( new_n5007 , new_n5005 , new_n5006 );
  xnor     g04631 ( new_n5008 , new_n5004 , new_n5007 );
  nand     g04632 ( new_n5009 , new_n4969 , new_n5008 );
  nand     g04633 ( new_n5010 , new_n4968 , new_n5009 );
  or       g04634 ( new_n5011 , new_n4933 , new_n4935 );
  nand     g04635 ( new_n5012 , pi020 , pi194 );
  nand     g04636 ( new_n5013 , pi143 , pi223 );
  nand     g04637 ( new_n5014 , pi057 , pi060 );
  xor      g04638 ( new_n5015 , new_n5013 , new_n5014 );
  xor      g04639 ( new_n5016 , new_n5012 , new_n5015 );
  nand     g04640 ( new_n5017 , pi085 , pi160 );
  nand     g04641 ( new_n5018 , new_n4930 , new_n4931 );
  nand     g04642 ( new_n5019 , new_n4929 , new_n4932 );
  nand     g04643 ( new_n5020 , new_n5018 , new_n5019 );
  xor      g04644 ( new_n5021 , new_n5017 , new_n5020 );
  xor      g04645 ( new_n5022 , new_n5016 , new_n5021 );
  xor      g04646 ( new_n5023 , new_n5011 , new_n5022 );
  nand g04647 ( new_n5024 , new_n5023 , new_n5023 );
  xor      g04648 ( new_n5025 , new_n5010 , new_n5024 );
  nand     g04649 ( new_n5026 , new_n4976 , new_n5003 );
  nand     g04650 ( new_n5027 , new_n5004 , new_n5007 );
  nand     g04651 ( new_n5028 , new_n5026 , new_n5027 );
  nand     g04652 ( new_n5029 , new_n4970 , new_n4975 );
  nand     g04653 ( new_n5030 , pi179 , pi182 );
  nand     g04654 ( new_n5031 , pi033 , pi041 );
  nand     g04655 ( new_n5032 , pi162 , pi216 );
  xor      g04656 ( new_n5033 , new_n5031 , new_n5032 );
  xor      g04657 ( new_n5034 , new_n5030 , new_n5033 );
  nand     g04658 ( new_n5035 , pi048 , pi138 );
  nand     g04659 ( new_n5036 , new_n4972 , new_n4973 );
  nand     g04660 ( new_n5037 , new_n4971 , new_n4974 );
  nand     g04661 ( new_n5038 , new_n5036 , new_n5037 );
  xor      g04662 ( new_n5039 , new_n5035 , new_n5038 );
  xor      g04663 ( new_n5040 , new_n5034 , new_n5039 );
  xnor     g04664 ( new_n5041 , new_n5029 , new_n5040 );
  xor      g04665 ( new_n5042 , new_n5028 , new_n5041 );
  nand     g04666 ( new_n5043 , new_n4992 , new_n4999 );
  nand     g04667 ( new_n5044 , pi123 , pi188 );
  nand     g04668 ( new_n5045 , pi061 , pi071 );
  nand     g04669 ( new_n5046 , pi169 , pi178 );
  xor      g04670 ( new_n5047 , new_n5045 , new_n5046 );
  xor      g04671 ( new_n5048 , new_n5044 , new_n5047 );
  nor      g04672 ( new_n5049 , new_n4996 , new_n4992 );
  or       g04673 ( new_n5050 , new_n4997 , new_n5049 );
  nand     g04674 ( new_n5051 , pi012 , pi142 );
  xnor     g04675 ( new_n5052 , new_n5050 , new_n5051 );
  xnor     g04676 ( new_n5053 , new_n5048 , new_n5052 );
  xnor     g04677 ( new_n5054 , new_n5043 , new_n5053 );
  and      g04678 ( new_n5055 , new_n4977 , new_n4985 );
  nand     g04679 ( new_n5056 , pi001 , pi051 );
  nand     g04680 ( new_n5057 , pi108 , pi219 );
  nand     g04681 ( new_n5058 , pi042 , pi102 );
  xor      g04682 ( new_n5059 , new_n5057 , new_n5058 );
  xor      g04683 ( new_n5060 , new_n5056 , new_n5059 );
  nand     g04684 ( new_n5061 , pi007 , pi087 );
  nor      g04685 ( new_n5062 , new_n4981 , new_n4977 );
  or       g04686 ( new_n5063 , new_n4983 , new_n5062 );
  xnor     g04687 ( new_n5064 , new_n5061 , new_n5063 );
  xnor     g04688 ( new_n5065 , new_n5060 , new_n5064 );
  xor      g04689 ( new_n5066 , new_n5055 , new_n5065 );
  xnor     g04690 ( new_n5067 , new_n5054 , new_n5066 );
  nand     g04691 ( new_n5068 , new_n4990 , new_n5001 );
  nand     g04692 ( new_n5069 , new_n4987 , new_n5002 );
  and      g04693 ( new_n5070 , new_n5068 , new_n5069 );
  xor      g04694 ( new_n5071 , new_n5067 , new_n5070 );
  xnor     g04695 ( new_n5072 , new_n5042 , new_n5071 );
  xor      g04696 ( po016 , new_n5025 , new_n5072 );
  nand     g04697 ( new_n5074 , pi132 , pi175 );
  nand     g04698 ( new_n5075 , pi107 , pi109 );
  nand     g04699 ( new_n5076 , pi163 , pi226 );
  xnor     g04700 ( new_n5077 , new_n5075 , new_n5076 );
  or       g04701 ( new_n5078 , new_n5074 , new_n5077 );
  nand     g04702 ( new_n5079 , pi134 , pi186 );
  or       g04703 ( new_n5080 , new_n5074 , new_n5079 );
  nand     g04704 ( new_n5081 , pi175 , pi186 );
  nand     g04705 ( new_n5082 , pi132 , pi134 );
  nand     g04706 ( new_n5083 , new_n5081 , new_n5082 );
  nand     g04707 ( new_n5084 , new_n5080 , new_n5083 );
  xor      g04708 ( new_n5085 , new_n5078 , new_n5084 );
  nand     g04709 ( new_n5086 , pi014 , pi171 );
  nor      g04710 ( new_n5087 , new_n5075 , new_n5086 );
  nand g04711 ( new_n5088 , pi107 , pi107 );
  nor      g04712 ( new_n5089 , new_n3916 , new_n5088 );
  nor      g04713 ( new_n5090 , new_n4033 , new_n2156 );
  nor      g04714 ( new_n5091 , new_n5089 , new_n5090 );
  or       g04715 ( new_n5092 , new_n5087 , new_n5091 );
  or       g04716 ( new_n5093 , new_n5075 , new_n5076 );
  nand     g04717 ( new_n5094 , pi148 , pi207 );
  or       g04718 ( new_n5095 , new_n5076 , new_n5094 );
  nand     g04719 ( new_n5096 , pi148 , pi226 );
  nand     g04720 ( new_n5097 , pi163 , pi207 );
  nand     g04721 ( new_n5098 , new_n5096 , new_n5097 );
  nand     g04722 ( new_n5099 , new_n5095 , new_n5098 );
  xnor     g04723 ( new_n5100 , new_n5093 , new_n5099 );
  xnor     g04724 ( new_n5101 , new_n5092 , new_n5100 );
  xor      g04725 ( new_n5102 , new_n5085 , new_n5101 );
  nand     g04726 ( new_n5103 , pi029 , pi103 );
  xnor     g04727 ( new_n5104 , new_n5074 , new_n5077 );
  nor      g04728 ( new_n5105 , new_n5103 , new_n5104 );
  nand     g04729 ( new_n5106 , pi029 , pi117 );
  nand     g04730 ( new_n5107 , pi069 , pi103 );
  xor      g04731 ( new_n5108 , new_n5106 , new_n5107 );
  xor      g04732 ( new_n5109 , new_n5105 , new_n5108 );
  nand g04733 ( new_n5110 , new_n5109 , new_n5109 );
  xor      g04734 ( po017 , new_n5102 , new_n5110 );
  xor      g04735 ( po018 , new_n3205 , new_n3206 );
  nand     g04736 ( new_n5113 , pi025 , pi213 );
  nand     g04737 ( new_n5114 , pi055 , pi212 );
  nand     g04738 ( new_n5115 , new_n3351 , new_n3352 );
  nand     g04739 ( new_n5116 , new_n3350 , new_n3353 );
  nand     g04740 ( new_n5117 , new_n5115 , new_n5116 );
  nand     g04741 ( new_n5118 , new_n5114 , new_n5117 );
  nand     g04742 ( new_n5119 , pi112 , pi226 );
  nand     g04743 ( new_n5120 , pi013 , pi207 );
  nand     g04744 ( new_n5121 , pi066 , pi104 );
  xor      g04745 ( new_n5122 , new_n5120 , new_n5121 );
  xor      g04746 ( new_n5123 , new_n5119 , new_n5122 );
  xor      g04747 ( new_n5124 , new_n5114 , new_n5117 );
  nand     g04748 ( new_n5125 , new_n5123 , new_n5124 );
  nand     g04749 ( new_n5126 , new_n5118 , new_n5125 );
  nand     g04750 ( new_n5127 , pi055 , pi104 );
  nand     g04751 ( new_n5128 , pi002 , pi212 );
  nand     g04752 ( new_n5129 , new_n5127 , new_n5128 );
  nand     g04753 ( new_n5130 , pi002 , pi104 );
  nor      g04754 ( new_n5131 , new_n5114 , new_n5130 );
  nand g04755 ( new_n5132 , new_n5131 , new_n5131 );
  nand     g04756 ( new_n5133 , new_n5129 , new_n5132 );
  nand     g04757 ( new_n5134 , pi013 , pi066 );
  nand     g04758 ( new_n5135 , new_n5120 , new_n5121 );
  nand     g04759 ( new_n5136 , new_n5119 , new_n5122 );
  nand     g04760 ( new_n5137 , new_n5135 , new_n5136 );
  nand     g04761 ( new_n5138 , pi105 , pi226 );
  nand     g04762 ( new_n5139 , pi112 , pi207 );
  nand     g04763 ( new_n5140 , new_n5138 , new_n5139 );
  nand     g04764 ( new_n5141 , pi105 , pi207 );
  or       g04765 ( new_n5142 , new_n5119 , new_n5141 );
  nand     g04766 ( new_n5143 , new_n5140 , new_n5142 );
  xor      g04767 ( new_n5144 , new_n5137 , new_n5143 );
  xor      g04768 ( new_n5145 , new_n5134 , new_n5144 );
  xor      g04769 ( new_n5146 , new_n5133 , new_n5145 );
  nand g04770 ( new_n5147 , new_n5146 , new_n5146 );
  xor      g04771 ( new_n5148 , new_n5126 , new_n5147 );
  nand     g04772 ( new_n5149 , pi002 , pi213 );
  nand     g04773 ( new_n5150 , new_n3355 , new_n3358 );
  nand g04774 ( new_n5151 , new_n5150 , new_n5150 );
  and      g04775 ( new_n5152 , new_n3354 , new_n3359 );
  nor      g04776 ( new_n5153 , new_n5151 , new_n5152 );
  nand g04777 ( new_n5154 , new_n5153 , new_n5153 );
  nor      g04778 ( new_n5155 , new_n5149 , new_n5154 );
  xor      g04779 ( new_n5156 , new_n5123 , new_n5124 );
  xor      g04780 ( new_n5157 , new_n5149 , new_n5153 );
  nor      g04781 ( new_n5158 , new_n5156 , new_n5157 );
  nor      g04782 ( new_n5159 , new_n5155 , new_n5158 );
  xor      g04783 ( new_n5160 , new_n5148 , new_n5159 );
  xnor     g04784 ( new_n5161 , new_n5113 , new_n5160 );
  nor      g04785 ( new_n5162 , new_n3349 , new_n3360 );
  xor      g04786 ( new_n5163 , new_n5156 , new_n5157 );
  nand     g04787 ( new_n5164 , new_n5162 , new_n5163 );
  xnor     g04788 ( new_n5165 , new_n5161 , new_n5164 );
  nand     g04789 ( new_n5166 , pi050 , pi236 );
  nand     g04790 ( new_n5167 , pi161 , pi173 );
  nand     g04791 ( new_n5168 , pi090 , pi109 );
  nand     g04792 ( new_n5169 , pi014 , pi141 );
  xor      g04793 ( new_n5170 , new_n5168 , new_n5169 );
  xor      g04794 ( new_n5171 , new_n5167 , new_n5170 );
  nand     g04795 ( new_n5172 , pi230 , pi241 );
  nand     g04796 ( new_n5173 , new_n3340 , new_n3341 );
  nand     g04797 ( new_n5174 , new_n3339 , new_n3342 );
  nand     g04798 ( new_n5175 , new_n5173 , new_n5174 );
  xor      g04799 ( new_n5176 , new_n5172 , new_n5175 );
  xor      g04800 ( new_n5177 , new_n5171 , new_n5176 );
  nor      g04801 ( new_n5178 , new_n5166 , new_n5177 );
  nor      g04802 ( new_n5179 , new_n3335 , new_n3337 );
  nand     g04803 ( new_n5180 , new_n3338 , new_n3344 );
  nand g04804 ( new_n5181 , new_n5180 , new_n5180 );
  nor      g04805 ( new_n5182 , new_n5179 , new_n5181 );
  xnor     g04806 ( new_n5183 , new_n5166 , new_n5177 );
  nor      g04807 ( new_n5184 , new_n5182 , new_n5183 );
  nor      g04808 ( new_n5185 , new_n5178 , new_n5184 );
  nand     g04809 ( new_n5186 , new_n5172 , new_n5175 );
  nand     g04810 ( new_n5187 , new_n5171 , new_n5176 );
  nand     g04811 ( new_n5188 , new_n5186 , new_n5187 );
  nand     g04812 ( new_n5189 , pi161 , pi230 );
  nand     g04813 ( new_n5190 , pi050 , pi241 );
  and      g04814 ( new_n5191 , new_n5189 , new_n5190 );
  nand     g04815 ( new_n5192 , pi050 , pi161 );
  nor      g04816 ( new_n5193 , new_n5172 , new_n5192 );
  or       g04817 ( new_n5194 , new_n5191 , new_n5193 );
  nand     g04818 ( new_n5195 , new_n5168 , new_n5169 );
  nand     g04819 ( new_n5196 , new_n5167 , new_n5170 );
  nand     g04820 ( new_n5197 , new_n5195 , new_n5196 );
  nand     g04821 ( new_n5198 , pi141 , pi173 );
  nand     g04822 ( new_n5199 , pi014 , pi090 );
  nand     g04823 ( new_n5200 , pi047 , pi109 );
  nand     g04824 ( new_n5201 , new_n5199 , new_n5200 );
  nand     g04825 ( new_n5202 , pi014 , pi047 );
  nor      g04826 ( new_n5203 , new_n5168 , new_n5202 );
  nand g04827 ( new_n5204 , new_n5203 , new_n5203 );
  nand     g04828 ( new_n5205 , new_n5201 , new_n5204 );
  xor      g04829 ( new_n5206 , new_n5198 , new_n5205 );
  xor      g04830 ( new_n5207 , new_n5197 , new_n5206 );
  xor      g04831 ( new_n5208 , new_n5194 , new_n5207 );
  xor      g04832 ( new_n5209 , new_n5188 , new_n5208 );
  xor      g04833 ( new_n5210 , new_n5185 , new_n5209 );
  nand     g04834 ( new_n5211 , pi236 , pi253 );
  nand     g04835 ( new_n5212 , new_n3277 , new_n3345 );
  xor      g04836 ( new_n5213 , new_n5182 , new_n5183 );
  nand g04837 ( new_n5214 , new_n5213 , new_n5213 );
  nor      g04838 ( new_n5215 , new_n5212 , new_n5214 );
  xor      g04839 ( new_n5216 , new_n5211 , new_n5215 );
  xor      g04840 ( new_n5217 , new_n5210 , new_n5216 );
  nor      g04841 ( new_n5218 , new_n5165 , new_n5217 );
  xor      g04842 ( new_n5219 , new_n5165 , new_n5217 );
  xor      g04843 ( new_n5220 , new_n5212 , new_n5213 );
  xnor     g04844 ( new_n5221 , new_n5162 , new_n5163 );
  nor      g04845 ( new_n5222 , new_n5220 , new_n5221 );
  nor      g04846 ( new_n5223 , new_n3334 , new_n3364 );
  or       g04847 ( new_n5224 , new_n3363 , new_n5223 );
  xnor     g04848 ( new_n5225 , new_n5220 , new_n5221 );
  nor      g04849 ( new_n5226 , new_n5224 , new_n5225 );
  or       g04850 ( new_n5227 , new_n5222 , new_n5226 );
  and      g04851 ( new_n5228 , new_n5219 , new_n5227 );
  nor      g04852 ( new_n5229 , new_n5218 , new_n5228 );
  nor      g04853 ( new_n5230 , new_n5113 , new_n5160 );
  nor      g04854 ( new_n5231 , new_n5161 , new_n5164 );
  nor      g04855 ( new_n5232 , new_n5230 , new_n5231 );
  nand g04856 ( new_n5233 , new_n5148 , new_n5148 );
  nor      g04857 ( new_n5234 , new_n5233 , new_n5159 );
  nor      g04858 ( new_n5235 , new_n5126 , new_n5147 );
  nand     g04859 ( new_n5236 , new_n5131 , new_n5235 );
  or       g04860 ( new_n5237 , new_n5133 , new_n5145 );
  nand     g04861 ( new_n5238 , new_n5132 , new_n5237 );
  or       g04862 ( new_n5239 , new_n5235 , new_n5238 );
  nand     g04863 ( new_n5240 , new_n5236 , new_n5239 );
  nand     g04864 ( new_n5241 , pi013 , pi055 );
  xnor     g04865 ( new_n5242 , new_n5142 , new_n5241 );
  nand     g04866 ( new_n5243 , pi183 , pi226 );
  nand     g04867 ( new_n5244 , pi066 , pi112 );
  xor      g04868 ( new_n5245 , new_n5243 , new_n5244 );
  xor      g04869 ( new_n5246 , new_n5141 , new_n5245 );
  xor      g04870 ( new_n5247 , new_n5242 , new_n5246 );
  nand     g04871 ( new_n5248 , new_n5137 , new_n5143 );
  nand     g04872 ( new_n5249 , new_n5134 , new_n5144 );
  nand     g04873 ( new_n5250 , new_n5248 , new_n5249 );
  nand     g04874 ( new_n5251 , pi025 , pi212 );
  nand     g04875 ( new_n5252 , pi213 , pi239 );
  xor      g04876 ( new_n5253 , new_n5251 , new_n5252 );
  xnor     g04877 ( new_n5254 , new_n5130 , new_n5253 );
  xor      g04878 ( new_n5255 , new_n5250 , new_n5254 );
  xor      g04879 ( new_n5256 , new_n5247 , new_n5255 );
  nand g04880 ( new_n5257 , new_n5256 , new_n5256 );
  xor      g04881 ( new_n5258 , new_n5240 , new_n5257 );
  xor      g04882 ( new_n5259 , new_n5234 , new_n5258 );
  xnor     g04883 ( new_n5260 , new_n5232 , new_n5259 );
  nor      g04884 ( new_n5261 , new_n5185 , new_n5209 );
  nand     g04885 ( new_n5262 , pi141 , pi230 );
  xor      g04886 ( new_n5263 , new_n5203 , new_n5262 );
  nand     g04887 ( new_n5264 , pi090 , pi173 );
  nand     g04888 ( new_n5265 , pi018 , pi109 );
  xor      g04889 ( new_n5266 , new_n5264 , new_n5265 );
  xor      g04890 ( new_n5267 , new_n5202 , new_n5266 );
  xnor     g04891 ( new_n5268 , new_n5263 , new_n5267 );
  nand     g04892 ( new_n5269 , new_n5198 , new_n5205 );
  nand     g04893 ( new_n5270 , new_n5197 , new_n5206 );
  nand     g04894 ( new_n5271 , new_n5269 , new_n5270 );
  nand     g04895 ( new_n5272 , pi241 , pi253 );
  nand     g04896 ( new_n5273 , pi074 , pi236 );
  xor      g04897 ( new_n5274 , new_n5272 , new_n5273 );
  xor      g04898 ( new_n5275 , new_n5192 , new_n5274 );
  xor      g04899 ( new_n5276 , new_n5271 , new_n5275 );
  xor      g04900 ( new_n5277 , new_n5268 , new_n5276 );
  nor      g04901 ( new_n5278 , new_n5194 , new_n5207 );
  nand g04902 ( new_n5279 , new_n5208 , new_n5208 );
  nor      g04903 ( new_n5280 , new_n5188 , new_n5279 );
  xor      g04904 ( new_n5281 , new_n5193 , new_n5280 );
  nor      g04905 ( new_n5282 , new_n5278 , new_n5281 );
  xor      g04906 ( new_n5283 , new_n5277 , new_n5282 );
  xor      g04907 ( new_n5284 , new_n5261 , new_n5283 );
  nand g04908 ( new_n5285 , new_n5211 , new_n5211 );
  nor      g04909 ( new_n5286 , new_n5285 , new_n5215 );
  nor      g04910 ( new_n5287 , new_n5210 , new_n5216 );
  nor      g04911 ( new_n5288 , new_n5286 , new_n5287 );
  xnor     g04912 ( new_n5289 , new_n5284 , new_n5288 );
  xor      g04913 ( new_n5290 , new_n5260 , new_n5289 );
  xor      g04914 ( new_n5291 , new_n5229 , new_n5290 );
  nand     g04915 ( new_n5292 , pi168 , pi199 );
  nand     g04916 ( new_n5293 , pi058 , pi139 );
  nand     g04917 ( new_n5294 , pi015 , pi132 );
  nand     g04918 ( new_n5295 , pi035 , pi186 );
  xor      g04919 ( new_n5296 , new_n5294 , new_n5295 );
  xor      g04920 ( new_n5297 , new_n5293 , new_n5296 );
  nand     g04921 ( new_n5298 , pi208 , pi211 );
  nand     g04922 ( new_n5299 , new_n3318 , new_n3319 );
  nand     g04923 ( new_n5300 , new_n3317 , new_n3320 );
  nand     g04924 ( new_n5301 , new_n5299 , new_n5300 );
  xor      g04925 ( new_n5302 , new_n5298 , new_n5301 );
  xor      g04926 ( new_n5303 , new_n5297 , new_n5302 );
  nor      g04927 ( new_n5304 , new_n5292 , new_n5303 );
  nor      g04928 ( new_n5305 , new_n3322 , new_n3325 );
  nor      g04929 ( new_n5306 , new_n3321 , new_n3327 );
  nor      g04930 ( new_n5307 , new_n5305 , new_n5306 );
  xor      g04931 ( new_n5308 , new_n5292 , new_n5303 );
  nand g04932 ( new_n5309 , new_n5308 , new_n5308 );
  nor      g04933 ( new_n5310 , new_n5307 , new_n5309 );
  nor      g04934 ( new_n5311 , new_n5304 , new_n5310 );
  nand     g04935 ( new_n5312 , pi139 , pi211 );
  nand     g04936 ( new_n5313 , pi199 , pi208 );
  and      g04937 ( new_n5314 , new_n5312 , new_n5313 );
  nand     g04938 ( new_n5315 , pi139 , pi199 );
  nor      g04939 ( new_n5316 , new_n5298 , new_n5315 );
  or       g04940 ( new_n5317 , new_n5314 , new_n5316 );
  nand     g04941 ( new_n5318 , new_n5294 , new_n5295 );
  nand     g04942 ( new_n5319 , new_n5293 , new_n5296 );
  nand     g04943 ( new_n5320 , new_n5318 , new_n5319 );
  nand     g04944 ( new_n5321 , pi035 , pi058 );
  nand     g04945 ( new_n5322 , pi015 , pi186 );
  nand     g04946 ( new_n5323 , pi132 , pi204 );
  nand     g04947 ( new_n5324 , new_n5322 , new_n5323 );
  nand     g04948 ( new_n5325 , pi186 , pi204 );
  nor      g04949 ( new_n5326 , new_n5294 , new_n5325 );
  nand g04950 ( new_n5327 , new_n5326 , new_n5326 );
  nand     g04951 ( new_n5328 , new_n5324 , new_n5327 );
  xor      g04952 ( new_n5329 , new_n5321 , new_n5328 );
  xor      g04953 ( new_n5330 , new_n5320 , new_n5329 );
  xor      g04954 ( new_n5331 , new_n5317 , new_n5330 );
  nand     g04955 ( new_n5332 , new_n5298 , new_n5301 );
  nand     g04956 ( new_n5333 , new_n5297 , new_n5302 );
  nand     g04957 ( new_n5334 , new_n5332 , new_n5333 );
  xor      g04958 ( new_n5335 , new_n5331 , new_n5334 );
  nor      g04959 ( new_n5336 , new_n5311 , new_n5335 );
  nand g04960 ( new_n5337 , new_n5336 , new_n5336 );
  nand     g04961 ( new_n5338 , new_n5321 , new_n5328 );
  nand     g04962 ( new_n5339 , new_n5320 , new_n5329 );
  nand     g04963 ( new_n5340 , new_n5338 , new_n5339 );
  nand g04964 ( new_n5341 , new_n5315 , new_n5315 );
  nand     g04965 ( new_n5342 , pi195 , pi208 );
  and      g04966 ( new_n5343 , pi168 , pi218 );
  xor      g04967 ( new_n5344 , new_n5342 , new_n5343 );
  xor      g04968 ( new_n5345 , new_n5341 , new_n5344 );
  xor      g04969 ( new_n5346 , new_n5340 , new_n5345 );
  nand     g04970 ( new_n5347 , pi132 , pi146 );
  nand     g04971 ( new_n5348 , pi015 , pi058 );
  xor      g04972 ( new_n5349 , new_n5347 , new_n5348 );
  xor      g04973 ( new_n5350 , new_n5325 , new_n5349 );
  nand     g04974 ( new_n5351 , pi035 , pi211 );
  xor      g04975 ( new_n5352 , new_n5326 , new_n5351 );
  xor      g04976 ( new_n5353 , new_n5350 , new_n5352 );
  nand g04977 ( new_n5354 , new_n5353 , new_n5353 );
  xor      g04978 ( new_n5355 , new_n5346 , new_n5354 );
  nor      g04979 ( new_n5356 , new_n5317 , new_n5330 );
  nand g04980 ( new_n5357 , new_n5334 , new_n5334 );
  nand     g04981 ( new_n5358 , new_n5331 , new_n5357 );
  xor      g04982 ( new_n5359 , new_n5316 , new_n5358 );
  nand g04983 ( new_n5360 , new_n5359 , new_n5359 );
  nor      g04984 ( new_n5361 , new_n5356 , new_n5360 );
  xor      g04985 ( new_n5362 , new_n5355 , new_n5361 );
  nand g04986 ( new_n5363 , new_n5362 , new_n5362 );
  nand     g04987 ( new_n5364 , pi168 , pi195 );
  nand g04988 ( new_n5365 , new_n3328 , new_n3328 );
  nor      g04989 ( new_n5366 , new_n3316 , new_n5365 );
  xor      g04990 ( new_n5367 , new_n5307 , new_n5309 );
  nand     g04991 ( new_n5368 , new_n5366 , new_n5367 );
  nand     g04992 ( new_n5369 , new_n5364 , new_n5368 );
  xor      g04993 ( new_n5370 , new_n5364 , new_n5368 );
  xnor     g04994 ( new_n5371 , new_n5311 , new_n5335 );
  nand     g04995 ( new_n5372 , new_n5370 , new_n5371 );
  nand     g04996 ( new_n5373 , new_n5369 , new_n5372 );
  xor      g04997 ( new_n5374 , new_n5363 , new_n5373 );
  xor      g04998 ( new_n5375 , new_n5337 , new_n5374 );
  xnor     g04999 ( new_n5376 , new_n5291 , new_n5375 );
  xor      g05000 ( new_n5377 , new_n5370 , new_n5371 );
  xnor     g05001 ( new_n5378 , new_n5219 , new_n5227 );
  nor      g05002 ( new_n5379 , new_n5377 , new_n5378 );
  xor      g05003 ( new_n5380 , new_n5366 , new_n5367 );
  nand g05004 ( new_n5381 , new_n5380 , new_n5380 );
  xnor     g05005 ( new_n5382 , new_n5224 , new_n5225 );
  nor      g05006 ( new_n5383 , new_n5381 , new_n5382 );
  nand     g05007 ( new_n5384 , new_n3314 , new_n3329 );
  nand     g05008 ( new_n5385 , new_n3330 , new_n3366 );
  nand     g05009 ( new_n5386 , new_n5384 , new_n5385 );
  xor      g05010 ( new_n5387 , new_n5380 , new_n5382 );
  nor      g05011 ( new_n5388 , new_n5386 , new_n5387 );
  nor      g05012 ( new_n5389 , new_n5383 , new_n5388 );
  xnor     g05013 ( new_n5390 , new_n5377 , new_n5378 );
  nor      g05014 ( new_n5391 , new_n5389 , new_n5390 );
  nor      g05015 ( new_n5392 , new_n5379 , new_n5391 );
  xor      g05016 ( new_n5393 , new_n5376 , new_n5392 );
  nand     g05017 ( new_n5394 , pi131 , pi196 );
  nor      g05018 ( new_n5395 , new_n3298 , new_n3309 );
  nand g05019 ( new_n5396 , new_n5395 , new_n5395 );
  nand     g05020 ( new_n5397 , pi131 , pi221 );
  nand     g05021 ( new_n5398 , new_n3304 , new_n3307 );
  nand     g05022 ( new_n5399 , new_n3303 , new_n3308 );
  nand     g05023 ( new_n5400 , new_n5398 , new_n5399 );
  xor      g05024 ( new_n5401 , new_n5397 , new_n5400 );
  nand     g05025 ( new_n5402 , pi029 , pi189 );
  nand     g05026 ( new_n5403 , pi077 , pi244 );
  nand     g05027 ( new_n5404 , pi069 , pi133 );
  xor      g05028 ( new_n5405 , new_n5403 , new_n5404 );
  xor      g05029 ( new_n5406 , new_n5402 , new_n5405 );
  nand     g05030 ( new_n5407 , pi052 , pi150 );
  nand     g05031 ( new_n5408 , new_n3300 , new_n3301 );
  nand     g05032 ( new_n5409 , new_n3299 , new_n3302 );
  nand     g05033 ( new_n5410 , new_n5408 , new_n5409 );
  xor      g05034 ( new_n5411 , new_n5407 , new_n5410 );
  xor      g05035 ( new_n5412 , new_n5406 , new_n5411 );
  xor      g05036 ( new_n5413 , new_n5401 , new_n5412 );
  nor      g05037 ( new_n5414 , new_n5396 , new_n5413 );
  nand g05038 ( new_n5415 , new_n5414 , new_n5414 );
  nand     g05039 ( new_n5416 , new_n5394 , new_n5415 );
  xor      g05040 ( new_n5417 , new_n5394 , new_n5415 );
  nand     g05041 ( new_n5418 , new_n5407 , new_n5410 );
  nand     g05042 ( new_n5419 , new_n5406 , new_n5411 );
  nand     g05043 ( new_n5420 , new_n5418 , new_n5419 );
  nand     g05044 ( new_n5421 , pi077 , pi150 );
  nand     g05045 ( new_n5422 , pi052 , pi221 );
  and      g05046 ( new_n5423 , new_n5421 , new_n5422 );
  nand     g05047 ( new_n5424 , pi077 , pi221 );
  nor      g05048 ( new_n5425 , new_n5407 , new_n5424 );
  or       g05049 ( new_n5426 , new_n5423 , new_n5425 );
  nand     g05050 ( new_n5427 , new_n5403 , new_n5404 );
  nand     g05051 ( new_n5428 , new_n5402 , new_n5405 );
  nand     g05052 ( new_n5429 , new_n5427 , new_n5428 );
  nand     g05053 ( new_n5430 , pi133 , pi244 );
  nand     g05054 ( new_n5431 , pi069 , pi189 );
  nand     g05055 ( new_n5432 , pi029 , pi064 );
  nand     g05056 ( new_n5433 , new_n5431 , new_n5432 );
  nand     g05057 ( new_n5434 , pi064 , pi069 );
  or       g05058 ( new_n5435 , new_n5402 , new_n5434 );
  nand     g05059 ( new_n5436 , new_n5433 , new_n5435 );
  xor      g05060 ( new_n5437 , new_n5430 , new_n5436 );
  xor      g05061 ( new_n5438 , new_n5429 , new_n5437 );
  xor      g05062 ( new_n5439 , new_n5426 , new_n5438 );
  nand g05063 ( new_n5440 , new_n5439 , new_n5439 );
  xor      g05064 ( new_n5441 , new_n5420 , new_n5440 );
  nor      g05065 ( new_n5442 , new_n5397 , new_n5400 );
  nand g05066 ( new_n5443 , new_n5412 , new_n5412 );
  nand     g05067 ( new_n5444 , new_n5401 , new_n5443 );
  nand g05068 ( new_n5445 , new_n5444 , new_n5444 );
  nor      g05069 ( new_n5446 , new_n5442 , new_n5445 );
  xor      g05070 ( new_n5447 , new_n5441 , new_n5446 );
  nand     g05071 ( new_n5448 , new_n5417 , new_n5447 );
  nand     g05072 ( new_n5449 , new_n5416 , new_n5448 );
  nand g05073 ( new_n5450 , new_n5441 , new_n5441 );
  nor      g05074 ( new_n5451 , new_n5450 , new_n5446 );
  nor      g05075 ( new_n5452 , new_n5426 , new_n5438 );
  nor      g05076 ( new_n5453 , new_n5420 , new_n5440 );
  xor      g05077 ( new_n5454 , new_n5425 , new_n5453 );
  nor      g05078 ( new_n5455 , new_n5452 , new_n5454 );
  nand     g05079 ( new_n5456 , pi133 , pi150 );
  xor      g05080 ( new_n5457 , new_n5435 , new_n5456 );
  nand     g05081 ( new_n5458 , pi029 , pi084 );
  and      g05082 ( new_n5459 , pi189 , pi244 );
  xor      g05083 ( new_n5460 , new_n5458 , new_n5459 );
  xor      g05084 ( new_n5461 , new_n5434 , new_n5460 );
  xor      g05085 ( new_n5462 , new_n5457 , new_n5461 );
  nand     g05086 ( new_n5463 , new_n5430 , new_n5436 );
  nand     g05087 ( new_n5464 , new_n5429 , new_n5437 );
  nand     g05088 ( new_n5465 , new_n5463 , new_n5464 );
  nand     g05089 ( new_n5466 , pi052 , pi196 );
  nand     g05090 ( new_n5467 , pi131 , pi184 );
  xor      g05091 ( new_n5468 , new_n5466 , new_n5467 );
  xnor     g05092 ( new_n5469 , new_n5424 , new_n5468 );
  xor      g05093 ( new_n5470 , new_n5465 , new_n5469 );
  xor      g05094 ( new_n5471 , new_n5462 , new_n5470 );
  xnor     g05095 ( new_n5472 , new_n5455 , new_n5471 );
  xor      g05096 ( new_n5473 , new_n5451 , new_n5472 );
  xor      g05097 ( new_n5474 , new_n5449 , new_n5473 );
  xnor     g05098 ( new_n5475 , new_n5393 , new_n5474 );
  xor      g05099 ( new_n5476 , new_n5389 , new_n5390 );
  xor      g05100 ( new_n5477 , new_n5396 , new_n5413 );
  nor      g05101 ( new_n5478 , new_n3296 , new_n3310 );
  and      g05102 ( new_n5479 , new_n3311 , new_n3367 );
  or       g05103 ( new_n5480 , new_n5478 , new_n5479 );
  nor      g05104 ( new_n5481 , new_n5477 , new_n5480 );
  xor      g05105 ( new_n5482 , new_n5386 , new_n5387 );
  xnor     g05106 ( new_n5483 , new_n5477 , new_n5480 );
  nor      g05107 ( new_n5484 , new_n5482 , new_n5483 );
  nor      g05108 ( new_n5485 , new_n5481 , new_n5484 );
  nand     g05109 ( new_n5486 , new_n5476 , new_n5485 );
  xor      g05110 ( new_n5487 , new_n5476 , new_n5485 );
  xor      g05111 ( new_n5488 , new_n5417 , new_n5447 );
  nand g05112 ( new_n5489 , new_n5488 , new_n5488 );
  nand     g05113 ( new_n5490 , new_n5487 , new_n5489 );
  nand     g05114 ( new_n5491 , new_n5486 , new_n5490 );
  xnor     g05115 ( po019 , new_n5475 , new_n5491 );
  xnor     g05116 ( po020 , new_n3263 , new_n3294 );
  nand     g05117 ( new_n5494 , pi079 , pi179 );
  nand     g05118 ( new_n5495 , pi142 , pi144 );
  nor      g05119 ( new_n5496 , new_n5050 , new_n5051 );
  nor      g05120 ( new_n5497 , new_n5048 , new_n5052 );
  nor      g05121 ( new_n5498 , new_n5496 , new_n5497 );
  or       g05122 ( new_n5499 , new_n5495 , new_n5498 );
  xor      g05123 ( new_n5500 , new_n5495 , new_n5498 );
  nand     g05124 ( new_n5501 , pi123 , pi178 );
  nand     g05125 ( new_n5502 , pi099 , pi188 );
  nand     g05126 ( new_n5503 , pi061 , pi169 );
  xor      g05127 ( new_n5504 , new_n5502 , new_n5503 );
  xor      g05128 ( new_n5505 , new_n5501 , new_n5504 );
  nand     g05129 ( new_n5506 , pi012 , pi071 );
  nand     g05130 ( new_n5507 , new_n5045 , new_n5046 );
  nand     g05131 ( new_n5508 , new_n5044 , new_n5047 );
  nand     g05132 ( new_n5509 , new_n5507 , new_n5508 );
  xor      g05133 ( new_n5510 , new_n5506 , new_n5509 );
  xnor     g05134 ( new_n5511 , new_n5505 , new_n5510 );
  nand     g05135 ( new_n5512 , new_n5500 , new_n5511 );
  nand     g05136 ( new_n5513 , new_n5499 , new_n5512 );
  nand g05137 ( new_n5514 , new_n5513 , new_n5513 );
  nand     g05138 ( new_n5515 , pi061 , pi123 );
  nand     g05139 ( new_n5516 , pi099 , pi178 );
  nand     g05140 ( new_n5517 , pi023 , pi188 );
  nand     g05141 ( new_n5518 , new_n5516 , new_n5517 );
  nand     g05142 ( new_n5519 , pi023 , pi178 );
  or       g05143 ( new_n5520 , new_n5502 , new_n5519 );
  nand     g05144 ( new_n5521 , new_n5518 , new_n5520 );
  xor      g05145 ( new_n5522 , new_n5515 , new_n5521 );
  nand     g05146 ( new_n5523 , new_n5502 , new_n5503 );
  nand     g05147 ( new_n5524 , new_n5501 , new_n5504 );
  nand     g05148 ( new_n5525 , new_n5523 , new_n5524 );
  xor      g05149 ( new_n5526 , new_n5522 , new_n5525 );
  nand     g05150 ( new_n5527 , pi144 , pi169 );
  nor      g05151 ( new_n5528 , new_n5506 , new_n5527 );
  nand     g05152 ( new_n5529 , pi012 , pi169 );
  nand     g05153 ( new_n5530 , pi071 , pi144 );
  and      g05154 ( new_n5531 , new_n5529 , new_n5530 );
  or       g05155 ( new_n5532 , new_n5528 , new_n5531 );
  xor      g05156 ( new_n5533 , new_n5526 , new_n5532 );
  nand     g05157 ( new_n5534 , new_n5506 , new_n5509 );
  nand     g05158 ( new_n5535 , new_n5505 , new_n5510 );
  nand     g05159 ( new_n5536 , new_n5534 , new_n5535 );
  xor      g05160 ( new_n5537 , new_n5533 , new_n5536 );
  or       g05161 ( new_n5538 , new_n5514 , new_n5537 );
  nor      g05162 ( new_n5539 , new_n5526 , new_n5532 );
  nand g05163 ( new_n5540 , new_n5533 , new_n5533 );
  nor      g05164 ( new_n5541 , new_n5540 , new_n5536 );
  xor      g05165 ( new_n5542 , new_n5528 , new_n5541 );
  nor      g05166 ( new_n5543 , new_n5539 , new_n5542 );
  nand     g05167 ( new_n5544 , pi071 , pi098 );
  nand     g05168 ( new_n5545 , pi043 , pi142 );
  xor      g05169 ( new_n5546 , new_n5544 , new_n5545 );
  xor      g05170 ( new_n5547 , new_n5527 , new_n5546 );
  nand     g05171 ( new_n5548 , new_n5515 , new_n5521 );
  nand     g05172 ( new_n5549 , new_n5522 , new_n5525 );
  nand     g05173 ( new_n5550 , new_n5548 , new_n5549 );
  xor      g05174 ( new_n5551 , new_n5547 , new_n5550 );
  nand     g05175 ( new_n5552 , pi012 , pi123 );
  xnor     g05176 ( new_n5553 , new_n5520 , new_n5552 );
  nand     g05177 ( new_n5554 , pi061 , pi099 );
  nand     g05178 ( new_n5555 , pi155 , pi188 );
  xor      g05179 ( new_n5556 , new_n5554 , new_n5555 );
  xor      g05180 ( new_n5557 , new_n5519 , new_n5556 );
  xnor     g05181 ( new_n5558 , new_n5553 , new_n5557 );
  xnor     g05182 ( new_n5559 , new_n5551 , new_n5558 );
  xor      g05183 ( new_n5560 , new_n5543 , new_n5559 );
  xor      g05184 ( new_n5561 , new_n5538 , new_n5560 );
  nand     g05185 ( new_n5562 , pi098 , pi142 );
  or       g05186 ( new_n5563 , new_n5043 , new_n5053 );
  xnor     g05187 ( new_n5564 , new_n5500 , new_n5511 );
  or       g05188 ( new_n5565 , new_n5563 , new_n5564 );
  nand     g05189 ( new_n5566 , new_n5562 , new_n5565 );
  xor      g05190 ( new_n5567 , new_n5513 , new_n5537 );
  nand g05191 ( new_n5568 , new_n5567 , new_n5567 );
  xnor     g05192 ( new_n5569 , new_n5562 , new_n5565 );
  or       g05193 ( new_n5570 , new_n5568 , new_n5569 );
  nand     g05194 ( new_n5571 , new_n5566 , new_n5570 );
  xor      g05195 ( new_n5572 , new_n5561 , new_n5571 );
  nand g05196 ( new_n5573 , new_n5572 , new_n5572 );
  nand     g05197 ( new_n5574 , pi118 , pi219 );
  nand     g05198 ( new_n5575 , pi007 , pi102 );
  and      g05199 ( new_n5576 , new_n5574 , new_n5575 );
  nand     g05200 ( new_n5577 , pi007 , pi219 );
  nand     g05201 ( new_n5578 , pi102 , pi118 );
  nor      g05202 ( new_n5579 , new_n5577 , new_n5578 );
  or       g05203 ( new_n5580 , new_n5576 , new_n5579 );
  nand     g05204 ( new_n5581 , pi102 , pi108 );
  nand     g05205 ( new_n5582 , pi001 , pi042 );
  nand     g05206 ( new_n5583 , new_n5581 , new_n5582 );
  nand     g05207 ( new_n5584 , pi051 , pi122 );
  xor      g05208 ( new_n5585 , new_n5581 , new_n5582 );
  nand     g05209 ( new_n5586 , new_n5584 , new_n5585 );
  nand     g05210 ( new_n5587 , new_n5583 , new_n5586 );
  nand     g05211 ( new_n5588 , pi001 , pi108 );
  nand     g05212 ( new_n5589 , pi042 , pi122 );
  nand     g05213 ( new_n5590 , pi051 , pi135 );
  nand     g05214 ( new_n5591 , new_n5589 , new_n5590 );
  nand     g05215 ( new_n5592 , pi042 , pi135 );
  or       g05216 ( new_n5593 , new_n5584 , new_n5592 );
  nand     g05217 ( new_n5594 , new_n5591 , new_n5593 );
  xor      g05218 ( new_n5595 , new_n5588 , new_n5594 );
  xor      g05219 ( new_n5596 , new_n5587 , new_n5595 );
  nor      g05220 ( new_n5597 , new_n5580 , new_n5596 );
  nand     g05221 ( new_n5598 , new_n5057 , new_n5058 );
  nand     g05222 ( new_n5599 , new_n5056 , new_n5059 );
  nand     g05223 ( new_n5600 , new_n5598 , new_n5599 );
  nand     g05224 ( new_n5601 , new_n5577 , new_n5600 );
  xor      g05225 ( new_n5602 , new_n5584 , new_n5585 );
  xor      g05226 ( new_n5603 , new_n5577 , new_n5600 );
  nand     g05227 ( new_n5604 , new_n5602 , new_n5603 );
  nand     g05228 ( new_n5605 , new_n5601 , new_n5604 );
  xnor     g05229 ( new_n5606 , new_n5580 , new_n5596 );
  nor      g05230 ( new_n5607 , new_n5605 , new_n5606 );
  xor      g05231 ( new_n5608 , new_n5579 , new_n5607 );
  nor      g05232 ( new_n5609 , new_n5597 , new_n5608 );
  nand     g05233 ( new_n5610 , new_n5588 , new_n5594 );
  nand     g05234 ( new_n5611 , new_n5587 , new_n5595 );
  nand     g05235 ( new_n5612 , new_n5610 , new_n5611 );
  nand     g05236 ( new_n5613 , pi038 , pi087 );
  nand     g05237 ( new_n5614 , pi113 , pi219 );
  xor      g05238 ( new_n5615 , new_n5613 , new_n5614 );
  xor      g05239 ( new_n5616 , new_n5578 , new_n5615 );
  xor      g05240 ( new_n5617 , new_n5612 , new_n5616 );
  nand     g05241 ( new_n5618 , pi001 , pi007 );
  xnor     g05242 ( new_n5619 , new_n5593 , new_n5618 );
  nand     g05243 ( new_n5620 , pi051 , pi059 );
  nand     g05244 ( new_n5621 , pi108 , pi122 );
  xor      g05245 ( new_n5622 , new_n5620 , new_n5621 );
  xor      g05246 ( new_n5623 , new_n5592 , new_n5622 );
  xor      g05247 ( new_n5624 , new_n5619 , new_n5623 );
  xor      g05248 ( new_n5625 , new_n5617 , new_n5624 );
  nand g05249 ( new_n5626 , new_n5625 , new_n5625 );
  xor      g05250 ( new_n5627 , new_n5609 , new_n5626 );
  xor      g05251 ( new_n5628 , new_n5605 , new_n5606 );
  nand     g05252 ( new_n5629 , pi087 , pi118 );
  nand g05253 ( new_n5630 , new_n5629 , new_n5629 );
  nor      g05254 ( new_n5631 , new_n5061 , new_n5063 );
  nor      g05255 ( new_n5632 , new_n5060 , new_n5064 );
  or       g05256 ( new_n5633 , new_n5631 , new_n5632 );
  nor      g05257 ( new_n5634 , new_n5630 , new_n5633 );
  and      g05258 ( new_n5635 , new_n5630 , new_n5633 );
  xnor     g05259 ( new_n5636 , new_n5602 , new_n5603 );
  nor      g05260 ( new_n5637 , new_n5635 , new_n5636 );
  nor      g05261 ( new_n5638 , new_n5634 , new_n5637 );
  and      g05262 ( new_n5639 , new_n5628 , new_n5638 );
  xor      g05263 ( new_n5640 , new_n5627 , new_n5639 );
  nand g05264 ( new_n5641 , new_n5640 , new_n5640 );
  nand     g05265 ( new_n5642 , pi087 , pi113 );
  xnor     g05266 ( new_n5643 , new_n5628 , new_n5638 );
  nor      g05267 ( new_n5644 , new_n5642 , new_n5643 );
  nand g05268 ( new_n5645 , new_n5055 , new_n5055 );
  nor      g05269 ( new_n5646 , new_n5645 , new_n5065 );
  nand g05270 ( new_n5647 , new_n5646 , new_n5646 );
  or       g05271 ( new_n5648 , new_n5634 , new_n5635 );
  xor      g05272 ( new_n5649 , new_n5636 , new_n5648 );
  or       g05273 ( new_n5650 , new_n5647 , new_n5649 );
  xnor     g05274 ( new_n5651 , new_n5642 , new_n5643 );
  nor      g05275 ( new_n5652 , new_n5650 , new_n5651 );
  nor      g05276 ( new_n5653 , new_n5644 , new_n5652 );
  xor      g05277 ( new_n5654 , new_n5641 , new_n5653 );
  xor      g05278 ( new_n5655 , new_n5573 , new_n5654 );
  xnor     g05279 ( new_n5656 , new_n5650 , new_n5651 );
  xor      g05280 ( new_n5657 , new_n5567 , new_n5569 );
  nand g05281 ( new_n5658 , new_n5657 , new_n5657 );
  nor      g05282 ( new_n5659 , new_n5656 , new_n5658 );
  xor      g05283 ( new_n5660 , new_n5646 , new_n5649 );
  xnor     g05284 ( new_n5661 , new_n5563 , new_n5564 );
  nand     g05285 ( new_n5662 , new_n5660 , new_n5661 );
  xor      g05286 ( new_n5663 , new_n5660 , new_n5661 );
  nor      g05287 ( new_n5664 , new_n5054 , new_n5066 );
  nor      g05288 ( new_n5665 , new_n5067 , new_n5070 );
  nor      g05289 ( new_n5666 , new_n5664 , new_n5665 );
  nand     g05290 ( new_n5667 , new_n5663 , new_n5666 );
  nand     g05291 ( new_n5668 , new_n5662 , new_n5667 );
  xor      g05292 ( new_n5669 , new_n5656 , new_n5657 );
  nor      g05293 ( new_n5670 , new_n5668 , new_n5669 );
  nor      g05294 ( new_n5671 , new_n5659 , new_n5670 );
  xor      g05295 ( new_n5672 , new_n5655 , new_n5671 );
  nand     g05296 ( new_n5673 , pi138 , pi237 );
  nand     g05297 ( new_n5674 , pi048 , pi182 );
  nand     g05298 ( new_n5675 , new_n5031 , new_n5032 );
  nand     g05299 ( new_n5676 , new_n5030 , new_n5033 );
  nand     g05300 ( new_n5677 , new_n5675 , new_n5676 );
  xor      g05301 ( new_n5678 , new_n5674 , new_n5677 );
  nand     g05302 ( new_n5679 , pi076 , pi162 );
  nand     g05303 ( new_n5680 , pi033 , pi216 );
  nand     g05304 ( new_n5681 , pi041 , pi179 );
  xor      g05305 ( new_n5682 , new_n5680 , new_n5681 );
  xor      g05306 ( new_n5683 , new_n5679 , new_n5682 );
  xnor     g05307 ( new_n5684 , new_n5678 , new_n5683 );
  nand g05308 ( new_n5685 , new_n5684 , new_n5684 );
  nor      g05309 ( new_n5686 , new_n5673 , new_n5685 );
  nand     g05310 ( new_n5687 , new_n5035 , new_n5038 );
  nand     g05311 ( new_n5688 , new_n5034 , new_n5039 );
  nand     g05312 ( new_n5689 , new_n5687 , new_n5688 );
  xor      g05313 ( new_n5690 , new_n5673 , new_n5684 );
  nor      g05314 ( new_n5691 , new_n5689 , new_n5690 );
  nor      g05315 ( new_n5692 , new_n5686 , new_n5691 );
  nand     g05316 ( new_n5693 , pi041 , pi048 );
  nand     g05317 ( new_n5694 , pi182 , pi237 );
  nand     g05318 ( new_n5695 , new_n5693 , new_n5694 );
  nand     g05319 ( new_n5696 , pi041 , pi237 );
  or       g05320 ( new_n5697 , new_n5674 , new_n5696 );
  nand     g05321 ( new_n5698 , new_n5695 , new_n5697 );
  nand     g05322 ( new_n5699 , new_n5680 , new_n5681 );
  nand     g05323 ( new_n5700 , new_n5679 , new_n5682 );
  nand     g05324 ( new_n5701 , new_n5699 , new_n5700 );
  nand     g05325 ( new_n5702 , pi179 , pi216 );
  nand     g05326 ( new_n5703 , pi033 , pi076 );
  nand     g05327 ( new_n5704 , pi079 , pi162 );
  nand     g05328 ( new_n5705 , new_n5703 , new_n5704 );
  nand     g05329 ( new_n5706 , pi033 , pi079 );
  nor      g05330 ( new_n5707 , new_n5679 , new_n5706 );
  nand g05331 ( new_n5708 , new_n5707 , new_n5707 );
  nand     g05332 ( new_n5709 , new_n5705 , new_n5708 );
  xor      g05333 ( new_n5710 , new_n5702 , new_n5709 );
  xor      g05334 ( new_n5711 , new_n5701 , new_n5710 );
  xor      g05335 ( new_n5712 , new_n5698 , new_n5711 );
  nand     g05336 ( new_n5713 , new_n5674 , new_n5677 );
  nand     g05337 ( new_n5714 , new_n5678 , new_n5683 );
  nand     g05338 ( new_n5715 , new_n5713 , new_n5714 );
  xor      g05339 ( new_n5716 , new_n5712 , new_n5715 );
  or       g05340 ( new_n5717 , new_n5692 , new_n5716 );
  nand     g05341 ( new_n5718 , new_n5698 , new_n5711 );
  nand     g05342 ( new_n5719 , new_n5712 , new_n5715 );
  nand     g05343 ( new_n5720 , new_n5718 , new_n5719 );
  xnor     g05344 ( new_n5721 , new_n5697 , new_n5720 );
  nand     g05345 ( new_n5722 , pi048 , pi216 );
  xor      g05346 ( new_n5723 , new_n5707 , new_n5722 );
  nand     g05347 ( new_n5724 , pi162 , pi251 );
  nand     g05348 ( new_n5725 , pi076 , pi179 );
  xor      g05349 ( new_n5726 , new_n5724 , new_n5725 );
  xor      g05350 ( new_n5727 , new_n5706 , new_n5726 );
  xor      g05351 ( new_n5728 , new_n5723 , new_n5727 );
  nand     g05352 ( new_n5729 , new_n5702 , new_n5709 );
  nand     g05353 ( new_n5730 , new_n5701 , new_n5710 );
  nand     g05354 ( new_n5731 , new_n5729 , new_n5730 );
  nand     g05355 ( new_n5732 , pi182 , pi238 );
  nand     g05356 ( new_n5733 , pi138 , pi193 );
  xor      g05357 ( new_n5734 , new_n5732 , new_n5733 );
  xor      g05358 ( new_n5735 , new_n5696 , new_n5734 );
  xor      g05359 ( new_n5736 , new_n5731 , new_n5735 );
  nand g05360 ( new_n5737 , new_n5736 , new_n5736 );
  xor      g05361 ( new_n5738 , new_n5728 , new_n5737 );
  xor      g05362 ( new_n5739 , new_n5721 , new_n5738 );
  nand g05363 ( new_n5740 , new_n5739 , new_n5739 );
  xor      g05364 ( new_n5741 , new_n5717 , new_n5740 );
  nand     g05365 ( new_n5742 , pi138 , pi238 );
  nor      g05366 ( new_n5743 , new_n5029 , new_n5040 );
  xor      g05367 ( new_n5744 , new_n5689 , new_n5690 );
  nand     g05368 ( new_n5745 , new_n5743 , new_n5744 );
  nand     g05369 ( new_n5746 , new_n5742 , new_n5745 );
  xor      g05370 ( new_n5747 , new_n5742 , new_n5745 );
  xor      g05371 ( new_n5748 , new_n5692 , new_n5716 );
  nand g05372 ( new_n5749 , new_n5748 , new_n5748 );
  nand     g05373 ( new_n5750 , new_n5747 , new_n5749 );
  nand     g05374 ( new_n5751 , new_n5746 , new_n5750 );
  xor      g05375 ( new_n5752 , new_n5741 , new_n5751 );
  nor      g05376 ( new_n5753 , new_n5672 , new_n5752 );
  xnor     g05377 ( new_n5754 , new_n5743 , new_n5744 );
  nand g05378 ( new_n5755 , new_n5028 , new_n5028 );
  and      g05379 ( new_n5756 , new_n5755 , new_n5041 );
  nor      g05380 ( new_n5757 , new_n5042 , new_n5071 );
  or       g05381 ( new_n5758 , new_n5756 , new_n5757 );
  nor      g05382 ( new_n5759 , new_n5754 , new_n5758 );
  xnor     g05383 ( new_n5760 , new_n5754 , new_n5758 );
  xor      g05384 ( new_n5761 , new_n5663 , new_n5666 );
  nor      g05385 ( new_n5762 , new_n5760 , new_n5761 );
  nor      g05386 ( new_n5763 , new_n5759 , new_n5762 );
  xnor     g05387 ( new_n5764 , new_n5668 , new_n5669 );
  nand     g05388 ( new_n5765 , new_n5763 , new_n5764 );
  xor      g05389 ( new_n5766 , new_n5747 , new_n5748 );
  xor      g05390 ( new_n5767 , new_n5763 , new_n5764 );
  nand g05391 ( new_n5768 , new_n5767 , new_n5767 );
  or       g05392 ( new_n5769 , new_n5766 , new_n5768 );
  nand     g05393 ( new_n5770 , new_n5765 , new_n5769 );
  xnor     g05394 ( new_n5771 , new_n5672 , new_n5752 );
  nor      g05395 ( new_n5772 , new_n5770 , new_n5771 );
  or       g05396 ( new_n5773 , new_n5753 , new_n5772 );
  xor      g05397 ( new_n5774 , new_n5494 , new_n5773 );
  nand     g05398 ( new_n5775 , pi155 , pi178 );
  xor      g05399 ( new_n5776 , new_n5774 , new_n5775 );
  nand     g05400 ( new_n5777 , pi194 , pi223 );
  nand     g05401 ( new_n5778 , pi143 , pi225 );
  nand     g05402 ( new_n5779 , pi057 , pi101 );
  nand     g05403 ( new_n5780 , new_n5778 , new_n5779 );
  nand     g05404 ( new_n5781 , pi101 , pi143 );
  nand     g05405 ( new_n5782 , pi057 , pi225 );
  nor      g05406 ( new_n5783 , new_n5781 , new_n5782 );
  nand g05407 ( new_n5784 , new_n5783 , new_n5783 );
  nand     g05408 ( new_n5785 , new_n5780 , new_n5784 );
  nand     g05409 ( new_n5786 , new_n5777 , new_n5785 );
  nand     g05410 ( new_n5787 , pi057 , pi223 );
  nand     g05411 ( new_n5788 , new_n5781 , new_n5787 );
  nand     g05412 ( new_n5789 , pi060 , pi194 );
  xor      g05413 ( new_n5790 , new_n5781 , new_n5787 );
  nand     g05414 ( new_n5791 , new_n5789 , new_n5790 );
  nand     g05415 ( new_n5792 , new_n5788 , new_n5791 );
  xor      g05416 ( new_n5793 , new_n5777 , new_n5785 );
  nand     g05417 ( new_n5794 , new_n5792 , new_n5793 );
  nand     g05418 ( new_n5795 , new_n5786 , new_n5794 );
  nand     g05419 ( new_n5796 , pi060 , pi180 );
  nand     g05420 ( new_n5797 , pi068 , pi160 );
  nand     g05421 ( new_n5798 , pi020 , pi036 );
  xor      g05422 ( new_n5799 , new_n5797 , new_n5798 );
  xor      g05423 ( new_n5800 , new_n5796 , new_n5799 );
  or       g05424 ( new_n5801 , new_n5795 , new_n5800 );
  nand     g05425 ( new_n5802 , pi143 , pi177 );
  nand     g05426 ( new_n5803 , pi101 , pi194 );
  xor      g05427 ( new_n5804 , new_n5802 , new_n5803 );
  xor      g05428 ( new_n5805 , new_n5782 , new_n5804 );
  nand     g05429 ( new_n5806 , pi085 , pi223 );
  xor      g05430 ( new_n5807 , new_n5783 , new_n5806 );
  xor      g05431 ( new_n5808 , new_n5805 , new_n5807 );
  xor      g05432 ( new_n5809 , new_n5795 , new_n5800 );
  nand     g05433 ( new_n5810 , new_n5808 , new_n5809 );
  nand     g05434 ( new_n5811 , new_n5801 , new_n5810 );
  nand     g05435 ( new_n5812 , new_n5528 , new_n5541 );
  nand g05436 ( new_n5813 , new_n5543 , new_n5543 );
  nand     g05437 ( new_n5814 , new_n5813 , new_n5559 );
  nand     g05438 ( new_n5815 , new_n5812 , new_n5814 );
  nor      g05439 ( new_n5816 , new_n5708 , new_n5722 );
  nor      g05440 ( new_n5817 , new_n5723 , new_n5727 );
  nor      g05441 ( new_n5818 , new_n5816 , new_n5817 );
  xor      g05442 ( new_n5819 , new_n5815 , new_n5818 );
  xor      g05443 ( new_n5820 , new_n5811 , new_n5819 );
  xor      g05444 ( new_n5821 , new_n5776 , new_n5820 );
  nand     g05445 ( new_n5822 , pi194 , pi225 );
  nand     g05446 ( new_n5823 , pi033 , pi251 );
  xor      g05447 ( new_n5824 , new_n5822 , new_n5823 );
  nand     g05448 ( new_n5825 , pi138 , pi159 );
  nand     g05449 ( new_n5826 , pi085 , pi101 );
  nand     g05450 ( new_n5827 , pi020 , pi068 );
  xor      g05451 ( new_n5828 , new_n5826 , new_n5827 );
  xor      g05452 ( new_n5829 , new_n5825 , new_n5828 );
  nand     g05453 ( new_n5830 , pi036 , pi060 );
  nand     g05454 ( new_n5831 , new_n5802 , new_n5803 );
  nand     g05455 ( new_n5832 , new_n5782 , new_n5804 );
  nand     g05456 ( new_n5833 , new_n5831 , new_n5832 );
  xor      g05457 ( new_n5834 , new_n5830 , new_n5833 );
  xor      g05458 ( new_n5835 , new_n5829 , new_n5834 );
  xor      g05459 ( new_n5836 , new_n5824 , new_n5835 );
  xor      g05460 ( new_n5837 , new_n5821 , new_n5836 );
  nand     g05461 ( new_n5838 , pi180 , pi223 );
  nor      g05462 ( new_n5839 , new_n5717 , new_n5740 );
  nand g05463 ( new_n5840 , new_n5741 , new_n5741 );
  nor      g05464 ( new_n5841 , new_n5840 , new_n5751 );
  nor      g05465 ( new_n5842 , new_n5839 , new_n5841 );
  xor      g05466 ( new_n5843 , new_n5838 , new_n5842 );
  nand     g05467 ( new_n5844 , new_n5797 , new_n5798 );
  nand     g05468 ( new_n5845 , new_n5796 , new_n5799 );
  nand     g05469 ( new_n5846 , new_n5844 , new_n5845 );
  nor      g05470 ( new_n5847 , new_n5697 , new_n5720 );
  nor      g05471 ( new_n5848 , new_n5721 , new_n5738 );
  nor      g05472 ( new_n5849 , new_n5847 , new_n5848 );
  xor      g05473 ( new_n5850 , new_n5846 , new_n5849 );
  xor      g05474 ( new_n5851 , new_n5843 , new_n5850 );
  nand     g05475 ( new_n5852 , new_n5547 , new_n5550 );
  nand     g05476 ( new_n5853 , new_n5551 , new_n5558 );
  nand     g05477 ( new_n5854 , new_n5852 , new_n5853 );
  nand     g05478 ( new_n5855 , pi012 , pi099 );
  nand     g05479 ( new_n5856 , pi098 , pi169 );
  xor      g05480 ( new_n5857 , new_n5855 , new_n5856 );
  xor      g05481 ( new_n5858 , new_n5854 , new_n5857 );
  and      g05482 ( new_n5859 , new_n5579 , new_n5607 );
  nor      g05483 ( new_n5860 , new_n5609 , new_n5626 );
  nor      g05484 ( new_n5861 , new_n5859 , new_n5860 );
  nand     g05485 ( new_n5862 , new_n5544 , new_n5545 );
  nand     g05486 ( new_n5863 , new_n5527 , new_n5546 );
  nand     g05487 ( new_n5864 , new_n5862 , new_n5863 );
  nand     g05488 ( new_n5865 , pi051 , pi094 );
  nor      g05489 ( new_n5866 , new_n5520 , new_n5552 );
  nor      g05490 ( new_n5867 , new_n5553 , new_n5557 );
  nor      g05491 ( new_n5868 , new_n5866 , new_n5867 );
  xor      g05492 ( new_n5869 , new_n5865 , new_n5868 );
  xor      g05493 ( new_n5870 , new_n5864 , new_n5869 );
  xor      g05494 ( new_n5871 , new_n5861 , new_n5870 );
  xor      g05495 ( new_n5872 , new_n5858 , new_n5871 );
  nand     g05496 ( new_n5873 , pi036 , pi160 );
  nor      g05497 ( new_n5874 , new_n5011 , new_n5022 );
  nand     g05498 ( new_n5875 , new_n5017 , new_n5020 );
  nand     g05499 ( new_n5876 , new_n5016 , new_n5021 );
  nand     g05500 ( new_n5877 , new_n5875 , new_n5876 );
  nand     g05501 ( new_n5878 , pi160 , pi180 );
  xor      g05502 ( new_n5879 , new_n5789 , new_n5790 );
  nand     g05503 ( new_n5880 , pi020 , pi085 );
  nand     g05504 ( new_n5881 , new_n5013 , new_n5014 );
  nand     g05505 ( new_n5882 , new_n5012 , new_n5015 );
  nand     g05506 ( new_n5883 , new_n5881 , new_n5882 );
  xor      g05507 ( new_n5884 , new_n5880 , new_n5883 );
  xor      g05508 ( new_n5885 , new_n5879 , new_n5884 );
  xnor     g05509 ( new_n5886 , new_n5878 , new_n5885 );
  xor      g05510 ( new_n5887 , new_n5877 , new_n5886 );
  nand     g05511 ( new_n5888 , new_n5874 , new_n5887 );
  xor      g05512 ( new_n5889 , new_n5873 , new_n5888 );
  nor      g05513 ( new_n5890 , new_n5878 , new_n5885 );
  nor      g05514 ( new_n5891 , new_n5877 , new_n5886 );
  nor      g05515 ( new_n5892 , new_n5890 , new_n5891 );
  nand     g05516 ( new_n5893 , new_n5880 , new_n5883 );
  nand     g05517 ( new_n5894 , new_n5879 , new_n5884 );
  nand     g05518 ( new_n5895 , new_n5893 , new_n5894 );
  nor      g05519 ( new_n5896 , new_n5796 , new_n5880 );
  nand g05520 ( new_n5897 , new_n5896 , new_n5896 );
  nand     g05521 ( new_n5898 , pi020 , pi180 );
  nand     g05522 ( new_n5899 , pi060 , pi085 );
  nand     g05523 ( new_n5900 , new_n5898 , new_n5899 );
  nand     g05524 ( new_n5901 , new_n5897 , new_n5900 );
  xor      g05525 ( new_n5902 , new_n5792 , new_n5793 );
  xnor     g05526 ( new_n5903 , new_n5901 , new_n5902 );
  xor      g05527 ( new_n5904 , new_n5895 , new_n5903 );
  xor      g05528 ( new_n5905 , new_n5892 , new_n5904 );
  xor      g05529 ( new_n5906 , new_n5889 , new_n5905 );
  nand g05530 ( new_n5907 , new_n5906 , new_n5906 );
  xor      g05531 ( new_n5908 , new_n5766 , new_n5767 );
  nor      g05532 ( new_n5909 , new_n5907 , new_n5908 );
  nor      g05533 ( new_n5910 , new_n5010 , new_n5024 );
  and      g05534 ( new_n5911 , new_n5025 , new_n5072 );
  nor      g05535 ( new_n5912 , new_n5910 , new_n5911 );
  xnor     g05536 ( new_n5913 , new_n5874 , new_n5887 );
  and      g05537 ( new_n5914 , new_n5912 , new_n5913 );
  xnor     g05538 ( new_n5915 , new_n5912 , new_n5913 );
  xor      g05539 ( new_n5916 , new_n5760 , new_n5761 );
  nor      g05540 ( new_n5917 , new_n5915 , new_n5916 );
  nor      g05541 ( new_n5918 , new_n5914 , new_n5917 );
  xor      g05542 ( new_n5919 , new_n5906 , new_n5908 );
  nor      g05543 ( new_n5920 , new_n5918 , new_n5919 );
  nor      g05544 ( new_n5921 , new_n5909 , new_n5920 );
  nand g05545 ( new_n5922 , new_n5904 , new_n5904 );
  nor      g05546 ( new_n5923 , new_n5892 , new_n5922 );
  nand     g05547 ( new_n5924 , new_n5873 , new_n5888 );
  nand     g05548 ( new_n5925 , new_n5889 , new_n5905 );
  nand     g05549 ( new_n5926 , new_n5924 , new_n5925 );
  xor      g05550 ( new_n5927 , new_n5808 , new_n5809 );
  nor      g05551 ( new_n5928 , new_n5901 , new_n5902 );
  nor      g05552 ( new_n5929 , new_n5895 , new_n5903 );
  xor      g05553 ( new_n5930 , new_n5897 , new_n5929 );
  nand g05554 ( new_n5931 , new_n5930 , new_n5930 );
  nor      g05555 ( new_n5932 , new_n5928 , new_n5931 );
  xor      g05556 ( new_n5933 , new_n5927 , new_n5932 );
  xor      g05557 ( new_n5934 , new_n5926 , new_n5933 );
  xor      g05558 ( new_n5935 , new_n5923 , new_n5934 );
  or       g05559 ( new_n5936 , new_n5921 , new_n5935 );
  xnor     g05560 ( new_n5937 , new_n5770 , new_n5771 );
  xor      g05561 ( new_n5938 , new_n5921 , new_n5935 );
  nand     g05562 ( new_n5939 , new_n5937 , new_n5938 );
  nand     g05563 ( new_n5940 , new_n5936 , new_n5939 );
  xor      g05564 ( new_n5941 , new_n5872 , new_n5940 );
  nand     g05565 ( new_n5942 , new_n5627 , new_n5639 );
  or       g05566 ( new_n5943 , new_n5641 , new_n5653 );
  nand     g05567 ( new_n5944 , new_n5942 , new_n5943 );
  nand     g05568 ( new_n5945 , new_n5732 , new_n5733 );
  nand     g05569 ( new_n5946 , new_n5696 , new_n5734 );
  nand     g05570 ( new_n5947 , new_n5945 , new_n5946 );
  xor      g05571 ( new_n5948 , new_n5944 , new_n5947 );
  nand     g05572 ( new_n5949 , pi057 , pi177 );
  nand     g05573 ( new_n5950 , pi182 , pi193 );
  xor      g05574 ( new_n5951 , new_n5949 , new_n5950 );
  nand     g05575 ( new_n5952 , pi048 , pi076 );
  nand     g05576 ( new_n5953 , new_n5731 , new_n5735 );
  or       g05577 ( new_n5954 , new_n5728 , new_n5737 );
  nand     g05578 ( new_n5955 , new_n5953 , new_n5954 );
  nand     g05579 ( new_n5956 , new_n5724 , new_n5725 );
  nand     g05580 ( new_n5957 , new_n5706 , new_n5726 );
  nand     g05581 ( new_n5958 , new_n5956 , new_n5957 );
  xor      g05582 ( new_n5959 , new_n5955 , new_n5958 );
  xor      g05583 ( new_n5960 , new_n5952 , new_n5959 );
  xor      g05584 ( new_n5961 , new_n5951 , new_n5960 );
  nand     g05585 ( new_n5962 , pi162 , pi192 );
  nor      g05586 ( new_n5963 , new_n5784 , new_n5806 );
  nor      g05587 ( new_n5964 , new_n5805 , new_n5807 );
  or       g05588 ( new_n5965 , new_n5963 , new_n5964 );
  xor      g05589 ( new_n5966 , new_n5962 , new_n5965 );
  xor      g05590 ( new_n5967 , new_n5961 , new_n5966 );
  nor      g05591 ( new_n5968 , new_n5573 , new_n5654 );
  and      g05592 ( new_n5969 , new_n5655 , new_n5671 );
  or       g05593 ( new_n5970 , new_n5968 , new_n5969 );
  nand     g05594 ( new_n5971 , pi086 , pi188 );
  nand     g05595 ( new_n5972 , new_n5538 , new_n5560 );
  nand     g05596 ( new_n5973 , new_n5561 , new_n5571 );
  nand     g05597 ( new_n5974 , new_n5972 , new_n5973 );
  xor      g05598 ( new_n5975 , new_n5971 , new_n5974 );
  xor      g05599 ( new_n5976 , new_n5970 , new_n5975 );
  xor      g05600 ( new_n5977 , new_n5967 , new_n5976 );
  nand     g05601 ( new_n5978 , pi216 , pi237 );
  xor      g05602 ( new_n5979 , new_n5977 , new_n5978 );
  xor      g05603 ( new_n5980 , new_n5948 , new_n5979 );
  xor      g05604 ( new_n5981 , new_n5941 , new_n5980 );
  nand     g05605 ( new_n5982 , pi001 , pi118 );
  nand     g05606 ( new_n5983 , pi123 , pi144 );
  nand     g05607 ( new_n5984 , pi007 , pi122 );
  xor      g05608 ( new_n5985 , new_n5983 , new_n5984 );
  nand     g05609 ( new_n5986 , pi108 , pi135 );
  nand     g05610 ( new_n5987 , pi043 , pi071 );
  xnor     g05611 ( new_n5988 , new_n5986 , new_n5987 );
  xor      g05612 ( new_n5989 , new_n5985 , new_n5988 );
  xor      g05613 ( new_n5990 , new_n5982 , new_n5989 );
  nand     g05614 ( new_n5991 , new_n5613 , new_n5614 );
  nand     g05615 ( new_n5992 , new_n5578 , new_n5615 );
  nand     g05616 ( new_n5993 , new_n5991 , new_n5992 );
  nand     g05617 ( new_n5994 , new_n5554 , new_n5555 );
  nand     g05618 ( new_n5995 , new_n5519 , new_n5556 );
  nand     g05619 ( new_n5996 , new_n5994 , new_n5995 );
  xnor     g05620 ( new_n5997 , new_n5993 , new_n5996 );
  xor      g05621 ( new_n5998 , new_n5990 , new_n5997 );
  nand     g05622 ( new_n5999 , new_n5896 , new_n5929 );
  nand g05623 ( new_n6000 , new_n5932 , new_n5932 );
  nand     g05624 ( new_n6001 , new_n5927 , new_n6000 );
  nand     g05625 ( new_n6002 , new_n5999 , new_n6001 );
  nand     g05626 ( new_n6003 , pi126 , pi142 );
  nand     g05627 ( new_n6004 , pi023 , pi061 );
  xnor     g05628 ( new_n6005 , new_n6003 , new_n6004 );
  nand     g05629 ( new_n6006 , pi038 , pi219 );
  xor      g05630 ( new_n6007 , new_n6005 , new_n6006 );
  xor      g05631 ( new_n6008 , new_n6002 , new_n6007 );
  nor      g05632 ( new_n6009 , new_n5612 , new_n5616 );
  and      g05633 ( new_n6010 , new_n5617 , new_n5624 );
  nor      g05634 ( new_n6011 , new_n6009 , new_n6010 );
  nand     g05635 ( new_n6012 , new_n5620 , new_n5621 );
  nand     g05636 ( new_n6013 , new_n5592 , new_n5622 );
  nand     g05637 ( new_n6014 , new_n6012 , new_n6013 );
  nand     g05638 ( new_n6015 , pi046 , pi160 );
  xor      g05639 ( new_n6016 , new_n6014 , new_n6015 );
  nor      g05640 ( new_n6017 , new_n5593 , new_n5618 );
  nor      g05641 ( new_n6018 , new_n5619 , new_n5623 );
  nor      g05642 ( new_n6019 , new_n6017 , new_n6018 );
  xor      g05643 ( new_n6020 , new_n6016 , new_n6019 );
  xor      g05644 ( new_n6021 , new_n6011 , new_n6020 );
  nand     g05645 ( new_n6022 , pi102 , pi113 );
  xor      g05646 ( new_n6023 , new_n6021 , new_n6022 );
  xor      g05647 ( new_n6024 , new_n6008 , new_n6023 );
  xor      g05648 ( new_n6025 , new_n5998 , new_n6024 );
  nand     g05649 ( new_n6026 , new_n5926 , new_n5933 );
  nand g05650 ( new_n6027 , new_n5923 , new_n5923 );
  nand     g05651 ( new_n6028 , new_n6027 , new_n5934 );
  nand     g05652 ( new_n6029 , new_n6026 , new_n6028 );
  nand     g05653 ( new_n6030 , pi042 , pi059 );
  xor      g05654 ( new_n6031 , new_n6029 , new_n6030 );
  nand     g05655 ( new_n6032 , pi041 , pi238 );
  nand     g05656 ( new_n6033 , pi137 , pi143 );
  nand     g05657 ( new_n6034 , pi028 , pi087 );
  xor      g05658 ( new_n6035 , new_n6033 , new_n6034 );
  xor      g05659 ( new_n6036 , new_n6032 , new_n6035 );
  xor      g05660 ( new_n6037 , new_n6031 , new_n6036 );
  xor      g05661 ( new_n6038 , new_n6025 , new_n6037 );
  xor      g05662 ( new_n6039 , new_n5981 , new_n6038 );
  xor      g05663 ( new_n6040 , new_n5851 , new_n6039 );
  xor      g05664 ( po021 , new_n5837 , new_n6040 );
  xor      g05665 ( po022 , new_n4914 , new_n4922 );
  xor      g05666 ( po023 , new_n2566 , new_n2604 );
  xnor     g05667 ( po024 , new_n1861 , new_n1868 );
  xnor     g05668 ( po025 , new_n4232 , new_n4233 );
  xor      g05669 ( po026 , new_n5487 , new_n5489 );
  nand     g05670 ( new_n6047 , pi153 , pi236 );
  nand     g05671 ( new_n6048 , pi120 , pi204 );
  nand     g05672 ( new_n6049 , pi053 , pi077 );
  nand     g05673 ( new_n6050 , pi030 , pi131 );
  nand     g05674 ( new_n6051 , new_n6049 , new_n6050 );
  nand     g05675 ( new_n6052 , pi052 , pi185 );
  xor      g05676 ( new_n6053 , new_n6049 , new_n6050 );
  nand     g05677 ( new_n6054 , new_n6052 , new_n6053 );
  nand     g05678 ( new_n6055 , new_n6051 , new_n6054 );
  xor      g05679 ( new_n6056 , new_n6048 , new_n6055 );
  nand     g05680 ( new_n6057 , pi212 , pi215 );
  nand     g05681 ( new_n6058 , pi165 , pi168 );
  or       g05682 ( new_n6059 , new_n3540 , new_n3543 );
  or       g05683 ( new_n6060 , new_n3544 , new_n3555 );
  nand     g05684 ( new_n6061 , new_n6059 , new_n6060 );
  nand     g05685 ( new_n6062 , new_n3552 , new_n3553 );
  nand     g05686 ( new_n6063 , new_n3549 , new_n3554 );
  nand     g05687 ( new_n6064 , new_n6062 , new_n6063 );
  nand     g05688 ( new_n6065 , pi139 , pi172 );
  nand     g05689 ( new_n6066 , pi198 , pi208 );
  nand     g05690 ( new_n6067 , new_n6065 , new_n6066 );
  nand     g05691 ( new_n6068 , pi139 , pi198 );
  nor      g05692 ( new_n6069 , new_n3553 , new_n6068 );
  nand g05693 ( new_n6070 , new_n6069 , new_n6069 );
  nand     g05694 ( new_n6071 , new_n6067 , new_n6070 );
  nand     g05695 ( new_n6072 , pi015 , pi062 );
  nand     g05696 ( new_n6073 , pi065 , pi204 );
  nand     g05697 ( new_n6074 , new_n6072 , new_n6073 );
  nand     g05698 ( new_n6075 , pi062 , pi204 );
  nor      g05699 ( new_n6076 , new_n3547 , new_n6075 );
  nand g05700 ( new_n6077 , new_n6076 , new_n6076 );
  nand     g05701 ( new_n6078 , new_n6074 , new_n6077 );
  nand     g05702 ( new_n6079 , pi035 , pi120 );
  nand     g05703 ( new_n6080 , new_n3546 , new_n3547 );
  nand     g05704 ( new_n6081 , new_n3545 , new_n3548 );
  nand     g05705 ( new_n6082 , new_n6080 , new_n6081 );
  xor      g05706 ( new_n6083 , new_n6079 , new_n6082 );
  xor      g05707 ( new_n6084 , new_n6078 , new_n6083 );
  xor      g05708 ( new_n6085 , new_n6071 , new_n6084 );
  xor      g05709 ( new_n6086 , new_n6064 , new_n6085 );
  xor      g05710 ( new_n6087 , new_n6061 , new_n6086 );
  nor      g05711 ( new_n6088 , new_n6058 , new_n6087 );
  nor      g05712 ( new_n6089 , new_n3539 , new_n3556 );
  xor      g05713 ( new_n6090 , new_n6058 , new_n6087 );
  and      g05714 ( new_n6091 , new_n6089 , new_n6090 );
  nor      g05715 ( new_n6092 , new_n6088 , new_n6091 );
  nand g05716 ( new_n6093 , new_n6061 , new_n6061 );
  nor      g05717 ( new_n6094 , new_n6093 , new_n6086 );
  nand     g05718 ( new_n6095 , new_n6079 , new_n6082 );
  nand     g05719 ( new_n6096 , new_n6078 , new_n6083 );
  nand     g05720 ( new_n6097 , new_n6095 , new_n6096 );
  nand     g05721 ( new_n6098 , pi168 , pi197 );
  nand     g05722 ( new_n6099 , pi165 , pi208 );
  xor      g05723 ( new_n6100 , new_n6098 , new_n6099 );
  xor      g05724 ( new_n6101 , new_n6068 , new_n6100 );
  xor      g05725 ( new_n6102 , new_n6097 , new_n6101 );
  nand     g05726 ( new_n6103 , pi035 , pi172 );
  xor      g05727 ( new_n6104 , new_n6077 , new_n6103 );
  nand     g05728 ( new_n6105 , pi015 , pi120 );
  nand     g05729 ( new_n6106 , pi065 , pi146 );
  xor      g05730 ( new_n6107 , new_n6105 , new_n6106 );
  xnor     g05731 ( new_n6108 , new_n6075 , new_n6107 );
  xnor     g05732 ( new_n6109 , new_n6104 , new_n6108 );
  xor      g05733 ( new_n6110 , new_n6102 , new_n6109 );
  nand     g05734 ( new_n6111 , new_n6071 , new_n6084 );
  nand     g05735 ( new_n6112 , new_n6064 , new_n6085 );
  nand     g05736 ( new_n6113 , new_n6111 , new_n6112 );
  xor      g05737 ( new_n6114 , new_n6070 , new_n6113 );
  xor      g05738 ( new_n6115 , new_n6110 , new_n6114 );
  xor      g05739 ( new_n6116 , new_n6094 , new_n6115 );
  xor      g05740 ( new_n6117 , new_n6092 , new_n6116 );
  nand g05741 ( new_n6118 , new_n6117 , new_n6117 );
  and      g05742 ( new_n6119 , new_n3585 , new_n3602 );
  nor      g05743 ( new_n6120 , new_n3586 , new_n3589 );
  and      g05744 ( new_n6121 , new_n3590 , new_n3601 );
  nor      g05745 ( new_n6122 , new_n6120 , new_n6121 );
  nand     g05746 ( new_n6123 , pi047 , pi254 );
  nand     g05747 ( new_n6124 , pi090 , pi158 );
  nand     g05748 ( new_n6125 , new_n6123 , new_n6124 );
  nand     g05749 ( new_n6126 , pi047 , pi158 );
  or       g05750 ( new_n6127 , new_n3593 , new_n6126 );
  nand     g05751 ( new_n6128 , new_n6125 , new_n6127 );
  nand     g05752 ( new_n6129 , pi089 , pi141 );
  nand     g05753 ( new_n6130 , new_n3592 , new_n3593 );
  nand     g05754 ( new_n6131 , new_n3591 , new_n3594 );
  nand     g05755 ( new_n6132 , new_n6130 , new_n6131 );
  xor      g05756 ( new_n6133 , new_n6129 , new_n6132 );
  xor      g05757 ( new_n6134 , new_n6128 , new_n6133 );
  and      g05758 ( new_n6135 , new_n3598 , new_n3599 );
  nor      g05759 ( new_n6136 , new_n3595 , new_n3600 );
  or       g05760 ( new_n6137 , new_n6135 , new_n6136 );
  nand     g05761 ( new_n6138 , pi154 , pi161 );
  nand     g05762 ( new_n6139 , pi095 , pi241 );
  and      g05763 ( new_n6140 , new_n6138 , new_n6139 );
  nand     g05764 ( new_n6141 , pi095 , pi161 );
  nor      g05765 ( new_n6142 , new_n3599 , new_n6141 );
  nor      g05766 ( new_n6143 , new_n6140 , new_n6142 );
  xor      g05767 ( new_n6144 , new_n6137 , new_n6143 );
  xor      g05768 ( new_n6145 , new_n6134 , new_n6144 );
  xor      g05769 ( new_n6146 , new_n6122 , new_n6145 );
  nand     g05770 ( new_n6147 , pi006 , pi236 );
  xor      g05771 ( new_n6148 , new_n6146 , new_n6147 );
  xnor     g05772 ( new_n6149 , new_n6119 , new_n6148 );
  nand     g05773 ( new_n6150 , new_n3563 , new_n3580 );
  nand     g05774 ( new_n6151 , pi124 , pi213 );
  nand     g05775 ( new_n6152 , new_n3575 , new_n3578 );
  nand     g05776 ( new_n6153 , new_n3574 , new_n3579 );
  nand     g05777 ( new_n6154 , new_n6152 , new_n6153 );
  nand     g05778 ( new_n6155 , new_n3569 , new_n3572 );
  nand     g05779 ( new_n6156 , new_n3568 , new_n3573 );
  nand     g05780 ( new_n6157 , new_n6155 , new_n6156 );
  nand     g05781 ( new_n6158 , pi130 , pi212 );
  nand     g05782 ( new_n6159 , pi003 , pi104 );
  and      g05783 ( new_n6160 , new_n6158 , new_n6159 );
  nand     g05784 ( new_n6161 , pi104 , pi130 );
  nor      g05785 ( new_n6162 , new_n3569 , new_n6161 );
  or       g05786 ( new_n6163 , new_n6160 , new_n6162 );
  nand     g05787 ( new_n6164 , new_n3565 , new_n3566 );
  nand     g05788 ( new_n6165 , new_n3564 , new_n3567 );
  nand     g05789 ( new_n6166 , new_n6164 , new_n6165 );
  nand     g05790 ( new_n6167 , pi013 , pi073 );
  nand     g05791 ( new_n6168 , pi004 , pi112 );
  nand     g05792 ( new_n6169 , pi105 , pi170 );
  nand     g05793 ( new_n6170 , new_n6168 , new_n6169 );
  nand     g05794 ( new_n6171 , pi004 , pi105 );
  or       g05795 ( new_n6172 , new_n3565 , new_n6171 );
  nand     g05796 ( new_n6173 , new_n6170 , new_n6172 );
  xor      g05797 ( new_n6174 , new_n6167 , new_n6173 );
  xor      g05798 ( new_n6175 , new_n6166 , new_n6174 );
  xor      g05799 ( new_n6176 , new_n6163 , new_n6175 );
  xor      g05800 ( new_n6177 , new_n6157 , new_n6176 );
  xnor     g05801 ( new_n6178 , new_n6154 , new_n6177 );
  xnor     g05802 ( new_n6179 , new_n6151 , new_n6178 );
  xnor     g05803 ( new_n6180 , new_n6150 , new_n6179 );
  nor      g05804 ( new_n6181 , new_n6149 , new_n6180 );
  nor      g05805 ( new_n6182 , new_n3584 , new_n3603 );
  nor      g05806 ( new_n6183 , new_n3581 , new_n3604 );
  or       g05807 ( new_n6184 , new_n6182 , new_n6183 );
  xnor     g05808 ( new_n6185 , new_n6149 , new_n6180 );
  nor      g05809 ( new_n6186 , new_n6184 , new_n6185 );
  nor      g05810 ( new_n6187 , new_n6181 , new_n6186 );
  nor      g05811 ( new_n6188 , new_n6154 , new_n6177 );
  nand     g05812 ( new_n6189 , pi213 , pi215 );
  nand     g05813 ( new_n6190 , pi124 , pi212 );
  xor      g05814 ( new_n6191 , new_n6161 , new_n6190 );
  xor      g05815 ( new_n6192 , new_n6189 , new_n6191 );
  nand     g05816 ( new_n6193 , new_n6167 , new_n6173 );
  nand     g05817 ( new_n6194 , new_n6166 , new_n6174 );
  nand     g05818 ( new_n6195 , new_n6193 , new_n6194 );
  xor      g05819 ( new_n6196 , new_n6192 , new_n6195 );
  nand     g05820 ( new_n6197 , pi170 , pi183 );
  nand     g05821 ( new_n6198 , pi073 , pi112 );
  xor      g05822 ( new_n6199 , new_n6197 , new_n6198 );
  xor      g05823 ( new_n6200 , new_n6171 , new_n6199 );
  nand     g05824 ( new_n6201 , pi003 , pi013 );
  xnor     g05825 ( new_n6202 , new_n6172 , new_n6201 );
  xnor     g05826 ( new_n6203 , new_n6200 , new_n6202 );
  xor      g05827 ( new_n6204 , new_n6196 , new_n6203 );
  nand g05828 ( new_n6205 , new_n6176 , new_n6176 );
  nor      g05829 ( new_n6206 , new_n6157 , new_n6205 );
  nand     g05830 ( new_n6207 , new_n6162 , new_n6206 );
  nor      g05831 ( new_n6208 , new_n6163 , new_n6175 );
  or       g05832 ( new_n6209 , new_n6162 , new_n6208 );
  or       g05833 ( new_n6210 , new_n6206 , new_n6209 );
  nand     g05834 ( new_n6211 , new_n6207 , new_n6210 );
  xor      g05835 ( new_n6212 , new_n6204 , new_n6211 );
  xor      g05836 ( new_n6213 , new_n6188 , new_n6212 );
  nor      g05837 ( new_n6214 , new_n6151 , new_n6178 );
  nor      g05838 ( new_n6215 , new_n6150 , new_n6179 );
  nor      g05839 ( new_n6216 , new_n6214 , new_n6215 );
  xor      g05840 ( new_n6217 , new_n6213 , new_n6216 );
  xor      g05841 ( new_n6218 , new_n6187 , new_n6217 );
  nor      g05842 ( new_n6219 , new_n6146 , new_n6147 );
  and      g05843 ( new_n6220 , new_n6119 , new_n6148 );
  nor      g05844 ( new_n6221 , new_n6219 , new_n6220 );
  nand g05845 ( new_n6222 , new_n6145 , new_n6145 );
  nor      g05846 ( new_n6223 , new_n6122 , new_n6222 );
  nand g05847 ( new_n6224 , new_n6143 , new_n6143 );
  nand     g05848 ( new_n6225 , new_n6137 , new_n6224 );
  nand g05849 ( new_n6226 , new_n6134 , new_n6134 );
  or       g05850 ( new_n6227 , new_n6226 , new_n6144 );
  nand     g05851 ( new_n6228 , new_n6225 , new_n6227 );
  xor      g05852 ( new_n6229 , new_n6142 , new_n6228 );
  nand     g05853 ( new_n6230 , pi006 , pi241 );
  nand     g05854 ( new_n6231 , pi209 , pi236 );
  xor      g05855 ( new_n6232 , new_n6230 , new_n6231 );
  xnor     g05856 ( new_n6233 , new_n6141 , new_n6232 );
  nand     g05857 ( new_n6234 , new_n6129 , new_n6132 );
  nand     g05858 ( new_n6235 , new_n6128 , new_n6133 );
  nand     g05859 ( new_n6236 , new_n6234 , new_n6235 );
  xor      g05860 ( new_n6237 , new_n6233 , new_n6236 );
  nand     g05861 ( new_n6238 , pi141 , pi154 );
  xor      g05862 ( new_n6239 , new_n6127 , new_n6238 );
  nand     g05863 ( new_n6240 , pi089 , pi090 );
  nand     g05864 ( new_n6241 , pi018 , pi254 );
  xor      g05865 ( new_n6242 , new_n6240 , new_n6241 );
  xor      g05866 ( new_n6243 , new_n6126 , new_n6242 );
  xor      g05867 ( new_n6244 , new_n6239 , new_n6243 );
  xor      g05868 ( new_n6245 , new_n6237 , new_n6244 );
  xor      g05869 ( new_n6246 , new_n6229 , new_n6245 );
  xor      g05870 ( new_n6247 , new_n6223 , new_n6246 );
  xor      g05871 ( new_n6248 , new_n6221 , new_n6247 );
  xnor     g05872 ( new_n6249 , new_n6218 , new_n6248 );
  nand     g05873 ( new_n6250 , new_n6118 , new_n6249 );
  xor      g05874 ( new_n6251 , new_n6117 , new_n6249 );
  nand g05875 ( new_n6252 , new_n6251 , new_n6251 );
  xnor     g05876 ( new_n6253 , new_n6089 , new_n6090 );
  xnor     g05877 ( new_n6254 , new_n6184 , new_n6185 );
  nor      g05878 ( new_n6255 , new_n6253 , new_n6254 );
  nand     g05879 ( new_n6256 , new_n3557 , new_n3560 );
  nand     g05880 ( new_n6257 , new_n3561 , new_n3605 );
  and      g05881 ( new_n6258 , new_n6256 , new_n6257 );
  xnor     g05882 ( new_n6259 , new_n6253 , new_n6254 );
  nor      g05883 ( new_n6260 , new_n6258 , new_n6259 );
  nor      g05884 ( new_n6261 , new_n6255 , new_n6260 );
  nand     g05885 ( new_n6262 , new_n6252 , new_n6261 );
  nand     g05886 ( new_n6263 , new_n6250 , new_n6262 );
  nand     g05887 ( new_n6264 , pi064 , pi229 );
  nand g05888 ( new_n6265 , new_n6094 , new_n6094 );
  nor      g05889 ( new_n6266 , new_n6265 , new_n6115 );
  nor      g05890 ( new_n6267 , new_n6092 , new_n6116 );
  or       g05891 ( new_n6268 , new_n6266 , new_n6267 );
  xor      g05892 ( new_n6269 , new_n6264 , new_n6268 );
  nand     g05893 ( new_n6270 , pi084 , pi092 );
  nand     g05894 ( new_n6271 , new_n6097 , new_n6101 );
  nand     g05895 ( new_n6272 , new_n6102 , new_n6109 );
  nand     g05896 ( new_n6273 , new_n6271 , new_n6272 );
  xor      g05897 ( new_n6274 , new_n6270 , new_n6273 );
  xnor     g05898 ( new_n6275 , new_n6269 , new_n6274 );
  xor      g05899 ( new_n6276 , new_n6263 , new_n6275 );
  xor      g05900 ( new_n6277 , new_n6057 , new_n6276 );
  nand     g05901 ( new_n6278 , pi133 , pi229 );
  nand     g05902 ( new_n6279 , new_n3520 , new_n3521 );
  nand     g05903 ( new_n6280 , new_n3519 , new_n3522 );
  nand     g05904 ( new_n6281 , new_n6279 , new_n6280 );
  nand     g05905 ( new_n6282 , new_n6278 , new_n6281 );
  nand     g05906 ( new_n6283 , pi064 , pi092 );
  or       g05907 ( new_n6284 , new_n3520 , new_n6283 );
  nand     g05908 ( new_n6285 , pi092 , pi189 );
  nand     g05909 ( new_n6286 , pi064 , pi190 );
  nand     g05910 ( new_n6287 , new_n6285 , new_n6286 );
  nand     g05911 ( new_n6288 , new_n6284 , new_n6287 );
  xor      g05912 ( new_n6289 , new_n6278 , new_n6281 );
  nand     g05913 ( new_n6290 , new_n6288 , new_n6289 );
  nand     g05914 ( new_n6291 , new_n6282 , new_n6290 );
  xor      g05915 ( new_n6292 , new_n6052 , new_n6053 );
  nand     g05916 ( new_n6293 , new_n6291 , new_n6292 );
  nand     g05917 ( new_n6294 , pi067 , pi133 );
  xor      g05918 ( new_n6295 , new_n6284 , new_n6294 );
  nand     g05919 ( new_n6296 , pi189 , pi229 );
  nand     g05920 ( new_n6297 , pi084 , pi190 );
  xor      g05921 ( new_n6298 , new_n6296 , new_n6297 );
  xnor     g05922 ( new_n6299 , new_n6283 , new_n6298 );
  xor      g05923 ( new_n6300 , new_n6295 , new_n6299 );
  xor      g05924 ( new_n6301 , new_n6291 , new_n6292 );
  nand g05925 ( new_n6302 , new_n6301 , new_n6301 );
  or       g05926 ( new_n6303 , new_n6300 , new_n6302 );
  nand     g05927 ( new_n6304 , new_n6293 , new_n6303 );
  nand     g05928 ( new_n6305 , pi062 , pi146 );
  xor      g05929 ( new_n6306 , new_n6304 , new_n6305 );
  nor      g05930 ( new_n6307 , new_n6070 , new_n6113 );
  nand g05931 ( new_n6308 , new_n6114 , new_n6114 );
  nor      g05932 ( new_n6309 , new_n6110 , new_n6308 );
  nor      g05933 ( new_n6310 , new_n6307 , new_n6309 );
  nand g05934 ( new_n6311 , new_n6223 , new_n6223 );
  nor      g05935 ( new_n6312 , new_n6311 , new_n6246 );
  nor      g05936 ( new_n6313 , new_n6221 , new_n6247 );
  or       g05937 ( new_n6314 , new_n6312 , new_n6313 );
  nand     g05938 ( new_n6315 , pi030 , pi052 );
  nand     g05939 ( new_n6316 , pi077 , pi185 );
  or       g05940 ( new_n6317 , new_n6284 , new_n6294 );
  nand     g05941 ( new_n6318 , new_n6295 , new_n6299 );
  nand     g05942 ( new_n6319 , new_n6317 , new_n6318 );
  xor      g05943 ( new_n6320 , new_n6316 , new_n6319 );
  xor      g05944 ( new_n6321 , new_n6315 , new_n6320 );
  xor      g05945 ( new_n6322 , new_n6314 , new_n6321 );
  xor      g05946 ( new_n6323 , new_n6310 , new_n6322 );
  xor      g05947 ( new_n6324 , new_n6306 , new_n6323 );
  xor      g05948 ( new_n6325 , new_n6277 , new_n6324 );
  xor      g05949 ( new_n6326 , new_n6056 , new_n6325 );
  xor      g05950 ( new_n6327 , new_n6047 , new_n6326 );
  nand     g05951 ( new_n6328 , pi018 , pi158 );
  nand     g05952 ( new_n6329 , pi006 , pi161 );
  nand     g05953 ( new_n6330 , pi088 , pi170 );
  xor      g05954 ( new_n6331 , new_n6329 , new_n6330 );
  xor      g05955 ( new_n6332 , new_n6328 , new_n6331 );
  or       g05956 ( new_n6333 , new_n6077 , new_n6103 );
  nand     g05957 ( new_n6334 , new_n6104 , new_n6108 );
  nand     g05958 ( new_n6335 , new_n6333 , new_n6334 );
  nand     g05959 ( new_n6336 , pi067 , pi189 );
  xor      g05960 ( new_n6337 , new_n6251 , new_n6261 );
  nand g05961 ( new_n6338 , new_n3518 , new_n3518 );
  nand     g05962 ( new_n6339 , new_n6338 , new_n3535 );
  nand     g05963 ( new_n6340 , pi131 , pi185 );
  nand     g05964 ( new_n6341 , new_n6339 , new_n6340 );
  nand g05965 ( new_n6342 , new_n6341 , new_n6341 );
  nor      g05966 ( new_n6343 , new_n3530 , new_n3533 );
  nor      g05967 ( new_n6344 , new_n3529 , new_n3534 );
  nor      g05968 ( new_n6345 , new_n6343 , new_n6344 );
  nand     g05969 ( new_n6346 , new_n3526 , new_n3527 );
  nand     g05970 ( new_n6347 , new_n3523 , new_n3528 );
  nand     g05971 ( new_n6348 , new_n6346 , new_n6347 );
  nand     g05972 ( new_n6349 , pi067 , pi077 );
  nand     g05973 ( new_n6350 , pi052 , pi053 );
  and      g05974 ( new_n6351 , new_n6349 , new_n6350 );
  nor      g05975 ( new_n6352 , new_n3527 , new_n6049 );
  or       g05976 ( new_n6353 , new_n6351 , new_n6352 );
  xor      g05977 ( new_n6354 , new_n6288 , new_n6289 );
  xor      g05978 ( new_n6355 , new_n6353 , new_n6354 );
  xor      g05979 ( new_n6356 , new_n6348 , new_n6355 );
  xor      g05980 ( new_n6357 , new_n6345 , new_n6356 );
  xnor     g05981 ( new_n6358 , new_n6339 , new_n6340 );
  nor      g05982 ( new_n6359 , new_n6357 , new_n6358 );
  nor      g05983 ( new_n6360 , new_n6342 , new_n6359 );
  nand g05984 ( new_n6361 , new_n6360 , new_n6360 );
  nor      g05985 ( new_n6362 , new_n6345 , new_n6356 );
  xor      g05986 ( new_n6363 , new_n6300 , new_n6302 );
  nor      g05987 ( new_n6364 , new_n6353 , new_n6354 );
  nand g05988 ( new_n6365 , new_n6355 , new_n6355 );
  nor      g05989 ( new_n6366 , new_n6348 , new_n6365 );
  xor      g05990 ( new_n6367 , new_n6352 , new_n6366 );
  nor      g05991 ( new_n6368 , new_n6364 , new_n6367 );
  xor      g05992 ( new_n6369 , new_n6363 , new_n6368 );
  or       g05993 ( new_n6370 , new_n6362 , new_n6369 );
  nand     g05994 ( new_n6371 , new_n6362 , new_n6369 );
  nand     g05995 ( new_n6372 , new_n6370 , new_n6371 );
  xor      g05996 ( new_n6373 , new_n6361 , new_n6372 );
  nand     g05997 ( new_n6374 , new_n6337 , new_n6373 );
  xor      g05998 ( new_n6375 , new_n6357 , new_n6358 );
  xnor     g05999 ( new_n6376 , new_n6258 , new_n6259 );
  or       g06000 ( new_n6377 , new_n6375 , new_n6376 );
  and      g06001 ( new_n6378 , new_n3516 , new_n3536 );
  nor      g06002 ( new_n6379 , new_n3537 , new_n3606 );
  nor      g06003 ( new_n6380 , new_n6378 , new_n6379 );
  xor      g06004 ( new_n6381 , new_n6375 , new_n6376 );
  nand     g06005 ( new_n6382 , new_n6380 , new_n6381 );
  nand     g06006 ( new_n6383 , new_n6377 , new_n6382 );
  xor      g06007 ( new_n6384 , new_n6337 , new_n6373 );
  nand     g06008 ( new_n6385 , new_n6383 , new_n6384 );
  nand     g06009 ( new_n6386 , new_n6374 , new_n6385 );
  xor      g06010 ( new_n6387 , new_n6336 , new_n6386 );
  and      g06011 ( new_n6388 , new_n6352 , new_n6366 );
  nor      g06012 ( new_n6389 , new_n6363 , new_n6368 );
  nor      g06013 ( new_n6390 , new_n6388 , new_n6389 );
  nand     g06014 ( new_n6391 , pi131 , pi220 );
  xor      g06015 ( new_n6392 , new_n6390 , new_n6391 );
  xor      g06016 ( new_n6393 , new_n6387 , new_n6392 );
  nand     g06017 ( new_n6394 , new_n6361 , new_n6371 );
  nand     g06018 ( new_n6395 , new_n6370 , new_n6394 );
  nand     g06019 ( new_n6396 , new_n6230 , new_n6231 );
  nand     g06020 ( new_n6397 , new_n6141 , new_n6232 );
  nand     g06021 ( new_n6398 , new_n6396 , new_n6397 );
  nand g06022 ( new_n6399 , new_n6236 , new_n6236 );
  nor      g06023 ( new_n6400 , new_n6233 , new_n6399 );
  nand g06024 ( new_n6401 , new_n6244 , new_n6244 );
  nor      g06025 ( new_n6402 , new_n6237 , new_n6401 );
  nor      g06026 ( new_n6403 , new_n6400 , new_n6402 );
  xor      g06027 ( new_n6404 , new_n6398 , new_n6403 );
  xor      g06028 ( new_n6405 , new_n6395 , new_n6404 );
  nand     g06029 ( new_n6406 , pi197 , pi208 );
  nand     g06030 ( new_n6407 , pi013 , pi130 );
  xor      g06031 ( new_n6408 , new_n6406 , new_n6407 );
  nand     g06032 ( new_n6409 , new_n6296 , new_n6297 );
  nand     g06033 ( new_n6410 , new_n6283 , new_n6298 );
  nand     g06034 ( new_n6411 , new_n6409 , new_n6410 );
  nand     g06035 ( new_n6412 , new_n6161 , new_n6190 );
  nand     g06036 ( new_n6413 , new_n6189 , new_n6191 );
  nand     g06037 ( new_n6414 , new_n6412 , new_n6413 );
  xor      g06038 ( new_n6415 , new_n6411 , new_n6414 );
  nand     g06039 ( new_n6416 , new_n6197 , new_n6198 );
  nand     g06040 ( new_n6417 , new_n6171 , new_n6199 );
  nand     g06041 ( new_n6418 , new_n6416 , new_n6417 );
  nor      g06042 ( new_n6419 , new_n6172 , new_n6201 );
  nor      g06043 ( new_n6420 , new_n6200 , new_n6202 );
  nor      g06044 ( new_n6421 , new_n6419 , new_n6420 );
  nand     g06045 ( new_n6422 , pi003 , pi112 );
  xor      g06046 ( new_n6423 , new_n6421 , new_n6422 );
  xor      g06047 ( new_n6424 , new_n6418 , new_n6423 );
  xor      g06048 ( new_n6425 , new_n6415 , new_n6424 );
  xor      g06049 ( new_n6426 , new_n6408 , new_n6425 );
  xor      g06050 ( new_n6427 , new_n6405 , new_n6426 );
  nand     g06051 ( new_n6428 , pi035 , pi198 );
  nand     g06052 ( new_n6429 , pi015 , pi172 );
  xor      g06053 ( new_n6430 , new_n6428 , new_n6429 );
  nand     g06054 ( new_n6431 , pi128 , pi254 );
  nand     g06055 ( new_n6432 , pi047 , pi089 );
  xor      g06056 ( new_n6433 , new_n6431 , new_n6432 );
  nor      g06057 ( new_n6434 , new_n6127 , new_n6238 );
  nand g06058 ( new_n6435 , new_n6239 , new_n6239 );
  nor      g06059 ( new_n6436 , new_n6435 , new_n6243 );
  nor      g06060 ( new_n6437 , new_n6434 , new_n6436 );
  nand     g06061 ( new_n6438 , pi004 , pi183 );
  xor      g06062 ( new_n6439 , new_n6437 , new_n6438 );
  xor      g06063 ( new_n6440 , new_n6433 , new_n6439 );
  xor      g06064 ( new_n6441 , new_n6430 , new_n6440 );
  xor      g06065 ( new_n6442 , new_n6427 , new_n6441 );
  and      g06066 ( new_n6443 , new_n6188 , new_n6212 );
  nand g06067 ( new_n6444 , new_n6213 , new_n6213 );
  nor      g06068 ( new_n6445 , new_n6444 , new_n6216 );
  nor      g06069 ( new_n6446 , new_n6443 , new_n6445 );
  xor      g06070 ( new_n6447 , new_n6442 , new_n6446 );
  nor      g06071 ( new_n6448 , new_n6187 , new_n6217 );
  and      g06072 ( new_n6449 , new_n6218 , new_n6248 );
  nor      g06073 ( new_n6450 , new_n6448 , new_n6449 );
  nand     g06074 ( new_n6451 , pi034 , pi190 );
  nand     g06075 ( new_n6452 , new_n6105 , new_n6106 );
  nand     g06076 ( new_n6453 , new_n6075 , new_n6107 );
  nand     g06077 ( new_n6454 , new_n6452 , new_n6453 );
  nand     g06078 ( new_n6455 , pi139 , pi165 );
  xor      g06079 ( new_n6456 , new_n6454 , new_n6455 );
  xor      g06080 ( new_n6457 , new_n6451 , new_n6456 );
  xor      g06081 ( new_n6458 , new_n6450 , new_n6457 );
  nand     g06082 ( new_n6459 , pi065 , pi152 );
  nand     g06083 ( new_n6460 , pi209 , pi241 );
  xor      g06084 ( new_n6461 , new_n6459 , new_n6460 );
  xor      g06085 ( new_n6462 , new_n6458 , new_n6461 );
  xor      g06086 ( new_n6463 , new_n6447 , new_n6462 );
  nand g06087 ( new_n6464 , new_n6204 , new_n6204 );
  nand     g06088 ( new_n6465 , new_n6464 , new_n6210 );
  nand     g06089 ( new_n6466 , new_n6207 , new_n6465 );
  nand     g06090 ( new_n6467 , pi095 , pi141 );
  nand     g06091 ( new_n6468 , pi090 , pi154 );
  xor      g06092 ( new_n6469 , new_n6467 , new_n6468 );
  xor      g06093 ( new_n6470 , new_n6466 , new_n6469 );
  nand g06094 ( new_n6471 , new_n6228 , new_n6228 );
  nand     g06095 ( new_n6472 , new_n6142 , new_n6471 );
  nand g06096 ( new_n6473 , new_n6229 , new_n6229 );
  nand     g06097 ( new_n6474 , new_n6473 , new_n6245 );
  nand     g06098 ( new_n6475 , new_n6472 , new_n6474 );
  nand     g06099 ( new_n6476 , new_n6192 , new_n6195 );
  nand     g06100 ( new_n6477 , new_n6196 , new_n6203 );
  nand     g06101 ( new_n6478 , new_n6476 , new_n6477 );
  nand     g06102 ( new_n6479 , pi053 , pi133 );
  nand     g06103 ( new_n6480 , pi073 , pi105 );
  xor      g06104 ( new_n6481 , new_n6479 , new_n6480 );
  nand     g06105 ( new_n6482 , pi078 , pi168 );
  nand     g06106 ( new_n6483 , new_n6098 , new_n6099 );
  nand     g06107 ( new_n6484 , new_n6068 , new_n6100 );
  nand     g06108 ( new_n6485 , new_n6483 , new_n6484 );
  xor      g06109 ( new_n6486 , new_n6482 , new_n6485 );
  xnor     g06110 ( new_n6487 , new_n6481 , new_n6486 );
  xor      g06111 ( new_n6488 , new_n6478 , new_n6487 );
  nand     g06112 ( new_n6489 , new_n6240 , new_n6241 );
  nand     g06113 ( new_n6490 , new_n6126 , new_n6242 );
  nand     g06114 ( new_n6491 , new_n6489 , new_n6490 );
  nand     g06115 ( new_n6492 , pi022 , pi213 );
  xnor     g06116 ( new_n6493 , new_n6491 , new_n6492 );
  nand     g06117 ( new_n6494 , pi104 , pi124 );
  xor      g06118 ( new_n6495 , new_n6493 , new_n6494 );
  xor      g06119 ( new_n6496 , new_n6488 , new_n6495 );
  xor      g06120 ( new_n6497 , new_n6475 , new_n6496 );
  xor      g06121 ( new_n6498 , new_n6470 , new_n6497 );
  xor      g06122 ( new_n6499 , new_n6463 , new_n6498 );
  xor      g06123 ( new_n6500 , new_n6393 , new_n6499 );
  xor      g06124 ( new_n6501 , new_n6335 , new_n6500 );
  xor      g06125 ( new_n6502 , new_n6332 , new_n6501 );
  xor      g06126 ( po027 , new_n6327 , new_n6502 );
  and      g06127 ( new_n6504 , new_n4881 , new_n4903 );
  nor      g06128 ( new_n6505 , new_n4841 , new_n4904 );
  nor      g06129 ( new_n6506 , new_n6504 , new_n6505 );
  nand     g06130 ( new_n6507 , new_n4867 , new_n4870 );
  nand     g06131 ( new_n6508 , new_n4866 , new_n4871 );
  nand     g06132 ( new_n6509 , new_n6507 , new_n6508 );
  nand     g06133 ( new_n6510 , pi048 , pi139 );
  nand     g06134 ( new_n6511 , pi208 , pi237 );
  and      g06135 ( new_n6512 , new_n6510 , new_n6511 );
  nand     g06136 ( new_n6513 , pi139 , pi237 );
  nor      g06137 ( new_n6514 , new_n4867 , new_n6513 );
  nor      g06138 ( new_n6515 , new_n6512 , new_n6514 );
  nand     g06139 ( new_n6516 , new_n4863 , new_n4864 );
  nand     g06140 ( new_n6517 , new_n4862 , new_n4865 );
  nand     g06141 ( new_n6518 , new_n6516 , new_n6517 );
  nand     g06142 ( new_n6519 , pi035 , pi179 );
  nand     g06143 ( new_n6520 , pi015 , pi033 );
  nand     g06144 ( new_n6521 , pi162 , pi204 );
  nand     g06145 ( new_n6522 , new_n6520 , new_n6521 );
  nand     g06146 ( new_n6523 , pi033 , pi204 );
  nor      g06147 ( new_n6524 , new_n4864 , new_n6523 );
  nand g06148 ( new_n6525 , new_n6524 , new_n6524 );
  nand     g06149 ( new_n6526 , new_n6522 , new_n6525 );
  xor      g06150 ( new_n6527 , new_n6519 , new_n6526 );
  xor      g06151 ( new_n6528 , new_n6518 , new_n6527 );
  xor      g06152 ( new_n6529 , new_n6515 , new_n6528 );
  xor      g06153 ( new_n6530 , new_n6509 , new_n6529 );
  nand g06154 ( new_n6531 , new_n6530 , new_n6530 );
  nor      g06155 ( new_n6532 , new_n4873 , new_n4878 );
  nor      g06156 ( new_n6533 , new_n4872 , new_n4879 );
  nor      g06157 ( new_n6534 , new_n6532 , new_n6533 );
  xor      g06158 ( new_n6535 , new_n6531 , new_n6534 );
  nand g06159 ( new_n6536 , new_n4861 , new_n4861 );
  or       g06160 ( new_n6537 , new_n6536 , new_n4880 );
  nand     g06161 ( new_n6538 , pi168 , pi238 );
  xnor     g06162 ( new_n6539 , new_n6537 , new_n6538 );
  xnor     g06163 ( new_n6540 , new_n6535 , new_n6539 );
  xor      g06164 ( new_n6541 , new_n6506 , new_n6540 );
  nand g06165 ( new_n6542 , new_n4839 , new_n4839 );
  nor      g06166 ( new_n6543 , new_n4820 , new_n6542 );
  nor      g06167 ( new_n6544 , new_n4801 , new_n4840 );
  or       g06168 ( new_n6545 , new_n6543 , new_n6544 );
  nor      g06169 ( new_n6546 , new_n4803 , new_n4806 );
  and      g06170 ( new_n6547 , new_n4807 , new_n4818 );
  nor      g06171 ( new_n6548 , new_n6546 , new_n6547 );
  nand     g06172 ( new_n6549 , new_n4813 , new_n4816 );
  nand     g06173 ( new_n6550 , new_n4812 , new_n4817 );
  nand     g06174 ( new_n6551 , new_n6549 , new_n6550 );
  nand     g06175 ( new_n6552 , pi108 , pi141 );
  nand     g06176 ( new_n6553 , new_n4809 , new_n4810 );
  nand     g06177 ( new_n6554 , new_n4808 , new_n4811 );
  nand     g06178 ( new_n6555 , new_n6553 , new_n6554 );
  xnor     g06179 ( new_n6556 , new_n6552 , new_n6555 );
  nand     g06180 ( new_n6557 , pi042 , pi090 );
  nand     g06181 ( new_n6558 , pi047 , pi051 );
  nand     g06182 ( new_n6559 , new_n6557 , new_n6558 );
  nand     g06183 ( new_n6560 , pi042 , pi047 );
  nor      g06184 ( new_n6561 , new_n4810 , new_n6560 );
  nand g06185 ( new_n6562 , new_n6561 , new_n6561 );
  nand     g06186 ( new_n6563 , new_n6559 , new_n6562 );
  xnor     g06187 ( new_n6564 , new_n6556 , new_n6563 );
  nand     g06188 ( new_n6565 , pi118 , pi161 );
  nor      g06189 ( new_n6566 , new_n4813 , new_n6565 );
  nand     g06190 ( new_n6567 , pi007 , pi161 );
  nand     g06191 ( new_n6568 , pi118 , pi241 );
  and      g06192 ( new_n6569 , new_n6567 , new_n6568 );
  or       g06193 ( new_n6570 , new_n6566 , new_n6569 );
  xnor     g06194 ( new_n6571 , new_n6564 , new_n6570 );
  xor      g06195 ( new_n6572 , new_n6551 , new_n6571 );
  nand g06196 ( new_n6573 , new_n6572 , new_n6572 );
  xor      g06197 ( new_n6574 , new_n6548 , new_n6573 );
  nand     g06198 ( new_n6575 , new_n4802 , new_n4819 );
  nand     g06199 ( new_n6576 , pi113 , pi236 );
  xnor     g06200 ( new_n6577 , new_n6575 , new_n6576 );
  xnor     g06201 ( new_n6578 , new_n6574 , new_n6577 );
  nand     g06202 ( new_n6579 , new_n4821 , new_n4838 );
  nand     g06203 ( new_n6580 , pi098 , pi213 );
  nand     g06204 ( new_n6581 , pi012 , pi104 );
  nand     g06205 ( new_n6582 , pi144 , pi212 );
  and      g06206 ( new_n6583 , new_n6581 , new_n6582 );
  nand     g06207 ( new_n6584 , pi104 , pi144 );
  nor      g06208 ( new_n6585 , new_n4832 , new_n6584 );
  or       g06209 ( new_n6586 , new_n6583 , new_n6585 );
  nand     g06210 ( new_n6587 , new_n4828 , new_n4829 );
  nand     g06211 ( new_n6588 , new_n4827 , new_n4830 );
  nand     g06212 ( new_n6589 , new_n6587 , new_n6588 );
  nand     g06213 ( new_n6590 , pi013 , pi061 );
  nand     g06214 ( new_n6591 , pi105 , pi188 );
  nand     g06215 ( new_n6592 , pi112 , pi178 );
  nand     g06216 ( new_n6593 , new_n6591 , new_n6592 );
  nand     g06217 ( new_n6594 , pi105 , pi178 );
  or       g06218 ( new_n6595 , new_n4827 , new_n6594 );
  nand     g06219 ( new_n6596 , new_n6593 , new_n6595 );
  xor      g06220 ( new_n6597 , new_n6590 , new_n6596 );
  xor      g06221 ( new_n6598 , new_n6589 , new_n6597 );
  xnor     g06222 ( new_n6599 , new_n6586 , new_n6598 );
  nand     g06223 ( new_n6600 , new_n4832 , new_n4835 );
  nand     g06224 ( new_n6601 , new_n4831 , new_n4836 );
  nand     g06225 ( new_n6602 , new_n6600 , new_n6601 );
  xor      g06226 ( new_n6603 , new_n6599 , new_n6602 );
  nor      g06227 ( new_n6604 , new_n4822 , new_n4825 );
  and      g06228 ( new_n6605 , new_n4826 , new_n4837 );
  or       g06229 ( new_n6606 , new_n6604 , new_n6605 );
  xnor     g06230 ( new_n6607 , new_n6603 , new_n6606 );
  xor      g06231 ( new_n6608 , new_n6580 , new_n6607 );
  xnor     g06232 ( new_n6609 , new_n6579 , new_n6608 );
  xnor     g06233 ( new_n6610 , new_n6578 , new_n6609 );
  xnor     g06234 ( new_n6611 , new_n6545 , new_n6610 );
  xnor     g06235 ( new_n6612 , new_n6541 , new_n6611 );
  nand     g06236 ( new_n6613 , new_n4739 , new_n4905 );
  nand     g06237 ( new_n6614 , new_n4906 , new_n4927 );
  nand     g06238 ( new_n6615 , new_n6613 , new_n6614 );
  nand     g06239 ( new_n6616 , new_n4730 , new_n4738 );
  nand     g06240 ( new_n6617 , pi036 , pi131 );
  xor      g06241 ( new_n6618 , new_n6616 , new_n6617 );
  nor      g06242 ( new_n6619 , new_n4716 , new_n4727 );
  nor      g06243 ( new_n6620 , new_n4715 , new_n4729 );
  nor      g06244 ( new_n6621 , new_n6619 , new_n6620 );
  nand     g06245 ( new_n6622 , pi077 , pi085 );
  nand     g06246 ( new_n6623 , pi052 , pi180 );
  nand     g06247 ( new_n6624 , new_n6622 , new_n6623 );
  nand     g06248 ( new_n6625 , pi077 , pi180 );
  nor      g06249 ( new_n6626 , new_n4722 , new_n6625 );
  nand g06250 ( new_n6627 , new_n6626 , new_n6626 );
  nand     g06251 ( new_n6628 , new_n6624 , new_n6627 );
  nand     g06252 ( new_n6629 , new_n4718 , new_n4719 );
  nand     g06253 ( new_n6630 , new_n4717 , new_n4720 );
  nand     g06254 ( new_n6631 , new_n6629 , new_n6630 );
  nand     g06255 ( new_n6632 , pi133 , pi194 );
  nand     g06256 ( new_n6633 , pi064 , pi143 );
  nand     g06257 ( new_n6634 , pi057 , pi189 );
  nand     g06258 ( new_n6635 , new_n6633 , new_n6634 );
  nand     g06259 ( new_n6636 , pi057 , pi064 );
  nor      g06260 ( new_n6637 , new_n4718 , new_n6636 );
  nand g06261 ( new_n6638 , new_n6637 , new_n6637 );
  nand     g06262 ( new_n6639 , new_n6635 , new_n6638 );
  xor      g06263 ( new_n6640 , new_n6632 , new_n6639 );
  xor      g06264 ( new_n6641 , new_n6631 , new_n6640 );
  xor      g06265 ( new_n6642 , new_n6628 , new_n6641 );
  nand     g06266 ( new_n6643 , new_n4722 , new_n4725 );
  nand     g06267 ( new_n6644 , new_n4721 , new_n4726 );
  nand     g06268 ( new_n6645 , new_n6643 , new_n6644 );
  xor      g06269 ( new_n6646 , new_n6642 , new_n6645 );
  xor      g06270 ( new_n6647 , new_n6621 , new_n6646 );
  xor      g06271 ( new_n6648 , new_n6618 , new_n6647 );
  xor      g06272 ( new_n6649 , new_n6615 , new_n6648 );
  xnor     g06273 ( po028 , new_n6612 , new_n6649 );
  xnor     g06274 ( po029 , new_n899 , new_n900 );
  xor      g06275 ( po030 , new_n1880 , new_n1881 );
  nand     g06276 ( new_n6653 , pi103 , pi217 );
  nand g06277 ( new_n6654 , new_n6653 , new_n6653 );
  and      g06278 ( new_n6655 , pi175 , pi249 );
  nand     g06279 ( new_n6656 , pi107 , pi242 );
  nand     g06280 ( new_n6657 , pi163 , pi210 );
  xor      g06281 ( new_n6658 , new_n6656 , new_n6657 );
  xor      g06282 ( new_n6659 , new_n6655 , new_n6658 );
  xor      g06283 ( po031 , new_n6654 , new_n6659 );
  xnor     g06284 ( po032 , new_n2573 , new_n2593 );
  or       g06285 ( new_n6662 , new_n6656 , new_n6657 );
  nand     g06286 ( new_n6663 , pi111 , pi148 );
  or       g06287 ( new_n6664 , new_n6657 , new_n6663 );
  nand     g06288 ( new_n6665 , pi148 , pi210 );
  nand     g06289 ( new_n6666 , pi111 , pi163 );
  nand     g06290 ( new_n6667 , new_n6665 , new_n6666 );
  nand     g06291 ( new_n6668 , new_n6664 , new_n6667 );
  nor      g06292 ( new_n6669 , new_n6662 , new_n6668 );
  xnor     g06293 ( new_n6670 , new_n6662 , new_n6668 );
  nand     g06294 ( new_n6671 , pi140 , pi171 );
  nor      g06295 ( new_n6672 , new_n6656 , new_n6671 );
  nand     g06296 ( new_n6673 , pi107 , pi140 );
  nand     g06297 ( new_n6674 , pi171 , pi242 );
  and      g06298 ( new_n6675 , new_n6673 , new_n6674 );
  or       g06299 ( new_n6676 , new_n6672 , new_n6675 );
  nor      g06300 ( new_n6677 , new_n6670 , new_n6676 );
  nor      g06301 ( new_n6678 , new_n6669 , new_n6677 );
  nand     g06302 ( new_n6679 , pi049 , pi242 );
  nand     g06303 ( new_n6680 , pi107 , pi252 );
  xor      g06304 ( new_n6681 , new_n6671 , new_n6680 );
  xnor     g06305 ( new_n6682 , new_n6679 , new_n6681 );
  xnor     g06306 ( new_n6683 , new_n6672 , new_n6682 );
  nand     g06307 ( new_n6684 , pi210 , pi228 );
  nand     g06308 ( new_n6685 , pi024 , pi163 );
  nand     g06309 ( new_n6686 , new_n6684 , new_n6685 );
  or       g06310 ( new_n6687 , new_n6684 , new_n6685 );
  and      g06311 ( new_n6688 , new_n6686 , new_n6687 );
  nand g06312 ( new_n6689 , new_n6657 , new_n6657 );
  nor      g06313 ( new_n6690 , new_n6689 , new_n6663 );
  or       g06314 ( new_n6691 , new_n6688 , new_n6690 );
  nand     g06315 ( new_n6692 , new_n6686 , new_n6690 );
  nand     g06316 ( new_n6693 , new_n6691 , new_n6692 );
  xnor     g06317 ( new_n6694 , new_n6683 , new_n6693 );
  xor      g06318 ( new_n6695 , new_n6678 , new_n6694 );
  nand     g06319 ( new_n6696 , new_n6655 , new_n6658 );
  nand     g06320 ( new_n6697 , pi134 , pi249 );
  nand     g06321 ( new_n6698 , pi175 , pi222 );
  xnor     g06322 ( new_n6699 , new_n6697 , new_n6698 );
  and      g06323 ( new_n6700 , new_n6696 , new_n6699 );
  xor      g06324 ( new_n6701 , new_n6670 , new_n6676 );
  xnor     g06325 ( new_n6702 , new_n6696 , new_n6699 );
  nor      g06326 ( new_n6703 , new_n6701 , new_n6702 );
  nor      g06327 ( new_n6704 , new_n6700 , new_n6703 );
  nand     g06328 ( new_n6705 , pi134 , pi222 );
  nor      g06329 ( new_n6706 , new_n6655 , new_n6705 );
  nand     g06330 ( new_n6707 , pi240 , pi249 );
  nand     g06331 ( new_n6708 , pi125 , pi175 );
  or       g06332 ( new_n6709 , new_n6707 , new_n6708 );
  nand     g06333 ( new_n6710 , new_n6707 , new_n6708 );
  and      g06334 ( new_n6711 , new_n6709 , new_n6710 );
  or       g06335 ( new_n6712 , new_n6706 , new_n6711 );
  nand     g06336 ( new_n6713 , new_n6710 , new_n6706 );
  nand     g06337 ( new_n6714 , new_n6712 , new_n6713 );
  xor      g06338 ( new_n6715 , new_n6704 , new_n6714 );
  xnor     g06339 ( new_n6716 , new_n6695 , new_n6715 );
  nand     g06340 ( new_n6717 , new_n6654 , new_n6659 );
  nand     g06341 ( new_n6718 , pi100 , pi117 );
  nand g06342 ( new_n6719 , new_n6718 , new_n6718 );
  nand     g06343 ( new_n6720 , new_n6654 , new_n6719 );
  nand     g06344 ( new_n6721 , pi100 , pi103 );
  nand     g06345 ( new_n6722 , pi117 , pi217 );
  nand     g06346 ( new_n6723 , new_n6721 , new_n6722 );
  nand     g06347 ( new_n6724 , new_n6720 , new_n6723 );
  or       g06348 ( new_n6725 , new_n6717 , new_n6724 );
  xor      g06349 ( new_n6726 , new_n6717 , new_n6724 );
  xnor     g06350 ( new_n6727 , new_n6701 , new_n6702 );
  nand     g06351 ( new_n6728 , new_n6726 , new_n6727 );
  and      g06352 ( new_n6729 , new_n6725 , new_n6728 );
  nand     g06353 ( new_n6730 , pi103 , pi227 );
  nand     g06354 ( new_n6731 , pi016 , pi217 );
  nor      g06355 ( new_n6732 , new_n6730 , new_n6731 );
  nand     g06356 ( new_n6733 , new_n6730 , new_n6731 );
  nor      g06357 ( new_n6734 , new_n6654 , new_n6718 );
  nor      g06358 ( new_n6735 , new_n6733 , new_n6734 );
  nor      g06359 ( new_n6736 , new_n6732 , new_n6735 );
  nand     g06360 ( new_n6737 , new_n6733 , new_n6734 );
  nand     g06361 ( new_n6738 , new_n6736 , new_n6737 );
  xnor     g06362 ( new_n6739 , new_n6729 , new_n6738 );
  xnor     g06363 ( po033 , new_n6716 , new_n6739 );
  xnor     g06364 ( po034 , new_n4409 , new_n4480 );
  xor      g06365 ( po035 , new_n4274 , new_n4283 );
  nand     g06366 ( new_n6743 , pi081 , pi117 );
  nand     g06367 ( new_n6744 , pi080 , pi217 );
  nand     g06368 ( new_n6745 , pi016 , pi100 );
  nand     g06369 ( new_n6746 , new_n6744 , new_n6745 );
  nand     g06370 ( new_n6747 , pi117 , pi227 );
  xor      g06371 ( new_n6748 , new_n6744 , new_n6745 );
  nand     g06372 ( new_n6749 , new_n6747 , new_n6748 );
  nand     g06373 ( new_n6750 , new_n6746 , new_n6749 );
  nand     g06374 ( new_n6751 , new_n6743 , new_n6750 );
  nand     g06375 ( new_n6752 , pi217 , pi247 );
  nand     g06376 ( new_n6753 , pi016 , pi227 );
  nand     g06377 ( new_n6754 , pi080 , pi100 );
  xor      g06378 ( new_n6755 , new_n6753 , new_n6754 );
  xor      g06379 ( new_n6756 , new_n6752 , new_n6755 );
  xor      g06380 ( new_n6757 , new_n6743 , new_n6750 );
  nand     g06381 ( new_n6758 , new_n6756 , new_n6757 );
  nand     g06382 ( new_n6759 , new_n6751 , new_n6758 );
  nand     g06383 ( new_n6760 , pi016 , pi106 );
  nor      g06384 ( new_n6761 , new_n6743 , new_n6760 );
  nand     g06385 ( new_n6762 , pi016 , pi081 );
  nand     g06386 ( new_n6763 , pi106 , pi117 );
  and      g06387 ( new_n6764 , new_n6762 , new_n6763 );
  nor      g06388 ( new_n6765 , new_n6761 , new_n6764 );
  nand     g06389 ( new_n6766 , new_n6753 , new_n6754 );
  nand     g06390 ( new_n6767 , new_n6752 , new_n6755 );
  nand     g06391 ( new_n6768 , new_n6766 , new_n6767 );
  nand     g06392 ( new_n6769 , pi080 , pi227 );
  nand     g06393 ( new_n6770 , pi100 , pi234 );
  nor      g06394 ( new_n6771 , new_n6752 , new_n6770 );
  nand g06395 ( new_n6772 , new_n6771 , new_n6771 );
  nand     g06396 ( new_n6773 , pi217 , pi234 );
  nand     g06397 ( new_n6774 , pi100 , pi247 );
  nand     g06398 ( new_n6775 , new_n6773 , new_n6774 );
  nand     g06399 ( new_n6776 , new_n6772 , new_n6775 );
  xor      g06400 ( new_n6777 , new_n6769 , new_n6776 );
  xor      g06401 ( new_n6778 , new_n6768 , new_n6777 );
  xor      g06402 ( new_n6779 , new_n6765 , new_n6778 );
  nor      g06403 ( new_n6780 , new_n6759 , new_n6779 );
  nand g06404 ( new_n6781 , new_n6780 , new_n6780 );
  nand g06405 ( new_n6782 , new_n6778 , new_n6778 );
  nand     g06406 ( new_n6783 , new_n6765 , new_n6782 );
  nand g06407 ( new_n6784 , new_n6783 , new_n6783 );
  nor      g06408 ( new_n6785 , new_n6761 , new_n6784 );
  nand     g06409 ( new_n6786 , new_n6781 , new_n6785 );
  nand     g06410 ( new_n6787 , pi214 , pi217 );
  nand     g06411 ( new_n6788 , pi227 , pi247 );
  xor      g06412 ( new_n6789 , new_n6787 , new_n6788 );
  xor      g06413 ( new_n6790 , new_n6770 , new_n6789 );
  nand     g06414 ( new_n6791 , pi080 , pi081 );
  xor      g06415 ( new_n6792 , new_n6771 , new_n6791 );
  xor      g06416 ( new_n6793 , new_n6790 , new_n6792 );
  nand     g06417 ( new_n6794 , new_n6769 , new_n6776 );
  nand     g06418 ( new_n6795 , new_n6768 , new_n6777 );
  nand     g06419 ( new_n6796 , new_n6794 , new_n6795 );
  nand     g06420 ( new_n6797 , pi117 , pi233 );
  nand     g06421 ( new_n6798 , pi103 , pi187 );
  xor      g06422 ( new_n6799 , new_n6797 , new_n6798 );
  xnor     g06423 ( new_n6800 , new_n6760 , new_n6799 );
  xor      g06424 ( new_n6801 , new_n6796 , new_n6800 );
  xor      g06425 ( new_n6802 , new_n6793 , new_n6801 );
  nand g06426 ( new_n6803 , new_n6802 , new_n6802 );
  nand     g06427 ( new_n6804 , new_n6761 , new_n6780 );
  nand     g06428 ( new_n6805 , new_n6786 , new_n6804 );
  or       g06429 ( new_n6806 , new_n6803 , new_n6805 );
  nand     g06430 ( new_n6807 , new_n6786 , new_n6806 );
  nand     g06431 ( new_n6808 , pi021 , pi171 );
  nand     g06432 ( new_n6809 , pi049 , pi231 );
  nand     g06433 ( new_n6810 , pi121 , pi171 );
  nor      g06434 ( new_n6811 , new_n6809 , new_n6810 );
  nand g06435 ( new_n6812 , new_n6811 , new_n6811 );
  nand     g06436 ( new_n6813 , pi171 , pi231 );
  nand     g06437 ( new_n6814 , pi049 , pi121 );
  nand     g06438 ( new_n6815 , new_n6813 , new_n6814 );
  nand     g06439 ( new_n6816 , new_n6812 , new_n6815 );
  nand     g06440 ( new_n6817 , pi140 , pi156 );
  nand     g06441 ( new_n6818 , pi201 , pi242 );
  nor      g06442 ( new_n6819 , new_n6817 , new_n6818 );
  nand g06443 ( new_n6820 , new_n6819 , new_n6819 );
  nand     g06444 ( new_n6821 , pi140 , pi201 );
  nand     g06445 ( new_n6822 , pi156 , pi242 );
  nand     g06446 ( new_n6823 , new_n6821 , new_n6822 );
  nand     g06447 ( new_n6824 , new_n6820 , new_n6823 );
  nand     g06448 ( new_n6825 , pi245 , pi252 );
  nand     g06449 ( new_n6826 , pi140 , pi245 );
  nand     g06450 ( new_n6827 , new_n6818 , new_n6826 );
  xor      g06451 ( new_n6828 , new_n6818 , new_n6826 );
  nand     g06452 ( new_n6829 , pi049 , pi252 );
  nand     g06453 ( new_n6830 , new_n6828 , new_n6829 );
  nand     g06454 ( new_n6831 , new_n6827 , new_n6830 );
  xor      g06455 ( new_n6832 , new_n6825 , new_n6831 );
  xor      g06456 ( new_n6833 , new_n6824 , new_n6832 );
  xor      g06457 ( new_n6834 , new_n6816 , new_n6833 );
  nand     g06458 ( new_n6835 , pi049 , pi140 );
  nand     g06459 ( new_n6836 , pi242 , pi245 );
  nand     g06460 ( new_n6837 , new_n6835 , new_n6836 );
  nand     g06461 ( new_n6838 , pi171 , pi252 );
  xor      g06462 ( new_n6839 , new_n6835 , new_n6836 );
  nand     g06463 ( new_n6840 , new_n6838 , new_n6839 );
  nand     g06464 ( new_n6841 , new_n6837 , new_n6840 );
  nand     g06465 ( new_n6842 , new_n6810 , new_n6841 );
  xor      g06466 ( new_n6843 , new_n6828 , new_n6829 );
  xor      g06467 ( new_n6844 , new_n6810 , new_n6841 );
  nand     g06468 ( new_n6845 , new_n6843 , new_n6844 );
  nand     g06469 ( new_n6846 , new_n6842 , new_n6845 );
  nand g06470 ( new_n6847 , new_n6846 , new_n6846 );
  nand     g06471 ( new_n6848 , new_n6834 , new_n6847 );
  nor      g06472 ( new_n6849 , new_n6816 , new_n6833 );
  nor      g06473 ( new_n6850 , new_n6811 , new_n6849 );
  nand     g06474 ( new_n6851 , new_n6848 , new_n6850 );
  nand     g06475 ( new_n6852 , pi063 , pi242 );
  nand     g06476 ( new_n6853 , pi201 , pi252 );
  xor      g06477 ( new_n6854 , new_n6852 , new_n6853 );
  xor      g06478 ( new_n6855 , new_n6817 , new_n6854 );
  nand     g06479 ( new_n6856 , pi121 , pi245 );
  xor      g06480 ( new_n6857 , new_n6819 , new_n6856 );
  xnor     g06481 ( new_n6858 , new_n6855 , new_n6857 );
  nand     g06482 ( new_n6859 , new_n6825 , new_n6831 );
  nand     g06483 ( new_n6860 , new_n6824 , new_n6832 );
  nand     g06484 ( new_n6861 , new_n6859 , new_n6860 );
  nand     g06485 ( new_n6862 , pi021 , pi107 );
  nand     g06486 ( new_n6863 , pi005 , pi171 );
  xor      g06487 ( new_n6864 , new_n6862 , new_n6863 );
  xor      g06488 ( new_n6865 , new_n6809 , new_n6864 );
  xnor     g06489 ( new_n6866 , new_n6861 , new_n6865 );
  xor      g06490 ( new_n6867 , new_n6858 , new_n6866 );
  or       g06491 ( new_n6868 , new_n6812 , new_n6848 );
  nand     g06492 ( new_n6869 , new_n6851 , new_n6868 );
  or       g06493 ( new_n6870 , new_n6867 , new_n6869 );
  nand     g06494 ( new_n6871 , new_n6851 , new_n6870 );
  xor      g06495 ( new_n6872 , new_n6808 , new_n6871 );
  nand     g06496 ( new_n6873 , pi163 , pi232 );
  nand     g06497 ( new_n6874 , pi127 , pi148 );
  nand     g06498 ( new_n6875 , new_n6873 , new_n6874 );
  nand     g06499 ( new_n6876 , pi228 , pi255 );
  xor      g06500 ( new_n6877 , new_n6873 , new_n6874 );
  nand     g06501 ( new_n6878 , new_n6876 , new_n6877 );
  nand     g06502 ( new_n6879 , new_n6875 , new_n6878 );
  nand     g06503 ( new_n6880 , new_n6709 , new_n6705 );
  nand     g06504 ( new_n6881 , new_n6710 , new_n6880 );
  nand     g06505 ( new_n6882 , pi175 , pi176 );
  nor      g06506 ( new_n6883 , new_n6881 , new_n6882 );
  xor      g06507 ( new_n6884 , new_n6881 , new_n6882 );
  nand g06508 ( new_n6885 , new_n6884 , new_n6884 );
  nand     g06509 ( new_n6886 , pi149 , pi249 );
  nand     g06510 ( new_n6887 , pi125 , pi134 );
  nand     g06511 ( new_n6888 , pi222 , pi240 );
  xor      g06512 ( new_n6889 , new_n6887 , new_n6888 );
  xor      g06513 ( new_n6890 , new_n6886 , new_n6889 );
  nor      g06514 ( new_n6891 , new_n6885 , new_n6890 );
  nor      g06515 ( new_n6892 , new_n6883 , new_n6891 );
  nand     g06516 ( new_n6893 , pi040 , pi175 );
  nand     g06517 ( new_n6894 , pi167 , pi249 );
  nand     g06518 ( new_n6895 , pi125 , pi240 );
  nand     g06519 ( new_n6896 , pi149 , pi222 );
  xor      g06520 ( new_n6897 , new_n6895 , new_n6896 );
  xor      g06521 ( new_n6898 , new_n6894 , new_n6897 );
  nand     g06522 ( new_n6899 , pi134 , pi176 );
  nand     g06523 ( new_n6900 , new_n6887 , new_n6888 );
  nand     g06524 ( new_n6901 , new_n6886 , new_n6889 );
  nand     g06525 ( new_n6902 , new_n6900 , new_n6901 );
  xor      g06526 ( new_n6903 , new_n6899 , new_n6902 );
  xor      g06527 ( new_n6904 , new_n6898 , new_n6903 );
  xor      g06528 ( new_n6905 , new_n6893 , new_n6904 );
  nand g06529 ( new_n6906 , new_n6905 , new_n6905 );
  xor      g06530 ( new_n6907 , new_n6892 , new_n6906 );
  nor      g06531 ( new_n6908 , new_n6705 , new_n6712 );
  xor      g06532 ( new_n6909 , new_n6884 , new_n6890 );
  nand g06533 ( new_n6910 , new_n6909 , new_n6909 );
  nand     g06534 ( new_n6911 , new_n6908 , new_n6910 );
  nand g06535 ( new_n6912 , new_n6911 , new_n6911 );
  nand     g06536 ( new_n6913 , new_n6907 , new_n6912 );
  nand     g06537 ( new_n6914 , pi174 , pi175 );
  nand     g06538 ( new_n6915 , new_n6913 , new_n6914 );
  xor      g06539 ( new_n6916 , new_n6913 , new_n6914 );
  nand g06540 ( new_n6917 , new_n6916 , new_n6916 );
  nand     g06541 ( new_n6918 , new_n6899 , new_n6902 );
  nand     g06542 ( new_n6919 , new_n6898 , new_n6903 );
  nand     g06543 ( new_n6920 , new_n6918 , new_n6919 );
  nand     g06544 ( new_n6921 , pi176 , pi240 );
  nand     g06545 ( new_n6922 , pi040 , pi134 );
  and      g06546 ( new_n6923 , new_n6921 , new_n6922 );
  nand     g06547 ( new_n6924 , pi040 , pi240 );
  nor      g06548 ( new_n6925 , new_n6899 , new_n6924 );
  or       g06549 ( new_n6926 , new_n6923 , new_n6925 );
  xor      g06550 ( new_n6927 , new_n6920 , new_n6926 );
  nand     g06551 ( new_n6928 , new_n6895 , new_n6896 );
  nand     g06552 ( new_n6929 , new_n6894 , new_n6897 );
  nand     g06553 ( new_n6930 , new_n6928 , new_n6929 );
  nand     g06554 ( new_n6931 , pi125 , pi149 );
  nand     g06555 ( new_n6932 , pi167 , pi222 );
  nand     g06556 ( new_n6933 , pi181 , pi249 );
  nand     g06557 ( new_n6934 , new_n6932 , new_n6933 );
  nand     g06558 ( new_n6935 , pi181 , pi222 );
  nor      g06559 ( new_n6936 , new_n6894 , new_n6935 );
  nand g06560 ( new_n6937 , new_n6936 , new_n6936 );
  nand     g06561 ( new_n6938 , new_n6934 , new_n6937 );
  xor      g06562 ( new_n6939 , new_n6931 , new_n6938 );
  xor      g06563 ( new_n6940 , new_n6930 , new_n6939 );
  xor      g06564 ( new_n6941 , new_n6927 , new_n6940 );
  nor      g06565 ( new_n6942 , new_n6893 , new_n6904 );
  nor      g06566 ( new_n6943 , new_n6892 , new_n6906 );
  nor      g06567 ( new_n6944 , new_n6942 , new_n6943 );
  xor      g06568 ( new_n6945 , new_n6941 , new_n6944 );
  or       g06569 ( new_n6946 , new_n6917 , new_n6945 );
  nand     g06570 ( new_n6947 , new_n6915 , new_n6946 );
  nor      g06571 ( new_n6948 , new_n6941 , new_n6944 );
  nand     g06572 ( new_n6949 , new_n6920 , new_n6926 );
  nand     g06573 ( new_n6950 , new_n6927 , new_n6940 );
  nand     g06574 ( new_n6951 , new_n6949 , new_n6950 );
  xor      g06575 ( new_n6952 , new_n6925 , new_n6951 );
  nand g06576 ( new_n6953 , new_n6952 , new_n6952 );
  nand     g06577 ( new_n6954 , pi149 , pi176 );
  xor      g06578 ( new_n6955 , new_n6936 , new_n6954 );
  nand     g06579 ( new_n6956 , pi200 , pi249 );
  nand     g06580 ( new_n6957 , pi125 , pi167 );
  xor      g06581 ( new_n6958 , new_n6956 , new_n6957 );
  xor      g06582 ( new_n6959 , new_n6935 , new_n6958 );
  xor      g06583 ( new_n6960 , new_n6955 , new_n6959 );
  nand     g06584 ( new_n6961 , new_n6931 , new_n6938 );
  nand     g06585 ( new_n6962 , new_n6930 , new_n6939 );
  nand     g06586 ( new_n6963 , new_n6961 , new_n6962 );
  nand     g06587 ( new_n6964 , pi157 , pi175 );
  nand     g06588 ( new_n6965 , pi134 , pi174 );
  xor      g06589 ( new_n6966 , new_n6964 , new_n6965 );
  xor      g06590 ( new_n6967 , new_n6924 , new_n6966 );
  xnor     g06591 ( new_n6968 , new_n6963 , new_n6967 );
  xor      g06592 ( new_n6969 , new_n6960 , new_n6968 );
  xor      g06593 ( new_n6970 , new_n6953 , new_n6969 );
  xor      g06594 ( new_n6971 , new_n6948 , new_n6970 );
  xnor     g06595 ( new_n6972 , new_n6947 , new_n6971 );
  nand     g06596 ( new_n6973 , pi107 , pi231 );
  nand     g06597 ( new_n6974 , pi107 , pi121 );
  nand     g06598 ( new_n6975 , new_n6671 , new_n6680 );
  nand     g06599 ( new_n6976 , new_n6679 , new_n6681 );
  nand     g06600 ( new_n6977 , new_n6975 , new_n6976 );
  nor      g06601 ( new_n6978 , new_n6974 , new_n6977 );
  xor      g06602 ( new_n6979 , new_n6838 , new_n6839 );
  xnor     g06603 ( new_n6980 , new_n6974 , new_n6977 );
  nor      g06604 ( new_n6981 , new_n6979 , new_n6980 );
  nor      g06605 ( new_n6982 , new_n6978 , new_n6981 );
  nor      g06606 ( new_n6983 , new_n6973 , new_n6982 );
  xor      g06607 ( new_n6984 , new_n6973 , new_n6982 );
  xor      g06608 ( new_n6985 , new_n6843 , new_n6844 );
  nand g06609 ( new_n6986 , new_n6985 , new_n6985 );
  and      g06610 ( new_n6987 , new_n6984 , new_n6986 );
  nor      g06611 ( new_n6988 , new_n6983 , new_n6987 );
  xor      g06612 ( new_n6989 , new_n6834 , new_n6846 );
  xor      g06613 ( new_n6990 , new_n6988 , new_n6989 );
  and      g06614 ( new_n6991 , pi005 , pi107 );
  and      g06615 ( new_n6992 , new_n6990 , new_n6991 );
  xor      g06616 ( new_n6993 , new_n6984 , new_n6986 );
  nand     g06617 ( new_n6994 , new_n6672 , new_n6682 );
  xnor     g06618 ( new_n6995 , new_n6979 , new_n6980 );
  nor      g06619 ( new_n6996 , new_n6994 , new_n6995 );
  and      g06620 ( new_n6997 , new_n6993 , new_n6996 );
  nand g06621 ( new_n6998 , new_n6997 , new_n6997 );
  xnor     g06622 ( new_n6999 , new_n6990 , new_n6991 );
  nor      g06623 ( new_n7000 , new_n6998 , new_n6999 );
  nor      g06624 ( new_n7001 , new_n6992 , new_n7000 );
  nor      g06625 ( new_n7002 , new_n6988 , new_n6989 );
  xor      g06626 ( new_n7003 , new_n6867 , new_n6869 );
  xor      g06627 ( new_n7004 , new_n7002 , new_n7003 );
  xor      g06628 ( new_n7005 , new_n7001 , new_n7004 );
  nand     g06629 ( new_n7006 , pi163 , pi255 );
  nand     g06630 ( new_n7007 , new_n6663 , new_n6687 );
  nand     g06631 ( new_n7008 , new_n6686 , new_n7007 );
  nand     g06632 ( new_n7009 , pi163 , pi224 );
  nand     g06633 ( new_n7010 , new_n7008 , new_n7009 );
  nand     g06634 ( new_n7011 , pi039 , pi210 );
  nand     g06635 ( new_n7012 , pi111 , pi228 );
  nand     g06636 ( new_n7013 , pi024 , pi148 );
  xor      g06637 ( new_n7014 , new_n7012 , new_n7013 );
  xor      g06638 ( new_n7015 , new_n7011 , new_n7014 );
  xor      g06639 ( new_n7016 , new_n7008 , new_n7009 );
  nand     g06640 ( new_n7017 , new_n7015 , new_n7016 );
  nand     g06641 ( new_n7018 , new_n7010 , new_n7017 );
  nor      g06642 ( new_n7019 , new_n7006 , new_n7018 );
  xor      g06643 ( new_n7020 , new_n7006 , new_n7018 );
  nand     g06644 ( new_n7021 , pi116 , pi210 );
  nand     g06645 ( new_n7022 , pi024 , pi228 );
  nand     g06646 ( new_n7023 , pi039 , pi111 );
  xor      g06647 ( new_n7024 , new_n7022 , new_n7023 );
  xor      g06648 ( new_n7025 , new_n7021 , new_n7024 );
  nand     g06649 ( new_n7026 , pi148 , pi224 );
  nand     g06650 ( new_n7027 , new_n7012 , new_n7013 );
  nand     g06651 ( new_n7028 , new_n7011 , new_n7014 );
  nand     g06652 ( new_n7029 , new_n7027 , new_n7028 );
  xnor     g06653 ( new_n7030 , new_n7026 , new_n7029 );
  xor      g06654 ( new_n7031 , new_n7025 , new_n7030 );
  and      g06655 ( new_n7032 , new_n7020 , new_n7031 );
  nor      g06656 ( new_n7033 , new_n7019 , new_n7032 );
  nand     g06657 ( new_n7034 , pi024 , pi039 );
  nand     g06658 ( new_n7035 , pi111 , pi116 );
  nand     g06659 ( new_n7036 , pi070 , pi210 );
  nand     g06660 ( new_n7037 , new_n7035 , new_n7036 );
  nand     g06661 ( new_n7038 , pi070 , pi111 );
  or       g06662 ( new_n7039 , new_n7021 , new_n7038 );
  nand     g06663 ( new_n7040 , new_n7037 , new_n7039 );
  xor      g06664 ( new_n7041 , new_n7034 , new_n7040 );
  nand     g06665 ( new_n7042 , new_n7022 , new_n7023 );
  nand     g06666 ( new_n7043 , new_n7021 , new_n7024 );
  nand     g06667 ( new_n7044 , new_n7042 , new_n7043 );
  xor      g06668 ( new_n7045 , new_n7041 , new_n7044 );
  nand     g06669 ( new_n7046 , pi224 , pi228 );
  nand     g06670 ( new_n7047 , pi148 , pi255 );
  and      g06671 ( new_n7048 , new_n7046 , new_n7047 );
  nor      g06672 ( new_n7049 , new_n6876 , new_n7026 );
  or       g06673 ( new_n7050 , new_n7048 , new_n7049 );
  xor      g06674 ( new_n7051 , new_n7045 , new_n7050 );
  nand     g06675 ( new_n7052 , new_n7026 , new_n7029 );
  nand g06676 ( new_n7053 , new_n7025 , new_n7025 );
  or       g06677 ( new_n7054 , new_n7053 , new_n7030 );
  nand     g06678 ( new_n7055 , new_n7052 , new_n7054 );
  xor      g06679 ( new_n7056 , new_n7051 , new_n7055 );
  xnor     g06680 ( new_n7057 , new_n7033 , new_n7056 );
  nand     g06681 ( new_n7058 , pi127 , pi163 );
  nor      g06682 ( new_n7059 , new_n7057 , new_n7058 );
  xor      g06683 ( new_n7060 , new_n7020 , new_n7031 );
  nor      g06684 ( new_n7061 , new_n6664 , new_n6688 );
  xnor     g06685 ( new_n7062 , new_n7015 , new_n7016 );
  and      g06686 ( new_n7063 , new_n7061 , new_n7062 );
  nand     g06687 ( new_n7064 , new_n7060 , new_n7063 );
  xnor     g06688 ( new_n7065 , new_n7057 , new_n7058 );
  nor      g06689 ( new_n7066 , new_n7064 , new_n7065 );
  nor      g06690 ( new_n7067 , new_n7059 , new_n7066 );
  or       g06691 ( new_n7068 , new_n7033 , new_n7056 );
  nand g06692 ( new_n7069 , new_n7051 , new_n7051 );
  nor      g06693 ( new_n7070 , new_n7069 , new_n7055 );
  and      g06694 ( new_n7071 , new_n7049 , new_n7070 );
  nor      g06695 ( new_n7072 , new_n7045 , new_n7050 );
  nor      g06696 ( new_n7073 , new_n7049 , new_n7072 );
  nand g06697 ( new_n7074 , new_n7073 , new_n7073 );
  nor      g06698 ( new_n7075 , new_n7070 , new_n7074 );
  or       g06699 ( new_n7076 , new_n7071 , new_n7075 );
  nand     g06700 ( new_n7077 , pi039 , pi224 );
  xnor     g06701 ( new_n7078 , new_n7039 , new_n7077 );
  nand     g06702 ( new_n7079 , pi115 , pi210 );
  nand     g06703 ( new_n7080 , pi024 , pi116 );
  xor      g06704 ( new_n7081 , new_n7079 , new_n7080 );
  xor      g06705 ( new_n7082 , new_n7038 , new_n7081 );
  xnor     g06706 ( new_n7083 , new_n7078 , new_n7082 );
  nand     g06707 ( new_n7084 , new_n7034 , new_n7040 );
  nand     g06708 ( new_n7085 , new_n7041 , new_n7044 );
  nand     g06709 ( new_n7086 , new_n7084 , new_n7085 );
  xor      g06710 ( new_n7087 , new_n6876 , new_n6877 );
  xnor     g06711 ( new_n7088 , new_n7086 , new_n7087 );
  xor      g06712 ( new_n7089 , new_n7083 , new_n7088 );
  xor      g06713 ( new_n7090 , new_n7076 , new_n7089 );
  xnor     g06714 ( new_n7091 , new_n7068 , new_n7090 );
  xor      g06715 ( new_n7092 , new_n7067 , new_n7091 );
  xor      g06716 ( new_n7093 , new_n7005 , new_n7092 );
  xnor     g06717 ( new_n7094 , new_n7064 , new_n7065 );
  xor      g06718 ( new_n7095 , new_n6997 , new_n6999 );
  nand     g06719 ( new_n7096 , new_n7094 , new_n7095 );
  or       g06720 ( new_n7097 , new_n7094 , new_n7095 );
  xor      g06721 ( new_n7098 , new_n7060 , new_n7063 );
  nor      g06722 ( new_n7099 , new_n6683 , new_n6693 );
  nor      g06723 ( new_n7100 , new_n6678 , new_n6694 );
  or       g06724 ( new_n7101 , new_n7099 , new_n7100 );
  xor      g06725 ( new_n7102 , new_n6994 , new_n6995 );
  nor      g06726 ( new_n7103 , new_n7101 , new_n7102 );
  xor      g06727 ( new_n7104 , new_n7061 , new_n7062 );
  xnor     g06728 ( new_n7105 , new_n7101 , new_n7102 );
  nor      g06729 ( new_n7106 , new_n7104 , new_n7105 );
  nor      g06730 ( new_n7107 , new_n7103 , new_n7106 );
  or       g06731 ( new_n7108 , new_n7098 , new_n7107 );
  xnor     g06732 ( new_n7109 , new_n6993 , new_n6996 );
  xor      g06733 ( new_n7110 , new_n7098 , new_n7107 );
  nand     g06734 ( new_n7111 , new_n7109 , new_n7110 );
  nand     g06735 ( new_n7112 , new_n7108 , new_n7111 );
  nand     g06736 ( new_n7113 , new_n7097 , new_n7112 );
  nand     g06737 ( new_n7114 , new_n7096 , new_n7113 );
  xor      g06738 ( new_n7115 , new_n7093 , new_n7114 );
  nor      g06739 ( new_n7116 , new_n6972 , new_n7115 );
  xor      g06740 ( new_n7117 , new_n6972 , new_n7115 );
  xor      g06741 ( new_n7118 , new_n6916 , new_n6945 );
  nand g06742 ( new_n7119 , new_n7118 , new_n7118 );
  xor      g06743 ( new_n7120 , new_n7094 , new_n7095 );
  xor      g06744 ( new_n7121 , new_n7112 , new_n7120 );
  nor      g06745 ( new_n7122 , new_n7119 , new_n7121 );
  xor      g06746 ( new_n7123 , new_n6907 , new_n6912 );
  xnor     g06747 ( new_n7124 , new_n7109 , new_n7110 );
  or       g06748 ( new_n7125 , new_n7123 , new_n7124 );
  xor      g06749 ( new_n7126 , new_n7123 , new_n7124 );
  xor      g06750 ( new_n7127 , new_n6908 , new_n6909 );
  nand g06751 ( new_n7128 , new_n7127 , new_n7127 );
  nand g06752 ( new_n7129 , new_n6714 , new_n6714 );
  nor      g06753 ( new_n7130 , new_n6704 , new_n7129 );
  nor      g06754 ( new_n7131 , new_n6695 , new_n6715 );
  nor      g06755 ( new_n7132 , new_n7130 , new_n7131 );
  nand     g06756 ( new_n7133 , new_n7128 , new_n7132 );
  xor      g06757 ( new_n7134 , new_n7128 , new_n7132 );
  xnor     g06758 ( new_n7135 , new_n7104 , new_n7105 );
  nand     g06759 ( new_n7136 , new_n7134 , new_n7135 );
  and      g06760 ( new_n7137 , new_n7133 , new_n7136 );
  nand     g06761 ( new_n7138 , new_n7126 , new_n7137 );
  nand     g06762 ( new_n7139 , new_n7125 , new_n7138 );
  xor      g06763 ( new_n7140 , new_n7118 , new_n7121 );
  nor      g06764 ( new_n7141 , new_n7139 , new_n7140 );
  or       g06765 ( new_n7142 , new_n7122 , new_n7141 );
  and      g06766 ( new_n7143 , new_n7117 , new_n7142 );
  nor      g06767 ( new_n7144 , new_n7116 , new_n7143 );
  nand     g06768 ( new_n7145 , new_n6852 , new_n6853 );
  nand     g06769 ( new_n7146 , new_n6817 , new_n6854 );
  nand     g06770 ( new_n7147 , new_n7145 , new_n7146 );
  xor      g06771 ( new_n7148 , new_n7144 , new_n7147 );
  xor      g06772 ( new_n7149 , new_n6879 , new_n7148 );
  nand     g06773 ( new_n7150 , pi039 , pi255 );
  nand     g06774 ( new_n7151 , pi156 , pi252 );
  xor      g06775 ( new_n7152 , new_n7150 , new_n7151 );
  nor      g06776 ( new_n7153 , new_n7039 , new_n7077 );
  nor      g06777 ( new_n7154 , new_n7078 , new_n7082 );
  nor      g06778 ( new_n7155 , new_n7153 , new_n7154 );
  xor      g06779 ( new_n7156 , new_n7152 , new_n7155 );
  xor      g06780 ( new_n7157 , new_n7149 , new_n7156 );
  xnor     g06781 ( new_n7158 , new_n6872 , new_n7157 );
  xor      g06782 ( new_n7159 , new_n6807 , new_n7158 );
  nand     g06783 ( new_n7160 , pi080 , pi106 );
  nand     g06784 ( new_n7161 , pi116 , pi224 );
  xor      g06785 ( new_n7162 , new_n7139 , new_n7140 );
  nand     g06786 ( new_n7163 , pi081 , pi103 );
  or       g06787 ( new_n7164 , new_n6719 , new_n6732 );
  nand     g06788 ( new_n7165 , new_n6733 , new_n7164 );
  nor      g06789 ( new_n7166 , new_n7163 , new_n7165 );
  xor      g06790 ( new_n7167 , new_n6747 , new_n6748 );
  xor      g06791 ( new_n7168 , new_n7163 , new_n7165 );
  nand g06792 ( new_n7169 , new_n7168 , new_n7168 );
  nor      g06793 ( new_n7170 , new_n7167 , new_n7169 );
  nor      g06794 ( new_n7171 , new_n7166 , new_n7170 );
  nand     g06795 ( new_n7172 , pi103 , pi106 );
  xor      g06796 ( new_n7173 , new_n6756 , new_n6757 );
  xnor     g06797 ( new_n7174 , new_n7172 , new_n7173 );
  xor      g06798 ( new_n7175 , new_n7171 , new_n7174 );
  nor      g06799 ( new_n7176 , new_n6720 , new_n6736 );
  nand g06800 ( new_n7177 , new_n7176 , new_n7176 );
  xor      g06801 ( new_n7178 , new_n7167 , new_n7168 );
  nor      g06802 ( new_n7179 , new_n7177 , new_n7178 );
  nand     g06803 ( new_n7180 , new_n7175 , new_n7179 );
  nand     g06804 ( new_n7181 , pi103 , pi233 );
  xor      g06805 ( new_n7182 , new_n7180 , new_n7181 );
  xor      g06806 ( new_n7183 , new_n6759 , new_n6779 );
  nor      g06807 ( new_n7184 , new_n7172 , new_n7173 );
  nor      g06808 ( new_n7185 , new_n7171 , new_n7174 );
  nor      g06809 ( new_n7186 , new_n7184 , new_n7185 );
  xor      g06810 ( new_n7187 , new_n7183 , new_n7186 );
  xnor     g06811 ( new_n7188 , new_n7182 , new_n7187 );
  and      g06812 ( new_n7189 , new_n7162 , new_n7188 );
  and      g06813 ( new_n7190 , new_n6729 , new_n6738 );
  nor      g06814 ( new_n7191 , new_n6716 , new_n6739 );
  nor      g06815 ( new_n7192 , new_n7190 , new_n7191 );
  xor      g06816 ( new_n7193 , new_n7177 , new_n7178 );
  or       g06817 ( new_n7194 , new_n7192 , new_n7193 );
  xnor     g06818 ( new_n7195 , new_n7134 , new_n7135 );
  xor      g06819 ( new_n7196 , new_n7192 , new_n7193 );
  nand     g06820 ( new_n7197 , new_n7195 , new_n7196 );
  nand     g06821 ( new_n7198 , new_n7194 , new_n7197 );
  xor      g06822 ( new_n7199 , new_n7175 , new_n7179 );
  nand g06823 ( new_n7200 , new_n7199 , new_n7199 );
  nor      g06824 ( new_n7201 , new_n7198 , new_n7200 );
  xor      g06825 ( new_n7202 , new_n7126 , new_n7137 );
  xor      g06826 ( new_n7203 , new_n7198 , new_n7199 );
  nor      g06827 ( new_n7204 , new_n7202 , new_n7203 );
  nor      g06828 ( new_n7205 , new_n7201 , new_n7204 );
  xnor     g06829 ( new_n7206 , new_n7162 , new_n7188 );
  nor      g06830 ( new_n7207 , new_n7205 , new_n7206 );
  nor      g06831 ( new_n7208 , new_n7189 , new_n7207 );
  nand     g06832 ( new_n7209 , new_n7180 , new_n7181 );
  nand     g06833 ( new_n7210 , new_n7182 , new_n7187 );
  nand     g06834 ( new_n7211 , new_n7209 , new_n7210 );
  nand g06835 ( new_n7212 , new_n7183 , new_n7183 );
  nor      g06836 ( new_n7213 , new_n7212 , new_n7186 );
  xor      g06837 ( new_n7214 , new_n6802 , new_n6805 );
  xor      g06838 ( new_n7215 , new_n7213 , new_n7214 );
  xor      g06839 ( new_n7216 , new_n7211 , new_n7215 );
  nand     g06840 ( new_n7217 , new_n7208 , new_n7216 );
  xor      g06841 ( new_n7218 , new_n7208 , new_n7216 );
  xnor     g06842 ( new_n7219 , new_n7117 , new_n7142 );
  nand     g06843 ( new_n7220 , new_n7218 , new_n7219 );
  nand     g06844 ( new_n7221 , new_n7217 , new_n7220 );
  xor      g06845 ( new_n7222 , new_n7161 , new_n7221 );
  xor      g06846 ( new_n7223 , new_n7160 , new_n7222 );
  nand     g06847 ( new_n7224 , new_n6787 , new_n6788 );
  nand     g06848 ( new_n7225 , new_n6770 , new_n6789 );
  nand     g06849 ( new_n7226 , new_n7224 , new_n7225 );
  nand     g06850 ( new_n7227 , pi203 , pi249 );
  nand     g06851 ( new_n7228 , pi081 , pi247 );
  xor      g06852 ( new_n7229 , new_n7227 , new_n7228 );
  nand g06853 ( new_n7230 , new_n6948 , new_n6948 );
  nor      g06854 ( new_n7231 , new_n7230 , new_n6970 );
  nor      g06855 ( new_n7232 , new_n6947 , new_n6971 );
  nor      g06856 ( new_n7233 , new_n7231 , new_n7232 );
  nand g06857 ( new_n7234 , new_n6951 , new_n6951 );
  nor      g06858 ( new_n7235 , new_n6925 , new_n7234 );
  and      g06859 ( new_n7236 , new_n6953 , new_n6969 );
  nor      g06860 ( new_n7237 , new_n7235 , new_n7236 );
  xor      g06861 ( new_n7238 , new_n7233 , new_n7237 );
  xor      g06862 ( new_n7239 , new_n7229 , new_n7238 );
  xor      g06863 ( new_n7240 , new_n7226 , new_n7239 );
  xor      g06864 ( new_n7241 , new_n7223 , new_n7240 );
  nand     g06865 ( new_n7242 , pi017 , pi175 );
  nand     g06866 ( new_n7243 , pi227 , pi234 );
  xor      g06867 ( new_n7244 , new_n7242 , new_n7243 );
  nand g06868 ( new_n7245 , new_n6796 , new_n6796 );
  nor      g06869 ( new_n7246 , new_n7245 , new_n6800 );
  nor      g06870 ( new_n7247 , new_n6793 , new_n6801 );
  nor      g06871 ( new_n7248 , new_n7246 , new_n7247 );
  nor      g06872 ( new_n7249 , new_n6861 , new_n6865 );
  nor      g06873 ( new_n7250 , new_n6858 , new_n6866 );
  nor      g06874 ( new_n7251 , new_n7249 , new_n7250 );
  xor      g06875 ( new_n7252 , new_n7248 , new_n7251 );
  nand     g06876 ( new_n7253 , pi231 , pi245 );
  nand     g06877 ( new_n7254 , pi082 , pi107 );
  xor      g06878 ( new_n7255 , new_n7253 , new_n7254 );
  xor      g06879 ( new_n7256 , new_n7252 , new_n7255 );
  nand     g06880 ( new_n7257 , new_n6862 , new_n6863 );
  nand     g06881 ( new_n7258 , new_n6809 , new_n6864 );
  nand     g06882 ( new_n7259 , new_n7257 , new_n7258 );
  nand     g06883 ( new_n7260 , new_n7079 , new_n7080 );
  nand     g06884 ( new_n7261 , new_n7038 , new_n7081 );
  nand     g06885 ( new_n7262 , new_n7260 , new_n7261 );
  xor      g06886 ( new_n7263 , new_n7259 , new_n7262 );
  xor      g06887 ( new_n7264 , new_n7256 , new_n7263 );
  xor      g06888 ( new_n7265 , new_n7244 , new_n7264 );
  xor      g06889 ( new_n7266 , new_n7241 , new_n7265 );
  nand     g06890 ( new_n7267 , pi040 , pi149 );
  nand     g06891 ( new_n7268 , pi100 , pi214 );
  xor      g06892 ( new_n7269 , new_n7267 , new_n7268 );
  nand     g06893 ( new_n7270 , pi005 , pi049 );
  nand     g06894 ( new_n7271 , pi111 , pi115 );
  xor      g06895 ( new_n7272 , new_n7270 , new_n7271 );
  nand     g06896 ( new_n7273 , pi083 , pi242 );
  nand     g06897 ( new_n7274 , new_n6797 , new_n6798 );
  nand     g06898 ( new_n7275 , new_n6760 , new_n6799 );
  nand     g06899 ( new_n7276 , new_n7274 , new_n7275 );
  xor      g06900 ( new_n7277 , new_n7273 , new_n7276 );
  nand     g06901 ( new_n7278 , pi016 , pi233 );
  nor      g06902 ( new_n7279 , new_n6963 , new_n6967 );
  nand g06903 ( new_n7280 , new_n6960 , new_n6960 );
  nor      g06904 ( new_n7281 , new_n7280 , new_n6968 );
  nor      g06905 ( new_n7282 , new_n7279 , new_n7281 );
  xor      g06906 ( new_n7283 , new_n7278 , new_n7282 );
  xor      g06907 ( new_n7284 , new_n7277 , new_n7283 );
  xor      g06908 ( new_n7285 , new_n7272 , new_n7284 );
  xor      g06909 ( new_n7286 , new_n7269 , new_n7285 );
  nand     g06910 ( new_n7287 , pi127 , pi228 );
  or       g06911 ( new_n7288 , new_n7005 , new_n7092 );
  nand     g06912 ( new_n7289 , new_n7093 , new_n7114 );
  nand     g06913 ( new_n7290 , new_n7288 , new_n7289 );
  xor      g06914 ( new_n7291 , new_n7287 , new_n7290 );
  nor      g06915 ( new_n7292 , new_n6772 , new_n6791 );
  nor      g06916 ( new_n7293 , new_n6790 , new_n6792 );
  nor      g06917 ( new_n7294 , new_n7292 , new_n7293 );
  nand     g06918 ( new_n7295 , pi125 , pi181 );
  xor      g06919 ( new_n7296 , new_n7294 , new_n7295 );
  nor      g06920 ( new_n7297 , new_n7068 , new_n7090 );
  nor      g06921 ( new_n7298 , new_n7067 , new_n7091 );
  nor      g06922 ( new_n7299 , new_n7297 , new_n7298 );
  xor      g06923 ( new_n7300 , new_n7296 , new_n7299 );
  nor      g06924 ( new_n7301 , new_n6820 , new_n6856 );
  nor      g06925 ( new_n7302 , new_n6855 , new_n6857 );
  nor      g06926 ( new_n7303 , new_n7301 , new_n7302 );
  nand     g06927 ( new_n7304 , new_n7213 , new_n7214 );
  nand g06928 ( new_n7305 , new_n7211 , new_n7211 );
  nand     g06929 ( new_n7306 , new_n7305 , new_n7215 );
  nand     g06930 ( new_n7307 , new_n7304 , new_n7306 );
  nor      g06931 ( new_n7308 , new_n7076 , new_n7089 );
  nor      g06932 ( new_n7309 , new_n7075 , new_n7308 );
  xor      g06933 ( new_n7310 , new_n7307 , new_n7309 );
  xor      g06934 ( new_n7311 , new_n7303 , new_n7310 );
  xor      g06935 ( new_n7312 , new_n7300 , new_n7311 );
  xor      g06936 ( new_n7313 , new_n7291 , new_n7312 );
  nor      g06937 ( new_n7314 , new_n6937 , new_n6954 );
  nor      g06938 ( new_n7315 , new_n6955 , new_n6959 );
  nor      g06939 ( new_n7316 , new_n7314 , new_n7315 );
  nand     g06940 ( new_n7317 , pi202 , pi217 );
  xor      g06941 ( new_n7318 , new_n7316 , new_n7317 );
  nand     g06942 ( new_n7319 , pi163 , pi191 );
  nand     g06943 ( new_n7320 , new_n6964 , new_n6965 );
  nand     g06944 ( new_n7321 , new_n6924 , new_n6966 );
  nand     g06945 ( new_n7322 , new_n7320 , new_n7321 );
  xor      g06946 ( new_n7323 , new_n7319 , new_n7322 );
  nand     g06947 ( new_n7324 , pi000 , pi210 );
  xor      g06948 ( new_n7325 , new_n7323 , new_n7324 );
  xor      g06949 ( new_n7326 , new_n7318 , new_n7325 );
  nand g06950 ( new_n7327 , new_n7002 , new_n7002 );
  nor      g06951 ( new_n7328 , new_n7327 , new_n7003 );
  nor      g06952 ( new_n7329 , new_n7001 , new_n7004 );
  nor      g06953 ( new_n7330 , new_n7328 , new_n7329 );
  nand     g06954 ( new_n7331 , pi103 , pi129 );
  xor      g06955 ( new_n7332 , new_n7330 , new_n7331 );
  nand     g06956 ( new_n7333 , pi167 , pi176 );
  nand     g06957 ( new_n7334 , pi200 , pi222 );
  nor      g06958 ( new_n7335 , new_n7086 , new_n7087 );
  nor      g06959 ( new_n7336 , new_n7083 , new_n7088 );
  nor      g06960 ( new_n7337 , new_n7335 , new_n7336 );
  nand     g06961 ( new_n7338 , pi134 , pi157 );
  xor      g06962 ( new_n7339 , new_n7337 , new_n7338 );
  xor      g06963 ( new_n7340 , new_n7334 , new_n7339 );
  xor      g06964 ( new_n7341 , new_n7333 , new_n7340 );
  xor      g06965 ( new_n7342 , new_n7332 , new_n7341 );
  nand     g06966 ( new_n7343 , new_n6956 , new_n6957 );
  nand     g06967 ( new_n7344 , new_n6935 , new_n6958 );
  nand     g06968 ( new_n7345 , new_n7343 , new_n7344 );
  nand     g06969 ( new_n7346 , pi063 , pi140 );
  xor      g06970 ( new_n7347 , new_n7345 , new_n7346 );
  nand     g06971 ( new_n7348 , pi117 , pi187 );
  nand     g06972 ( new_n7349 , pi174 , pi240 );
  xor      g06973 ( new_n7350 , new_n7348 , new_n7349 );
  xor      g06974 ( new_n7351 , new_n7347 , new_n7350 );
  xor      g06975 ( new_n7352 , new_n7342 , new_n7351 );
  xor      g06976 ( new_n7353 , new_n7326 , new_n7352 );
  xor      g06977 ( new_n7354 , new_n7313 , new_n7353 );
  xor      g06978 ( new_n7355 , new_n7286 , new_n7354 );
  nand     g06979 ( new_n7356 , pi024 , pi070 );
  nand     g06980 ( new_n7357 , pi148 , pi232 );
  nand     g06981 ( new_n7358 , pi121 , pi201 );
  xor      g06982 ( new_n7359 , new_n7357 , new_n7358 );
  xor      g06983 ( new_n7360 , new_n7356 , new_n7359 );
  xor      g06984 ( new_n7361 , new_n7355 , new_n7360 );
  xor      g06985 ( new_n7362 , new_n7266 , new_n7361 );
  xor      g06986 ( po036 , new_n7159 , new_n7362 );
  xor      g06987 ( po037 , new_n7205 , new_n7206 );
  xor      g06988 ( po038 , new_n3252 , new_n3253 );
  nand     g06989 ( new_n7366 , pi044 , pi052 );
  nand     g06990 ( new_n7367 , pi119 , pi133 );
  nand     g06991 ( new_n7368 , pi045 , pi077 );
  nand     g06992 ( new_n7369 , new_n7367 , new_n7368 );
  nand     g06993 ( new_n7370 , pi052 , pi250 );
  xor      g06994 ( new_n7371 , new_n7367 , new_n7368 );
  nand     g06995 ( new_n7372 , new_n7370 , new_n7371 );
  nand     g06996 ( new_n7373 , new_n7369 , new_n7372 );
  nand     g06997 ( new_n7374 , new_n7366 , new_n7373 );
  nand     g06998 ( new_n7375 , pi045 , pi133 );
  nand     g06999 ( new_n7376 , pi119 , pi189 );
  nand g07000 ( new_n7377 , new_n7376 , new_n7376 );
  nand     g07001 ( new_n7378 , pi077 , pi250 );
  xor      g07002 ( new_n7379 , new_n7377 , new_n7378 );
  xor      g07003 ( new_n7380 , new_n7375 , new_n7379 );
  nand g07004 ( new_n7381 , new_n7380 , new_n7380 );
  xor      g07005 ( new_n7382 , new_n7366 , new_n7373 );
  nand     g07006 ( new_n7383 , new_n7381 , new_n7382 );
  nand     g07007 ( new_n7384 , new_n7374 , new_n7383 );
  nand     g07008 ( new_n7385 , pi044 , pi077 );
  nand     g07009 ( new_n7386 , pi052 , pi054 );
  and      g07010 ( new_n7387 , new_n7385 , new_n7386 );
  nand     g07011 ( new_n7388 , pi054 , pi077 );
  nor      g07012 ( new_n7389 , new_n7366 , new_n7388 );
  nor      g07013 ( new_n7390 , new_n7387 , new_n7389 );
  nand     g07014 ( new_n7391 , new_n7376 , new_n7378 );
  nand g07015 ( new_n7392 , new_n7379 , new_n7379 );
  nand     g07016 ( new_n7393 , new_n7375 , new_n7392 );
  nand     g07017 ( new_n7394 , new_n7391 , new_n7393 );
  nand     g07018 ( new_n7395 , pi133 , pi250 );
  nand     g07019 ( new_n7396 , pi045 , pi064 );
  nand g07020 ( new_n7397 , new_n7396 , new_n7396 );
  nand     g07021 ( new_n7398 , new_n7377 , new_n7397 );
  nand     g07022 ( new_n7399 , pi045 , pi189 );
  nand     g07023 ( new_n7400 , pi064 , pi119 );
  nand     g07024 ( new_n7401 , new_n7399 , new_n7400 );
  nand     g07025 ( new_n7402 , new_n7398 , new_n7401 );
  xor      g07026 ( new_n7403 , new_n7395 , new_n7402 );
  xor      g07027 ( new_n7404 , new_n7394 , new_n7403 );
  xor      g07028 ( new_n7405 , new_n7390 , new_n7404 );
  xor      g07029 ( new_n7406 , new_n7384 , new_n7405 );
  nand     g07030 ( new_n7407 , pi054 , pi131 );
  nand     g07031 ( new_n7408 , pi044 , pi131 );
  nand     g07032 ( new_n7409 , pi131 , pi250 );
  nand     g07033 ( new_n7410 , pi045 , pi052 );
  nand     g07034 ( new_n7411 , new_n7409 , new_n7410 );
  nand     g07035 ( new_n7412 , pi077 , pi119 );
  xor      g07036 ( new_n7413 , new_n7409 , new_n7410 );
  nand     g07037 ( new_n7414 , new_n7412 , new_n7413 );
  nand     g07038 ( new_n7415 , new_n7411 , new_n7414 );
  nand     g07039 ( new_n7416 , new_n7408 , new_n7415 );
  xor      g07040 ( new_n7417 , new_n7370 , new_n7371 );
  xor      g07041 ( new_n7418 , new_n7408 , new_n7415 );
  nand     g07042 ( new_n7419 , new_n7417 , new_n7418 );
  nand     g07043 ( new_n7420 , new_n7416 , new_n7419 );
  nor      g07044 ( new_n7421 , new_n7407 , new_n7420 );
  xor      g07045 ( new_n7422 , new_n7407 , new_n7420 );
  xor      g07046 ( new_n7423 , new_n7380 , new_n7382 );
  nand     g07047 ( new_n7424 , new_n7422 , new_n7423 );
  nand g07048 ( new_n7425 , new_n7424 , new_n7424 );
  nor      g07049 ( new_n7426 , new_n7421 , new_n7425 );
  xor      g07050 ( new_n7427 , new_n7406 , new_n7426 );
  nand g07051 ( new_n7428 , new_n7427 , new_n7427 );
  nand     g07052 ( new_n7429 , pi072 , pi131 );
  xor      g07053 ( new_n7430 , new_n7417 , new_n7418 );
  nand g07054 ( new_n7431 , new_n7430 , new_n7430 );
  xor      g07055 ( new_n7432 , new_n7412 , new_n7413 );
  nand g07056 ( new_n7433 , new_n7432 , new_n7432 );
  nand     g07057 ( new_n7434 , pi045 , pi131 );
  nand     g07058 ( new_n7435 , pi052 , pi119 );
  nor      g07059 ( new_n7436 , new_n7434 , new_n7435 );
  nand     g07060 ( new_n7437 , new_n7433 , new_n7436 );
  nand g07061 ( new_n7438 , new_n7437 , new_n7437 );
  nand     g07062 ( new_n7439 , new_n7431 , new_n7438 );
  nand g07063 ( new_n7440 , new_n7439 , new_n7439 );
  xor      g07064 ( new_n7441 , new_n7422 , new_n7423 );
  nand     g07065 ( new_n7442 , new_n7440 , new_n7441 );
  xnor     g07066 ( new_n7443 , new_n7429 , new_n7442 );
  xor      g07067 ( new_n7444 , new_n7428 , new_n7443 );
  nand     g07068 ( new_n7445 , pi151 , pi208 );
  nand     g07069 ( new_n7446 , pi019 , pi168 );
  nand     g07070 ( new_n7447 , pi139 , pi147 );
  or       g07071 ( new_n7448 , new_n7446 , new_n7447 );
  nand g07072 ( new_n7449 , new_n7445 , new_n7445 );
  nand     g07073 ( new_n7450 , new_n378 , new_n7449 );
  nand g07074 ( new_n7451 , new_n7450 , new_n7450 );
  nand     g07075 ( new_n7452 , new_n7446 , new_n7447 );
  or       g07076 ( new_n7453 , new_n7451 , new_n7452 );
  nand     g07077 ( new_n7454 , new_n7448 , new_n7453 );
  nand g07078 ( new_n7455 , new_n7454 , new_n7454 );
  nor      g07079 ( new_n7456 , new_n7445 , new_n7455 );
  nand     g07080 ( new_n7457 , new_n7445 , new_n7448 );
  nand     g07081 ( new_n7458 , new_n7452 , new_n7457 );
  nand     g07082 ( new_n7459 , pi097 , pi168 );
  xor      g07083 ( new_n7460 , new_n7458 , new_n7459 );
  nand     g07084 ( new_n7461 , pi035 , pi147 );
  nand     g07085 ( new_n7462 , pi019 , pi208 );
  nand     g07086 ( new_n7463 , pi139 , pi151 );
  xor      g07087 ( new_n7464 , new_n7462 , new_n7463 );
  xor      g07088 ( new_n7465 , new_n7461 , new_n7464 );
  xor      g07089 ( new_n7466 , new_n7460 , new_n7465 );
  nand g07090 ( new_n7467 , new_n7466 , new_n7466 );
  xor      g07091 ( new_n7468 , new_n7456 , new_n7467 );
  nand     g07092 ( new_n7469 , pi104 , pi164 );
  nand     g07093 ( new_n7470 , pi206 , pi212 );
  nand     g07094 ( new_n7471 , pi032 , pi213 );
  xor      g07095 ( new_n7472 , new_n7470 , new_n7471 );
  xor      g07096 ( new_n7473 , new_n7469 , new_n7472 );
  nor      g07097 ( new_n7474 , new_n379 , new_n7470 );
  xor      g07098 ( new_n7475 , new_n7473 , new_n7474 );
  nand     g07099 ( new_n7476 , pi027 , pi161 );
  nand     g07100 ( new_n7477 , pi008 , pi236 );
  nor      g07101 ( new_n7478 , new_n7476 , new_n7477 );
  nand     g07102 ( new_n7479 , new_n7476 , new_n7477 );
  nand     g07103 ( new_n7480 , pi026 , pi241 );
  nor      g07104 ( new_n7481 , new_n381 , new_n7480 );
  nor      g07105 ( new_n7482 , new_n7479 , new_n7481 );
  nor      g07106 ( new_n7483 , new_n7478 , new_n7482 );
  nand     g07107 ( new_n7484 , new_n7479 , new_n7481 );
  nand     g07108 ( new_n7485 , new_n7483 , new_n7484 );
  or       g07109 ( new_n7486 , new_n7475 , new_n7485 );
  nor      g07110 ( new_n7487 , new_n379 , new_n380 );
  nand     g07111 ( new_n7488 , pi027 , pi241 );
  nand     g07112 ( new_n7489 , pi026 , pi236 );
  xor      g07113 ( new_n7490 , new_n7488 , new_n7489 );
  nand     g07114 ( new_n7491 , new_n7487 , new_n7490 );
  nand     g07115 ( new_n7492 , pi206 , pi213 );
  nand     g07116 ( new_n7493 , pi164 , pi212 );
  and      g07117 ( new_n7494 , new_n7492 , new_n7493 );
  nor      g07118 ( new_n7495 , new_n7474 , new_n7494 );
  xor      g07119 ( new_n7496 , new_n7487 , new_n7490 );
  nand     g07120 ( new_n7497 , new_n7495 , new_n7496 );
  nand     g07121 ( new_n7498 , new_n7491 , new_n7497 );
  xor      g07122 ( new_n7499 , new_n7475 , new_n7485 );
  nand     g07123 ( new_n7500 , new_n7498 , new_n7499 );
  nand     g07124 ( new_n7501 , new_n7486 , new_n7500 );
  nor      g07125 ( new_n7502 , new_n7480 , new_n7483 );
  nand     g07126 ( new_n7503 , pi026 , pi161 );
  nand     g07127 ( new_n7504 , pi008 , pi241 );
  nand     g07128 ( new_n7505 , pi027 , pi141 );
  xnor     g07129 ( new_n7506 , new_n7504 , new_n7505 );
  nand g07130 ( new_n7507 , new_n7506 , new_n7506 );
  xor      g07131 ( new_n7508 , new_n7503 , new_n7507 );
  nand g07132 ( new_n7509 , new_n7479 , new_n7479 );
  nand g07133 ( new_n7510 , new_n7480 , new_n7480 );
  nor      g07134 ( new_n7511 , new_n7510 , new_n7478 );
  nor      g07135 ( new_n7512 , new_n7509 , new_n7511 );
  nand     g07136 ( new_n7513 , pi056 , pi236 );
  xor      g07137 ( new_n7514 , new_n7512 , new_n7513 );
  xor      g07138 ( new_n7515 , new_n7508 , new_n7514 );
  xor      g07139 ( new_n7516 , new_n7502 , new_n7515 );
  xnor     g07140 ( new_n7517 , new_n7501 , new_n7516 );
  nand g07141 ( new_n7518 , new_n7473 , new_n7473 );
  nand     g07142 ( new_n7519 , new_n7518 , new_n7474 );
  nand     g07143 ( new_n7520 , pi145 , pi213 );
  nand     g07144 ( new_n7521 , new_n7470 , new_n7471 );
  nand     g07145 ( new_n7522 , new_n7469 , new_n7472 );
  nand     g07146 ( new_n7523 , new_n7521 , new_n7522 );
  xor      g07147 ( new_n7524 , new_n7520 , new_n7523 );
  nand     g07148 ( new_n7525 , pi032 , pi212 );
  nand     g07149 ( new_n7526 , pi104 , pi206 );
  nand     g07150 ( new_n7527 , pi013 , pi164 );
  xor      g07151 ( new_n7528 , new_n7526 , new_n7527 );
  xor      g07152 ( new_n7529 , new_n7525 , new_n7528 );
  xor      g07153 ( new_n7530 , new_n7524 , new_n7529 );
  xor      g07154 ( new_n7531 , new_n7519 , new_n7530 );
  xnor     g07155 ( new_n7532 , new_n7517 , new_n7531 );
  nor      g07156 ( new_n7533 , new_n7468 , new_n7532 );
  xnor     g07157 ( new_n7534 , new_n7468 , new_n7532 );
  xor      g07158 ( new_n7535 , new_n7498 , new_n7499 );
  nand     g07159 ( new_n7536 , new_n7451 , new_n7452 );
  nand     g07160 ( new_n7537 , new_n7455 , new_n7536 );
  nand g07161 ( new_n7538 , new_n7537 , new_n7537 );
  nor      g07162 ( new_n7539 , new_n7535 , new_n7538 );
  nor      g07163 ( new_n7540 , new_n378 , new_n382 );
  nand     g07164 ( new_n7541 , pi151 , pi168 );
  nand     g07165 ( new_n7542 , pi147 , pi208 );
  xor      g07166 ( new_n7543 , new_n7541 , new_n7542 );
  nor      g07167 ( new_n7544 , new_n7540 , new_n7543 );
  xor      g07168 ( new_n7545 , new_n7540 , new_n7543 );
  xnor     g07169 ( new_n7546 , new_n7495 , new_n7496 );
  and      g07170 ( new_n7547 , new_n7545 , new_n7546 );
  nor      g07171 ( new_n7548 , new_n7544 , new_n7547 );
  xor      g07172 ( new_n7549 , new_n7535 , new_n7537 );
  nor      g07173 ( new_n7550 , new_n7548 , new_n7549 );
  nor      g07174 ( new_n7551 , new_n7539 , new_n7550 );
  nor      g07175 ( new_n7552 , new_n7534 , new_n7551 );
  or       g07176 ( new_n7553 , new_n7533 , new_n7552 );
  nor      g07177 ( new_n7554 , new_n7501 , new_n7516 );
  nor      g07178 ( new_n7555 , new_n7517 , new_n7531 );
  nor      g07179 ( new_n7556 , new_n7554 , new_n7555 );
  nand     g07180 ( new_n7557 , new_n7502 , new_n7515 );
  nand g07181 ( new_n7558 , new_n7512 , new_n7512 );
  nor      g07182 ( new_n7559 , new_n7558 , new_n7513 );
  nor      g07183 ( new_n7560 , new_n7508 , new_n7514 );
  nor      g07184 ( new_n7561 , new_n7559 , new_n7560 );
  nand     g07185 ( new_n7562 , pi136 , pi236 );
  nand     g07186 ( new_n7563 , pi008 , pi161 );
  nand     g07187 ( new_n7564 , pi027 , pi090 );
  nand     g07188 ( new_n7565 , pi026 , pi141 );
  xor      g07189 ( new_n7566 , new_n7564 , new_n7565 );
  xor      g07190 ( new_n7567 , new_n7563 , new_n7566 );
  nand g07191 ( new_n7568 , new_n7567 , new_n7567 );
  nand     g07192 ( new_n7569 , new_n7504 , new_n7505 );
  nand     g07193 ( new_n7570 , new_n7503 , new_n7507 );
  nand     g07194 ( new_n7571 , new_n7569 , new_n7570 );
  nand     g07195 ( new_n7572 , pi056 , pi241 );
  xnor     g07196 ( new_n7573 , new_n7571 , new_n7572 );
  xor      g07197 ( new_n7574 , new_n7568 , new_n7573 );
  xnor     g07198 ( new_n7575 , new_n7562 , new_n7574 );
  xnor     g07199 ( new_n7576 , new_n7561 , new_n7575 );
  xor      g07200 ( new_n7577 , new_n7557 , new_n7576 );
  xnor     g07201 ( new_n7578 , new_n7556 , new_n7577 );
  nor      g07202 ( new_n7579 , new_n7519 , new_n7530 );
  nand     g07203 ( new_n7580 , pi145 , pi212 );
  nand     g07204 ( new_n7581 , new_n7526 , new_n7527 );
  nand     g07205 ( new_n7582 , new_n7525 , new_n7528 );
  nand     g07206 ( new_n7583 , new_n7581 , new_n7582 );
  xor      g07207 ( new_n7584 , new_n7580 , new_n7583 );
  nand     g07208 ( new_n7585 , pi112 , pi164 );
  nand     g07209 ( new_n7586 , pi013 , pi206 );
  nand     g07210 ( new_n7587 , pi032 , pi104 );
  xor      g07211 ( new_n7588 , new_n7586 , new_n7587 );
  xor      g07212 ( new_n7589 , new_n7585 , new_n7588 );
  xor      g07213 ( new_n7590 , new_n7584 , new_n7589 );
  nand     g07214 ( new_n7591 , pi213 , pi246 );
  xnor     g07215 ( new_n7592 , new_n7590 , new_n7591 );
  nand     g07216 ( new_n7593 , new_n7520 , new_n7523 );
  nand     g07217 ( new_n7594 , new_n7524 , new_n7529 );
  nand     g07218 ( new_n7595 , new_n7593 , new_n7594 );
  xor      g07219 ( new_n7596 , new_n7592 , new_n7595 );
  xor      g07220 ( new_n7597 , new_n7579 , new_n7596 );
  xor      g07221 ( new_n7598 , new_n7578 , new_n7597 );
  nand     g07222 ( new_n7599 , new_n7456 , new_n7467 );
  nand     g07223 ( new_n7600 , pi075 , pi168 );
  nor      g07224 ( new_n7601 , new_n7458 , new_n7459 );
  nand g07225 ( new_n7602 , new_n7460 , new_n7460 );
  nor      g07226 ( new_n7603 , new_n7602 , new_n7465 );
  nor      g07227 ( new_n7604 , new_n7601 , new_n7603 );
  xor      g07228 ( new_n7605 , new_n7600 , new_n7604 );
  nand     g07229 ( new_n7606 , pi019 , pi139 );
  nand     g07230 ( new_n7607 , pi015 , pi147 );
  nand     g07231 ( new_n7608 , pi035 , pi151 );
  xor      g07232 ( new_n7609 , new_n7607 , new_n7608 );
  xor      g07233 ( new_n7610 , new_n7606 , new_n7609 );
  nand     g07234 ( new_n7611 , pi097 , pi208 );
  nand     g07235 ( new_n7612 , new_n7462 , new_n7463 );
  nand     g07236 ( new_n7613 , new_n7461 , new_n7464 );
  nand     g07237 ( new_n7614 , new_n7612 , new_n7613 );
  xor      g07238 ( new_n7615 , new_n7611 , new_n7614 );
  xnor     g07239 ( new_n7616 , new_n7610 , new_n7615 );
  xor      g07240 ( new_n7617 , new_n7605 , new_n7616 );
  xor      g07241 ( new_n7618 , new_n7599 , new_n7617 );
  xor      g07242 ( new_n7619 , new_n7598 , new_n7618 );
  xor      g07243 ( new_n7620 , new_n7553 , new_n7619 );
  xor      g07244 ( new_n7621 , new_n7439 , new_n7441 );
  nor      g07245 ( new_n7622 , new_n7620 , new_n7621 );
  xor      g07246 ( new_n7623 , new_n7534 , new_n7551 );
  xor      g07247 ( new_n7624 , new_n7430 , new_n7438 );
  nor      g07248 ( new_n7625 , new_n7623 , new_n7624 );
  nor      g07249 ( new_n7626 , new_n377 , new_n384 );
  xor      g07250 ( new_n7627 , new_n7434 , new_n7435 );
  or       g07251 ( new_n7628 , new_n7626 , new_n7627 );
  xor      g07252 ( new_n7629 , new_n7545 , new_n7546 );
  xor      g07253 ( new_n7630 , new_n7626 , new_n7627 );
  nand     g07254 ( new_n7631 , new_n7629 , new_n7630 );
  nand     g07255 ( new_n7632 , new_n7628 , new_n7631 );
  xor      g07256 ( new_n7633 , new_n7548 , new_n7549 );
  nand     g07257 ( new_n7634 , new_n7632 , new_n7633 );
  xor      g07258 ( new_n7635 , new_n7433 , new_n7436 );
  nand g07259 ( new_n7636 , new_n7635 , new_n7635 );
  xor      g07260 ( new_n7637 , new_n7632 , new_n7633 );
  nand     g07261 ( new_n7638 , new_n7636 , new_n7637 );
  nand     g07262 ( new_n7639 , new_n7634 , new_n7638 );
  xnor     g07263 ( new_n7640 , new_n7623 , new_n7624 );
  nor      g07264 ( new_n7641 , new_n7639 , new_n7640 );
  nor      g07265 ( new_n7642 , new_n7625 , new_n7641 );
  xnor     g07266 ( new_n7643 , new_n7620 , new_n7621 );
  nor      g07267 ( new_n7644 , new_n7642 , new_n7643 );
  nor      g07268 ( new_n7645 , new_n7622 , new_n7644 );
  nor      g07269 ( new_n7646 , new_n7444 , new_n7645 );
  nand     g07270 ( new_n7647 , new_n7598 , new_n7618 );
  nand     g07271 ( new_n7648 , new_n7553 , new_n7619 );
  and      g07272 ( new_n7649 , new_n7647 , new_n7648 );
  nand g07273 ( new_n7650 , new_n7617 , new_n7617 );
  nor      g07274 ( new_n7651 , new_n7599 , new_n7650 );
  nand g07275 ( new_n7652 , new_n7651 , new_n7651 );
  nand     g07276 ( new_n7653 , pi093 , pi168 );
  xor      g07277 ( new_n7654 , new_n7652 , new_n7653 );
  nand     g07278 ( new_n7655 , pi075 , pi139 );
  nor      g07279 ( new_n7656 , new_n7611 , new_n7655 );
  nand     g07280 ( new_n7657 , pi097 , pi139 );
  nand     g07281 ( new_n7658 , pi075 , pi208 );
  and      g07282 ( new_n7659 , new_n7657 , new_n7658 );
  or       g07283 ( new_n7660 , new_n7656 , new_n7659 );
  nand     g07284 ( new_n7661 , pi015 , pi151 );
  nand     g07285 ( new_n7662 , pi147 , pi204 );
  nand     g07286 ( new_n7663 , new_n7661 , new_n7662 );
  nand     g07287 ( new_n7664 , pi151 , pi204 );
  nor      g07288 ( new_n7665 , new_n7607 , new_n7664 );
  nand g07289 ( new_n7666 , new_n7665 , new_n7665 );
  nand     g07290 ( new_n7667 , new_n7663 , new_n7666 );
  nand     g07291 ( new_n7668 , pi019 , pi035 );
  nand     g07292 ( new_n7669 , new_n7607 , new_n7608 );
  nand     g07293 ( new_n7670 , new_n7606 , new_n7609 );
  nand     g07294 ( new_n7671 , new_n7669 , new_n7670 );
  xor      g07295 ( new_n7672 , new_n7668 , new_n7671 );
  xor      g07296 ( new_n7673 , new_n7667 , new_n7672 );
  xor      g07297 ( new_n7674 , new_n7660 , new_n7673 );
  nand     g07298 ( new_n7675 , new_n7611 , new_n7614 );
  nand     g07299 ( new_n7676 , new_n7610 , new_n7615 );
  nand     g07300 ( new_n7677 , new_n7675 , new_n7676 );
  xor      g07301 ( new_n7678 , new_n7674 , new_n7677 );
  nor      g07302 ( new_n7679 , new_n7600 , new_n7604 );
  nand     g07303 ( new_n7680 , new_n7605 , new_n7616 );
  nand g07304 ( new_n7681 , new_n7680 , new_n7680 );
  nor      g07305 ( new_n7682 , new_n7679 , new_n7681 );
  xor      g07306 ( new_n7683 , new_n7678 , new_n7682 );
  xor      g07307 ( new_n7684 , new_n7654 , new_n7683 );
  nor      g07308 ( new_n7685 , new_n7556 , new_n7577 );
  nor      g07309 ( new_n7686 , new_n7578 , new_n7597 );
  nor      g07310 ( new_n7687 , new_n7685 , new_n7686 );
  nor      g07311 ( new_n7688 , new_n7590 , new_n7591 );
  nor      g07312 ( new_n7689 , new_n7592 , new_n7595 );
  nor      g07313 ( new_n7690 , new_n7688 , new_n7689 );
  nand     g07314 ( new_n7691 , pi104 , pi246 );
  nor      g07315 ( new_n7692 , new_n7580 , new_n7691 );
  nand     g07316 ( new_n7693 , pi104 , pi145 );
  nand     g07317 ( new_n7694 , pi212 , pi246 );
  and      g07318 ( new_n7695 , new_n7693 , new_n7694 );
  or       g07319 ( new_n7696 , new_n7692 , new_n7695 );
  nand     g07320 ( new_n7697 , new_n7586 , new_n7587 );
  nand     g07321 ( new_n7698 , new_n7585 , new_n7588 );
  nand     g07322 ( new_n7699 , new_n7697 , new_n7698 );
  nand     g07323 ( new_n7700 , pi112 , pi206 );
  nand     g07324 ( new_n7701 , pi105 , pi164 );
  nand     g07325 ( new_n7702 , new_n7700 , new_n7701 );
  nand     g07326 ( new_n7703 , pi105 , pi206 );
  nor      g07327 ( new_n7704 , new_n7585 , new_n7703 );
  nand g07328 ( new_n7705 , new_n7704 , new_n7704 );
  nand     g07329 ( new_n7706 , new_n7702 , new_n7705 );
  nand     g07330 ( new_n7707 , pi013 , pi032 );
  xor      g07331 ( new_n7708 , new_n7706 , new_n7707 );
  xor      g07332 ( new_n7709 , new_n7699 , new_n7708 );
  xor      g07333 ( new_n7710 , new_n7696 , new_n7709 );
  nand     g07334 ( new_n7711 , new_n7580 , new_n7583 );
  nand     g07335 ( new_n7712 , new_n7584 , new_n7589 );
  nand     g07336 ( new_n7713 , new_n7711 , new_n7712 );
  xor      g07337 ( new_n7714 , new_n7710 , new_n7713 );
  xnor     g07338 ( new_n7715 , new_n7690 , new_n7714 );
  nand     g07339 ( new_n7716 , new_n7579 , new_n7596 );
  nand     g07340 ( new_n7717 , pi114 , pi213 );
  xor      g07341 ( new_n7718 , new_n7716 , new_n7717 );
  xnor     g07342 ( new_n7719 , new_n7715 , new_n7718 );
  or       g07343 ( new_n7720 , new_n7557 , new_n7576 );
  nand     g07344 ( new_n7721 , pi096 , pi236 );
  xor      g07345 ( new_n7722 , new_n7720 , new_n7721 );
  nand     g07346 ( new_n7723 , new_n7571 , new_n7572 );
  or       g07347 ( new_n7724 , new_n7568 , new_n7573 );
  nand     g07348 ( new_n7725 , new_n7723 , new_n7724 );
  nand     g07349 ( new_n7726 , pi136 , pi241 );
  nand     g07350 ( new_n7727 , pi056 , pi161 );
  nand     g07351 ( new_n7728 , new_n7726 , new_n7727 );
  nand     g07352 ( new_n7729 , pi136 , pi161 );
  nor      g07353 ( new_n7730 , new_n7572 , new_n7729 );
  nand g07354 ( new_n7731 , new_n7730 , new_n7730 );
  nand     g07355 ( new_n7732 , new_n7728 , new_n7731 );
  nand     g07356 ( new_n7733 , new_n7564 , new_n7565 );
  nand     g07357 ( new_n7734 , new_n7563 , new_n7566 );
  nand     g07358 ( new_n7735 , new_n7733 , new_n7734 );
  nand     g07359 ( new_n7736 , pi008 , pi141 );
  nand     g07360 ( new_n7737 , pi026 , pi090 );
  nand     g07361 ( new_n7738 , pi027 , pi047 );
  nand     g07362 ( new_n7739 , new_n7737 , new_n7738 );
  nand     g07363 ( new_n7740 , pi026 , pi047 );
  nor      g07364 ( new_n7741 , new_n7564 , new_n7740 );
  nand g07365 ( new_n7742 , new_n7741 , new_n7741 );
  nand     g07366 ( new_n7743 , new_n7739 , new_n7742 );
  xor      g07367 ( new_n7744 , new_n7736 , new_n7743 );
  xor      g07368 ( new_n7745 , new_n7735 , new_n7744 );
  xnor     g07369 ( new_n7746 , new_n7732 , new_n7745 );
  xor      g07370 ( new_n7747 , new_n7725 , new_n7746 );
  nor      g07371 ( new_n7748 , new_n7562 , new_n7574 );
  nor      g07372 ( new_n7749 , new_n7561 , new_n7575 );
  nor      g07373 ( new_n7750 , new_n7748 , new_n7749 );
  xor      g07374 ( new_n7751 , new_n7747 , new_n7750 );
  xnor     g07375 ( new_n7752 , new_n7722 , new_n7751 );
  nor      g07376 ( new_n7753 , new_n7719 , new_n7752 );
  and      g07377 ( new_n7754 , new_n7719 , new_n7752 );
  nor      g07378 ( new_n7755 , new_n7753 , new_n7754 );
  xor      g07379 ( new_n7756 , new_n7687 , new_n7755 );
  xnor     g07380 ( new_n7757 , new_n7684 , new_n7756 );
  xor      g07381 ( new_n7758 , new_n7649 , new_n7757 );
  xnor     g07382 ( new_n7759 , new_n7444 , new_n7645 );
  nor      g07383 ( new_n7760 , new_n7758 , new_n7759 );
  nor      g07384 ( new_n7761 , new_n7646 , new_n7760 );
  nand     g07385 ( new_n7762 , new_n7429 , new_n7442 );
  nand g07386 ( new_n7763 , new_n7762 , new_n7762 );
  nor      g07387 ( new_n7764 , new_n7428 , new_n7443 );
  nor      g07388 ( new_n7765 , new_n7763 , new_n7764 );
  nand g07389 ( new_n7766 , new_n7406 , new_n7406 );
  nor      g07390 ( new_n7767 , new_n7766 , new_n7426 );
  nand g07391 ( new_n7768 , new_n7767 , new_n7767 );
  nand g07392 ( new_n7769 , new_n7404 , new_n7404 );
  nand     g07393 ( new_n7770 , new_n7390 , new_n7769 );
  nand g07394 ( new_n7771 , new_n7770 , new_n7770 );
  nor      g07395 ( new_n7772 , new_n7384 , new_n7405 );
  xor      g07396 ( new_n7773 , new_n7389 , new_n7772 );
  nor      g07397 ( new_n7774 , new_n7771 , new_n7773 );
  nand     g07398 ( new_n7775 , pi044 , pi133 );
  xor      g07399 ( new_n7776 , new_n7398 , new_n7775 );
  nand     g07400 ( new_n7777 , pi189 , pi250 );
  and      g07401 ( new_n7778 , pi084 , pi119 );
  xor      g07402 ( new_n7779 , new_n7777 , new_n7778 );
  xor      g07403 ( new_n7780 , new_n7396 , new_n7779 );
  xor      g07404 ( new_n7781 , new_n7776 , new_n7780 );
  nand     g07405 ( new_n7782 , new_n7395 , new_n7402 );
  nand     g07406 ( new_n7783 , new_n7394 , new_n7403 );
  nand     g07407 ( new_n7784 , new_n7782 , new_n7783 );
  nand     g07408 ( new_n7785 , pi052 , pi072 );
  nand     g07409 ( new_n7786 , pi131 , pi248 );
  xor      g07410 ( new_n7787 , new_n7785 , new_n7786 );
  xor      g07411 ( new_n7788 , new_n7388 , new_n7787 );
  xor      g07412 ( new_n7789 , new_n7784 , new_n7788 );
  xor      g07413 ( new_n7790 , new_n7781 , new_n7789 );
  xor      g07414 ( new_n7791 , new_n7774 , new_n7790 );
  nor      g07415 ( new_n7792 , new_n7768 , new_n7791 );
  and      g07416 ( new_n7793 , new_n7768 , new_n7791 );
  or       g07417 ( new_n7794 , new_n7792 , new_n7793 );
  xor      g07418 ( new_n7795 , new_n7765 , new_n7794 );
  nand     g07419 ( new_n7796 , new_n7761 , new_n7795 );
  xor      g07420 ( new_n7797 , new_n7761 , new_n7795 );
  nand     g07421 ( new_n7798 , new_n7716 , new_n7717 );
  nand     g07422 ( new_n7799 , new_n7715 , new_n7718 );
  nand     g07423 ( new_n7800 , new_n7798 , new_n7799 );
  nor      g07424 ( new_n7801 , new_n7690 , new_n7714 );
  nand     g07425 ( new_n7802 , pi114 , pi212 );
  nand     g07426 ( new_n7803 , pi091 , pi213 );
  xor      g07427 ( new_n7804 , new_n7802 , new_n7803 );
  xor      g07428 ( new_n7805 , new_n7691 , new_n7804 );
  nand     g07429 ( new_n7806 , new_n7706 , new_n7707 );
  nand     g07430 ( new_n7807 , new_n7699 , new_n7708 );
  nand     g07431 ( new_n7808 , new_n7806 , new_n7807 );
  xor      g07432 ( new_n7809 , new_n7805 , new_n7808 );
  nand     g07433 ( new_n7810 , pi164 , pi183 );
  nand     g07434 ( new_n7811 , pi032 , pi112 );
  xor      g07435 ( new_n7812 , new_n7810 , new_n7811 );
  xor      g07436 ( new_n7813 , new_n7703 , new_n7812 );
  nand     g07437 ( new_n7814 , pi013 , pi145 );
  xor      g07438 ( new_n7815 , new_n7704 , new_n7814 );
  xnor     g07439 ( new_n7816 , new_n7813 , new_n7815 );
  xor      g07440 ( new_n7817 , new_n7809 , new_n7816 );
  nor      g07441 ( new_n7818 , new_n7696 , new_n7709 );
  nand g07442 ( new_n7819 , new_n7710 , new_n7710 );
  nor      g07443 ( new_n7820 , new_n7819 , new_n7713 );
  xor      g07444 ( new_n7821 , new_n7692 , new_n7820 );
  nor      g07445 ( new_n7822 , new_n7818 , new_n7821 );
  xor      g07446 ( new_n7823 , new_n7817 , new_n7822 );
  xnor     g07447 ( new_n7824 , new_n7801 , new_n7823 );
  xnor     g07448 ( new_n7825 , new_n7800 , new_n7824 );
  nand g07449 ( new_n7826 , new_n7747 , new_n7747 );
  nor      g07450 ( new_n7827 , new_n7826 , new_n7750 );
  nand g07451 ( new_n7828 , new_n7827 , new_n7827 );
  nand     g07452 ( new_n7829 , pi056 , pi141 );
  xor      g07453 ( new_n7830 , new_n7741 , new_n7829 );
  nand     g07454 ( new_n7831 , pi018 , pi027 );
  nand     g07455 ( new_n7832 , pi008 , pi090 );
  xor      g07456 ( new_n7833 , new_n7831 , new_n7832 );
  xor      g07457 ( new_n7834 , new_n7740 , new_n7833 );
  xor      g07458 ( new_n7835 , new_n7830 , new_n7834 );
  nand     g07459 ( new_n7836 , new_n7736 , new_n7743 );
  nand     g07460 ( new_n7837 , new_n7735 , new_n7744 );
  nand     g07461 ( new_n7838 , new_n7836 , new_n7837 );
  nand     g07462 ( new_n7839 , pi096 , pi241 );
  nand     g07463 ( new_n7840 , pi235 , pi236 );
  xor      g07464 ( new_n7841 , new_n7839 , new_n7840 );
  xnor     g07465 ( new_n7842 , new_n7729 , new_n7841 );
  xor      g07466 ( new_n7843 , new_n7838 , new_n7842 );
  xnor     g07467 ( new_n7844 , new_n7835 , new_n7843 );
  nor      g07468 ( new_n7845 , new_n7732 , new_n7745 );
  nor      g07469 ( new_n7846 , new_n7725 , new_n7746 );
  xor      g07470 ( new_n7847 , new_n7730 , new_n7846 );
  nor      g07471 ( new_n7848 , new_n7845 , new_n7847 );
  xor      g07472 ( new_n7849 , new_n7844 , new_n7848 );
  nand     g07473 ( new_n7850 , new_n7828 , new_n7849 );
  or       g07474 ( new_n7851 , new_n7828 , new_n7849 );
  nand     g07475 ( new_n7852 , new_n7850 , new_n7851 );
  nand     g07476 ( new_n7853 , new_n7720 , new_n7721 );
  nand     g07477 ( new_n7854 , new_n7722 , new_n7751 );
  nand     g07478 ( new_n7855 , new_n7853 , new_n7854 );
  xor      g07479 ( new_n7856 , new_n7852 , new_n7855 );
  xor      g07480 ( new_n7857 , new_n7825 , new_n7856 );
  nor      g07481 ( new_n7858 , new_n7687 , new_n7754 );
  nor      g07482 ( new_n7859 , new_n7753 , new_n7858 );
  xnor     g07483 ( new_n7860 , new_n7857 , new_n7859 );
  nand     g07484 ( new_n7861 , new_n7652 , new_n7653 );
  nand g07485 ( new_n7862 , new_n7683 , new_n7683 );
  nand     g07486 ( new_n7863 , new_n7654 , new_n7862 );
  nand     g07487 ( new_n7864 , new_n7861 , new_n7863 );
  nor      g07488 ( new_n7865 , new_n7678 , new_n7682 );
  nand g07489 ( new_n7866 , new_n7865 , new_n7865 );
  nand     g07490 ( new_n7867 , pi146 , pi147 );
  nand     g07491 ( new_n7868 , pi015 , pi019 );
  xor      g07492 ( new_n7869 , new_n7867 , new_n7868 );
  xor      g07493 ( new_n7870 , new_n7664 , new_n7869 );
  nand     g07494 ( new_n7871 , pi035 , pi097 );
  xor      g07495 ( new_n7872 , new_n7665 , new_n7871 );
  xor      g07496 ( new_n7873 , new_n7870 , new_n7872 );
  nand     g07497 ( new_n7874 , new_n7668 , new_n7671 );
  nand     g07498 ( new_n7875 , new_n7667 , new_n7672 );
  nand     g07499 ( new_n7876 , new_n7874 , new_n7875 );
  nand     g07500 ( new_n7877 , pi093 , pi208 );
  nand     g07501 ( new_n7878 , pi166 , pi168 );
  xor      g07502 ( new_n7879 , new_n7877 , new_n7878 );
  xor      g07503 ( new_n7880 , new_n7655 , new_n7879 );
  xor      g07504 ( new_n7881 , new_n7876 , new_n7880 );
  xor      g07505 ( new_n7882 , new_n7873 , new_n7881 );
  nand     g07506 ( new_n7883 , new_n7660 , new_n7673 );
  nand     g07507 ( new_n7884 , new_n7674 , new_n7677 );
  nand     g07508 ( new_n7885 , new_n7883 , new_n7884 );
  xor      g07509 ( new_n7886 , new_n7656 , new_n7885 );
  xor      g07510 ( new_n7887 , new_n7882 , new_n7886 );
  xor      g07511 ( new_n7888 , new_n7866 , new_n7887 );
  xor      g07512 ( new_n7889 , new_n7864 , new_n7888 );
  xor      g07513 ( new_n7890 , new_n7860 , new_n7889 );
  nor      g07514 ( new_n7891 , new_n7684 , new_n7756 );
  nor      g07515 ( new_n7892 , new_n7649 , new_n7757 );
  nor      g07516 ( new_n7893 , new_n7891 , new_n7892 );
  xor      g07517 ( new_n7894 , new_n7890 , new_n7893 );
  nand     g07518 ( new_n7895 , new_n7797 , new_n7894 );
  nand     g07519 ( new_n7896 , new_n7796 , new_n7895 );
  nand     g07520 ( new_n7897 , pi146 , pi151 );
  xor      g07521 ( new_n7898 , new_n7896 , new_n7897 );
  nand g07522 ( new_n7899 , new_n7885 , new_n7885 );
  nand     g07523 ( new_n7900 , new_n7656 , new_n7899 );
  nand g07524 ( new_n7901 , new_n7886 , new_n7886 );
  nand     g07525 ( new_n7902 , new_n7882 , new_n7901 );
  nand     g07526 ( new_n7903 , new_n7900 , new_n7902 );
  nand     g07527 ( new_n7904 , pi093 , pi139 );
  xor      g07528 ( new_n7905 , new_n7903 , new_n7904 );
  nand     g07529 ( new_n7906 , pi166 , pi208 );
  nand     g07530 ( new_n7907 , pi072 , pi077 );
  xor      g07531 ( new_n7908 , new_n7906 , new_n7907 );
  nor      g07532 ( new_n7909 , new_n7666 , new_n7871 );
  nor      g07533 ( new_n7910 , new_n7870 , new_n7872 );
  nor      g07534 ( new_n7911 , new_n7909 , new_n7910 );
  xor      g07535 ( new_n7912 , new_n7908 , new_n7911 );
  xor      g07536 ( new_n7913 , new_n7905 , new_n7912 );
  xor      g07537 ( new_n7914 , new_n7898 , new_n7913 );
  or       g07538 ( new_n7915 , new_n7398 , new_n7775 );
  nand     g07539 ( new_n7916 , new_n7776 , new_n7780 );
  nand     g07540 ( new_n7917 , new_n7915 , new_n7916 );
  nand     g07541 ( new_n7918 , pi110 , pi236 );
  nand     g07542 ( new_n7919 , pi056 , pi090 );
  xor      g07543 ( new_n7920 , new_n7918 , new_n7919 );
  xor      g07544 ( new_n7921 , new_n7917 , new_n7920 );
  nand     g07545 ( new_n7922 , pi008 , pi047 );
  nand g07546 ( new_n7923 , new_n7777 , new_n7777 );
  nor      g07547 ( new_n7924 , new_n7923 , new_n7778 );
  nor      g07548 ( new_n7925 , new_n7397 , new_n7779 );
  nor      g07549 ( new_n7926 , new_n7924 , new_n7925 );
  xor      g07550 ( new_n7927 , new_n7922 , new_n7926 );
  xor      g07551 ( new_n7928 , new_n7921 , new_n7927 );
  nand     g07552 ( new_n7929 , pi019 , pi204 );
  nand     g07553 ( new_n7930 , new_n7801 , new_n7823 );
  or       g07554 ( new_n7931 , new_n7800 , new_n7824 );
  nand     g07555 ( new_n7932 , new_n7930 , new_n7931 );
  xor      g07556 ( new_n7933 , new_n7929 , new_n7932 );
  nand g07557 ( new_n7934 , new_n7825 , new_n7825 );
  nor      g07558 ( new_n7935 , new_n7934 , new_n7856 );
  nor      g07559 ( new_n7936 , new_n7857 , new_n7859 );
  nor      g07560 ( new_n7937 , new_n7935 , new_n7936 );
  xor      g07561 ( new_n7938 , new_n7933 , new_n7937 );
  nand     g07562 ( new_n7939 , pi235 , pi241 );
  nand     g07563 ( new_n7940 , new_n7692 , new_n7820 );
  or       g07564 ( new_n7941 , new_n7817 , new_n7822 );
  nand     g07565 ( new_n7942 , new_n7940 , new_n7941 );
  xor      g07566 ( new_n7943 , new_n7939 , new_n7942 );
  nand     g07567 ( new_n7944 , pi183 , pi206 );
  nand     g07568 ( new_n7945 , pi052 , pi248 );
  xor      g07569 ( new_n7946 , new_n7944 , new_n7945 );
  nand     g07570 ( new_n7947 , pi035 , pi075 );
  xor      g07571 ( new_n7948 , new_n7946 , new_n7947 );
  xor      g07572 ( new_n7949 , new_n7943 , new_n7948 );
  xor      g07573 ( new_n7950 , new_n7938 , new_n7949 );
  nand     g07574 ( new_n7951 , new_n7876 , new_n7880 );
  nand g07575 ( new_n7952 , new_n7873 , new_n7873 );
  nand     g07576 ( new_n7953 , new_n7952 , new_n7881 );
  nand     g07577 ( new_n7954 , new_n7951 , new_n7953 );
  nand     g07578 ( new_n7955 , new_n7867 , new_n7868 );
  nand     g07579 ( new_n7956 , new_n7664 , new_n7869 );
  nand     g07580 ( new_n7957 , new_n7955 , new_n7956 );
  nand     g07581 ( new_n7958 , pi011 , pi168 );
  nand     g07582 ( new_n7959 , pi088 , pi164 );
  xnor     g07583 ( new_n7960 , new_n7958 , new_n7959 );
  xor      g07584 ( new_n7961 , new_n7957 , new_n7960 );
  xor      g07585 ( new_n7962 , new_n7954 , new_n7961 );
  nand     g07586 ( new_n7963 , pi015 , pi097 );
  nand     g07587 ( new_n7964 , pi031 , pi213 );
  nand     g07588 ( new_n7965 , pi032 , pi105 );
  nand     g07589 ( new_n7966 , new_n7877 , new_n7878 );
  nand     g07590 ( new_n7967 , new_n7655 , new_n7879 );
  nand     g07591 ( new_n7968 , new_n7966 , new_n7967 );
  xnor     g07592 ( new_n7969 , new_n7965 , new_n7968 );
  xor      g07593 ( new_n7970 , new_n7964 , new_n7969 );
  xor      g07594 ( new_n7971 , new_n7963 , new_n7970 );
  xnor     g07595 ( new_n7972 , new_n7962 , new_n7971 );
  nand     g07596 ( new_n7973 , pi045 , pi084 );
  xor      g07597 ( new_n7974 , new_n7972 , new_n7973 );
  xor      g07598 ( new_n7975 , new_n7950 , new_n7974 );
  xor      g07599 ( new_n7976 , new_n7928 , new_n7975 );
  xor      g07600 ( new_n7977 , new_n7914 , new_n7976 );
  nand g07601 ( new_n7978 , new_n7889 , new_n7889 );
  nor      g07602 ( new_n7979 , new_n7860 , new_n7978 );
  nor      g07603 ( new_n7980 , new_n7890 , new_n7893 );
  nor      g07604 ( new_n7981 , new_n7979 , new_n7980 );
  nand     g07605 ( new_n7982 , new_n7805 , new_n7808 );
  nand     g07606 ( new_n7983 , new_n7809 , new_n7816 );
  nand     g07607 ( new_n7984 , new_n7982 , new_n7983 );
  nand     g07608 ( new_n7985 , pi091 , pi212 );
  nand     g07609 ( new_n7986 , pi013 , pi246 );
  nand     g07610 ( new_n7987 , pi018 , pi026 );
  xnor     g07611 ( new_n7988 , new_n7986 , new_n7987 );
  xor      g07612 ( new_n7989 , new_n7985 , new_n7988 );
  xor      g07613 ( new_n7990 , new_n7984 , new_n7989 );
  xor      g07614 ( new_n7991 , new_n7981 , new_n7990 );
  nand     g07615 ( new_n7992 , pi147 , pi152 );
  nand     g07616 ( new_n7993 , pi009 , pi131 );
  nand     g07617 ( new_n7994 , new_n7389 , new_n7772 );
  nand g07618 ( new_n7995 , new_n7774 , new_n7774 );
  nand     g07619 ( new_n7996 , new_n7995 , new_n7790 );
  nand     g07620 ( new_n7997 , new_n7994 , new_n7996 );
  nand g07621 ( new_n7998 , new_n7838 , new_n7838 );
  nor      g07622 ( new_n7999 , new_n7998 , new_n7842 );
  nor      g07623 ( new_n8000 , new_n7835 , new_n7843 );
  or       g07624 ( new_n8001 , new_n7999 , new_n8000 );
  xor      g07625 ( new_n8002 , new_n7997 , new_n8001 );
  xor      g07626 ( new_n8003 , new_n7993 , new_n8002 );
  nand     g07627 ( new_n8004 , new_n7785 , new_n7786 );
  nand     g07628 ( new_n8005 , new_n7388 , new_n7787 );
  nand     g07629 ( new_n8006 , new_n8004 , new_n8005 );
  nand     g07630 ( new_n8007 , pi064 , pi250 );
  xor      g07631 ( new_n8008 , new_n8006 , new_n8007 );
  nand     g07632 ( new_n8009 , pi096 , pi161 );
  nand     g07633 ( new_n8010 , new_n7839 , new_n7840 );
  nand     g07634 ( new_n8011 , new_n7729 , new_n7841 );
  nand     g07635 ( new_n8012 , new_n8010 , new_n8011 );
  nor      g07636 ( new_n8013 , new_n7705 , new_n7814 );
  nor      g07637 ( new_n8014 , new_n7813 , new_n7815 );
  nor      g07638 ( new_n8015 , new_n8013 , new_n8014 );
  xor      g07639 ( new_n8016 , new_n8012 , new_n8015 );
  xor      g07640 ( new_n8017 , new_n8009 , new_n8016 );
  xor      g07641 ( new_n8018 , new_n8008 , new_n8017 );
  nand     g07642 ( new_n8019 , new_n7784 , new_n7788 );
  nand g07643 ( new_n8020 , new_n7781 , new_n7781 );
  nand     g07644 ( new_n8021 , new_n8020 , new_n7789 );
  nand     g07645 ( new_n8022 , new_n8019 , new_n8021 );
  nor      g07646 ( new_n8023 , new_n7742 , new_n7829 );
  nor      g07647 ( new_n8024 , new_n7830 , new_n7834 );
  nor      g07648 ( new_n8025 , new_n8023 , new_n8024 );
  nand     g07649 ( new_n8026 , pi034 , pi119 );
  xor      g07650 ( new_n8027 , new_n8025 , new_n8026 );
  xor      g07651 ( new_n8028 , new_n8022 , new_n8027 );
  xor      g07652 ( new_n8029 , new_n8018 , new_n8028 );
  xor      g07653 ( new_n8030 , new_n8003 , new_n8029 );
  xor      g07654 ( new_n8031 , new_n7992 , new_n8030 );
  nand     g07655 ( new_n8032 , pi044 , pi189 );
  nand     g07656 ( new_n8033 , pi054 , pi133 );
  nor      g07657 ( new_n8034 , new_n7765 , new_n7792 );
  nor      g07658 ( new_n8035 , new_n7793 , new_n8034 );
  nand     g07659 ( new_n8036 , new_n7831 , new_n7832 );
  nand     g07660 ( new_n8037 , new_n7740 , new_n7833 );
  nand     g07661 ( new_n8038 , new_n8036 , new_n8037 );
  xor      g07662 ( new_n8039 , new_n8035 , new_n8038 );
  xor      g07663 ( new_n8040 , new_n8033 , new_n8039 );
  xor      g07664 ( new_n8041 , new_n8032 , new_n8040 );
  or       g07665 ( new_n8042 , new_n7866 , new_n7887 );
  nand g07666 ( new_n8043 , new_n7864 , new_n7864 );
  nand     g07667 ( new_n8044 , new_n8043 , new_n7888 );
  nand     g07668 ( new_n8045 , new_n8042 , new_n8044 );
  nand     g07669 ( new_n8046 , new_n7810 , new_n7811 );
  nand     g07670 ( new_n8047 , new_n7703 , new_n7812 );
  nand     g07671 ( new_n8048 , new_n8046 , new_n8047 );
  xor      g07672 ( new_n8049 , new_n8045 , new_n8048 );
  xor      g07673 ( new_n8050 , new_n8041 , new_n8049 );
  xor      g07674 ( new_n8051 , new_n8031 , new_n8050 );
  nand     g07675 ( new_n8052 , pi112 , pi145 );
  nand     g07676 ( new_n8053 , new_n7851 , new_n7855 );
  nand     g07677 ( new_n8054 , new_n7850 , new_n8053 );
  xor      g07678 ( new_n8055 , new_n8052 , new_n8054 );
  nand     g07679 ( new_n8056 , pi136 , pi141 );
  nand     g07680 ( new_n8057 , pi104 , pi114 );
  nand     g07681 ( new_n8058 , pi027 , pi128 );
  nand     g07682 ( new_n8059 , new_n7730 , new_n7846 );
  nand g07683 ( new_n8060 , new_n7848 , new_n7848 );
  nand     g07684 ( new_n8061 , new_n7844 , new_n8060 );
  nand     g07685 ( new_n8062 , new_n8059 , new_n8061 );
  nand     g07686 ( new_n8063 , new_n7802 , new_n7803 );
  nand     g07687 ( new_n8064 , new_n7691 , new_n7804 );
  nand     g07688 ( new_n8065 , new_n8063 , new_n8064 );
  xor      g07689 ( new_n8066 , new_n8062 , new_n8065 );
  xor      g07690 ( new_n8067 , new_n8058 , new_n8066 );
  xor      g07691 ( new_n8068 , new_n8057 , new_n8067 );
  xor      g07692 ( new_n8069 , new_n8056 , new_n8068 );
  xor      g07693 ( new_n8070 , new_n8055 , new_n8069 );
  xor      g07694 ( new_n8071 , new_n8051 , new_n8070 );
  xor      g07695 ( new_n8072 , new_n7991 , new_n8071 );
  xor      g07696 ( po039 , new_n7977 , new_n8072 );
  xor      g07697 ( po040 , new_n7758 , new_n7759 );
  nand     g07698 ( new_n8075 , pi103 , pi150 );
  nand     g07699 ( new_n8076 , pi069 , pi117 );
  nand     g07700 ( new_n8077 , pi103 , pi244 );
  nand     g07701 ( new_n8078 , pi016 , pi029 );
  or       g07702 ( new_n8079 , new_n8077 , new_n8078 );
  nand     g07703 ( new_n8080 , new_n8076 , new_n8079 );
  nand     g07704 ( new_n8081 , new_n8077 , new_n8078 );
  nand     g07705 ( new_n8082 , new_n8080 , new_n8081 );
  xor      g07706 ( new_n8083 , new_n8075 , new_n8082 );
  nand     g07707 ( new_n8084 , pi016 , pi069 );
  nand     g07708 ( new_n8085 , pi029 , pi080 );
  nand     g07709 ( new_n8086 , pi117 , pi244 );
  xor      g07710 ( new_n8087 , new_n8085 , new_n8086 );
  xor      g07711 ( new_n8088 , new_n8084 , new_n8087 );
  nand g07712 ( new_n8089 , new_n8088 , new_n8088 );
  xor      g07713 ( new_n8090 , new_n8083 , new_n8089 );
  nand g07714 ( new_n8091 , new_n5103 , new_n5103 );
  nor      g07715 ( new_n8092 , new_n8091 , new_n8076 );
  and      g07716 ( new_n8093 , new_n8079 , new_n8081 );
  or       g07717 ( new_n8094 , new_n8092 , new_n8093 );
  nor      g07718 ( new_n8095 , new_n8076 , new_n8094 );
  nand     g07719 ( new_n8096 , new_n8090 , new_n8095 );
  nand g07720 ( new_n8097 , new_n8096 , new_n8096 );
  nand     g07721 ( new_n8098 , pi016 , pi244 );
  nand     g07722 ( new_n8099 , pi029 , pi247 );
  nand     g07723 ( new_n8100 , pi069 , pi080 );
  xor      g07724 ( new_n8101 , new_n8099 , new_n8100 );
  xor      g07725 ( new_n8102 , new_n8098 , new_n8101 );
  nand     g07726 ( new_n8103 , pi117 , pi150 );
  nand     g07727 ( new_n8104 , new_n8085 , new_n8086 );
  nand     g07728 ( new_n8105 , new_n8084 , new_n8087 );
  nand     g07729 ( new_n8106 , new_n8104 , new_n8105 );
  xor      g07730 ( new_n8107 , new_n8103 , new_n8106 );
  xor      g07731 ( new_n8108 , new_n8102 , new_n8107 );
  nand     g07732 ( new_n8109 , pi103 , pi221 );
  nor      g07733 ( new_n8110 , new_n8075 , new_n8082 );
  nand     g07734 ( new_n8111 , new_n8083 , new_n8089 );
  nand g07735 ( new_n8112 , new_n8111 , new_n8111 );
  nor      g07736 ( new_n8113 , new_n8110 , new_n8112 );
  xor      g07737 ( new_n8114 , new_n8109 , new_n8113 );
  xnor     g07738 ( new_n8115 , new_n8108 , new_n8114 );
  xor      g07739 ( new_n8116 , new_n8097 , new_n8115 );
  xor      g07740 ( new_n8117 , new_n8090 , new_n8095 );
  nand     g07741 ( new_n8118 , new_n8081 , new_n8092 );
  nand     g07742 ( new_n8119 , new_n8094 , new_n8118 );
  nand     g07743 ( new_n8120 , new_n5105 , new_n5108 );
  or       g07744 ( new_n8121 , new_n5102 , new_n5110 );
  and      g07745 ( new_n8122 , new_n8120 , new_n8121 );
  nor      g07746 ( new_n8123 , new_n8119 , new_n8122 );
  nand     g07747 ( new_n8124 , pi049 , pi109 );
  nand     g07748 ( new_n8125 , pi107 , pi173 );
  xor      g07749 ( new_n8126 , new_n5086 , new_n8125 );
  xor      g07750 ( new_n8127 , new_n8124 , new_n8126 );
  xor      g07751 ( new_n8128 , new_n5087 , new_n8127 );
  nor      g07752 ( new_n8129 , new_n5093 , new_n5099 );
  nor      g07753 ( new_n8130 , new_n5092 , new_n5100 );
  nor      g07754 ( new_n8131 , new_n8129 , new_n8130 );
  xor      g07755 ( new_n8132 , new_n8128 , new_n8131 );
  nand     g07756 ( new_n8133 , pi066 , pi163 );
  xor      g07757 ( new_n8134 , new_n5094 , new_n8133 );
  nand     g07758 ( new_n8135 , pi226 , pi228 );
  xor      g07759 ( new_n8136 , new_n8134 , new_n8135 );
  xnor     g07760 ( new_n8137 , new_n5095 , new_n8136 );
  xor      g07761 ( new_n8138 , new_n8132 , new_n8137 );
  nand     g07762 ( new_n8139 , new_n5078 , new_n5084 );
  nand     g07763 ( new_n8140 , new_n5085 , new_n5101 );
  nand     g07764 ( new_n8141 , new_n8139 , new_n8140 );
  nand     g07765 ( new_n8142 , pi058 , pi175 );
  xor      g07766 ( new_n8143 , new_n5079 , new_n8142 );
  nand     g07767 ( new_n8144 , pi132 , pi240 );
  xor      g07768 ( new_n8145 , new_n8143 , new_n8144 );
  xor      g07769 ( new_n8146 , new_n5080 , new_n8145 );
  xor      g07770 ( new_n8147 , new_n8141 , new_n8146 );
  xnor     g07771 ( new_n8148 , new_n8138 , new_n8147 );
  xnor     g07772 ( new_n8149 , new_n8119 , new_n8122 );
  nor      g07773 ( new_n8150 , new_n8148 , new_n8149 );
  or       g07774 ( new_n8151 , new_n8123 , new_n8150 );
  nor      g07775 ( new_n8152 , new_n8117 , new_n8151 );
  xnor     g07776 ( new_n8153 , new_n8117 , new_n8151 );
  nand g07777 ( new_n8154 , new_n8146 , new_n8146 );
  nor      g07778 ( new_n8155 , new_n8141 , new_n8154 );
  nor      g07779 ( new_n8156 , new_n8138 , new_n8147 );
  or       g07780 ( new_n8157 , new_n8155 , new_n8156 );
  nor      g07781 ( new_n8158 , new_n5080 , new_n8145 );
  nand     g07782 ( new_n8159 , pi175 , pi211 );
  nand     g07783 ( new_n8160 , new_n5079 , new_n8142 );
  nand     g07784 ( new_n8161 , new_n8143 , new_n8144 );
  nand     g07785 ( new_n8162 , new_n8160 , new_n8161 );
  xor      g07786 ( new_n8163 , new_n8159 , new_n8162 );
  nand     g07787 ( new_n8164 , pi058 , pi134 );
  nand     g07788 ( new_n8165 , pi132 , pi149 );
  nand     g07789 ( new_n8166 , pi186 , pi240 );
  xor      g07790 ( new_n8167 , new_n8165 , new_n8166 );
  xor      g07791 ( new_n8168 , new_n8164 , new_n8167 );
  nand g07792 ( new_n8169 , new_n8168 , new_n8168 );
  xor      g07793 ( new_n8170 , new_n8163 , new_n8169 );
  xor      g07794 ( new_n8171 , new_n8158 , new_n8170 );
  nand g07795 ( new_n8172 , new_n8171 , new_n8171 );
  nand     g07796 ( new_n8173 , new_n8128 , new_n8131 );
  nand     g07797 ( new_n8174 , new_n8132 , new_n8137 );
  nand     g07798 ( new_n8175 , new_n8173 , new_n8174 );
  nor      g07799 ( new_n8176 , new_n5095 , new_n8136 );
  nand     g07800 ( new_n8177 , pi055 , pi163 );
  nand     g07801 ( new_n8178 , new_n5094 , new_n8133 );
  nand     g07802 ( new_n8179 , new_n8134 , new_n8135 );
  nand     g07803 ( new_n8180 , new_n8178 , new_n8179 );
  xor      g07804 ( new_n8181 , new_n8177 , new_n8180 );
  nand     g07805 ( new_n8182 , pi207 , pi228 );
  nand     g07806 ( new_n8183 , pi066 , pi148 );
  nand     g07807 ( new_n8184 , pi039 , pi226 );
  xor      g07808 ( new_n8185 , new_n8183 , new_n8184 );
  xor      g07809 ( new_n8186 , new_n8182 , new_n8185 );
  xor      g07810 ( new_n8187 , new_n8181 , new_n8186 );
  xor      g07811 ( new_n8188 , new_n8176 , new_n8187 );
  nand g07812 ( new_n8189 , new_n8127 , new_n8127 );
  nand     g07813 ( new_n8190 , new_n5087 , new_n8189 );
  nand     g07814 ( new_n8191 , pi107 , pi230 );
  nand     g07815 ( new_n8192 , new_n5086 , new_n8125 );
  nand     g07816 ( new_n8193 , new_n8124 , new_n8126 );
  nand     g07817 ( new_n8194 , new_n8192 , new_n8193 );
  xor      g07818 ( new_n8195 , new_n8191 , new_n8194 );
  nand     g07819 ( new_n8196 , pi171 , pi173 );
  nand     g07820 ( new_n8197 , pi109 , pi245 );
  nand     g07821 ( new_n8198 , pi014 , pi049 );
  xor      g07822 ( new_n8199 , new_n8197 , new_n8198 );
  xor      g07823 ( new_n8200 , new_n8196 , new_n8199 );
  xor      g07824 ( new_n8201 , new_n8195 , new_n8200 );
  xnor     g07825 ( new_n8202 , new_n8190 , new_n8201 );
  xnor     g07826 ( new_n8203 , new_n8188 , new_n8202 );
  xnor     g07827 ( new_n8204 , new_n8175 , new_n8203 );
  xor      g07828 ( new_n8205 , new_n8172 , new_n8204 );
  xor      g07829 ( new_n8206 , new_n8157 , new_n8205 );
  nor      g07830 ( new_n8207 , new_n8153 , new_n8206 );
  nor      g07831 ( new_n8208 , new_n8152 , new_n8207 );
  xnor     g07832 ( new_n8209 , new_n8116 , new_n8208 );
  nor      g07833 ( new_n8210 , new_n8172 , new_n8204 );
  and      g07834 ( new_n8211 , new_n8157 , new_n8205 );
  nor      g07835 ( new_n8212 , new_n8210 , new_n8211 );
  nor      g07836 ( new_n8213 , new_n8190 , new_n8201 );
  nand     g07837 ( new_n8214 , pi050 , pi107 );
  nand     g07838 ( new_n8215 , new_n8191 , new_n8194 );
  nand     g07839 ( new_n8216 , new_n8195 , new_n8200 );
  nand     g07840 ( new_n8217 , new_n8215 , new_n8216 );
  xor      g07841 ( new_n8218 , new_n8214 , new_n8217 );
  nand     g07842 ( new_n8219 , pi171 , pi230 );
  nand     g07843 ( new_n8220 , new_n8197 , new_n8198 );
  nand     g07844 ( new_n8221 , new_n8196 , new_n8199 );
  nand     g07845 ( new_n8222 , new_n8220 , new_n8221 );
  xor      g07846 ( new_n8223 , new_n8219 , new_n8222 );
  nand     g07847 ( new_n8224 , pi049 , pi173 );
  nand     g07848 ( new_n8225 , pi109 , pi201 );
  nand     g07849 ( new_n8226 , pi014 , pi245 );
  xor      g07850 ( new_n8227 , new_n8225 , new_n8226 );
  xor      g07851 ( new_n8228 , new_n8224 , new_n8227 );
  xnor     g07852 ( new_n8229 , new_n8223 , new_n8228 );
  xor      g07853 ( new_n8230 , new_n8218 , new_n8229 );
  xor      g07854 ( new_n8231 , new_n8213 , new_n8230 );
  nand g07855 ( new_n8232 , new_n8176 , new_n8176 );
  or       g07856 ( new_n8233 , new_n8232 , new_n8187 );
  nand     g07857 ( new_n8234 , pi002 , pi163 );
  nand     g07858 ( new_n8235 , new_n8177 , new_n8180 );
  nand     g07859 ( new_n8236 , new_n8181 , new_n8186 );
  nand     g07860 ( new_n8237 , new_n8235 , new_n8236 );
  xnor     g07861 ( new_n8238 , new_n8234 , new_n8237 );
  nand     g07862 ( new_n8239 , pi055 , pi148 );
  nand     g07863 ( new_n8240 , new_n8183 , new_n8184 );
  nand     g07864 ( new_n8241 , new_n8182 , new_n8185 );
  nand     g07865 ( new_n8242 , new_n8240 , new_n8241 );
  xor      g07866 ( new_n8243 , new_n8239 , new_n8242 );
  nand     g07867 ( new_n8244 , pi116 , pi226 );
  nand     g07868 ( new_n8245 , pi066 , pi228 );
  nand     g07869 ( new_n8246 , pi039 , pi207 );
  xor      g07870 ( new_n8247 , new_n8245 , new_n8246 );
  xor      g07871 ( new_n8248 , new_n8244 , new_n8247 );
  xor      g07872 ( new_n8249 , new_n8243 , new_n8248 );
  xnor     g07873 ( new_n8250 , new_n8238 , new_n8249 );
  xor      g07874 ( new_n8251 , new_n8233 , new_n8250 );
  xnor     g07875 ( new_n8252 , new_n8231 , new_n8251 );
  nor      g07876 ( new_n8253 , new_n8188 , new_n8202 );
  nor      g07877 ( new_n8254 , new_n8175 , new_n8203 );
  nor      g07878 ( new_n8255 , new_n8253 , new_n8254 );
  xnor     g07879 ( new_n8256 , new_n8252 , new_n8255 );
  nand     g07880 ( new_n8257 , new_n8158 , new_n8170 );
  nand     g07881 ( new_n8258 , pi058 , pi240 );
  nand     g07882 ( new_n8259 , pi149 , pi186 );
  nand     g07883 ( new_n8260 , pi132 , pi167 );
  xor      g07884 ( new_n8261 , new_n8259 , new_n8260 );
  xor      g07885 ( new_n8262 , new_n8258 , new_n8261 );
  nand     g07886 ( new_n8263 , new_n8165 , new_n8166 );
  nand     g07887 ( new_n8264 , new_n8164 , new_n8167 );
  nand     g07888 ( new_n8265 , new_n8263 , new_n8264 );
  nand     g07889 ( new_n8266 , pi134 , pi211 );
  xor      g07890 ( new_n8267 , new_n8265 , new_n8266 );
  xor      g07891 ( new_n8268 , new_n8262 , new_n8267 );
  nand     g07892 ( new_n8269 , pi175 , pi199 );
  nor      g07893 ( new_n8270 , new_n8159 , new_n8162 );
  nand     g07894 ( new_n8271 , new_n8163 , new_n8169 );
  nand g07895 ( new_n8272 , new_n8271 , new_n8271 );
  or       g07896 ( new_n8273 , new_n8270 , new_n8272 );
  xor      g07897 ( new_n8274 , new_n8269 , new_n8273 );
  xnor     g07898 ( new_n8275 , new_n8268 , new_n8274 );
  xnor     g07899 ( new_n8276 , new_n8257 , new_n8275 );
  xnor     g07900 ( new_n8277 , new_n8256 , new_n8276 );
  xor      g07901 ( new_n8278 , new_n8212 , new_n8277 );
  xnor     g07902 ( po041 , new_n8209 , new_n8278 );
  xnor     g07903 ( po042 , new_n7195 , new_n7196 );
  xnor     g07904 ( po043 , new_n4969 , new_n5008 );
  xor      g07905 ( po044 , new_n925 , new_n930 );
  xor      g07906 ( po045 , new_n2601 , new_n2602 );
  xor      g07907 ( po046 , new_n4934 , new_n4943 );
  nand     g07908 ( new_n8285 , pi150 , pi247 );
  nand     g07909 ( new_n8286 , pi058 , pi181 );
  xor      g07910 ( new_n8287 , new_n8285 , new_n8286 );
  nand     g07911 ( new_n8288 , pi049 , pi253 );
  nand     g07912 ( new_n8289 , pi037 , pi175 );
  xor      g07913 ( new_n8290 , new_n8288 , new_n8289 );
  xor      g07914 ( new_n8291 , new_n8287 , new_n8290 );
  nand     g07915 ( new_n8292 , pi186 , pi200 );
  nand     g07916 ( new_n8293 , pi010 , pi103 );
  xor      g07917 ( new_n8294 , new_n8292 , new_n8293 );
  nand     g07918 ( new_n8295 , pi016 , pi221 );
  nor      g07919 ( new_n8296 , new_n8103 , new_n8295 );
  nand     g07920 ( new_n8297 , pi016 , pi150 );
  nand     g07921 ( new_n8298 , pi117 , pi221 );
  and      g07922 ( new_n8299 , new_n8297 , new_n8298 );
  nor      g07923 ( new_n8300 , new_n8296 , new_n8299 );
  nand g07924 ( new_n8301 , new_n8300 , new_n8300 );
  nand     g07925 ( new_n8302 , pi069 , pi247 );
  nand     g07926 ( new_n8303 , pi029 , pi234 );
  nand     g07927 ( new_n8304 , new_n8302 , new_n8303 );
  nand     g07928 ( new_n8305 , pi069 , pi234 );
  nor      g07929 ( new_n8306 , new_n8099 , new_n8305 );
  nand g07930 ( new_n8307 , new_n8306 , new_n8306 );
  nand     g07931 ( new_n8308 , new_n8304 , new_n8307 );
  nand     g07932 ( new_n8309 , pi080 , pi244 );
  nand     g07933 ( new_n8310 , new_n8099 , new_n8100 );
  nand     g07934 ( new_n8311 , new_n8098 , new_n8101 );
  nand     g07935 ( new_n8312 , new_n8310 , new_n8311 );
  xor      g07936 ( new_n8313 , new_n8309 , new_n8312 );
  xor      g07937 ( new_n8314 , new_n8308 , new_n8313 );
  nand     g07938 ( new_n8315 , new_n8301 , new_n8314 );
  nand     g07939 ( new_n8316 , new_n8103 , new_n8106 );
  nand     g07940 ( new_n8317 , new_n8102 , new_n8107 );
  nand     g07941 ( new_n8318 , new_n8316 , new_n8317 );
  xor      g07942 ( new_n8319 , new_n8300 , new_n8314 );
  nand g07943 ( new_n8320 , new_n8319 , new_n8319 );
  nand     g07944 ( new_n8321 , new_n8318 , new_n8320 );
  nand     g07945 ( new_n8322 , new_n8315 , new_n8321 );
  nand g07946 ( new_n8323 , new_n8322 , new_n8322 );
  nand     g07947 ( new_n8324 , new_n8296 , new_n8323 );
  nand     g07948 ( new_n8325 , pi080 , pi150 );
  xor      g07949 ( new_n8326 , new_n8306 , new_n8325 );
  nand     g07950 ( new_n8327 , pi244 , pi247 );
  nand     g07951 ( new_n8328 , pi029 , pi214 );
  xor      g07952 ( new_n8329 , new_n8305 , new_n8328 );
  xor      g07953 ( new_n8330 , new_n8327 , new_n8329 );
  xor      g07954 ( new_n8331 , new_n8326 , new_n8330 );
  nand     g07955 ( new_n8332 , new_n8309 , new_n8312 );
  nand     g07956 ( new_n8333 , new_n8308 , new_n8313 );
  nand     g07957 ( new_n8334 , new_n8332 , new_n8333 );
  nand     g07958 ( new_n8335 , pi117 , pi196 );
  nand     g07959 ( new_n8336 , pi103 , pi184 );
  xor      g07960 ( new_n8337 , new_n8335 , new_n8336 );
  xnor     g07961 ( new_n8338 , new_n8295 , new_n8337 );
  xor      g07962 ( new_n8339 , new_n8334 , new_n8338 );
  xor      g07963 ( new_n8340 , new_n8331 , new_n8339 );
  xor      g07964 ( new_n8341 , new_n8296 , new_n8322 );
  or       g07965 ( new_n8342 , new_n8340 , new_n8341 );
  nand     g07966 ( new_n8343 , new_n8324 , new_n8342 );
  xor      g07967 ( new_n8344 , new_n8294 , new_n8343 );
  nand     g07968 ( new_n8345 , pi163 , pi243 );
  nand     g07969 ( new_n8346 , pi016 , pi196 );
  xnor     g07970 ( new_n8347 , new_n8345 , new_n8346 );
  nand     g07971 ( new_n8348 , pi074 , pi171 );
  xor      g07972 ( new_n8349 , new_n8347 , new_n8348 );
  xor      g07973 ( new_n8350 , new_n8344 , new_n8349 );
  nand     g07974 ( new_n8351 , pi000 , pi226 );
  nand     g07975 ( new_n8352 , pi115 , pi207 );
  nand     g07976 ( new_n8353 , pi066 , pi070 );
  xor      g07977 ( new_n8354 , new_n8352 , new_n8353 );
  xor      g07978 ( new_n8355 , new_n8351 , new_n8354 );
  nand g07979 ( new_n8356 , new_n8273 , new_n8273 );
  nor      g07980 ( new_n8357 , new_n8269 , new_n8356 );
  nor      g07981 ( new_n8358 , new_n8268 , new_n8274 );
  nor      g07982 ( new_n8359 , new_n8357 , new_n8358 );
  nand     g07983 ( new_n8360 , new_n8265 , new_n8266 );
  nand     g07984 ( new_n8361 , new_n8262 , new_n8267 );
  nand     g07985 ( new_n8362 , new_n8360 , new_n8361 );
  nand     g07986 ( new_n8363 , pi211 , pi240 );
  nand     g07987 ( new_n8364 , pi134 , pi199 );
  and      g07988 ( new_n8365 , new_n8363 , new_n8364 );
  nand     g07989 ( new_n8366 , pi199 , pi240 );
  nor      g07990 ( new_n8367 , new_n8266 , new_n8366 );
  nor      g07991 ( new_n8368 , new_n8365 , new_n8367 );
  nand     g07992 ( new_n8369 , pi167 , pi186 );
  nand     g07993 ( new_n8370 , pi132 , pi181 );
  nand     g07994 ( new_n8371 , new_n8369 , new_n8370 );
  nand     g07995 ( new_n8372 , pi181 , pi186 );
  nor      g07996 ( new_n8373 , new_n8260 , new_n8372 );
  nand g07997 ( new_n8374 , new_n8373 , new_n8373 );
  nand     g07998 ( new_n8375 , new_n8371 , new_n8374 );
  nand     g07999 ( new_n8376 , pi058 , pi149 );
  nand     g08000 ( new_n8377 , new_n8259 , new_n8260 );
  nand     g08001 ( new_n8378 , new_n8258 , new_n8261 );
  nand     g08002 ( new_n8379 , new_n8377 , new_n8378 );
  xor      g08003 ( new_n8380 , new_n8376 , new_n8379 );
  xor      g08004 ( new_n8381 , new_n8375 , new_n8380 );
  xor      g08005 ( new_n8382 , new_n8368 , new_n8381 );
  xnor     g08006 ( new_n8383 , new_n8362 , new_n8382 );
  nor      g08007 ( new_n8384 , new_n8359 , new_n8383 );
  nand     g08008 ( new_n8385 , pi134 , pi195 );
  nand     g08009 ( new_n8386 , pi175 , pi218 );
  xor      g08010 ( new_n8387 , new_n8385 , new_n8386 );
  xnor     g08011 ( new_n8388 , new_n8366 , new_n8387 );
  nand     g08012 ( new_n8389 , new_n8376 , new_n8379 );
  nand     g08013 ( new_n8390 , new_n8375 , new_n8380 );
  nand     g08014 ( new_n8391 , new_n8389 , new_n8390 );
  nand g08015 ( new_n8392 , new_n8391 , new_n8391 );
  xor      g08016 ( new_n8393 , new_n8388 , new_n8392 );
  nand     g08017 ( new_n8394 , pi149 , pi211 );
  xor      g08018 ( new_n8395 , new_n8373 , new_n8394 );
  nand     g08019 ( new_n8396 , pi132 , pi200 );
  nand     g08020 ( new_n8397 , pi058 , pi167 );
  xor      g08021 ( new_n8398 , new_n8396 , new_n8397 );
  xor      g08022 ( new_n8399 , new_n8372 , new_n8398 );
  xor      g08023 ( new_n8400 , new_n8395 , new_n8399 );
  xor      g08024 ( new_n8401 , new_n8393 , new_n8400 );
  nand g08025 ( new_n8402 , new_n8401 , new_n8401 );
  nand g08026 ( new_n8403 , new_n8381 , new_n8381 );
  nand     g08027 ( new_n8404 , new_n8368 , new_n8403 );
  nand g08028 ( new_n8405 , new_n8404 , new_n8404 );
  nor      g08029 ( new_n8406 , new_n8362 , new_n8382 );
  xor      g08030 ( new_n8407 , new_n8367 , new_n8406 );
  nor      g08031 ( new_n8408 , new_n8405 , new_n8407 );
  xor      g08032 ( new_n8409 , new_n8402 , new_n8408 );
  nor      g08033 ( new_n8410 , new_n8384 , new_n8409 );
  nor      g08034 ( new_n8411 , new_n8257 , new_n8275 );
  nand g08035 ( new_n8412 , new_n8411 , new_n8411 );
  nand     g08036 ( new_n8413 , pi175 , pi195 );
  nand     g08037 ( new_n8414 , new_n8412 , new_n8413 );
  nand g08038 ( new_n8415 , new_n8414 , new_n8414 );
  xor      g08039 ( new_n8416 , new_n8411 , new_n8413 );
  xor      g08040 ( new_n8417 , new_n8359 , new_n8383 );
  nor      g08041 ( new_n8418 , new_n8416 , new_n8417 );
  nor      g08042 ( new_n8419 , new_n8415 , new_n8418 );
  xnor     g08043 ( new_n8420 , new_n8384 , new_n8409 );
  nor      g08044 ( new_n8421 , new_n8419 , new_n8420 );
  nor      g08045 ( new_n8422 , new_n8410 , new_n8421 );
  xor      g08046 ( new_n8423 , new_n8355 , new_n8422 );
  xor      g08047 ( new_n8424 , new_n8350 , new_n8423 );
  xor      g08048 ( new_n8425 , new_n8291 , new_n8424 );
  nand     g08049 ( new_n8426 , pi002 , pi039 );
  nand     g08050 ( new_n8427 , pi132 , pi203 );
  xor      g08051 ( new_n8428 , new_n8426 , new_n8427 );
  xor      g08052 ( new_n8429 , new_n8425 , new_n8428 );
  nand     g08053 ( new_n8430 , pi039 , pi066 );
  nand     g08054 ( new_n8431 , pi116 , pi207 );
  nand     g08055 ( new_n8432 , pi070 , pi226 );
  nand     g08056 ( new_n8433 , new_n8431 , new_n8432 );
  nand     g08057 ( new_n8434 , pi070 , pi207 );
  nor      g08058 ( new_n8435 , new_n8244 , new_n8434 );
  nand g08059 ( new_n8436 , new_n8435 , new_n8435 );
  nand     g08060 ( new_n8437 , new_n8433 , new_n8436 );
  nand     g08061 ( new_n8438 , new_n8430 , new_n8437 );
  nand     g08062 ( new_n8439 , new_n8245 , new_n8246 );
  nand     g08063 ( new_n8440 , new_n8244 , new_n8247 );
  nand     g08064 ( new_n8441 , new_n8439 , new_n8440 );
  xor      g08065 ( new_n8442 , new_n8430 , new_n8437 );
  nand     g08066 ( new_n8443 , new_n8441 , new_n8442 );
  nand     g08067 ( new_n8444 , new_n8438 , new_n8443 );
  nand     g08068 ( new_n8445 , pi002 , pi228 );
  nand     g08069 ( new_n8446 , pi163 , pi239 );
  nand     g08070 ( new_n8447 , pi025 , pi148 );
  xor      g08071 ( new_n8448 , new_n8446 , new_n8447 );
  xor      g08072 ( new_n8449 , new_n8445 , new_n8448 );
  nand     g08073 ( new_n8450 , new_n8444 , new_n8449 );
  xor      g08074 ( new_n8451 , new_n8444 , new_n8449 );
  nand     g08075 ( new_n8452 , pi039 , pi055 );
  xor      g08076 ( new_n8453 , new_n8435 , new_n8452 );
  nand     g08077 ( new_n8454 , pi115 , pi226 );
  nand     g08078 ( new_n8455 , pi066 , pi116 );
  xor      g08079 ( new_n8456 , new_n8454 , new_n8455 );
  xor      g08080 ( new_n8457 , new_n8434 , new_n8456 );
  xnor     g08081 ( new_n8458 , new_n8453 , new_n8457 );
  nand     g08082 ( new_n8459 , new_n8451 , new_n8458 );
  nand     g08083 ( new_n8460 , new_n8450 , new_n8459 );
  nand     g08084 ( new_n8461 , new_n8454 , new_n8455 );
  nand     g08085 ( new_n8462 , new_n8434 , new_n8456 );
  nand     g08086 ( new_n8463 , new_n8461 , new_n8462 );
  nand     g08087 ( new_n8464 , new_n8305 , new_n8328 );
  nand     g08088 ( new_n8465 , new_n8327 , new_n8329 );
  nand     g08089 ( new_n8466 , new_n8464 , new_n8465 );
  xor      g08090 ( new_n8467 , new_n8463 , new_n8466 );
  nand     g08091 ( new_n8468 , pi063 , pi109 );
  nand     g08092 ( new_n8469 , pi173 , pi201 );
  nand     g08093 ( new_n8470 , new_n8468 , new_n8469 );
  nand     g08094 ( new_n8471 , pi014 , pi156 );
  xor      g08095 ( new_n8472 , new_n8468 , new_n8469 );
  nand     g08096 ( new_n8473 , new_n8471 , new_n8472 );
  nand     g08097 ( new_n8474 , new_n8470 , new_n8473 );
  nand     g08098 ( new_n8475 , pi029 , pi202 );
  xor      g08099 ( new_n8476 , new_n8474 , new_n8475 );
  xor      g08100 ( new_n8477 , new_n8467 , new_n8476 );
  xor      g08101 ( new_n8478 , new_n8460 , new_n8477 );
  nand     g08102 ( new_n8479 , pi014 , pi063 );
  nor      g08103 ( new_n8480 , new_n8225 , new_n8471 );
  nand g08104 ( new_n8481 , new_n8480 , new_n8480 );
  nand     g08105 ( new_n8482 , pi230 , pi245 );
  nor      g08106 ( new_n8483 , new_n8481 , new_n8482 );
  xor      g08107 ( new_n8484 , new_n8471 , new_n8472 );
  xor      g08108 ( new_n8485 , new_n8480 , new_n8482 );
  nor      g08109 ( new_n8486 , new_n8484 , new_n8485 );
  or       g08110 ( new_n8487 , new_n8483 , new_n8486 );
  nand     g08111 ( new_n8488 , pi083 , pi109 );
  xor      g08112 ( new_n8489 , new_n8487 , new_n8488 );
  xor      g08113 ( new_n8490 , new_n8479 , new_n8489 );
  nand     g08114 ( new_n8491 , new_n8446 , new_n8447 );
  nand     g08115 ( new_n8492 , new_n8445 , new_n8448 );
  nand     g08116 ( new_n8493 , new_n8491 , new_n8492 );
  xor      g08117 ( new_n8494 , new_n8490 , new_n8493 );
  nand     g08118 ( new_n8495 , pi171 , pi253 );
  nand     g08119 ( new_n8496 , pi074 , pi107 );
  nand     g08120 ( new_n8497 , new_n8495 , new_n8496 );
  nand     g08121 ( new_n8498 , pi049 , pi050 );
  xor      g08122 ( new_n8499 , new_n8495 , new_n8496 );
  nand     g08123 ( new_n8500 , new_n8498 , new_n8499 );
  nand     g08124 ( new_n8501 , new_n8497 , new_n8500 );
  nor      g08125 ( new_n8502 , new_n8436 , new_n8452 );
  nor      g08126 ( new_n8503 , new_n8453 , new_n8457 );
  nor      g08127 ( new_n8504 , new_n8502 , new_n8503 );
  xor      g08128 ( new_n8505 , new_n8501 , new_n8504 );
  nand     g08129 ( new_n8506 , new_n8367 , new_n8406 );
  or       g08130 ( new_n8507 , new_n8402 , new_n8408 );
  nand     g08131 ( new_n8508 , new_n8506 , new_n8507 );
  nor      g08132 ( new_n8509 , new_n8307 , new_n8325 );
  nor      g08133 ( new_n8510 , new_n8326 , new_n8330 );
  nor      g08134 ( new_n8511 , new_n8509 , new_n8510 );
  nand     g08135 ( new_n8512 , pi201 , pi230 );
  xor      g08136 ( new_n8513 , new_n8511 , new_n8512 );
  xor      g08137 ( new_n8514 , new_n8508 , new_n8513 );
  xor      g08138 ( new_n8515 , new_n8505 , new_n8514 );
  nand     g08139 ( new_n8516 , pi025 , pi228 );
  nand     g08140 ( new_n8517 , pi050 , pi245 );
  nand     g08141 ( new_n8518 , pi173 , pi245 );
  nand     g08142 ( new_n8519 , pi014 , pi201 );
  nand     g08143 ( new_n8520 , pi109 , pi156 );
  nand     g08144 ( new_n8521 , new_n8519 , new_n8520 );
  nand     g08145 ( new_n8522 , new_n8521 , new_n8481 );
  nand     g08146 ( new_n8523 , new_n8518 , new_n8522 );
  nand     g08147 ( new_n8524 , new_n8225 , new_n8226 );
  nand     g08148 ( new_n8525 , new_n8224 , new_n8227 );
  nand     g08149 ( new_n8526 , new_n8524 , new_n8525 );
  xor      g08150 ( new_n8527 , new_n8518 , new_n8522 );
  nand     g08151 ( new_n8528 , new_n8526 , new_n8527 );
  nand     g08152 ( new_n8529 , new_n8523 , new_n8528 );
  xor      g08153 ( new_n8530 , new_n8498 , new_n8499 );
  nand     g08154 ( new_n8531 , new_n8529 , new_n8530 );
  xor      g08155 ( new_n8532 , new_n8529 , new_n8530 );
  xor      g08156 ( new_n8533 , new_n8484 , new_n8485 );
  nand g08157 ( new_n8534 , new_n8533 , new_n8533 );
  nand     g08158 ( new_n8535 , new_n8532 , new_n8534 );
  nand     g08159 ( new_n8536 , new_n8531 , new_n8535 );
  xor      g08160 ( new_n8537 , new_n8517 , new_n8536 );
  xor      g08161 ( new_n8538 , new_n8516 , new_n8537 );
  xor      g08162 ( new_n8539 , new_n8515 , new_n8538 );
  xor      g08163 ( new_n8540 , new_n8494 , new_n8539 );
  nor      g08164 ( new_n8541 , new_n8219 , new_n8498 );
  nand     g08165 ( new_n8542 , new_n8219 , new_n8222 );
  nand     g08166 ( new_n8543 , new_n8223 , new_n8228 );
  nand     g08167 ( new_n8544 , new_n8542 , new_n8543 );
  nand     g08168 ( new_n8545 , pi049 , pi230 );
  nand     g08169 ( new_n8546 , pi050 , pi171 );
  and      g08170 ( new_n8547 , new_n8545 , new_n8546 );
  or       g08171 ( new_n8548 , new_n8541 , new_n8547 );
  xor      g08172 ( new_n8549 , new_n8526 , new_n8527 );
  xor      g08173 ( new_n8550 , new_n8548 , new_n8549 );
  nand g08174 ( new_n8551 , new_n8550 , new_n8550 );
  nor      g08175 ( new_n8552 , new_n8544 , new_n8551 );
  nand     g08176 ( new_n8553 , new_n8541 , new_n8552 );
  nor      g08177 ( new_n8554 , new_n8548 , new_n8549 );
  xor      g08178 ( new_n8555 , new_n8541 , new_n8552 );
  nor      g08179 ( new_n8556 , new_n8554 , new_n8555 );
  nand g08180 ( new_n8557 , new_n8556 , new_n8556 );
  xor      g08181 ( new_n8558 , new_n8532 , new_n8533 );
  nand     g08182 ( new_n8559 , new_n8557 , new_n8558 );
  nand     g08183 ( new_n8560 , new_n8553 , new_n8559 );
  nand     g08184 ( new_n8561 , pi148 , pi239 );
  nand     g08185 ( new_n8562 , pi156 , pi173 );
  xor      g08186 ( new_n8563 , new_n8561 , new_n8562 );
  xor      g08187 ( new_n8564 , new_n8560 , new_n8563 );
  nor      g08188 ( new_n8565 , new_n8214 , new_n8217 );
  and      g08189 ( new_n8566 , new_n8218 , new_n8229 );
  nor      g08190 ( new_n8567 , new_n8565 , new_n8566 );
  xor      g08191 ( new_n8568 , new_n8544 , new_n8550 );
  nor      g08192 ( new_n8569 , new_n8567 , new_n8568 );
  nand g08193 ( new_n8570 , new_n8569 , new_n8569 );
  xor      g08194 ( new_n8571 , new_n8556 , new_n8558 );
  nand     g08195 ( new_n8572 , new_n8570 , new_n8571 );
  nor      g08196 ( new_n8573 , new_n8570 , new_n8571 );
  nand     g08197 ( new_n8574 , new_n8213 , new_n8230 );
  nand     g08198 ( new_n8575 , pi107 , pi253 );
  or       g08199 ( new_n8576 , new_n8574 , new_n8575 );
  nand     g08200 ( new_n8577 , new_n8574 , new_n8575 );
  xor      g08201 ( new_n8578 , new_n8567 , new_n8568 );
  nand     g08202 ( new_n8579 , new_n8577 , new_n8578 );
  nand     g08203 ( new_n8580 , new_n8576 , new_n8579 );
  or       g08204 ( new_n8581 , new_n8573 , new_n8580 );
  nand     g08205 ( new_n8582 , new_n8572 , new_n8581 );
  xor      g08206 ( new_n8583 , new_n8318 , new_n8320 );
  nand     g08207 ( new_n8584 , new_n8109 , new_n8113 );
  nand     g08208 ( new_n8585 , new_n8108 , new_n8114 );
  nand     g08209 ( new_n8586 , new_n8584 , new_n8585 );
  nor      g08210 ( new_n8587 , new_n8583 , new_n8586 );
  xor      g08211 ( new_n8588 , new_n8340 , new_n8341 );
  nand     g08212 ( new_n8589 , new_n8587 , new_n8588 );
  xor      g08213 ( new_n8590 , new_n8583 , new_n8586 );
  nand g08214 ( new_n8591 , new_n8590 , new_n8590 );
  nand     g08215 ( new_n8592 , pi103 , pi196 );
  nor      g08216 ( new_n8593 , new_n8591 , new_n8592 );
  nand     g08217 ( new_n8594 , new_n8097 , new_n8115 );
  xor      g08218 ( new_n8595 , new_n8590 , new_n8592 );
  nor      g08219 ( new_n8596 , new_n8594 , new_n8595 );
  nor      g08220 ( new_n8597 , new_n8593 , new_n8596 );
  xor      g08221 ( new_n8598 , new_n8587 , new_n8588 );
  nand g08222 ( new_n8599 , new_n8598 , new_n8598 );
  or       g08223 ( new_n8600 , new_n8597 , new_n8599 );
  nand     g08224 ( new_n8601 , new_n8589 , new_n8600 );
  xor      g08225 ( new_n8602 , new_n8582 , new_n8601 );
  xor      g08226 ( new_n8603 , new_n8564 , new_n8602 );
  xor      g08227 ( new_n8604 , new_n8540 , new_n8603 );
  xor      g08228 ( new_n8605 , new_n8478 , new_n8604 );
  xor      g08229 ( new_n8606 , new_n8597 , new_n8599 );
  xnor     g08230 ( new_n8607 , new_n8419 , new_n8420 );
  xor      g08231 ( new_n8608 , new_n8416 , new_n8417 );
  nor      g08232 ( new_n8609 , new_n8256 , new_n8276 );
  nor      g08233 ( new_n8610 , new_n8212 , new_n8277 );
  nor      g08234 ( new_n8611 , new_n8609 , new_n8610 );
  or       g08235 ( new_n8612 , new_n8608 , new_n8611 );
  xor      g08236 ( new_n8613 , new_n8608 , new_n8611 );
  and      g08237 ( new_n8614 , new_n8231 , new_n8251 );
  nor      g08238 ( new_n8615 , new_n8252 , new_n8255 );
  or       g08239 ( new_n8616 , new_n8614 , new_n8615 );
  nor      g08240 ( new_n8617 , new_n8234 , new_n8237 );
  nor      g08241 ( new_n8618 , new_n8238 , new_n8249 );
  nor      g08242 ( new_n8619 , new_n8617 , new_n8618 );
  xor      g08243 ( new_n8620 , new_n8441 , new_n8442 );
  nand     g08244 ( new_n8621 , new_n8239 , new_n8242 );
  nand     g08245 ( new_n8622 , new_n8243 , new_n8248 );
  and      g08246 ( new_n8623 , new_n8621 , new_n8622 );
  nand     g08247 ( new_n8624 , pi055 , pi228 );
  nand     g08248 ( new_n8625 , pi002 , pi148 );
  and      g08249 ( new_n8626 , new_n8624 , new_n8625 );
  nor      g08250 ( new_n8627 , new_n8239 , new_n8445 );
  nor      g08251 ( new_n8628 , new_n8626 , new_n8627 );
  xnor     g08252 ( new_n8629 , new_n8623 , new_n8628 );
  xor      g08253 ( new_n8630 , new_n8620 , new_n8629 );
  xor      g08254 ( new_n8631 , new_n8619 , new_n8630 );
  or       g08255 ( new_n8632 , new_n8233 , new_n8250 );
  nand     g08256 ( new_n8633 , pi025 , pi163 );
  xor      g08257 ( new_n8634 , new_n8632 , new_n8633 );
  xnor     g08258 ( new_n8635 , new_n8631 , new_n8634 );
  xnor     g08259 ( new_n8636 , new_n8616 , new_n8635 );
  nand     g08260 ( new_n8637 , new_n8576 , new_n8577 );
  xor      g08261 ( new_n8638 , new_n8578 , new_n8637 );
  xor      g08262 ( new_n8639 , new_n8636 , new_n8638 );
  nand     g08263 ( new_n8640 , new_n8613 , new_n8639 );
  nand     g08264 ( new_n8641 , new_n8612 , new_n8640 );
  and      g08265 ( new_n8642 , new_n8616 , new_n8635 );
  nor      g08266 ( new_n8643 , new_n8636 , new_n8638 );
  nor      g08267 ( new_n8644 , new_n8642 , new_n8643 );
  nand g08268 ( new_n8645 , new_n8619 , new_n8619 );
  and      g08269 ( new_n8646 , new_n8645 , new_n8630 );
  nor      g08270 ( new_n8647 , new_n8623 , new_n8628 );
  nand g08271 ( new_n8648 , new_n8620 , new_n8620 );
  nor      g08272 ( new_n8649 , new_n8648 , new_n8629 );
  nor      g08273 ( new_n8650 , new_n8647 , new_n8649 );
  xnor     g08274 ( new_n8651 , new_n8627 , new_n8650 );
  nand g08275 ( new_n8652 , new_n8651 , new_n8651 );
  xnor     g08276 ( new_n8653 , new_n8451 , new_n8458 );
  xor      g08277 ( new_n8654 , new_n8652 , new_n8653 );
  xor      g08278 ( new_n8655 , new_n8646 , new_n8654 );
  nand     g08279 ( new_n8656 , new_n8632 , new_n8633 );
  nand     g08280 ( new_n8657 , new_n8631 , new_n8634 );
  nand     g08281 ( new_n8658 , new_n8656 , new_n8657 );
  xor      g08282 ( new_n8659 , new_n8655 , new_n8658 );
  xor      g08283 ( new_n8660 , new_n8570 , new_n8571 );
  xor      g08284 ( new_n8661 , new_n8580 , new_n8660 );
  xor      g08285 ( new_n8662 , new_n8659 , new_n8661 );
  xor      g08286 ( new_n8663 , new_n8644 , new_n8662 );
  xor      g08287 ( new_n8664 , new_n8641 , new_n8663 );
  xor      g08288 ( new_n8665 , new_n8607 , new_n8664 );
  nand     g08289 ( new_n8666 , new_n8606 , new_n8665 );
  xor      g08290 ( new_n8667 , new_n8594 , new_n8595 );
  nor      g08291 ( new_n8668 , new_n8116 , new_n8208 );
  nor      g08292 ( new_n8669 , new_n8209 , new_n8278 );
  nor      g08293 ( new_n8670 , new_n8668 , new_n8669 );
  nor      g08294 ( new_n8671 , new_n8667 , new_n8670 );
  xnor     g08295 ( new_n8672 , new_n8667 , new_n8670 );
  xor      g08296 ( new_n8673 , new_n8613 , new_n8639 );
  nor      g08297 ( new_n8674 , new_n8672 , new_n8673 );
  nor      g08298 ( new_n8675 , new_n8671 , new_n8674 );
  xor      g08299 ( new_n8676 , new_n8606 , new_n8665 );
  nand     g08300 ( new_n8677 , new_n8675 , new_n8676 );
  nand     g08301 ( new_n8678 , new_n8666 , new_n8677 );
  nand     g08302 ( new_n8679 , pi107 , pi205 );
  xor      g08303 ( new_n8680 , new_n8678 , new_n8679 );
  nand     g08304 ( new_n8681 , pi080 , pi221 );
  nand     g08305 ( new_n8682 , pi234 , pi244 );
  nand     g08306 ( new_n8683 , pi055 , pi116 );
  xor      g08307 ( new_n8684 , new_n8682 , new_n8683 );
  xor      g08308 ( new_n8685 , new_n8681 , new_n8684 );
  xor      g08309 ( new_n8686 , new_n8680 , new_n8685 );
  xor      g08310 ( new_n8687 , new_n8605 , new_n8686 );
  xor      g08311 ( new_n8688 , new_n8429 , new_n8687 );
  nor      g08312 ( new_n8689 , new_n8641 , new_n8663 );
  nand g08313 ( new_n8690 , new_n8664 , new_n8664 );
  nor      g08314 ( new_n8691 , new_n8607 , new_n8690 );
  nor      g08315 ( new_n8692 , new_n8689 , new_n8691 );
  nor      g08316 ( new_n8693 , new_n8374 , new_n8394 );
  nor      g08317 ( new_n8694 , new_n8395 , new_n8399 );
  nor      g08318 ( new_n8695 , new_n8693 , new_n8694 );
  nand     g08319 ( new_n8696 , pi134 , pi218 );
  xor      g08320 ( new_n8697 , new_n8695 , new_n8696 );
  nand     g08321 ( new_n8698 , pi167 , pi211 );
  or       g08322 ( new_n8699 , new_n8646 , new_n8654 );
  nand     g08323 ( new_n8700 , new_n8655 , new_n8658 );
  nand     g08324 ( new_n8701 , new_n8699 , new_n8700 );
  xor      g08325 ( new_n8702 , new_n8698 , new_n8701 );
  nor      g08326 ( new_n8703 , new_n8388 , new_n8392 );
  nand g08327 ( new_n8704 , new_n8393 , new_n8393 );
  nor      g08328 ( new_n8705 , new_n8704 , new_n8400 );
  nor      g08329 ( new_n8706 , new_n8703 , new_n8705 );
  nand     g08330 ( new_n8707 , new_n8627 , new_n8650 );
  nand     g08331 ( new_n8708 , new_n8652 , new_n8653 );
  nand     g08332 ( new_n8709 , new_n8707 , new_n8708 );
  nand     g08333 ( new_n8710 , new_n8396 , new_n8397 );
  nand     g08334 ( new_n8711 , new_n8372 , new_n8398 );
  nand     g08335 ( new_n8712 , new_n8710 , new_n8711 );
  nand     g08336 ( new_n8713 , new_n8385 , new_n8386 );
  nand     g08337 ( new_n8714 , new_n8366 , new_n8387 );
  nand     g08338 ( new_n8715 , new_n8713 , new_n8714 );
  xor      g08339 ( new_n8716 , new_n8712 , new_n8715 );
  xor      g08340 ( new_n8717 , new_n8709 , new_n8716 );
  xor      g08341 ( new_n8718 , new_n8706 , new_n8717 );
  xor      g08342 ( new_n8719 , new_n8702 , new_n8718 );
  xor      g08343 ( new_n8720 , new_n8697 , new_n8719 );
  xor      g08344 ( new_n8721 , new_n8692 , new_n8720 );
  nand     g08345 ( new_n8722 , pi117 , pi184 );
  nand g08346 ( new_n8723 , new_n8659 , new_n8659 );
  nor      g08347 ( new_n8724 , new_n8723 , new_n8661 );
  nand g08348 ( new_n8725 , new_n8644 , new_n8644 );
  nor      g08349 ( new_n8726 , new_n8725 , new_n8662 );
  nor      g08350 ( new_n8727 , new_n8724 , new_n8726 );
  xor      g08351 ( new_n8728 , new_n8722 , new_n8727 );
  nand     g08352 ( new_n8729 , new_n8335 , new_n8336 );
  nand     g08353 ( new_n8730 , new_n8295 , new_n8337 );
  nand     g08354 ( new_n8731 , new_n8729 , new_n8730 );
  xor      g08355 ( new_n8732 , new_n8728 , new_n8731 );
  xor      g08356 ( new_n8733 , new_n8721 , new_n8732 );
  nand     g08357 ( new_n8734 , pi069 , pi214 );
  nand     g08358 ( new_n8735 , pi195 , pi240 );
  nand g08359 ( new_n8736 , new_n8334 , new_n8334 );
  nor      g08360 ( new_n8737 , new_n8736 , new_n8338 );
  nor      g08361 ( new_n8738 , new_n8331 , new_n8339 );
  nor      g08362 ( new_n8739 , new_n8737 , new_n8738 );
  nand     g08363 ( new_n8740 , pi149 , pi199 );
  xor      g08364 ( new_n8741 , new_n8739 , new_n8740 );
  xor      g08365 ( new_n8742 , new_n8735 , new_n8741 );
  xor      g08366 ( new_n8743 , new_n8734 , new_n8742 );
  xor      g08367 ( new_n8744 , new_n8733 , new_n8743 );
  xor      g08368 ( po047 , new_n8688 , new_n8744 );
  xnor     g08369 ( po048 , new_n4924 , new_n4925 );
  xor      g08370 ( po049 , new_n3184 , new_n3185 );
  nand     g08371 ( new_n8748 , new_n1191 , new_n1201 );
  nand g08372 ( new_n8749 , new_n8748 , new_n8748 );
  nand     g08373 ( new_n8750 , pi231 , pi236 );
  nor      g08374 ( new_n8751 , new_n1198 , new_n1199 );
  nor      g08375 ( new_n8752 , new_n1196 , new_n1200 );
  nor      g08376 ( new_n8753 , new_n8751 , new_n8752 );
  xor      g08377 ( new_n8754 , new_n8750 , new_n8753 );
  nand     g08378 ( new_n8755 , pi161 , pi252 );
  nand     g08379 ( new_n8756 , pi090 , pi242 );
  nand     g08380 ( new_n8757 , pi140 , pi141 );
  xor      g08381 ( new_n8758 , new_n8756 , new_n8757 );
  xor      g08382 ( new_n8759 , new_n8755 , new_n8758 );
  nand     g08383 ( new_n8760 , pi121 , pi241 );
  nand     g08384 ( new_n8761 , new_n1193 , new_n1194 );
  nand     g08385 ( new_n8762 , new_n1192 , new_n1195 );
  nand     g08386 ( new_n8763 , new_n8761 , new_n8762 );
  xor      g08387 ( new_n8764 , new_n8760 , new_n8763 );
  xnor     g08388 ( new_n8765 , new_n8759 , new_n8764 );
  xor      g08389 ( new_n8766 , new_n8754 , new_n8765 );
  xor      g08390 ( new_n8767 , new_n8749 , new_n8766 );
  nand g08391 ( new_n8768 , new_n1204 , new_n1204 );
  nor      g08392 ( new_n8769 , new_n8768 , new_n1214 );
  nand     g08393 ( new_n8770 , pi213 , pi255 );
  nand     g08394 ( new_n8771 , new_n1211 , new_n1212 );
  nand     g08395 ( new_n8772 , new_n1209 , new_n1213 );
  nand     g08396 ( new_n8773 , new_n8771 , new_n8772 );
  xor      g08397 ( new_n8774 , new_n8770 , new_n8773 );
  nand     g08398 ( new_n8775 , pi024 , pi104 );
  nand     g08399 ( new_n8776 , pi013 , pi111 );
  nand     g08400 ( new_n8777 , pi112 , pi210 );
  xor      g08401 ( new_n8778 , new_n8776 , new_n8777 );
  xor      g08402 ( new_n8779 , new_n8775 , new_n8778 );
  nand     g08403 ( new_n8780 , pi212 , pi224 );
  nand     g08404 ( new_n8781 , new_n1206 , new_n1207 );
  nand     g08405 ( new_n8782 , new_n1205 , new_n1208 );
  nand     g08406 ( new_n8783 , new_n8781 , new_n8782 );
  xor      g08407 ( new_n8784 , new_n8780 , new_n8783 );
  xnor     g08408 ( new_n8785 , new_n8779 , new_n8784 );
  xor      g08409 ( new_n8786 , new_n8774 , new_n8785 );
  xor      g08410 ( new_n8787 , new_n8769 , new_n8786 );
  nor      g08411 ( new_n8788 , new_n1202 , new_n1215 );
  and      g08412 ( new_n8789 , new_n1216 , new_n1219 );
  nor      g08413 ( new_n8790 , new_n8788 , new_n8789 );
  xor      g08414 ( new_n8791 , new_n8787 , new_n8790 );
  xor      g08415 ( new_n8792 , new_n8767 , new_n8791 );
  nand     g08416 ( new_n8793 , new_n1220 , new_n1233 );
  nand     g08417 ( new_n8794 , new_n1190 , new_n1234 );
  and      g08418 ( new_n8795 , new_n8793 , new_n8794 );
  nand     g08419 ( new_n8796 , new_n1221 , new_n1232 );
  nand     g08420 ( new_n8797 , pi040 , pi168 );
  nand     g08421 ( new_n8798 , new_n1227 , new_n1230 );
  nand     g08422 ( new_n8799 , new_n1226 , new_n1231 );
  nand     g08423 ( new_n8800 , new_n8798 , new_n8799 );
  xor      g08424 ( new_n8801 , new_n8797 , new_n8800 );
  nand     g08425 ( new_n8802 , pi015 , pi249 );
  nand     g08426 ( new_n8803 , pi035 , pi222 );
  nand     g08427 ( new_n8804 , pi125 , pi139 );
  xor      g08428 ( new_n8805 , new_n8803 , new_n8804 );
  xor      g08429 ( new_n8806 , new_n8802 , new_n8805 );
  nand     g08430 ( new_n8807 , pi176 , pi208 );
  nand     g08431 ( new_n8808 , new_n1223 , new_n1224 );
  nand     g08432 ( new_n8809 , new_n1222 , new_n1225 );
  nand     g08433 ( new_n8810 , new_n8808 , new_n8809 );
  xor      g08434 ( new_n8811 , new_n8807 , new_n8810 );
  xor      g08435 ( new_n8812 , new_n8806 , new_n8811 );
  nand g08436 ( new_n8813 , new_n8812 , new_n8812 );
  xor      g08437 ( new_n8814 , new_n8801 , new_n8813 );
  xor      g08438 ( new_n8815 , new_n8796 , new_n8814 );
  xnor     g08439 ( new_n8816 , new_n8795 , new_n8815 );
  xnor     g08440 ( new_n8817 , new_n8792 , new_n8816 );
  nand g08441 ( new_n8818 , new_n1184 , new_n1184 );
  nand     g08442 ( new_n8819 , new_n8818 , new_n1185 );
  nand     g08443 ( new_n8820 , pi106 , pi131 );
  nand     g08444 ( new_n8821 , new_n1176 , new_n1177 );
  nand     g08445 ( new_n8822 , new_n1178 , new_n1183 );
  nand     g08446 ( new_n8823 , new_n8821 , new_n8822 );
  xor      g08447 ( new_n8824 , new_n8820 , new_n8823 );
  nand     g08448 ( new_n8825 , pi100 , pi133 );
  nand     g08449 ( new_n8826 , pi077 , pi227 );
  nand     g08450 ( new_n8827 , pi189 , pi217 );
  xor      g08451 ( new_n8828 , new_n8826 , new_n8827 );
  xor      g08452 ( new_n8829 , new_n8825 , new_n8828 );
  nand     g08453 ( new_n8830 , new_n1180 , new_n1181 );
  nand     g08454 ( new_n8831 , new_n1179 , new_n1182 );
  nand     g08455 ( new_n8832 , new_n8830 , new_n8831 );
  nand     g08456 ( new_n8833 , pi052 , pi081 );
  xor      g08457 ( new_n8834 , new_n8832 , new_n8833 );
  xor      g08458 ( new_n8835 , new_n8829 , new_n8834 );
  xor      g08459 ( new_n8836 , new_n8824 , new_n8835 );
  xor      g08460 ( new_n8837 , new_n8819 , new_n8836 );
  xor      g08461 ( new_n8838 , new_n8817 , new_n8837 );
  nand     g08462 ( new_n8839 , new_n1173 , new_n1186 );
  nand g08463 ( new_n8840 , new_n1235 , new_n1235 );
  nand     g08464 ( new_n8841 , new_n1187 , new_n8840 );
  nand     g08465 ( new_n8842 , new_n8839 , new_n8841 );
  xor      g08466 ( po050 , new_n8838 , new_n8842 );
  nand     g08467 ( new_n8844 , pi176 , pi216 );
  nand     g08468 ( new_n8845 , pi076 , pi249 );
  nand g08469 ( new_n8846 , new_n8845 , new_n8845 );
  nand     g08470 ( new_n8847 , pi079 , pi222 );
  nand g08471 ( new_n8848 , new_n8847 , new_n8847 );
  nand     g08472 ( new_n8849 , new_n8846 , new_n8848 );
  nor      g08473 ( new_n8850 , new_n8844 , new_n8849 );
  xnor     g08474 ( new_n8851 , new_n8844 , new_n8849 );
  nand     g08475 ( new_n8852 , pi076 , pi125 );
  nand     g08476 ( new_n8853 , pi249 , pi251 );
  xor      g08477 ( new_n8854 , new_n8852 , new_n8853 );
  xor      g08478 ( new_n8855 , new_n8847 , new_n8854 );
  nor      g08479 ( new_n8856 , new_n8851 , new_n8855 );
  nor      g08480 ( new_n8857 , new_n8850 , new_n8856 );
  nand     g08481 ( new_n8858 , pi020 , pi081 );
  nand     g08482 ( new_n8859 , pi060 , pi106 );
  nor      g08483 ( new_n8860 , new_n8858 , new_n8859 );
  nand     g08484 ( new_n8861 , pi217 , pi223 );
  nand     g08485 ( new_n8862 , pi060 , pi100 );
  nand     g08486 ( new_n8863 , new_n8861 , new_n8862 );
  nand     g08487 ( new_n8864 , pi020 , pi227 );
  xor      g08488 ( new_n8865 , new_n8861 , new_n8862 );
  nand     g08489 ( new_n8866 , new_n8864 , new_n8865 );
  nand     g08490 ( new_n8867 , new_n8863 , new_n8866 );
  nand     g08491 ( new_n8868 , new_n8858 , new_n8867 );
  nand     g08492 ( new_n8869 , pi060 , pi227 );
  nand     g08493 ( new_n8870 , pi101 , pi217 );
  nand     g08494 ( new_n8871 , pi100 , pi223 );
  xor      g08495 ( new_n8872 , new_n8870 , new_n8871 );
  xor      g08496 ( new_n8873 , new_n8869 , new_n8872 );
  xor      g08497 ( new_n8874 , new_n8858 , new_n8867 );
  nand     g08498 ( new_n8875 , new_n8873 , new_n8874 );
  nand     g08499 ( new_n8876 , new_n8868 , new_n8875 );
  nand     g08500 ( new_n8877 , pi060 , pi081 );
  nand     g08501 ( new_n8878 , pi020 , pi106 );
  and      g08502 ( new_n8879 , new_n8877 , new_n8878 );
  or       g08503 ( new_n8880 , new_n8860 , new_n8879 );
  nand     g08504 ( new_n8881 , new_n8870 , new_n8871 );
  nand     g08505 ( new_n8882 , new_n8869 , new_n8872 );
  nand     g08506 ( new_n8883 , new_n8881 , new_n8882 );
  nand     g08507 ( new_n8884 , pi223 , pi227 );
  nand     g08508 ( new_n8885 , pi217 , pi225 );
  nand     g08509 ( new_n8886 , pi100 , pi101 );
  nand     g08510 ( new_n8887 , new_n8885 , new_n8886 );
  nand     g08511 ( new_n8888 , pi100 , pi225 );
  or       g08512 ( new_n8889 , new_n8870 , new_n8888 );
  nand     g08513 ( new_n8890 , new_n8887 , new_n8889 );
  xor      g08514 ( new_n8891 , new_n8884 , new_n8890 );
  xor      g08515 ( new_n8892 , new_n8883 , new_n8891 );
  xor      g08516 ( new_n8893 , new_n8880 , new_n8892 );
  nand g08517 ( new_n8894 , new_n8893 , new_n8893 );
  nor      g08518 ( new_n8895 , new_n8876 , new_n8894 );
  and      g08519 ( new_n8896 , new_n8860 , new_n8895 );
  nand     g08520 ( new_n8897 , pi020 , pi233 );
  nand     g08521 ( new_n8898 , pi160 , pi187 );
  xor      g08522 ( new_n8899 , new_n8897 , new_n8898 );
  xor      g08523 ( new_n8900 , new_n8859 , new_n8899 );
  nand     g08524 ( new_n8901 , new_n8884 , new_n8890 );
  nand     g08525 ( new_n8902 , new_n8883 , new_n8891 );
  nand     g08526 ( new_n8903 , new_n8901 , new_n8902 );
  xor      g08527 ( new_n8904 , new_n8900 , new_n8903 );
  nand     g08528 ( new_n8905 , pi081 , pi223 );
  xor      g08529 ( new_n8906 , new_n8889 , new_n8905 );
  nand     g08530 ( new_n8907 , pi101 , pi227 );
  nand     g08531 ( new_n8908 , pi177 , pi217 );
  xor      g08532 ( new_n8909 , new_n8907 , new_n8908 );
  xnor     g08533 ( new_n8910 , new_n8888 , new_n8909 );
  xnor     g08534 ( new_n8911 , new_n8906 , new_n8910 );
  xor      g08535 ( new_n8912 , new_n8904 , new_n8911 );
  nor      g08536 ( new_n8913 , new_n8880 , new_n8892 );
  xor      g08537 ( new_n8914 , new_n8860 , new_n8895 );
  nor      g08538 ( new_n8915 , new_n8913 , new_n8914 );
  nor      g08539 ( new_n8916 , new_n8912 , new_n8915 );
  nor      g08540 ( new_n8917 , new_n8896 , new_n8916 );
  xor      g08541 ( new_n8918 , new_n8857 , new_n8917 );
  nand     g08542 ( new_n8919 , pi142 , pi255 );
  nand     g08543 ( new_n8920 , pi071 , pi111 );
  nand g08544 ( new_n8921 , new_n8920 , new_n8920 );
  nand     g08545 ( new_n8922 , pi169 , pi210 );
  nand     g08546 ( new_n8923 , pi024 , pi142 );
  nor      g08547 ( new_n8924 , new_n8922 , new_n8923 );
  nor      g08548 ( new_n8925 , new_n8921 , new_n8924 );
  nand     g08549 ( new_n8926 , new_n8922 , new_n8923 );
  nand g08550 ( new_n8927 , new_n8926 , new_n8926 );
  nor      g08551 ( new_n8928 , new_n8925 , new_n8927 );
  nand g08552 ( new_n8929 , new_n8928 , new_n8928 );
  nand     g08553 ( new_n8930 , pi142 , pi224 );
  nor      g08554 ( new_n8931 , new_n8929 , new_n8930 );
  nand     g08555 ( new_n8932 , pi123 , pi210 );
  nand     g08556 ( new_n8933 , pi111 , pi169 );
  nand     g08557 ( new_n8934 , pi024 , pi071 );
  xor      g08558 ( new_n8935 , new_n8933 , new_n8934 );
  xor      g08559 ( new_n8936 , new_n8932 , new_n8935 );
  xor      g08560 ( new_n8937 , new_n8928 , new_n8930 );
  nor      g08561 ( new_n8938 , new_n8936 , new_n8937 );
  nor      g08562 ( new_n8939 , new_n8931 , new_n8938 );
  xor      g08563 ( new_n8940 , new_n8919 , new_n8939 );
  nand     g08564 ( new_n8941 , pi099 , pi210 );
  nand     g08565 ( new_n8942 , pi024 , pi169 );
  nand     g08566 ( new_n8943 , pi111 , pi123 );
  xor      g08567 ( new_n8944 , new_n8942 , new_n8943 );
  xor      g08568 ( new_n8945 , new_n8941 , new_n8944 );
  nand     g08569 ( new_n8946 , pi071 , pi224 );
  nand     g08570 ( new_n8947 , new_n8933 , new_n8934 );
  nand     g08571 ( new_n8948 , new_n8932 , new_n8935 );
  nand     g08572 ( new_n8949 , new_n8947 , new_n8948 );
  xor      g08573 ( new_n8950 , new_n8946 , new_n8949 );
  xnor     g08574 ( new_n8951 , new_n8945 , new_n8950 );
  xor      g08575 ( new_n8952 , new_n8940 , new_n8951 );
  xnor     g08576 ( new_n8953 , new_n8936 , new_n8937 );
  nand     g08577 ( new_n8954 , pi142 , pi210 );
  and      g08578 ( new_n8955 , new_n8921 , new_n8954 );
  nor      g08579 ( new_n8956 , new_n8926 , new_n8955 );
  nor      g08580 ( new_n8957 , new_n8924 , new_n8956 );
  nor      g08581 ( new_n8958 , new_n8920 , new_n8957 );
  nand g08582 ( new_n8959 , new_n8958 , new_n8958 );
  nor      g08583 ( new_n8960 , new_n8953 , new_n8959 );
  nand     g08584 ( new_n8961 , new_n8952 , new_n8960 );
  nand     g08585 ( new_n8962 , pi127 , pi142 );
  nand     g08586 ( new_n8963 , new_n8961 , new_n8962 );
  xor      g08587 ( new_n8964 , new_n8961 , new_n8962 );
  nand     g08588 ( new_n8965 , new_n8946 , new_n8949 );
  nand     g08589 ( new_n8966 , new_n8945 , new_n8950 );
  nand     g08590 ( new_n8967 , new_n8965 , new_n8966 );
  nand     g08591 ( new_n8968 , pi169 , pi224 );
  nand     g08592 ( new_n8969 , pi071 , pi255 );
  and      g08593 ( new_n8970 , new_n8968 , new_n8969 );
  nand     g08594 ( new_n8971 , pi169 , pi255 );
  nor      g08595 ( new_n8972 , new_n8946 , new_n8971 );
  nor      g08596 ( new_n8973 , new_n8970 , new_n8972 );
  nand     g08597 ( new_n8974 , new_n8942 , new_n8943 );
  nand     g08598 ( new_n8975 , new_n8941 , new_n8944 );
  nand     g08599 ( new_n8976 , new_n8974 , new_n8975 );
  nand     g08600 ( new_n8977 , pi024 , pi123 );
  nand     g08601 ( new_n8978 , pi023 , pi210 );
  nand     g08602 ( new_n8979 , pi099 , pi111 );
  nand     g08603 ( new_n8980 , new_n8978 , new_n8979 );
  nand     g08604 ( new_n8981 , pi023 , pi111 );
  nor      g08605 ( new_n8982 , new_n8941 , new_n8981 );
  nand g08606 ( new_n8983 , new_n8982 , new_n8982 );
  nand     g08607 ( new_n8984 , new_n8980 , new_n8983 );
  xor      g08608 ( new_n8985 , new_n8977 , new_n8984 );
  xor      g08609 ( new_n8986 , new_n8976 , new_n8985 );
  xor      g08610 ( new_n8987 , new_n8973 , new_n8986 );
  xor      g08611 ( new_n8988 , new_n8967 , new_n8987 );
  nor      g08612 ( new_n8989 , new_n8919 , new_n8939 );
  and      g08613 ( new_n8990 , new_n8940 , new_n8951 );
  nor      g08614 ( new_n8991 , new_n8989 , new_n8990 );
  xor      g08615 ( new_n8992 , new_n8988 , new_n8991 );
  nand     g08616 ( new_n8993 , new_n8964 , new_n8992 );
  nand     g08617 ( new_n8994 , new_n8963 , new_n8993 );
  nand g08618 ( new_n8995 , new_n8988 , new_n8988 );
  nor      g08619 ( new_n8996 , new_n8995 , new_n8991 );
  nor      g08620 ( new_n8997 , new_n8967 , new_n8987 );
  nand     g08621 ( new_n8998 , new_n8972 , new_n8997 );
  nand g08622 ( new_n8999 , new_n8997 , new_n8997 );
  nand g08623 ( new_n9000 , new_n8973 , new_n8973 );
  nor      g08624 ( new_n9001 , new_n9000 , new_n8986 );
  nor      g08625 ( new_n9002 , new_n8972 , new_n9001 );
  nand     g08626 ( new_n9003 , new_n8999 , new_n9002 );
  nand     g08627 ( new_n9004 , new_n8998 , new_n9003 );
  nand     g08628 ( new_n9005 , pi071 , pi127 );
  nand     g08629 ( new_n9006 , pi142 , pi232 );
  xor      g08630 ( new_n9007 , new_n9005 , new_n9006 );
  xor      g08631 ( new_n9008 , new_n8971 , new_n9007 );
  nand     g08632 ( new_n9009 , new_n8977 , new_n8984 );
  nand     g08633 ( new_n9010 , new_n8976 , new_n8985 );
  nand     g08634 ( new_n9011 , new_n9009 , new_n9010 );
  xor      g08635 ( new_n9012 , new_n9008 , new_n9011 );
  nand     g08636 ( new_n9013 , pi024 , pi099 );
  nand     g08637 ( new_n9014 , pi155 , pi210 );
  xor      g08638 ( new_n9015 , new_n8981 , new_n9014 );
  xor      g08639 ( new_n9016 , new_n9013 , new_n9015 );
  nand     g08640 ( new_n9017 , pi123 , pi224 );
  xor      g08641 ( new_n9018 , new_n8982 , new_n9017 );
  xnor     g08642 ( new_n9019 , new_n9016 , new_n9018 );
  xnor     g08643 ( new_n9020 , new_n9012 , new_n9019 );
  xor      g08644 ( new_n9021 , new_n9004 , new_n9020 );
  xor      g08645 ( new_n9022 , new_n8996 , new_n9021 );
  xor      g08646 ( new_n9023 , new_n8994 , new_n9022 );
  nand     g08647 ( new_n9024 , pi121 , pi219 );
  nand     g08648 ( new_n9025 , pi102 , pi231 );
  nor      g08649 ( new_n9026 , new_n9024 , new_n9025 );
  nand     g08650 ( new_n9027 , pi001 , pi242 );
  nand     g08651 ( new_n9028 , pi219 , pi252 );
  nand     g08652 ( new_n9029 , new_n9027 , new_n9028 );
  nand     g08653 ( new_n9030 , pi102 , pi140 );
  xor      g08654 ( new_n9031 , new_n9027 , new_n9028 );
  nand     g08655 ( new_n9032 , new_n9030 , new_n9031 );
  nand     g08656 ( new_n9033 , new_n9029 , new_n9032 );
  and      g08657 ( new_n9034 , new_n9024 , new_n9033 );
  nand     g08658 ( new_n9035 , pi102 , pi252 );
  nand     g08659 ( new_n9036 , pi001 , pi140 );
  nand     g08660 ( new_n9037 , pi122 , pi242 );
  xor      g08661 ( new_n9038 , new_n9036 , new_n9037 );
  xor      g08662 ( new_n9039 , new_n9035 , new_n9038 );
  xor      g08663 ( new_n9040 , new_n9024 , new_n9033 );
  and      g08664 ( new_n9041 , new_n9039 , new_n9040 );
  nor      g08665 ( new_n9042 , new_n9034 , new_n9041 );
  nand     g08666 ( new_n9043 , pi102 , pi121 );
  nand     g08667 ( new_n9044 , pi219 , pi231 );
  and      g08668 ( new_n9045 , new_n9043 , new_n9044 );
  nor      g08669 ( new_n9046 , new_n9026 , new_n9045 );
  or       g08670 ( new_n9047 , new_n9042 , new_n9046 );
  nand g08671 ( new_n9048 , new_n9047 , new_n9047 );
  nand     g08672 ( new_n9049 , new_n9036 , new_n9037 );
  nand     g08673 ( new_n9050 , new_n9035 , new_n9038 );
  nand     g08674 ( new_n9051 , new_n9049 , new_n9050 );
  nand     g08675 ( new_n9052 , pi001 , pi252 );
  nand     g08676 ( new_n9053 , pi122 , pi140 );
  nand     g08677 ( new_n9054 , pi135 , pi242 );
  nand     g08678 ( new_n9055 , new_n9053 , new_n9054 );
  nand     g08679 ( new_n9056 , pi135 , pi140 );
  or       g08680 ( new_n9057 , new_n9037 , new_n9056 );
  nand     g08681 ( new_n9058 , new_n9055 , new_n9057 );
  xor      g08682 ( new_n9059 , new_n9052 , new_n9058 );
  xor      g08683 ( new_n9060 , new_n9051 , new_n9059 );
  nand g08684 ( new_n9061 , new_n9060 , new_n9060 );
  xnor     g08685 ( new_n9062 , new_n9042 , new_n9046 );
  nor      g08686 ( new_n9063 , new_n9061 , new_n9062 );
  or       g08687 ( new_n9064 , new_n9048 , new_n9063 );
  xor      g08688 ( new_n9065 , new_n9026 , new_n9064 );
  nand     g08689 ( new_n9066 , pi001 , pi121 );
  xor      g08690 ( new_n9067 , new_n9057 , new_n9066 );
  nand     g08691 ( new_n9068 , pi122 , pi252 );
  nand     g08692 ( new_n9069 , pi059 , pi242 );
  xor      g08693 ( new_n9070 , new_n9068 , new_n9069 );
  xnor     g08694 ( new_n9071 , new_n9056 , new_n9070 );
  xor      g08695 ( new_n9072 , new_n9067 , new_n9071 );
  nand     g08696 ( new_n9073 , new_n9052 , new_n9058 );
  nand     g08697 ( new_n9074 , new_n9051 , new_n9059 );
  nand     g08698 ( new_n9075 , new_n9073 , new_n9074 );
  nand     g08699 ( new_n9076 , pi021 , pi087 );
  nand     g08700 ( new_n9077 , pi005 , pi219 );
  xor      g08701 ( new_n9078 , new_n9076 , new_n9077 );
  xor      g08702 ( new_n9079 , new_n9025 , new_n9078 );
  xor      g08703 ( new_n9080 , new_n9075 , new_n9079 );
  xor      g08704 ( new_n9081 , new_n9072 , new_n9080 );
  xnor     g08705 ( new_n9082 , new_n9065 , new_n9081 );
  nand     g08706 ( new_n9083 , pi087 , pi231 );
  nand     g08707 ( new_n9084 , pi102 , pi242 );
  nand     g08708 ( new_n9085 , pi087 , pi252 );
  nand     g08709 ( new_n9086 , new_n9084 , new_n9085 );
  nand     g08710 ( new_n9087 , pi140 , pi219 );
  or       g08711 ( new_n9088 , new_n9084 , new_n9085 );
  nand     g08712 ( new_n9089 , new_n9087 , new_n9088 );
  nand     g08713 ( new_n9090 , new_n9086 , new_n9089 );
  nand     g08714 ( new_n9091 , pi087 , pi121 );
  nor      g08715 ( new_n9092 , new_n9090 , new_n9091 );
  xor      g08716 ( new_n9093 , new_n9090 , new_n9091 );
  xnor     g08717 ( new_n9094 , new_n9030 , new_n9031 );
  and      g08718 ( new_n9095 , new_n9093 , new_n9094 );
  nor      g08719 ( new_n9096 , new_n9092 , new_n9095 );
  nor      g08720 ( new_n9097 , new_n9083 , new_n9096 );
  xor      g08721 ( new_n9098 , new_n9039 , new_n9040 );
  xnor     g08722 ( new_n9099 , new_n9083 , new_n9096 );
  nor      g08723 ( new_n9100 , new_n9098 , new_n9099 );
  nor      g08724 ( new_n9101 , new_n9097 , new_n9100 );
  xor      g08725 ( new_n9102 , new_n9061 , new_n9062 );
  or       g08726 ( new_n9103 , new_n9101 , new_n9102 );
  nand     g08727 ( new_n9104 , pi087 , pi242 );
  nand g08728 ( new_n9105 , new_n9104 , new_n9104 );
  nor      g08729 ( new_n9106 , new_n9087 , new_n9105 );
  and      g08730 ( new_n9107 , new_n9088 , new_n9086 );
  or       g08731 ( new_n9108 , new_n9106 , new_n9107 );
  nor      g08732 ( new_n9109 , new_n9087 , new_n9108 );
  xor      g08733 ( new_n9110 , new_n9093 , new_n9094 );
  nand     g08734 ( new_n9111 , new_n9109 , new_n9110 );
  xnor     g08735 ( new_n9112 , new_n9098 , new_n9099 );
  nor      g08736 ( new_n9113 , new_n9111 , new_n9112 );
  nand     g08737 ( new_n9114 , pi005 , pi087 );
  xnor     g08738 ( new_n9115 , new_n9101 , new_n9102 );
  xor      g08739 ( new_n9116 , new_n9114 , new_n9115 );
  nand     g08740 ( new_n9117 , new_n9113 , new_n9116 );
  nor      g08741 ( new_n9118 , new_n9103 , new_n9117 );
  nand g08742 ( new_n9119 , new_n9117 , new_n9117 );
  or       g08743 ( new_n9120 , new_n9114 , new_n9115 );
  nand     g08744 ( new_n9121 , new_n9103 , new_n9120 );
  nor      g08745 ( new_n9122 , new_n9119 , new_n9121 );
  or       g08746 ( new_n9123 , new_n9118 , new_n9122 );
  xnor     g08747 ( new_n9124 , new_n9082 , new_n9123 );
  and      g08748 ( new_n9125 , new_n9023 , new_n9124 );
  xnor     g08749 ( new_n9126 , new_n9113 , new_n9116 );
  xor      g08750 ( new_n9127 , new_n8964 , new_n8992 );
  nor      g08751 ( new_n9128 , new_n9126 , new_n9127 );
  xnor     g08752 ( new_n9129 , new_n9111 , new_n9112 );
  xor      g08753 ( new_n9130 , new_n8952 , new_n8960 );
  nand g08754 ( new_n9131 , new_n9130 , new_n9130 );
  nor      g08755 ( new_n9132 , new_n9129 , new_n9131 );
  xor      g08756 ( new_n9133 , new_n9129 , new_n9130 );
  xor      g08757 ( new_n9134 , new_n9109 , new_n9110 );
  nand     g08758 ( new_n9135 , new_n8926 , new_n8955 );
  nand     g08759 ( new_n9136 , new_n8957 , new_n9135 );
  nand     g08760 ( new_n9137 , new_n9086 , new_n9106 );
  nand     g08761 ( new_n9138 , new_n9108 , new_n9137 );
  and      g08762 ( new_n9139 , new_n9136 , new_n9138 );
  nor      g08763 ( new_n9140 , new_n9136 , new_n9138 );
  nand     g08764 ( new_n9141 , pi111 , pi142 );
  nand     g08765 ( new_n9142 , pi071 , pi210 );
  xor      g08766 ( new_n9143 , new_n9141 , new_n9142 );
  nor      g08767 ( new_n9144 , new_n9104 , new_n8954 );
  nand     g08768 ( new_n9145 , new_n9143 , new_n9144 );
  nand     g08769 ( new_n9146 , pi219 , pi242 );
  nand     g08770 ( new_n9147 , pi087 , pi140 );
  xor      g08771 ( new_n9148 , new_n9146 , new_n9147 );
  xor      g08772 ( new_n9149 , new_n9143 , new_n9144 );
  nand     g08773 ( new_n9150 , new_n9148 , new_n9149 );
  nand     g08774 ( new_n9151 , new_n9145 , new_n9150 );
  nor      g08775 ( new_n9152 , new_n9140 , new_n9151 );
  nor      g08776 ( new_n9153 , new_n9139 , new_n9152 );
  or       g08777 ( new_n9154 , new_n9134 , new_n9153 );
  xnor     g08778 ( new_n9155 , new_n9134 , new_n9153 );
  xor      g08779 ( new_n9156 , new_n8953 , new_n8959 );
  or       g08780 ( new_n9157 , new_n9155 , new_n9156 );
  nand     g08781 ( new_n9158 , new_n9154 , new_n9157 );
  nor      g08782 ( new_n9159 , new_n9133 , new_n9158 );
  nor      g08783 ( new_n9160 , new_n9132 , new_n9159 );
  nand g08784 ( new_n9161 , new_n9160 , new_n9160 );
  xor      g08785 ( new_n9162 , new_n9126 , new_n9127 );
  and      g08786 ( new_n9163 , new_n9161 , new_n9162 );
  nor      g08787 ( new_n9164 , new_n9128 , new_n9163 );
  xor      g08788 ( new_n9165 , new_n9023 , new_n9124 );
  nand g08789 ( new_n9166 , new_n9165 , new_n9165 );
  nor      g08790 ( new_n9167 , new_n9164 , new_n9166 );
  nor      g08791 ( new_n9168 , new_n9125 , new_n9167 );
  nand     g08792 ( new_n9169 , pi192 , pi249 );
  nand     g08793 ( new_n9170 , new_n8900 , new_n8903 );
  nand     g08794 ( new_n9171 , new_n8904 , new_n8911 );
  nand     g08795 ( new_n9172 , new_n9170 , new_n9171 );
  nand     g08796 ( new_n9173 , pi040 , pi138 );
  nand     g08797 ( new_n9174 , pi216 , pi222 );
  nand     g08798 ( new_n9175 , pi041 , pi125 );
  xor      g08799 ( new_n9176 , new_n8846 , new_n9175 );
  xor      g08800 ( new_n9177 , new_n9174 , new_n9176 );
  nand     g08801 ( new_n9178 , pi176 , pi182 );
  nand     g08802 ( new_n9179 , pi041 , pi222 );
  nand     g08803 ( new_n9180 , pi216 , pi249 );
  nand     g08804 ( new_n9181 , new_n9179 , new_n9180 );
  nand     g08805 ( new_n9182 , pi125 , pi182 );
  xor      g08806 ( new_n9183 , new_n9179 , new_n9180 );
  nand     g08807 ( new_n9184 , new_n9182 , new_n9183 );
  nand     g08808 ( new_n9185 , new_n9181 , new_n9184 );
  xor      g08809 ( new_n9186 , new_n9178 , new_n9185 );
  xor      g08810 ( new_n9187 , new_n9177 , new_n9186 );
  nand g08811 ( new_n9188 , new_n9187 , new_n9187 );
  nor      g08812 ( new_n9189 , new_n9173 , new_n9188 );
  nand     g08813 ( new_n9190 , pi182 , pi222 );
  nand g08814 ( new_n9191 , new_n9190 , new_n9190 );
  nand     g08815 ( new_n9192 , pi041 , pi249 );
  nand     g08816 ( new_n9193 , pi125 , pi138 );
  nor      g08817 ( new_n9194 , new_n9192 , new_n9193 );
  or       g08818 ( new_n9195 , new_n9191 , new_n9194 );
  nand     g08819 ( new_n9196 , new_n9192 , new_n9193 );
  nand     g08820 ( new_n9197 , new_n9195 , new_n9196 );
  nand     g08821 ( new_n9198 , pi138 , pi176 );
  nor      g08822 ( new_n9199 , new_n9197 , new_n9198 );
  xor      g08823 ( new_n9200 , new_n9197 , new_n9198 );
  nand g08824 ( new_n9201 , new_n9200 , new_n9200 );
  xor      g08825 ( new_n9202 , new_n9182 , new_n9183 );
  nor      g08826 ( new_n9203 , new_n9201 , new_n9202 );
  nor      g08827 ( new_n9204 , new_n9199 , new_n9203 );
  xor      g08828 ( new_n9205 , new_n9173 , new_n9187 );
  nor      g08829 ( new_n9206 , new_n9204 , new_n9205 );
  nor      g08830 ( new_n9207 , new_n9189 , new_n9206 );
  nand     g08831 ( new_n9208 , new_n8845 , new_n9175 );
  nand g08832 ( new_n9209 , new_n9176 , new_n9176 );
  nand     g08833 ( new_n9210 , new_n9174 , new_n9209 );
  nand     g08834 ( new_n9211 , new_n9208 , new_n9210 );
  nand     g08835 ( new_n9212 , pi125 , pi216 );
  nand     g08836 ( new_n9213 , pi076 , pi222 );
  nand     g08837 ( new_n9214 , pi079 , pi249 );
  nand     g08838 ( new_n9215 , new_n9213 , new_n9214 );
  nand     g08839 ( new_n9216 , new_n8849 , new_n9215 );
  xor      g08840 ( new_n9217 , new_n9212 , new_n9216 );
  xor      g08841 ( new_n9218 , new_n9211 , new_n9217 );
  nand     g08842 ( new_n9219 , new_n9178 , new_n9185 );
  nand g08843 ( new_n9220 , new_n9177 , new_n9177 );
  nand     g08844 ( new_n9221 , new_n9220 , new_n9186 );
  nand     g08845 ( new_n9222 , new_n9219 , new_n9221 );
  nand     g08846 ( new_n9223 , pi040 , pi041 );
  nor      g08847 ( new_n9224 , new_n9178 , new_n9223 );
  nand     g08848 ( new_n9225 , pi041 , pi176 );
  nand     g08849 ( new_n9226 , pi040 , pi182 );
  nand     g08850 ( new_n9227 , new_n9225 , new_n9226 );
  nand g08851 ( new_n9228 , new_n9227 , new_n9227 );
  nor      g08852 ( new_n9229 , new_n9224 , new_n9228 );
  xor      g08853 ( new_n9230 , new_n9222 , new_n9229 );
  xor      g08854 ( new_n9231 , new_n9218 , new_n9230 );
  nand g08855 ( new_n9232 , new_n9231 , new_n9231 );
  nor      g08856 ( new_n9233 , new_n9207 , new_n9232 );
  nand g08857 ( new_n9234 , new_n9229 , new_n9229 );
  nand     g08858 ( new_n9235 , new_n9222 , new_n9234 );
  nand g08859 ( new_n9236 , new_n9235 , new_n9235 );
  nand g08860 ( new_n9237 , new_n9218 , new_n9218 );
  nor      g08861 ( new_n9238 , new_n9237 , new_n9230 );
  nor      g08862 ( new_n9239 , new_n9236 , new_n9238 );
  xor      g08863 ( new_n9240 , new_n9224 , new_n9239 );
  xnor     g08864 ( new_n9241 , new_n8851 , new_n8855 );
  nand     g08865 ( new_n9242 , new_n9212 , new_n9216 );
  nand     g08866 ( new_n9243 , new_n9211 , new_n9217 );
  nand     g08867 ( new_n9244 , new_n9242 , new_n9243 );
  nand     g08868 ( new_n9245 , pi174 , pi182 );
  nand     g08869 ( new_n9246 , pi138 , pi157 );
  xor      g08870 ( new_n9247 , new_n9245 , new_n9246 );
  xor      g08871 ( new_n9248 , new_n9223 , new_n9247 );
  xor      g08872 ( new_n9249 , new_n9244 , new_n9248 );
  xnor     g08873 ( new_n9250 , new_n9241 , new_n9249 );
  xor      g08874 ( new_n9251 , new_n9240 , new_n9250 );
  nand     g08875 ( new_n9252 , new_n9233 , new_n9251 );
  nand     g08876 ( new_n9253 , pi138 , pi174 );
  xor      g08877 ( new_n9254 , new_n9204 , new_n9205 );
  nand     g08878 ( new_n9255 , pi138 , pi249 );
  nand g08879 ( new_n9256 , new_n9255 , new_n9255 );
  nor      g08880 ( new_n9257 , new_n9190 , new_n9256 );
  nor      g08881 ( new_n9258 , new_n9196 , new_n9257 );
  nor      g08882 ( new_n9259 , new_n9194 , new_n9258 );
  nor      g08883 ( new_n9260 , new_n9190 , new_n9259 );
  xor      g08884 ( new_n9261 , new_n9200 , new_n9202 );
  nand g08885 ( new_n9262 , new_n9261 , new_n9261 );
  nand     g08886 ( new_n9263 , new_n9260 , new_n9262 );
  nand g08887 ( new_n9264 , new_n9263 , new_n9263 );
  nand     g08888 ( new_n9265 , new_n9254 , new_n9264 );
  nand     g08889 ( new_n9266 , new_n9253 , new_n9265 );
  xor      g08890 ( new_n9267 , new_n9253 , new_n9265 );
  xor      g08891 ( new_n9268 , new_n9207 , new_n9231 );
  nand     g08892 ( new_n9269 , new_n9267 , new_n9268 );
  nand     g08893 ( new_n9270 , new_n9266 , new_n9269 );
  nand g08894 ( new_n9271 , new_n9270 , new_n9270 );
  xor      g08895 ( new_n9272 , new_n9233 , new_n9251 );
  nand     g08896 ( new_n9273 , new_n9271 , new_n9272 );
  nand     g08897 ( new_n9274 , new_n9252 , new_n9273 );
  nand     g08898 ( new_n9275 , pi017 , pi138 );
  nand     g08899 ( new_n9276 , pi142 , pi191 );
  xor      g08900 ( new_n9277 , new_n9275 , new_n9276 );
  xor      g08901 ( new_n9278 , new_n9274 , new_n9277 );
  xor      g08902 ( new_n9279 , new_n9172 , new_n9278 );
  xor      g08903 ( new_n9280 , new_n9169 , new_n9279 );
  xor      g08904 ( new_n9281 , new_n9168 , new_n9280 );
  nand     g08905 ( new_n9282 , pi106 , pi223 );
  or       g08906 ( new_n9283 , new_n8889 , new_n8905 );
  nand     g08907 ( new_n9284 , new_n8906 , new_n8910 );
  nand     g08908 ( new_n9285 , new_n9283 , new_n9284 );
  nand     g08909 ( new_n9286 , pi081 , pi101 );
  nand     g08910 ( new_n9287 , pi100 , pi177 );
  xor      g08911 ( new_n9288 , new_n9286 , new_n9287 );
  xor      g08912 ( new_n9289 , new_n9285 , new_n9288 );
  xor      g08913 ( new_n9290 , new_n9282 , new_n9289 );
  nand     g08914 ( new_n9291 , pi086 , pi210 );
  nand     g08915 ( new_n9292 , new_n8897 , new_n8898 );
  nand     g08916 ( new_n9293 , new_n8859 , new_n8899 );
  nand     g08917 ( new_n9294 , new_n9292 , new_n9293 );
  nand     g08918 ( new_n9295 , new_n9224 , new_n9239 );
  nand     g08919 ( new_n9296 , new_n9240 , new_n9250 );
  nand     g08920 ( new_n9297 , new_n9295 , new_n9296 );
  nand     g08921 ( new_n9298 , new_n8907 , new_n8908 );
  nand     g08922 ( new_n9299 , new_n8888 , new_n8909 );
  nand     g08923 ( new_n9300 , new_n9298 , new_n9299 );
  nand     g08924 ( new_n9301 , pi222 , pi251 );
  xor      g08925 ( new_n9302 , new_n9300 , new_n9301 );
  xor      g08926 ( new_n9303 , new_n9297 , new_n9302 );
  xor      g08927 ( new_n9304 , new_n9294 , new_n9303 );
  xor      g08928 ( new_n9305 , new_n9291 , new_n9304 );
  xor      g08929 ( new_n9306 , new_n9290 , new_n9305 );
  xor      g08930 ( new_n9307 , new_n9270 , new_n9272 );
  xor      g08931 ( new_n9308 , new_n9164 , new_n9165 );
  nand     g08932 ( new_n9309 , new_n9307 , new_n9308 );
  xor      g08933 ( new_n9310 , new_n9267 , new_n9268 );
  xor      g08934 ( new_n9311 , new_n9160 , new_n9162 );
  nor      g08935 ( new_n9312 , new_n9310 , new_n9311 );
  xnor     g08936 ( new_n9313 , new_n9155 , new_n9156 );
  xor      g08937 ( new_n9314 , new_n9260 , new_n9261 );
  nand g08938 ( new_n9315 , new_n9314 , new_n9314 );
  nor      g08939 ( new_n9316 , new_n9313 , new_n9315 );
  xor      g08940 ( new_n9317 , new_n9104 , new_n8954 );
  nand     g08941 ( new_n9318 , new_n9256 , new_n9317 );
  nand g08942 ( new_n9319 , new_n9318 , new_n9318 );
  nand     g08943 ( new_n9320 , pi138 , pi222 );
  nand     g08944 ( new_n9321 , pi182 , pi249 );
  xor      g08945 ( new_n9322 , new_n9320 , new_n9321 );
  nor      g08946 ( new_n9323 , new_n9319 , new_n9322 );
  xor      g08947 ( new_n9324 , new_n9148 , new_n9149 );
  xor      g08948 ( new_n9325 , new_n9318 , new_n9322 );
  nor      g08949 ( new_n9326 , new_n9324 , new_n9325 );
  nor      g08950 ( new_n9327 , new_n9323 , new_n9326 );
  nor      g08951 ( new_n9328 , new_n9139 , new_n9140 );
  xor      g08952 ( new_n9329 , new_n9151 , new_n9328 );
  nand     g08953 ( new_n9330 , new_n9327 , new_n9329 );
  xnor     g08954 ( new_n9331 , new_n9327 , new_n9329 );
  nand     g08955 ( new_n9332 , new_n9196 , new_n9257 );
  nand     g08956 ( new_n9333 , new_n9259 , new_n9332 );
  or       g08957 ( new_n9334 , new_n9331 , new_n9333 );
  nand     g08958 ( new_n9335 , new_n9330 , new_n9334 );
  xor      g08959 ( new_n9336 , new_n9313 , new_n9314 );
  nor      g08960 ( new_n9337 , new_n9335 , new_n9336 );
  or       g08961 ( new_n9338 , new_n9316 , new_n9337 );
  xor      g08962 ( new_n9339 , new_n9254 , new_n9263 );
  nand     g08963 ( new_n9340 , new_n9338 , new_n9339 );
  xor      g08964 ( new_n9341 , new_n9133 , new_n9158 );
  xnor     g08965 ( new_n9342 , new_n9338 , new_n9339 );
  or       g08966 ( new_n9343 , new_n9341 , new_n9342 );
  nand     g08967 ( new_n9344 , new_n9340 , new_n9343 );
  xnor     g08968 ( new_n9345 , new_n9310 , new_n9311 );
  nor      g08969 ( new_n9346 , new_n9344 , new_n9345 );
  or       g08970 ( new_n9347 , new_n9312 , new_n9346 );
  xnor     g08971 ( new_n9348 , new_n9307 , new_n9308 );
  or       g08972 ( new_n9349 , new_n9347 , new_n9348 );
  nand     g08973 ( new_n9350 , new_n9309 , new_n9349 );
  or       g08974 ( new_n9351 , new_n9004 , new_n9020 );
  nand     g08975 ( new_n9352 , new_n9003 , new_n9351 );
  nand     g08976 ( new_n9353 , new_n9245 , new_n9246 );
  nand     g08977 ( new_n9354 , new_n9223 , new_n9247 );
  nand     g08978 ( new_n9355 , new_n9353 , new_n9354 );
  xnor     g08979 ( new_n9356 , new_n9352 , new_n9355 );
  xor      g08980 ( new_n9357 , new_n9350 , new_n9356 );
  xor      g08981 ( new_n9358 , new_n9306 , new_n9357 );
  xor      g08982 ( new_n9359 , new_n9281 , new_n9358 );
  xor      g08983 ( new_n9360 , new_n8918 , new_n9359 );
  nand     g08984 ( new_n9361 , pi123 , pi255 );
  nand     g08985 ( new_n9362 , pi041 , pi174 );
  nand     g08986 ( new_n9363 , new_n9244 , new_n9248 );
  nand     g08987 ( new_n9364 , new_n9241 , new_n9249 );
  nand     g08988 ( new_n9365 , new_n9363 , new_n9364 );
  xor      g08989 ( new_n9366 , new_n9362 , new_n9365 );
  nand     g08990 ( new_n9367 , pi157 , pi182 );
  nand     g08991 ( new_n9368 , pi111 , pi155 );
  nand     g08992 ( new_n9369 , pi040 , pi216 );
  xnor     g08993 ( new_n9370 , new_n9368 , new_n9369 );
  xor      g08994 ( new_n9371 , new_n9367 , new_n9370 );
  xor      g08995 ( new_n9372 , new_n9366 , new_n9371 );
  xor      g08996 ( new_n9373 , new_n9361 , new_n9372 );
  nand     g08997 ( new_n9374 , pi160 , pi233 );
  nand     g08998 ( new_n9375 , pi106 , pi160 );
  xor      g08999 ( new_n9376 , new_n8873 , new_n8874 );
  xor      g09000 ( new_n9377 , new_n9375 , new_n9376 );
  nand g09001 ( new_n9378 , new_n9377 , new_n9377 );
  nand     g09002 ( new_n9379 , pi081 , pi160 );
  nand     g09003 ( new_n9380 , pi160 , pi227 );
  nand     g09004 ( new_n9381 , pi020 , pi100 );
  nand     g09005 ( new_n9382 , new_n9380 , new_n9381 );
  nand     g09006 ( new_n9383 , pi060 , pi217 );
  xor      g09007 ( new_n9384 , new_n9380 , new_n9381 );
  nand     g09008 ( new_n9385 , new_n9383 , new_n9384 );
  nand     g09009 ( new_n9386 , new_n9382 , new_n9385 );
  nor      g09010 ( new_n9387 , new_n9379 , new_n9386 );
  xor      g09011 ( new_n9388 , new_n8864 , new_n8865 );
  xnor     g09012 ( new_n9389 , new_n9379 , new_n9386 );
  nor      g09013 ( new_n9390 , new_n9388 , new_n9389 );
  nor      g09014 ( new_n9391 , new_n9387 , new_n9390 );
  xor      g09015 ( new_n9392 , new_n9378 , new_n9391 );
  xor      g09016 ( new_n9393 , new_n9383 , new_n9384 );
  nand g09017 ( new_n9394 , new_n9393 , new_n9393 );
  nand     g09018 ( new_n9395 , pi100 , pi160 );
  nand     g09019 ( new_n9396 , pi020 , pi217 );
  nor      g09020 ( new_n9397 , new_n9395 , new_n9396 );
  nand     g09021 ( new_n9398 , new_n9394 , new_n9397 );
  nand g09022 ( new_n9399 , new_n9398 , new_n9398 );
  xor      g09023 ( new_n9400 , new_n9388 , new_n9389 );
  nand     g09024 ( new_n9401 , new_n9399 , new_n9400 );
  nand g09025 ( new_n9402 , new_n9401 , new_n9401 );
  nand     g09026 ( new_n9403 , new_n9392 , new_n9402 );
  nand     g09027 ( new_n9404 , new_n9374 , new_n9403 );
  xor      g09028 ( new_n9405 , new_n9374 , new_n9403 );
  nor      g09029 ( new_n9406 , new_n9375 , new_n9376 );
  nor      g09030 ( new_n9407 , new_n9378 , new_n9391 );
  nor      g09031 ( new_n9408 , new_n9406 , new_n9407 );
  xor      g09032 ( new_n9409 , new_n8876 , new_n8893 );
  xor      g09033 ( new_n9410 , new_n9408 , new_n9409 );
  nand g09034 ( new_n9411 , new_n9410 , new_n9410 );
  nand     g09035 ( new_n9412 , new_n9405 , new_n9411 );
  nand     g09036 ( new_n9413 , new_n9404 , new_n9412 );
  or       g09037 ( new_n9414 , new_n9408 , new_n9409 );
  xnor     g09038 ( new_n9415 , new_n8912 , new_n8915 );
  xor      g09039 ( new_n9416 , new_n9414 , new_n9415 );
  xor      g09040 ( new_n9417 , new_n9413 , new_n9416 );
  xor      g09041 ( new_n9418 , new_n9347 , new_n9348 );
  nor      g09042 ( new_n9419 , new_n9417 , new_n9418 );
  xnor     g09043 ( new_n9420 , new_n9344 , new_n9345 );
  xor      g09044 ( new_n9421 , new_n9405 , new_n9410 );
  nand g09045 ( new_n9422 , new_n9421 , new_n9421 );
  nor      g09046 ( new_n9423 , new_n9420 , new_n9422 );
  xor      g09047 ( new_n9424 , new_n9394 , new_n9397 );
  nand     g09048 ( new_n9425 , pi160 , pi217 );
  xor      g09049 ( new_n9426 , new_n9255 , new_n9317 );
  nor      g09050 ( new_n9427 , new_n9425 , new_n9426 );
  xor      g09051 ( new_n9428 , new_n9395 , new_n9396 );
  nor      g09052 ( new_n9429 , new_n9427 , new_n9428 );
  xor      g09053 ( new_n9430 , new_n9427 , new_n9428 );
  nand g09054 ( new_n9431 , new_n9430 , new_n9430 );
  xnor     g09055 ( new_n9432 , new_n9324 , new_n9325 );
  nor      g09056 ( new_n9433 , new_n9431 , new_n9432 );
  nor      g09057 ( new_n9434 , new_n9429 , new_n9433 );
  nor      g09058 ( new_n9435 , new_n9424 , new_n9434 );
  xnor     g09059 ( new_n9436 , new_n9424 , new_n9434 );
  xor      g09060 ( new_n9437 , new_n9331 , new_n9333 );
  nor      g09061 ( new_n9438 , new_n9436 , new_n9437 );
  or       g09062 ( new_n9439 , new_n9435 , new_n9438 );
  xor      g09063 ( new_n9440 , new_n9335 , new_n9336 );
  nand     g09064 ( new_n9441 , new_n9439 , new_n9440 );
  xnor     g09065 ( new_n9442 , new_n9439 , new_n9440 );
  xor      g09066 ( new_n9443 , new_n9398 , new_n9400 );
  nand g09067 ( new_n9444 , new_n9443 , new_n9443 );
  or       g09068 ( new_n9445 , new_n9442 , new_n9444 );
  nand     g09069 ( new_n9446 , new_n9441 , new_n9445 );
  xor      g09070 ( new_n9447 , new_n9392 , new_n9401 );
  nor      g09071 ( new_n9448 , new_n9446 , new_n9447 );
  xor      g09072 ( new_n9449 , new_n9341 , new_n9342 );
  xnor     g09073 ( new_n9450 , new_n9446 , new_n9447 );
  nor      g09074 ( new_n9451 , new_n9449 , new_n9450 );
  nor      g09075 ( new_n9452 , new_n9448 , new_n9451 );
  xor      g09076 ( new_n9453 , new_n9420 , new_n9421 );
  nor      g09077 ( new_n9454 , new_n9452 , new_n9453 );
  nor      g09078 ( new_n9455 , new_n9423 , new_n9454 );
  xnor     g09079 ( new_n9456 , new_n9417 , new_n9418 );
  nor      g09080 ( new_n9457 , new_n9455 , new_n9456 );
  nor      g09081 ( new_n9458 , new_n9419 , new_n9457 );
  nand     g09082 ( new_n9459 , new_n9008 , new_n9011 );
  nand     g09083 ( new_n9460 , new_n9012 , new_n9019 );
  nand     g09084 ( new_n9461 , new_n9459 , new_n9460 );
  nand     g09085 ( new_n9462 , pi020 , pi187 );
  xor      g09086 ( new_n9463 , new_n9461 , new_n9462 );
  nand     g09087 ( new_n9464 , pi225 , pi227 );
  xor      g09088 ( new_n9465 , new_n9463 , new_n9464 );
  xor      g09089 ( new_n9466 , new_n9458 , new_n9465 );
  nand     g09090 ( new_n9467 , new_n9068 , new_n9069 );
  nand     g09091 ( new_n9468 , new_n9056 , new_n9070 );
  nand     g09092 ( new_n9469 , new_n9467 , new_n9468 );
  nand     g09093 ( new_n9470 , pi001 , pi231 );
  xor      g09094 ( new_n9471 , new_n9469 , new_n9470 );
  nand     g09095 ( new_n9472 , pi023 , pi024 );
  nand     g09096 ( new_n9473 , pi060 , pi233 );
  nand     g09097 ( new_n9474 , pi082 , pi087 );
  nand g09098 ( new_n9475 , new_n8996 , new_n8996 );
  nor      g09099 ( new_n9476 , new_n9475 , new_n9021 );
  nor      g09100 ( new_n9477 , new_n8994 , new_n9022 );
  nor      g09101 ( new_n9478 , new_n9476 , new_n9477 );
  xor      g09102 ( new_n9479 , new_n9474 , new_n9478 );
  xor      g09103 ( new_n9480 , new_n9473 , new_n9479 );
  nand     g09104 ( new_n9481 , pi005 , pi102 );
  or       g09105 ( new_n9482 , new_n9075 , new_n9079 );
  nand     g09106 ( new_n9483 , new_n9072 , new_n9080 );
  nand     g09107 ( new_n9484 , new_n9482 , new_n9483 );
  xor      g09108 ( new_n9485 , new_n9481 , new_n9484 );
  nor      g09109 ( new_n9486 , new_n8983 , new_n9017 );
  nor      g09110 ( new_n9487 , new_n9016 , new_n9018 );
  nor      g09111 ( new_n9488 , new_n9486 , new_n9487 );
  xor      g09112 ( new_n9489 , new_n9485 , new_n9488 );
  xor      g09113 ( new_n9490 , new_n9480 , new_n9489 );
  nand     g09114 ( new_n9491 , pi127 , pi169 );
  nor      g09115 ( new_n9492 , new_n9082 , new_n9123 );
  or       g09116 ( new_n9493 , new_n9122 , new_n9492 );
  xor      g09117 ( new_n9494 , new_n9491 , new_n9493 );
  nand     g09118 ( new_n9495 , pi071 , pi232 );
  nand g09119 ( new_n9496 , new_n9064 , new_n9064 );
  nor      g09120 ( new_n9497 , new_n9026 , new_n9496 );
  nor      g09121 ( new_n9498 , new_n9065 , new_n9081 );
  nor      g09122 ( new_n9499 , new_n9497 , new_n9498 );
  xor      g09123 ( new_n9500 , new_n9495 , new_n9499 );
  xor      g09124 ( new_n9501 , new_n9494 , new_n9500 );
  xor      g09125 ( new_n9502 , new_n9490 , new_n9501 );
  nand     g09126 ( new_n9503 , pi059 , pi140 );
  nand     g09127 ( new_n9504 , pi135 , pi252 );
  xor      g09128 ( new_n9505 , new_n9503 , new_n9504 );
  nand     g09129 ( new_n9506 , pi121 , pi122 );
  xor      g09130 ( new_n9507 , new_n9505 , new_n9506 );
  xor      g09131 ( new_n9508 , new_n9502 , new_n9507 );
  xor      g09132 ( new_n9509 , new_n9472 , new_n9508 );
  nand     g09133 ( new_n9510 , new_n9414 , new_n9415 );
  nand     g09134 ( new_n9511 , new_n9413 , new_n9416 );
  nand     g09135 ( new_n9512 , new_n9510 , new_n9511 );
  nand     g09136 ( new_n9513 , pi129 , pi160 );
  nand     g09137 ( new_n9514 , new_n8852 , new_n8853 );
  nand     g09138 ( new_n9515 , new_n8847 , new_n8854 );
  nand     g09139 ( new_n9516 , new_n9514 , new_n9515 );
  xnor     g09140 ( new_n9517 , new_n9513 , new_n9516 );
  nand     g09141 ( new_n9518 , pi079 , pi125 );
  nand     g09142 ( new_n9519 , pi076 , pi176 );
  xor      g09143 ( new_n9520 , new_n9518 , new_n9519 );
  xor      g09144 ( new_n9521 , new_n9517 , new_n9520 );
  xor      g09145 ( new_n9522 , new_n9512 , new_n9521 );
  nand     g09146 ( new_n9523 , new_n9076 , new_n9077 );
  nand     g09147 ( new_n9524 , new_n9025 , new_n9078 );
  nand     g09148 ( new_n9525 , new_n9523 , new_n9524 );
  nand     g09149 ( new_n9526 , new_n9005 , new_n9006 );
  nand     g09150 ( new_n9527 , new_n8971 , new_n9007 );
  nand     g09151 ( new_n9528 , new_n9526 , new_n9527 );
  nand     g09152 ( new_n9529 , pi094 , pi242 );
  nand     g09153 ( new_n9530 , new_n8981 , new_n9014 );
  nand     g09154 ( new_n9531 , new_n9013 , new_n9015 );
  nand     g09155 ( new_n9532 , new_n9530 , new_n9531 );
  nand     g09156 ( new_n9533 , pi099 , pi224 );
  xor      g09157 ( new_n9534 , new_n9532 , new_n9533 );
  nand     g09158 ( new_n9535 , pi021 , pi219 );
  nand     g09159 ( new_n9536 , pi137 , pi217 );
  xor      g09160 ( new_n9537 , new_n9535 , new_n9536 );
  or       g09161 ( new_n9538 , new_n9057 , new_n9066 );
  nand     g09162 ( new_n9539 , new_n9067 , new_n9071 );
  nand     g09163 ( new_n9540 , new_n9538 , new_n9539 );
  xor      g09164 ( new_n9541 , new_n9537 , new_n9540 );
  xor      g09165 ( new_n9542 , new_n9534 , new_n9541 );
  xor      g09166 ( new_n9543 , new_n9529 , new_n9542 );
  xor      g09167 ( new_n9544 , new_n9528 , new_n9543 );
  xor      g09168 ( new_n9545 , new_n9525 , new_n9544 );
  xor      g09169 ( new_n9546 , new_n9522 , new_n9545 );
  xor      g09170 ( new_n9547 , new_n9509 , new_n9546 );
  xor      g09171 ( new_n9548 , new_n9471 , new_n9547 );
  xor      g09172 ( new_n9549 , new_n9466 , new_n9548 );
  xor      g09173 ( new_n9550 , new_n9373 , new_n9549 );
  xor      g09174 ( po051 , new_n9360 , new_n9550 );
  xor      g09175 ( po052 , new_n3213 , new_n3218 );
  xor      g09176 ( po053 , new_n3492 , new_n3497 );
  xor      g09177 ( po054 , new_n393 , new_n890 );
  xor      g09178 ( po055 , new_n7639 , new_n7640 );
  xor      g09179 ( po056 , new_n4269 , new_n4270 );
  xor      g09180 ( po057 , new_n1855 , new_n1857 );
  xor      g09181 ( po058 , new_n4247 , new_n4248 );
  xnor     g09182 ( po059 , new_n5482 , new_n5483 );
  nand     g09183 ( new_n9560 , new_n2598 , new_n2600 );
  xor      g09184 ( po060 , new_n2595 , new_n9560 );
  xor      g09185 ( po061 , new_n2589 , new_n2591 );
  nor      g09186 ( new_n9563 , new_n8820 , new_n8823 );
  nand g09187 ( new_n9564 , new_n8824 , new_n8824 );
  nor      g09188 ( new_n9565 , new_n9564 , new_n8835 );
  nor      g09189 ( new_n9566 , new_n9563 , new_n9565 );
  nand     g09190 ( new_n9567 , new_n8832 , new_n8833 );
  nand     g09191 ( new_n9568 , new_n8829 , new_n8834 );
  nand     g09192 ( new_n9569 , new_n9567 , new_n9568 );
  nand     g09193 ( new_n9570 , pi077 , pi081 );
  nand     g09194 ( new_n9571 , pi052 , pi106 );
  and      g09195 ( new_n9572 , new_n9570 , new_n9571 );
  nand     g09196 ( new_n9573 , pi077 , pi106 );
  nor      g09197 ( new_n9574 , new_n8833 , new_n9573 );
  nor      g09198 ( new_n9575 , new_n9572 , new_n9574 );
  nand g09199 ( new_n9576 , new_n9575 , new_n9575 );
  nand     g09200 ( new_n9577 , pi133 , pi227 );
  nand     g09201 ( new_n9578 , new_n8826 , new_n8827 );
  nand     g09202 ( new_n9579 , new_n8825 , new_n8828 );
  nand     g09203 ( new_n9580 , new_n9578 , new_n9579 );
  nand     g09204 ( new_n9581 , pi100 , pi189 );
  nand     g09205 ( new_n9582 , pi064 , pi217 );
  nand     g09206 ( new_n9583 , new_n9581 , new_n9582 );
  nand     g09207 ( new_n9584 , pi064 , pi100 );
  or       g09208 ( new_n9585 , new_n8827 , new_n9584 );
  nand     g09209 ( new_n9586 , new_n9583 , new_n9585 );
  xor      g09210 ( new_n9587 , new_n9580 , new_n9586 );
  xor      g09211 ( new_n9588 , new_n9577 , new_n9587 );
  xor      g09212 ( new_n9589 , new_n9576 , new_n9588 );
  xor      g09213 ( new_n9590 , new_n9569 , new_n9589 );
  xor      g09214 ( new_n9591 , new_n9566 , new_n9590 );
  nor      g09215 ( new_n9592 , new_n8819 , new_n8836 );
  nand     g09216 ( new_n9593 , pi131 , pi233 );
  xor      g09217 ( new_n9594 , new_n9592 , new_n9593 );
  xor      g09218 ( new_n9595 , new_n9591 , new_n9594 );
  nand g09219 ( new_n9596 , new_n8817 , new_n8817 );
  nor      g09220 ( new_n9597 , new_n9596 , new_n8837 );
  nand g09221 ( new_n9598 , new_n8842 , new_n8842 );
  nor      g09222 ( new_n9599 , new_n8838 , new_n9598 );
  nor      g09223 ( new_n9600 , new_n9597 , new_n9599 );
  nand g09224 ( new_n9601 , new_n9600 , new_n9600 );
  nor      g09225 ( new_n9602 , new_n9595 , new_n9601 );
  nor      g09226 ( new_n9603 , new_n8795 , new_n8815 );
  nor      g09227 ( new_n9604 , new_n8792 , new_n8816 );
  nor      g09228 ( new_n9605 , new_n9603 , new_n9604 );
  nand g09229 ( new_n9606 , new_n8814 , new_n8814 );
  nor      g09230 ( new_n9607 , new_n8796 , new_n9606 );
  nand     g09231 ( new_n9608 , pi168 , pi174 );
  nor      g09232 ( new_n9609 , new_n8797 , new_n8800 );
  and      g09233 ( new_n9610 , new_n8801 , new_n8813 );
  nor      g09234 ( new_n9611 , new_n9609 , new_n9610 );
  nand     g09235 ( new_n9612 , pi139 , pi176 );
  nand     g09236 ( new_n9613 , pi040 , pi208 );
  nand     g09237 ( new_n9614 , new_n9612 , new_n9613 );
  nand     g09238 ( new_n9615 , pi040 , pi139 );
  nor      g09239 ( new_n9616 , new_n8807 , new_n9615 );
  nand g09240 ( new_n9617 , new_n9616 , new_n9616 );
  nand     g09241 ( new_n9618 , new_n9614 , new_n9617 );
  nand     g09242 ( new_n9619 , new_n8807 , new_n8810 );
  nand     g09243 ( new_n9620 , new_n8806 , new_n8811 );
  nand     g09244 ( new_n9621 , new_n9619 , new_n9620 );
  nand     g09245 ( new_n9622 , pi035 , pi125 );
  nand     g09246 ( new_n9623 , new_n8803 , new_n8804 );
  nand     g09247 ( new_n9624 , new_n8802 , new_n8805 );
  nand     g09248 ( new_n9625 , new_n9623 , new_n9624 );
  nand     g09249 ( new_n9626 , pi204 , pi249 );
  nand     g09250 ( new_n9627 , pi015 , pi222 );
  nand     g09251 ( new_n9628 , new_n9626 , new_n9627 );
  nand     g09252 ( new_n9629 , pi204 , pi222 );
  or       g09253 ( new_n9630 , new_n8802 , new_n9629 );
  nand     g09254 ( new_n9631 , new_n9628 , new_n9630 );
  xor      g09255 ( new_n9632 , new_n9625 , new_n9631 );
  xor      g09256 ( new_n9633 , new_n9622 , new_n9632 );
  xor      g09257 ( new_n9634 , new_n9621 , new_n9633 );
  xor      g09258 ( new_n9635 , new_n9618 , new_n9634 );
  xnor     g09259 ( new_n9636 , new_n9611 , new_n9635 );
  xor      g09260 ( new_n9637 , new_n9608 , new_n9636 );
  xnor     g09261 ( new_n9638 , new_n9607 , new_n9637 );
  xor      g09262 ( new_n9639 , new_n9605 , new_n9638 );
  nand g09263 ( new_n9640 , new_n8787 , new_n8787 );
  nand     g09264 ( new_n9641 , new_n9640 , new_n8790 );
  or       g09265 ( new_n9642 , new_n8767 , new_n8791 );
  nand     g09266 ( new_n9643 , new_n9641 , new_n9642 );
  nand     g09267 ( new_n9644 , new_n8749 , new_n8766 );
  nand     g09268 ( new_n9645 , pi005 , pi236 );
  nand     g09269 ( new_n9646 , new_n8760 , new_n8763 );
  nand     g09270 ( new_n9647 , new_n8759 , new_n8764 );
  nand     g09271 ( new_n9648 , new_n9646 , new_n9647 );
  nand     g09272 ( new_n9649 , pi121 , pi161 );
  nand     g09273 ( new_n9650 , pi231 , pi241 );
  and      g09274 ( new_n9651 , new_n9649 , new_n9650 );
  nand     g09275 ( new_n9652 , pi161 , pi231 );
  nor      g09276 ( new_n9653 , new_n8760 , new_n9652 );
  nor      g09277 ( new_n9654 , new_n9651 , new_n9653 );
  nand     g09278 ( new_n9655 , new_n8756 , new_n8757 );
  nand     g09279 ( new_n9656 , new_n8755 , new_n8758 );
  nand     g09280 ( new_n9657 , new_n9655 , new_n9656 );
  nand     g09281 ( new_n9658 , pi141 , pi252 );
  nand     g09282 ( new_n9659 , pi090 , pi140 );
  nand     g09283 ( new_n9660 , pi047 , pi242 );
  nand     g09284 ( new_n9661 , new_n9659 , new_n9660 );
  nand     g09285 ( new_n9662 , pi047 , pi140 );
  or       g09286 ( new_n9663 , new_n8756 , new_n9662 );
  nand     g09287 ( new_n9664 , new_n9661 , new_n9663 );
  xor      g09288 ( new_n9665 , new_n9658 , new_n9664 );
  xor      g09289 ( new_n9666 , new_n9657 , new_n9665 );
  xor      g09290 ( new_n9667 , new_n9654 , new_n9666 );
  xor      g09291 ( new_n9668 , new_n9648 , new_n9667 );
  nor      g09292 ( new_n9669 , new_n8750 , new_n8753 );
  and      g09293 ( new_n9670 , new_n8754 , new_n8765 );
  nor      g09294 ( new_n9671 , new_n9669 , new_n9670 );
  xor      g09295 ( new_n9672 , new_n9668 , new_n9671 );
  xor      g09296 ( new_n9673 , new_n9645 , new_n9672 );
  xor      g09297 ( new_n9674 , new_n9644 , new_n9673 );
  nand     g09298 ( new_n9675 , new_n8769 , new_n8786 );
  nand     g09299 ( new_n9676 , pi127 , pi213 );
  xor      g09300 ( new_n9677 , new_n9675 , new_n9676 );
  nand     g09301 ( new_n9678 , pi104 , pi224 );
  nand     g09302 ( new_n9679 , pi212 , pi255 );
  nand     g09303 ( new_n9680 , new_n9678 , new_n9679 );
  nand     g09304 ( new_n9681 , pi104 , pi255 );
  or       g09305 ( new_n9682 , new_n8780 , new_n9681 );
  nand     g09306 ( new_n9683 , new_n9680 , new_n9682 );
  nand     g09307 ( new_n9684 , pi013 , pi024 );
  nand     g09308 ( new_n9685 , new_n8776 , new_n8777 );
  nand     g09309 ( new_n9686 , new_n8775 , new_n8778 );
  nand     g09310 ( new_n9687 , new_n9685 , new_n9686 );
  nand     g09311 ( new_n9688 , pi111 , pi112 );
  nand     g09312 ( new_n9689 , pi105 , pi210 );
  nand     g09313 ( new_n9690 , new_n9688 , new_n9689 );
  nand     g09314 ( new_n9691 , pi105 , pi111 );
  nor      g09315 ( new_n9692 , new_n8777 , new_n9691 );
  nand g09316 ( new_n9693 , new_n9692 , new_n9692 );
  nand     g09317 ( new_n9694 , new_n9690 , new_n9693 );
  xor      g09318 ( new_n9695 , new_n9687 , new_n9694 );
  xor      g09319 ( new_n9696 , new_n9684 , new_n9695 );
  xor      g09320 ( new_n9697 , new_n9683 , new_n9696 );
  nand     g09321 ( new_n9698 , new_n8780 , new_n8783 );
  nand     g09322 ( new_n9699 , new_n8779 , new_n8784 );
  nand     g09323 ( new_n9700 , new_n9698 , new_n9699 );
  xor      g09324 ( new_n9701 , new_n9697 , new_n9700 );
  nor      g09325 ( new_n9702 , new_n8770 , new_n8773 );
  nand     g09326 ( new_n9703 , new_n8774 , new_n8785 );
  nand g09327 ( new_n9704 , new_n9703 , new_n9703 );
  nor      g09328 ( new_n9705 , new_n9702 , new_n9704 );
  xnor     g09329 ( new_n9706 , new_n9701 , new_n9705 );
  xor      g09330 ( new_n9707 , new_n9677 , new_n9706 );
  xor      g09331 ( new_n9708 , new_n9674 , new_n9707 );
  xor      g09332 ( new_n9709 , new_n9643 , new_n9708 );
  xor      g09333 ( new_n9710 , new_n9639 , new_n9709 );
  xor      g09334 ( new_n9711 , new_n9595 , new_n9600 );
  nor      g09335 ( new_n9712 , new_n9710 , new_n9711 );
  nor      g09336 ( new_n9713 , new_n9602 , new_n9712 );
  nand     g09337 ( new_n9714 , new_n9674 , new_n9707 );
  nand     g09338 ( new_n9715 , new_n9643 , new_n9708 );
  and      g09339 ( new_n9716 , new_n9714 , new_n9715 );
  nor      g09340 ( new_n9717 , new_n9645 , new_n9672 );
  nand g09341 ( new_n9718 , new_n9673 , new_n9673 );
  nor      g09342 ( new_n9719 , new_n9644 , new_n9718 );
  nor      g09343 ( new_n9720 , new_n9717 , new_n9719 );
  nand g09344 ( new_n9721 , new_n9668 , new_n9668 );
  nor      g09345 ( new_n9722 , new_n9721 , new_n9671 );
  nor      g09346 ( new_n9723 , new_n9648 , new_n9667 );
  and      g09347 ( new_n9724 , new_n9653 , new_n9723 );
  nand g09348 ( new_n9725 , new_n9666 , new_n9666 );
  nand     g09349 ( new_n9726 , new_n9654 , new_n9725 );
  nand g09350 ( new_n9727 , new_n9726 , new_n9726 );
  nor      g09351 ( new_n9728 , new_n9653 , new_n9727 );
  nand g09352 ( new_n9729 , new_n9728 , new_n9728 );
  nor      g09353 ( new_n9730 , new_n9723 , new_n9729 );
  or       g09354 ( new_n9731 , new_n9724 , new_n9730 );
  nand     g09355 ( new_n9732 , pi121 , pi141 );
  xor      g09356 ( new_n9733 , new_n9663 , new_n9732 );
  nand     g09357 ( new_n9734 , pi018 , pi242 );
  nand     g09358 ( new_n9735 , pi090 , pi252 );
  xor      g09359 ( new_n9736 , new_n9734 , new_n9735 );
  xnor     g09360 ( new_n9737 , new_n9662 , new_n9736 );
  xor      g09361 ( new_n9738 , new_n9733 , new_n9737 );
  nand     g09362 ( new_n9739 , new_n9658 , new_n9664 );
  nand     g09363 ( new_n9740 , new_n9657 , new_n9665 );
  nand     g09364 ( new_n9741 , new_n9739 , new_n9740 );
  nand     g09365 ( new_n9742 , pi021 , pi236 );
  nand     g09366 ( new_n9743 , pi005 , pi241 );
  xor      g09367 ( new_n9744 , new_n9742 , new_n9743 );
  xor      g09368 ( new_n9745 , new_n9652 , new_n9744 );
  xor      g09369 ( new_n9746 , new_n9741 , new_n9745 );
  xor      g09370 ( new_n9747 , new_n9738 , new_n9746 );
  xor      g09371 ( new_n9748 , new_n9731 , new_n9747 );
  xor      g09372 ( new_n9749 , new_n9722 , new_n9748 );
  xor      g09373 ( new_n9750 , new_n9720 , new_n9749 );
  nand     g09374 ( new_n9751 , new_n9675 , new_n9676 );
  nand g09375 ( new_n9752 , new_n9751 , new_n9751 );
  and      g09376 ( new_n9753 , new_n9677 , new_n9706 );
  nor      g09377 ( new_n9754 , new_n9752 , new_n9753 );
  nor      g09378 ( new_n9755 , new_n9701 , new_n9705 );
  nand     g09379 ( new_n9756 , new_n9683 , new_n9696 );
  nand     g09380 ( new_n9757 , new_n9697 , new_n9700 );
  nand     g09381 ( new_n9758 , new_n9756 , new_n9757 );
  xor      g09382 ( new_n9759 , new_n9682 , new_n9758 );
  nand     g09383 ( new_n9760 , pi183 , pi210 );
  nand     g09384 ( new_n9761 , pi024 , pi112 );
  xor      g09385 ( new_n9762 , new_n9760 , new_n9761 );
  xor      g09386 ( new_n9763 , new_n9691 , new_n9762 );
  nand     g09387 ( new_n9764 , pi013 , pi224 );
  xor      g09388 ( new_n9765 , new_n9692 , new_n9764 );
  xor      g09389 ( new_n9766 , new_n9763 , new_n9765 );
  nand     g09390 ( new_n9767 , new_n9687 , new_n9694 );
  nand     g09391 ( new_n9768 , new_n9684 , new_n9695 );
  nand     g09392 ( new_n9769 , new_n9767 , new_n9768 );
  nand     g09393 ( new_n9770 , pi127 , pi212 );
  nand     g09394 ( new_n9771 , pi213 , pi232 );
  xor      g09395 ( new_n9772 , new_n9770 , new_n9771 );
  xnor     g09396 ( new_n9773 , new_n9681 , new_n9772 );
  xor      g09397 ( new_n9774 , new_n9769 , new_n9773 );
  xor      g09398 ( new_n9775 , new_n9766 , new_n9774 );
  xor      g09399 ( new_n9776 , new_n9759 , new_n9775 );
  nand g09400 ( new_n9777 , new_n9776 , new_n9776 );
  and      g09401 ( new_n9778 , new_n9755 , new_n9777 );
  nor      g09402 ( new_n9779 , new_n9755 , new_n9777 );
  nor      g09403 ( new_n9780 , new_n9778 , new_n9779 );
  xor      g09404 ( new_n9781 , new_n9754 , new_n9780 );
  xor      g09405 ( new_n9782 , new_n9750 , new_n9781 );
  xor      g09406 ( new_n9783 , new_n9716 , new_n9782 );
  nand     g09407 ( new_n9784 , new_n9605 , new_n9638 );
  nand     g09408 ( new_n9785 , new_n9639 , new_n9709 );
  and      g09409 ( new_n9786 , new_n9784 , new_n9785 );
  nor      g09410 ( new_n9787 , new_n9608 , new_n9636 );
  nand     g09411 ( new_n9788 , new_n9607 , new_n9637 );
  nand g09412 ( new_n9789 , new_n9788 , new_n9788 );
  nor      g09413 ( new_n9790 , new_n9787 , new_n9789 );
  nor      g09414 ( new_n9791 , new_n9611 , new_n9635 );
  nand     g09415 ( new_n9792 , pi174 , pi208 );
  nand     g09416 ( new_n9793 , pi157 , pi168 );
  xor      g09417 ( new_n9794 , new_n9792 , new_n9793 );
  xnor     g09418 ( new_n9795 , new_n9615 , new_n9794 );
  nand     g09419 ( new_n9796 , new_n9625 , new_n9631 );
  nand     g09420 ( new_n9797 , new_n9622 , new_n9632 );
  nand     g09421 ( new_n9798 , new_n9796 , new_n9797 );
  xor      g09422 ( new_n9799 , new_n9795 , new_n9798 );
  nand     g09423 ( new_n9800 , pi035 , pi176 );
  xor      g09424 ( new_n9801 , new_n9630 , new_n9800 );
  nand     g09425 ( new_n9802 , pi146 , pi249 );
  nand     g09426 ( new_n9803 , pi015 , pi125 );
  xor      g09427 ( new_n9804 , new_n9802 , new_n9803 );
  xor      g09428 ( new_n9805 , new_n9629 , new_n9804 );
  xor      g09429 ( new_n9806 , new_n9801 , new_n9805 );
  xor      g09430 ( new_n9807 , new_n9799 , new_n9806 );
  nor      g09431 ( new_n9808 , new_n9621 , new_n9633 );
  xor      g09432 ( new_n9809 , new_n9617 , new_n9808 );
  nand     g09433 ( new_n9810 , new_n9614 , new_n9634 );
  nand     g09434 ( new_n9811 , new_n9809 , new_n9810 );
  xor      g09435 ( new_n9812 , new_n9807 , new_n9811 );
  xor      g09436 ( new_n9813 , new_n9791 , new_n9812 );
  nand g09437 ( new_n9814 , new_n9813 , new_n9813 );
  xor      g09438 ( new_n9815 , new_n9790 , new_n9814 );
  xnor     g09439 ( new_n9816 , new_n9786 , new_n9815 );
  xor      g09440 ( new_n9817 , new_n9783 , new_n9816 );
  nor      g09441 ( new_n9818 , new_n9566 , new_n9590 );
  nand g09442 ( new_n9819 , new_n9593 , new_n9593 );
  nor      g09443 ( new_n9820 , new_n9592 , new_n9819 );
  nand g09444 ( new_n9821 , new_n9820 , new_n9820 );
  or       g09445 ( new_n9822 , new_n9591 , new_n9594 );
  nand     g09446 ( new_n9823 , new_n9821 , new_n9822 );
  nand     g09447 ( new_n9824 , pi131 , pi187 );
  nand     g09448 ( new_n9825 , pi052 , pi233 );
  xor      g09449 ( new_n9826 , new_n9824 , new_n9825 );
  xnor     g09450 ( new_n9827 , new_n9573 , new_n9826 );
  nand     g09451 ( new_n9828 , new_n9580 , new_n9586 );
  nand     g09452 ( new_n9829 , new_n9577 , new_n9587 );
  nand     g09453 ( new_n9830 , new_n9828 , new_n9829 );
  nand g09454 ( new_n9831 , new_n9830 , new_n9830 );
  xor      g09455 ( new_n9832 , new_n9827 , new_n9831 );
  nand     g09456 ( new_n9833 , pi081 , pi133 );
  xor      g09457 ( new_n9834 , new_n9585 , new_n9833 );
  nand     g09458 ( new_n9835 , pi189 , pi227 );
  nand     g09459 ( new_n9836 , pi084 , pi217 );
  xor      g09460 ( new_n9837 , new_n9835 , new_n9836 );
  xor      g09461 ( new_n9838 , new_n9584 , new_n9837 );
  xor      g09462 ( new_n9839 , new_n9834 , new_n9838 );
  xor      g09463 ( new_n9840 , new_n9832 , new_n9839 );
  nand     g09464 ( new_n9841 , new_n9576 , new_n9588 );
  nand     g09465 ( new_n9842 , new_n9569 , new_n9589 );
  nand     g09466 ( new_n9843 , new_n9841 , new_n9842 );
  xor      g09467 ( new_n9844 , new_n9574 , new_n9843 );
  xor      g09468 ( new_n9845 , new_n9840 , new_n9844 );
  nand g09469 ( new_n9846 , new_n9845 , new_n9845 );
  xor      g09470 ( new_n9847 , new_n9823 , new_n9846 );
  xnor     g09471 ( new_n9848 , new_n9818 , new_n9847 );
  xnor     g09472 ( new_n9849 , new_n9817 , new_n9848 );
  xor      g09473 ( po062 , new_n9713 , new_n9849 );
  xor      g09474 ( po063 , new_n9425 , new_n9426 );
  nor      g09475 ( new_n9852 , new_n3015 , new_n3019 );
  nor      g09476 ( new_n9853 , new_n3012 , new_n3020 );
  nor      g09477 ( new_n9854 , new_n9852 , new_n9853 );
  nand     g09478 ( new_n9855 , pi023 , pi073 );
  xor      g09479 ( new_n9856 , new_n9854 , new_n9855 );
  nand     g09480 ( new_n9857 , new_n2995 , new_n3062 );
  nand     g09481 ( new_n9858 , new_n2961 , new_n3063 );
  nand     g09482 ( new_n9859 , new_n9857 , new_n9858 );
  nand g09483 ( new_n9860 , new_n3036 , new_n3036 );
  nor      g09484 ( new_n9861 , new_n9860 , new_n3058 );
  nor      g09485 ( new_n9862 , new_n3035 , new_n3059 );
  or       g09486 ( new_n9863 , new_n9861 , new_n9862 );
  nor      g09487 ( new_n9864 , new_n2986 , new_n2990 );
  and      g09488 ( new_n9865 , new_n2983 , new_n2991 );
  nor      g09489 ( new_n9866 , new_n9864 , new_n9865 );
  xor      g09490 ( new_n9867 , new_n9863 , new_n9866 );
  xor      g09491 ( new_n9868 , new_n9859 , new_n9867 );
  nand     g09492 ( new_n9869 , pi060 , pi185 );
  or       g09493 ( new_n9870 , new_n3005 , new_n3028 );
  nand g09494 ( new_n9871 , new_n3002 , new_n3002 );
  nand     g09495 ( new_n9872 , new_n9871 , new_n3029 );
  nand     g09496 ( new_n9873 , new_n9870 , new_n9872 );
  xor      g09497 ( new_n9874 , new_n9869 , new_n9873 );
  nand     g09498 ( new_n9875 , pi078 , pi138 );
  nand     g09499 ( new_n9876 , new_n3079 , new_n3096 );
  nand     g09500 ( new_n9877 , new_n3074 , new_n3097 );
  nand     g09501 ( new_n9878 , new_n9876 , new_n9877 );
  xor      g09502 ( new_n9879 , new_n9875 , new_n9878 );
  nand     g09503 ( new_n9880 , new_n2979 , new_n2980 );
  nand     g09504 ( new_n9881 , new_n2899 , new_n2981 );
  nand     g09505 ( new_n9882 , new_n9880 , new_n9881 );
  xor      g09506 ( new_n9883 , new_n9879 , new_n9882 );
  xor      g09507 ( new_n9884 , new_n9874 , new_n9883 );
  xor      g09508 ( new_n9885 , new_n9868 , new_n9884 );
  xor      g09509 ( new_n9886 , new_n9856 , new_n9885 );
  nand     g09510 ( new_n9887 , pi182 , pi197 );
  nand     g09511 ( new_n9888 , new_n3070 , new_n3071 );
  nand     g09512 ( new_n9889 , new_n3066 , new_n3072 );
  nand     g09513 ( new_n9890 , new_n9888 , new_n9889 );
  xor      g09514 ( new_n9891 , new_n9887 , new_n9890 );
  xor      g09515 ( new_n9892 , new_n9886 , new_n9891 );
  or       g09516 ( new_n9893 , new_n3098 , new_n3126 );
  nand     g09517 ( new_n9894 , new_n3123 , new_n9893 );
  nand     g09518 ( new_n9895 , new_n2785 , new_n3017 );
  nand     g09519 ( new_n9896 , new_n3016 , new_n3018 );
  nand     g09520 ( new_n9897 , new_n9895 , new_n9896 );
  xnor     g09521 ( new_n9898 , new_n9894 , new_n9897 );
  or       g09522 ( new_n9899 , new_n3021 , new_n3027 );
  nand     g09523 ( new_n9900 , new_n3026 , new_n9899 );
  nand     g09524 ( new_n9901 , pi094 , pi254 );
  xnor     g09525 ( new_n9902 , new_n9900 , new_n9901 );
  nand     g09526 ( new_n9903 , pi123 , pi130 );
  nand     g09527 ( new_n9904 , new_n3051 , new_n3052 );
  nand     g09528 ( new_n9905 , new_n2830 , new_n3053 );
  nand     g09529 ( new_n9906 , new_n9904 , new_n9905 );
  xor      g09530 ( new_n9907 , new_n9903 , new_n9906 );
  nor      g09531 ( new_n9908 , new_n3043 , new_n3047 );
  nor      g09532 ( new_n9909 , new_n3048 , new_n3055 );
  nor      g09533 ( new_n9910 , new_n9908 , new_n9909 );
  nand     g09534 ( new_n9911 , new_n3008 , new_n3009 );
  nand     g09535 ( new_n9912 , new_n2792 , new_n3010 );
  nand     g09536 ( new_n9913 , new_n9911 , new_n9912 );
  nand     g09537 ( new_n9914 , pi022 , pi142 );
  xor      g09538 ( new_n9915 , new_n9913 , new_n9914 );
  xor      g09539 ( new_n9916 , new_n9910 , new_n9915 );
  xor      g09540 ( new_n9917 , new_n9907 , new_n9916 );
  xor      g09541 ( new_n9918 , new_n9902 , new_n9917 );
  xor      g09542 ( new_n9919 , new_n9898 , new_n9918 );
  nand     g09543 ( new_n9920 , pi062 , pi251 );
  nand     g09544 ( new_n9921 , new_n3076 , new_n3077 );
  nand     g09545 ( new_n9922 , new_n3075 , new_n3078 );
  nand     g09546 ( new_n9923 , new_n9921 , new_n9922 );
  nand     g09547 ( new_n9924 , pi160 , pi220 );
  xor      g09548 ( new_n9925 , new_n9923 , new_n9924 );
  xor      g09549 ( new_n9926 , new_n9920 , new_n9925 );
  nand     g09550 ( new_n9927 , pi020 , pi030 );
  nor      g09551 ( new_n9928 , new_n2968 , new_n2993 );
  nor      g09552 ( new_n9929 , new_n2966 , new_n2994 );
  nor      g09553 ( new_n9930 , new_n9928 , new_n9929 );
  xor      g09554 ( new_n9931 , new_n9927 , new_n9930 );
  nand     g09555 ( new_n9932 , pi079 , pi120 );
  xor      g09556 ( new_n9933 , new_n9931 , new_n9932 );
  xor      g09557 ( new_n9934 , new_n9926 , new_n9933 );
  nand     g09558 ( new_n9935 , pi001 , pi095 );
  nand     g09559 ( new_n9936 , new_n3044 , new_n3045 );
  nand     g09560 ( new_n9937 , new_n2823 , new_n3046 );
  nand     g09561 ( new_n9938 , new_n9936 , new_n9937 );
  nor      g09562 ( new_n9939 , new_n2832 , new_n3049 );
  nor      g09563 ( new_n9940 , new_n3050 , new_n3054 );
  nor      g09564 ( new_n9941 , new_n9939 , new_n9940 );
  xor      g09565 ( new_n9942 , new_n9938 , new_n9941 );
  xor      g09566 ( new_n9943 , new_n9935 , new_n9942 );
  xor      g09567 ( new_n9944 , new_n9934 , new_n9943 );
  xor      g09568 ( new_n9945 , new_n9919 , new_n9944 );
  nand     g09569 ( new_n9946 , pi041 , pi165 );
  nand     g09570 ( new_n9947 , pi071 , pi215 );
  nand     g09571 ( new_n9948 , pi059 , pi158 );
  xor      g09572 ( new_n9949 , new_n9947 , new_n9948 );
  xor      g09573 ( new_n9950 , new_n9946 , new_n9949 );
  xor      g09574 ( new_n9951 , new_n9945 , new_n9950 );
  nand     g09575 ( new_n9952 , new_n2987 , new_n2988 );
  nand     g09576 ( new_n9953 , new_n2889 , new_n2989 );
  nand     g09577 ( new_n9954 , new_n9952 , new_n9953 );
  nand     g09578 ( new_n9955 , pi003 , pi099 );
  xor      g09579 ( new_n9956 , new_n9954 , new_n9955 );
  nand     g09580 ( new_n9957 , pi209 , pi219 );
  nand     g09581 ( new_n9958 , pi089 , pi135 );
  nand g09582 ( new_n9959 , new_n3150 , new_n3150 );
  nor      g09583 ( new_n9960 , new_n3127 , new_n9959 );
  nor      g09584 ( new_n9961 , new_n3151 , new_n3171 );
  nor      g09585 ( new_n9962 , new_n9960 , new_n9961 );
  xor      g09586 ( new_n9963 , new_n9958 , new_n9962 );
  xor      g09587 ( new_n9964 , new_n9957 , new_n9963 );
  nand     g09588 ( new_n9965 , pi198 , pi216 );
  nor      g09589 ( new_n9966 , new_n2901 , new_n2977 );
  nor      g09590 ( new_n9967 , new_n2978 , new_n2982 );
  nor      g09591 ( new_n9968 , new_n9966 , new_n9967 );
  xor      g09592 ( new_n9969 , new_n9965 , new_n9968 );
  xor      g09593 ( new_n9970 , new_n9964 , new_n9969 );
  nor      g09594 ( new_n9971 , new_n3030 , new_n3060 );
  nor      g09595 ( new_n9972 , new_n2999 , new_n3061 );
  nor      g09596 ( new_n9973 , new_n9971 , new_n9972 );
  nor      g09597 ( new_n9974 , new_n3086 , new_n3068 );
  nor      g09598 ( new_n9975 , new_n3069 , new_n3073 );
  nor      g09599 ( new_n9976 , new_n9974 , new_n9975 );
  nand     g09600 ( new_n9977 , pi137 , pi190 );
  nand     g09601 ( new_n9978 , pi076 , pi172 );
  xor      g09602 ( new_n9979 , new_n9977 , new_n9978 );
  xor      g09603 ( new_n9980 , new_n9976 , new_n9979 );
  xor      g09604 ( new_n9981 , new_n9973 , new_n9980 );
  nand     g09605 ( new_n9982 , new_n2825 , new_n3039 );
  nand     g09606 ( new_n9983 , new_n3040 , new_n3057 );
  nand     g09607 ( new_n9984 , new_n9982 , new_n9983 );
  nand     g09608 ( new_n9985 , pi004 , pi155 );
  xor      g09609 ( new_n9986 , new_n9984 , new_n9985 );
  nand     g09610 ( new_n9987 , pi092 , pi177 );
  nand     g09611 ( new_n9988 , pi065 , pi192 );
  nand     g09612 ( new_n9989 , pi067 , pi101 );
  xor      g09613 ( new_n9990 , new_n9988 , new_n9989 );
  nand     g09614 ( new_n9991 , pi225 , pi229 );
  xor      g09615 ( new_n9992 , new_n9990 , new_n9991 );
  xor      g09616 ( new_n9993 , new_n9987 , new_n9992 );
  xor      g09617 ( new_n9994 , new_n9986 , new_n9993 );
  xor      g09618 ( new_n9995 , new_n9981 , new_n9994 );
  nand     g09619 ( new_n9996 , pi006 , pi102 );
  nand     g09620 ( new_n9997 , pi086 , pi170 );
  xor      g09621 ( new_n9998 , new_n9996 , new_n9997 );
  nor      g09622 ( new_n9999 , new_n2976 , new_n2992 );
  nor      g09623 ( new_n10000 , new_n2975 , new_n9999 );
  nand     g09624 ( new_n10001 , pi053 , pi223 );
  xor      g09625 ( new_n10002 , new_n10000 , new_n10001 );
  xor      g09626 ( new_n10003 , new_n9998 , new_n10002 );
  xor      g09627 ( new_n10004 , new_n9995 , new_n10003 );
  xor      g09628 ( new_n10005 , new_n9970 , new_n10004 );
  nand     g09629 ( new_n10006 , pi122 , pi154 );
  nand     g09630 ( new_n10007 , pi124 , pi169 );
  xor      g09631 ( new_n10008 , new_n10006 , new_n10007 );
  xor      g09632 ( new_n10009 , new_n10005 , new_n10008 );
  xor      g09633 ( new_n10010 , new_n9956 , new_n10009 );
  xor      g09634 ( new_n10011 , new_n9951 , new_n10010 );
  nand     g09635 ( new_n10012 , new_n3064 , new_n3172 );
  nand     g09636 ( new_n10013 , new_n3173 , new_n3211 );
  nand     g09637 ( new_n10014 , new_n10012 , new_n10013 );
  nor      g09638 ( new_n10015 , new_n2794 , new_n3006 );
  nor      g09639 ( new_n10016 , new_n3007 , new_n3011 );
  nor      g09640 ( new_n10017 , new_n10015 , new_n10016 );
  nand     g09641 ( new_n10018 , pi087 , pi153 );
  xor      g09642 ( new_n10019 , new_n10017 , new_n10018 );
  xor      g09643 ( new_n10020 , new_n10014 , new_n10019 );
  xor      g09644 ( new_n10021 , new_n10011 , new_n10020 );
  xor      g09645 ( po064 , new_n9892 , new_n10021 );
  xnor     g09646 ( po065 , new_n9436 , new_n9437 );
  xnor     g09647 ( po066 , new_n3192 , new_n3193 );
  xor      g09648 ( po067 , new_n5103 , new_n5104 );
  xor      g09649 ( po068 , new_n7202 , new_n7203 );
  xnor     g09650 ( po069 , new_n4252 , new_n4259 );
  xnor     g09651 ( po070 , new_n1132 , new_n1171 );
  xor      g09652 ( po071 , new_n9442 , new_n9443 );
  nand     g09653 ( new_n10030 , pi068 , pi131 );
  nand     g09654 ( new_n10031 , pi036 , pi052 );
  nand     g09655 ( new_n10032 , new_n10030 , new_n10031 );
  xor      g09656 ( new_n10033 , new_n10030 , new_n10031 );
  nand     g09657 ( new_n10034 , new_n6625 , new_n10033 );
  nand     g09658 ( new_n10035 , new_n10032 , new_n10034 );
  or       g09659 ( new_n10036 , new_n6531 , new_n6534 );
  nand     g09660 ( new_n10037 , pi015 , pi179 );
  nand     g09661 ( new_n10038 , pi146 , pi162 );
  xor      g09662 ( new_n10039 , new_n10037 , new_n10038 );
  xnor     g09663 ( new_n10040 , new_n6523 , new_n10039 );
  nand     g09664 ( new_n10041 , pi035 , pi048 );
  xor      g09665 ( new_n10042 , new_n6524 , new_n10041 );
  xor      g09666 ( new_n10043 , new_n10040 , new_n10042 );
  nand     g09667 ( new_n10044 , new_n6519 , new_n6526 );
  nand     g09668 ( new_n10045 , new_n6518 , new_n6527 );
  nand     g09669 ( new_n10046 , new_n10044 , new_n10045 );
  nand     g09670 ( new_n10047 , pi168 , pi193 );
  nand     g09671 ( new_n10048 , pi208 , pi238 );
  xor      g09672 ( new_n10049 , new_n10047 , new_n10048 );
  xor      g09673 ( new_n10050 , new_n6513 , new_n10049 );
  xnor     g09674 ( new_n10051 , new_n10046 , new_n10050 );
  xor      g09675 ( new_n10052 , new_n10043 , new_n10051 );
  nor      g09676 ( new_n10053 , new_n6509 , new_n6529 );
  nand     g09677 ( new_n10054 , new_n6514 , new_n10053 );
  nand g09678 ( new_n10055 , new_n10053 , new_n10053 );
  nand g09679 ( new_n10056 , new_n6528 , new_n6528 );
  nand     g09680 ( new_n10057 , new_n6515 , new_n10056 );
  nand g09681 ( new_n10058 , new_n10057 , new_n10057 );
  nor      g09682 ( new_n10059 , new_n6514 , new_n10058 );
  nand     g09683 ( new_n10060 , new_n10055 , new_n10059 );
  nand     g09684 ( new_n10061 , new_n10054 , new_n10060 );
  xor      g09685 ( new_n10062 , new_n10052 , new_n10061 );
  nor      g09686 ( new_n10063 , new_n10036 , new_n10062 );
  nand     g09687 ( new_n10064 , new_n6537 , new_n6538 );
  or       g09688 ( new_n10065 , new_n6535 , new_n6539 );
  and      g09689 ( new_n10066 , new_n10064 , new_n10065 );
  xor      g09690 ( new_n10067 , new_n10036 , new_n10062 );
  and      g09691 ( new_n10068 , new_n10066 , new_n10067 );
  nor      g09692 ( new_n10069 , new_n10063 , new_n10068 );
  xor      g09693 ( new_n10070 , new_n10035 , new_n10069 );
  nor      g09694 ( new_n10071 , new_n6548 , new_n6573 );
  nand     g09695 ( new_n10072 , pi018 , pi051 );
  nand     g09696 ( new_n10073 , pi090 , pi108 );
  xor      g09697 ( new_n10074 , new_n10072 , new_n10073 );
  xor      g09698 ( new_n10075 , new_n6560 , new_n10074 );
  nand     g09699 ( new_n10076 , pi007 , pi141 );
  xor      g09700 ( new_n10077 , new_n6561 , new_n10076 );
  xnor     g09701 ( new_n10078 , new_n10075 , new_n10077 );
  nor      g09702 ( new_n10079 , new_n6552 , new_n6555 );
  nor      g09703 ( new_n10080 , new_n6556 , new_n6563 );
  nor      g09704 ( new_n10081 , new_n10079 , new_n10080 );
  nand     g09705 ( new_n10082 , pi113 , pi241 );
  nand     g09706 ( new_n10083 , pi038 , pi236 );
  xor      g09707 ( new_n10084 , new_n10082 , new_n10083 );
  xor      g09708 ( new_n10085 , new_n6565 , new_n10084 );
  xor      g09709 ( new_n10086 , new_n10081 , new_n10085 );
  xor      g09710 ( new_n10087 , new_n10078 , new_n10086 );
  nor      g09711 ( new_n10088 , new_n6564 , new_n6570 );
  nor      g09712 ( new_n10089 , new_n6551 , new_n6571 );
  xor      g09713 ( new_n10090 , new_n6566 , new_n10089 );
  nor      g09714 ( new_n10091 , new_n10088 , new_n10090 );
  xor      g09715 ( new_n10092 , new_n10087 , new_n10091 );
  xnor     g09716 ( new_n10093 , new_n10071 , new_n10092 );
  nand     g09717 ( new_n10094 , new_n6575 , new_n6576 );
  or       g09718 ( new_n10095 , new_n6574 , new_n6577 );
  nand     g09719 ( new_n10096 , new_n10094 , new_n10095 );
  nand g09720 ( new_n10097 , new_n10096 , new_n10096 );
  xor      g09721 ( new_n10098 , new_n10093 , new_n10097 );
  nand     g09722 ( new_n10099 , new_n6580 , new_n6607 );
  nand     g09723 ( new_n10100 , new_n6579 , new_n6608 );
  nand     g09724 ( new_n10101 , new_n10099 , new_n10100 );
  nand     g09725 ( new_n10102 , new_n6603 , new_n6606 );
  nand     g09726 ( new_n10103 , new_n6590 , new_n6596 );
  nand     g09727 ( new_n10104 , new_n6589 , new_n6597 );
  nand     g09728 ( new_n10105 , new_n10103 , new_n10104 );
  nand     g09729 ( new_n10106 , pi098 , pi212 );
  nand     g09730 ( new_n10107 , pi043 , pi213 );
  xor      g09731 ( new_n10108 , new_n10106 , new_n10107 );
  xor      g09732 ( new_n10109 , new_n6584 , new_n10108 );
  xor      g09733 ( new_n10110 , new_n10105 , new_n10109 );
  nand     g09734 ( new_n10111 , pi012 , pi013 );
  xor      g09735 ( new_n10112 , new_n6595 , new_n10111 );
  nand     g09736 ( new_n10113 , pi183 , pi188 );
  nand     g09737 ( new_n10114 , pi061 , pi112 );
  xor      g09738 ( new_n10115 , new_n10113 , new_n10114 );
  xor      g09739 ( new_n10116 , new_n6594 , new_n10115 );
  xor      g09740 ( new_n10117 , new_n10112 , new_n10116 );
  xor      g09741 ( new_n10118 , new_n10110 , new_n10117 );
  nor      g09742 ( new_n10119 , new_n6586 , new_n6598 );
  nor      g09743 ( new_n10120 , new_n6599 , new_n6602 );
  xor      g09744 ( new_n10121 , new_n6585 , new_n10120 );
  nor      g09745 ( new_n10122 , new_n10119 , new_n10121 );
  xor      g09746 ( new_n10123 , new_n10118 , new_n10122 );
  nand g09747 ( new_n10124 , new_n10123 , new_n10123 );
  xor      g09748 ( new_n10125 , new_n10102 , new_n10124 );
  xor      g09749 ( new_n10126 , new_n10101 , new_n10125 );
  xor      g09750 ( new_n10127 , new_n10098 , new_n10126 );
  nor      g09751 ( new_n10128 , new_n6578 , new_n6609 );
  nor      g09752 ( new_n10129 , new_n6545 , new_n6610 );
  nor      g09753 ( new_n10130 , new_n10128 , new_n10129 );
  xnor     g09754 ( new_n10131 , new_n10127 , new_n10130 );
  xnor     g09755 ( new_n10132 , new_n10066 , new_n10067 );
  nand     g09756 ( new_n10133 , new_n10131 , new_n10132 );
  nand     g09757 ( new_n10134 , new_n6506 , new_n6540 );
  nand     g09758 ( new_n10135 , new_n6541 , new_n6611 );
  and      g09759 ( new_n10136 , new_n10134 , new_n10135 );
  xor      g09760 ( new_n10137 , new_n10131 , new_n10132 );
  nand     g09761 ( new_n10138 , new_n10136 , new_n10137 );
  nand     g09762 ( new_n10139 , new_n10133 , new_n10138 );
  nand     g09763 ( new_n10140 , pi064 , pi194 );
  xor      g09764 ( new_n10141 , new_n10139 , new_n10140 );
  nand     g09765 ( new_n10142 , pi057 , pi084 );
  nand     g09766 ( new_n10143 , pi028 , pi236 );
  xor      g09767 ( new_n10144 , new_n10142 , new_n10143 );
  xor      g09768 ( new_n10145 , new_n10141 , new_n10144 );
  xor      g09769 ( new_n10146 , new_n10070 , new_n10145 );
  nand     g09770 ( new_n10147 , pi052 , pi068 );
  nand     g09771 ( new_n10148 , pi012 , pi112 );
  nor      g09772 ( new_n10149 , new_n10102 , new_n10124 );
  nand g09773 ( new_n10150 , new_n10125 , new_n10125 );
  nor      g09774 ( new_n10151 , new_n10101 , new_n10150 );
  nor      g09775 ( new_n10152 , new_n10149 , new_n10151 );
  xor      g09776 ( new_n10153 , new_n10148 , new_n10152 );
  xor      g09777 ( new_n10154 , new_n10147 , new_n10153 );
  nand     g09778 ( new_n10155 , pi043 , pi212 );
  nand     g09779 ( new_n10156 , pi047 , pi108 );
  xor      g09780 ( new_n10157 , new_n10155 , new_n10156 );
  nand     g09781 ( new_n10158 , pi098 , pi104 );
  nand     g09782 ( new_n10159 , pi013 , pi144 );
  nand     g09783 ( new_n10160 , pi133 , pi180 );
  xnor     g09784 ( new_n10161 , new_n10159 , new_n10160 );
  xor      g09785 ( new_n10162 , new_n10158 , new_n10161 );
  xor      g09786 ( new_n10163 , new_n10157 , new_n10162 );
  nand     g09787 ( new_n10164 , new_n10047 , new_n10048 );
  nand     g09788 ( new_n10165 , new_n6513 , new_n10049 );
  nand     g09789 ( new_n10166 , new_n10164 , new_n10165 );
  xor      g09790 ( new_n10167 , new_n10163 , new_n10166 );
  xor      g09791 ( new_n10168 , new_n10154 , new_n10167 );
  nand     g09792 ( new_n10169 , pi085 , pi189 );
  nand     g09793 ( new_n10170 , pi036 , pi077 );
  xor      g09794 ( new_n10171 , new_n10169 , new_n10170 );
  nand     g09795 ( new_n10172 , pi113 , pi161 );
  nand     g09796 ( new_n10173 , pi035 , pi237 );
  xor      g09797 ( new_n10174 , new_n10172 , new_n10173 );
  xor      g09798 ( new_n10175 , new_n10171 , new_n10174 );
  xor      g09799 ( new_n10176 , new_n10168 , new_n10175 );
  xor      g09800 ( new_n10177 , new_n10146 , new_n10176 );
  nand     g09801 ( new_n10178 , pi007 , pi090 );
  nand     g09802 ( new_n10179 , pi051 , pi128 );
  nand     g09803 ( new_n10180 , new_n10082 , new_n10083 );
  nand     g09804 ( new_n10181 , new_n6565 , new_n10084 );
  nand     g09805 ( new_n10182 , new_n10180 , new_n10181 );
  nand     g09806 ( new_n10183 , pi189 , pi194 );
  nand     g09807 ( new_n10184 , pi084 , pi143 );
  nand     g09808 ( new_n10185 , new_n10183 , new_n10184 );
  xor      g09809 ( new_n10186 , new_n10183 , new_n10184 );
  nand     g09810 ( new_n10187 , new_n6636 , new_n10186 );
  nand     g09811 ( new_n10188 , new_n10185 , new_n10187 );
  xor      g09812 ( new_n10189 , new_n10182 , new_n10188 );
  xor      g09813 ( new_n10190 , new_n10179 , new_n10189 );
  xor      g09814 ( new_n10191 , new_n10178 , new_n10190 );
  nor      g09815 ( new_n10192 , new_n6621 , new_n6646 );
  nand g09816 ( new_n10193 , new_n10192 , new_n10192 );
  xor      g09817 ( new_n10194 , new_n6636 , new_n10186 );
  nand     g09818 ( new_n10195 , pi085 , pi133 );
  xor      g09819 ( new_n10196 , new_n6637 , new_n10195 );
  xnor     g09820 ( new_n10197 , new_n10194 , new_n10196 );
  nand     g09821 ( new_n10198 , new_n6632 , new_n6639 );
  nand     g09822 ( new_n10199 , new_n6631 , new_n6640 );
  nand     g09823 ( new_n10200 , new_n10198 , new_n10199 );
  xor      g09824 ( new_n10201 , new_n6625 , new_n10033 );
  xnor     g09825 ( new_n10202 , new_n10200 , new_n10201 );
  xnor     g09826 ( new_n10203 , new_n10197 , new_n10202 );
  nand g09827 ( new_n10204 , new_n6645 , new_n6645 );
  nand     g09828 ( new_n10205 , new_n6642 , new_n10204 );
  nor      g09829 ( new_n10206 , new_n6628 , new_n6641 );
  nor      g09830 ( new_n10207 , new_n6626 , new_n10206 );
  nand     g09831 ( new_n10208 , new_n10205 , new_n10207 );
  nand g09832 ( new_n10209 , new_n10208 , new_n10208 );
  nor      g09833 ( new_n10210 , new_n6627 , new_n10205 );
  nor      g09834 ( new_n10211 , new_n10209 , new_n10210 );
  xor      g09835 ( new_n10212 , new_n10203 , new_n10211 );
  nor      g09836 ( new_n10213 , new_n10193 , new_n10212 );
  xor      g09837 ( new_n10214 , new_n10193 , new_n10212 );
  nand g09838 ( new_n10215 , new_n10214 , new_n10214 );
  nand     g09839 ( new_n10216 , new_n6616 , new_n6617 );
  nand g09840 ( new_n10217 , new_n6647 , new_n6647 );
  nand     g09841 ( new_n10218 , new_n6618 , new_n10217 );
  nand     g09842 ( new_n10219 , new_n10216 , new_n10218 );
  nor      g09843 ( new_n10220 , new_n10215 , new_n10219 );
  or       g09844 ( new_n10221 , new_n10213 , new_n10220 );
  nand     g09845 ( new_n10222 , pi033 , pi146 );
  xor      g09846 ( new_n10223 , new_n10221 , new_n10222 );
  xor      g09847 ( new_n10224 , new_n10191 , new_n10223 );
  nand     g09848 ( new_n10225 , new_n10081 , new_n10085 );
  nand     g09849 ( new_n10226 , new_n10078 , new_n10086 );
  nand     g09850 ( new_n10227 , new_n10225 , new_n10226 );
  nor      g09851 ( new_n10228 , new_n6638 , new_n10195 );
  nor      g09852 ( new_n10229 , new_n10194 , new_n10196 );
  nor      g09853 ( new_n10230 , new_n10228 , new_n10229 );
  nand     g09854 ( new_n10231 , new_n10203 , new_n10211 );
  nand     g09855 ( new_n10232 , new_n10208 , new_n10231 );
  xor      g09856 ( new_n10233 , new_n10230 , new_n10232 );
  nand     g09857 ( new_n10234 , pi139 , pi238 );
  xor      g09858 ( new_n10235 , new_n10233 , new_n10234 );
  xor      g09859 ( new_n10236 , new_n10227 , new_n10235 );
  nor      g09860 ( new_n10237 , new_n6595 , new_n10111 );
  nand g09861 ( new_n10238 , new_n10112 , new_n10112 );
  nor      g09862 ( new_n10239 , new_n10238 , new_n10116 );
  nor      g09863 ( new_n10240 , new_n10237 , new_n10239 );
  nand     g09864 ( new_n10241 , pi193 , pi208 );
  xor      g09865 ( new_n10242 , new_n10240 , new_n10241 );
  xor      g09866 ( new_n10243 , new_n10236 , new_n10242 );
  xor      g09867 ( new_n10244 , new_n10224 , new_n10243 );
  nand     g09868 ( new_n10245 , new_n10113 , new_n10114 );
  nand     g09869 ( new_n10246 , new_n6594 , new_n10115 );
  nand     g09870 ( new_n10247 , new_n10245 , new_n10246 );
  nor      g09871 ( new_n10248 , new_n10098 , new_n10126 );
  and      g09872 ( new_n10249 , new_n10127 , new_n10130 );
  nor      g09873 ( new_n10250 , new_n10248 , new_n10249 );
  nand     g09874 ( new_n10251 , pi046 , pi131 );
  and      g09875 ( new_n10252 , new_n6585 , new_n10120 );
  nor      g09876 ( new_n10253 , new_n10118 , new_n10122 );
  nor      g09877 ( new_n10254 , new_n10252 , new_n10253 );
  nand     g09878 ( new_n10255 , pi126 , pi213 );
  nand     g09879 ( new_n10256 , pi015 , pi048 );
  xor      g09880 ( new_n10257 , new_n10255 , new_n10256 );
  xor      g09881 ( new_n10258 , new_n10254 , new_n10257 );
  xor      g09882 ( new_n10259 , new_n10251 , new_n10258 );
  xor      g09883 ( new_n10260 , new_n10250 , new_n10259 );
  xor      g09884 ( new_n10261 , new_n10247 , new_n10260 );
  nor      g09885 ( new_n10262 , new_n10046 , new_n10050 );
  nor      g09886 ( new_n10263 , new_n10043 , new_n10051 );
  nor      g09887 ( new_n10264 , new_n10262 , new_n10263 );
  nand     g09888 ( new_n10265 , pi061 , pi105 );
  nand     g09889 ( new_n10266 , pi034 , pi143 );
  xor      g09890 ( new_n10267 , new_n10265 , new_n10266 );
  xor      g09891 ( new_n10268 , new_n10264 , new_n10267 );
  nand     g09892 ( new_n10269 , new_n10072 , new_n10073 );
  nand     g09893 ( new_n10270 , new_n6560 , new_n10074 );
  nand     g09894 ( new_n10271 , new_n10269 , new_n10270 );
  nand     g09895 ( new_n10272 , pi038 , pi241 );
  nand     g09896 ( new_n10273 , pi018 , pi042 );
  xnor     g09897 ( new_n10274 , new_n10272 , new_n10273 );
  xor      g09898 ( new_n10275 , new_n10271 , new_n10274 );
  xor      g09899 ( new_n10276 , new_n10268 , new_n10275 );
  xor      g09900 ( new_n10277 , new_n10261 , new_n10276 );
  xor      g09901 ( new_n10278 , new_n10215 , new_n10219 );
  xnor     g09902 ( new_n10279 , new_n10136 , new_n10137 );
  and      g09903 ( new_n10280 , new_n10278 , new_n10279 );
  xnor     g09904 ( new_n10281 , new_n10278 , new_n10279 );
  or       g09905 ( new_n10282 , new_n6615 , new_n6648 );
  nand     g09906 ( new_n10283 , new_n6612 , new_n6649 );
  nand     g09907 ( new_n10284 , new_n10282 , new_n10283 );
  nor      g09908 ( new_n10285 , new_n10281 , new_n10284 );
  nor      g09909 ( new_n10286 , new_n10280 , new_n10285 );
  nand     g09910 ( new_n10287 , pi088 , pi188 );
  nand     g09911 ( new_n10288 , pi159 , pi168 );
  or       g09912 ( new_n10289 , new_n10052 , new_n10061 );
  nand     g09913 ( new_n10290 , new_n10060 , new_n10289 );
  xnor     g09914 ( new_n10291 , new_n10288 , new_n10290 );
  xor      g09915 ( new_n10292 , new_n10287 , new_n10291 );
  xor      g09916 ( new_n10293 , new_n10286 , new_n10292 );
  xor      g09917 ( new_n10294 , new_n10277 , new_n10293 );
  nand     g09918 ( new_n10295 , pi118 , pi141 );
  nand     g09919 ( new_n10296 , new_n10037 , new_n10038 );
  nand     g09920 ( new_n10297 , new_n6523 , new_n10039 );
  nand     g09921 ( new_n10298 , new_n10296 , new_n10297 );
  nand     g09922 ( new_n10299 , pi178 , pi183 );
  xor      g09923 ( new_n10300 , new_n10298 , new_n10299 );
  nor      g09924 ( new_n10301 , new_n10071 , new_n10092 );
  nor      g09925 ( new_n10302 , new_n10093 , new_n10097 );
  nor      g09926 ( new_n10303 , new_n10301 , new_n10302 );
  nand     g09927 ( new_n10304 , new_n10105 , new_n10109 );
  nand     g09928 ( new_n10305 , new_n10110 , new_n10117 );
  nand     g09929 ( new_n10306 , new_n10304 , new_n10305 );
  nand     g09930 ( new_n10307 , new_n10106 , new_n10107 );
  nand     g09931 ( new_n10308 , new_n6584 , new_n10108 );
  nand     g09932 ( new_n10309 , new_n10307 , new_n10308 );
  xnor     g09933 ( new_n10310 , new_n10306 , new_n10309 );
  xor      g09934 ( new_n10311 , new_n10303 , new_n10310 );
  xor      g09935 ( new_n10312 , new_n10300 , new_n10311 );
  xor      g09936 ( new_n10313 , new_n10295 , new_n10312 );
  nor      g09937 ( new_n10314 , new_n6562 , new_n10076 );
  nor      g09938 ( new_n10315 , new_n10075 , new_n10077 );
  nor      g09939 ( new_n10316 , new_n10314 , new_n10315 );
  nor      g09940 ( new_n10317 , new_n10200 , new_n10201 );
  nor      g09941 ( new_n10318 , new_n10197 , new_n10202 );
  nor      g09942 ( new_n10319 , new_n10317 , new_n10318 );
  xor      g09943 ( new_n10320 , new_n10316 , new_n10319 );
  or       g09944 ( new_n10321 , new_n6525 , new_n10041 );
  nand g09945 ( new_n10322 , new_n10042 , new_n10042 );
  nand     g09946 ( new_n10323 , new_n10040 , new_n10322 );
  nand     g09947 ( new_n10324 , new_n10321 , new_n10323 );
  nand     g09948 ( new_n10325 , pi179 , pi204 );
  xor      g09949 ( new_n10326 , new_n10324 , new_n10325 );
  and      g09950 ( new_n10327 , new_n6566 , new_n10089 );
  nor      g09951 ( new_n10328 , new_n10087 , new_n10091 );
  nor      g09952 ( new_n10329 , new_n10327 , new_n10328 );
  nand     g09953 ( new_n10330 , pi152 , pi162 );
  xor      g09954 ( new_n10331 , new_n10329 , new_n10330 );
  xor      g09955 ( new_n10332 , new_n10326 , new_n10331 );
  xor      g09956 ( new_n10333 , new_n10320 , new_n10332 );
  xor      g09957 ( new_n10334 , new_n10313 , new_n10333 );
  xor      g09958 ( new_n10335 , new_n10294 , new_n10334 );
  xor      g09959 ( new_n10336 , new_n10244 , new_n10335 );
  xor      g09960 ( po072 , new_n10177 , new_n10336 );
  xor      g09961 ( po073 , new_n913 , new_n914 );
  xor      g09962 ( po074 , new_n6380 , new_n6381 );
  xor      g09963 ( po075 , new_n7642 , new_n7643 );
  xor      g09964 ( po076 , new_n6726 , new_n6727 );
  xor      g09965 ( po077 , new_n1085 , new_n1091 );
  xor      g09966 ( po078 , new_n1898 , new_n1905 );
  xnor     g09967 ( po079 , new_n5915 , new_n5916 );
  xor      g09968 ( po080 , new_n9430 , new_n9432 );
  xor      g09969 ( po081 , new_n7635 , new_n7637 );
  xor      g09970 ( po082 , new_n6383 , new_n6384 );
  xnor     g09971 ( po083 , new_n1116 , new_n1117 );
  nand     g09972 ( new_n10349 , new_n816 , new_n880 );
  or       g09973 ( new_n10350 , new_n787 , new_n881 );
  nand     g09974 ( new_n10351 , new_n10349 , new_n10350 );
  nor      g09975 ( new_n10352 , new_n736 , new_n803 );
  nand g09976 ( new_n10353 , new_n804 , new_n804 );
  nor      g09977 ( new_n10354 , new_n10353 , new_n808 );
  nor      g09978 ( new_n10355 , new_n10352 , new_n10354 );
  xor      g09979 ( new_n10356 , new_n10351 , new_n10355 );
  nand     g09980 ( new_n10357 , new_n552 , new_n873 );
  or       g09981 ( new_n10358 , new_n871 , new_n875 );
  nand     g09982 ( new_n10359 , new_n10357 , new_n10358 );
  nand     g09983 ( new_n10360 , pi097 , pi167 );
  nand     g09984 ( new_n10361 , pi011 , pi175 );
  xnor     g09985 ( new_n10362 , new_n10360 , new_n10361 );
  nand     g09986 ( new_n10363 , pi075 , pi149 );
  xor      g09987 ( new_n10364 , new_n10362 , new_n10363 );
  xor      g09988 ( new_n10365 , new_n10359 , new_n10364 );
  xor      g09989 ( new_n10366 , new_n10356 , new_n10365 );
  nand     g09990 ( new_n10367 , new_n789 , new_n811 );
  nand g09991 ( new_n10368 , new_n815 , new_n815 );
  nand     g09992 ( new_n10369 , new_n812 , new_n10368 );
  nand     g09993 ( new_n10370 , new_n10367 , new_n10369 );
  nand     g09994 ( new_n10371 , pi117 , pi248 );
  nand     g09995 ( new_n10372 , new_n438 , new_n483 );
  nand     g09996 ( new_n10373 , new_n482 , new_n484 );
  nand     g09997 ( new_n10374 , new_n10372 , new_n10373 );
  xnor     g09998 ( new_n10375 , new_n10371 , new_n10374 );
  xor      g09999 ( new_n10376 , new_n10370 , new_n10375 );
  or       g10000 ( new_n10377 , new_n471 , new_n488 );
  nand     g10001 ( new_n10378 , new_n469 , new_n10377 );
  nand     g10002 ( new_n10379 , pi044 , pi247 );
  nand     g10003 ( new_n10380 , pi054 , pi080 );
  xor      g10004 ( new_n10381 , new_n10379 , new_n10380 );
  xor      g10005 ( new_n10382 , new_n10378 , new_n10381 );
  xor      g10006 ( new_n10383 , new_n10376 , new_n10382 );
  xor      g10007 ( new_n10384 , new_n10366 , new_n10383 );
  nand     g10008 ( new_n10385 , pi016 , pi072 );
  nand     g10009 ( new_n10386 , pi031 , pi163 );
  xor      g10010 ( new_n10387 , new_n10385 , new_n10386 );
  and      g10011 ( new_n10388 , new_n726 , new_n791 );
  nor      g10012 ( new_n10389 , new_n793 , new_n810 );
  nor      g10013 ( new_n10390 , new_n10388 , new_n10389 );
  nand     g10014 ( new_n10391 , pi045 , pi214 );
  nand     g10015 ( new_n10392 , new_n842 , new_n843 );
  nand     g10016 ( new_n10393 , new_n615 , new_n844 );
  nand     g10017 ( new_n10394 , new_n10392 , new_n10393 );
  xor      g10018 ( new_n10395 , new_n10391 , new_n10394 );
  xor      g10019 ( new_n10396 , new_n10390 , new_n10395 );
  xor      g10020 ( new_n10397 , new_n10387 , new_n10396 );
  xor      g10021 ( new_n10398 , new_n10384 , new_n10397 );
  nand     g10022 ( new_n10399 , pi147 , pi203 );
  nand     g10023 ( new_n10400 , pi151 , pi200 );
  xor      g10024 ( new_n10401 , new_n10399 , new_n10400 );
  nand     g10025 ( new_n10402 , pi027 , pi083 );
  nor      g10026 ( new_n10403 , new_n463 , new_n489 );
  nor      g10027 ( new_n10404 , new_n462 , new_n490 );
  nor      g10028 ( new_n10405 , new_n10403 , new_n10404 );
  xor      g10029 ( new_n10406 , new_n10402 , new_n10405 );
  nand     g10030 ( new_n10407 , pi049 , pi096 );
  nor      g10031 ( new_n10408 , new_n617 , new_n840 );
  nor      g10032 ( new_n10409 , new_n841 , new_n845 );
  nor      g10033 ( new_n10410 , new_n10408 , new_n10409 );
  xor      g10034 ( new_n10411 , new_n10407 , new_n10410 );
  nand     g10035 ( new_n10412 , new_n832 , new_n833 );
  nand     g10036 ( new_n10413 , new_n627 , new_n834 );
  nand     g10037 ( new_n10414 , new_n10412 , new_n10413 );
  nand     g10038 ( new_n10415 , pi119 , pi202 );
  xor      g10039 ( new_n10416 , new_n10414 , new_n10415 );
  xor      g10040 ( new_n10417 , new_n10411 , new_n10416 );
  xor      g10041 ( new_n10418 , new_n10406 , new_n10417 );
  xor      g10042 ( new_n10419 , new_n10401 , new_n10418 );
  xor      g10043 ( new_n10420 , new_n10398 , new_n10419 );
  nor      g10044 ( new_n10421 , new_n446 , new_n476 );
  nor      g10045 ( new_n10422 , new_n475 , new_n477 );
  nor      g10046 ( new_n10423 , new_n10421 , new_n10422 );
  nand     g10047 ( new_n10424 , new_n472 , new_n473 );
  nand     g10048 ( new_n10425 , new_n444 , new_n474 );
  nand     g10049 ( new_n10426 , new_n10424 , new_n10425 );
  xor      g10050 ( new_n10427 , new_n10423 , new_n10426 );
  nand g10051 ( new_n10428 , new_n878 , new_n878 );
  nor      g10052 ( new_n10429 , new_n850 , new_n10428 );
  nand g10053 ( new_n10430 , new_n879 , new_n879 );
  nor      g10054 ( new_n10431 , new_n823 , new_n10430 );
  nor      g10055 ( new_n10432 , new_n10429 , new_n10431 );
  nor      g10056 ( new_n10433 , new_n481 , new_n485 );
  nand g10057 ( new_n10434 , new_n478 , new_n478 );
  nor      g10058 ( new_n10435 , new_n10434 , new_n486 );
  nor      g10059 ( new_n10436 , new_n10433 , new_n10435 );
  xor      g10060 ( new_n10437 , new_n10432 , new_n10436 );
  nand     g10061 ( new_n10438 , pi039 , pi246 );
  nor      g10062 ( new_n10439 , new_n827 , new_n848 );
  nor      g10063 ( new_n10440 , new_n826 , new_n849 );
  nor      g10064 ( new_n10441 , new_n10439 , new_n10440 );
  nand     g10065 ( new_n10442 , pi056 , pi201 );
  nand     g10066 ( new_n10443 , new_n866 , new_n867 );
  nand     g10067 ( new_n10444 , new_n551 , new_n868 );
  nand     g10068 ( new_n10445 , new_n10443 , new_n10444 );
  xor      g10069 ( new_n10446 , new_n10442 , new_n10445 );
  xor      g10070 ( new_n10447 , new_n10441 , new_n10446 );
  nand     g10071 ( new_n10448 , pi136 , pi245 );
  nand     g10072 ( new_n10449 , pi116 , pi145 );
  nand     g10073 ( new_n10450 , new_n858 , new_n859 );
  nand     g10074 ( new_n10451 , new_n540 , new_n860 );
  nand     g10075 ( new_n10452 , new_n10450 , new_n10451 );
  xor      g10076 ( new_n10453 , new_n10449 , new_n10452 );
  xor      g10077 ( new_n10454 , new_n10448 , new_n10453 );
  xor      g10078 ( new_n10455 , new_n10447 , new_n10454 );
  xor      g10079 ( new_n10456 , new_n10438 , new_n10455 );
  xor      g10080 ( new_n10457 , new_n10437 , new_n10456 );
  xor      g10081 ( new_n10458 , new_n10427 , new_n10457 );
  xor      g10082 ( new_n10459 , new_n10420 , new_n10458 );
  nor      g10083 ( new_n10460 , new_n629 , new_n830 );
  nand g10084 ( new_n10461 , new_n847 , new_n847 );
  nor      g10085 ( new_n10462 , new_n831 , new_n10461 );
  nor      g10086 ( new_n10463 , new_n10460 , new_n10462 );
  nand     g10087 ( new_n10464 , new_n865 , new_n869 );
  nand     g10088 ( new_n10465 , new_n862 , new_n870 );
  nand     g10089 ( new_n10466 , new_n10464 , new_n10465 );
  nand     g10090 ( new_n10467 , pi171 , pi235 );
  nor      g10091 ( new_n10468 , new_n541 , new_n856 );
  nor      g10092 ( new_n10469 , new_n857 , new_n861 );
  nor      g10093 ( new_n10470 , new_n10468 , new_n10469 );
  xor      g10094 ( new_n10471 , new_n10467 , new_n10470 );
  xor      g10095 ( new_n10472 , new_n10466 , new_n10471 );
  xor      g10096 ( new_n10473 , new_n10463 , new_n10472 );
  xor      g10097 ( new_n10474 , new_n10459 , new_n10473 );
  nand     g10098 ( new_n10475 , new_n855 , new_n876 );
  nand     g10099 ( new_n10476 , new_n854 , new_n877 );
  nand     g10100 ( new_n10477 , new_n10475 , new_n10476 );
  nand     g10101 ( new_n10478 , pi026 , pi063 );
  nand     g10102 ( new_n10479 , new_n835 , new_n838 );
  nand g10103 ( new_n10480 , new_n839 , new_n839 );
  nand     g10104 ( new_n10481 , new_n10480 , new_n846 );
  nand     g10105 ( new_n10482 , new_n10479 , new_n10481 );
  nand     g10106 ( new_n10483 , new_n798 , new_n801 );
  nand     g10107 ( new_n10484 , new_n802 , new_n809 );
  nand     g10108 ( new_n10485 , new_n10483 , new_n10484 );
  xnor     g10109 ( new_n10486 , new_n10482 , new_n10485 );
  xor      g10110 ( new_n10487 , new_n10478 , new_n10486 );
  xor      g10111 ( new_n10488 , new_n10477 , new_n10487 );
  xor      g10112 ( new_n10489 , new_n10474 , new_n10488 );
  nand     g10113 ( new_n10490 , pi107 , pi110 );
  nand     g10114 ( new_n10491 , pi091 , pi148 );
  nand g10115 ( new_n10492 , new_n882 , new_n882 );
  nor      g10116 ( new_n10493 , new_n491 , new_n10492 );
  nor      g10117 ( new_n10494 , new_n883 , new_n923 );
  nor      g10118 ( new_n10495 , new_n10493 , new_n10494 );
  xor      g10119 ( new_n10496 , new_n10491 , new_n10495 );
  xor      g10120 ( new_n10497 , new_n10490 , new_n10496 );
  nand     g10121 ( new_n10498 , pi008 , pi156 );
  nand     g10122 ( new_n10499 , pi000 , pi164 );
  xor      g10123 ( new_n10500 , new_n10498 , new_n10499 );
  nand     g10124 ( new_n10501 , pi019 , pi181 );
  nand     g10125 ( new_n10502 , new_n805 , new_n806 );
  nand     g10126 ( new_n10503 , new_n735 , new_n807 );
  nand     g10127 ( new_n10504 , new_n10502 , new_n10503 );
  xor      g10128 ( new_n10505 , new_n10501 , new_n10504 );
  nand     g10129 ( new_n10506 , pi134 , pi166 );
  nand g10130 ( new_n10507 , new_n795 , new_n795 );
  nor      g10131 ( new_n10508 , new_n10507 , new_n796 );
  nor      g10132 ( new_n10509 , new_n794 , new_n797 );
  nor      g10133 ( new_n10510 , new_n10508 , new_n10509 );
  nand     g10134 ( new_n10511 , pi032 , pi070 );
  xor      g10135 ( new_n10512 , new_n10510 , new_n10511 );
  xor      g10136 ( new_n10513 , new_n10506 , new_n10512 );
  xor      g10137 ( new_n10514 , new_n10505 , new_n10513 );
  nand     g10138 ( new_n10515 , pi114 , pi228 );
  nand     g10139 ( new_n10516 , pi009 , pi103 );
  xor      g10140 ( new_n10517 , new_n10515 , new_n10516 );
  nand     g10141 ( new_n10518 , pi115 , pi206 );
  nand     g10142 ( new_n10519 , pi093 , pi240 );
  nand     g10143 ( new_n10520 , pi234 , pi250 );
  xnor     g10144 ( new_n10521 , new_n10519 , new_n10520 );
  xor      g10145 ( new_n10522 , new_n10518 , new_n10521 );
  xor      g10146 ( new_n10523 , new_n10517 , new_n10522 );
  xor      g10147 ( new_n10524 , new_n10514 , new_n10523 );
  xor      g10148 ( new_n10525 , new_n10500 , new_n10524 );
  xor      g10149 ( new_n10526 , new_n10497 , new_n10525 );
  xor      g10150 ( po084 , new_n10489 , new_n10526 );
  xor      g10151 ( po085 , new_n10281 , new_n10284 );
  nor      g10152 ( new_n10529 , new_n9750 , new_n9781 );
  nand g10153 ( new_n10530 , new_n9782 , new_n9782 );
  nor      g10154 ( new_n10531 , new_n9716 , new_n10530 );
  nor      g10155 ( new_n10532 , new_n10529 , new_n10531 );
  nor      g10156 ( new_n10533 , new_n9817 , new_n9848 );
  nor      g10157 ( new_n10534 , new_n9713 , new_n9849 );
  nor      g10158 ( new_n10535 , new_n10533 , new_n10534 );
  xor      g10159 ( new_n10536 , new_n10532 , new_n10535 );
  nand     g10160 ( new_n10537 , pi081 , pi189 );
  xor      g10161 ( new_n10538 , new_n10536 , new_n10537 );
  nand     g10162 ( new_n10539 , new_n9791 , new_n9812 );
  or       g10163 ( new_n10540 , new_n9790 , new_n9814 );
  nand     g10164 ( new_n10541 , new_n10539 , new_n10540 );
  nand     g10165 ( new_n10542 , new_n9786 , new_n9815 );
  nand g10166 ( new_n10543 , new_n9783 , new_n9783 );
  or       g10167 ( new_n10544 , new_n10543 , new_n9816 );
  nand     g10168 ( new_n10545 , new_n10542 , new_n10544 );
  nand     g10169 ( new_n10546 , pi104 , pi127 );
  xor      g10170 ( new_n10547 , new_n10545 , new_n10546 );
  nand     g10171 ( new_n10548 , new_n9835 , new_n9836 );
  nand     g10172 ( new_n10549 , new_n9584 , new_n9837 );
  nand     g10173 ( new_n10550 , new_n10548 , new_n10549 );
  nand g10174 ( new_n10551 , new_n9798 , new_n9798 );
  nor      g10175 ( new_n10552 , new_n9795 , new_n10551 );
  nand g10176 ( new_n10553 , new_n9806 , new_n9806 );
  nor      g10177 ( new_n10554 , new_n9799 , new_n10553 );
  nor      g10178 ( new_n10555 , new_n10552 , new_n10554 );
  nand     g10179 ( new_n10556 , pi157 , pi208 );
  xor      g10180 ( new_n10557 , new_n10555 , new_n10556 );
  xor      g10181 ( new_n10558 , new_n10550 , new_n10557 );
  nand     g10182 ( new_n10559 , pi052 , pi187 );
  or       g10183 ( new_n10560 , new_n9823 , new_n9846 );
  nand     g10184 ( new_n10561 , new_n9818 , new_n9847 );
  nand     g10185 ( new_n10562 , new_n10560 , new_n10561 );
  xor      g10186 ( new_n10563 , new_n10559 , new_n10562 );
  nand     g10187 ( new_n10564 , pi084 , pi100 );
  nor      g10188 ( new_n10565 , new_n9585 , new_n9833 );
  nand g10189 ( new_n10566 , new_n9834 , new_n9834 );
  nor      g10190 ( new_n10567 , new_n10566 , new_n9838 );
  nor      g10191 ( new_n10568 , new_n10565 , new_n10567 );
  xor      g10192 ( new_n10569 , new_n10564 , new_n10568 );
  xor      g10193 ( new_n10570 , new_n10563 , new_n10569 );
  xor      g10194 ( new_n10571 , new_n10558 , new_n10570 );
  nand     g10195 ( new_n10572 , pi035 , pi040 );
  nand     g10196 ( new_n10573 , new_n9792 , new_n9793 );
  nand     g10197 ( new_n10574 , new_n9615 , new_n9794 );
  nand     g10198 ( new_n10575 , new_n10573 , new_n10574 );
  xor      g10199 ( new_n10576 , new_n10572 , new_n10575 );
  nand     g10200 ( new_n10577 , new_n9616 , new_n9808 );
  nand     g10201 ( new_n10578 , new_n9807 , new_n9811 );
  nand     g10202 ( new_n10579 , new_n10577 , new_n10578 );
  nand     g10203 ( new_n10580 , pi152 , pi249 );
  xor      g10204 ( new_n10581 , new_n10579 , new_n10580 );
  nand     g10205 ( new_n10582 , pi064 , pi227 );
  nor      g10206 ( new_n10583 , new_n9754 , new_n9778 );
  nor      g10207 ( new_n10584 , new_n9779 , new_n10583 );
  nor      g10208 ( new_n10585 , new_n9682 , new_n9758 );
  nand g10209 ( new_n10586 , new_n9759 , new_n9759 );
  nor      g10210 ( new_n10587 , new_n10586 , new_n9775 );
  nor      g10211 ( new_n10588 , new_n10585 , new_n10587 );
  nand     g10212 ( new_n10589 , pi015 , pi176 );
  xor      g10213 ( new_n10590 , new_n10588 , new_n10589 );
  xor      g10214 ( new_n10591 , new_n10584 , new_n10590 );
  xor      g10215 ( new_n10592 , new_n10582 , new_n10591 );
  xor      g10216 ( new_n10593 , new_n10581 , new_n10592 );
  xor      g10217 ( new_n10594 , new_n10576 , new_n10593 );
  xor      g10218 ( new_n10595 , new_n10571 , new_n10594 );
  xor      g10219 ( new_n10596 , new_n10547 , new_n10595 );
  nand     g10220 ( new_n10597 , pi047 , pi252 );
  nand g10221 ( new_n10598 , new_n9722 , new_n9722 );
  nor      g10222 ( new_n10599 , new_n10598 , new_n9748 );
  nor      g10223 ( new_n10600 , new_n9720 , new_n9749 );
  nor      g10224 ( new_n10601 , new_n10599 , new_n10600 );
  nor      g10225 ( new_n10602 , new_n9693 , new_n9764 );
  nor      g10226 ( new_n10603 , new_n9763 , new_n9765 );
  or       g10227 ( new_n10604 , new_n10602 , new_n10603 );
  nand g10228 ( new_n10605 , new_n9843 , new_n9843 );
  nor      g10229 ( new_n10606 , new_n9574 , new_n10605 );
  nand g10230 ( new_n10607 , new_n9840 , new_n9840 );
  nor      g10231 ( new_n10608 , new_n10607 , new_n9844 );
  nor      g10232 ( new_n10609 , new_n10606 , new_n10608 );
  xor      g10233 ( new_n10610 , new_n10604 , new_n10609 );
  xor      g10234 ( new_n10611 , new_n10601 , new_n10610 );
  xor      g10235 ( new_n10612 , new_n10597 , new_n10611 );
  nand     g10236 ( new_n10613 , pi212 , pi232 );
  nand     g10237 ( new_n10614 , pi128 , pi242 );
  nand     g10238 ( new_n10615 , pi018 , pi140 );
  xnor     g10239 ( new_n10616 , new_n10614 , new_n10615 );
  nand     g10240 ( new_n10617 , new_n9742 , new_n9743 );
  nand     g10241 ( new_n10618 , new_n9652 , new_n9744 );
  nand     g10242 ( new_n10619 , new_n10617 , new_n10618 );
  xor      g10243 ( new_n10620 , new_n10616 , new_n10619 );
  xor      g10244 ( new_n10621 , new_n10613 , new_n10620 );
  nand     g10245 ( new_n10622 , pi082 , pi236 );
  nand     g10246 ( new_n10623 , new_n9760 , new_n9761 );
  nand     g10247 ( new_n10624 , new_n9691 , new_n9762 );
  nand     g10248 ( new_n10625 , new_n10623 , new_n10624 );
  xor      g10249 ( new_n10626 , new_n10622 , new_n10625 );
  nor      g10250 ( new_n10627 , new_n9731 , new_n9747 );
  nor      g10251 ( new_n10628 , new_n9730 , new_n10627 );
  nand     g10252 ( new_n10629 , pi088 , pi210 );
  xor      g10253 ( new_n10630 , new_n10628 , new_n10629 );
  xor      g10254 ( new_n10631 , new_n10626 , new_n10630 );
  xor      g10255 ( new_n10632 , new_n10621 , new_n10631 );
  nand     g10256 ( new_n10633 , new_n9734 , new_n9735 );
  nand     g10257 ( new_n10634 , new_n9662 , new_n9736 );
  nand     g10258 ( new_n10635 , new_n10633 , new_n10634 );
  nand     g10259 ( new_n10636 , pi112 , pi224 );
  nand     g10260 ( new_n10637 , pi013 , pi255 );
  xor      g10261 ( new_n10638 , new_n10636 , new_n10637 );
  xor      g10262 ( new_n10639 , new_n10635 , new_n10638 );
  xor      g10263 ( new_n10640 , new_n10632 , new_n10639 );
  xor      g10264 ( new_n10641 , new_n10612 , new_n10640 );
  nand     g10265 ( new_n10642 , pi129 , pi131 );
  nand     g10266 ( new_n10643 , pi005 , pi161 );
  nand g10267 ( new_n10644 , new_n9769 , new_n9769 );
  nor      g10268 ( new_n10645 , new_n10644 , new_n9773 );
  nor      g10269 ( new_n10646 , new_n9766 , new_n9774 );
  nor      g10270 ( new_n10647 , new_n10645 , new_n10646 );
  xor      g10271 ( new_n10648 , new_n10643 , new_n10647 );
  or       g10272 ( new_n10649 , new_n9663 , new_n9732 );
  nand     g10273 ( new_n10650 , new_n9733 , new_n9737 );
  nand     g10274 ( new_n10651 , new_n10649 , new_n10650 );
  nand     g10275 ( new_n10652 , new_n9770 , new_n9771 );
  nand     g10276 ( new_n10653 , new_n9681 , new_n9772 );
  nand     g10277 ( new_n10654 , new_n10652 , new_n10653 );
  or       g10278 ( new_n10655 , new_n9741 , new_n9745 );
  nand     g10279 ( new_n10656 , new_n9738 , new_n9746 );
  nand     g10280 ( new_n10657 , new_n10655 , new_n10656 );
  nand     g10281 ( new_n10658 , pi034 , pi217 );
  nand     g10282 ( new_n10659 , pi021 , pi241 );
  xor      g10283 ( new_n10660 , new_n10658 , new_n10659 );
  xor      g10284 ( new_n10661 , new_n10657 , new_n10660 );
  xor      g10285 ( new_n10662 , new_n10654 , new_n10661 );
  xor      g10286 ( new_n10663 , new_n10651 , new_n10662 );
  xor      g10287 ( new_n10664 , new_n10648 , new_n10663 );
  xor      g10288 ( new_n10665 , new_n10642 , new_n10664 );
  xor      g10289 ( new_n10666 , new_n10641 , new_n10665 );
  xor      g10290 ( new_n10667 , new_n10596 , new_n10666 );
  xor      g10291 ( new_n10668 , new_n10541 , new_n10667 );
  nand     g10292 ( new_n10669 , new_n9802 , new_n9803 );
  nand     g10293 ( new_n10670 , new_n9629 , new_n9804 );
  nand     g10294 ( new_n10671 , new_n10669 , new_n10670 );
  nor      g10295 ( new_n10672 , new_n9630 , new_n9800 );
  nand g10296 ( new_n10673 , new_n9801 , new_n9801 );
  nor      g10297 ( new_n10674 , new_n10673 , new_n9805 );
  nor      g10298 ( new_n10675 , new_n10672 , new_n10674 );
  xor      g10299 ( new_n10676 , new_n10671 , new_n10675 );
  nand     g10300 ( new_n10677 , pi139 , pi174 );
  nand     g10301 ( new_n10678 , pi077 , pi233 );
  nand     g10302 ( new_n10679 , pi141 , pi231 );
  nand     g10303 ( new_n10680 , pi111 , pi183 );
  xor      g10304 ( new_n10681 , new_n10679 , new_n10680 );
  nand     g10305 ( new_n10682 , pi125 , pi204 );
  nand     g10306 ( new_n10683 , pi146 , pi222 );
  nand     g10307 ( new_n10684 , pi024 , pi105 );
  xor      g10308 ( new_n10685 , new_n10683 , new_n10684 );
  xor      g10309 ( new_n10686 , new_n10682 , new_n10685 );
  nand     g10310 ( new_n10687 , pi090 , pi121 );
  nand     g10311 ( new_n10688 , new_n9824 , new_n9825 );
  nand     g10312 ( new_n10689 , new_n9573 , new_n9826 );
  nand     g10313 ( new_n10690 , new_n10688 , new_n10689 );
  nand     g10314 ( new_n10691 , pi106 , pi133 );
  xor      g10315 ( new_n10692 , new_n10690 , new_n10691 );
  xor      g10316 ( new_n10693 , new_n10687 , new_n10692 );
  xor      g10317 ( new_n10694 , new_n10686 , new_n10693 );
  xor      g10318 ( new_n10695 , new_n10681 , new_n10694 );
  nand     g10319 ( new_n10696 , pi017 , pi168 );
  nand     g10320 ( new_n10697 , pi191 , pi213 );
  nor      g10321 ( new_n10698 , new_n9827 , new_n9831 );
  and      g10322 ( new_n10699 , new_n9832 , new_n9839 );
  nor      g10323 ( new_n10700 , new_n10698 , new_n10699 );
  xor      g10324 ( new_n10701 , new_n10697 , new_n10700 );
  xor      g10325 ( new_n10702 , new_n10696 , new_n10701 );
  xor      g10326 ( new_n10703 , new_n10695 , new_n10702 );
  xor      g10327 ( new_n10704 , new_n10678 , new_n10703 );
  xor      g10328 ( new_n10705 , new_n10677 , new_n10704 );
  xor      g10329 ( new_n10706 , new_n10676 , new_n10705 );
  xor      g10330 ( new_n10707 , new_n10668 , new_n10706 );
  xor      g10331 ( po086 , new_n10538 , new_n10707 );
  xnor     g10332 ( po087 , new_n7629 , new_n7630 );
  xnor     g10333 ( po088 , new_n4918 , new_n4919 );
  xor      g10334 ( po089 , new_n3154 , new_n3178 );
  xor      g10335 ( po090 , new_n2582 , new_n2584 );
  xnor     g10336 ( po091 , new_n3504 , new_n3505 );
  xnor     g10337 ( po092 , new_n5918 , new_n5919 );
  xor      g10338 ( po093 , new_n9452 , new_n9453 );
  xnor     g10339 ( po094 , new_n920 , new_n921 );
  xor      g10340 ( po095 , new_n976 , new_n1009 );
  xor      g10341 ( po096 , new_n3510 , new_n3511 );
  nand     g10342 ( new_n10719 , pi205 , pi236 );
  nand     g10343 ( new_n10720 , pi090 , pi230 );
  nand g10344 ( new_n10721 , new_n5250 , new_n5250 );
  nor      g10345 ( new_n10722 , new_n10721 , new_n5254 );
  nor      g10346 ( new_n10723 , new_n5247 , new_n5255 );
  nor      g10347 ( new_n10724 , new_n10722 , new_n10723 );
  xor      g10348 ( new_n10725 , new_n10720 , new_n10724 );
  xor      g10349 ( new_n10726 , new_n10719 , new_n10725 );
  nand     g10350 ( new_n10727 , new_n5243 , new_n5244 );
  nand     g10351 ( new_n10728 , new_n5141 , new_n5245 );
  nand     g10352 ( new_n10729 , new_n10727 , new_n10728 );
  nor      g10353 ( new_n10730 , new_n5142 , new_n5241 );
  nor      g10354 ( new_n10731 , new_n5242 , new_n5246 );
  nor      g10355 ( new_n10732 , new_n10730 , new_n10731 );
  xor      g10356 ( new_n10733 , new_n10729 , new_n10732 );
  xor      g10357 ( new_n10734 , new_n10726 , new_n10733 );
  nand     g10358 ( new_n10735 , pi055 , pi112 );
  nand     g10359 ( new_n10736 , new_n5251 , new_n5252 );
  nand     g10360 ( new_n10737 , new_n5130 , new_n5253 );
  nand     g10361 ( new_n10738 , new_n10736 , new_n10737 );
  xor      g10362 ( new_n10739 , new_n10735 , new_n10738 );
  xor      g10363 ( new_n10740 , new_n10734 , new_n10739 );
  nand     g10364 ( new_n10741 , pi050 , pi141 );
  nand     g10365 ( new_n10742 , pi212 , pi239 );
  nand     g10366 ( new_n10743 , pi025 , pi104 );
  xor      g10367 ( new_n10744 , new_n10742 , new_n10743 );
  xor      g10368 ( new_n10745 , new_n10741 , new_n10744 );
  xor      g10369 ( new_n10746 , new_n10740 , new_n10745 );
  nor      g10370 ( new_n10747 , new_n5393 , new_n5474 );
  nor      g10371 ( new_n10748 , new_n5475 , new_n5491 );
  nor      g10372 ( new_n10749 , new_n10747 , new_n10748 );
  nand     g10373 ( new_n10750 , pi002 , pi013 );
  nand     g10374 ( new_n10751 , new_n5261 , new_n5283 );
  nand     g10375 ( new_n10752 , new_n5284 , new_n5288 );
  nand     g10376 ( new_n10753 , new_n10751 , new_n10752 );
  xor      g10377 ( new_n10754 , new_n10750 , new_n10753 );
  xor      g10378 ( new_n10755 , new_n10749 , new_n10754 );
  xor      g10379 ( new_n10756 , new_n10746 , new_n10755 );
  nand     g10380 ( new_n10757 , pi064 , pi244 );
  nand     g10381 ( new_n10758 , pi150 , pi189 );
  nand     g10382 ( new_n10759 , new_n5340 , new_n5345 );
  nand     g10383 ( new_n10760 , new_n5346 , new_n5354 );
  nand     g10384 ( new_n10761 , new_n10759 , new_n10760 );
  nand     g10385 ( new_n10762 , pi035 , pi199 );
  xnor     g10386 ( new_n10763 , new_n10761 , new_n10762 );
  xor      g10387 ( new_n10764 , new_n10758 , new_n10763 );
  nand     g10388 ( new_n10765 , new_n5466 , new_n5467 );
  nand     g10389 ( new_n10766 , new_n5424 , new_n5468 );
  nand     g10390 ( new_n10767 , new_n10765 , new_n10766 );
  nand g10391 ( new_n10768 , new_n5358 , new_n5358 );
  nand     g10392 ( new_n10769 , new_n5316 , new_n10768 );
  or       g10393 ( new_n10770 , new_n5355 , new_n5361 );
  nand     g10394 ( new_n10771 , new_n10769 , new_n10770 );
  nand     g10395 ( new_n10772 , pi146 , pi186 );
  nand     g10396 ( new_n10773 , pi132 , pi152 );
  xor      g10397 ( new_n10774 , new_n10772 , new_n10773 );
  nand     g10398 ( new_n10775 , pi037 , pi168 );
  nand g10399 ( new_n10776 , new_n5465 , new_n5465 );
  nor      g10400 ( new_n10777 , new_n10776 , new_n5469 );
  nor      g10401 ( new_n10778 , new_n5462 , new_n5470 );
  nor      g10402 ( new_n10779 , new_n10777 , new_n10778 );
  xor      g10403 ( new_n10780 , new_n10775 , new_n10779 );
  xor      g10404 ( new_n10781 , new_n10774 , new_n10780 );
  nand     g10405 ( new_n10782 , pi077 , pi196 );
  nand     g10406 ( new_n10783 , pi052 , pi184 );
  xor      g10407 ( new_n10784 , new_n10782 , new_n10783 );
  xor      g10408 ( new_n10785 , new_n10781 , new_n10784 );
  xor      g10409 ( new_n10786 , new_n10771 , new_n10785 );
  xor      g10410 ( new_n10787 , new_n10767 , new_n10786 );
  xor      g10411 ( new_n10788 , new_n10764 , new_n10787 );
  xor      g10412 ( new_n10789 , new_n10757 , new_n10788 );
  xor      g10413 ( new_n10790 , new_n10756 , new_n10789 );
  nand     g10414 ( new_n10791 , pi133 , pi221 );
  nand     g10415 ( new_n10792 , pi015 , pi211 );
  xor      g10416 ( new_n10793 , new_n10791 , new_n10792 );
  nand     g10417 ( new_n10794 , pi010 , pi131 );
  nand     g10418 ( new_n10795 , new_n5272 , new_n5273 );
  nand     g10419 ( new_n10796 , new_n5192 , new_n5274 );
  nand     g10420 ( new_n10797 , new_n10795 , new_n10796 );
  xor      g10421 ( new_n10798 , new_n10794 , new_n10797 );
  xor      g10422 ( new_n10799 , new_n10793 , new_n10798 );
  nand     g10423 ( new_n10800 , pi109 , pi128 );
  nand     g10424 ( new_n10801 , pi069 , pi084 );
  xor      g10425 ( new_n10802 , new_n10800 , new_n10801 );
  or       g10426 ( new_n10803 , new_n5435 , new_n5456 );
  nand     g10427 ( new_n10804 , new_n5457 , new_n5461 );
  nand     g10428 ( new_n10805 , new_n10803 , new_n10804 );
  nand g10429 ( new_n10806 , new_n5234 , new_n5234 );
  nor      g10430 ( new_n10807 , new_n10806 , new_n5258 );
  nor      g10431 ( new_n10808 , new_n5232 , new_n5259 );
  nor      g10432 ( new_n10809 , new_n10807 , new_n10808 );
  xor      g10433 ( new_n10810 , new_n10805 , new_n10809 );
  xor      g10434 ( new_n10811 , new_n10802 , new_n10810 );
  nand     g10435 ( new_n10812 , pi047 , pi173 );
  nand     g10436 ( new_n10813 , pi074 , pi241 );
  xor      g10437 ( new_n10814 , new_n10812 , new_n10813 );
  nand     g10438 ( new_n10815 , pi029 , pi034 );
  nand g10439 ( new_n10816 , new_n5342 , new_n5342 );
  nor      g10440 ( new_n10817 , new_n10816 , new_n5343 );
  nor      g10441 ( new_n10818 , new_n5341 , new_n5344 );
  nor      g10442 ( new_n10819 , new_n10817 , new_n10818 );
  xor      g10443 ( new_n10820 , new_n10815 , new_n10819 );
  xor      g10444 ( new_n10821 , new_n10814 , new_n10820 );
  nor      g10445 ( new_n10822 , new_n5204 , new_n5262 );
  nor      g10446 ( new_n10823 , new_n5263 , new_n5267 );
  nor      g10447 ( new_n10824 , new_n10822 , new_n10823 );
  nand     g10448 ( new_n10825 , new_n5271 , new_n5275 );
  nand     g10449 ( new_n10826 , new_n5268 , new_n5276 );
  nand     g10450 ( new_n10827 , new_n10825 , new_n10826 );
  xor      g10451 ( new_n10828 , new_n10824 , new_n10827 );
  nand     g10452 ( new_n10829 , pi161 , pi253 );
  nand     g10453 ( new_n10830 , pi058 , pi204 );
  xor      g10454 ( new_n10831 , new_n10829 , new_n10830 );
  xor      g10455 ( new_n10832 , new_n10828 , new_n10831 );
  xor      g10456 ( new_n10833 , new_n10821 , new_n10832 );
  nand     g10457 ( new_n10834 , new_n5193 , new_n5280 );
  or       g10458 ( new_n10835 , new_n5277 , new_n5282 );
  nand     g10459 ( new_n10836 , new_n10834 , new_n10835 );
  nand     g10460 ( new_n10837 , pi014 , pi018 );
  xor      g10461 ( new_n10838 , new_n10836 , new_n10837 );
  nand g10462 ( new_n10839 , new_n5451 , new_n5451 );
  nor      g10463 ( new_n10840 , new_n10839 , new_n5472 );
  nor      g10464 ( new_n10841 , new_n5449 , new_n5473 );
  nor      g10465 ( new_n10842 , new_n10840 , new_n10841 );
  nand     g10466 ( new_n10843 , pi066 , pi105 );
  nand     g10467 ( new_n10844 , pi208 , pi218 );
  nor      g10468 ( new_n10845 , new_n5327 , new_n5351 );
  nor      g10469 ( new_n10846 , new_n5350 , new_n5352 );
  nor      g10470 ( new_n10847 , new_n10845 , new_n10846 );
  xor      g10471 ( new_n10848 , new_n10844 , new_n10847 );
  xor      g10472 ( new_n10849 , new_n10843 , new_n10848 );
  xor      g10473 ( new_n10850 , new_n10842 , new_n10849 );
  and      g10474 ( new_n10851 , new_n5425 , new_n5453 );
  nor      g10475 ( new_n10852 , new_n5455 , new_n5471 );
  nor      g10476 ( new_n10853 , new_n10851 , new_n10852 );
  nand     g10477 ( new_n10854 , new_n5347 , new_n5348 );
  nand     g10478 ( new_n10855 , new_n5325 , new_n5349 );
  nand     g10479 ( new_n10856 , new_n10854 , new_n10855 );
  nand     g10480 ( new_n10857 , pi213 , pi243 );
  nand     g10481 ( new_n10858 , pi183 , pi207 );
  xor      g10482 ( new_n10859 , new_n10857 , new_n10858 );
  xor      g10483 ( new_n10860 , new_n10856 , new_n10859 );
  xor      g10484 ( new_n10861 , new_n10853 , new_n10860 );
  xor      g10485 ( new_n10862 , new_n10850 , new_n10861 );
  xor      g10486 ( new_n10863 , new_n10838 , new_n10862 );
  xor      g10487 ( new_n10864 , new_n10833 , new_n10863 );
  xor      g10488 ( new_n10865 , new_n10811 , new_n10864 );
  xor      g10489 ( new_n10866 , new_n10799 , new_n10865 );
  nand     g10490 ( new_n10867 , new_n5291 , new_n5375 );
  nand g10491 ( new_n10868 , new_n5376 , new_n5376 );
  nand     g10492 ( new_n10869 , new_n10868 , new_n5392 );
  nand     g10493 ( new_n10870 , new_n10867 , new_n10869 );
  nand     g10494 ( new_n10871 , new_n5363 , new_n5373 );
  nand     g10495 ( new_n10872 , new_n5337 , new_n5374 );
  nand     g10496 ( new_n10873 , new_n10871 , new_n10872 );
  xnor     g10497 ( new_n10874 , new_n10870 , new_n10873 );
  or       g10498 ( new_n10875 , new_n5240 , new_n5257 );
  nand     g10499 ( new_n10876 , new_n5239 , new_n10875 );
  nand     g10500 ( new_n10877 , pi139 , pi195 );
  xor      g10501 ( new_n10878 , new_n10876 , new_n10877 );
  nand     g10502 ( new_n10879 , new_n5264 , new_n5265 );
  nand     g10503 ( new_n10880 , new_n5202 , new_n5266 );
  nand     g10504 ( new_n10881 , new_n10879 , new_n10880 );
  nand g10505 ( new_n10882 , new_n5458 , new_n5458 );
  nor      g10506 ( new_n10883 , new_n10882 , new_n5459 );
  nand g10507 ( new_n10884 , new_n5434 , new_n5434 );
  nor      g10508 ( new_n10885 , new_n10884 , new_n5460 );
  nor      g10509 ( new_n10886 , new_n10883 , new_n10885 );
  xor      g10510 ( new_n10887 , new_n10881 , new_n10886 );
  nand     g10511 ( new_n10888 , pi088 , pi226 );
  nand     g10512 ( new_n10889 , new_n5260 , new_n5289 );
  nand     g10513 ( new_n10890 , new_n5229 , new_n5290 );
  nand     g10514 ( new_n10891 , new_n10889 , new_n10890 );
  xor      g10515 ( new_n10892 , new_n10888 , new_n10891 );
  xor      g10516 ( new_n10893 , new_n10887 , new_n10892 );
  xor      g10517 ( new_n10894 , new_n10878 , new_n10893 );
  xor      g10518 ( new_n10895 , new_n10874 , new_n10894 );
  xor      g10519 ( new_n10896 , new_n10866 , new_n10895 );
  xor      g10520 ( po097 , new_n10790 , new_n10896 );
  xnor     g10521 ( po098 , new_n1850 , new_n1851 );
  xnor     g10522 ( po099 , new_n7797 , new_n7894 );
  xnor     g10523 ( po100 , new_n908 , new_n909 );
  xnor     g10524 ( po101 , new_n905 , new_n906 );
  xnor     g10525 ( po102 , new_n939 , new_n965 );
  xor      g10526 ( po103 , new_n3208 , new_n3209 );
  xor      g10527 ( po104 , new_n2454 , new_n2574 );
  xnor     g10528 ( po105 , new_n4223 , new_n4235 );
  xnor     g10529 ( po106 , new_n5937 , new_n5938 );
  xor      g10530 ( po107 , new_n9455 , new_n9456 );
  xor      g10531 ( po108 , new_n4180 , new_n4225 );
  nand     g10532 ( new_n10909 , pi028 , pi107 );
  nand     g10533 ( new_n10910 , pi098 , pi228 );
  xor      g10534 ( new_n10911 , new_n10909 , new_n10910 );
  or       g10535 ( new_n10912 , new_n4628 , new_n4649 );
  nand     g10536 ( new_n10913 , new_n4650 , new_n4654 );
  nand     g10537 ( new_n10914 , new_n10912 , new_n10913 );
  nand     g10538 ( new_n10915 , new_n4344 , new_n4379 );
  nand g10539 ( new_n10916 , new_n4382 , new_n4382 );
  nand     g10540 ( new_n10917 , new_n10916 , new_n4399 );
  nand     g10541 ( new_n10918 , new_n10915 , new_n10917 );
  nor      g10542 ( new_n10919 , new_n4360 , new_n4383 );
  nor      g10543 ( new_n10920 , new_n4384 , new_n4388 );
  nor      g10544 ( new_n10921 , new_n10919 , new_n10920 );
  xor      g10545 ( new_n10922 , new_n10918 , new_n10921 );
  xor      g10546 ( new_n10923 , new_n10914 , new_n10922 );
  xor      g10547 ( new_n10924 , new_n10911 , new_n10923 );
  nand     g10548 ( new_n10925 , pi108 , pi156 );
  nand     g10549 ( new_n10926 , pi118 , pi245 );
  xor      g10550 ( new_n10927 , new_n10925 , new_n10926 );
  nand     g10551 ( new_n10928 , pi043 , pi148 );
  xor      g10552 ( new_n10929 , new_n10927 , new_n10928 );
  nand     g10553 ( new_n10930 , new_n4608 , new_n4609 );
  nand     g10554 ( new_n10931 , new_n4534 , new_n4610 );
  nand     g10555 ( new_n10932 , new_n10930 , new_n10931 );
  nand     g10556 ( new_n10933 , pi039 , pi144 );
  nand     g10557 ( new_n10934 , pi012 , pi116 );
  nor      g10558 ( new_n10935 , new_n4611 , new_n4615 );
  and      g10559 ( new_n10936 , new_n4616 , new_n4623 );
  nor      g10560 ( new_n10937 , new_n10935 , new_n10936 );
  nand     g10561 ( new_n10938 , new_n4619 , new_n4620 );
  nand     g10562 ( new_n10939 , new_n4541 , new_n4621 );
  nand     g10563 ( new_n10940 , new_n10938 , new_n10939 );
  xor      g10564 ( new_n10941 , new_n10937 , new_n10940 );
  xor      g10565 ( new_n10942 , new_n10934 , new_n10941 );
  xor      g10566 ( new_n10943 , new_n10933 , new_n10942 );
  nand     g10567 ( new_n10944 , pi046 , pi103 );
  nor      g10568 ( new_n10945 , new_n4542 , new_n4617 );
  nand g10569 ( new_n10946 , new_n4618 , new_n4618 );
  nor      g10570 ( new_n10947 , new_n10946 , new_n4622 );
  nor      g10571 ( new_n10948 , new_n10945 , new_n10947 );
  nand     g10572 ( new_n10949 , pi042 , pi063 );
  xor      g10573 ( new_n10950 , new_n10948 , new_n10949 );
  xor      g10574 ( new_n10951 , new_n10944 , new_n10950 );
  xor      g10575 ( new_n10952 , new_n10943 , new_n10951 );
  xor      g10576 ( new_n10953 , new_n10932 , new_n10952 );
  xor      g10577 ( new_n10954 , new_n10929 , new_n10953 );
  and      g10578 ( new_n10955 , new_n4499 , new_n4630 );
  nor      g10579 ( new_n10956 , new_n4632 , new_n4648 );
  nor      g10580 ( new_n10957 , new_n10955 , new_n10956 );
  nand     g10581 ( new_n10958 , pi051 , pi083 );
  xor      g10582 ( new_n10959 , new_n10957 , new_n10958 );
  xor      g10583 ( new_n10960 , new_n10954 , new_n10959 );
  xor      g10584 ( new_n10961 , new_n10924 , new_n10960 );
  nand     g10585 ( new_n10962 , pi085 , pi247 );
  nand     g10586 ( new_n10963 , new_n4627 , new_n4655 );
  nand     g10587 ( new_n10964 , new_n4656 , new_n4660 );
  nand     g10588 ( new_n10965 , new_n10963 , new_n10964 );
  xor      g10589 ( new_n10966 , new_n10962 , new_n10965 );
  xor      g10590 ( new_n10967 , new_n10961 , new_n10966 );
  nand     g10591 ( new_n10968 , new_n4666 , new_n4667 );
  nand     g10592 ( new_n10969 , new_n4579 , new_n4668 );
  nand     g10593 ( new_n10970 , new_n10968 , new_n10969 );
  nand     g10594 ( new_n10971 , pi194 , pi234 );
  nand     g10595 ( new_n10972 , pi238 , pi240 );
  nand     g10596 ( new_n10973 , new_n4390 , new_n4391 );
  nand     g10597 ( new_n10974 , new_n4343 , new_n4392 );
  nand     g10598 ( new_n10975 , new_n10973 , new_n10974 );
  xor      g10599 ( new_n10976 , new_n10972 , new_n10975 );
  xor      g10600 ( new_n10977 , new_n10971 , new_n10976 );
  nand     g10601 ( new_n10978 , pi162 , pi203 );
  nand     g10602 ( new_n10979 , pi080 , pi180 );
  xor      g10603 ( new_n10980 , new_n10978 , new_n10979 );
  xor      g10604 ( new_n10981 , new_n10977 , new_n10980 );
  xor      g10605 ( new_n10982 , new_n10970 , new_n10981 );
  nor      g10606 ( new_n10983 , new_n4661 , new_n4692 );
  nor      g10607 ( new_n10984 , new_n4693 , new_n4696 );
  nor      g10608 ( new_n10985 , new_n10983 , new_n10984 );
  nor      g10609 ( new_n10986 , new_n4642 , new_n4646 );
  nand g10610 ( new_n10987 , new_n4647 , new_n4647 );
  nor      g10611 ( new_n10988 , new_n4639 , new_n10987 );
  nor      g10612 ( new_n10989 , new_n10986 , new_n10988 );
  xor      g10613 ( new_n10990 , new_n10985 , new_n10989 );
  nor      g10614 ( new_n10991 , new_n4565 , new_n4675 );
  nor      g10615 ( new_n10992 , new_n4674 , new_n4676 );
  nor      g10616 ( new_n10993 , new_n10991 , new_n10992 );
  xor      g10617 ( new_n10994 , new_n10990 , new_n10993 );
  xor      g10618 ( new_n10995 , new_n10982 , new_n10994 );
  xor      g10619 ( new_n10996 , new_n10967 , new_n10995 );
  nand     g10620 ( new_n10997 , new_n4643 , new_n4644 );
  nand     g10621 ( new_n10998 , new_n4498 , new_n4645 );
  nand     g10622 ( new_n10999 , new_n10997 , new_n10998 );
  nand     g10623 ( new_n11000 , new_n4635 , new_n4636 );
  nand     g10624 ( new_n11001 , new_n4508 , new_n4637 );
  nand     g10625 ( new_n11002 , new_n11000 , new_n11001 );
  xor      g10626 ( new_n11003 , new_n10999 , new_n11002 );
  nand     g10627 ( new_n11004 , new_n4393 , new_n4397 );
  nand g10628 ( new_n11005 , new_n4389 , new_n4389 );
  nand     g10629 ( new_n11006 , new_n11005 , new_n4398 );
  nand     g10630 ( new_n11007 , new_n11004 , new_n11006 );
  nand     g10631 ( new_n11008 , pi061 , pi070 );
  nand     g10632 ( new_n11009 , pi000 , pi188 );
  nand     g10633 ( new_n11010 , pi149 , pi237 );
  xor      g10634 ( new_n11011 , new_n11009 , new_n11010 );
  xor      g10635 ( new_n11012 , new_n11008 , new_n11011 );
  xor      g10636 ( new_n11013 , new_n11007 , new_n11012 );
  nand     g10637 ( new_n11014 , new_n4671 , new_n4672 );
  nand     g10638 ( new_n11015 , new_n4563 , new_n4673 );
  nand     g10639 ( new_n11016 , new_n11014 , new_n11015 );
  nand     g10640 ( new_n11017 , pi134 , pi193 );
  xor      g10641 ( new_n11018 , new_n11016 , new_n11017 );
  xor      g10642 ( new_n11019 , new_n11013 , new_n11018 );
  xor      g10643 ( new_n11020 , new_n11003 , new_n11019 );
  nand g10644 ( new_n11021 , new_n4377 , new_n4377 );
  nor      g10645 ( new_n11022 , new_n11021 , new_n4400 );
  nor      g10646 ( new_n11023 , new_n4376 , new_n4401 );
  or       g10647 ( new_n11024 , new_n11022 , new_n11023 );
  nor      g10648 ( new_n11025 , new_n4402 , new_n4597 );
  nor      g10649 ( new_n11026 , new_n4598 , new_n4697 );
  nor      g10650 ( new_n11027 , new_n11025 , new_n11026 );
  xor      g10651 ( new_n11028 , new_n11024 , new_n11027 );
  xor      g10652 ( new_n11029 , new_n11020 , new_n11028 );
  nand     g10653 ( new_n11030 , new_n4685 , new_n4691 );
  nand     g10654 ( new_n11031 , new_n4686 , new_n11030 );
  nand     g10655 ( new_n11032 , pi007 , pi201 );
  nand     g10656 ( new_n11033 , pi049 , pi113 );
  xor      g10657 ( new_n11034 , new_n11032 , new_n11033 );
  nand     g10658 ( new_n11035 , pi038 , pi171 );
  nand     g10659 ( new_n11036 , pi143 , pi202 );
  nand     g10660 ( new_n11037 , pi159 , pi175 );
  xor      g10661 ( new_n11038 , new_n11036 , new_n11037 );
  xor      g10662 ( new_n11039 , new_n11035 , new_n11038 );
  xor      g10663 ( new_n11040 , new_n11034 , new_n11039 );
  nand     g10664 ( new_n11041 , pi115 , pi178 );
  nand     g10665 ( new_n11042 , pi126 , pi163 );
  nand     g10666 ( new_n11043 , pi033 , pi200 );
  xor      g10667 ( new_n11044 , new_n11042 , new_n11043 );
  xor      g10668 ( new_n11045 , new_n11041 , new_n11044 );
  xor      g10669 ( new_n11046 , new_n11040 , new_n11045 );
  xor      g10670 ( new_n11047 , new_n11031 , new_n11046 );
  xor      g10671 ( new_n11048 , new_n11029 , new_n11047 );
  nand     g10672 ( new_n11049 , new_n4603 , new_n4625 );
  nand g10673 ( new_n11050 , new_n4601 , new_n4601 );
  nand     g10674 ( new_n11051 , new_n11050 , new_n4626 );
  nand     g10675 ( new_n11052 , new_n11049 , new_n11051 );
  nand     g10676 ( new_n11053 , pi016 , pi036 );
  nor      g10677 ( new_n11054 , new_n4510 , new_n4633 );
  nor      g10678 ( new_n11055 , new_n4634 , new_n4638 );
  nor      g10679 ( new_n11056 , new_n11054 , new_n11055 );
  xor      g10680 ( new_n11057 , new_n11053 , new_n11056 );
  xor      g10681 ( new_n11058 , new_n11052 , new_n11057 );
  nand     g10682 ( new_n11059 , pi057 , pi214 );
  and      g10683 ( new_n11060 , new_n4535 , new_n4605 );
  nor      g10684 ( new_n11061 , new_n4607 , new_n4624 );
  nor      g10685 ( new_n11062 , new_n11060 , new_n11061 );
  xor      g10686 ( new_n11063 , new_n11059 , new_n11062 );
  nand     g10687 ( new_n11064 , pi068 , pi117 );
  nand     g10688 ( new_n11065 , pi179 , pi181 );
  xor      g10689 ( new_n11066 , new_n11064 , new_n11065 );
  nand     g10690 ( new_n11067 , new_n4665 , new_n4669 );
  nand     g10691 ( new_n11068 , new_n4670 , new_n4677 );
  nand     g10692 ( new_n11069 , new_n11067 , new_n11068 );
  and      g10693 ( new_n11070 , new_n4580 , new_n4681 );
  nor      g10694 ( new_n11071 , new_n4678 , new_n4683 );
  nor      g10695 ( new_n11072 , new_n11070 , new_n11071 );
  xor      g10696 ( new_n11073 , new_n11069 , new_n11072 );
  nand     g10697 ( new_n11074 , pi048 , pi167 );
  nand     g10698 ( new_n11075 , new_n4385 , new_n4386 );
  nand     g10699 ( new_n11076 , new_n4358 , new_n4387 );
  nand     g10700 ( new_n11077 , new_n11075 , new_n11076 );
  xor      g10701 ( new_n11078 , new_n11074 , new_n11077 );
  xor      g10702 ( new_n11079 , new_n11073 , new_n11078 );
  xor      g10703 ( new_n11080 , new_n11066 , new_n11079 );
  xor      g10704 ( new_n11081 , new_n11063 , new_n11080 );
  xor      g10705 ( new_n11082 , new_n11058 , new_n11081 );
  xor      g10706 ( new_n11083 , new_n11048 , new_n11082 );
  xor      g10707 ( po109 , new_n10996 , new_n11083 );
  xor      g10708 ( po110 , new_n4950 , new_n4965 );
  xor      g10709 ( po111 , new_n3197 , new_n3199 );
  xor      g10710 ( po112 , new_n8148 , new_n8149 );
  xnor     g10711 ( po113 , new_n8153 , new_n8206 );
  xnor     g10712 ( po114 , new_n8672 , new_n8673 );
  xnor     g10713 ( po115 , new_n7218 , new_n7219 );
  xor      g10714 ( po116 , new_n9449 , new_n9450 );
  xor      g10715 ( po117 , new_n9710 , new_n9711 );
  xor      g10716 ( po118 , new_n8675 , new_n8676 );
  xnor     g10717 ( po119 , new_n4485 , new_n4595 );
endmodule


