 module top_809960632_810038711_1598227639_893650103 (a, b, o);

      input a, b; output o; nor_6 g0(a,b,o); endmodule