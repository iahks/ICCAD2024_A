 module top_809568696_809776567_809698999_863110837_1234615 (a, o);

      input a, b; output o; buf_7 g0(a,o); endmodule