// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Wed Aug 14 19:23:49 2024

module top_810026173_826291639_946996917_1246901 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83,
    pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81,
    pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181;
  wire new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n908, new_n910, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1161,
    new_n1162, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211, new_n1213, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1426, new_n1428, new_n1430, new_n1431, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1468, new_n1470, new_n1471, new_n1472, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1483, new_n1484,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1497,
    new_n1498, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1518,
    new_n1520, new_n1522, new_n1527, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1537, new_n1542, new_n1546, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556, new_n1559,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1567, new_n1568,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1579,
    new_n1587, new_n1592, new_n1599, new_n1602, new_n1604, new_n1605,
    new_n1611, new_n1617, new_n1618, new_n1621, new_n1624, new_n1625,
    new_n1631, new_n1636, new_n1640, new_n1645, new_n1649;
  not_8  g0000(.A(pi25), .Y(new_n276));
  nand_5 g0001(.A(pi85), .B(pi03), .Y(new_n277));
  or_6   g0002(.A(pi85), .B(pi03), .Y(new_n278));
  nand_5 g0003(.A(pi47), .B(pi30), .Y(new_n279));
  xor_4  g0004(.A(pi47), .B(pi30), .Y(new_n280));
  nand_5 g0005(.A(pi45), .B(pi19), .Y(new_n281));
  xor_4  g0006(.A(pi45), .B(pi19), .Y(new_n282));
  or_6   g0007(.A(pi56), .B(pi17), .Y(new_n283));
  xor_4  g0008(.A(pi56), .B(pi17), .Y(new_n284));
  nand_5 g0009(.A(pi63), .B(pi55), .Y(new_n285));
  nand_5 g0010(.A(new_n285), .B(new_n284), .Y(new_n286));
  nand_5 g0011(.A(new_n286), .B(new_n283), .Y(new_n287));
  not_8  g0012(.A(new_n287), .Y(new_n288));
  nand_5 g0013(.A(new_n288), .B(new_n282), .Y(new_n289));
  nand_5 g0014(.A(new_n289), .B(new_n281), .Y(new_n290));
  nand_5 g0015(.A(new_n290), .B(new_n280), .Y(new_n291));
  nand_5 g0016(.A(new_n291), .B(new_n279), .Y(new_n292));
  nand_5 g0017(.A(new_n292), .B(new_n278), .Y(new_n293));
  nand_5 g0018(.A(new_n293), .B(new_n277), .Y(new_n294));
  nand_5 g0019(.A(new_n294), .B(pi77), .Y(new_n295));
  xor_4  g0020(.A(new_n295), .B(new_n276), .Y(new_n296));
  not_8  g0021(.A(new_n296), .Y(new_n297));
  not_8  g0022(.A(pi39), .Y(new_n298));
  not_8  g0023(.A(pi60), .Y(new_n299));
  nand_5 g0024(.A(new_n299), .B(new_n298), .Y(new_n300));
  or_6   g0025(.A(pi86), .B(new_n299), .Y(new_n301));
  nand_5 g0026(.A(new_n301), .B(new_n300), .Y(new_n302));
  nand_5 g0027(.A(pi60), .B(pi51), .Y(new_n303));
  nand_5 g0028(.A(new_n299), .B(pi06), .Y(new_n304));
  nand_5 g0029(.A(new_n304), .B(new_n303), .Y(new_n305));
  nand_5 g0030(.A(new_n305), .B(pi41), .Y(new_n306));
  xor_4  g0031(.A(new_n305), .B(pi41), .Y(new_n307));
  nand_5 g0032(.A(pi76), .B(pi60), .Y(new_n308));
  nand_5 g0033(.A(new_n299), .B(pi18), .Y(new_n309));
  nand_5 g0034(.A(new_n309), .B(new_n308), .Y(new_n310));
  nand_5 g0035(.A(new_n310), .B(pi79), .Y(new_n311));
  not_8  g0036(.A(new_n311), .Y(new_n312));
  not_8  g0037(.A(pi91), .Y(new_n313));
  nand_5 g0038(.A(pi60), .B(pi32), .Y(new_n314));
  nand_5 g0039(.A(new_n299), .B(pi59), .Y(new_n315));
  nand_5 g0040(.A(new_n315), .B(new_n314), .Y(new_n316));
  not_8  g0041(.A(new_n316), .Y(new_n317));
  nand_5 g0042(.A(new_n317), .B(new_n313), .Y(new_n318));
  nor_5  g0043(.A(new_n318), .B(new_n312), .Y(new_n319));
  nor_5  g0044(.A(new_n317), .B(new_n313), .Y(new_n320));
  and_6  g0045(.A(new_n320), .B(new_n312), .Y(new_n321));
  or_6   g0046(.A(new_n321), .B(new_n319), .Y(new_n322));
  nand_5 g0047(.A(new_n322), .B(new_n307), .Y(new_n323));
  nand_5 g0048(.A(new_n323), .B(new_n306), .Y(new_n324));
  nand_5 g0049(.A(pi60), .B(pi08), .Y(new_n325));
  nand_5 g0050(.A(pi75), .B(new_n299), .Y(new_n326));
  nand_5 g0051(.A(new_n326), .B(new_n325), .Y(new_n327));
  not_8  g0052(.A(new_n327), .Y(new_n328));
  nand_5 g0053(.A(new_n328), .B(new_n319), .Y(new_n329));
  nor_5  g0054(.A(new_n329), .B(new_n324), .Y(new_n330));
  nor_5  g0055(.A(new_n330), .B(new_n302), .Y(new_n331));
  nor_5  g0056(.A(new_n328), .B(new_n319), .Y(new_n332));
  nand_5 g0057(.A(new_n332), .B(new_n324), .Y(new_n333));
  nand_5 g0058(.A(new_n333), .B(new_n302), .Y(new_n334));
  nand_5 g0059(.A(pi60), .B(pi34), .Y(new_n335));
  not_8  g0060(.A(pi82), .Y(new_n336));
  nand_5 g0061(.A(new_n336), .B(new_n299), .Y(new_n337));
  nand_5 g0062(.A(new_n337), .B(new_n335), .Y(new_n338));
  nand_5 g0063(.A(new_n338), .B(new_n334), .Y(new_n339));
  nor_5  g0064(.A(new_n339), .B(new_n331), .Y(new_n340));
  nand_5 g0065(.A(new_n336), .B(new_n298), .Y(new_n341));
  xor_4  g0066(.A(new_n341), .B(pi04), .Y(new_n342));
  nor_5  g0067(.A(new_n342), .B(pi60), .Y(new_n343));
  not_8  g0068(.A(pi02), .Y(new_n344));
  nand_5 g0069(.A(pi86), .B(pi34), .Y(new_n345));
  nand_5 g0070(.A(new_n345), .B(new_n344), .Y(new_n346));
  not_8  g0071(.A(new_n346), .Y(new_n347));
  nor_5  g0072(.A(new_n345), .B(new_n344), .Y(new_n348));
  not_8  g0073(.A(new_n348), .Y(new_n349));
  nand_5 g0074(.A(new_n349), .B(pi60), .Y(new_n350));
  nor_5  g0075(.A(new_n350), .B(new_n347), .Y(new_n351));
  nor_5  g0076(.A(new_n351), .B(new_n343), .Y(new_n352));
  xor_4  g0077(.A(new_n352), .B(new_n340), .Y(new_n353));
  xor_4  g0078(.A(new_n353), .B(new_n297), .Y(new_n354));
  xor_4  g0079(.A(new_n294), .B(pi77), .Y(new_n355));
  not_8  g0080(.A(new_n355), .Y(new_n356));
  not_8  g0081(.A(new_n330), .Y(new_n357));
  nand_5 g0082(.A(new_n334), .B(new_n357), .Y(new_n358));
  xor_4  g0083(.A(new_n358), .B(new_n338), .Y(new_n359));
  nand_5 g0084(.A(new_n359), .B(new_n356), .Y(new_n360));
  not_8  g0085(.A(new_n360), .Y(new_n361));
  nand_5 g0086(.A(new_n278), .B(new_n277), .Y(new_n362));
  xor_4  g0087(.A(new_n362), .B(new_n292), .Y(new_n363));
  not_8  g0088(.A(new_n363), .Y(new_n364));
  nand_5 g0089(.A(new_n333), .B(new_n357), .Y(new_n365));
  xor_4  g0090(.A(new_n365), .B(new_n302), .Y(new_n366));
  nand_5 g0091(.A(new_n366), .B(new_n364), .Y(new_n367));
  xor_4  g0092(.A(new_n290), .B(new_n280), .Y(new_n368));
  not_8  g0093(.A(new_n368), .Y(new_n369));
  xor_4  g0094(.A(new_n288), .B(new_n282), .Y(new_n370));
  not_8  g0095(.A(new_n370), .Y(new_n371));
  xor_4  g0096(.A(new_n316), .B(new_n313), .Y(new_n372));
  nand_5 g0097(.A(new_n372), .B(new_n312), .Y(new_n373));
  xor_4  g0098(.A(new_n285), .B(new_n284), .Y(new_n374));
  not_8  g0099(.A(new_n374), .Y(new_n375));
  nand_5 g0100(.A(new_n375), .B(new_n372), .Y(new_n376));
  xor_4  g0101(.A(new_n375), .B(new_n372), .Y(new_n377));
  or_6   g0102(.A(pi63), .B(pi55), .Y(new_n378));
  nand_5 g0103(.A(new_n378), .B(new_n285), .Y(new_n379));
  not_8  g0104(.A(new_n379), .Y(new_n380));
  xor_4  g0105(.A(new_n310), .B(pi79), .Y(new_n381));
  nand_5 g0106(.A(new_n381), .B(new_n380), .Y(new_n382));
  nand_5 g0107(.A(new_n382), .B(new_n311), .Y(new_n383));
  nand_5 g0108(.A(new_n383), .B(new_n377), .Y(new_n384));
  nand_5 g0109(.A(new_n384), .B(new_n376), .Y(new_n385));
  nand_5 g0110(.A(new_n385), .B(new_n373), .Y(new_n386));
  nand_5 g0111(.A(new_n386), .B(new_n371), .Y(new_n387));
  xor_4  g0112(.A(new_n322), .B(new_n307), .Y(new_n388));
  xor_4  g0113(.A(new_n386), .B(new_n370), .Y(new_n389));
  or_6   g0114(.A(new_n389), .B(new_n388), .Y(new_n390));
  nand_5 g0115(.A(new_n390), .B(new_n387), .Y(new_n391));
  nand_5 g0116(.A(new_n391), .B(new_n369), .Y(new_n392));
  xor_4  g0117(.A(new_n391), .B(new_n368), .Y(new_n393));
  xor_4  g0118(.A(new_n328), .B(new_n319), .Y(new_n394));
  xor_4  g0119(.A(new_n394), .B(new_n324), .Y(new_n395));
  not_8  g0120(.A(new_n395), .Y(new_n396));
  or_6   g0121(.A(new_n396), .B(new_n393), .Y(new_n397));
  nand_5 g0122(.A(new_n397), .B(new_n392), .Y(new_n398));
  xor_4  g0123(.A(new_n366), .B(new_n363), .Y(new_n399));
  or_6   g0124(.A(new_n399), .B(new_n398), .Y(new_n400));
  nand_5 g0125(.A(new_n400), .B(new_n367), .Y(new_n401));
  xor_4  g0126(.A(new_n359), .B(new_n355), .Y(new_n402));
  nor_5  g0127(.A(new_n402), .B(new_n401), .Y(new_n403));
  nor_5  g0128(.A(new_n403), .B(new_n361), .Y(new_n404));
  xor_4  g0129(.A(new_n404), .B(new_n354), .Y(po000));
  not_8  g0130(.A(pi73), .Y(new_n406));
  nand_5 g0131(.A(new_n406), .B(pi22), .Y(new_n407));
  nand_5 g0132(.A(new_n407), .B(pi76), .Y(new_n408));
  not_8  g0133(.A(new_n407), .Y(new_n409));
  nand_5 g0134(.A(new_n409), .B(pi18), .Y(new_n410));
  nand_5 g0135(.A(new_n410), .B(new_n408), .Y(new_n411));
  xor_4  g0136(.A(new_n411), .B(pi16), .Y(new_n412));
  nand_5 g0137(.A(new_n412), .B(new_n380), .Y(new_n413));
  nand_5 g0138(.A(new_n413), .B(new_n374), .Y(new_n414));
  nand_5 g0139(.A(new_n411), .B(pi16), .Y(new_n415));
  nand_5 g0140(.A(new_n407), .B(pi32), .Y(new_n416));
  nand_5 g0141(.A(new_n409), .B(pi59), .Y(new_n417));
  nand_5 g0142(.A(new_n417), .B(new_n416), .Y(new_n418));
  xor_4  g0143(.A(new_n418), .B(pi57), .Y(new_n419));
  xor_4  g0144(.A(new_n419), .B(new_n415), .Y(new_n420));
  not_8  g0145(.A(new_n420), .Y(new_n421));
  not_8  g0146(.A(new_n412), .Y(new_n422));
  nand_5 g0147(.A(new_n378), .B(new_n284), .Y(new_n423));
  nor_5  g0148(.A(new_n423), .B(new_n422), .Y(new_n424));
  or_6   g0149(.A(new_n424), .B(new_n421), .Y(new_n425));
  nand_5 g0150(.A(new_n425), .B(new_n414), .Y(new_n426));
  xor_4  g0151(.A(new_n426), .B(new_n371), .Y(new_n427));
  nand_5 g0152(.A(new_n407), .B(pi51), .Y(new_n428));
  nand_5 g0153(.A(new_n409), .B(pi06), .Y(new_n429));
  nand_5 g0154(.A(new_n429), .B(new_n428), .Y(new_n430));
  xor_4  g0155(.A(new_n430), .B(pi07), .Y(new_n431));
  not_8  g0156(.A(new_n431), .Y(new_n432));
  nand_5 g0157(.A(new_n418), .B(pi57), .Y(new_n433));
  not_8  g0158(.A(new_n415), .Y(new_n434));
  nand_5 g0159(.A(new_n419), .B(new_n434), .Y(new_n435));
  nand_5 g0160(.A(new_n435), .B(new_n433), .Y(new_n436));
  xor_4  g0161(.A(new_n436), .B(new_n432), .Y(new_n437));
  not_8  g0162(.A(new_n437), .Y(new_n438));
  xor_4  g0163(.A(new_n438), .B(new_n427), .Y(po001));
  not_8  g0164(.A(pi04), .Y(new_n440));
  not_8  g0165(.A(pi78), .Y(new_n441));
  nand_5 g0166(.A(new_n441), .B(new_n440), .Y(new_n442));
  xor_4  g0167(.A(new_n442), .B(pi20), .Y(new_n443));
  nor_5  g0168(.A(new_n443), .B(new_n407), .Y(new_n444));
  not_8  g0169(.A(pi84), .Y(new_n445));
  not_8  g0170(.A(pi13), .Y(new_n446));
  not_8  g0171(.A(pi34), .Y(new_n447));
  nand_5 g0172(.A(new_n447), .B(new_n344), .Y(new_n448));
  nor_5  g0173(.A(new_n448), .B(new_n406), .Y(new_n449));
  nand_5 g0174(.A(new_n449), .B(new_n446), .Y(new_n450));
  not_8  g0175(.A(new_n450), .Y(new_n451));
  nand_5 g0176(.A(new_n451), .B(new_n445), .Y(new_n452));
  nor_5  g0177(.A(new_n409), .B(new_n445), .Y(new_n453));
  nand_5 g0178(.A(new_n453), .B(new_n450), .Y(new_n454));
  nand_5 g0179(.A(new_n454), .B(new_n452), .Y(new_n455));
  nor_5  g0180(.A(new_n455), .B(new_n444), .Y(new_n456));
  not_8  g0181(.A(new_n442), .Y(new_n457));
  nand_5 g0182(.A(pi78), .B(pi04), .Y(new_n458));
  nand_5 g0183(.A(new_n458), .B(new_n409), .Y(new_n459));
  nor_5  g0184(.A(new_n459), .B(new_n457), .Y(new_n460));
  nand_5 g0185(.A(new_n407), .B(new_n446), .Y(new_n461));
  not_8  g0186(.A(new_n461), .Y(new_n462));
  nor_5  g0187(.A(new_n462), .B(new_n449), .Y(new_n463));
  not_8  g0188(.A(new_n463), .Y(new_n464));
  nor_5  g0189(.A(new_n464), .B(new_n460), .Y(new_n465));
  nor_5  g0190(.A(new_n465), .B(new_n451), .Y(new_n466));
  not_8  g0191(.A(new_n466), .Y(new_n467));
  xor_4  g0192(.A(pi34), .B(pi02), .Y(new_n468));
  or_6   g0193(.A(new_n468), .B(new_n406), .Y(new_n469));
  not_8  g0194(.A(new_n469), .Y(new_n470));
  nand_5 g0195(.A(new_n409), .B(new_n440), .Y(new_n471));
  nor_5  g0196(.A(pi73), .B(pi22), .Y(new_n472));
  nand_5 g0197(.A(new_n472), .B(pi02), .Y(new_n473));
  nand_5 g0198(.A(new_n473), .B(new_n471), .Y(new_n474));
  nor_5  g0199(.A(new_n474), .B(new_n470), .Y(new_n475));
  nand_5 g0200(.A(new_n409), .B(new_n336), .Y(new_n476));
  not_8  g0201(.A(new_n476), .Y(new_n477));
  nand_5 g0202(.A(new_n472), .B(new_n447), .Y(new_n478));
  nand_5 g0203(.A(pi73), .B(pi34), .Y(new_n479));
  nand_5 g0204(.A(new_n479), .B(new_n478), .Y(new_n480));
  nor_5  g0205(.A(new_n480), .B(new_n477), .Y(new_n481));
  not_8  g0206(.A(new_n481), .Y(new_n482));
  not_8  g0207(.A(pi85), .Y(new_n483));
  nand_5 g0208(.A(new_n407), .B(pi86), .Y(new_n484));
  nand_5 g0209(.A(new_n409), .B(pi39), .Y(new_n485));
  nand_5 g0210(.A(new_n485), .B(new_n484), .Y(new_n486));
  not_8  g0211(.A(new_n486), .Y(new_n487));
  nand_5 g0212(.A(new_n487), .B(new_n483), .Y(new_n488));
  xor_4  g0213(.A(new_n486), .B(pi85), .Y(new_n489));
  nand_5 g0214(.A(new_n407), .B(pi08), .Y(new_n490));
  nand_5 g0215(.A(new_n409), .B(pi75), .Y(new_n491));
  nand_5 g0216(.A(new_n491), .B(new_n490), .Y(new_n492));
  and_6  g0217(.A(new_n492), .B(pi30), .Y(new_n493));
  or_6   g0218(.A(new_n430), .B(pi19), .Y(new_n494));
  or_6   g0219(.A(new_n418), .B(pi56), .Y(new_n495));
  nand_5 g0220(.A(new_n411), .B(pi63), .Y(new_n496));
  nand_5 g0221(.A(new_n418), .B(pi56), .Y(new_n497));
  nand_5 g0222(.A(new_n497), .B(new_n495), .Y(new_n498));
  not_8  g0223(.A(new_n498), .Y(new_n499));
  nand_5 g0224(.A(new_n499), .B(new_n496), .Y(new_n500));
  nand_5 g0225(.A(new_n500), .B(new_n495), .Y(new_n501));
  xor_4  g0226(.A(new_n430), .B(pi19), .Y(new_n502));
  nand_5 g0227(.A(new_n502), .B(new_n501), .Y(new_n503));
  nand_5 g0228(.A(new_n503), .B(new_n494), .Y(new_n504));
  not_8  g0229(.A(pi30), .Y(new_n505));
  xor_4  g0230(.A(new_n492), .B(new_n505), .Y(new_n506));
  nor_5  g0231(.A(new_n506), .B(new_n504), .Y(new_n507));
  nor_5  g0232(.A(new_n507), .B(new_n493), .Y(new_n508));
  nand_5 g0233(.A(new_n508), .B(new_n489), .Y(new_n509));
  nand_5 g0234(.A(new_n509), .B(new_n488), .Y(new_n510));
  nand_5 g0235(.A(new_n510), .B(new_n482), .Y(new_n511));
  nor_5  g0236(.A(new_n510), .B(new_n482), .Y(new_n512));
  not_8  g0237(.A(new_n512), .Y(new_n513));
  xor_4  g0238(.A(new_n508), .B(new_n489), .Y(new_n514));
  xor_4  g0239(.A(new_n502), .B(new_n501), .Y(new_n515));
  nor_5  g0240(.A(new_n411), .B(pi63), .Y(new_n516));
  nand_5 g0241(.A(new_n516), .B(new_n495), .Y(new_n517));
  not_8  g0242(.A(new_n516), .Y(new_n518));
  nand_5 g0243(.A(new_n518), .B(new_n497), .Y(new_n519));
  nand_5 g0244(.A(new_n519), .B(new_n517), .Y(new_n520));
  xnor_4 g0245(.A(new_n520), .B(new_n502), .Y(po053));
  nand_5 g0246(.A(po053), .B(new_n515), .Y(new_n522));
  xor_4  g0247(.A(new_n506), .B(new_n504), .Y(po176));
  nor_5  g0248(.A(po176), .B(new_n522), .Y(new_n524));
  or_6   g0249(.A(new_n524), .B(new_n514), .Y(new_n525));
  nand_5 g0250(.A(new_n525), .B(new_n513), .Y(new_n526));
  nand_5 g0251(.A(new_n526), .B(new_n511), .Y(new_n527));
  nor_5  g0252(.A(new_n527), .B(new_n475), .Y(new_n528));
  nand_5 g0253(.A(new_n528), .B(new_n467), .Y(new_n529));
  xor_4  g0254(.A(new_n529), .B(new_n456), .Y(po002));
  xor_4  g0255(.A(new_n381), .B(new_n380), .Y(po003));
  not_8  g0256(.A(pi14), .Y(new_n532));
  xor_4  g0257(.A(pi86), .B(pi34), .Y(new_n533));
  nor_5  g0258(.A(new_n533), .B(new_n532), .Y(new_n534));
  nand_5 g0259(.A(pi82), .B(pi39), .Y(new_n535));
  not_8  g0260(.A(new_n535), .Y(new_n536));
  nand_5 g0261(.A(new_n341), .B(new_n532), .Y(new_n537));
  nor_5  g0262(.A(new_n537), .B(new_n536), .Y(new_n538));
  nor_5  g0263(.A(new_n538), .B(new_n534), .Y(new_n539));
  nand_5 g0264(.A(pi86), .B(pi14), .Y(new_n540));
  nand_5 g0265(.A(pi39), .B(new_n532), .Y(new_n541));
  nand_5 g0266(.A(new_n541), .B(new_n540), .Y(new_n542));
  not_8  g0267(.A(new_n542), .Y(new_n543));
  nand_5 g0268(.A(pi14), .B(pi08), .Y(new_n544));
  nand_5 g0269(.A(pi75), .B(new_n532), .Y(new_n545));
  nand_5 g0270(.A(new_n545), .B(new_n544), .Y(new_n546));
  nand_5 g0271(.A(new_n546), .B(pi12), .Y(new_n547));
  nor_5  g0272(.A(new_n546), .B(pi12), .Y(new_n548));
  nand_5 g0273(.A(pi32), .B(pi14), .Y(new_n549));
  nand_5 g0274(.A(pi59), .B(new_n532), .Y(new_n550));
  nand_5 g0275(.A(new_n550), .B(new_n549), .Y(new_n551));
  nand_5 g0276(.A(new_n551), .B(pi28), .Y(new_n552));
  not_8  g0277(.A(new_n552), .Y(new_n553));
  nand_5 g0278(.A(pi51), .B(pi14), .Y(new_n554));
  nand_5 g0279(.A(new_n532), .B(pi06), .Y(new_n555));
  nand_5 g0280(.A(new_n555), .B(new_n554), .Y(new_n556));
  or_6   g0281(.A(new_n556), .B(pi26), .Y(new_n557));
  nor_5  g0282(.A(new_n557), .B(new_n553), .Y(new_n558));
  nand_5 g0283(.A(new_n556), .B(pi26), .Y(new_n559));
  nor_5  g0284(.A(new_n559), .B(new_n552), .Y(new_n560));
  nor_5  g0285(.A(new_n560), .B(new_n558), .Y(new_n561));
  or_6   g0286(.A(new_n561), .B(new_n548), .Y(new_n562));
  nand_5 g0287(.A(new_n562), .B(new_n547), .Y(new_n563));
  nor_5  g0288(.A(new_n563), .B(new_n543), .Y(new_n564));
  not_8  g0289(.A(new_n548), .Y(new_n565));
  nand_5 g0290(.A(new_n558), .B(new_n565), .Y(new_n566));
  not_8  g0291(.A(new_n566), .Y(new_n567));
  nor_5  g0292(.A(new_n558), .B(new_n542), .Y(new_n568));
  nor_5  g0293(.A(new_n568), .B(new_n567), .Y(new_n569));
  not_8  g0294(.A(new_n569), .Y(new_n570));
  nor_5  g0295(.A(new_n570), .B(new_n564), .Y(new_n571));
  not_8  g0296(.A(new_n571), .Y(new_n572));
  nor_5  g0297(.A(new_n572), .B(new_n539), .Y(new_n573));
  not_8  g0298(.A(new_n573), .Y(new_n574));
  nand_5 g0299(.A(new_n468), .B(pi14), .Y(new_n575));
  nand_5 g0300(.A(new_n532), .B(pi04), .Y(new_n576));
  nand_5 g0301(.A(new_n576), .B(new_n575), .Y(new_n577));
  nor_5  g0302(.A(new_n577), .B(new_n574), .Y(new_n578));
  nand_5 g0303(.A(new_n441), .B(new_n532), .Y(new_n579));
  nand_5 g0304(.A(new_n336), .B(new_n532), .Y(new_n580));
  not_8  g0305(.A(new_n580), .Y(new_n581));
  nand_5 g0306(.A(new_n581), .B(new_n440), .Y(new_n582));
  nand_5 g0307(.A(new_n582), .B(new_n579), .Y(new_n583));
  nand_5 g0308(.A(new_n457), .B(new_n336), .Y(new_n584));
  nand_5 g0309(.A(new_n584), .B(new_n583), .Y(new_n585));
  nand_5 g0310(.A(pi14), .B(new_n446), .Y(new_n586));
  nand_5 g0311(.A(new_n586), .B(new_n585), .Y(new_n587));
  not_8  g0312(.A(new_n587), .Y(new_n588));
  xor_4  g0313(.A(new_n588), .B(new_n578), .Y(new_n589));
  xor_4  g0314(.A(new_n589), .B(pi81), .Y(new_n590));
  nand_5 g0315(.A(pi14), .B(pi02), .Y(new_n591));
  not_8  g0316(.A(new_n582), .Y(new_n592));
  nor_5  g0317(.A(new_n576), .B(new_n336), .Y(new_n593));
  nor_5  g0318(.A(new_n593), .B(new_n592), .Y(new_n594));
  nand_5 g0319(.A(new_n594), .B(new_n591), .Y(new_n595));
  not_8  g0320(.A(new_n595), .Y(new_n596));
  xor_4  g0321(.A(new_n596), .B(new_n573), .Y(new_n597));
  not_8  g0322(.A(new_n597), .Y(new_n598));
  nand_5 g0323(.A(new_n598), .B(pi21), .Y(new_n599));
  not_8  g0324(.A(new_n599), .Y(new_n600));
  nand_5 g0325(.A(pi34), .B(pi14), .Y(new_n601));
  nand_5 g0326(.A(new_n601), .B(new_n580), .Y(new_n602));
  not_8  g0327(.A(new_n602), .Y(new_n603));
  xor_4  g0328(.A(new_n603), .B(new_n571), .Y(new_n604));
  not_8  g0329(.A(new_n604), .Y(new_n605));
  nand_5 g0330(.A(new_n605), .B(pi69), .Y(new_n606));
  nor_5  g0331(.A(new_n563), .B(new_n558), .Y(new_n607));
  nor_5  g0332(.A(new_n607), .B(new_n567), .Y(new_n608));
  xor_4  g0333(.A(new_n608), .B(new_n543), .Y(new_n609));
  nor_5  g0334(.A(pi71), .B(pi19), .Y(new_n610));
  not_8  g0335(.A(new_n610), .Y(new_n611));
  nand_5 g0336(.A(pi71), .B(pi19), .Y(new_n612));
  or_6   g0337(.A(pi56), .B(pi43), .Y(new_n613));
  nand_5 g0338(.A(pi56), .B(pi43), .Y(new_n614));
  nand_5 g0339(.A(pi63), .B(pi40), .Y(new_n615));
  nand_5 g0340(.A(new_n615), .B(new_n614), .Y(new_n616));
  nand_5 g0341(.A(new_n616), .B(new_n613), .Y(new_n617));
  nand_5 g0342(.A(new_n617), .B(new_n612), .Y(new_n618));
  nand_5 g0343(.A(new_n618), .B(new_n611), .Y(new_n619));
  nor_5  g0344(.A(pi62), .B(pi30), .Y(new_n620));
  or_6   g0345(.A(new_n620), .B(new_n619), .Y(new_n621));
  nand_5 g0346(.A(pi62), .B(pi30), .Y(new_n622));
  nand_5 g0347(.A(new_n622), .B(new_n621), .Y(new_n623));
  not_8  g0348(.A(new_n623), .Y(new_n624));
  or_6   g0349(.A(pi87), .B(pi85), .Y(new_n625));
  nand_5 g0350(.A(pi87), .B(pi85), .Y(new_n626));
  nand_5 g0351(.A(new_n626), .B(new_n625), .Y(new_n627));
  xor_4  g0352(.A(new_n627), .B(new_n624), .Y(new_n628));
  not_8  g0353(.A(new_n628), .Y(new_n629));
  nor_5  g0354(.A(new_n629), .B(new_n609), .Y(new_n630));
  xor_4  g0355(.A(new_n629), .B(new_n609), .Y(new_n631));
  xor_4  g0356(.A(pi62), .B(new_n505), .Y(new_n632));
  xor_4  g0357(.A(new_n632), .B(new_n619), .Y(new_n633));
  nand_5 g0358(.A(new_n565), .B(new_n547), .Y(new_n634));
  xor_4  g0359(.A(new_n634), .B(new_n561), .Y(new_n635));
  nor_5  g0360(.A(new_n635), .B(new_n633), .Y(new_n636));
  xnor_4 g0361(.A(new_n635), .B(new_n633), .Y(new_n637));
  nand_5 g0362(.A(new_n559), .B(new_n557), .Y(new_n638));
  xor_4  g0363(.A(new_n638), .B(new_n553), .Y(new_n639));
  nand_5 g0364(.A(new_n611), .B(new_n612), .Y(new_n640));
  xor_4  g0365(.A(new_n640), .B(new_n617), .Y(new_n641));
  nand_5 g0366(.A(new_n641), .B(new_n639), .Y(new_n642));
  nor_5  g0367(.A(new_n641), .B(new_n639), .Y(new_n643));
  not_8  g0368(.A(new_n551), .Y(new_n644));
  xor_4  g0369(.A(new_n644), .B(pi28), .Y(new_n645));
  nand_5 g0370(.A(new_n614), .B(new_n613), .Y(new_n646));
  xor_4  g0371(.A(new_n646), .B(new_n615), .Y(new_n647));
  not_8  g0372(.A(new_n647), .Y(new_n648));
  nor_5  g0373(.A(new_n648), .B(new_n645), .Y(new_n649));
  nand_5 g0374(.A(pi76), .B(pi14), .Y(new_n650));
  nand_5 g0375(.A(pi18), .B(new_n532), .Y(new_n651));
  nand_5 g0376(.A(new_n651), .B(new_n650), .Y(new_n652));
  nand_5 g0377(.A(new_n652), .B(pi48), .Y(new_n653));
  not_8  g0378(.A(new_n653), .Y(new_n654));
  nor_5  g0379(.A(new_n652), .B(pi48), .Y(new_n655));
  not_8  g0380(.A(pi63), .Y(new_n656));
  not_8  g0381(.A(new_n652), .Y(new_n657));
  nand_5 g0382(.A(new_n657), .B(new_n656), .Y(new_n658));
  nand_5 g0383(.A(new_n652), .B(pi63), .Y(new_n659));
  nand_5 g0384(.A(new_n659), .B(new_n658), .Y(po125));
  not_8  g0385(.A(po125), .Y(po058));
  xor_4  g0386(.A(pi48), .B(pi40), .Y(new_n662));
  xor_4  g0387(.A(new_n662), .B(po058), .Y(po037));
  nor_5  g0388(.A(po037), .B(new_n655), .Y(new_n664));
  nor_5  g0389(.A(new_n664), .B(new_n654), .Y(new_n665));
  not_8  g0390(.A(new_n665), .Y(new_n666));
  xor_4  g0391(.A(new_n648), .B(new_n645), .Y(new_n667));
  nand_5 g0392(.A(new_n667), .B(new_n666), .Y(new_n668));
  not_8  g0393(.A(new_n668), .Y(new_n669));
  nor_5  g0394(.A(new_n669), .B(new_n649), .Y(new_n670));
  or_6   g0395(.A(new_n670), .B(new_n643), .Y(new_n671));
  nand_5 g0396(.A(new_n671), .B(new_n642), .Y(new_n672));
  nor_5  g0397(.A(new_n672), .B(new_n637), .Y(new_n673));
  nor_5  g0398(.A(new_n673), .B(new_n636), .Y(new_n674));
  nand_5 g0399(.A(new_n674), .B(new_n631), .Y(new_n675));
  not_8  g0400(.A(new_n675), .Y(new_n676));
  nor_5  g0401(.A(new_n676), .B(new_n630), .Y(new_n677));
  not_8  g0402(.A(new_n677), .Y(new_n678));
  not_8  g0403(.A(pi69), .Y(new_n679));
  nand_5 g0404(.A(new_n604), .B(new_n679), .Y(new_n680));
  nand_5 g0405(.A(new_n680), .B(new_n606), .Y(new_n681));
  nand_5 g0406(.A(new_n626), .B(new_n624), .Y(new_n682));
  nand_5 g0407(.A(new_n682), .B(new_n625), .Y(new_n683));
  xor_4  g0408(.A(new_n683), .B(new_n681), .Y(new_n684));
  nand_5 g0409(.A(new_n684), .B(new_n678), .Y(new_n685));
  nor_5  g0410(.A(new_n685), .B(new_n606), .Y(new_n686));
  nand_5 g0411(.A(new_n686), .B(new_n600), .Y(new_n687));
  not_8  g0412(.A(new_n685), .Y(new_n688));
  not_8  g0413(.A(new_n680), .Y(new_n689));
  not_8  g0414(.A(new_n683), .Y(new_n690));
  nor_5  g0415(.A(new_n690), .B(new_n681), .Y(new_n691));
  nor_5  g0416(.A(new_n691), .B(new_n689), .Y(new_n692));
  nor_5  g0417(.A(new_n692), .B(new_n688), .Y(new_n693));
  or_6   g0418(.A(new_n693), .B(new_n686), .Y(new_n694));
  xor_4  g0419(.A(new_n597), .B(pi21), .Y(new_n695));
  not_8  g0420(.A(new_n695), .Y(new_n696));
  nor_5  g0421(.A(new_n696), .B(new_n694), .Y(new_n697));
  nor_5  g0422(.A(new_n697), .B(new_n693), .Y(new_n698));
  nor_5  g0423(.A(new_n698), .B(new_n600), .Y(new_n699));
  not_8  g0424(.A(new_n699), .Y(new_n700));
  nand_5 g0425(.A(new_n700), .B(new_n687), .Y(new_n701));
  xnor_4 g0426(.A(new_n701), .B(new_n590), .Y(po004));
  not_8  g0427(.A(new_n578), .Y(new_n703));
  xor_4  g0428(.A(new_n603), .B(new_n587), .Y(new_n704));
  nor_5  g0429(.A(new_n704), .B(new_n703), .Y(new_n705));
  not_8  g0430(.A(pi20), .Y(new_n706));
  nand_5 g0431(.A(new_n457), .B(new_n706), .Y(new_n707));
  not_8  g0432(.A(new_n707), .Y(new_n708));
  nand_5 g0433(.A(new_n581), .B(new_n708), .Y(new_n709));
  not_8  g0434(.A(new_n709), .Y(new_n710));
  nor_5  g0435(.A(new_n706), .B(pi14), .Y(new_n711));
  nand_5 g0436(.A(new_n711), .B(new_n584), .Y(new_n712));
  nand_5 g0437(.A(pi84), .B(pi14), .Y(new_n713));
  nand_5 g0438(.A(new_n713), .B(new_n712), .Y(new_n714));
  nor_5  g0439(.A(new_n714), .B(new_n710), .Y(new_n715));
  nand_5 g0440(.A(new_n715), .B(new_n705), .Y(new_n716));
  nor_5  g0441(.A(new_n716), .B(new_n602), .Y(new_n717));
  nor_5  g0442(.A(new_n603), .B(new_n587), .Y(new_n718));
  not_8  g0443(.A(new_n715), .Y(new_n719));
  nand_5 g0444(.A(new_n719), .B(new_n718), .Y(new_n720));
  nor_5  g0445(.A(new_n720), .B(new_n703), .Y(new_n721));
  nor_5  g0446(.A(new_n721), .B(new_n717), .Y(new_n722));
  nand_5 g0447(.A(new_n709), .B(new_n532), .Y(new_n723));
  not_8  g0448(.A(new_n723), .Y(new_n724));
  nand_5 g0449(.A(new_n724), .B(pi66), .Y(new_n725));
  not_8  g0450(.A(new_n725), .Y(new_n726));
  not_8  g0451(.A(pi66), .Y(new_n727));
  nand_5 g0452(.A(new_n710), .B(new_n727), .Y(new_n728));
  nand_5 g0453(.A(pi14), .B(pi09), .Y(new_n729));
  nand_5 g0454(.A(new_n729), .B(new_n728), .Y(new_n730));
  nor_5  g0455(.A(new_n730), .B(new_n726), .Y(new_n731));
  not_8  g0456(.A(new_n731), .Y(new_n732));
  xor_4  g0457(.A(new_n732), .B(new_n722), .Y(new_n733));
  nand_5 g0458(.A(new_n589), .B(pi81), .Y(new_n734));
  nor_5  g0459(.A(new_n687), .B(new_n734), .Y(new_n735));
  not_8  g0460(.A(new_n734), .Y(new_n736));
  nor_5  g0461(.A(new_n701), .B(new_n590), .Y(new_n737));
  nor_5  g0462(.A(new_n737), .B(new_n699), .Y(new_n738));
  nor_5  g0463(.A(new_n738), .B(new_n736), .Y(new_n739));
  nor_5  g0464(.A(new_n739), .B(new_n735), .Y(new_n740));
  not_8  g0465(.A(new_n740), .Y(new_n741));
  not_8  g0466(.A(pi35), .Y(new_n742));
  xor_4  g0467(.A(new_n719), .B(new_n705), .Y(new_n743));
  xor_4  g0468(.A(new_n743), .B(new_n742), .Y(new_n744));
  nor_5  g0469(.A(new_n744), .B(new_n741), .Y(new_n745));
  not_8  g0470(.A(new_n735), .Y(new_n746));
  nand_5 g0471(.A(new_n743), .B(pi35), .Y(new_n747));
  nand_5 g0472(.A(new_n747), .B(new_n746), .Y(new_n748));
  nor_5  g0473(.A(new_n748), .B(new_n745), .Y(new_n749));
  or_6   g0474(.A(new_n749), .B(new_n733), .Y(new_n750));
  not_8  g0475(.A(new_n733), .Y(new_n751));
  nor_5  g0476(.A(new_n747), .B(new_n746), .Y(new_n752));
  or_6   g0477(.A(new_n752), .B(new_n751), .Y(new_n753));
  nand_5 g0478(.A(new_n753), .B(new_n750), .Y(new_n754));
  nor_5  g0479(.A(new_n732), .B(new_n721), .Y(new_n755));
  nor_5  g0480(.A(new_n755), .B(new_n717), .Y(new_n756));
  nand_5 g0481(.A(new_n708), .B(new_n727), .Y(new_n757));
  nand_5 g0482(.A(new_n757), .B(pi74), .Y(new_n758));
  nand_5 g0483(.A(new_n758), .B(new_n532), .Y(new_n759));
  not_8  g0484(.A(pi31), .Y(new_n760));
  nand_5 g0485(.A(new_n760), .B(pi14), .Y(new_n761));
  nand_5 g0486(.A(new_n761), .B(new_n759), .Y(new_n762));
  not_8  g0487(.A(new_n762), .Y(new_n763));
  nand_5 g0488(.A(new_n727), .B(new_n706), .Y(new_n764));
  nor_5  g0489(.A(new_n764), .B(pi74), .Y(new_n765));
  nand_5 g0490(.A(new_n765), .B(new_n710), .Y(new_n766));
  nand_5 g0491(.A(new_n724), .B(pi74), .Y(new_n767));
  nand_5 g0492(.A(new_n767), .B(new_n766), .Y(new_n768));
  nor_5  g0493(.A(new_n768), .B(new_n763), .Y(new_n769));
  xor_4  g0494(.A(new_n769), .B(new_n756), .Y(new_n770));
  xor_4  g0495(.A(new_n770), .B(new_n754), .Y(po005));
  xor_4  g0496(.A(pi85), .B(pi27), .Y(new_n772));
  or_6   g0497(.A(pi54), .B(pi30), .Y(new_n773));
  not_8  g0498(.A(new_n773), .Y(new_n774));
  nand_5 g0499(.A(pi54), .B(pi30), .Y(new_n775));
  not_8  g0500(.A(new_n775), .Y(new_n776));
  nor_5  g0501(.A(pi37), .B(pi19), .Y(new_n777));
  xor_4  g0502(.A(pi37), .B(pi19), .Y(new_n778));
  nand_5 g0503(.A(pi56), .B(pi36), .Y(new_n779));
  nand_5 g0504(.A(new_n779), .B(new_n778), .Y(new_n780));
  not_8  g0505(.A(new_n780), .Y(new_n781));
  nor_5  g0506(.A(new_n781), .B(new_n777), .Y(new_n782));
  nor_5  g0507(.A(new_n782), .B(new_n776), .Y(new_n783));
  nor_5  g0508(.A(new_n783), .B(new_n774), .Y(new_n784));
  xor_4  g0509(.A(new_n784), .B(new_n772), .Y(new_n785));
  xor_4  g0510(.A(new_n785), .B(new_n366), .Y(new_n786));
  nor_5  g0511(.A(new_n776), .B(new_n774), .Y(new_n787));
  xor_4  g0512(.A(new_n787), .B(new_n782), .Y(new_n788));
  or_6   g0513(.A(new_n788), .B(new_n396), .Y(new_n789));
  xor_4  g0514(.A(new_n788), .B(new_n396), .Y(new_n790));
  or_6   g0515(.A(pi56), .B(pi36), .Y(new_n791));
  nand_5 g0516(.A(new_n791), .B(new_n779), .Y(new_n792));
  xor_4  g0517(.A(new_n372), .B(new_n312), .Y(new_n793));
  nand_5 g0518(.A(pi92), .B(pi63), .Y(new_n794));
  xor_4  g0519(.A(pi92), .B(pi63), .Y(new_n795));
  nand_5 g0520(.A(new_n795), .B(new_n381), .Y(new_n796));
  nand_5 g0521(.A(new_n796), .B(new_n794), .Y(new_n797));
  xor_4  g0522(.A(new_n797), .B(new_n793), .Y(new_n798));
  or_6   g0523(.A(new_n798), .B(new_n792), .Y(new_n799));
  nand_5 g0524(.A(new_n799), .B(new_n791), .Y(new_n800));
  xor_4  g0525(.A(new_n800), .B(new_n778), .Y(new_n801));
  not_8  g0526(.A(new_n388), .Y(new_n802));
  nand_5 g0527(.A(new_n797), .B(new_n793), .Y(new_n803));
  nand_5 g0528(.A(new_n803), .B(new_n802), .Y(new_n804));
  nor_5  g0529(.A(new_n804), .B(new_n801), .Y(new_n805));
  nor_5  g0530(.A(new_n800), .B(new_n778), .Y(new_n806));
  or_6   g0531(.A(new_n803), .B(new_n802), .Y(new_n807));
  nand_5 g0532(.A(new_n807), .B(new_n780), .Y(new_n808));
  nor_5  g0533(.A(new_n808), .B(new_n806), .Y(new_n809));
  or_6   g0534(.A(new_n809), .B(new_n805), .Y(new_n810));
  nand_5 g0535(.A(new_n810), .B(new_n790), .Y(new_n811));
  nand_5 g0536(.A(new_n811), .B(new_n789), .Y(new_n812));
  xnor_4 g0537(.A(new_n812), .B(new_n786), .Y(po006));
  not_8  g0538(.A(pi09), .Y(new_n814));
  not_8  g0539(.A(new_n452), .Y(new_n815));
  nand_5 g0540(.A(new_n815), .B(new_n814), .Y(new_n816));
  or_6   g0541(.A(new_n816), .B(pi31), .Y(new_n817));
  nor_5  g0542(.A(new_n471), .B(pi78), .Y(new_n818));
  nand_5 g0543(.A(new_n818), .B(new_n765), .Y(new_n819));
  nand_5 g0544(.A(new_n819), .B(new_n817), .Y(new_n820));
  nand_5 g0545(.A(new_n758), .B(new_n409), .Y(new_n821));
  not_8  g0546(.A(new_n821), .Y(new_n822));
  nand_5 g0547(.A(new_n407), .B(new_n760), .Y(new_n823));
  nand_5 g0548(.A(new_n823), .B(new_n816), .Y(new_n824));
  nor_5  g0549(.A(new_n824), .B(new_n822), .Y(new_n825));
  nor_5  g0550(.A(new_n825), .B(new_n820), .Y(new_n826));
  not_8  g0551(.A(new_n826), .Y(new_n827));
  or_6   g0552(.A(new_n529), .B(new_n456), .Y(new_n828));
  nand_5 g0553(.A(new_n407), .B(new_n814), .Y(new_n829));
  nand_5 g0554(.A(new_n829), .B(new_n452), .Y(new_n830));
  nand_5 g0555(.A(new_n830), .B(new_n816), .Y(new_n831));
  not_8  g0556(.A(new_n831), .Y(new_n832));
  nand_5 g0557(.A(new_n707), .B(pi66), .Y(new_n833));
  not_8  g0558(.A(new_n833), .Y(new_n834));
  nand_5 g0559(.A(new_n757), .B(new_n409), .Y(new_n835));
  nor_5  g0560(.A(new_n835), .B(new_n834), .Y(new_n836));
  nor_5  g0561(.A(new_n836), .B(new_n832), .Y(new_n837));
  not_8  g0562(.A(new_n837), .Y(new_n838));
  nor_5  g0563(.A(new_n838), .B(new_n828), .Y(new_n839));
  xor_4  g0564(.A(new_n839), .B(new_n827), .Y(po007));
  xor_4  g0565(.A(new_n527), .B(new_n475), .Y(po008));
  xor_4  g0566(.A(new_n674), .B(new_n631), .Y(po009));
  nand_5 g0567(.A(new_n542), .B(pi85), .Y(new_n843));
  not_8  g0568(.A(new_n843), .Y(new_n844));
  xor_4  g0569(.A(new_n542), .B(pi85), .Y(new_n845));
  not_8  g0570(.A(new_n845), .Y(new_n846));
  nand_5 g0571(.A(new_n546), .B(pi30), .Y(new_n847));
  not_8  g0572(.A(new_n847), .Y(new_n848));
  or_6   g0573(.A(new_n556), .B(pi19), .Y(new_n849));
  xor_4  g0574(.A(new_n556), .B(pi19), .Y(new_n850));
  not_8  g0575(.A(pi56), .Y(new_n851));
  nand_5 g0576(.A(new_n644), .B(new_n851), .Y(new_n852));
  nand_5 g0577(.A(new_n551), .B(pi56), .Y(new_n853));
  nand_5 g0578(.A(new_n853), .B(new_n659), .Y(new_n854));
  nand_5 g0579(.A(new_n854), .B(new_n852), .Y(new_n855));
  nand_5 g0580(.A(new_n855), .B(new_n850), .Y(new_n856));
  nand_5 g0581(.A(new_n856), .B(new_n849), .Y(new_n857));
  xor_4  g0582(.A(new_n546), .B(new_n505), .Y(new_n858));
  nor_5  g0583(.A(new_n858), .B(new_n857), .Y(new_n859));
  nor_5  g0584(.A(new_n859), .B(new_n848), .Y(new_n860));
  nor_5  g0585(.A(new_n860), .B(new_n846), .Y(new_n861));
  nor_5  g0586(.A(new_n861), .B(new_n844), .Y(new_n862));
  not_8  g0587(.A(new_n862), .Y(new_n863));
  nand_5 g0588(.A(new_n863), .B(new_n602), .Y(new_n864));
  xor_4  g0589(.A(new_n864), .B(new_n596), .Y(po010));
  not_8  g0590(.A(new_n475), .Y(new_n866));
  nand_5 g0591(.A(new_n512), .B(new_n866), .Y(new_n867));
  not_8  g0592(.A(new_n867), .Y(new_n868));
  nand_5 g0593(.A(new_n868), .B(new_n467), .Y(new_n869));
  or_6   g0594(.A(new_n869), .B(new_n456), .Y(new_n870));
  nor_5  g0595(.A(new_n870), .B(new_n838), .Y(new_n871));
  xor_4  g0596(.A(new_n871), .B(new_n827), .Y(po011));
  xor_4  g0597(.A(new_n380), .B(pi18), .Y(po012));
  xor_4  g0598(.A(new_n355), .B(pi82), .Y(new_n874));
  nand_5 g0599(.A(new_n364), .B(pi39), .Y(new_n875));
  nand_5 g0600(.A(new_n363), .B(new_n298), .Y(new_n876));
  nand_5 g0601(.A(new_n368), .B(pi75), .Y(new_n877));
  or_6   g0602(.A(new_n368), .B(pi75), .Y(new_n878));
  nand_5 g0603(.A(new_n370), .B(pi06), .Y(new_n879));
  not_8  g0604(.A(new_n879), .Y(new_n880));
  nand_5 g0605(.A(new_n380), .B(pi18), .Y(new_n881));
  not_8  g0606(.A(new_n881), .Y(new_n882));
  nand_5 g0607(.A(new_n882), .B(pi59), .Y(new_n883));
  xor_4  g0608(.A(new_n882), .B(pi59), .Y(new_n884));
  nand_5 g0609(.A(new_n884), .B(new_n375), .Y(new_n885));
  nand_5 g0610(.A(new_n885), .B(new_n883), .Y(new_n886));
  not_8  g0611(.A(new_n886), .Y(new_n887));
  xor_4  g0612(.A(new_n371), .B(pi06), .Y(new_n888));
  nor_5  g0613(.A(new_n888), .B(new_n887), .Y(new_n889));
  nor_5  g0614(.A(new_n889), .B(new_n880), .Y(new_n890));
  not_8  g0615(.A(new_n890), .Y(new_n891));
  nand_5 g0616(.A(new_n891), .B(new_n878), .Y(new_n892));
  nand_5 g0617(.A(new_n892), .B(new_n877), .Y(new_n893));
  nand_5 g0618(.A(new_n893), .B(new_n876), .Y(new_n894));
  nand_5 g0619(.A(new_n894), .B(new_n875), .Y(new_n895));
  xor_4  g0620(.A(new_n895), .B(new_n874), .Y(new_n896));
  xor_4  g0621(.A(new_n888), .B(new_n887), .Y(po145));
  not_8  g0622(.A(po145), .Y(po047));
  nor_5  g0623(.A(po047), .B(new_n896), .Y(new_n899));
  nor_5  g0624(.A(new_n890), .B(new_n877), .Y(new_n900));
  nor_5  g0625(.A(new_n891), .B(new_n878), .Y(new_n901));
  nor_5  g0626(.A(new_n901), .B(new_n893), .Y(new_n902));
  nor_5  g0627(.A(new_n902), .B(new_n900), .Y(po162));
  nand_5 g0628(.A(new_n875), .B(new_n876), .Y(new_n904));
  or_6   g0629(.A(new_n901), .B(new_n900), .Y(new_n905));
  xor_4  g0630(.A(new_n905), .B(new_n904), .Y(new_n906));
  not_8  g0631(.A(new_n906), .Y(po147));
  nand_5 g0632(.A(po147), .B(po162), .Y(new_n908));
  xnor_4 g0633(.A(new_n908), .B(new_n896), .Y(po099));
  nor_5  g0634(.A(po099), .B(po145), .Y(new_n910));
  nor_5  g0635(.A(new_n910), .B(new_n899), .Y(po013));
  xor_4  g0636(.A(new_n389), .B(new_n802), .Y(po014));
  and_6  g0637(.A(pi72), .B(pi30), .Y(new_n913));
  and_6  g0638(.A(pi29), .B(pi19), .Y(new_n914));
  and_6  g0639(.A(pi56), .B(pi23), .Y(new_n915));
  xor_4  g0640(.A(pi56), .B(pi23), .Y(new_n916));
  not_8  g0641(.A(new_n916), .Y(new_n917));
  nand_5 g0642(.A(pi63), .B(pi10), .Y(new_n918));
  nor_5  g0643(.A(new_n918), .B(new_n917), .Y(new_n919));
  nor_5  g0644(.A(new_n919), .B(new_n915), .Y(new_n920));
  not_8  g0645(.A(pi19), .Y(new_n921));
  xor_4  g0646(.A(pi29), .B(new_n921), .Y(new_n922));
  nor_5  g0647(.A(new_n922), .B(new_n920), .Y(new_n923));
  nor_5  g0648(.A(new_n923), .B(new_n914), .Y(new_n924));
  xor_4  g0649(.A(pi72), .B(new_n505), .Y(new_n925));
  nor_5  g0650(.A(new_n925), .B(new_n924), .Y(new_n926));
  nor_5  g0651(.A(new_n926), .B(new_n913), .Y(new_n927));
  not_8  g0652(.A(new_n546), .Y(new_n928));
  or_6   g0653(.A(new_n556), .B(pi11), .Y(new_n929));
  nand_5 g0654(.A(new_n551), .B(pi88), .Y(new_n930));
  xor_4  g0655(.A(new_n556), .B(pi11), .Y(new_n931));
  nand_5 g0656(.A(new_n931), .B(new_n930), .Y(new_n932));
  nand_5 g0657(.A(new_n932), .B(new_n929), .Y(new_n933));
  nor_5  g0658(.A(new_n933), .B(new_n928), .Y(new_n934));
  xor_4  g0659(.A(new_n934), .B(new_n542), .Y(new_n935));
  nand_5 g0660(.A(pi85), .B(pi24), .Y(new_n936));
  or_6   g0661(.A(pi85), .B(pi24), .Y(new_n937));
  nand_5 g0662(.A(new_n937), .B(new_n936), .Y(new_n938));
  xor_4  g0663(.A(new_n938), .B(new_n935), .Y(new_n939));
  nor_5  g0664(.A(new_n939), .B(new_n927), .Y(new_n940));
  xor_4  g0665(.A(new_n933), .B(new_n928), .Y(new_n941));
  xor_4  g0666(.A(new_n925), .B(new_n924), .Y(new_n942));
  or_6   g0667(.A(new_n942), .B(new_n941), .Y(new_n943));
  xor_4  g0668(.A(new_n922), .B(new_n920), .Y(new_n944));
  xnor_4 g0669(.A(new_n931), .B(new_n930), .Y(new_n945));
  nor_5  g0670(.A(new_n945), .B(new_n944), .Y(new_n946));
  xnor_4 g0671(.A(new_n945), .B(new_n944), .Y(new_n947));
  xor_4  g0672(.A(new_n551), .B(pi88), .Y(new_n948));
  nand_5 g0673(.A(pi33), .B(pi10), .Y(new_n949));
  or_6   g0674(.A(new_n949), .B(new_n659), .Y(new_n950));
  not_8  g0675(.A(new_n950), .Y(new_n951));
  xor_4  g0676(.A(pi33), .B(pi10), .Y(new_n952));
  nand_5 g0677(.A(new_n952), .B(po058), .Y(new_n953));
  not_8  g0678(.A(new_n953), .Y(new_n954));
  nand_5 g0679(.A(new_n949), .B(new_n659), .Y(new_n955));
  nor_5  g0680(.A(new_n955), .B(new_n954), .Y(new_n956));
  nor_5  g0681(.A(new_n956), .B(new_n951), .Y(new_n957));
  xor_4  g0682(.A(new_n957), .B(new_n916), .Y(new_n958));
  nand_5 g0683(.A(new_n958), .B(new_n948), .Y(new_n959));
  nand_5 g0684(.A(new_n957), .B(new_n917), .Y(new_n960));
  nor_5  g0685(.A(new_n956), .B(new_n919), .Y(new_n961));
  nand_5 g0686(.A(new_n961), .B(new_n960), .Y(new_n962));
  nand_5 g0687(.A(new_n962), .B(new_n959), .Y(new_n963));
  nor_5  g0688(.A(new_n963), .B(new_n947), .Y(new_n964));
  or_6   g0689(.A(new_n964), .B(new_n946), .Y(new_n965));
  xor_4  g0690(.A(new_n942), .B(new_n941), .Y(new_n966));
  nand_5 g0691(.A(new_n966), .B(new_n965), .Y(new_n967));
  nand_5 g0692(.A(new_n967), .B(new_n943), .Y(new_n968));
  xor_4  g0693(.A(new_n939), .B(new_n927), .Y(new_n969));
  not_8  g0694(.A(new_n969), .Y(new_n970));
  nor_5  g0695(.A(new_n970), .B(new_n968), .Y(new_n971));
  or_6   g0696(.A(new_n971), .B(new_n940), .Y(new_n972));
  nand_5 g0697(.A(new_n934), .B(new_n542), .Y(new_n973));
  not_8  g0698(.A(new_n973), .Y(new_n974));
  nand_5 g0699(.A(new_n974), .B(new_n602), .Y(new_n975));
  nand_5 g0700(.A(new_n973), .B(new_n603), .Y(new_n976));
  nand_5 g0701(.A(new_n976), .B(new_n975), .Y(new_n977));
  xnor_4 g0702(.A(new_n977), .B(pi01), .Y(new_n978));
  nand_5 g0703(.A(new_n937), .B(new_n935), .Y(new_n979));
  nand_5 g0704(.A(new_n979), .B(new_n936), .Y(new_n980));
  xnor_4 g0705(.A(new_n980), .B(new_n978), .Y(new_n981));
  xnor_4 g0706(.A(new_n981), .B(new_n972), .Y(po015));
  xnor_4 g0707(.A(new_n963), .B(new_n947), .Y(po016));
  nor_5  g0708(.A(new_n752), .B(new_n749), .Y(new_n984));
  xor_4  g0709(.A(new_n984), .B(new_n751), .Y(po017));
  xor_4  g0710(.A(new_n719), .B(pi89), .Y(new_n986));
  xor_4  g0711(.A(new_n588), .B(pi44), .Y(new_n987));
  nand_5 g0712(.A(new_n595), .B(pi58), .Y(new_n988));
  nor_5  g0713(.A(new_n980), .B(new_n978), .Y(new_n989));
  nor_5  g0714(.A(new_n981), .B(new_n972), .Y(new_n990));
  nor_5  g0715(.A(new_n990), .B(new_n989), .Y(new_n991));
  nand_5 g0716(.A(new_n976), .B(pi01), .Y(new_n992));
  nand_5 g0717(.A(new_n992), .B(new_n975), .Y(new_n993));
  nand_5 g0718(.A(new_n993), .B(new_n991), .Y(new_n994));
  xor_4  g0719(.A(new_n994), .B(new_n988), .Y(new_n995));
  xor_4  g0720(.A(new_n596), .B(pi58), .Y(new_n996));
  xor_4  g0721(.A(new_n993), .B(new_n991), .Y(new_n997));
  not_8  g0722(.A(new_n997), .Y(new_n998));
  nor_5  g0723(.A(new_n998), .B(new_n996), .Y(new_n999));
  or_6   g0724(.A(new_n999), .B(new_n995), .Y(new_n1000));
  nand_5 g0725(.A(new_n1000), .B(new_n987), .Y(new_n1001));
  nand_5 g0726(.A(new_n588), .B(pi44), .Y(new_n1002));
  nor_5  g0727(.A(new_n994), .B(new_n988), .Y(new_n1003));
  xor_4  g0728(.A(new_n1003), .B(new_n1002), .Y(new_n1004));
  nand_5 g0729(.A(new_n1004), .B(new_n1001), .Y(new_n1005));
  xor_4  g0730(.A(new_n1005), .B(new_n986), .Y(po018));
  nor_5  g0731(.A(new_n295), .B(new_n276), .Y(new_n1007));
  xor_4  g0732(.A(new_n1007), .B(pi80), .Y(new_n1008));
  not_8  g0733(.A(new_n1008), .Y(new_n1009));
  nand_5 g0734(.A(new_n1009), .B(new_n441), .Y(new_n1010));
  xor_4  g0735(.A(new_n1008), .B(pi78), .Y(new_n1011));
  not_8  g0736(.A(new_n1011), .Y(new_n1012));
  nand_5 g0737(.A(new_n296), .B(pi04), .Y(new_n1013));
  nand_5 g0738(.A(new_n356), .B(new_n336), .Y(new_n1014));
  not_8  g0739(.A(new_n874), .Y(new_n1015));
  or_6   g0740(.A(new_n895), .B(new_n1015), .Y(new_n1016));
  nand_5 g0741(.A(new_n1016), .B(new_n1014), .Y(new_n1017));
  xor_4  g0742(.A(new_n296), .B(new_n440), .Y(new_n1018));
  or_6   g0743(.A(new_n1018), .B(new_n1017), .Y(new_n1019));
  nand_5 g0744(.A(new_n1019), .B(new_n1013), .Y(new_n1020));
  or_6   g0745(.A(new_n1020), .B(new_n1012), .Y(new_n1021));
  nand_5 g0746(.A(new_n1021), .B(new_n1010), .Y(new_n1022));
  nand_5 g0747(.A(new_n1007), .B(pi80), .Y(new_n1023));
  not_8  g0748(.A(new_n1023), .Y(new_n1024));
  nand_5 g0749(.A(new_n1024), .B(pi38), .Y(new_n1025));
  or_6   g0750(.A(new_n1024), .B(pi38), .Y(new_n1026));
  nand_5 g0751(.A(new_n1026), .B(new_n1025), .Y(new_n1027));
  xor_4  g0752(.A(new_n1027), .B(pi20), .Y(new_n1028));
  or_6   g0753(.A(new_n1028), .B(new_n1022), .Y(new_n1029));
  nand_5 g0754(.A(new_n1029), .B(new_n727), .Y(new_n1030));
  or_6   g0755(.A(new_n1029), .B(new_n727), .Y(new_n1031));
  nand_5 g0756(.A(new_n1031), .B(new_n1030), .Y(new_n1032));
  nand_5 g0757(.A(new_n1025), .B(new_n706), .Y(new_n1033));
  nand_5 g0758(.A(new_n1033), .B(new_n1026), .Y(new_n1034));
  xor_4  g0759(.A(new_n1034), .B(new_n1032), .Y(new_n1035));
  nor_5  g0760(.A(new_n908), .B(new_n896), .Y(new_n1036));
  not_8  g0761(.A(new_n1036), .Y(new_n1037));
  xor_4  g0762(.A(new_n1018), .B(new_n1017), .Y(new_n1038));
  nor_5  g0763(.A(new_n1038), .B(new_n1037), .Y(new_n1039));
  not_8  g0764(.A(new_n1039), .Y(new_n1040));
  xor_4  g0765(.A(new_n1020), .B(new_n1011), .Y(new_n1041));
  nor_5  g0766(.A(new_n1041), .B(new_n1040), .Y(new_n1042));
  not_8  g0767(.A(new_n1042), .Y(new_n1043));
  xor_4  g0768(.A(new_n1028), .B(new_n1022), .Y(new_n1044));
  nor_5  g0769(.A(new_n1044), .B(new_n1043), .Y(new_n1045));
  not_8  g0770(.A(new_n1045), .Y(new_n1046));
  nor_5  g0771(.A(new_n1046), .B(new_n1035), .Y(new_n1047));
  nand_5 g0772(.A(new_n1047), .B(po047), .Y(new_n1048));
  nand_5 g0773(.A(new_n1045), .B(po047), .Y(new_n1049));
  nand_5 g0774(.A(new_n1049), .B(new_n1035), .Y(new_n1050));
  nand_5 g0775(.A(new_n1050), .B(new_n1048), .Y(po019));
  xor_4  g0776(.A(new_n609), .B(new_n363), .Y(new_n1052));
  or_6   g0777(.A(new_n639), .B(new_n370), .Y(new_n1053));
  xor_4  g0778(.A(new_n639), .B(new_n370), .Y(new_n1054));
  nand_5 g0779(.A(new_n645), .B(new_n374), .Y(new_n1055));
  xor_4  g0780(.A(new_n645), .B(new_n374), .Y(new_n1056));
  nand_5 g0781(.A(new_n657), .B(new_n379), .Y(new_n1057));
  not_8  g0782(.A(pi48), .Y(new_n1058));
  nand_5 g0783(.A(new_n652), .B(new_n380), .Y(new_n1059));
  nand_5 g0784(.A(new_n1059), .B(new_n1057), .Y(new_n1060));
  not_8  g0785(.A(new_n1060), .Y(new_n1061));
  nand_5 g0786(.A(new_n1061), .B(new_n1058), .Y(new_n1062));
  nand_5 g0787(.A(new_n1062), .B(new_n1057), .Y(new_n1063));
  nand_5 g0788(.A(new_n1063), .B(new_n1056), .Y(new_n1064));
  nand_5 g0789(.A(new_n1064), .B(new_n1055), .Y(new_n1065));
  nand_5 g0790(.A(new_n1065), .B(new_n1054), .Y(new_n1066));
  nand_5 g0791(.A(new_n1066), .B(new_n1053), .Y(new_n1067));
  and_6  g0792(.A(new_n1067), .B(new_n369), .Y(new_n1068));
  nor_5  g0793(.A(new_n1067), .B(new_n369), .Y(new_n1069));
  nor_5  g0794(.A(new_n1069), .B(new_n635), .Y(new_n1070));
  or_6   g0795(.A(new_n1070), .B(new_n1068), .Y(new_n1071));
  xnor_4 g0796(.A(new_n1071), .B(new_n1052), .Y(po020));
  xor_4  g0797(.A(new_n795), .B(new_n381), .Y(po021));
  xor_4  g0798(.A(new_n884), .B(new_n375), .Y(po022));
  not_8  g0799(.A(new_n1002), .Y(new_n1075));
  nand_5 g0800(.A(new_n1003), .B(new_n1075), .Y(new_n1076));
  nand_5 g0801(.A(new_n1076), .B(new_n731), .Y(new_n1077));
  not_8  g0802(.A(new_n1077), .Y(new_n1078));
  xor_4  g0803(.A(new_n1076), .B(new_n731), .Y(new_n1079));
  not_8  g0804(.A(new_n1079), .Y(new_n1080));
  nor_5  g0805(.A(new_n719), .B(pi89), .Y(new_n1081));
  not_8  g0806(.A(new_n986), .Y(new_n1082));
  nor_5  g0807(.A(new_n1005), .B(new_n1082), .Y(new_n1083));
  nor_5  g0808(.A(new_n1083), .B(new_n1081), .Y(new_n1084));
  nor_5  g0809(.A(new_n1084), .B(new_n1080), .Y(new_n1085));
  nor_5  g0810(.A(new_n1085), .B(new_n1078), .Y(new_n1086));
  nor_5  g0811(.A(new_n1086), .B(new_n766), .Y(po023));
  not_8  g0812(.A(pi46), .Y(new_n1088));
  nand_5 g0813(.A(new_n483), .B(new_n1088), .Y(new_n1089));
  not_8  g0814(.A(new_n1089), .Y(new_n1090));
  nor_5  g0815(.A(pi64), .B(pi30), .Y(new_n1091));
  xor_4  g0816(.A(pi64), .B(pi30), .Y(new_n1092));
  not_8  g0817(.A(new_n1092), .Y(new_n1093));
  nor_5  g0818(.A(pi42), .B(pi19), .Y(new_n1094));
  nand_5 g0819(.A(pi67), .B(pi56), .Y(new_n1095));
  not_8  g0820(.A(new_n1095), .Y(new_n1096));
  xor_4  g0821(.A(pi42), .B(new_n921), .Y(new_n1097));
  nor_5  g0822(.A(new_n1097), .B(new_n1096), .Y(new_n1098));
  nor_5  g0823(.A(new_n1098), .B(new_n1094), .Y(new_n1099));
  nor_5  g0824(.A(new_n1099), .B(new_n1093), .Y(new_n1100));
  nor_5  g0825(.A(new_n1100), .B(new_n1091), .Y(new_n1101));
  xor_4  g0826(.A(pi85), .B(new_n1088), .Y(new_n1102));
  nor_5  g0827(.A(new_n1102), .B(new_n1101), .Y(new_n1103));
  nor_5  g0828(.A(new_n1103), .B(new_n1090), .Y(new_n1104));
  nand_5 g0829(.A(new_n1104), .B(pi50), .Y(new_n1105));
  nor_5  g0830(.A(new_n492), .B(pi70), .Y(new_n1106));
  xor_4  g0831(.A(new_n492), .B(pi70), .Y(new_n1107));
  not_8  g0832(.A(new_n1107), .Y(new_n1108));
  nor_5  g0833(.A(new_n430), .B(pi07), .Y(new_n1109));
  nor_5  g0834(.A(new_n436), .B(new_n432), .Y(new_n1110));
  nor_5  g0835(.A(new_n1110), .B(new_n1109), .Y(new_n1111));
  nor_5  g0836(.A(new_n1111), .B(new_n1108), .Y(new_n1112));
  or_6   g0837(.A(new_n1112), .B(new_n1106), .Y(new_n1113));
  nor_5  g0838(.A(new_n1113), .B(new_n487), .Y(new_n1114));
  xor_4  g0839(.A(new_n1114), .B(new_n481), .Y(new_n1115));
  xor_4  g0840(.A(new_n1113), .B(new_n487), .Y(new_n1116));
  xor_4  g0841(.A(new_n1102), .B(new_n1101), .Y(new_n1117));
  not_8  g0842(.A(new_n1117), .Y(new_n1118));
  nand_5 g0843(.A(new_n1118), .B(new_n1116), .Y(new_n1119));
  xor_4  g0844(.A(new_n1118), .B(new_n1116), .Y(new_n1120));
  xor_4  g0845(.A(new_n1111), .B(new_n1107), .Y(new_n1121));
  xor_4  g0846(.A(new_n1099), .B(new_n1092), .Y(new_n1122));
  nor_5  g0847(.A(new_n1122), .B(new_n1121), .Y(new_n1123));
  xnor_4 g0848(.A(new_n1122), .B(new_n1121), .Y(new_n1124));
  xor_4  g0849(.A(new_n1097), .B(new_n1096), .Y(new_n1125));
  xor_4  g0850(.A(pi67), .B(pi56), .Y(new_n1126));
  or_6   g0851(.A(new_n1126), .B(new_n421), .Y(new_n1127));
  xor_4  g0852(.A(new_n1126), .B(new_n421), .Y(new_n1128));
  nor_5  g0853(.A(pi63), .B(pi61), .Y(new_n1129));
  xor_4  g0854(.A(new_n656), .B(pi61), .Y(new_n1130));
  nor_5  g0855(.A(new_n1130), .B(new_n412), .Y(new_n1131));
  or_6   g0856(.A(new_n1131), .B(new_n1129), .Y(new_n1132));
  nand_5 g0857(.A(new_n1132), .B(new_n1128), .Y(new_n1133));
  nand_5 g0858(.A(new_n1133), .B(new_n1127), .Y(new_n1134));
  nor_5  g0859(.A(new_n1134), .B(new_n1125), .Y(new_n1135));
  xor_4  g0860(.A(new_n1134), .B(new_n1125), .Y(new_n1136));
  nand_5 g0861(.A(new_n1136), .B(new_n438), .Y(new_n1137));
  not_8  g0862(.A(new_n1137), .Y(new_n1138));
  nor_5  g0863(.A(new_n1138), .B(new_n1135), .Y(new_n1139));
  not_8  g0864(.A(new_n1139), .Y(new_n1140));
  nor_5  g0865(.A(new_n1140), .B(new_n1124), .Y(new_n1141));
  nor_5  g0866(.A(new_n1141), .B(new_n1123), .Y(new_n1142));
  nand_5 g0867(.A(new_n1142), .B(new_n1120), .Y(new_n1143));
  nand_5 g0868(.A(new_n1143), .B(new_n1119), .Y(new_n1144));
  nand_5 g0869(.A(new_n1144), .B(new_n1115), .Y(new_n1145));
  nor_5  g0870(.A(new_n1145), .B(new_n1105), .Y(new_n1146));
  or_6   g0871(.A(new_n1144), .B(new_n1115), .Y(new_n1147));
  nand_5 g0872(.A(new_n1147), .B(new_n1145), .Y(new_n1148));
  xor_4  g0873(.A(new_n1104), .B(pi50), .Y(new_n1149));
  or_6   g0874(.A(new_n1149), .B(new_n1148), .Y(new_n1150));
  nand_5 g0875(.A(new_n1150), .B(new_n1147), .Y(new_n1151));
  and_6  g0876(.A(new_n1151), .B(new_n1105), .Y(new_n1152));
  or_6   g0877(.A(new_n1152), .B(new_n1146), .Y(new_n1153));
  nand_5 g0878(.A(new_n1114), .B(new_n481), .Y(new_n1154));
  xor_4  g0879(.A(new_n1154), .B(new_n475), .Y(new_n1155));
  not_8  g0880(.A(new_n1155), .Y(new_n1156));
  xor_4  g0881(.A(new_n1156), .B(pi65), .Y(new_n1157));
  xor_4  g0882(.A(new_n1157), .B(new_n1153), .Y(po024));
  xor_4  g0883(.A(new_n1130), .B(new_n422), .Y(po025));
  xnor_4 g0884(.A(new_n810), .B(new_n790), .Y(po026));
  not_8  g0885(.A(new_n766), .Y(new_n1161));
  nand_5 g0886(.A(new_n862), .B(new_n1161), .Y(new_n1162));
  not_8  g0887(.A(new_n1162), .Y(po076));
  xor_4  g0888(.A(new_n858), .B(new_n857), .Y(po172));
  xor_4  g0889(.A(new_n855), .B(new_n850), .Y(new_n1165));
  not_8  g0890(.A(new_n658), .Y(new_n1166));
  nor_5  g0891(.A(new_n853), .B(new_n1166), .Y(new_n1167));
  nor_5  g0892(.A(new_n852), .B(new_n658), .Y(new_n1168));
  or_6   g0893(.A(new_n1168), .B(new_n1167), .Y(new_n1169));
  xor_4  g0894(.A(new_n1169), .B(new_n850), .Y(po066));
  nand_5 g0895(.A(po066), .B(new_n1165), .Y(new_n1171));
  nand_5 g0896(.A(new_n1171), .B(po172), .Y(new_n1172));
  xor_4  g0897(.A(new_n860), .B(new_n845), .Y(new_n1173));
  or_6   g0898(.A(new_n1173), .B(new_n1172), .Y(new_n1174));
  nand_5 g0899(.A(new_n1174), .B(po076), .Y(new_n1175));
  nand_5 g0900(.A(new_n862), .B(new_n603), .Y(new_n1176));
  nand_5 g0901(.A(new_n1174), .B(new_n864), .Y(new_n1177));
  nand_5 g0902(.A(new_n1177), .B(new_n1176), .Y(new_n1178));
  nor_5  g0903(.A(new_n1178), .B(new_n596), .Y(new_n1179));
  nand_5 g0904(.A(new_n1179), .B(new_n588), .Y(new_n1180));
  nor_5  g0905(.A(new_n1180), .B(new_n715), .Y(new_n1181));
  and_6  g0906(.A(new_n1181), .B(new_n732), .Y(new_n1182));
  nand_5 g0907(.A(new_n1182), .B(new_n763), .Y(new_n1183));
  nand_5 g0908(.A(new_n1183), .B(new_n1175), .Y(po027));
  nor_5  g0909(.A(new_n1154), .B(new_n475), .Y(new_n1185));
  xor_4  g0910(.A(new_n1185), .B(new_n467), .Y(new_n1186));
  xor_4  g0911(.A(new_n1186), .B(pi90), .Y(new_n1187));
  nor_5  g0912(.A(new_n1157), .B(new_n1153), .Y(new_n1188));
  nand_5 g0913(.A(new_n1155), .B(pi65), .Y(new_n1189));
  not_8  g0914(.A(new_n1189), .Y(new_n1190));
  xor_4  g0915(.A(new_n1190), .B(new_n1146), .Y(new_n1191));
  nor_5  g0916(.A(new_n1191), .B(new_n1188), .Y(new_n1192));
  xnor_4 g0917(.A(new_n1192), .B(new_n1187), .Y(po028));
  not_8  g0918(.A(new_n515), .Y(po029));
  nand_5 g0919(.A(new_n807), .B(new_n804), .Y(new_n1195));
  xor_4  g0920(.A(new_n1195), .B(new_n801), .Y(po030));
  or_6   g0921(.A(new_n426), .B(new_n371), .Y(new_n1197));
  nand_5 g0922(.A(new_n438), .B(new_n427), .Y(new_n1198));
  nand_5 g0923(.A(new_n1198), .B(new_n1197), .Y(new_n1199));
  xor_4  g0924(.A(new_n1199), .B(new_n368), .Y(new_n1200));
  xor_4  g0925(.A(new_n1200), .B(new_n1121), .Y(po031));
  not_8  g0926(.A(new_n769), .Y(new_n1202));
  xor_4  g0927(.A(new_n1182), .B(new_n1202), .Y(po032));
  and_6  g0928(.A(new_n1176), .B(new_n864), .Y(po071));
  xnor_4 g0929(.A(po071), .B(new_n1174), .Y(po033));
  xor_4  g0930(.A(new_n1116), .B(new_n364), .Y(new_n1206));
  nand_5 g0931(.A(new_n1199), .B(new_n368), .Y(new_n1207));
  nand_5 g0932(.A(new_n1200), .B(new_n1121), .Y(new_n1208));
  nand_5 g0933(.A(new_n1208), .B(new_n1207), .Y(new_n1209));
  xor_4  g0934(.A(new_n1209), .B(new_n1206), .Y(po034));
  nor_5  g0935(.A(new_n1038), .B(po047), .Y(new_n1211));
  xor_4  g0936(.A(new_n1038), .B(new_n1036), .Y(po113));
  nor_5  g0937(.A(po113), .B(po145), .Y(new_n1213));
  nor_5  g0938(.A(new_n1213), .B(new_n1211), .Y(po035));
  xor_4  g0939(.A(new_n1084), .B(new_n1079), .Y(po036));
  xor_4  g0940(.A(new_n395), .B(new_n393), .Y(po038));
  or_6   g0941(.A(new_n864), .B(new_n596), .Y(new_n1217));
  nor_5  g0942(.A(new_n1217), .B(new_n587), .Y(new_n1218));
  nand_5 g0943(.A(new_n1218), .B(new_n719), .Y(new_n1219));
  nor_5  g0944(.A(new_n1219), .B(new_n731), .Y(new_n1220));
  xor_4  g0945(.A(new_n1220), .B(new_n1202), .Y(po040));
  nand_5 g0946(.A(new_n1185), .B(new_n467), .Y(new_n1222));
  not_8  g0947(.A(new_n1222), .Y(new_n1223));
  nand_5 g0948(.A(new_n1156), .B(new_n297), .Y(new_n1224));
  xor_4  g0949(.A(new_n1155), .B(new_n296), .Y(new_n1225));
  nor_5  g0950(.A(new_n1115), .B(new_n355), .Y(new_n1226));
  nor_5  g0951(.A(new_n1116), .B(new_n364), .Y(new_n1227));
  not_8  g0952(.A(new_n1206), .Y(new_n1228));
  nor_5  g0953(.A(new_n1209), .B(new_n1228), .Y(new_n1229));
  nor_5  g0954(.A(new_n1229), .B(new_n1227), .Y(new_n1230));
  xor_4  g0955(.A(new_n1115), .B(new_n356), .Y(new_n1231));
  nor_5  g0956(.A(new_n1231), .B(new_n1230), .Y(new_n1232));
  or_6   g0957(.A(new_n1232), .B(new_n1226), .Y(new_n1233));
  nand_5 g0958(.A(new_n1233), .B(new_n1225), .Y(new_n1234));
  nand_5 g0959(.A(new_n1234), .B(new_n1224), .Y(new_n1235));
  xor_4  g0960(.A(new_n1186), .B(new_n1009), .Y(new_n1236));
  nor_5  g0961(.A(new_n1236), .B(new_n1235), .Y(new_n1237));
  nand_5 g0962(.A(new_n1237), .B(new_n1223), .Y(new_n1238));
  nand_5 g0963(.A(new_n1238), .B(new_n1025), .Y(new_n1239));
  xor_4  g0964(.A(new_n1239), .B(new_n837), .Y(new_n1240));
  nand_5 g0965(.A(new_n1027), .B(new_n456), .Y(new_n1241));
  not_8  g0966(.A(new_n1241), .Y(new_n1242));
  xor_4  g0967(.A(new_n1027), .B(new_n456), .Y(new_n1243));
  not_8  g0968(.A(new_n1243), .Y(new_n1244));
  nand_5 g0969(.A(new_n1186), .B(new_n1008), .Y(new_n1245));
  xor_4  g0970(.A(new_n1237), .B(new_n1222), .Y(new_n1246));
  nand_5 g0971(.A(new_n1246), .B(new_n1245), .Y(new_n1247));
  nor_5  g0972(.A(new_n1247), .B(new_n1244), .Y(new_n1248));
  nor_5  g0973(.A(new_n1248), .B(new_n1242), .Y(new_n1249));
  xor_4  g0974(.A(new_n1249), .B(new_n1240), .Y(po041));
  xor_4  g0975(.A(new_n1027), .B(new_n715), .Y(new_n1251));
  xor_4  g0976(.A(new_n1008), .B(new_n588), .Y(new_n1252));
  xor_4  g0977(.A(new_n595), .B(new_n296), .Y(new_n1253));
  or_6   g0978(.A(new_n941), .B(new_n368), .Y(new_n1254));
  xor_4  g0979(.A(new_n941), .B(new_n368), .Y(new_n1255));
  or_6   g0980(.A(new_n945), .B(new_n370), .Y(new_n1256));
  xor_4  g0981(.A(new_n945), .B(new_n370), .Y(new_n1257));
  not_8  g0982(.A(new_n948), .Y(new_n1258));
  nand_5 g0983(.A(new_n1258), .B(new_n374), .Y(new_n1259));
  xor_4  g0984(.A(new_n1258), .B(new_n374), .Y(new_n1260));
  not_8  g0985(.A(new_n1260), .Y(new_n1261));
  nand_5 g0986(.A(new_n1061), .B(pi33), .Y(new_n1262));
  nand_5 g0987(.A(new_n1262), .B(new_n1059), .Y(new_n1263));
  or_6   g0988(.A(new_n1263), .B(new_n1261), .Y(new_n1264));
  nand_5 g0989(.A(new_n1264), .B(new_n1259), .Y(new_n1265));
  nand_5 g0990(.A(new_n1265), .B(new_n1257), .Y(new_n1266));
  nand_5 g0991(.A(new_n1266), .B(new_n1256), .Y(new_n1267));
  nand_5 g0992(.A(new_n1267), .B(new_n1255), .Y(new_n1268));
  nand_5 g0993(.A(new_n1268), .B(new_n1254), .Y(new_n1269));
  xor_4  g0994(.A(new_n935), .B(new_n363), .Y(new_n1270));
  nor_5  g0995(.A(new_n1270), .B(new_n1269), .Y(new_n1271));
  or_6   g0996(.A(new_n1271), .B(new_n974), .Y(new_n1272));
  nand_5 g0997(.A(new_n935), .B(new_n364), .Y(new_n1273));
  nand_5 g0998(.A(new_n602), .B(new_n355), .Y(new_n1274));
  nand_5 g0999(.A(new_n1274), .B(new_n1273), .Y(new_n1275));
  nor_5  g1000(.A(new_n1275), .B(new_n1272), .Y(new_n1276));
  nand_5 g1001(.A(new_n1271), .B(new_n974), .Y(new_n1277));
  nor_5  g1002(.A(new_n1277), .B(new_n1274), .Y(new_n1278));
  not_8  g1003(.A(new_n1278), .Y(new_n1279));
  nor_5  g1004(.A(new_n602), .B(new_n355), .Y(new_n1280));
  nand_5 g1005(.A(new_n1280), .B(new_n1277), .Y(new_n1281));
  nand_5 g1006(.A(new_n1281), .B(new_n1279), .Y(new_n1282));
  nor_5  g1007(.A(new_n1282), .B(new_n1276), .Y(new_n1283));
  nand_5 g1008(.A(new_n1283), .B(new_n1253), .Y(new_n1284));
  nand_5 g1009(.A(new_n595), .B(new_n296), .Y(new_n1285));
  xor_4  g1010(.A(new_n1278), .B(new_n1285), .Y(new_n1286));
  nand_5 g1011(.A(new_n1286), .B(new_n1284), .Y(new_n1287));
  nand_5 g1012(.A(new_n1287), .B(new_n1252), .Y(new_n1288));
  nand_5 g1013(.A(new_n1008), .B(new_n588), .Y(new_n1289));
  nor_5  g1014(.A(new_n1279), .B(new_n1285), .Y(new_n1290));
  xor_4  g1015(.A(new_n1290), .B(new_n1289), .Y(new_n1291));
  nand_5 g1016(.A(new_n1291), .B(new_n1288), .Y(new_n1292));
  xor_4  g1017(.A(new_n1292), .B(new_n1251), .Y(po042));
  nand_5 g1018(.A(new_n597), .B(new_n297), .Y(new_n1294));
  not_8  g1019(.A(new_n1294), .Y(new_n1295));
  xor_4  g1020(.A(new_n597), .B(new_n296), .Y(new_n1296));
  nand_5 g1021(.A(new_n605), .B(new_n355), .Y(new_n1297));
  not_8  g1022(.A(new_n1297), .Y(new_n1298));
  nand_5 g1023(.A(new_n609), .B(new_n363), .Y(new_n1299));
  nand_5 g1024(.A(new_n1071), .B(new_n1052), .Y(new_n1300));
  nand_5 g1025(.A(new_n1300), .B(new_n1299), .Y(new_n1301));
  xor_4  g1026(.A(new_n604), .B(new_n355), .Y(new_n1302));
  nor_5  g1027(.A(new_n1302), .B(new_n1301), .Y(new_n1303));
  nor_5  g1028(.A(new_n1303), .B(new_n1298), .Y(new_n1304));
  not_8  g1029(.A(new_n1304), .Y(new_n1305));
  nor_5  g1030(.A(new_n1305), .B(new_n1296), .Y(new_n1306));
  nor_5  g1031(.A(new_n1306), .B(new_n1295), .Y(new_n1307));
  xor_4  g1032(.A(new_n1252), .B(new_n703), .Y(new_n1308));
  nor_5  g1033(.A(new_n1308), .B(new_n1307), .Y(new_n1309));
  nor_5  g1034(.A(new_n1008), .B(new_n589), .Y(new_n1310));
  or_6   g1035(.A(new_n1310), .B(new_n1309), .Y(new_n1311));
  xor_4  g1036(.A(new_n1027), .B(new_n743), .Y(new_n1312));
  xor_4  g1037(.A(new_n1312), .B(new_n1311), .Y(po043));
  xor_4  g1038(.A(new_n1044), .B(new_n1042), .Y(po044));
  nor_5  g1039(.A(new_n299), .B(pi02), .Y(new_n1315));
  nor_5  g1040(.A(pi60), .B(new_n440), .Y(new_n1316));
  nor_5  g1041(.A(new_n1316), .B(new_n1315), .Y(new_n1317));
  nand_5 g1042(.A(new_n1317), .B(new_n340), .Y(new_n1318));
  or_6   g1043(.A(new_n341), .B(pi04), .Y(new_n1319));
  nand_5 g1044(.A(new_n1319), .B(pi78), .Y(new_n1320));
  not_8  g1045(.A(new_n1320), .Y(new_n1321));
  nor_5  g1046(.A(new_n584), .B(pi39), .Y(new_n1322));
  nor_5  g1047(.A(new_n1322), .B(new_n1321), .Y(new_n1323));
  nor_5  g1048(.A(new_n1323), .B(pi60), .Y(new_n1324));
  nand_5 g1049(.A(new_n349), .B(new_n446), .Y(new_n1325));
  not_8  g1050(.A(new_n1325), .Y(new_n1326));
  nand_5 g1051(.A(new_n348), .B(pi13), .Y(new_n1327));
  nand_5 g1052(.A(new_n1327), .B(pi60), .Y(new_n1328));
  nor_5  g1053(.A(new_n1328), .B(new_n1326), .Y(new_n1329));
  nor_5  g1054(.A(new_n1329), .B(new_n1324), .Y(new_n1330));
  not_8  g1055(.A(new_n1330), .Y(new_n1331));
  xor_4  g1056(.A(new_n1331), .B(new_n324), .Y(new_n1332));
  nor_5  g1057(.A(new_n1332), .B(new_n1318), .Y(new_n1333));
  xor_4  g1058(.A(new_n1327), .B(new_n445), .Y(new_n1334));
  nand_5 g1059(.A(new_n1334), .B(pi60), .Y(new_n1335));
  xor_4  g1060(.A(new_n1322), .B(pi20), .Y(new_n1336));
  nand_5 g1061(.A(new_n1336), .B(new_n299), .Y(new_n1337));
  nand_5 g1062(.A(new_n1337), .B(new_n1335), .Y(new_n1338));
  xor_4  g1063(.A(new_n1338), .B(new_n1333), .Y(new_n1339));
  not_8  g1064(.A(new_n1339), .Y(new_n1340));
  nand_5 g1065(.A(new_n1340), .B(pi84), .Y(new_n1341));
  or_6   g1066(.A(new_n1341), .B(pi09), .Y(new_n1342));
  nand_5 g1067(.A(new_n1342), .B(pi60), .Y(new_n1343));
  not_8  g1068(.A(new_n1343), .Y(new_n1344));
  nand_5 g1069(.A(new_n1341), .B(pi09), .Y(new_n1345));
  nand_5 g1070(.A(new_n1345), .B(new_n1344), .Y(new_n1346));
  not_8  g1071(.A(new_n1346), .Y(new_n1347));
  nand_5 g1072(.A(new_n1339), .B(new_n706), .Y(new_n1348));
  nand_5 g1073(.A(new_n1348), .B(pi66), .Y(new_n1349));
  nand_5 g1074(.A(new_n1349), .B(new_n299), .Y(new_n1350));
  nor_5  g1075(.A(new_n1348), .B(pi66), .Y(new_n1351));
  nor_5  g1076(.A(new_n1351), .B(new_n1350), .Y(new_n1352));
  nor_5  g1077(.A(new_n1352), .B(new_n1347), .Y(new_n1353));
  not_8  g1078(.A(new_n1353), .Y(new_n1354));
  xor_4  g1079(.A(new_n1339), .B(pi15), .Y(new_n1355));
  xor_4  g1080(.A(new_n1331), .B(new_n1318), .Y(new_n1356));
  not_8  g1081(.A(new_n1356), .Y(new_n1357));
  nand_5 g1082(.A(new_n1357), .B(pi53), .Y(new_n1358));
  xor_4  g1083(.A(new_n353), .B(pi83), .Y(new_n1359));
  not_8  g1084(.A(new_n1359), .Y(new_n1360));
  nand_5 g1085(.A(pi85), .B(pi27), .Y(new_n1361));
  nand_5 g1086(.A(new_n784), .B(new_n772), .Y(new_n1362));
  nand_5 g1087(.A(new_n1362), .B(new_n1361), .Y(new_n1363));
  nand_5 g1088(.A(new_n1363), .B(pi05), .Y(new_n1364));
  not_8  g1089(.A(new_n1364), .Y(new_n1365));
  or_6   g1090(.A(new_n785), .B(new_n366), .Y(new_n1366));
  nand_5 g1091(.A(new_n812), .B(new_n786), .Y(new_n1367));
  nand_5 g1092(.A(new_n1367), .B(new_n1366), .Y(new_n1368));
  nand_5 g1093(.A(new_n1368), .B(new_n359), .Y(new_n1369));
  nor_5  g1094(.A(new_n1369), .B(new_n1365), .Y(new_n1370));
  nor_5  g1095(.A(new_n1368), .B(new_n359), .Y(new_n1371));
  not_8  g1096(.A(new_n1371), .Y(new_n1372));
  nor_5  g1097(.A(new_n1363), .B(pi05), .Y(new_n1373));
  nand_5 g1098(.A(new_n1373), .B(new_n1372), .Y(new_n1374));
  nand_5 g1099(.A(new_n1365), .B(new_n1371), .Y(new_n1375));
  nand_5 g1100(.A(new_n1375), .B(new_n1374), .Y(new_n1376));
  nor_5  g1101(.A(new_n1376), .B(new_n1370), .Y(new_n1377));
  nand_5 g1102(.A(new_n1377), .B(new_n1360), .Y(new_n1378));
  not_8  g1103(.A(new_n1378), .Y(new_n1379));
  not_8  g1104(.A(new_n353), .Y(new_n1380));
  nand_5 g1105(.A(new_n1380), .B(pi83), .Y(new_n1381));
  nand_5 g1106(.A(new_n1375), .B(new_n1381), .Y(new_n1382));
  nor_5  g1107(.A(new_n1382), .B(new_n1379), .Y(new_n1383));
  nand_5 g1108(.A(new_n1383), .B(new_n1358), .Y(new_n1384));
  nor_5  g1109(.A(new_n1375), .B(new_n1381), .Y(new_n1385));
  not_8  g1110(.A(new_n1385), .Y(new_n1386));
  nor_5  g1111(.A(new_n1386), .B(new_n1358), .Y(new_n1387));
  or_6   g1112(.A(new_n1357), .B(pi53), .Y(new_n1388));
  nor_5  g1113(.A(new_n1388), .B(new_n1385), .Y(new_n1389));
  nor_5  g1114(.A(new_n1389), .B(new_n1387), .Y(new_n1390));
  nand_5 g1115(.A(new_n1390), .B(new_n1384), .Y(new_n1391));
  not_8  g1116(.A(new_n1391), .Y(new_n1392));
  nand_5 g1117(.A(new_n1392), .B(new_n1355), .Y(new_n1393));
  not_8  g1118(.A(new_n1393), .Y(new_n1394));
  nand_5 g1119(.A(new_n1339), .B(pi15), .Y(new_n1395));
  not_8  g1120(.A(new_n1387), .Y(new_n1396));
  nand_5 g1121(.A(new_n1396), .B(new_n1395), .Y(new_n1397));
  nor_5  g1122(.A(new_n1397), .B(new_n1394), .Y(new_n1398));
  or_6   g1123(.A(new_n1398), .B(new_n1354), .Y(new_n1399));
  nor_5  g1124(.A(new_n1396), .B(new_n1395), .Y(new_n1400));
  or_6   g1125(.A(new_n1400), .B(new_n1353), .Y(new_n1401));
  nand_5 g1126(.A(new_n1401), .B(new_n1399), .Y(new_n1402));
  nand_5 g1127(.A(new_n765), .B(new_n299), .Y(new_n1403));
  nor_5  g1128(.A(new_n1403), .B(new_n1402), .Y(po045));
  xnor_4 g1129(.A(po176), .B(new_n522), .Y(po046));
  not_8  g1130(.A(new_n1289), .Y(new_n1406));
  nand_5 g1131(.A(new_n1290), .B(new_n1406), .Y(new_n1407));
  nand_5 g1132(.A(new_n1407), .B(new_n1025), .Y(new_n1408));
  or_6   g1133(.A(new_n1408), .B(new_n732), .Y(new_n1409));
  not_8  g1134(.A(new_n1409), .Y(new_n1410));
  nand_5 g1135(.A(new_n1027), .B(new_n715), .Y(new_n1411));
  not_8  g1136(.A(new_n1411), .Y(new_n1412));
  not_8  g1137(.A(new_n1251), .Y(new_n1413));
  nor_5  g1138(.A(new_n1292), .B(new_n1413), .Y(new_n1414));
  nor_5  g1139(.A(new_n1414), .B(new_n1412), .Y(new_n1415));
  xor_4  g1140(.A(new_n1408), .B(new_n731), .Y(new_n1416));
  nor_5  g1141(.A(new_n1416), .B(new_n1415), .Y(new_n1417));
  nor_5  g1142(.A(new_n1417), .B(new_n1410), .Y(new_n1418));
  nor_5  g1143(.A(new_n1418), .B(new_n766), .Y(po048));
  xor_4  g1144(.A(new_n1304), .B(new_n1296), .Y(po049));
  not_8  g1145(.A(new_n1173), .Y(po050));
  xor_4  g1146(.A(new_n1270), .B(new_n1269), .Y(po051));
  xnor_4 g1147(.A(new_n1416), .B(new_n1415), .Y(po052));
  not_8  g1148(.A(new_n1175), .Y(po054));
  xor_4  g1149(.A(new_n1086), .B(new_n1202), .Y(po055));
  not_8  g1150(.A(new_n820), .Y(new_n1426));
  nor_5  g1151(.A(new_n871), .B(new_n1426), .Y(po056));
  nand_5 g1152(.A(new_n853), .B(new_n852), .Y(new_n1428));
  xor_4  g1153(.A(new_n1428), .B(new_n659), .Y(po057));
  nand_5 g1154(.A(new_n1369), .B(new_n1372), .Y(new_n1430));
  or_6   g1155(.A(new_n1365), .B(new_n1373), .Y(new_n1431));
  xor_4  g1156(.A(new_n1431), .B(new_n1430), .Y(po059));
  xor_4  g1157(.A(new_n684), .B(new_n678), .Y(po060));
  xor_4  g1158(.A(new_n1000), .B(new_n987), .Y(po061));
  nand_5 g1159(.A(new_n1344), .B(new_n814), .Y(new_n1435));
  nand_5 g1160(.A(new_n1435), .B(new_n1350), .Y(new_n1436));
  nand_5 g1161(.A(pi60), .B(pi31), .Y(new_n1437));
  nand_5 g1162(.A(pi74), .B(new_n299), .Y(new_n1438));
  nand_5 g1163(.A(new_n1438), .B(new_n1437), .Y(new_n1439));
  not_8  g1164(.A(new_n1439), .Y(new_n1440));
  nand_5 g1165(.A(new_n1440), .B(new_n1436), .Y(new_n1441));
  not_8  g1166(.A(new_n1025), .Y(new_n1442));
  not_8  g1167(.A(new_n1027), .Y(new_n1443));
  xor_4  g1168(.A(new_n1339), .B(new_n1443), .Y(new_n1444));
  nand_5 g1169(.A(new_n1357), .B(new_n1008), .Y(new_n1445));
  xor_4  g1170(.A(new_n1356), .B(new_n1009), .Y(new_n1446));
  nand_5 g1171(.A(new_n1380), .B(new_n296), .Y(new_n1447));
  nand_5 g1172(.A(new_n404), .B(new_n354), .Y(new_n1448));
  nand_5 g1173(.A(new_n1448), .B(new_n1447), .Y(new_n1449));
  nand_5 g1174(.A(new_n1449), .B(new_n1446), .Y(new_n1450));
  nand_5 g1175(.A(new_n1450), .B(new_n1445), .Y(new_n1451));
  nand_5 g1176(.A(new_n1451), .B(new_n1444), .Y(new_n1452));
  nand_5 g1177(.A(new_n1452), .B(new_n1442), .Y(new_n1453));
  nor_5  g1178(.A(new_n1452), .B(new_n1442), .Y(new_n1454));
  nand_5 g1179(.A(new_n1339), .B(new_n1443), .Y(new_n1455));
  nand_5 g1180(.A(new_n1453), .B(new_n1455), .Y(new_n1456));
  nor_5  g1181(.A(new_n1456), .B(new_n1454), .Y(new_n1457));
  nand_5 g1182(.A(new_n1457), .B(new_n1353), .Y(new_n1458));
  nand_5 g1183(.A(new_n1458), .B(new_n1453), .Y(new_n1459));
  not_8  g1184(.A(new_n1459), .Y(new_n1460));
  nor_5  g1185(.A(new_n1460), .B(new_n1441), .Y(po062));
  xnor_4 g1186(.A(new_n798), .B(new_n792), .Y(po063));
  not_8  g1187(.A(new_n514), .Y(po064));
  xor_4  g1188(.A(new_n1178), .B(new_n596), .Y(po065));
  xnor_4 g1189(.A(new_n1308), .B(new_n1307), .Y(po067));
  xor_4  g1190(.A(new_n1449), .B(new_n1446), .Y(po068));
  xor_4  g1191(.A(new_n1236), .B(new_n1235), .Y(po069));
  nand_5 g1192(.A(new_n1047), .B(new_n765), .Y(new_n1468));
  not_8  g1193(.A(new_n1468), .Y(po070));
  xor_4  g1194(.A(new_n602), .B(new_n355), .Y(new_n1470));
  nand_5 g1195(.A(new_n1277), .B(new_n1272), .Y(new_n1471));
  nand_5 g1196(.A(new_n1471), .B(new_n1273), .Y(new_n1472));
  xor_4  g1197(.A(new_n1472), .B(new_n1470), .Y(po072));
  xor_4  g1198(.A(new_n1025), .B(new_n733), .Y(new_n1474));
  not_8  g1199(.A(new_n1474), .Y(new_n1475));
  nand_5 g1200(.A(new_n1443), .B(new_n743), .Y(new_n1476));
  not_8  g1201(.A(new_n1476), .Y(new_n1477));
  nor_5  g1202(.A(new_n1312), .B(new_n1311), .Y(new_n1478));
  nor_5  g1203(.A(new_n1478), .B(new_n1477), .Y(new_n1479));
  xor_4  g1204(.A(new_n1479), .B(new_n1475), .Y(po073));
  xor_4  g1205(.A(new_n970), .B(new_n968), .Y(po074));
  xor_4  g1206(.A(new_n1136), .B(new_n438), .Y(po075));
  nand_5 g1207(.A(new_n424), .B(new_n285), .Y(new_n1483));
  nand_5 g1208(.A(new_n1483), .B(new_n414), .Y(new_n1484));
  xor_4  g1209(.A(new_n1484), .B(new_n420), .Y(po077));
  xor_4  g1210(.A(new_n1451), .B(new_n1444), .Y(po078));
  xnor_4 g1211(.A(new_n1149), .B(new_n1148), .Y(po079));
  xor_4  g1212(.A(new_n1218), .B(new_n719), .Y(po080));
  xor_4  g1213(.A(new_n1287), .B(new_n1252), .Y(po081));
  nor_5  g1214(.A(new_n1239), .B(new_n837), .Y(new_n1490));
  not_8  g1215(.A(new_n1249), .Y(new_n1491));
  nand_5 g1216(.A(new_n1491), .B(new_n1240), .Y(new_n1492));
  not_8  g1217(.A(new_n1492), .Y(new_n1493));
  nor_5  g1218(.A(new_n1493), .B(new_n1490), .Y(new_n1494));
  xor_4  g1219(.A(new_n1494), .B(new_n827), .Y(po082));
  xor_4  g1220(.A(new_n695), .B(new_n694), .Y(po083));
  not_8  g1221(.A(new_n456), .Y(new_n1497));
  nand_5 g1222(.A(new_n1497), .B(pi49), .Y(new_n1498));
  xor_4  g1223(.A(new_n1497), .B(pi49), .Y(new_n1499));
  nand_5 g1224(.A(new_n1190), .B(new_n1146), .Y(new_n1500));
  nand_5 g1225(.A(new_n1500), .B(new_n1222), .Y(new_n1501));
  nand_5 g1226(.A(new_n1501), .B(new_n1499), .Y(new_n1502));
  nand_5 g1227(.A(new_n1502), .B(new_n1498), .Y(new_n1503));
  nor_5  g1228(.A(new_n1503), .B(new_n837), .Y(new_n1504));
  xor_4  g1229(.A(new_n1501), .B(new_n1499), .Y(new_n1505));
  nor_5  g1230(.A(new_n1186), .B(pi90), .Y(new_n1506));
  nand_5 g1231(.A(new_n1192), .B(new_n1187), .Y(new_n1507));
  not_8  g1232(.A(new_n1507), .Y(new_n1508));
  nor_5  g1233(.A(new_n1508), .B(new_n1506), .Y(new_n1509));
  nand_5 g1234(.A(new_n1509), .B(new_n1505), .Y(new_n1510));
  not_8  g1235(.A(new_n1510), .Y(new_n1511));
  xor_4  g1236(.A(new_n1503), .B(new_n838), .Y(new_n1512));
  nor_5  g1237(.A(new_n1512), .B(new_n1511), .Y(new_n1513));
  nor_5  g1238(.A(new_n1513), .B(new_n1504), .Y(new_n1514));
  xor_4  g1239(.A(new_n1514), .B(new_n827), .Y(po084));
  nor_5  g1240(.A(new_n1514), .B(new_n1426), .Y(po085));
  xor_4  g1241(.A(new_n952), .B(po058), .Y(po086));
  nor_5  g1242(.A(new_n1069), .B(new_n1068), .Y(new_n1518));
  xor_4  g1243(.A(new_n1518), .B(new_n635), .Y(po087));
  nor_5  g1244(.A(new_n1041), .B(po047), .Y(new_n1520));
  xor_4  g1245(.A(new_n1041), .B(new_n1039), .Y(po117));
  nor_5  g1246(.A(po117), .B(po145), .Y(new_n1522));
  nor_5  g1247(.A(new_n1522), .B(new_n1520), .Y(po088));
  xor_4  g1248(.A(new_n838), .B(new_n828), .Y(po089));
  xor_4  g1249(.A(new_n1179), .B(new_n588), .Y(po090));
  xor_4  g1250(.A(new_n998), .B(new_n996), .Y(po091));
  not_8  g1251(.A(new_n765), .Y(new_n1527));
  nor_5  g1252(.A(new_n1048), .B(new_n1527), .Y(po092));
  xnor_4 g1253(.A(new_n402), .B(new_n401), .Y(po093));
  nand_5 g1254(.A(new_n769), .B(pi35), .Y(new_n1530));
  not_8  g1255(.A(new_n770), .Y(new_n1531));
  nand_5 g1256(.A(new_n1531), .B(new_n742), .Y(new_n1532));
  nand_5 g1257(.A(new_n1532), .B(new_n1530), .Y(new_n1533));
  nor_5  g1258(.A(new_n1533), .B(new_n754), .Y(new_n1534));
  and_6  g1259(.A(new_n1534), .B(new_n762), .Y(po094));
  xor_4  g1260(.A(new_n1283), .B(new_n1253), .Y(po095));
  xor_4  g1261(.A(new_n1440), .B(new_n1436), .Y(new_n1537));
  xor_4  g1262(.A(new_n1537), .B(new_n1459), .Y(po096));
  xor_4  g1263(.A(new_n1509), .B(new_n1505), .Y(po097));
  xor_4  g1264(.A(new_n1247), .B(new_n1243), .Y(po098));
  not_8  g1265(.A(new_n1165), .Y(po100));
  nand_5 g1266(.A(new_n763), .B(new_n756), .Y(new_n1542));
  xnor_4 g1267(.A(new_n1542), .B(new_n1534), .Y(po101));
  xor_4  g1268(.A(new_n1512), .B(new_n1510), .Y(po102));
  xor_4  g1269(.A(new_n744), .B(new_n741), .Y(po103));
  and_6  g1270(.A(new_n1514), .B(new_n825), .Y(new_n1546));
  or_6   g1271(.A(new_n1546), .B(po085), .Y(po104));
  xor_4  g1272(.A(new_n524), .B(new_n514), .Y(po105));
  xor_4  g1273(.A(new_n422), .B(new_n379), .Y(po106));
  xor_4  g1274(.A(new_n1217), .B(new_n587), .Y(po107));
  not_8  g1275(.A(new_n1047), .Y(new_n1551));
  not_8  g1276(.A(pi74), .Y(new_n1552));
  nand_5 g1277(.A(new_n1034), .B(new_n1031), .Y(new_n1553));
  nand_5 g1278(.A(new_n1553), .B(new_n1030), .Y(new_n1554));
  nor_5  g1279(.A(new_n1554), .B(new_n1552), .Y(new_n1555));
  nand_5 g1280(.A(new_n1555), .B(new_n1551), .Y(new_n1556));
  nand_5 g1281(.A(new_n1556), .B(new_n1468), .Y(po108));
  xor_4  g1282(.A(new_n867), .B(new_n466), .Y(po109));
  xor_4  g1283(.A(new_n1537), .B(new_n1402), .Y(new_n1559));
  not_8  g1284(.A(new_n1559), .Y(po135));
  not_8  g1285(.A(new_n1438), .Y(new_n1561));
  nand_5 g1286(.A(new_n1561), .B(new_n764), .Y(new_n1562));
  and_6  g1287(.A(new_n1562), .B(new_n1437), .Y(new_n1563));
  nor_5  g1288(.A(new_n1563), .B(po135), .Y(new_n1564));
  or_6   g1289(.A(new_n1564), .B(po045), .Y(po110));
  xor_4  g1290(.A(new_n870), .B(new_n838), .Y(po111));
  or_6   g1291(.A(new_n1440), .B(new_n1436), .Y(new_n1567));
  nor_5  g1292(.A(new_n1567), .B(new_n1459), .Y(new_n1568));
  or_6   g1293(.A(new_n1568), .B(po062), .Y(po112));
  xor_4  g1294(.A(new_n1180), .B(new_n715), .Y(po114));
  nand_5 g1295(.A(new_n518), .B(new_n496), .Y(po123));
  not_8  g1296(.A(po123), .Y(po115));
  nand_5 g1297(.A(new_n1025), .B(new_n733), .Y(new_n1573));
  not_8  g1298(.A(new_n1573), .Y(new_n1574));
  nor_5  g1299(.A(new_n1479), .B(new_n1475), .Y(new_n1575));
  nor_5  g1300(.A(new_n1575), .B(new_n1574), .Y(new_n1576));
  nand_5 g1301(.A(new_n1576), .B(new_n770), .Y(new_n1577));
  nor_5  g1302(.A(new_n1577), .B(new_n763), .Y(po165));
  nor_5  g1303(.A(new_n1576), .B(new_n1542), .Y(new_n1579));
  or_6   g1304(.A(new_n1579), .B(po165), .Y(po116));
  xor_4  g1305(.A(new_n399), .B(new_n398), .Y(po118));
  xnor_4 g1306(.A(new_n1265), .B(new_n1257), .Y(po119));
  xor_4  g1307(.A(new_n1428), .B(new_n658), .Y(po120));
  xor_4  g1308(.A(new_n1173), .B(new_n1172), .Y(po121));
  xor_4  g1309(.A(new_n1045), .B(new_n1035), .Y(po122));
  xor_4  g1310(.A(new_n1219), .B(new_n731), .Y(po124));
  and_6  g1311(.A(new_n1086), .B(new_n763), .Y(new_n1587));
  or_6   g1312(.A(new_n1587), .B(po023), .Y(po126));
  xor_4  g1313(.A(new_n1181), .B(new_n732), .Y(po127));
  nor_5  g1314(.A(new_n1494), .B(new_n1426), .Y(po128));
  xor_4  g1315(.A(new_n383), .B(new_n377), .Y(po129));
  and_6  g1316(.A(new_n1555), .B(new_n1048), .Y(new_n1592));
  or_6   g1317(.A(new_n1592), .B(po092), .Y(po130));
  and_6  g1318(.A(new_n513), .B(new_n511), .Y(po177));
  xnor_4 g1319(.A(po177), .B(new_n525), .Y(po131));
  xor_4  g1320(.A(new_n1392), .B(new_n1355), .Y(po132));
  xor_4  g1321(.A(new_n1302), .B(new_n1301), .Y(po133));
  xor_4  g1322(.A(new_n667), .B(new_n666), .Y(po134));
  and_6  g1323(.A(new_n871), .B(new_n825), .Y(new_n1599));
  or_6   g1324(.A(new_n1599), .B(po056), .Y(po136));
  xor_4  g1325(.A(new_n1142), .B(new_n1120), .Y(po137));
  xor_4  g1326(.A(new_n1554), .B(new_n1552), .Y(new_n1602));
  xor_4  g1327(.A(new_n1602), .B(new_n1047), .Y(po138));
  nand_5 g1328(.A(po138), .B(po047), .Y(new_n1604));
  nand_5 g1329(.A(new_n1602), .B(po145), .Y(new_n1605));
  nand_5 g1330(.A(new_n1605), .B(new_n1604), .Y(po139));
  xor_4  g1331(.A(new_n512), .B(new_n866), .Y(po140));
  xor_4  g1332(.A(new_n1377), .B(new_n1360), .Y(po141));
  xor_4  g1333(.A(new_n1263), .B(new_n1260), .Y(po142));
  xnor_4 g1334(.A(new_n1065), .B(new_n1054), .Y(po143));
  nand_5 g1335(.A(new_n1220), .B(new_n763), .Y(new_n1611));
  nand_5 g1336(.A(new_n1611), .B(new_n1162), .Y(po144));
  nor_5  g1337(.A(new_n839), .B(new_n1426), .Y(po146));
  xor_4  g1338(.A(new_n498), .B(new_n496), .Y(po148));
  xnor_4 g1339(.A(new_n1063), .B(new_n1056), .Y(po149));
  xor_4  g1340(.A(new_n1576), .B(new_n1531), .Y(po150));
  nor_5  g1341(.A(new_n1044), .B(po047), .Y(new_n1617));
  nor_5  g1342(.A(po044), .B(po145), .Y(new_n1618));
  nor_5  g1343(.A(new_n1618), .B(new_n1617), .Y(po151));
  xor_4  g1344(.A(new_n1061), .B(pi33), .Y(po152));
  xor_4  g1345(.A(new_n641), .B(new_n639), .Y(new_n1621));
  xnor_4 g1346(.A(new_n1621), .B(new_n670), .Y(po153));
  xnor_4 g1347(.A(new_n966), .B(new_n965), .Y(po154));
  nand_5 g1348(.A(new_n1388), .B(new_n1358), .Y(new_n1624));
  or_6   g1349(.A(new_n1385), .B(new_n1383), .Y(new_n1625));
  xor_4  g1350(.A(new_n1625), .B(new_n1624), .Y(po155));
  xor_4  g1351(.A(new_n1139), .B(new_n1124), .Y(po156));
  xor_4  g1352(.A(new_n1171), .B(po172), .Y(po157));
  xnor_4 g1353(.A(new_n672), .B(new_n637), .Y(po158));
  xor_4  g1354(.A(po162), .B(po145), .Y(po159));
  and_6  g1355(.A(new_n839), .B(new_n825), .Y(new_n1631));
  or_6   g1356(.A(new_n1631), .B(po146), .Y(po160));
  xnor_4 g1357(.A(new_n1267), .B(new_n1255), .Y(po161));
  xor_4  g1358(.A(new_n518), .B(new_n498), .Y(po163));
  xnor_4 g1359(.A(new_n1132), .B(new_n1128), .Y(po164));
  nand_5 g1360(.A(po162), .B(po145), .Y(new_n1636));
  xor_4  g1361(.A(new_n1636), .B(new_n906), .Y(po166));
  xnor_4 g1362(.A(new_n1233), .B(new_n1225), .Y(po167));
  xor_4  g1363(.A(new_n528), .B(new_n467), .Y(po168));
  and_6  g1364(.A(new_n1494), .B(new_n825), .Y(new_n1640));
  or_6   g1365(.A(new_n1640), .B(po128), .Y(po169));
  xor_4  g1366(.A(new_n958), .B(new_n948), .Y(po170));
  xor_4  g1367(.A(new_n1418), .B(new_n1202), .Y(po173));
  xor_4  g1368(.A(new_n1060), .B(new_n1058), .Y(po174));
  nor_5  g1369(.A(new_n1400), .B(new_n1398), .Y(new_n1645));
  xor_4  g1370(.A(new_n1645), .B(new_n1353), .Y(po175));
  xor_4  g1371(.A(new_n1457), .B(new_n1354), .Y(po178));
  xor_4  g1372(.A(new_n869), .B(new_n456), .Y(po179));
  and_6  g1373(.A(new_n1418), .B(new_n763), .Y(new_n1649));
  or_6   g1374(.A(new_n1649), .B(po048), .Y(po180));
  xnor_4 g1375(.A(new_n1231), .B(new_n1230), .Y(po181));
  buf_8  g1376(.A(po012), .Y(po039));
  buf_8  g1377(.A(po022), .Y(po171));
endmodule


