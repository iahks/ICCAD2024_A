// Benchmark "top_809568696_809776567_809698999_863110837_1234615" written by ABC on Mon Aug 19 00:27:35 2024

module top_809568696_809776567_809698999_863110837_1234615 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128;
  wire new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1955, new_n1956, new_n1957, new_n1958, new_n1959, new_n1960,
    new_n1961, new_n1962, new_n1963, new_n1964, new_n1965, new_n1966,
    new_n1967, new_n1968, new_n1969, new_n1970, new_n1971, new_n1972,
    new_n1973, new_n1974, new_n1975, new_n1976, new_n1977, new_n1978,
    new_n1979, new_n1980, new_n1981, new_n1982, new_n1983, new_n1984,
    new_n1985, new_n1986, new_n1987, new_n1988, new_n1989, new_n1990,
    new_n1991, new_n1992, new_n1993, new_n1994, new_n1995, new_n1996,
    new_n1997, new_n1998, new_n1999, new_n2000, new_n2001, new_n2002,
    new_n2003, new_n2004, new_n2005, new_n2006, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2154, new_n2155, new_n2156,
    new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252,
    new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2347, new_n2348, new_n2349, new_n2350,
    new_n2351, new_n2352, new_n2353, new_n2354, new_n2355, new_n2356,
    new_n2357, new_n2358, new_n2359, new_n2360, new_n2361, new_n2362,
    new_n2363, new_n2364, new_n2365, new_n2366, new_n2367, new_n2368,
    new_n2369, new_n2370, new_n2371, new_n2372, new_n2373, new_n2374,
    new_n2375, new_n2376, new_n2377, new_n2378, new_n2379, new_n2381,
    new_n2382, new_n2383, new_n2384, new_n2385, new_n2386, new_n2387,
    new_n2388, new_n2389, new_n2390, new_n2391, new_n2392, new_n2393,
    new_n2394, new_n2395, new_n2396, new_n2397, new_n2398, new_n2399,
    new_n2400, new_n2401, new_n2402, new_n2403, new_n2404, new_n2405,
    new_n2406, new_n2407, new_n2408, new_n2409, new_n2410, new_n2411,
    new_n2412, new_n2413, new_n2414, new_n2415, new_n2416, new_n2417,
    new_n2418, new_n2419, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430,
    new_n2431, new_n2432, new_n2434, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2509, new_n2510, new_n2511, new_n2512,
    new_n2513, new_n2514, new_n2515, new_n2516, new_n2517, new_n2518,
    new_n2519, new_n2520, new_n2522, new_n2523, new_n2524, new_n2525,
    new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2532,
    new_n2533, new_n2534, new_n2535, new_n2536, new_n2537, new_n2538,
    new_n2539, new_n2540, new_n2541, new_n2542, new_n2543, new_n2544,
    new_n2545, new_n2546, new_n2548, new_n2549, new_n2550, new_n2551,
    new_n2553, new_n2554, new_n2555, new_n2557, new_n2559, new_n2560,
    new_n2561, new_n2562, new_n2563, new_n2564, new_n2565, new_n2566,
    new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2573,
    new_n2574, new_n2575, new_n2576, new_n2577, new_n2578, new_n2580,
    new_n2581, new_n2582, new_n2583, new_n2584, new_n2586, new_n2587,
    new_n2588, new_n2589, new_n2590, new_n2591, new_n2592, new_n2593,
    new_n2594, new_n2595, new_n2596, new_n2597, new_n2598, new_n2599,
    new_n2600, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2644, new_n2645,
    new_n2646, new_n2647, new_n2650, new_n2651, new_n2652, new_n2653,
    new_n2654, new_n2656, new_n2657, new_n2659, new_n2660, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2683, new_n2684, new_n2686, new_n2687, new_n2688,
    new_n2689, new_n2690, new_n2692, new_n2693, new_n2694, new_n2695,
    new_n2696, new_n2697, new_n2698, new_n2699, new_n2700, new_n2701,
    new_n2702, new_n2703, new_n2704, new_n2705, new_n2706, new_n2707,
    new_n2708, new_n2709, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2716, new_n2717, new_n2718, new_n2719, new_n2721, new_n2722,
    new_n2723, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2739, new_n2740, new_n2741, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2768, new_n2769,
    new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775,
    new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781,
    new_n2782, new_n2783, new_n2784, new_n2785, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2793, new_n2794, new_n2795, new_n2796,
    new_n2797, new_n2798, new_n2799, new_n2800, new_n2801, new_n2802,
    new_n2803, new_n2804, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2816, new_n2817,
    new_n2818, new_n2819, new_n2820, new_n2821, new_n2822, new_n2823,
    new_n2824, new_n2825, new_n2826, new_n2827, new_n2828, new_n2829,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2838, new_n2839, new_n2841, new_n2842, new_n2844, new_n2845,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2852, new_n2853,
    new_n2854, new_n2855, new_n2856, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2881, new_n2882, new_n2883, new_n2884, new_n2886,
    new_n2888, new_n2889, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2896, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2920, new_n2922, new_n2924, new_n2925,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2941, new_n2942, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2956, new_n2957, new_n2958, new_n2959,
    new_n2960, new_n2962, new_n2964, new_n2965, new_n2966, new_n2968,
    new_n2969, new_n2970, new_n2972, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2979, new_n2980, new_n2983, new_n2984, new_n2986,
    new_n2988, new_n2990, new_n2991, new_n2993, new_n2994, new_n2996,
    new_n2997, new_n2999, new_n3000, new_n3001, new_n3003, new_n3005,
    new_n3006, new_n3008, new_n3010, new_n3011, new_n3012, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3020, new_n3021,
    new_n3022, new_n3025, new_n3026, new_n3027, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3034, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3042, new_n3044, new_n3045, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3055,
    new_n3056, new_n3058, new_n3060, new_n3061, new_n3062, new_n3064,
    new_n3066, new_n3067, new_n3069, new_n3071, new_n3073, new_n3074,
    new_n3076, new_n3077, new_n3078, new_n3081, new_n3082, new_n3084,
    new_n3085, new_n3086, new_n3088, new_n3089, new_n3092, new_n3095,
    new_n3096, new_n3098, new_n3101, new_n3102, new_n3106, new_n3108,
    new_n3109, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115;
  nand_5 g0000(.A(pi238), .B(pi238), .Y(new_n386));
  nand_5 g0001(.A(pi060), .B(pi060), .Y(new_n387));
  nand_5 g0002(.A(pi200), .B(pi200), .Y(new_n388));
  nand_5     g0003(.A(new_n388), .B(new_n387), .Y(new_n389));
  nand_5 g0004(.A(new_n389), .B(new_n389), .Y(new_n390));
  nand_5 g0005(.A(pi094), .B(pi094), .Y(new_n391));
  nand_5 g0006(.A(pi146), .B(pi146), .Y(new_n392));
  nand_5     g0007(.A(new_n392), .B(pi128), .Y(new_n393));
  nand_5     g0008(.A(new_n393), .B(new_n391), .Y(new_n394));
  nand_5 g0009(.A(new_n394), .B(new_n394), .Y(new_n395));
  nand_5     g0010(.A(new_n395), .B(new_n390), .Y(new_n396));
  nand_5 g0011(.A(new_n396), .B(new_n396), .Y(new_n397));
  nand_5 g0012(.A(pi246), .B(pi246), .Y(new_n398));
  nand_5     g0013(.A(new_n398), .B(new_n392), .Y(new_n399));
  nand_5 g0014(.A(new_n399), .B(new_n399), .Y(new_n400));
  nand_5     g0015(.A(new_n400), .B(pi117), .Y(new_n401));
  nand_5     g0016(.A(new_n401), .B(new_n397), .Y(new_n402));
  nand_5 g0017(.A(pi171), .B(pi171), .Y(new_n403));
  nand_5     g0018(.A(pi226), .B(new_n388), .Y(new_n404));
  nand_5     g0019(.A(new_n404), .B(new_n403), .Y(new_n405));
  nand_5 g0020(.A(new_n405), .B(new_n405), .Y(new_n406));
  nand_5     g0021(.A(new_n406), .B(new_n402), .Y(new_n407));
  nand_5 g0022(.A(pi103), .B(pi103), .Y(new_n408));
  nand_5 g0023(.A(pi153), .B(pi153), .Y(new_n409));
  nand_5     g0024(.A(new_n409), .B(new_n408), .Y(new_n410));
  nand_5 g0025(.A(pi021), .B(pi021), .Y(new_n411));
  nand_5     g0026(.A(new_n387), .B(new_n411), .Y(new_n412));
  nor_5      g0027(.A(new_n412), .B(new_n410), .Y(new_n413));
  nand_5 g0028(.A(new_n413), .B(new_n413), .Y(new_n414));
  nand_5 g0029(.A(pi182), .B(pi182), .Y(new_n415));
  nand_5 g0030(.A(pi144), .B(pi144), .Y(new_n416));
  nand_5 g0031(.A(pi077), .B(pi077), .Y(new_n417));
  nand_5 g0032(.A(pi090), .B(pi090), .Y(new_n418));
  nand_5     g0033(.A(new_n418), .B(new_n417), .Y(new_n419));
  nand_5 g0034(.A(new_n419), .B(new_n419), .Y(new_n420));
  nand_5     g0035(.A(new_n420), .B(new_n416), .Y(new_n421));
  nand_5 g0036(.A(new_n421), .B(new_n421), .Y(new_n422));
  nand_5     g0037(.A(new_n422), .B(new_n415), .Y(new_n423));
  nor_5      g0038(.A(new_n423), .B(new_n414), .Y(new_n424));
  nand_5     g0039(.A(new_n424), .B(new_n407), .Y(new_n425));
  nand_5 g0040(.A(new_n425), .B(new_n425), .Y(new_n426));
  nor_5      g0041(.A(pi098), .B(pi069), .Y(new_n427));
  nand_5 g0042(.A(pi223), .B(pi223), .Y(new_n428));
  nand_5 g0043(.A(pi069), .B(pi069), .Y(new_n429));
  nand_5     g0044(.A(pi220), .B(new_n429), .Y(new_n430));
  nand_5     g0045(.A(new_n430), .B(new_n428), .Y(new_n431));
  nor_5      g0046(.A(new_n431), .B(new_n427), .Y(new_n432));
  nor_5      g0047(.A(new_n432), .B(pi120), .Y(new_n433));
  nand_5 g0048(.A(pi156), .B(pi156), .Y(new_n434));
  nor_5      g0049(.A(pi076), .B(pi049), .Y(new_n435));
  nand_5     g0050(.A(new_n435), .B(new_n434), .Y(new_n436));
  nand_5 g0051(.A(new_n436), .B(new_n436), .Y(new_n437));
  nand_5 g0052(.A(pi239), .B(pi239), .Y(new_n438));
  nand_5 g0053(.A(pi204), .B(pi204), .Y(new_n439));
  nand_5     g0054(.A(new_n439), .B(pi010), .Y(new_n440));
  nand_5     g0055(.A(new_n440), .B(new_n438), .Y(new_n441));
  nand_5     g0056(.A(new_n441), .B(new_n437), .Y(new_n442));
  nand_5 g0057(.A(pi237), .B(pi237), .Y(new_n443));
  nor_5      g0058(.A(new_n443), .B(pi049), .Y(new_n444));
  nor_5      g0059(.A(new_n444), .B(pi030), .Y(new_n445));
  nor_5      g0060(.A(new_n445), .B(pi156), .Y(new_n446));
  nand_5 g0061(.A(pi159), .B(pi159), .Y(new_n447));
  nand_5 g0062(.A(pi220), .B(pi220), .Y(new_n448));
  nand_5     g0063(.A(new_n448), .B(new_n447), .Y(new_n449));
  nand_5 g0064(.A(new_n449), .B(new_n449), .Y(new_n450));
  nand_5     g0065(.A(new_n450), .B(new_n428), .Y(new_n451));
  nor_5      g0066(.A(new_n451), .B(new_n446), .Y(new_n452));
  nand_5     g0067(.A(new_n452), .B(new_n442), .Y(new_n453));
  nand_5     g0068(.A(new_n453), .B(new_n433), .Y(new_n454));
  nand_5 g0069(.A(pi016), .B(pi016), .Y(new_n455));
  nand_5 g0070(.A(pi056), .B(pi056), .Y(new_n456));
  nand_5     g0071(.A(new_n456), .B(new_n455), .Y(new_n457));
  nand_5 g0072(.A(pi126), .B(pi126), .Y(new_n458));
  nand_5 g0073(.A(pi139), .B(pi139), .Y(new_n459));
  nand_5 g0074(.A(pi232), .B(pi232), .Y(new_n460));
  nand_5     g0075(.A(new_n460), .B(new_n459), .Y(new_n461));
  nand_5 g0076(.A(new_n461), .B(new_n461), .Y(new_n462));
  nand_5     g0077(.A(new_n462), .B(new_n458), .Y(new_n463));
  nor_5      g0078(.A(new_n463), .B(new_n457), .Y(new_n464));
  nand_5     g0079(.A(new_n464), .B(new_n454), .Y(new_n465));
  nand_5 g0080(.A(pi178), .B(pi178), .Y(new_n466));
  nor_5      g0081(.A(new_n461), .B(new_n466), .Y(new_n467));
  nand_5 g0082(.A(pi012), .B(pi012), .Y(new_n468));
  nand_5     g0083(.A(pi207), .B(new_n459), .Y(new_n469));
  nand_5     g0084(.A(new_n469), .B(new_n468), .Y(new_n470));
  nor_5      g0085(.A(new_n470), .B(new_n467), .Y(new_n471));
  nor_5      g0086(.A(new_n471), .B(new_n457), .Y(new_n472));
  nand_5 g0087(.A(pi082), .B(pi082), .Y(new_n473));
  nand_5 g0088(.A(pi011), .B(pi011), .Y(new_n474));
  nand_5     g0089(.A(pi056), .B(new_n474), .Y(new_n475));
  nand_5 g0090(.A(pi152), .B(pi152), .Y(new_n476));
  nand_5     g0091(.A(new_n476), .B(new_n474), .Y(new_n477));
  nand_5     g0092(.A(new_n477), .B(new_n475), .Y(new_n478));
  nand_5     g0093(.A(new_n478), .B(new_n473), .Y(new_n479));
  nor_5      g0094(.A(new_n479), .B(new_n472), .Y(new_n480));
  nand_5     g0095(.A(new_n480), .B(new_n465), .Y(new_n481));
  nor_5      g0096(.A(pi253), .B(pi227), .Y(new_n482));
  nand_5 g0097(.A(pi255), .B(pi255), .Y(new_n483));
  nand_5     g0098(.A(new_n483), .B(pi252), .Y(new_n484));
  nand_5 g0099(.A(pi125), .B(pi125), .Y(new_n485));
  nand_5 g0100(.A(pi251), .B(pi251), .Y(new_n486));
  nand_5     g0101(.A(new_n486), .B(new_n485), .Y(new_n487));
  nand_5 g0102(.A(new_n487), .B(new_n487), .Y(new_n488));
  nand_5     g0103(.A(new_n488), .B(new_n484), .Y(new_n489));
  nor_5      g0104(.A(new_n489), .B(pi176), .Y(new_n490));
  nand_5     g0105(.A(new_n490), .B(new_n482), .Y(new_n491));
  nand_5 g0106(.A(new_n491), .B(new_n491), .Y(new_n492));
  nor_5      g0107(.A(pi190), .B(pi025), .Y(new_n493));
  nand_5 g0108(.A(pi165), .B(pi165), .Y(new_n494));
  nor_5      g0109(.A(pi190), .B(new_n494), .Y(new_n495));
  nor_5      g0110(.A(new_n495), .B(new_n493), .Y(new_n496));
  nor_5      g0111(.A(new_n496), .B(pi007), .Y(new_n497));
  nand_5 g0112(.A(pi155), .B(pi155), .Y(new_n498));
  nor_5      g0113(.A(pi141), .B(pi047), .Y(new_n499));
  nand_5     g0114(.A(new_n499), .B(new_n498), .Y(new_n500));
  nand_5     g0115(.A(new_n499), .B(pi198), .Y(new_n501));
  nand_5     g0116(.A(new_n501), .B(new_n500), .Y(new_n502));
  nand_5     g0117(.A(new_n502), .B(new_n497), .Y(new_n503));
  nand_5 g0118(.A(pi143), .B(pi143), .Y(new_n504));
  nand_5     g0119(.A(new_n494), .B(new_n504), .Y(new_n505));
  nand_5     g0120(.A(new_n505), .B(new_n497), .Y(new_n506));
  nand_5 g0121(.A(pi066), .B(pi066), .Y(new_n507));
  nand_5 g0122(.A(pi007), .B(pi007), .Y(new_n508));
  nand_5     g0123(.A(pi199), .B(new_n508), .Y(new_n509));
  nand_5     g0124(.A(new_n509), .B(new_n507), .Y(new_n510));
  nand_5 g0125(.A(new_n510), .B(new_n510), .Y(new_n511));
  nand_5     g0126(.A(new_n511), .B(new_n506), .Y(new_n512));
  nand_5 g0127(.A(pi092), .B(pi092), .Y(new_n513));
  nor_5      g0128(.A(pi141), .B(new_n513), .Y(new_n514));
  nand_5     g0129(.A(new_n514), .B(new_n497), .Y(new_n515));
  nor_5      g0130(.A(pi215), .B(pi041), .Y(new_n516));
  nand_5 g0131(.A(pi050), .B(pi050), .Y(new_n517));
  nand_5 g0132(.A(pi079), .B(pi079), .Y(new_n518));
  nand_5     g0133(.A(new_n518), .B(new_n517), .Y(new_n519));
  nand_5 g0134(.A(new_n519), .B(new_n519), .Y(new_n520));
  nand_5     g0135(.A(new_n520), .B(new_n516), .Y(new_n521));
  nand_5 g0136(.A(new_n521), .B(new_n521), .Y(new_n522));
  nand_5     g0137(.A(new_n522), .B(new_n515), .Y(new_n523));
  nor_5      g0138(.A(new_n523), .B(new_n512), .Y(new_n524));
  nand_5     g0139(.A(new_n524), .B(new_n503), .Y(new_n525));
  nand_5 g0140(.A(new_n525), .B(new_n525), .Y(new_n526));
  nand_5     g0141(.A(new_n526), .B(new_n492), .Y(new_n527));
  nand_5 g0142(.A(pi067), .B(pi067), .Y(new_n528));
  nand_5     g0143(.A(pi079), .B(new_n528), .Y(new_n529));
  nand_5 g0144(.A(pi109), .B(pi109), .Y(new_n530));
  nand_5     g0145(.A(new_n530), .B(new_n528), .Y(new_n531));
  nand_5     g0146(.A(new_n531), .B(new_n529), .Y(new_n532));
  nand_5     g0147(.A(new_n532), .B(new_n483), .Y(new_n533));
  nand_5 g0148(.A(new_n516), .B(new_n516), .Y(new_n534));
  nand_5 g0149(.A(pi228), .B(pi228), .Y(new_n535));
  nor_5      g0150(.A(new_n535), .B(pi215), .Y(new_n536));
  nor_5      g0151(.A(new_n536), .B(pi105), .Y(new_n537));
  nand_5     g0152(.A(new_n537), .B(new_n534), .Y(new_n538));
  nand_5     g0153(.A(new_n538), .B(new_n520), .Y(new_n539));
  nand_5 g0154(.A(pi105), .B(pi105), .Y(new_n540));
  nand_5 g0155(.A(pi183), .B(pi183), .Y(new_n541));
  nand_5     g0156(.A(new_n535), .B(new_n541), .Y(new_n542));
  nand_5 g0157(.A(new_n542), .B(new_n542), .Y(new_n543));
  nand_5     g0158(.A(new_n543), .B(new_n540), .Y(new_n544));
  nand_5 g0159(.A(new_n544), .B(new_n544), .Y(new_n545));
  nor_5      g0160(.A(new_n545), .B(new_n539), .Y(new_n546));
  nor_5      g0161(.A(new_n546), .B(new_n533), .Y(new_n547));
  nor_5      g0162(.A(new_n547), .B(new_n491), .Y(new_n548));
  nand_5 g0163(.A(pi120), .B(pi120), .Y(new_n549));
  nand_5     g0164(.A(new_n427), .B(new_n434), .Y(new_n550));
  nand_5 g0165(.A(new_n550), .B(new_n550), .Y(new_n551));
  nand_5     g0166(.A(new_n551), .B(new_n435), .Y(new_n552));
  nand_5 g0167(.A(new_n552), .B(new_n552), .Y(new_n553));
  nand_5     g0168(.A(new_n553), .B(new_n549), .Y(new_n554));
  nor_5      g0169(.A(pi210), .B(pi138), .Y(new_n555));
  nand_5 g0170(.A(new_n555), .B(new_n555), .Y(new_n556));
  nor_5      g0171(.A(new_n556), .B(pi242), .Y(new_n557));
  nand_5 g0172(.A(new_n557), .B(new_n557), .Y(new_n558));
  nand_5     g0173(.A(new_n555), .B(pi125), .Y(new_n559));
  nand_5 g0174(.A(new_n559), .B(new_n559), .Y(new_n560));
  nand_5 g0175(.A(pi176), .B(pi176), .Y(new_n561));
  nor_5      g0176(.A(new_n561), .B(pi138), .Y(new_n562));
  nand_5 g0177(.A(new_n562), .B(new_n562), .Y(new_n563));
  nand_5     g0178(.A(new_n563), .B(new_n482), .Y(new_n564));
  nor_5      g0179(.A(new_n564), .B(new_n560), .Y(new_n565));
  nand_5     g0180(.A(new_n565), .B(new_n558), .Y(new_n566));
  nand_5 g0181(.A(pi115), .B(pi115), .Y(new_n567));
  nand_5 g0182(.A(pi227), .B(pi227), .Y(new_n568));
  nand_5     g0183(.A(new_n568), .B(pi214), .Y(new_n569));
  nand_5     g0184(.A(new_n569), .B(new_n567), .Y(new_n570));
  nor_5      g0185(.A(new_n570), .B(pi204), .Y(new_n571));
  nand_5     g0186(.A(new_n571), .B(new_n566), .Y(new_n572));
  nor_5      g0187(.A(new_n572), .B(new_n554), .Y(new_n573));
  nand_5     g0188(.A(new_n573), .B(new_n480), .Y(new_n574));
  nor_5      g0189(.A(new_n574), .B(new_n548), .Y(new_n575));
  nand_5     g0190(.A(new_n575), .B(new_n527), .Y(new_n576));
  nand_5 g0191(.A(new_n576), .B(new_n576), .Y(new_n577));
  nand_5 g0192(.A(pi219), .B(pi219), .Y(new_n578));
  nand_5 g0193(.A(pi163), .B(pi163), .Y(new_n579));
  nand_5 g0194(.A(pi248), .B(pi248), .Y(new_n580));
  nand_5     g0195(.A(new_n580), .B(new_n579), .Y(new_n581));
  nand_5 g0196(.A(new_n581), .B(new_n581), .Y(new_n582));
  nand_5     g0197(.A(new_n582), .B(new_n578), .Y(new_n583));
  nand_5 g0198(.A(new_n583), .B(new_n583), .Y(new_n584));
  nand_5 g0199(.A(pi166), .B(pi166), .Y(new_n585));
  nand_5 g0200(.A(pi123), .B(pi123), .Y(new_n586));
  nand_5     g0201(.A(pi187), .B(new_n586), .Y(new_n587));
  nand_5     g0202(.A(new_n587), .B(new_n585), .Y(new_n588));
  nand_5 g0203(.A(new_n588), .B(new_n588), .Y(new_n589));
  nor_5      g0204(.A(pi189), .B(pi129), .Y(new_n590));
  nand_5 g0205(.A(new_n590), .B(new_n590), .Y(new_n591));
  nor_5      g0206(.A(pi123), .B(pi057), .Y(new_n592));
  nand_5 g0207(.A(new_n592), .B(new_n592), .Y(new_n593));
  nand_5 g0208(.A(pi194), .B(pi194), .Y(new_n594));
  nor_5      g0209(.A(new_n594), .B(pi129), .Y(new_n595));
  nor_5      g0210(.A(new_n595), .B(new_n593), .Y(new_n596));
  nand_5     g0211(.A(new_n596), .B(new_n591), .Y(new_n597));
  nand_5     g0212(.A(new_n597), .B(new_n589), .Y(new_n598));
  nor_5      g0213(.A(new_n598), .B(pi136), .Y(new_n599));
  nand_5 g0214(.A(pi164), .B(pi164), .Y(new_n600));
  nand_5     g0215(.A(new_n594), .B(new_n600), .Y(new_n601));
  nand_5 g0216(.A(new_n601), .B(new_n601), .Y(new_n602));
  nand_5     g0217(.A(new_n602), .B(new_n592), .Y(new_n603));
  nand_5 g0218(.A(new_n603), .B(new_n603), .Y(new_n604));
  nand_5 g0219(.A(pi111), .B(pi111), .Y(new_n605));
  nand_5 g0220(.A(pi224), .B(pi224), .Y(new_n606));
  nand_5     g0221(.A(new_n606), .B(new_n605), .Y(new_n607));
  nand_5 g0222(.A(pi108), .B(pi108), .Y(new_n608));
  nand_5     g0223(.A(pi185), .B(new_n605), .Y(new_n609));
  nand_5     g0224(.A(new_n609), .B(new_n608), .Y(new_n610));
  nand_5 g0225(.A(new_n610), .B(new_n610), .Y(new_n611));
  nand_5     g0226(.A(new_n611), .B(new_n607), .Y(new_n612));
  nand_5     g0227(.A(new_n612), .B(new_n604), .Y(new_n613));
  nand_5     g0228(.A(new_n613), .B(new_n599), .Y(new_n614));
  nand_5 g0229(.A(new_n614), .B(new_n614), .Y(new_n615));
  nand_5     g0230(.A(new_n615), .B(new_n584), .Y(new_n616));
  nand_5 g0231(.A(pi169), .B(pi169), .Y(new_n617));
  nand_5 g0232(.A(pi192), .B(pi192), .Y(new_n618));
  nand_5     g0233(.A(new_n618), .B(pi118), .Y(new_n619));
  nor_5      g0234(.A(pi217), .B(pi192), .Y(new_n620));
  nand_5 g0235(.A(new_n620), .B(new_n620), .Y(new_n621));
  nand_5     g0236(.A(new_n621), .B(new_n619), .Y(new_n622));
  nand_5     g0237(.A(new_n622), .B(new_n617), .Y(new_n623));
  nand_5 g0238(.A(pi100), .B(pi100), .Y(new_n624));
  nor_5      g0239(.A(pi167), .B(pi017), .Y(new_n625));
  nor_5      g0240(.A(pi113), .B(pi068), .Y(new_n626));
  nand_5     g0241(.A(new_n626), .B(new_n625), .Y(new_n627));
  nand_5 g0242(.A(new_n627), .B(new_n627), .Y(new_n628));
  nand_5     g0243(.A(new_n628), .B(new_n624), .Y(new_n629));
  nand_5 g0244(.A(new_n629), .B(new_n629), .Y(new_n630));
  nand_5     g0245(.A(new_n580), .B(pi026), .Y(new_n631));
  nand_5     g0246(.A(new_n631), .B(new_n630), .Y(new_n632));
  nand_5 g0247(.A(new_n632), .B(new_n632), .Y(new_n633));
  nand_5 g0248(.A(pi089), .B(pi089), .Y(new_n634));
  nor_5      g0249(.A(pi102), .B(pi042), .Y(new_n635));
  nand_5 g0250(.A(new_n635), .B(new_n635), .Y(new_n636));
  nand_5 g0251(.A(pi136), .B(pi136), .Y(new_n637));
  nor_5      g0252(.A(new_n637), .B(pi042), .Y(new_n638));
  nand_5 g0253(.A(new_n638), .B(new_n638), .Y(new_n639));
  nand_5     g0254(.A(new_n639), .B(new_n636), .Y(new_n640));
  nand_5     g0255(.A(new_n640), .B(new_n634), .Y(new_n641));
  nand_5     g0256(.A(pi219), .B(new_n634), .Y(new_n642));
  nand_5     g0257(.A(new_n642), .B(new_n582), .Y(new_n643));
  nand_5 g0258(.A(new_n643), .B(new_n643), .Y(new_n644));
  nand_5     g0259(.A(new_n644), .B(new_n641), .Y(new_n645));
  nand_5     g0260(.A(new_n645), .B(new_n633), .Y(new_n646));
  nor_5      g0261(.A(new_n646), .B(new_n623), .Y(new_n647));
  nand_5     g0262(.A(new_n647), .B(new_n616), .Y(new_n648));
  nand_5 g0263(.A(pi221), .B(pi221), .Y(new_n649));
  nand_5 g0264(.A(pi062), .B(pi062), .Y(new_n650));
  nand_5 g0265(.A(pi071), .B(pi071), .Y(new_n651));
  nand_5 g0266(.A(pi172), .B(pi172), .Y(new_n652));
  nand_5     g0267(.A(pi181), .B(new_n652), .Y(new_n653));
  nand_5     g0268(.A(new_n653), .B(new_n651), .Y(new_n654));
  nand_5     g0269(.A(new_n654), .B(new_n650), .Y(new_n655));
  nand_5     g0270(.A(new_n655), .B(new_n649), .Y(new_n656));
  nand_5     g0271(.A(new_n652), .B(new_n650), .Y(new_n657));
  nor_5      g0272(.A(new_n657), .B(pi247), .Y(new_n658));
  nand_5 g0273(.A(pi196), .B(pi196), .Y(new_n659));
  nand_5     g0274(.A(new_n659), .B(pi078), .Y(new_n660));
  nand_5 g0275(.A(pi201), .B(pi201), .Y(new_n661));
  nand_5     g0276(.A(new_n661), .B(new_n659), .Y(new_n662));
  nand_5     g0277(.A(new_n662), .B(new_n660), .Y(new_n663));
  nand_5 g0278(.A(new_n663), .B(new_n663), .Y(new_n664));
  nand_5     g0279(.A(new_n664), .B(new_n658), .Y(new_n665));
  nor_5      g0280(.A(pi185), .B(pi108), .Y(new_n666));
  nand_5 g0281(.A(pi187), .B(pi187), .Y(new_n667));
  nand_5     g0282(.A(new_n667), .B(new_n585), .Y(new_n668));
  nor_5      g0283(.A(new_n668), .B(new_n591), .Y(new_n669));
  nand_5     g0284(.A(new_n669), .B(new_n666), .Y(new_n670));
  nor_5      g0285(.A(new_n670), .B(pi136), .Y(new_n671));
  nand_5     g0286(.A(new_n671), .B(new_n665), .Y(new_n672));
  nor_5      g0287(.A(new_n672), .B(new_n656), .Y(new_n673));
  nand_5 g0288(.A(new_n607), .B(new_n607), .Y(new_n674));
  nand_5     g0289(.A(new_n658), .B(new_n674), .Y(new_n675));
  nand_5 g0290(.A(new_n675), .B(new_n675), .Y(new_n676));
  nand_5     g0291(.A(new_n676), .B(new_n604), .Y(new_n677));
  nand_5 g0292(.A(new_n677), .B(new_n677), .Y(new_n678));
  nand_5 g0293(.A(pi039), .B(pi039), .Y(new_n679));
  nor_5      g0294(.A(pi195), .B(pi078), .Y(new_n680));
  nand_5     g0295(.A(new_n680), .B(new_n679), .Y(new_n681));
  nand_5     g0296(.A(new_n680), .B(pi104), .Y(new_n682));
  nand_5     g0297(.A(new_n682), .B(new_n681), .Y(new_n683));
  nand_5     g0298(.A(new_n683), .B(new_n678), .Y(new_n684));
  nand_5 g0299(.A(new_n684), .B(new_n684), .Y(new_n685));
  nor_5      g0300(.A(new_n685), .B(new_n583), .Y(new_n686));
  nand_5     g0301(.A(new_n686), .B(new_n673), .Y(new_n687));
  nand_5 g0302(.A(pi013), .B(pi013), .Y(new_n688));
  nand_5 g0303(.A(pi168), .B(pi168), .Y(new_n689));
  nand_5     g0304(.A(new_n689), .B(new_n688), .Y(new_n690));
  nor_5      g0305(.A(new_n690), .B(pi070), .Y(new_n691));
  nand_5 g0306(.A(pi051), .B(pi051), .Y(new_n692));
  nand_5     g0307(.A(pi074), .B(new_n688), .Y(new_n693));
  nand_5     g0308(.A(new_n693), .B(new_n692), .Y(new_n694));
  nand_5     g0309(.A(new_n694), .B(new_n689), .Y(new_n695));
  nor_5      g0310(.A(pi179), .B(pi114), .Y(new_n696));
  nand_5     g0311(.A(new_n696), .B(new_n695), .Y(new_n697));
  nor_5      g0312(.A(new_n697), .B(new_n691), .Y(new_n698));
  nand_5 g0313(.A(new_n698), .B(new_n698), .Y(new_n699));
  nand_5 g0314(.A(pi147), .B(pi147), .Y(new_n700));
  nand_5     g0315(.A(new_n700), .B(pi009), .Y(new_n701));
  nor_5      g0316(.A(pi074), .B(pi051), .Y(new_n702));
  nor_5      g0317(.A(pi240), .B(pi179), .Y(new_n703));
  nand_5     g0318(.A(new_n703), .B(new_n702), .Y(new_n704));
  nor_5      g0319(.A(new_n704), .B(pi114), .Y(new_n705));
  nand_5     g0320(.A(new_n705), .B(new_n701), .Y(new_n706));
  nand_5     g0321(.A(new_n706), .B(new_n699), .Y(new_n707));
  nand_5     g0322(.A(new_n707), .B(new_n687), .Y(new_n708));
  nor_5      g0323(.A(new_n708), .B(new_n648), .Y(new_n709));
  nand_5 g0324(.A(pi154), .B(pi154), .Y(new_n710));
  nand_5     g0325(.A(new_n710), .B(pi055), .Y(new_n711));
  nand_5 g0326(.A(new_n711), .B(new_n711), .Y(new_n712));
  nand_5 g0327(.A(pi035), .B(pi035), .Y(new_n713));
  nand_5 g0328(.A(pi132), .B(pi132), .Y(new_n714));
  nand_5     g0329(.A(new_n714), .B(new_n713), .Y(new_n715));
  nor_5      g0330(.A(new_n715), .B(new_n712), .Y(new_n716));
  nand_5 g0331(.A(pi243), .B(pi243), .Y(new_n717));
  nor_5      g0332(.A(pi145), .B(pi083), .Y(new_n718));
  nand_5     g0333(.A(new_n718), .B(new_n717), .Y(new_n719));
  nand_5 g0334(.A(pi059), .B(pi059), .Y(new_n720));
  nand_5 g0335(.A(pi208), .B(pi208), .Y(new_n721));
  nand_5     g0336(.A(new_n721), .B(new_n720), .Y(new_n722));
  nor_5      g0337(.A(new_n722), .B(new_n719), .Y(new_n723));
  nand_5 g0338(.A(pi001), .B(pi001), .Y(new_n724));
  nand_5 g0339(.A(pi151), .B(pi151), .Y(new_n725));
  nand_5     g0340(.A(new_n725), .B(new_n724), .Y(new_n726));
  nand_5 g0341(.A(pi061), .B(pi061), .Y(new_n727));
  nand_5 g0342(.A(pi173), .B(pi173), .Y(new_n728));
  nand_5     g0343(.A(new_n728), .B(new_n727), .Y(new_n729));
  nor_5      g0344(.A(new_n729), .B(new_n726), .Y(new_n730));
  nand_5     g0345(.A(new_n730), .B(new_n723), .Y(new_n731));
  nand_5 g0346(.A(new_n731), .B(new_n731), .Y(new_n732));
  nand_5     g0347(.A(new_n732), .B(new_n716), .Y(new_n733));
  nand_5 g0348(.A(pi086), .B(pi086), .Y(new_n734));
  nand_5 g0349(.A(pi148), .B(pi148), .Y(new_n735));
  nand_5 g0350(.A(pi188), .B(pi188), .Y(new_n736));
  nand_5     g0351(.A(new_n736), .B(pi084), .Y(new_n737));
  nand_5 g0352(.A(new_n737), .B(new_n737), .Y(new_n738));
  nand_5 g0353(.A(pi048), .B(pi048), .Y(new_n739));
  nand_5 g0354(.A(pi052), .B(pi052), .Y(new_n740));
  nand_5     g0355(.A(new_n740), .B(new_n739), .Y(new_n741));
  nor_5      g0356(.A(new_n741), .B(new_n738), .Y(new_n742));
  nand_5 g0357(.A(pi015), .B(pi015), .Y(new_n743));
  nand_5     g0358(.A(pi235), .B(new_n740), .Y(new_n744));
  nand_5     g0359(.A(new_n744), .B(new_n743), .Y(new_n745));
  nor_5      g0360(.A(new_n745), .B(new_n742), .Y(new_n746));
  nand_5 g0361(.A(new_n746), .B(new_n746), .Y(new_n747));
  nand_5     g0362(.A(new_n747), .B(new_n735), .Y(new_n748));
  nand_5     g0363(.A(new_n748), .B(new_n734), .Y(new_n749));
  nand_5 g0364(.A(pi091), .B(pi091), .Y(new_n750));
  nand_5 g0365(.A(pi142), .B(pi142), .Y(new_n751));
  nand_5     g0366(.A(new_n751), .B(new_n750), .Y(new_n752));
  nand_5 g0367(.A(new_n752), .B(new_n752), .Y(new_n753));
  nand_5     g0368(.A(new_n753), .B(new_n749), .Y(new_n754));
  nand_5 g0369(.A(pi216), .B(pi216), .Y(new_n755));
  nand_5 g0370(.A(pi045), .B(pi045), .Y(new_n756));
  nand_5 g0371(.A(pi058), .B(pi058), .Y(new_n757));
  nand_5     g0372(.A(new_n757), .B(new_n756), .Y(new_n758));
  nand_5 g0373(.A(new_n758), .B(new_n758), .Y(new_n759));
  nand_5     g0374(.A(new_n759), .B(new_n755), .Y(new_n760));
  nand_5 g0375(.A(new_n760), .B(new_n760), .Y(new_n761));
  nand_5     g0376(.A(pi064), .B(new_n757), .Y(new_n762));
  nand_5     g0377(.A(new_n762), .B(new_n758), .Y(new_n763));
  nor_5      g0378(.A(pi191), .B(pi064), .Y(new_n764));
  nand_5 g0379(.A(new_n764), .B(new_n764), .Y(new_n765));
  nand_5     g0380(.A(new_n765), .B(new_n763), .Y(new_n766));
  nand_5 g0381(.A(pi046), .B(pi046), .Y(new_n767));
  nand_5 g0382(.A(pi112), .B(pi112), .Y(new_n768));
  nand_5     g0383(.A(new_n768), .B(new_n767), .Y(new_n769));
  nand_5 g0384(.A(new_n769), .B(new_n769), .Y(new_n770));
  nand_5     g0385(.A(new_n770), .B(new_n766), .Y(new_n771));
  nor_5      g0386(.A(new_n771), .B(new_n761), .Y(new_n772));
  nand_5 g0387(.A(pi222), .B(pi222), .Y(new_n773));
  nand_5     g0388(.A(new_n764), .B(new_n773), .Y(new_n774));
  nand_5 g0389(.A(pi004), .B(pi004), .Y(new_n775));
  nand_5     g0390(.A(pi150), .B(new_n775), .Y(new_n776));
  nand_5     g0391(.A(new_n776), .B(new_n770), .Y(new_n777));
  nor_5      g0392(.A(new_n777), .B(new_n774), .Y(new_n778));
  nor_5      g0393(.A(new_n778), .B(new_n772), .Y(new_n779));
  nand_5 g0394(.A(new_n779), .B(new_n779), .Y(new_n780));
  nand_5 g0395(.A(pi133), .B(pi133), .Y(new_n781));
  nand_5 g0396(.A(pi175), .B(pi175), .Y(new_n782));
  nand_5     g0397(.A(new_n782), .B(new_n781), .Y(new_n783));
  nand_5 g0398(.A(new_n783), .B(new_n783), .Y(new_n784));
  nand_5 g0399(.A(pi053), .B(pi053), .Y(new_n785));
  nand_5     g0400(.A(pi184), .B(new_n785), .Y(new_n786));
  nand_5     g0401(.A(new_n786), .B(new_n784), .Y(new_n787));
  nand_5 g0402(.A(pi110), .B(pi110), .Y(new_n788));
  nand_5 g0403(.A(pi093), .B(pi093), .Y(new_n789));
  nand_5     g0404(.A(pi244), .B(new_n789), .Y(new_n790));
  nand_5     g0405(.A(new_n790), .B(new_n788), .Y(new_n791));
  nor_5      g0406(.A(new_n791), .B(pi053), .Y(new_n792));
  nor_5      g0407(.A(new_n792), .B(new_n787), .Y(new_n793));
  nand_5 g0408(.A(pi008), .B(pi008), .Y(new_n794));
  nand_5 g0409(.A(pi229), .B(pi229), .Y(new_n795));
  nand_5     g0410(.A(new_n781), .B(pi124), .Y(new_n796));
  nand_5     g0411(.A(new_n796), .B(new_n795), .Y(new_n797));
  nand_5 g0412(.A(new_n797), .B(new_n797), .Y(new_n798));
  nand_5     g0413(.A(new_n798), .B(new_n794), .Y(new_n799));
  nor_5      g0414(.A(new_n799), .B(new_n793), .Y(new_n800));
  nand_5     g0415(.A(new_n800), .B(new_n780), .Y(new_n801));
  nor_5      g0416(.A(new_n801), .B(new_n754), .Y(new_n802));
  nor_5      g0417(.A(pi209), .B(pi160), .Y(new_n803));
  nand_5 g0418(.A(new_n803), .B(new_n803), .Y(new_n804));
  nand_5 g0419(.A(pi160), .B(pi160), .Y(new_n805));
  nand_5     g0420(.A(new_n805), .B(pi008), .Y(new_n806));
  nand_5     g0421(.A(new_n806), .B(new_n804), .Y(new_n807));
  nand_5     g0422(.A(new_n807), .B(new_n775), .Y(new_n808));
  nand_5 g0423(.A(new_n808), .B(new_n808), .Y(new_n809));
  nand_5     g0424(.A(new_n809), .B(new_n761), .Y(new_n810));
  nand_5     g0425(.A(new_n810), .B(new_n780), .Y(new_n811));
  nand_5     g0426(.A(new_n811), .B(new_n801), .Y(new_n812));
  nor_5      g0427(.A(new_n810), .B(new_n787), .Y(new_n813));
  nor_5      g0428(.A(pi093), .B(pi031), .Y(new_n814));
  nand_5     g0429(.A(pi249), .B(new_n750), .Y(new_n815));
  nand_5     g0430(.A(new_n815), .B(new_n814), .Y(new_n816));
  nand_5 g0431(.A(new_n816), .B(new_n816), .Y(new_n817));
  nand_5     g0432(.A(new_n817), .B(new_n813), .Y(new_n818));
  nand_5     g0433(.A(new_n818), .B(new_n812), .Y(new_n819));
  nand_5 g0434(.A(new_n819), .B(new_n819), .Y(new_n820));
  nor_5      g0435(.A(new_n820), .B(new_n802), .Y(new_n821));
  nor_5      g0436(.A(new_n821), .B(new_n733), .Y(new_n822));
  nand_5 g0437(.A(new_n681), .B(new_n681), .Y(new_n823));
  nand_5 g0438(.A(new_n733), .B(new_n733), .Y(new_n824));
  nor_5      g0439(.A(pi203), .B(pi135), .Y(new_n825));
  nand_5 g0440(.A(new_n825), .B(new_n825), .Y(new_n826));
  nor_5      g0441(.A(pi177), .B(pi087), .Y(new_n827));
  nand_5 g0442(.A(pi177), .B(pi177), .Y(new_n828));
  nand_5     g0443(.A(new_n828), .B(pi059), .Y(new_n829));
  nand_5     g0444(.A(new_n829), .B(new_n721), .Y(new_n830));
  nor_5      g0445(.A(new_n830), .B(new_n827), .Y(new_n831));
  nor_5      g0446(.A(new_n831), .B(new_n826), .Y(new_n832));
  nor_5      g0447(.A(pi203), .B(new_n727), .Y(new_n833));
  nand_5 g0448(.A(new_n833), .B(new_n833), .Y(new_n834));
  nand_5     g0449(.A(new_n834), .B(new_n728), .Y(new_n835));
  nor_5      g0450(.A(new_n835), .B(new_n832), .Y(new_n836));
  nand_5 g0451(.A(pi211), .B(pi211), .Y(new_n837));
  nand_5 g0452(.A(pi225), .B(pi225), .Y(new_n838));
  nand_5     g0453(.A(new_n838), .B(new_n837), .Y(new_n839));
  nor_5      g0454(.A(new_n839), .B(new_n836), .Y(new_n840));
  nor_5      g0455(.A(pi040), .B(pi024), .Y(new_n841));
  nand_5     g0456(.A(new_n841), .B(new_n827), .Y(new_n842));
  nand_5 g0457(.A(pi024), .B(pi024), .Y(new_n843));
  nand_5     g0458(.A(pi145), .B(new_n843), .Y(new_n844));
  nand_5     g0459(.A(new_n844), .B(new_n717), .Y(new_n845));
  nand_5     g0460(.A(new_n845), .B(new_n827), .Y(new_n846));
  nand_5     g0461(.A(new_n846), .B(new_n842), .Y(new_n847));
  nand_5     g0462(.A(new_n847), .B(new_n719), .Y(new_n848));
  nor_5      g0463(.A(new_n830), .B(pi061), .Y(new_n849));
  nand_5     g0464(.A(new_n849), .B(new_n848), .Y(new_n850));
  nand_5 g0465(.A(new_n850), .B(new_n850), .Y(new_n851));
  nand_5     g0466(.A(new_n851), .B(new_n728), .Y(new_n852));
  nand_5 g0467(.A(new_n852), .B(new_n852), .Y(new_n853));
  nand_5 g0468(.A(pi014), .B(pi014), .Y(new_n854));
  nand_5     g0469(.A(new_n854), .B(pi001), .Y(new_n855));
  nor_5      g0470(.A(pi140), .B(pi014), .Y(new_n856));
  nand_5 g0471(.A(pi134), .B(pi134), .Y(new_n857));
  nand_5     g0472(.A(pi250), .B(new_n714), .Y(new_n858));
  nand_5     g0473(.A(new_n858), .B(new_n857), .Y(new_n859));
  nand_5     g0474(.A(new_n859), .B(new_n725), .Y(new_n860));
  nand_5     g0475(.A(new_n860), .B(new_n856), .Y(new_n861));
  nand_5     g0476(.A(new_n861), .B(new_n855), .Y(new_n862));
  nand_5     g0477(.A(new_n862), .B(new_n841), .Y(new_n863));
  nand_5     g0478(.A(new_n863), .B(new_n853), .Y(new_n864));
  nand_5     g0479(.A(new_n864), .B(new_n840), .Y(new_n865));
  nor_5      g0480(.A(new_n865), .B(new_n824), .Y(new_n866));
  nand_5     g0481(.A(new_n866), .B(new_n823), .Y(new_n867));
  nor_5      g0482(.A(new_n839), .B(new_n681), .Y(new_n868));
  nand_5 g0483(.A(pi197), .B(pi197), .Y(new_n869));
  nand_5     g0484(.A(new_n768), .B(pi006), .Y(new_n870));
  nand_5     g0485(.A(new_n870), .B(new_n869), .Y(new_n871));
  nand_5 g0486(.A(new_n871), .B(new_n871), .Y(new_n872));
  nand_5     g0487(.A(new_n872), .B(new_n710), .Y(new_n873));
  nand_5 g0488(.A(new_n873), .B(new_n873), .Y(new_n874));
  nand_5 g0489(.A(new_n842), .B(new_n842), .Y(new_n875));
  nand_5     g0490(.A(new_n856), .B(new_n875), .Y(new_n876));
  nand_5 g0491(.A(pi250), .B(pi250), .Y(new_n877));
  nand_5     g0492(.A(new_n877), .B(new_n857), .Y(new_n878));
  nand_5 g0493(.A(new_n878), .B(new_n878), .Y(new_n879));
  nand_5     g0494(.A(new_n879), .B(new_n825), .Y(new_n880));
  nor_5      g0495(.A(new_n880), .B(new_n876), .Y(new_n881));
  nand_5     g0496(.A(new_n881), .B(new_n874), .Y(new_n882));
  nand_5 g0497(.A(new_n882), .B(new_n882), .Y(new_n883));
  nand_5     g0498(.A(new_n883), .B(new_n868), .Y(new_n884));
  nand_5     g0499(.A(new_n884), .B(new_n867), .Y(new_n885));
  nand_5     g0500(.A(new_n676), .B(new_n600), .Y(new_n886));
  nand_5 g0501(.A(new_n886), .B(new_n886), .Y(new_n887));
  nand_5     g0502(.A(new_n887), .B(new_n885), .Y(new_n888));
  nor_5      g0503(.A(new_n888), .B(new_n822), .Y(new_n889));
  nand_5     g0504(.A(new_n656), .B(new_n674), .Y(new_n890));
  nand_5     g0505(.A(new_n890), .B(new_n611), .Y(new_n891));
  nand_5 g0506(.A(new_n891), .B(new_n891), .Y(new_n892));
  nand_5     g0507(.A(new_n892), .B(new_n675), .Y(new_n893));
  nand_5     g0508(.A(new_n893), .B(new_n600), .Y(new_n894));
  nand_5     g0509(.A(new_n894), .B(new_n590), .Y(new_n895));
  nand_5     g0510(.A(new_n682), .B(new_n663), .Y(new_n896));
  nand_5 g0511(.A(new_n896), .B(new_n896), .Y(new_n897));
  nand_5 g0512(.A(pi054), .B(pi054), .Y(new_n898));
  nand_5     g0513(.A(pi211), .B(new_n898), .Y(new_n899));
  nand_5     g0514(.A(new_n899), .B(new_n823), .Y(new_n900));
  nand_5     g0515(.A(new_n900), .B(new_n897), .Y(new_n901));
  nand_5 g0516(.A(new_n662), .B(new_n662), .Y(new_n902));
  nand_5 g0517(.A(pi104), .B(pi104), .Y(new_n903));
  nand_5 g0518(.A(pi158), .B(pi158), .Y(new_n904));
  nand_5     g0519(.A(new_n904), .B(new_n898), .Y(new_n905));
  nand_5 g0520(.A(new_n905), .B(new_n905), .Y(new_n906));
  nand_5     g0521(.A(new_n906), .B(new_n903), .Y(new_n907));
  nand_5 g0522(.A(new_n907), .B(new_n907), .Y(new_n908));
  nand_5     g0523(.A(new_n908), .B(new_n902), .Y(new_n909));
  nand_5     g0524(.A(new_n909), .B(new_n901), .Y(new_n910));
  nand_5     g0525(.A(new_n674), .B(pi221), .Y(new_n911));
  nand_5     g0526(.A(new_n911), .B(new_n611), .Y(new_n912));
  nand_5 g0527(.A(pi181), .B(pi181), .Y(new_n913));
  nand_5     g0528(.A(new_n913), .B(new_n651), .Y(new_n914));
  nand_5 g0529(.A(new_n914), .B(new_n914), .Y(new_n915));
  nand_5     g0530(.A(new_n915), .B(new_n590), .Y(new_n916));
  nor_5      g0531(.A(new_n916), .B(new_n912), .Y(new_n917));
  nand_5     g0532(.A(new_n917), .B(new_n910), .Y(new_n918));
  nand_5     g0533(.A(new_n918), .B(new_n895), .Y(new_n919));
  nand_5 g0534(.A(new_n919), .B(new_n919), .Y(new_n920));
  nor_5      g0535(.A(new_n920), .B(new_n889), .Y(new_n921));
  nand_5 g0536(.A(new_n787), .B(new_n787), .Y(new_n922));
  nor_5      g0537(.A(pi249), .B(new_n751), .Y(new_n923));
  nor_5      g0538(.A(new_n923), .B(pi091), .Y(new_n924));
  nor_5      g0539(.A(pi249), .B(pi086), .Y(new_n925));
  nand_5     g0540(.A(new_n925), .B(pi148), .Y(new_n926));
  nand_5     g0541(.A(new_n926), .B(new_n924), .Y(new_n927));
  nand_5     g0542(.A(new_n927), .B(new_n814), .Y(new_n928));
  nand_5     g0543(.A(new_n925), .B(new_n743), .Y(new_n929));
  nand_5     g0544(.A(new_n814), .B(new_n744), .Y(new_n930));
  nor_5      g0545(.A(new_n930), .B(new_n929), .Y(new_n931));
  nand_5 g0546(.A(new_n931), .B(new_n931), .Y(new_n932));
  nand_5     g0547(.A(new_n932), .B(new_n928), .Y(new_n933));
  nand_5     g0548(.A(new_n933), .B(new_n922), .Y(new_n934));
  nand_5     g0549(.A(new_n934), .B(new_n800), .Y(new_n935));
  nand_5     g0550(.A(new_n935), .B(new_n809), .Y(new_n936));
  nand_5 g0551(.A(new_n936), .B(new_n936), .Y(new_n937));
  nand_5 g0552(.A(new_n840), .B(new_n840), .Y(new_n938));
  nand_5 g0553(.A(new_n772), .B(new_n772), .Y(new_n939));
  nand_5     g0554(.A(new_n883), .B(new_n939), .Y(new_n940));
  nor_5      g0555(.A(new_n940), .B(new_n938), .Y(new_n941));
  nand_5     g0556(.A(new_n941), .B(new_n937), .Y(new_n942));
  nand_5 g0557(.A(pi193), .B(pi193), .Y(new_n943));
  nor_5      g0558(.A(pi162), .B(pi096), .Y(new_n944));
  nand_5 g0559(.A(pi002), .B(pi002), .Y(new_n945));
  nand_5 g0560(.A(pi095), .B(pi095), .Y(new_n946));
  nand_5     g0561(.A(new_n946), .B(pi034), .Y(new_n947));
  nand_5     g0562(.A(new_n947), .B(new_n945), .Y(new_n948));
  nand_5     g0563(.A(new_n948), .B(new_n944), .Y(new_n949));
  nand_5 g0564(.A(pi044), .B(pi044), .Y(new_n950));
  nor_5      g0565(.A(pi162), .B(new_n950), .Y(new_n951));
  nor_5      g0566(.A(new_n951), .B(pi205), .Y(new_n952));
  nand_5     g0567(.A(new_n952), .B(new_n949), .Y(new_n953));
  nand_5     g0568(.A(new_n953), .B(new_n943), .Y(new_n954));
  nor_5      g0569(.A(pi116), .B(pi084), .Y(new_n955));
  nand_5     g0570(.A(new_n955), .B(new_n954), .Y(new_n956));
  nand_5 g0571(.A(pi245), .B(pi245), .Y(new_n957));
  nand_5     g0572(.A(new_n957), .B(pi023), .Y(new_n958));
  nor_5      g0573(.A(pi101), .B(pi095), .Y(new_n959));
  nand_5     g0574(.A(new_n959), .B(new_n958), .Y(new_n960));
  nand_5     g0575(.A(new_n944), .B(new_n943), .Y(new_n961));
  nor_5      g0576(.A(new_n961), .B(new_n960), .Y(new_n962));
  nor_5      g0577(.A(new_n962), .B(new_n956), .Y(new_n963));
  nand_5 g0578(.A(pi130), .B(pi130), .Y(new_n964));
  nor_5      g0579(.A(new_n964), .B(pi084), .Y(new_n965));
  nand_5 g0580(.A(pi235), .B(pi235), .Y(new_n966));
  nand_5     g0581(.A(new_n966), .B(new_n736), .Y(new_n967));
  nor_5      g0582(.A(new_n967), .B(new_n965), .Y(new_n968));
  nand_5 g0583(.A(new_n968), .B(new_n968), .Y(new_n969));
  nor_5      g0584(.A(new_n969), .B(new_n963), .Y(new_n970));
  nand_5 g0585(.A(new_n970), .B(new_n970), .Y(new_n971));
  nor_5      g0586(.A(new_n971), .B(new_n942), .Y(new_n972));
  nand_5     g0587(.A(new_n584), .B(new_n637), .Y(new_n973));
  nand_5 g0588(.A(new_n973), .B(new_n973), .Y(new_n974));
  nand_5     g0589(.A(new_n974), .B(new_n589), .Y(new_n975));
  nor_5      g0590(.A(new_n975), .B(new_n972), .Y(new_n976));
  nand_5     g0591(.A(new_n976), .B(new_n921), .Y(new_n977));
  nand_5     g0592(.A(new_n977), .B(new_n709), .Y(new_n978));
  nand_5 g0593(.A(new_n623), .B(new_n623), .Y(new_n979));
  nand_5 g0594(.A(pi174), .B(pi174), .Y(new_n980));
  nand_5 g0595(.A(pi068), .B(pi068), .Y(new_n981));
  nand_5     g0596(.A(pi180), .B(new_n981), .Y(new_n982));
  nand_5     g0597(.A(new_n982), .B(new_n980), .Y(new_n983));
  nand_5     g0598(.A(new_n983), .B(new_n625), .Y(new_n984));
  nand_5 g0599(.A(pi005), .B(pi005), .Y(new_n985));
  nor_5      g0600(.A(pi167), .B(new_n985), .Y(new_n986));
  nor_5      g0601(.A(new_n986), .B(pi107), .Y(new_n987));
  nand_5     g0602(.A(new_n987), .B(new_n984), .Y(new_n988));
  nand_5 g0603(.A(new_n988), .B(new_n988), .Y(new_n989));
  nand_5     g0604(.A(new_n628), .B(pi063), .Y(new_n990));
  nand_5     g0605(.A(new_n990), .B(new_n989), .Y(new_n991));
  nor_5      g0606(.A(new_n991), .B(pi118), .Y(new_n992));
  nand_5 g0607(.A(new_n992), .B(new_n992), .Y(new_n993));
  nand_5     g0608(.A(new_n993), .B(new_n979), .Y(new_n994));
  nand_5     g0609(.A(new_n617), .B(pi019), .Y(new_n995));
  nand_5 g0610(.A(pi037), .B(pi037), .Y(new_n996));
  nand_5     g0611(.A(new_n700), .B(new_n996), .Y(new_n997));
  nand_5 g0612(.A(new_n997), .B(new_n997), .Y(new_n998));
  nand_5     g0613(.A(new_n998), .B(new_n995), .Y(new_n999));
  nand_5 g0614(.A(new_n999), .B(new_n999), .Y(new_n1000));
  nand_5     g0615(.A(new_n1000), .B(new_n691), .Y(new_n1001));
  nand_5 g0616(.A(new_n1001), .B(new_n1001), .Y(new_n1002));
  nand_5     g0617(.A(new_n1002), .B(new_n994), .Y(new_n1003));
  nand_5     g0618(.A(new_n1003), .B(new_n707), .Y(new_n1004));
  nand_5 g0619(.A(pi043), .B(pi043), .Y(new_n1005));
  nand_5 g0620(.A(pi198), .B(pi198), .Y(new_n1006));
  nand_5     g0621(.A(new_n1006), .B(new_n513), .Y(new_n1007));
  nand_5 g0622(.A(new_n1007), .B(new_n1007), .Y(new_n1008));
  nand_5     g0623(.A(new_n1008), .B(new_n1005), .Y(new_n1009));
  nand_5 g0624(.A(new_n505), .B(new_n505), .Y(new_n1010));
  nor_5      g0625(.A(pi199), .B(pi066), .Y(new_n1011));
  nand_5     g0626(.A(new_n1011), .B(new_n1010), .Y(new_n1012));
  nor_5      g0627(.A(new_n1012), .B(new_n1009), .Y(new_n1013));
  nand_5 g0628(.A(new_n1013), .B(new_n1013), .Y(new_n1014));
  nand_5 g0629(.A(pi114), .B(pi114), .Y(new_n1015));
  nand_5     g0630(.A(new_n1015), .B(pi106), .Y(new_n1016));
  nand_5     g0631(.A(new_n1016), .B(new_n522), .Y(new_n1017));
  nor_5      g0632(.A(new_n1017), .B(new_n1014), .Y(new_n1018));
  and_6      g0633(.A(new_n1018), .B(new_n492), .Y(new_n1019));
  nand_5     g0634(.A(new_n1019), .B(new_n1004), .Y(new_n1020));
  nand_5 g0635(.A(new_n1020), .B(new_n1020), .Y(new_n1021));
  nand_5     g0636(.A(new_n1021), .B(new_n978), .Y(new_n1022));
  nand_5     g0637(.A(new_n1022), .B(new_n577), .Y(new_n1023));
  nand_5     g0638(.A(new_n1023), .B(new_n481), .Y(new_n1024));
  nand_5     g0639(.A(new_n1024), .B(new_n426), .Y(new_n1025));
  nand_5 g0640(.A(new_n1025), .B(new_n1025), .Y(new_n1026));
  nand_5 g0641(.A(pi184), .B(pi184), .Y(new_n1027));
  nand_5     g0642(.A(new_n814), .B(new_n1027), .Y(new_n1028));
  nand_5     g0643(.A(new_n925), .B(new_n782), .Y(new_n1029));
  nor_5      g0644(.A(new_n1029), .B(new_n1028), .Y(new_n1030));
  nand_5     g0645(.A(new_n959), .B(new_n944), .Y(new_n1031));
  nand_5 g0646(.A(new_n1031), .B(new_n1031), .Y(new_n1032));
  nor_5      g0647(.A(new_n1032), .B(new_n953), .Y(new_n1033));
  nand_5 g0648(.A(pi034), .B(pi034), .Y(new_n1034));
  nand_5     g0649(.A(new_n1034), .B(new_n945), .Y(new_n1035));
  nor_5      g0650(.A(pi205), .B(pi044), .Y(new_n1036));
  nand_5     g0651(.A(new_n1036), .B(new_n957), .Y(new_n1037));
  nor_5      g0652(.A(new_n1037), .B(new_n1035), .Y(new_n1038));
  nor_5      g0653(.A(new_n1038), .B(new_n1033), .Y(new_n1039));
  nor_5      g0654(.A(new_n1039), .B(pi116), .Y(new_n1040));
  nor_5      g0655(.A(pi170), .B(pi085), .Y(new_n1041));
  nand_5 g0656(.A(pi233), .B(pi233), .Y(new_n1042));
  nand_5     g0657(.A(new_n1042), .B(pi119), .Y(new_n1043));
  nor_5      g0658(.A(pi233), .B(pi157), .Y(new_n1044));
  nor_5      g0659(.A(new_n1044), .B(pi202), .Y(new_n1045));
  nand_5     g0660(.A(new_n1045), .B(new_n1043), .Y(new_n1046));
  nand_5     g0661(.A(new_n1046), .B(new_n1041), .Y(new_n1047));
  nand_5 g0662(.A(pi137), .B(pi137), .Y(new_n1048));
  nor_5      g0663(.A(pi170), .B(new_n1048), .Y(new_n1049));
  nor_5      g0664(.A(new_n1049), .B(pi023), .Y(new_n1050));
  nand_5     g0665(.A(new_n1050), .B(new_n1047), .Y(new_n1051));
  nand_5 g0666(.A(pi119), .B(pi119), .Y(new_n1052));
  nand_5 g0667(.A(pi234), .B(pi234), .Y(new_n1053));
  nand_5     g0668(.A(new_n1053), .B(new_n1052), .Y(new_n1054));
  nand_5 g0669(.A(pi023), .B(pi023), .Y(new_n1055));
  nor_5      g0670(.A(pi202), .B(pi137), .Y(new_n1056));
  nand_5     g0671(.A(new_n1056), .B(new_n1055), .Y(new_n1057));
  nor_5      g0672(.A(new_n1057), .B(new_n1054), .Y(new_n1058));
  nor_5      g0673(.A(new_n1058), .B(pi245), .Y(new_n1059));
  nand_5     g0674(.A(new_n1059), .B(new_n1051), .Y(new_n1060));
  nand_5     g0675(.A(new_n1060), .B(new_n1032), .Y(new_n1061));
  nand_5     g0676(.A(new_n1061), .B(new_n1040), .Y(new_n1062));
  nand_5 g0677(.A(new_n1062), .B(new_n1062), .Y(new_n1063));
  nand_5 g0678(.A(new_n1047), .B(new_n1047), .Y(new_n1064));
  nor_5      g0679(.A(pi231), .B(pi000), .Y(new_n1065));
  nand_5 g0680(.A(new_n1065), .B(new_n1065), .Y(new_n1066));
  nand_5 g0681(.A(pi161), .B(pi161), .Y(new_n1067));
  nor_5      g0682(.A(pi231), .B(new_n1067), .Y(new_n1068));
  nand_5 g0683(.A(new_n1068), .B(new_n1068), .Y(new_n1069));
  nand_5     g0684(.A(new_n1069), .B(new_n1066), .Y(new_n1070));
  nand_5     g0685(.A(new_n1070), .B(new_n1064), .Y(new_n1071));
  nand_5 g0686(.A(new_n1071), .B(new_n1071), .Y(new_n1072));
  nand_5     g0687(.A(new_n1072), .B(new_n1040), .Y(new_n1073));
  nand_5     g0688(.A(new_n943), .B(new_n964), .Y(new_n1074));
  nand_5     g0689(.A(new_n964), .B(pi116), .Y(new_n1075));
  nand_5     g0690(.A(new_n1075), .B(new_n1074), .Y(new_n1076));
  nand_5     g0691(.A(new_n734), .B(new_n743), .Y(new_n1077));
  nor_5      g0692(.A(new_n1077), .B(new_n967), .Y(new_n1078));
  nand_5     g0693(.A(new_n1078), .B(new_n1076), .Y(new_n1079));
  nand_5 g0694(.A(new_n1079), .B(new_n1079), .Y(new_n1080));
  nand_5     g0695(.A(new_n1080), .B(new_n1073), .Y(new_n1081));
  nor_5      g0696(.A(new_n1081), .B(new_n1063), .Y(new_n1082));
  nand_5 g0697(.A(new_n1082), .B(new_n1082), .Y(new_n1083));
  nand_5 g0698(.A(pi073), .B(pi073), .Y(new_n1084));
  nand_5     g0699(.A(new_n1067), .B(new_n1084), .Y(new_n1085));
  nand_5 g0700(.A(new_n1085), .B(new_n1085), .Y(new_n1086));
  nand_5 g0701(.A(pi065), .B(pi065), .Y(new_n1087));
  nand_5     g0702(.A(pi072), .B(new_n1087), .Y(new_n1088));
  nand_5     g0703(.A(new_n1088), .B(new_n1086), .Y(new_n1089));
  nor_5      g0704(.A(new_n1089), .B(new_n1031), .Y(new_n1090));
  nand_5     g0705(.A(new_n1090), .B(new_n1058), .Y(new_n1091));
  nor_5      g0706(.A(new_n1091), .B(new_n1079), .Y(new_n1092));
  nor_5      g0707(.A(new_n1092), .B(new_n746), .Y(new_n1093));
  nand_5     g0708(.A(new_n1093), .B(new_n1083), .Y(new_n1094));
  nand_5     g0709(.A(new_n1094), .B(new_n1030), .Y(new_n1095));
  nor_5      g0710(.A(pi229), .B(pi124), .Y(new_n1096));
  nand_5 g0711(.A(pi031), .B(pi031), .Y(new_n1097));
  nand_5     g0712(.A(new_n789), .B(new_n1097), .Y(new_n1098));
  nor_5      g0713(.A(new_n1098), .B(pi184), .Y(new_n1099));
  nand_5     g0714(.A(new_n929), .B(new_n926), .Y(new_n1100));
  nand_5     g0715(.A(new_n1100), .B(new_n1099), .Y(new_n1101));
  nor_5      g0716(.A(pi148), .B(pi052), .Y(new_n1102));
  nor_5      g0717(.A(new_n1102), .B(new_n1101), .Y(new_n1103));
  nand_5     g0718(.A(new_n791), .B(new_n1027), .Y(new_n1104));
  nand_5 g0719(.A(pi249), .B(pi249), .Y(new_n1105));
  nand_5     g0720(.A(new_n1105), .B(pi142), .Y(new_n1106));
  nand_5     g0721(.A(new_n1106), .B(new_n750), .Y(new_n1107));
  nand_5     g0722(.A(new_n1099), .B(new_n1107), .Y(new_n1108));
  nand_5     g0723(.A(new_n1108), .B(new_n1104), .Y(new_n1109));
  nor_5      g0724(.A(new_n1109), .B(new_n1103), .Y(new_n1110));
  nand_5     g0725(.A(new_n1110), .B(new_n785), .Y(new_n1111));
  nand_5     g0726(.A(new_n1111), .B(new_n782), .Y(new_n1112));
  nand_5     g0727(.A(new_n1112), .B(new_n1096), .Y(new_n1113));
  nand_5 g0728(.A(new_n1113), .B(new_n1113), .Y(new_n1114));
  nand_5     g0729(.A(new_n1114), .B(new_n1095), .Y(new_n1115));
  nand_5     g0730(.A(new_n795), .B(pi133), .Y(new_n1116));
  nand_5 g0731(.A(new_n876), .B(new_n876), .Y(new_n1117));
  nand_5     g0732(.A(pi222), .B(new_n755), .Y(new_n1118));
  nand_5     g0733(.A(new_n755), .B(new_n775), .Y(new_n1119));
  nand_5     g0734(.A(new_n1119), .B(new_n1118), .Y(new_n1120));
  nand_5     g0735(.A(new_n869), .B(new_n710), .Y(new_n1121));
  nand_5 g0736(.A(pi006), .B(pi006), .Y(new_n1122));
  nand_5     g0737(.A(new_n759), .B(new_n1122), .Y(new_n1123));
  nor_5      g0738(.A(new_n1123), .B(new_n1121), .Y(new_n1124));
  nand_5     g0739(.A(new_n1124), .B(new_n1120), .Y(new_n1125));
  nor_5      g0740(.A(new_n1125), .B(new_n878), .Y(new_n1126));
  nand_5     g0741(.A(new_n1126), .B(new_n1117), .Y(new_n1127));
  nand_5 g0742(.A(new_n1127), .B(new_n1127), .Y(new_n1128));
  nand_5     g0743(.A(new_n1128), .B(new_n803), .Y(new_n1129));
  nand_5 g0744(.A(new_n1129), .B(new_n1129), .Y(new_n1130));
  nand_5     g0745(.A(new_n1130), .B(new_n1116), .Y(new_n1131));
  nand_5 g0746(.A(new_n1131), .B(new_n1131), .Y(new_n1132));
  nand_5     g0747(.A(new_n1132), .B(new_n1115), .Y(new_n1133));
  nand_5 g0748(.A(new_n1133), .B(new_n1133), .Y(new_n1134));
  nand_5     g0749(.A(new_n1061), .B(new_n949), .Y(new_n1135));
  nand_5     g0750(.A(new_n1076), .B(new_n736), .Y(new_n1136));
  nand_5 g0751(.A(new_n1136), .B(new_n1136), .Y(new_n1137));
  nand_5     g0752(.A(new_n1137), .B(new_n1135), .Y(new_n1138));
  nand_5 g0753(.A(new_n1138), .B(new_n1138), .Y(new_n1139));
  nand_5 g0754(.A(pi072), .B(pi072), .Y(new_n1140));
  nand_5     g0755(.A(pi080), .B(new_n1140), .Y(new_n1141));
  nand_5     g0756(.A(new_n1141), .B(new_n1087), .Y(new_n1142));
  nand_5     g0757(.A(new_n1142), .B(new_n1086), .Y(new_n1143));
  nand_5     g0758(.A(new_n1143), .B(new_n1070), .Y(new_n1144));
  nand_5     g0759(.A(new_n1086), .B(new_n1140), .Y(new_n1145));
  nand_5 g0760(.A(new_n1145), .B(new_n1145), .Y(new_n1146));
  nand_5 g0761(.A(pi213), .B(pi213), .Y(new_n1147));
  nand_5     g0762(.A(new_n1147), .B(pi027), .Y(new_n1148));
  nand_5 g0763(.A(new_n1148), .B(new_n1148), .Y(new_n1149));
  nand_5     g0764(.A(new_n1149), .B(new_n1146), .Y(new_n1150));
  nand_5     g0765(.A(new_n1041), .B(new_n957), .Y(new_n1151));
  nand_5 g0766(.A(new_n1035), .B(new_n1035), .Y(new_n1152));
  nand_5     g0767(.A(new_n1044), .B(new_n1152), .Y(new_n1153));
  nor_5      g0768(.A(new_n1153), .B(new_n1151), .Y(new_n1154));
  nand_5     g0769(.A(new_n1154), .B(new_n1150), .Y(new_n1155));
  nor_5      g0770(.A(new_n1155), .B(new_n1144), .Y(new_n1156));
  nor_5      g0771(.A(pi213), .B(pi097), .Y(new_n1157));
  nand_5     g0772(.A(new_n1157), .B(pi236), .Y(new_n1158));
  nand_5 g0773(.A(pi036), .B(pi036), .Y(new_n1159));
  nand_5     g0774(.A(new_n1157), .B(new_n1159), .Y(new_n1160));
  nand_5     g0775(.A(new_n1160), .B(new_n1158), .Y(new_n1161));
  nand_5     g0776(.A(new_n1161), .B(new_n1146), .Y(new_n1162));
  nand_5     g0777(.A(new_n1162), .B(new_n1156), .Y(new_n1163));
  nand_5     g0778(.A(new_n1163), .B(new_n1139), .Y(new_n1164));
  nand_5     g0779(.A(new_n1051), .B(new_n1038), .Y(new_n1165));
  nand_5     g0780(.A(new_n955), .B(new_n739), .Y(new_n1166));
  nor_5      g0781(.A(new_n1166), .B(new_n1165), .Y(new_n1167));
  nand_5 g0782(.A(new_n1167), .B(new_n1167), .Y(new_n1168));
  nor_5      g0783(.A(new_n1168), .B(new_n754), .Y(new_n1169));
  nand_5     g0784(.A(new_n1169), .B(new_n1164), .Y(new_n1170));
  nand_5     g0785(.A(new_n1170), .B(new_n1134), .Y(new_n1171));
  nand_5     g0786(.A(new_n874), .B(new_n811), .Y(new_n1172));
  nand_5 g0787(.A(new_n1172), .B(new_n1172), .Y(new_n1173));
  nand_5     g0788(.A(new_n1173), .B(new_n801), .Y(new_n1174));
  nand_5     g0789(.A(new_n975), .B(new_n645), .Y(new_n1175));
  nand_5 g0790(.A(new_n1175), .B(new_n1175), .Y(new_n1176));
  nand_5     g0791(.A(new_n1176), .B(new_n633), .Y(new_n1177));
  nand_5     g0792(.A(new_n1177), .B(new_n992), .Y(new_n1178));
  nand_5     g0793(.A(new_n1018), .B(new_n1002), .Y(new_n1179));
  nor_5      g0794(.A(new_n1179), .B(new_n1178), .Y(new_n1180));
  nand_5 g0795(.A(new_n1180), .B(new_n1180), .Y(new_n1181));
  nand_5 g0796(.A(new_n918), .B(new_n918), .Y(new_n1182));
  nand_5     g0797(.A(new_n1182), .B(new_n824), .Y(new_n1183));
  nor_5      g0798(.A(new_n1183), .B(new_n1181), .Y(new_n1184));
  nand_5     g0799(.A(new_n1184), .B(new_n1174), .Y(new_n1185));
  nand_5 g0800(.A(new_n1185), .B(new_n1185), .Y(new_n1186));
  nand_5     g0801(.A(new_n1186), .B(new_n1171), .Y(new_n1187));
  nand_5 g0802(.A(new_n868), .B(new_n868), .Y(new_n1188));
  nand_5     g0803(.A(new_n1182), .B(new_n1188), .Y(new_n1189));
  nand_5     g0804(.A(new_n893), .B(new_n604), .Y(new_n1190));
  nand_5     g0805(.A(new_n1190), .B(new_n597), .Y(new_n1191));
  nand_5 g0806(.A(new_n1191), .B(new_n1191), .Y(new_n1192));
  nand_5 g0807(.A(new_n641), .B(new_n641), .Y(new_n1193));
  nand_5     g0808(.A(new_n1193), .B(new_n633), .Y(new_n1194));
  nor_5      g0809(.A(new_n1194), .B(new_n1192), .Y(new_n1195));
  nand_5     g0810(.A(new_n1195), .B(new_n1189), .Y(new_n1196));
  nand_5     g0811(.A(new_n1196), .B(new_n1180), .Y(new_n1197));
  nand_5 g0812(.A(new_n1197), .B(new_n1197), .Y(new_n1198));
  nor_5      g0813(.A(new_n847), .B(new_n830), .Y(new_n1199));
  nor_5      g0814(.A(new_n1199), .B(new_n826), .Y(new_n1200));
  nand_5     g0815(.A(new_n855), .B(new_n723), .Y(new_n1201));
  nand_5     g0816(.A(new_n1201), .B(new_n1200), .Y(new_n1202));
  nand_5     g0817(.A(new_n725), .B(pi134), .Y(new_n1203));
  nand_5     g0818(.A(new_n1203), .B(new_n856), .Y(new_n1204));
  nand_5 g0819(.A(new_n1204), .B(new_n1204), .Y(new_n1205));
  nand_5     g0820(.A(new_n1205), .B(new_n1200), .Y(new_n1206));
  nand_5 g0821(.A(new_n1206), .B(new_n1206), .Y(new_n1207));
  nand_5     g0822(.A(new_n877), .B(pi035), .Y(new_n1208));
  nand_5     g0823(.A(new_n725), .B(new_n714), .Y(new_n1209));
  nand_5 g0824(.A(new_n1209), .B(new_n1209), .Y(new_n1210));
  and_6      g0825(.A(new_n1210), .B(new_n1208), .Y(new_n1211));
  nand_5 g0826(.A(new_n1211), .B(new_n1211), .Y(new_n1212));
  nand_5     g0827(.A(new_n1212), .B(new_n1207), .Y(new_n1213));
  nand_5     g0828(.A(new_n1213), .B(new_n1202), .Y(new_n1214));
  nand_5 g0829(.A(new_n835), .B(new_n835), .Y(new_n1215));
  nand_5     g0830(.A(new_n1182), .B(new_n1215), .Y(new_n1216));
  nor_5      g0831(.A(new_n1216), .B(new_n1214), .Y(new_n1217));
  nand_5     g0832(.A(new_n1121), .B(new_n711), .Y(new_n1218));
  nand_5     g0833(.A(new_n1218), .B(new_n877), .Y(new_n1219));
  nand_5 g0834(.A(new_n1219), .B(new_n1219), .Y(new_n1220));
  nand_5     g0835(.A(new_n1220), .B(new_n1207), .Y(new_n1221));
  nand_5     g0836(.A(new_n1221), .B(new_n1180), .Y(new_n1222));
  nand_5 g0837(.A(new_n1222), .B(new_n1222), .Y(new_n1223));
  nand_5     g0838(.A(new_n1223), .B(new_n1217), .Y(new_n1224));
  nor_5      g0839(.A(new_n542), .B(new_n503), .Y(new_n1225));
  nand_5 g0840(.A(new_n706), .B(new_n706), .Y(new_n1226));
  nand_5     g0841(.A(new_n1000), .B(new_n623), .Y(new_n1227));
  nand_5     g0842(.A(new_n1227), .B(new_n1226), .Y(new_n1228));
  nand_5     g0843(.A(new_n1228), .B(new_n699), .Y(new_n1229));
  nand_5     g0844(.A(new_n1229), .B(new_n1225), .Y(new_n1230));
  nor_5      g0845(.A(new_n1018), .B(new_n546), .Y(new_n1231));
  nand_5     g0846(.A(new_n1231), .B(new_n525), .Y(new_n1232));
  nand_5     g0847(.A(new_n1232), .B(new_n1230), .Y(new_n1233));
  nand_5     g0848(.A(new_n1233), .B(new_n1224), .Y(new_n1234));
  nor_5      g0849(.A(new_n1234), .B(new_n1198), .Y(new_n1235));
  nand_5     g0850(.A(new_n1235), .B(new_n1187), .Y(new_n1236));
  nand_5 g0851(.A(new_n1073), .B(new_n1073), .Y(new_n1237));
  nand_5 g0852(.A(new_n1089), .B(new_n1089), .Y(new_n1238));
  nand_5 g0853(.A(pi186), .B(pi186), .Y(new_n1239));
  nand_5     g0854(.A(pi230), .B(new_n1239), .Y(new_n1240));
  nand_5 g0855(.A(new_n1240), .B(new_n1240), .Y(new_n1241));
  nand_5 g0856(.A(pi122), .B(pi122), .Y(new_n1242));
  nand_5 g0857(.A(pi236), .B(pi236), .Y(new_n1243));
  nand_5     g0858(.A(new_n1243), .B(new_n1242), .Y(new_n1244));
  nor_5      g0859(.A(new_n1244), .B(new_n1241), .Y(new_n1245));
  nand_5 g0860(.A(new_n1245), .B(new_n1245), .Y(new_n1246));
  nand_5     g0861(.A(new_n1246), .B(new_n1161), .Y(new_n1247));
  nor_5      g0862(.A(pi080), .B(pi065), .Y(new_n1248));
  nand_5 g0863(.A(new_n1248), .B(new_n1248), .Y(new_n1249));
  nor_5      g0864(.A(new_n1249), .B(new_n1149), .Y(new_n1250));
  nand_5     g0865(.A(new_n1250), .B(new_n1247), .Y(new_n1251));
  nand_5     g0866(.A(new_n1251), .B(new_n1238), .Y(new_n1252));
  nand_5 g0867(.A(new_n1252), .B(new_n1252), .Y(new_n1253));
  nor_5      g0868(.A(new_n1253), .B(new_n754), .Y(new_n1254));
  nand_5     g0869(.A(new_n1254), .B(new_n1237), .Y(new_n1255));
  nor_5      g0870(.A(new_n1255), .B(new_n1185), .Y(new_n1256));
  nand_5     g0871(.A(new_n1144), .B(new_n1053), .Y(new_n1257));
  nand_5     g0872(.A(new_n1257), .B(new_n1044), .Y(new_n1258));
  nand_5 g0873(.A(new_n1258), .B(new_n1258), .Y(new_n1259));
  nand_5 g0874(.A(pi020), .B(pi020), .Y(new_n1260));
  nand_5 g0875(.A(pi028), .B(pi028), .Y(new_n1261));
  nand_5     g0876(.A(new_n1261), .B(new_n1260), .Y(new_n1262));
  nor_5      g0877(.A(new_n1262), .B(pi127), .Y(new_n1263));
  nand_5 g0878(.A(new_n1263), .B(new_n1263), .Y(new_n1264));
  nor_5      g0879(.A(new_n1264), .B(pi206), .Y(new_n1265));
  nand_5 g0880(.A(pi029), .B(pi029), .Y(new_n1266));
  nand_5     g0881(.A(pi099), .B(new_n1266), .Y(new_n1267));
  nand_5     g0882(.A(new_n1267), .B(new_n1265), .Y(new_n1268));
  nand_5 g0883(.A(pi230), .B(pi230), .Y(new_n1269));
  nand_5     g0884(.A(new_n1269), .B(new_n1242), .Y(new_n1270));
  nand_5 g0885(.A(new_n1270), .B(new_n1270), .Y(new_n1271));
  nor_5      g0886(.A(pi236), .B(pi027), .Y(new_n1272));
  nand_5     g0887(.A(new_n1272), .B(new_n1271), .Y(new_n1273));
  nor_5      g0888(.A(new_n1273), .B(new_n1268), .Y(new_n1274));
  nor_5      g0889(.A(pi032), .B(pi029), .Y(new_n1275));
  nand_5 g0890(.A(pi033), .B(pi033), .Y(new_n1276));
  nand_5     g0891(.A(pi131), .B(new_n1276), .Y(new_n1277));
  nand_5     g0892(.A(new_n1277), .B(new_n1275), .Y(new_n1278));
  nand_5     g0893(.A(new_n1278), .B(new_n1274), .Y(new_n1279));
  nand_5     g0894(.A(new_n1158), .B(new_n1148), .Y(new_n1280));
  nand_5     g0895(.A(new_n1280), .B(new_n1140), .Y(new_n1281));
  nand_5 g0896(.A(new_n1281), .B(new_n1281), .Y(new_n1282));
  nand_5     g0897(.A(new_n1263), .B(pi018), .Y(new_n1283));
  nor_5      g0898(.A(new_n1283), .B(new_n1270), .Y(new_n1284));
  nand_5 g0899(.A(pi254), .B(pi254), .Y(new_n1285));
  nand_5 g0900(.A(pi241), .B(pi241), .Y(new_n1286));
  nand_5     g0901(.A(new_n1286), .B(pi127), .Y(new_n1287));
  nor_5      g0902(.A(pi241), .B(pi212), .Y(new_n1288));
  nand_5 g0903(.A(new_n1288), .B(new_n1288), .Y(new_n1289));
  nand_5     g0904(.A(new_n1289), .B(new_n1261), .Y(new_n1290));
  nand_5 g0905(.A(new_n1290), .B(new_n1290), .Y(new_n1291));
  nand_5     g0906(.A(new_n1291), .B(new_n1287), .Y(new_n1292));
  nand_5     g0907(.A(new_n1292), .B(new_n1285), .Y(new_n1293));
  nand_5     g0908(.A(new_n1293), .B(new_n1271), .Y(new_n1294));
  nor_5      g0909(.A(new_n1160), .B(pi072), .Y(new_n1295));
  nand_5 g0910(.A(new_n1295), .B(new_n1295), .Y(new_n1296));
  nor_5      g0911(.A(new_n1239), .B(pi122), .Y(new_n1297));
  nor_5      g0912(.A(new_n1297), .B(new_n1296), .Y(new_n1298));
  nand_5     g0913(.A(new_n1298), .B(new_n1294), .Y(new_n1299));
  nor_5      g0914(.A(new_n1299), .B(new_n1284), .Y(new_n1300));
  nor_5      g0915(.A(new_n1300), .B(new_n1282), .Y(new_n1301));
  nand_5     g0916(.A(new_n1086), .B(new_n1053), .Y(new_n1302));
  nor_5      g0917(.A(new_n1302), .B(new_n1301), .Y(new_n1303));
  nand_5     g0918(.A(new_n1303), .B(new_n1279), .Y(new_n1304));
  nand_5     g0919(.A(new_n1304), .B(new_n1259), .Y(new_n1305));
  nand_5 g0920(.A(new_n1305), .B(new_n1305), .Y(new_n1306));
  nand_5     g0921(.A(new_n1306), .B(new_n1256), .Y(new_n1307));
  nand_5 g0922(.A(new_n1307), .B(new_n1307), .Y(new_n1308));
  nor_5      g0923(.A(new_n1308), .B(new_n1236), .Y(new_n1309));
  nand_5     g0924(.A(new_n1309), .B(new_n1026), .Y(new_n1310));
  nand_5 g0925(.A(new_n465), .B(new_n465), .Y(new_n1311));
  nand_5     g0926(.A(new_n492), .B(new_n1311), .Y(new_n1312));
  nor_5      g0927(.A(new_n573), .B(new_n465), .Y(new_n1313));
  nand_5     g0928(.A(new_n480), .B(new_n426), .Y(new_n1314));
  nor_5      g0929(.A(new_n1314), .B(new_n1313), .Y(new_n1315));
  nand_5     g0930(.A(new_n1315), .B(new_n1312), .Y(new_n1316));
  nand_5 g0931(.A(pi218), .B(pi218), .Y(new_n1317));
  nor_5      g0932(.A(new_n1317), .B(pi090), .Y(new_n1318));
  nor_5      g0933(.A(new_n1318), .B(new_n420), .Y(new_n1319));
  nor_5      g0934(.A(new_n1319), .B(pi182), .Y(new_n1320));
  nand_5 g0935(.A(pi003), .B(pi003), .Y(new_n1321));
  nand_5     g0936(.A(pi103), .B(new_n1321), .Y(new_n1322));
  nand_5     g0937(.A(new_n1322), .B(new_n409), .Y(new_n1323));
  nand_5 g0938(.A(new_n1323), .B(new_n1323), .Y(new_n1324));
  nand_5     g0939(.A(new_n1324), .B(new_n411), .Y(new_n1325));
  nand_5 g0940(.A(new_n1325), .B(new_n1325), .Y(new_n1326));
  nand_5 g0941(.A(pi081), .B(pi081), .Y(new_n1327));
  nand_5     g0942(.A(new_n1327), .B(new_n1321), .Y(new_n1328));
  nand_5     g0943(.A(new_n1328), .B(new_n1326), .Y(new_n1329));
  nand_5 g0944(.A(new_n1329), .B(new_n1329), .Y(new_n1330));
  nand_5     g0945(.A(new_n1330), .B(new_n416), .Y(new_n1331));
  nand_5 g0946(.A(pi149), .B(pi149), .Y(new_n1332));
  nand_5 g0947(.A(pi075), .B(pi075), .Y(new_n1333));
  nand_5     g0948(.A(new_n1333), .B(pi021), .Y(new_n1334));
  nand_5     g0949(.A(new_n1334), .B(new_n416), .Y(new_n1335));
  nand_5 g0950(.A(new_n1335), .B(new_n1335), .Y(new_n1336));
  nor_5      g0951(.A(pi075), .B(pi022), .Y(new_n1337));
  nand_5 g0952(.A(new_n1337), .B(new_n1337), .Y(new_n1338));
  nand_5     g0953(.A(new_n1338), .B(new_n1336), .Y(new_n1339));
  nand_5     g0954(.A(new_n1339), .B(new_n1332), .Y(new_n1340));
  nand_5 g0955(.A(new_n1340), .B(new_n1340), .Y(new_n1341));
  nand_5     g0956(.A(new_n1341), .B(new_n1317), .Y(new_n1342));
  nand_5 g0957(.A(new_n1342), .B(new_n1342), .Y(new_n1343));
  nand_5     g0958(.A(new_n1343), .B(new_n1331), .Y(new_n1344));
  nand_5     g0959(.A(new_n1344), .B(new_n1320), .Y(new_n1345));
  nand_5     g0960(.A(new_n1345), .B(new_n425), .Y(new_n1346));
  nand_5 g0961(.A(new_n1346), .B(new_n1346), .Y(new_n1347));
  nand_5     g0962(.A(new_n403), .B(new_n392), .Y(new_n1348));
  nor_5      g0963(.A(new_n1348), .B(pi226), .Y(new_n1349));
  nand_5     g0964(.A(pi088), .B(new_n473), .Y(new_n1350));
  nand_5 g0965(.A(pi121), .B(pi121), .Y(new_n1351));
  nand_5     g0966(.A(new_n398), .B(new_n1351), .Y(new_n1352));
  nand_5 g0967(.A(new_n1352), .B(new_n1352), .Y(new_n1353));
  nand_5     g0968(.A(new_n1353), .B(new_n1350), .Y(new_n1354));
  nand_5 g0969(.A(new_n1354), .B(new_n1354), .Y(new_n1355));
  nand_5     g0970(.A(new_n1355), .B(new_n1349), .Y(new_n1356));
  nor_5      g0971(.A(new_n1356), .B(new_n1344), .Y(new_n1357));
  nor_5      g0972(.A(new_n1357), .B(new_n1347), .Y(new_n1358));
  nand_5 g0973(.A(new_n1358), .B(new_n1358), .Y(new_n1359));
  nand_5     g0974(.A(new_n1359), .B(new_n1316), .Y(new_n1360));
  nand_5     g0975(.A(new_n415), .B(pi038), .Y(new_n1361));
  nand_5 g0976(.A(new_n1361), .B(new_n1361), .Y(new_n1362));
  nor_5      g0977(.A(new_n1362), .B(new_n1360), .Y(new_n1363));
  nand_5     g0978(.A(new_n1363), .B(new_n1310), .Y(new_n1364));
  nor_5      g0979(.A(new_n1364), .B(new_n386), .Y(po000));
  nand_5     g0980(.A(new_n928), .B(new_n792), .Y(new_n1366));
  nand_5 g0981(.A(new_n1366), .B(new_n1366), .Y(new_n1367));
  nand_5     g0982(.A(new_n874), .B(new_n813), .Y(new_n1368));
  nor_5      g0983(.A(new_n1368), .B(new_n1367), .Y(new_n1369));
  nand_5 g0984(.A(new_n799), .B(new_n799), .Y(new_n1370));
  nand_5     g0985(.A(new_n1370), .B(new_n780), .Y(new_n1371));
  nand_5     g0986(.A(new_n1371), .B(new_n1173), .Y(new_n1372));
  nand_5     g0987(.A(new_n1372), .B(new_n716), .Y(new_n1373));
  nor_5      g0988(.A(new_n1373), .B(new_n1369), .Y(new_n1374));
  nand_5     g0989(.A(new_n908), .B(new_n732), .Y(new_n1375));
  nand_5 g0990(.A(new_n1375), .B(new_n1375), .Y(new_n1376));
  nand_5     g0991(.A(new_n1376), .B(new_n1374), .Y(new_n1377));
  nand_5     g0992(.A(new_n908), .B(new_n1215), .Y(new_n1378));
  nand_5     g0993(.A(pi225), .B(new_n904), .Y(new_n1379));
  nand_5     g0994(.A(new_n1379), .B(new_n837), .Y(new_n1380));
  nor_5      g0995(.A(new_n1380), .B(pi039), .Y(new_n1381));
  nand_5     g0996(.A(pi054), .B(new_n679), .Y(new_n1382));
  nand_5     g0997(.A(new_n1382), .B(new_n903), .Y(new_n1383));
  nor_5      g0998(.A(new_n1383), .B(new_n1381), .Y(new_n1384));
  nand_5 g0999(.A(new_n1384), .B(new_n1384), .Y(new_n1385));
  nand_5     g1000(.A(new_n1385), .B(new_n1378), .Y(new_n1386));
  nand_5     g1001(.A(new_n1386), .B(new_n865), .Y(new_n1387));
  nand_5     g1002(.A(new_n1387), .B(new_n685), .Y(new_n1388));
  nand_5 g1003(.A(new_n1388), .B(new_n1388), .Y(new_n1389));
  nand_5     g1004(.A(new_n1389), .B(new_n1377), .Y(new_n1390));
  nor_5      g1005(.A(new_n673), .B(new_n615), .Y(new_n1391));
  nand_5 g1006(.A(new_n1391), .B(new_n1391), .Y(new_n1392));
  nand_5     g1007(.A(new_n1392), .B(new_n1390), .Y(new_n1393));
  nand_5 g1008(.A(pi116), .B(pi116), .Y(new_n1394));
  nand_5     g1009(.A(new_n952), .B(new_n1394), .Y(new_n1395));
  nand_5     g1010(.A(new_n1395), .B(new_n1137), .Y(new_n1396));
  nand_5     g1011(.A(new_n1396), .B(new_n742), .Y(new_n1397));
  nand_5 g1012(.A(new_n1397), .B(new_n1397), .Y(new_n1398));
  nand_5     g1013(.A(new_n1398), .B(new_n1138), .Y(new_n1399));
  nor_5      g1014(.A(new_n1368), .B(new_n932), .Y(new_n1400));
  nand_5     g1015(.A(new_n1400), .B(new_n1399), .Y(new_n1401));
  nand_5 g1016(.A(new_n1401), .B(new_n1401), .Y(new_n1402));
  nand_5     g1017(.A(new_n1402), .B(new_n1389), .Y(new_n1403));
  nand_5 g1018(.A(new_n1403), .B(new_n1403), .Y(new_n1404));
  nand_5 g1019(.A(new_n1162), .B(new_n1162), .Y(new_n1405));
  nand_5 g1020(.A(pi131), .B(pi131), .Y(new_n1406));
  nand_5     g1021(.A(new_n415), .B(new_n1406), .Y(new_n1407));
  nand_5 g1022(.A(new_n1407), .B(new_n1407), .Y(new_n1408));
  nand_5 g1023(.A(pi018), .B(pi018), .Y(new_n1409));
  nand_5     g1024(.A(new_n1275), .B(new_n1409), .Y(new_n1410));
  nand_5 g1025(.A(new_n1410), .B(new_n1410), .Y(new_n1411));
  nand_5     g1026(.A(new_n1411), .B(new_n1288), .Y(new_n1412));
  nand_5 g1027(.A(new_n1412), .B(new_n1412), .Y(new_n1413));
  nand_5     g1028(.A(new_n1413), .B(new_n1408), .Y(new_n1414));
  nand_5     g1029(.A(new_n1283), .B(new_n1268), .Y(new_n1415));
  nor_5      g1030(.A(pi238), .B(pi033), .Y(new_n1416));
  nand_5 g1031(.A(new_n1416), .B(new_n1416), .Y(new_n1417));
  nand_5     g1032(.A(new_n1417), .B(new_n1277), .Y(new_n1418));
  nand_5 g1033(.A(new_n1418), .B(new_n1418), .Y(new_n1419));
  nand_5     g1034(.A(new_n1419), .B(new_n1411), .Y(new_n1420));
  nand_5     g1035(.A(new_n1420), .B(new_n1415), .Y(new_n1421));
  nand_5 g1036(.A(new_n1421), .B(new_n1421), .Y(new_n1422));
  nand_5     g1037(.A(new_n1422), .B(new_n1414), .Y(new_n1423));
  nand_5     g1038(.A(new_n1285), .B(new_n1239), .Y(new_n1424));
  nand_5 g1039(.A(new_n1424), .B(new_n1424), .Y(new_n1425));
  nand_5     g1040(.A(new_n1425), .B(new_n1292), .Y(new_n1426));
  nand_5 g1041(.A(new_n1426), .B(new_n1426), .Y(new_n1427));
  nand_5     g1042(.A(new_n1427), .B(new_n1423), .Y(new_n1428));
  nand_5 g1043(.A(new_n1428), .B(new_n1428), .Y(new_n1429));
  nor_5      g1044(.A(new_n1318), .B(pi038), .Y(new_n1430));
  nand_5     g1045(.A(new_n1430), .B(new_n1416), .Y(new_n1431));
  nor_5      g1046(.A(new_n1431), .B(new_n1268), .Y(new_n1432));
  nand_5 g1047(.A(new_n1432), .B(new_n1432), .Y(new_n1433));
  nand_5     g1048(.A(new_n1433), .B(new_n1429), .Y(new_n1434));
  nand_5     g1049(.A(new_n1434), .B(new_n1245), .Y(new_n1435));
  nand_5     g1050(.A(new_n1435), .B(new_n1405), .Y(new_n1436));
  and_6      g1051(.A(new_n1398), .B(new_n1156), .Y(new_n1437));
  nand_5     g1052(.A(new_n1437), .B(new_n1436), .Y(new_n1438));
  and_6      g1053(.A(new_n1438), .B(new_n1404), .Y(new_n1439));
  nor_5      g1054(.A(new_n1439), .B(new_n1393), .Y(new_n1440));
  nand_5 g1055(.A(new_n1228), .B(new_n1228), .Y(new_n1441));
  nand_5 g1056(.A(new_n625), .B(new_n625), .Y(new_n1442));
  nand_5     g1057(.A(new_n987), .B(new_n1442), .Y(new_n1443));
  nand_5 g1058(.A(new_n1443), .B(new_n1443), .Y(new_n1444));
  nor_5      g1059(.A(pi037), .B(pi019), .Y(new_n1445));
  nand_5 g1060(.A(new_n1445), .B(new_n1445), .Y(new_n1446));
  nand_5 g1061(.A(pi118), .B(pi118), .Y(new_n1447));
  nand_5     g1062(.A(new_n700), .B(new_n1447), .Y(new_n1448));
  nor_5      g1063(.A(new_n1448), .B(new_n1446), .Y(new_n1449));
  nand_5     g1064(.A(new_n1449), .B(new_n1444), .Y(new_n1450));
  nand_5     g1065(.A(new_n1450), .B(new_n1441), .Y(new_n1451));
  nand_5 g1066(.A(new_n480), .B(new_n480), .Y(new_n1452));
  nand_5 g1067(.A(new_n464), .B(new_n464), .Y(new_n1453));
  nor_5      g1068(.A(new_n1453), .B(new_n433), .Y(new_n1454));
  nor_5      g1069(.A(new_n1454), .B(new_n1452), .Y(new_n1455));
  nor_5      g1070(.A(new_n1455), .B(new_n1354), .Y(new_n1456));
  nand_5 g1071(.A(pi088), .B(pi088), .Y(new_n1457));
  nand_5     g1072(.A(new_n464), .B(new_n1457), .Y(new_n1458));
  nand_5 g1073(.A(new_n451), .B(new_n451), .Y(new_n1459));
  nand_5     g1074(.A(new_n1353), .B(new_n1459), .Y(new_n1460));
  nor_5      g1075(.A(new_n1460), .B(new_n1458), .Y(new_n1461));
  nand_5 g1076(.A(new_n1461), .B(new_n1461), .Y(new_n1462));
  nand_5 g1077(.A(new_n446), .B(new_n446), .Y(new_n1463));
  nand_5     g1078(.A(new_n1463), .B(new_n436), .Y(new_n1464));
  nor_5      g1079(.A(new_n1464), .B(new_n1462), .Y(new_n1465));
  nor_5      g1080(.A(new_n1465), .B(new_n1456), .Y(new_n1466));
  nand_5 g1081(.A(new_n1466), .B(new_n1466), .Y(new_n1467));
  nand_5 g1082(.A(new_n441), .B(new_n441), .Y(new_n1468));
  nand_5 g1083(.A(new_n482), .B(new_n482), .Y(new_n1469));
  nand_5     g1084(.A(new_n571), .B(new_n1469), .Y(new_n1470));
  nand_5     g1085(.A(new_n1470), .B(new_n1468), .Y(new_n1471));
  nand_5 g1086(.A(new_n1471), .B(new_n1471), .Y(new_n1472));
  nand_5 g1087(.A(pi214), .B(pi214), .Y(new_n1473));
  nand_5     g1088(.A(new_n1473), .B(new_n567), .Y(new_n1474));
  nor_5      g1089(.A(new_n1474), .B(pi204), .Y(new_n1475));
  nand_5     g1090(.A(new_n1475), .B(new_n562), .Y(new_n1476));
  nand_5     g1091(.A(new_n1476), .B(new_n1472), .Y(new_n1477));
  nor_5      g1092(.A(pi237), .B(pi030), .Y(new_n1478));
  nand_5     g1093(.A(new_n1478), .B(new_n1461), .Y(new_n1479));
  nor_5      g1094(.A(new_n1479), .B(new_n1477), .Y(new_n1480));
  nor_5      g1095(.A(new_n1480), .B(new_n1467), .Y(new_n1481));
  nand_5 g1096(.A(new_n1481), .B(new_n1481), .Y(new_n1482));
  nand_5 g1097(.A(new_n1328), .B(new_n1328), .Y(new_n1483));
  nand_5     g1098(.A(new_n405), .B(new_n387), .Y(new_n1484));
  nand_5     g1099(.A(new_n1484), .B(new_n1483), .Y(new_n1485));
  nand_5     g1100(.A(new_n1337), .B(new_n1332), .Y(new_n1486));
  nand_5 g1101(.A(pi038), .B(pi038), .Y(new_n1487));
  nand_5     g1102(.A(new_n1317), .B(new_n1487), .Y(new_n1488));
  nand_5 g1103(.A(new_n1488), .B(new_n1488), .Y(new_n1489));
  nand_5     g1104(.A(new_n1489), .B(new_n1416), .Y(new_n1490));
  nor_5      g1105(.A(new_n1490), .B(new_n1486), .Y(new_n1491));
  nand_5     g1106(.A(new_n1491), .B(new_n392), .Y(new_n1492));
  nor_5      g1107(.A(new_n1492), .B(new_n1485), .Y(new_n1493));
  nand_5     g1108(.A(new_n1493), .B(new_n1482), .Y(new_n1494));
  nand_5 g1109(.A(new_n1494), .B(new_n1494), .Y(new_n1495));
  nand_5 g1110(.A(pi252), .B(pi252), .Y(new_n1496));
  nand_5     g1111(.A(new_n488), .B(new_n1496), .Y(new_n1497));
  nand_5 g1112(.A(new_n1497), .B(new_n1497), .Y(new_n1498));
  nand_5     g1113(.A(new_n1498), .B(new_n1018), .Y(new_n1499));
  nor_5      g1114(.A(new_n1499), .B(new_n698), .Y(new_n1500));
  nand_5     g1115(.A(new_n1500), .B(new_n1495), .Y(new_n1501));
  nand_5 g1116(.A(new_n1501), .B(new_n1501), .Y(new_n1502));
  nand_5     g1117(.A(new_n1502), .B(new_n1451), .Y(new_n1503));
  nand_5     g1118(.A(new_n1495), .B(new_n576), .Y(new_n1504));
  nand_5     g1119(.A(new_n1416), .B(new_n1361), .Y(new_n1505));
  nand_5 g1120(.A(new_n1505), .B(new_n1505), .Y(new_n1506));
  nand_5     g1121(.A(new_n1506), .B(new_n1347), .Y(new_n1507));
  nand_5 g1122(.A(new_n1302), .B(new_n1302), .Y(new_n1508));
  nand_5     g1123(.A(new_n1424), .B(new_n1240), .Y(new_n1509));
  nand_5     g1124(.A(new_n1509), .B(new_n1508), .Y(new_n1510));
  nor_5      g1125(.A(new_n1510), .B(new_n1296), .Y(new_n1511));
  nand_5 g1126(.A(new_n1511), .B(new_n1511), .Y(new_n1512));
  nand_5     g1127(.A(new_n1413), .B(new_n1277), .Y(new_n1513));
  nor_5      g1128(.A(new_n1513), .B(new_n1512), .Y(new_n1514));
  nand_5 g1129(.A(new_n1514), .B(new_n1514), .Y(new_n1515));
  nand_5     g1130(.A(new_n1056), .B(new_n1052), .Y(new_n1516));
  nor_5      g1131(.A(new_n1516), .B(new_n1515), .Y(new_n1517));
  nand_5     g1132(.A(new_n1517), .B(new_n1507), .Y(new_n1518));
  nand_5 g1133(.A(new_n1518), .B(new_n1518), .Y(new_n1519));
  nand_5     g1134(.A(new_n1519), .B(new_n1504), .Y(new_n1520));
  nand_5 g1135(.A(new_n1520), .B(new_n1520), .Y(new_n1521));
  nand_5     g1136(.A(new_n1521), .B(new_n1503), .Y(new_n1522));
  nand_5     g1137(.A(new_n1522), .B(new_n1440), .Y(new_n1523));
  nand_5 g1138(.A(new_n1221), .B(new_n1221), .Y(new_n1524));
  nand_5 g1139(.A(pi026), .B(pi026), .Y(new_n1525));
  nand_5     g1140(.A(new_n634), .B(new_n1525), .Y(new_n1526));
  nand_5 g1141(.A(new_n1526), .B(new_n1526), .Y(new_n1527));
  nand_5     g1142(.A(new_n1527), .B(new_n635), .Y(new_n1528));
  nand_5 g1143(.A(new_n1528), .B(new_n1528), .Y(new_n1529));
  nand_5     g1144(.A(new_n1529), .B(new_n868), .Y(new_n1530));
  nor_5      g1145(.A(new_n1530), .B(new_n677), .Y(new_n1531));
  nand_5     g1146(.A(new_n1531), .B(new_n1524), .Y(new_n1532));
  nand_5 g1147(.A(new_n956), .B(new_n956), .Y(new_n1533));
  nand_5     g1148(.A(new_n1048), .B(pi085), .Y(new_n1534));
  nand_5 g1149(.A(new_n1534), .B(new_n1534), .Y(new_n1535));
  nand_5 g1150(.A(pi170), .B(pi170), .Y(new_n1536));
  nand_5     g1151(.A(new_n957), .B(new_n1536), .Y(new_n1537));
  nor_5      g1152(.A(new_n1537), .B(new_n1535), .Y(new_n1538));
  nand_5     g1153(.A(new_n1056), .B(new_n1043), .Y(new_n1539));
  nand_5 g1154(.A(new_n1539), .B(new_n1539), .Y(new_n1540));
  nand_5     g1155(.A(new_n1295), .B(pi122), .Y(new_n1541));
  nand_5     g1156(.A(new_n1541), .B(new_n1281), .Y(new_n1542));
  nand_5     g1157(.A(new_n1542), .B(new_n1508), .Y(new_n1543));
  nor_5      g1158(.A(new_n1511), .B(new_n1258), .Y(new_n1544));
  nand_5     g1159(.A(new_n1544), .B(new_n1543), .Y(new_n1545));
  nand_5     g1160(.A(new_n1545), .B(new_n1540), .Y(new_n1546));
  nand_5     g1161(.A(new_n1546), .B(new_n1538), .Y(new_n1547));
  nand_5 g1162(.A(new_n1415), .B(new_n1415), .Y(new_n1548));
  nand_5     g1163(.A(new_n1548), .B(new_n1292), .Y(new_n1549));
  nand_5     g1164(.A(new_n1065), .B(new_n1044), .Y(new_n1550));
  nor_5      g1165(.A(new_n1550), .B(new_n1249), .Y(new_n1551));
  nor_5      g1166(.A(new_n1270), .B(new_n1151), .Y(new_n1552));
  nand_5     g1167(.A(new_n1552), .B(new_n1551), .Y(new_n1553));
  nor_5      g1168(.A(new_n1553), .B(new_n1282), .Y(new_n1554));
  nand_5     g1169(.A(new_n1554), .B(new_n1549), .Y(new_n1555));
  nand_5     g1170(.A(new_n1555), .B(new_n1547), .Y(new_n1556));
  nand_5     g1171(.A(new_n1556), .B(new_n1533), .Y(new_n1557));
  nor_5      g1172(.A(new_n1299), .B(pi073), .Y(new_n1558));
  nand_5     g1173(.A(new_n1410), .B(new_n1271), .Y(new_n1559));
  nand_5 g1174(.A(new_n1559), .B(new_n1559), .Y(new_n1560));
  nand_5     g1175(.A(new_n1560), .B(new_n1415), .Y(new_n1561));
  nand_5     g1176(.A(new_n1561), .B(new_n1558), .Y(new_n1562));
  nand_5     g1177(.A(pi090), .B(new_n1487), .Y(new_n1563));
  nand_5     g1178(.A(new_n1563), .B(new_n1408), .Y(new_n1564));
  nand_5 g1179(.A(new_n1564), .B(new_n1564), .Y(new_n1565));
  nand_5     g1180(.A(new_n1336), .B(new_n417), .Y(new_n1566));
  nand_5 g1181(.A(new_n1566), .B(new_n1566), .Y(new_n1567));
  nand_5     g1182(.A(new_n1567), .B(new_n1565), .Y(new_n1568));
  nand_5     g1183(.A(pi149), .B(new_n417), .Y(new_n1569));
  nand_5     g1184(.A(new_n1569), .B(new_n1489), .Y(new_n1570));
  nand_5     g1185(.A(new_n1570), .B(new_n1565), .Y(new_n1571));
  nand_5 g1186(.A(pi099), .B(pi099), .Y(new_n1572));
  nand_5     g1187(.A(new_n1271), .B(new_n1572), .Y(new_n1573));
  nor_5      g1188(.A(new_n1573), .B(new_n1419), .Y(new_n1574));
  nand_5     g1189(.A(new_n1574), .B(new_n1265), .Y(new_n1575));
  nand_5 g1190(.A(new_n1575), .B(new_n1575), .Y(new_n1576));
  nand_5     g1191(.A(new_n1576), .B(new_n1571), .Y(new_n1577));
  nand_5 g1192(.A(new_n1577), .B(new_n1577), .Y(new_n1578));
  nand_5     g1193(.A(new_n1578), .B(new_n1568), .Y(new_n1579));
  nor_5      g1194(.A(new_n1074), .B(new_n1031), .Y(new_n1580));
  nand_5 g1195(.A(new_n1580), .B(new_n1580), .Y(new_n1581));
  nand_5     g1196(.A(new_n1058), .B(new_n1067), .Y(new_n1582));
  nor_5      g1197(.A(new_n1582), .B(new_n1581), .Y(new_n1583));
  nand_5     g1198(.A(new_n1583), .B(new_n1579), .Y(new_n1584));
  nor_5      g1199(.A(new_n1584), .B(new_n1562), .Y(new_n1585));
  nor_5      g1200(.A(new_n1585), .B(new_n1557), .Y(new_n1586));
  nand_5 g1201(.A(new_n967), .B(new_n967), .Y(new_n1587));
  nand_5     g1202(.A(new_n1587), .B(new_n1055), .Y(new_n1588));
  nor_5      g1203(.A(new_n1588), .B(new_n1539), .Y(new_n1589));
  nand_5     g1204(.A(new_n1589), .B(new_n1580), .Y(new_n1590));
  nand_5     g1205(.A(new_n1538), .B(new_n1533), .Y(new_n1591));
  nand_5     g1206(.A(new_n1591), .B(new_n970), .Y(new_n1592));
  nand_5     g1207(.A(new_n966), .B(pi048), .Y(new_n1593));
  nand_5     g1208(.A(new_n1593), .B(new_n1102), .Y(new_n1594));
  nand_5 g1209(.A(new_n1594), .B(new_n1594), .Y(new_n1595));
  and_6      g1210(.A(new_n1595), .B(new_n1592), .Y(new_n1596));
  nand_5     g1211(.A(new_n1596), .B(new_n1590), .Y(new_n1597));
  nand_5     g1212(.A(new_n763), .B(new_n1122), .Y(new_n1598));
  nand_5 g1213(.A(new_n1598), .B(new_n1598), .Y(new_n1599));
  nand_5 g1214(.A(pi150), .B(pi150), .Y(new_n1600));
  nand_5     g1215(.A(pi160), .B(new_n1600), .Y(new_n1601));
  nand_5 g1216(.A(new_n1601), .B(new_n1601), .Y(new_n1602));
  nor_5      g1217(.A(new_n1602), .B(new_n1119), .Y(new_n1603));
  nand_5     g1218(.A(new_n1603), .B(new_n1599), .Y(new_n1604));
  nand_5 g1219(.A(new_n1604), .B(new_n1604), .Y(new_n1605));
  nand_5 g1220(.A(pi209), .B(pi209), .Y(new_n1606));
  nand_5     g1221(.A(new_n784), .B(new_n1606), .Y(new_n1607));
  nor_5      g1222(.A(new_n1607), .B(new_n1101), .Y(new_n1608));
  nand_5     g1223(.A(new_n1608), .B(new_n1605), .Y(new_n1609));
  nand_5 g1224(.A(new_n1609), .B(new_n1609), .Y(new_n1610));
  nand_5     g1225(.A(new_n1610), .B(new_n1597), .Y(new_n1611));
  nor_5      g1226(.A(new_n1611), .B(new_n1586), .Y(new_n1612));
  nand_5     g1227(.A(new_n1118), .B(new_n764), .Y(new_n1613));
  nand_5     g1228(.A(new_n1613), .B(new_n1599), .Y(new_n1614));
  nand_5     g1229(.A(pi046), .B(new_n1122), .Y(new_n1615));
  nand_5 g1230(.A(new_n1615), .B(new_n1615), .Y(new_n1616));
  nand_5 g1231(.A(pi055), .B(pi055), .Y(new_n1617));
  nand_5     g1232(.A(new_n768), .B(new_n1617), .Y(new_n1618));
  nor_5      g1233(.A(new_n1618), .B(new_n1616), .Y(new_n1619));
  nand_5     g1234(.A(new_n1619), .B(new_n1614), .Y(new_n1620));
  nand_5 g1235(.A(new_n1620), .B(new_n1620), .Y(new_n1621));
  nand_5     g1236(.A(new_n807), .B(new_n799), .Y(new_n1622));
  nand_5 g1237(.A(new_n1622), .B(new_n1622), .Y(new_n1623));
  nand_5     g1238(.A(new_n1607), .B(new_n1600), .Y(new_n1624));
  nor_5      g1239(.A(new_n1624), .B(new_n1623), .Y(new_n1625));
  nor_5      g1240(.A(new_n1625), .B(new_n1604), .Y(new_n1626));
  nand_5     g1241(.A(new_n785), .B(new_n794), .Y(new_n1627));
  nor_5      g1242(.A(new_n1627), .B(pi150), .Y(new_n1628));
  nand_5     g1243(.A(new_n1628), .B(new_n1096), .Y(new_n1629));
  nor_5      g1244(.A(new_n1593), .B(new_n1101), .Y(new_n1630));
  nor_5      g1245(.A(new_n1630), .B(new_n1629), .Y(new_n1631));
  nand_5     g1246(.A(new_n1631), .B(new_n1110), .Y(new_n1632));
  nand_5     g1247(.A(new_n1632), .B(new_n1626), .Y(new_n1633));
  nand_5     g1248(.A(new_n1633), .B(new_n1621), .Y(new_n1634));
  nor_5      g1249(.A(new_n1634), .B(new_n1612), .Y(new_n1635));
  nor_5      g1250(.A(new_n1635), .B(new_n1532), .Y(new_n1636));
  nand_5     g1251(.A(new_n1636), .B(new_n1523), .Y(new_n1637));
  nand_5     g1252(.A(new_n676), .B(new_n660), .Y(new_n1638));
  nand_5     g1253(.A(new_n1638), .B(new_n892), .Y(new_n1639));
  nand_5 g1254(.A(new_n1639), .B(new_n1639), .Y(new_n1640));
  nand_5 g1255(.A(pi195), .B(pi195), .Y(new_n1641));
  nand_5     g1256(.A(new_n1385), .B(new_n1641), .Y(new_n1642));
  nand_5     g1257(.A(new_n915), .B(new_n649), .Y(new_n1643));
  nand_5     g1258(.A(new_n666), .B(new_n902), .Y(new_n1644));
  nor_5      g1259(.A(new_n1644), .B(new_n1643), .Y(new_n1645));
  nand_5     g1260(.A(new_n1645), .B(new_n1642), .Y(new_n1646));
  nand_5     g1261(.A(new_n1646), .B(new_n602), .Y(new_n1647));
  nor_5      g1262(.A(new_n1647), .B(new_n1640), .Y(new_n1648));
  nand_5     g1263(.A(new_n1648), .B(new_n592), .Y(new_n1649));
  nand_5     g1264(.A(new_n1649), .B(new_n597), .Y(new_n1650));
  nor_5      g1265(.A(new_n1528), .B(new_n1217), .Y(new_n1651));
  nand_5     g1266(.A(new_n1651), .B(new_n1650), .Y(new_n1652));
  nand_5 g1267(.A(pi063), .B(pi063), .Y(new_n1653));
  nand_5     g1268(.A(new_n580), .B(new_n1653), .Y(new_n1654));
  nand_5 g1269(.A(new_n1654), .B(new_n1654), .Y(new_n1655));
  nand_5     g1270(.A(new_n1176), .B(new_n1525), .Y(new_n1656));
  nand_5     g1271(.A(new_n1656), .B(new_n1655), .Y(new_n1657));
  nand_5 g1272(.A(new_n1657), .B(new_n1657), .Y(new_n1658));
  nand_5     g1273(.A(new_n1658), .B(new_n1652), .Y(new_n1659));
  nand_5 g1274(.A(new_n1659), .B(new_n1659), .Y(new_n1660));
  nand_5     g1275(.A(new_n1660), .B(new_n1637), .Y(new_n1661));
  nand_5 g1276(.A(new_n626), .B(new_n626), .Y(new_n1662));
  nor_5      g1277(.A(new_n624), .B(pi063), .Y(new_n1663));
  nor_5      g1278(.A(new_n1663), .B(new_n1662), .Y(new_n1664));
  nand_5     g1279(.A(new_n1664), .B(new_n1661), .Y(new_n1665));
  and_6      g1280(.A(new_n982), .B(pi174), .Y(new_n1666));
  nand_5     g1281(.A(new_n1666), .B(new_n1665), .Y(new_n1667));
  nand_5 g1282(.A(new_n1667), .B(new_n1667), .Y(po001));
  nand_5 g1283(.A(new_n1626), .B(new_n1626), .Y(new_n1669));
  and_6      g1284(.A(new_n1669), .B(new_n1614), .Y(new_n1670));
  nand_5 g1285(.A(new_n1670), .B(new_n1670), .Y(new_n1671));
  nand_5 g1286(.A(new_n1109), .B(new_n1109), .Y(new_n1672));
  nor_5      g1287(.A(new_n1629), .B(new_n774), .Y(new_n1673));
  nand_5     g1288(.A(new_n1673), .B(new_n1672), .Y(new_n1674));
  nand_5     g1289(.A(new_n1674), .B(new_n1671), .Y(new_n1675));
  nand_5     g1290(.A(new_n1675), .B(new_n1619), .Y(new_n1676));
  nand_5     g1291(.A(new_n1676), .B(new_n1220), .Y(new_n1677));
  nand_5     g1292(.A(new_n1677), .B(new_n1211), .Y(new_n1678));
  nor_5      g1293(.A(new_n1522), .B(new_n1198), .Y(new_n1679));
  nand_5     g1294(.A(new_n1514), .B(new_n1360), .Y(new_n1680));
  nand_5     g1295(.A(new_n1506), .B(new_n1274), .Y(new_n1681));
  and_6      g1296(.A(new_n1681), .B(new_n1279), .Y(new_n1682));
  nand_5     g1297(.A(new_n1682), .B(new_n1303), .Y(new_n1683));
  nand_5 g1298(.A(new_n1683), .B(new_n1683), .Y(new_n1684));
  nand_5     g1299(.A(new_n1102), .B(new_n1041), .Y(new_n1685));
  nor_5      g1300(.A(new_n1685), .B(new_n1166), .Y(new_n1686));
  nand_5     g1301(.A(new_n1686), .B(new_n1038), .Y(new_n1687));
  nand_5 g1302(.A(new_n1687), .B(new_n1687), .Y(new_n1688));
  nand_5     g1303(.A(new_n1688), .B(new_n1259), .Y(new_n1689));
  nor_5      g1304(.A(new_n1689), .B(new_n1684), .Y(new_n1690));
  nand_5     g1305(.A(new_n1690), .B(new_n1680), .Y(new_n1691));
  nor_5      g1306(.A(new_n1691), .B(new_n1679), .Y(new_n1692));
  nand_5 g1307(.A(new_n1611), .B(new_n1611), .Y(new_n1693));
  nand_5     g1308(.A(new_n1693), .B(new_n1220), .Y(new_n1694));
  nor_5      g1309(.A(new_n1694), .B(new_n1692), .Y(new_n1695));
  nor_5      g1310(.A(new_n1695), .B(new_n1678), .Y(new_n1696));
  nand_5 g1311(.A(new_n1696), .B(new_n1696), .Y(new_n1697));
  nand_5     g1312(.A(new_n1697), .B(new_n1207), .Y(new_n1698));
  nand_5     g1313(.A(new_n1698), .B(new_n1202), .Y(new_n1699));
  nand_5     g1314(.A(new_n1215), .B(new_n904), .Y(new_n1700));
  nor_5      g1315(.A(new_n1700), .B(new_n1699), .Y(new_n1701));
  nor_5      g1316(.A(new_n1701), .B(new_n1380), .Y(new_n1702));
  nor_5      g1317(.A(new_n1702), .B(new_n898), .Y(po002));
  nand_5 g1318(.A(pi040), .B(pi040), .Y(new_n1704));
  nand_5 g1319(.A(pi083), .B(pi083), .Y(new_n1705));
  nand_5 g1320(.A(new_n1691), .B(new_n1691), .Y(new_n1706));
  nand_5 g1321(.A(new_n975), .B(new_n975), .Y(new_n1707));
  nor_5      g1322(.A(pi107), .B(pi005), .Y(new_n1708));
  nand_5     g1323(.A(new_n980), .B(new_n1653), .Y(new_n1709));
  nor_5      g1324(.A(new_n1709), .B(pi180), .Y(new_n1710));
  nand_5     g1325(.A(new_n1710), .B(new_n1708), .Y(new_n1711));
  nand_5     g1326(.A(new_n1002), .B(new_n1447), .Y(new_n1712));
  nor_5      g1327(.A(new_n1712), .B(new_n1711), .Y(new_n1713));
  and_6      g1328(.A(new_n1713), .B(new_n1707), .Y(new_n1714));
  nand_5 g1329(.A(new_n1714), .B(new_n1714), .Y(new_n1715));
  nor_5      g1330(.A(new_n1715), .B(new_n1216), .Y(new_n1716));
  nand_5     g1331(.A(new_n1716), .B(new_n1232), .Y(new_n1717));
  nor_5      g1332(.A(new_n1717), .B(new_n1678), .Y(new_n1718));
  nand_5     g1333(.A(new_n1718), .B(new_n1706), .Y(new_n1719));
  nand_5     g1334(.A(new_n1719), .B(new_n1205), .Y(new_n1720));
  nor_5      g1335(.A(new_n1720), .B(new_n1696), .Y(new_n1721));
  nand_5     g1336(.A(new_n1698), .B(new_n855), .Y(new_n1722));
  nor_5      g1337(.A(new_n1722), .B(new_n1721), .Y(new_n1723));
  nand_5     g1338(.A(new_n1723), .B(new_n1705), .Y(new_n1724));
  nand_5     g1339(.A(new_n1724), .B(new_n1704), .Y(new_n1725));
  nor_5      g1340(.A(new_n1725), .B(pi024), .Y(new_n1726));
  nor_5      g1341(.A(new_n1726), .B(new_n845), .Y(new_n1727));
  nor_5      g1342(.A(new_n1727), .B(pi087), .Y(new_n1728));
  nor_5      g1343(.A(new_n1728), .B(new_n720), .Y(po003));
  nand_5 g1344(.A(pi215), .B(pi215), .Y(new_n1730));
  nand_5     g1345(.A(new_n535), .B(pi041), .Y(new_n1731));
  nand_5     g1346(.A(new_n901), .B(new_n676), .Y(new_n1732));
  nand_5     g1347(.A(new_n1732), .B(new_n890), .Y(new_n1733));
  nand_5     g1348(.A(new_n635), .B(new_n604), .Y(new_n1734));
  nand_5 g1349(.A(new_n640), .B(new_n640), .Y(new_n1735));
  nor_5      g1350(.A(new_n1735), .B(new_n599), .Y(new_n1736));
  nor_5      g1351(.A(new_n1736), .B(pi219), .Y(new_n1737));
  nand_5     g1352(.A(new_n1737), .B(new_n1734), .Y(new_n1738));
  nand_5 g1353(.A(new_n1738), .B(new_n1738), .Y(new_n1739));
  nand_5 g1354(.A(pi009), .B(pi009), .Y(new_n1740));
  nand_5     g1355(.A(new_n617), .B(new_n1740), .Y(new_n1741));
  nor_5      g1356(.A(new_n1741), .B(new_n621), .Y(new_n1742));
  nand_5 g1357(.A(new_n1742), .B(new_n1742), .Y(new_n1743));
  nand_5     g1358(.A(new_n1664), .B(new_n625), .Y(new_n1744));
  nor_5      g1359(.A(new_n1744), .B(new_n1743), .Y(new_n1745));
  nand_5     g1360(.A(new_n1745), .B(new_n1527), .Y(new_n1746));
  nor_5      g1361(.A(new_n1746), .B(new_n1739), .Y(new_n1747));
  nand_5     g1362(.A(new_n1747), .B(new_n1733), .Y(new_n1748));
  nand_5 g1363(.A(new_n514), .B(new_n514), .Y(new_n1749));
  nand_5     g1364(.A(new_n1749), .B(new_n501), .Y(new_n1750));
  nand_5 g1365(.A(new_n1750), .B(new_n1750), .Y(new_n1751));
  nand_5     g1366(.A(new_n1751), .B(new_n1010), .Y(new_n1752));
  nand_5 g1367(.A(new_n1752), .B(new_n1752), .Y(new_n1753));
  nor_5      g1368(.A(new_n1753), .B(new_n496), .Y(new_n1754));
  nand_5 g1369(.A(new_n1754), .B(new_n1754), .Y(new_n1755));
  nand_5     g1370(.A(new_n1755), .B(new_n1011), .Y(new_n1756));
  nand_5 g1371(.A(new_n1756), .B(new_n1756), .Y(new_n1757));
  nand_5 g1372(.A(pi106), .B(pi106), .Y(new_n1758));
  nand_5     g1373(.A(new_n691), .B(new_n1758), .Y(new_n1759));
  nor_5      g1374(.A(new_n1759), .B(pi147), .Y(new_n1760));
  nand_5     g1375(.A(new_n1760), .B(new_n1005), .Y(new_n1761));
  nand_5     g1376(.A(new_n1664), .B(new_n1654), .Y(new_n1762));
  nand_5 g1377(.A(new_n1762), .B(new_n1762), .Y(new_n1763));
  nor_5      g1378(.A(new_n1763), .B(new_n983), .Y(new_n1764));
  nand_5     g1379(.A(new_n1764), .B(new_n1708), .Y(new_n1765));
  nand_5     g1380(.A(new_n1443), .B(new_n620), .Y(new_n1766));
  nand_5 g1381(.A(new_n1766), .B(new_n1766), .Y(new_n1767));
  nand_5     g1382(.A(new_n1767), .B(new_n1765), .Y(new_n1768));
  nand_5     g1383(.A(new_n1445), .B(new_n619), .Y(new_n1769));
  nand_5     g1384(.A(pi163), .B(new_n1525), .Y(new_n1770));
  nand_5     g1385(.A(new_n1770), .B(new_n1526), .Y(new_n1771));
  nand_5     g1386(.A(new_n1771), .B(new_n620), .Y(new_n1772));
  nor_5      g1387(.A(new_n1772), .B(new_n629), .Y(new_n1773));
  nand_5 g1388(.A(new_n1773), .B(new_n1773), .Y(new_n1774));
  nand_5     g1389(.A(new_n578), .B(new_n579), .Y(new_n1775));
  nor_5      g1390(.A(new_n1775), .B(new_n638), .Y(new_n1776));
  nor_5      g1391(.A(new_n1776), .B(new_n1774), .Y(new_n1777));
  nor_5      g1392(.A(new_n1777), .B(new_n1769), .Y(new_n1778));
  nand_5     g1393(.A(new_n1778), .B(new_n1768), .Y(new_n1779));
  nor_5      g1394(.A(new_n1779), .B(new_n1761), .Y(new_n1780));
  nand_5     g1395(.A(new_n1780), .B(new_n1757), .Y(new_n1781));
  nand_5     g1396(.A(new_n610), .B(new_n604), .Y(new_n1782));
  nand_5 g1397(.A(new_n1782), .B(new_n1782), .Y(new_n1783));
  nor_5      g1398(.A(new_n1783), .B(new_n598), .Y(new_n1784));
  nand_5     g1399(.A(new_n1773), .B(new_n635), .Y(new_n1785));
  nor_5      g1400(.A(new_n1785), .B(new_n1784), .Y(new_n1786));
  nor_5      g1401(.A(new_n1786), .B(new_n1781), .Y(new_n1787));
  nand_5     g1402(.A(new_n1787), .B(new_n1748), .Y(new_n1788));
  nand_5 g1403(.A(new_n500), .B(new_n500), .Y(new_n1789));
  nand_5     g1404(.A(new_n707), .B(new_n1789), .Y(new_n1790));
  nand_5     g1405(.A(new_n1016), .B(new_n1005), .Y(new_n1791));
  nand_5     g1406(.A(new_n1791), .B(new_n1789), .Y(new_n1792));
  nand_5     g1407(.A(new_n1792), .B(new_n1790), .Y(new_n1793));
  nand_5     g1408(.A(new_n1793), .B(new_n493), .Y(new_n1794));
  nand_5     g1409(.A(pi169), .B(new_n996), .Y(new_n1795));
  nor_5      g1410(.A(new_n1795), .B(new_n1761), .Y(new_n1796));
  nor_5      g1411(.A(new_n1796), .B(new_n1794), .Y(new_n1797));
  nor_5      g1412(.A(new_n1797), .B(new_n1756), .Y(new_n1798));
  nand_5     g1413(.A(new_n507), .B(pi007), .Y(new_n1799));
  nand_5     g1414(.A(new_n1799), .B(new_n543), .Y(new_n1800));
  nor_5      g1415(.A(new_n1800), .B(new_n1798), .Y(new_n1801));
  nand_5     g1416(.A(new_n1801), .B(new_n1788), .Y(new_n1802));
  nand_5 g1417(.A(new_n1802), .B(new_n1802), .Y(new_n1803));
  nand_5     g1418(.A(new_n773), .B(new_n1600), .Y(new_n1804));
  nand_5 g1419(.A(new_n1804), .B(new_n1804), .Y(new_n1805));
  nand_5     g1420(.A(new_n1805), .B(new_n1622), .Y(new_n1806));
  nand_5     g1421(.A(new_n803), .B(new_n781), .Y(new_n1807));
  nor_5      g1422(.A(new_n1807), .B(new_n1112), .Y(new_n1808));
  nor_5      g1423(.A(new_n1808), .B(new_n1806), .Y(new_n1809));
  nand_5 g1424(.A(new_n1030), .B(new_n1030), .Y(new_n1810));
  nand_5     g1425(.A(new_n1593), .B(new_n967), .Y(new_n1811));
  nor_5      g1426(.A(new_n1807), .B(pi015), .Y(new_n1812));
  nand_5     g1427(.A(new_n1812), .B(new_n1811), .Y(new_n1813));
  nor_5      g1428(.A(new_n1813), .B(new_n1810), .Y(new_n1814));
  nand_5 g1429(.A(new_n1814), .B(new_n1814), .Y(new_n1815));
  nand_5     g1430(.A(new_n1815), .B(new_n1809), .Y(new_n1816));
  nand_5     g1431(.A(new_n834), .B(new_n826), .Y(new_n1817));
  nand_5     g1432(.A(new_n1817), .B(new_n838), .Y(new_n1818));
  nor_5      g1433(.A(new_n1818), .B(new_n1127), .Y(new_n1819));
  nand_5     g1434(.A(new_n1819), .B(new_n1816), .Y(new_n1820));
  nand_5 g1435(.A(new_n1806), .B(new_n1806), .Y(new_n1821));
  nand_5 g1436(.A(new_n1112), .B(new_n1112), .Y(new_n1822));
  nand_5 g1437(.A(new_n1807), .B(new_n1807), .Y(new_n1823));
  nand_5     g1438(.A(new_n1823), .B(new_n1822), .Y(new_n1824));
  nand_5     g1439(.A(new_n1824), .B(new_n1821), .Y(new_n1825));
  nor_5      g1440(.A(new_n970), .B(pi048), .Y(new_n1826));
  nand_5     g1441(.A(new_n1069), .B(new_n1058), .Y(new_n1827));
  nand_5     g1442(.A(new_n1827), .B(new_n1167), .Y(new_n1828));
  nand_5     g1443(.A(new_n1828), .B(new_n1814), .Y(new_n1829));
  nor_5      g1444(.A(new_n1829), .B(new_n1826), .Y(new_n1830));
  nor_5      g1445(.A(new_n1830), .B(new_n1825), .Y(new_n1831));
  nor_5      g1446(.A(new_n1831), .B(new_n1820), .Y(new_n1832));
  nand_5 g1447(.A(new_n1142), .B(new_n1142), .Y(new_n1833));
  nand_5     g1448(.A(new_n1281), .B(new_n1833), .Y(new_n1834));
  nand_5     g1449(.A(new_n1834), .B(new_n1084), .Y(new_n1835));
  nand_5     g1450(.A(new_n1835), .B(new_n1065), .Y(new_n1836));
  nor_5      g1451(.A(new_n1836), .B(new_n1168), .Y(new_n1837));
  nand_5     g1452(.A(new_n1837), .B(new_n1809), .Y(new_n1838));
  nand_5     g1453(.A(new_n1838), .B(new_n1832), .Y(new_n1839));
  nand_5 g1454(.A(new_n849), .B(new_n849), .Y(new_n1840));
  nand_5 g1455(.A(new_n1818), .B(new_n1818), .Y(new_n1841));
  nand_5     g1456(.A(new_n1841), .B(new_n1840), .Y(new_n1842));
  nand_5     g1457(.A(new_n838), .B(pi173), .Y(new_n1843));
  nand_5     g1458(.A(new_n1843), .B(new_n906), .Y(new_n1844));
  nand_5 g1459(.A(new_n1844), .B(new_n1844), .Y(new_n1845));
  nand_5     g1460(.A(new_n1845), .B(new_n1842), .Y(new_n1846));
  nand_5 g1461(.A(new_n1846), .B(new_n1846), .Y(new_n1847));
  nand_5     g1462(.A(new_n1847), .B(new_n1839), .Y(new_n1848));
  nand_5 g1463(.A(new_n719), .B(new_n719), .Y(new_n1849));
  nand_5     g1464(.A(new_n874), .B(new_n771), .Y(new_n1850));
  nand_5 g1465(.A(new_n726), .B(new_n726), .Y(new_n1851));
  nand_5     g1466(.A(new_n1851), .B(new_n716), .Y(new_n1852));
  nand_5 g1467(.A(new_n1852), .B(new_n1852), .Y(new_n1853));
  nand_5     g1468(.A(new_n1853), .B(new_n1850), .Y(new_n1854));
  nand_5     g1469(.A(new_n1854), .B(new_n862), .Y(new_n1855));
  nand_5     g1470(.A(new_n1855), .B(new_n1849), .Y(new_n1856));
  nand_5     g1471(.A(new_n1856), .B(new_n847), .Y(new_n1857));
  nor_5      g1472(.A(new_n1857), .B(new_n1818), .Y(new_n1858));
  nor_5      g1473(.A(new_n1858), .B(new_n1848), .Y(new_n1859));
  nor_5      g1474(.A(new_n1643), .B(new_n896), .Y(new_n1860));
  nand_5 g1475(.A(new_n1860), .B(new_n1860), .Y(new_n1861));
  nor_5      g1476(.A(new_n1861), .B(new_n670), .Y(new_n1862));
  nand_5     g1477(.A(new_n1862), .B(new_n1859), .Y(new_n1863));
  nor_5      g1478(.A(new_n1863), .B(new_n1781), .Y(new_n1864));
  nand_5 g1479(.A(new_n1585), .B(new_n1585), .Y(new_n1865));
  nor_5      g1480(.A(new_n1820), .B(new_n1865), .Y(new_n1866));
  nand_5     g1481(.A(new_n1551), .B(new_n1265), .Y(new_n1867));
  nand_5 g1482(.A(new_n1867), .B(new_n1867), .Y(new_n1868));
  nand_5 g1483(.A(new_n1273), .B(new_n1273), .Y(new_n1869));
  nand_5     g1484(.A(new_n1869), .B(new_n1572), .Y(new_n1870));
  nor_5      g1485(.A(new_n1870), .B(new_n1505), .Y(new_n1871));
  nand_5     g1486(.A(new_n1871), .B(new_n1868), .Y(new_n1872));
  nor_5      g1487(.A(new_n1872), .B(new_n1358), .Y(new_n1873));
  nand_5 g1488(.A(new_n1873), .B(new_n1873), .Y(new_n1874));
  nor_5      g1489(.A(new_n1874), .B(new_n1315), .Y(new_n1875));
  nor_5      g1490(.A(new_n1590), .B(new_n929), .Y(new_n1876));
  nand_5     g1491(.A(new_n1876), .B(new_n1305), .Y(new_n1877));
  nor_5      g1492(.A(new_n1877), .B(new_n1875), .Y(new_n1878));
  nand_5     g1493(.A(new_n1485), .B(new_n1324), .Y(new_n1879));
  nand_5     g1494(.A(new_n1879), .B(new_n1337), .Y(new_n1880));
  nand_5 g1495(.A(new_n1880), .B(new_n1880), .Y(new_n1881));
  nor_5      g1496(.A(new_n410), .B(new_n396), .Y(new_n1882));
  nand_5 g1497(.A(pi117), .B(pi117), .Y(new_n1883));
  nand_5     g1498(.A(pi121), .B(new_n1883), .Y(new_n1884));
  nand_5 g1499(.A(new_n1884), .B(new_n1884), .Y(new_n1885));
  nor_5      g1500(.A(new_n1885), .B(new_n399), .Y(new_n1886));
  nand_5 g1501(.A(new_n1886), .B(new_n1886), .Y(new_n1887));
  nand_5     g1502(.A(new_n1887), .B(new_n1882), .Y(new_n1888));
  nand_5     g1503(.A(new_n1888), .B(new_n1881), .Y(new_n1889));
  nand_5 g1504(.A(new_n1889), .B(new_n1889), .Y(new_n1890));
  nand_5 g1505(.A(new_n432), .B(new_n432), .Y(new_n1891));
  nand_5     g1506(.A(new_n451), .B(new_n1891), .Y(new_n1892));
  nand_5     g1507(.A(new_n1892), .B(new_n458), .Y(new_n1893));
  nand_5     g1508(.A(new_n458), .B(pi120), .Y(new_n1894));
  nand_5     g1509(.A(new_n1894), .B(new_n466), .Y(new_n1895));
  nand_5 g1510(.A(new_n1895), .B(new_n1895), .Y(new_n1896));
  nand_5     g1511(.A(new_n1896), .B(new_n1893), .Y(new_n1897));
  nand_5 g1512(.A(pi207), .B(pi207), .Y(new_n1898));
  nand_5     g1513(.A(new_n1898), .B(new_n468), .Y(new_n1899));
  nand_5 g1514(.A(new_n1899), .B(new_n1899), .Y(new_n1900));
  nand_5 g1515(.A(new_n477), .B(new_n477), .Y(new_n1901));
  nand_5     g1516(.A(new_n1883), .B(new_n473), .Y(new_n1902));
  nand_5 g1517(.A(new_n1902), .B(new_n1902), .Y(new_n1903));
  nand_5     g1518(.A(new_n1903), .B(new_n1901), .Y(new_n1904));
  nand_5 g1519(.A(new_n1904), .B(new_n1904), .Y(new_n1905));
  nand_5     g1520(.A(new_n1905), .B(new_n1900), .Y(new_n1906));
  nand_5 g1521(.A(new_n1906), .B(new_n1906), .Y(new_n1907));
  nand_5     g1522(.A(new_n1907), .B(new_n1882), .Y(new_n1908));
  nor_5      g1523(.A(new_n1908), .B(new_n1897), .Y(new_n1909));
  nand_5     g1524(.A(new_n475), .B(new_n1457), .Y(new_n1910));
  nand_5 g1525(.A(new_n1910), .B(new_n1910), .Y(new_n1911));
  nand_5     g1526(.A(pi232), .B(new_n1898), .Y(new_n1912));
  nand_5     g1527(.A(new_n1912), .B(new_n459), .Y(new_n1913));
  nand_5 g1528(.A(new_n1913), .B(new_n1913), .Y(new_n1914));
  nand_5     g1529(.A(new_n1914), .B(new_n455), .Y(new_n1915));
  nand_5     g1530(.A(new_n455), .B(pi012), .Y(new_n1916));
  nand_5     g1531(.A(new_n1916), .B(new_n1901), .Y(new_n1917));
  nand_5 g1532(.A(new_n1917), .B(new_n1917), .Y(new_n1918));
  nand_5     g1533(.A(new_n1918), .B(new_n1915), .Y(new_n1919));
  nand_5     g1534(.A(new_n1919), .B(new_n1911), .Y(new_n1920));
  nand_5     g1535(.A(new_n1903), .B(new_n1882), .Y(new_n1921));
  nand_5 g1536(.A(new_n1921), .B(new_n1921), .Y(new_n1922));
  nand_5     g1537(.A(new_n1922), .B(new_n1920), .Y(new_n1923));
  nand_5 g1538(.A(new_n1923), .B(new_n1923), .Y(new_n1924));
  nor_5      g1539(.A(new_n1924), .B(new_n1909), .Y(new_n1925));
  nand_5     g1540(.A(new_n1925), .B(new_n1890), .Y(new_n1926));
  nor_5      g1541(.A(pi239), .B(pi010), .Y(new_n1927));
  nand_5 g1542(.A(new_n1927), .B(new_n1927), .Y(new_n1928));
  nand_5     g1543(.A(new_n1478), .B(new_n482), .Y(new_n1929));
  nor_5      g1544(.A(new_n1929), .B(new_n1928), .Y(new_n1930));
  nand_5     g1545(.A(new_n1930), .B(new_n1578), .Y(new_n1931));
  nor_5      g1546(.A(new_n1931), .B(new_n1926), .Y(new_n1932));
  nor_5      g1547(.A(new_n531), .B(pi105), .Y(new_n1933));
  nand_5     g1548(.A(new_n1475), .B(new_n435), .Y(new_n1934));
  nand_5     g1549(.A(pi255), .B(new_n486), .Y(new_n1935));
  nand_5     g1550(.A(new_n1935), .B(new_n557), .Y(new_n1936));
  nor_5      g1551(.A(new_n1936), .B(new_n1934), .Y(new_n1937));
  nand_5     g1552(.A(new_n1937), .B(new_n1933), .Y(new_n1938));
  nand_5 g1553(.A(new_n489), .B(new_n489), .Y(new_n1939));
  nand_5 g1554(.A(new_n533), .B(new_n533), .Y(new_n1940));
  nand_5     g1555(.A(new_n1940), .B(new_n519), .Y(new_n1941));
  nand_5     g1556(.A(new_n1941), .B(new_n1939), .Y(new_n1942));
  nand_5     g1557(.A(new_n559), .B(new_n558), .Y(new_n1943));
  nand_5     g1558(.A(new_n1943), .B(new_n1942), .Y(new_n1944));
  nand_5     g1559(.A(new_n1944), .B(new_n563), .Y(new_n1945));
  nand_5     g1560(.A(new_n1945), .B(new_n1473), .Y(new_n1946));
  and_6      g1561(.A(new_n1946), .B(new_n1938), .Y(new_n1947));
  nand_5     g1562(.A(new_n1947), .B(new_n1932), .Y(new_n1948));
  and_6      g1563(.A(new_n1948), .B(new_n1878), .Y(new_n1949));
  nand_5     g1564(.A(new_n1949), .B(new_n1866), .Y(new_n1950));
  nand_5     g1565(.A(new_n1950), .B(new_n1864), .Y(new_n1951));
  nand_5     g1566(.A(new_n1951), .B(new_n1803), .Y(new_n1952));
  nand_5     g1567(.A(new_n1952), .B(new_n1731), .Y(new_n1953));
  nor_5      g1568(.A(new_n1953), .B(new_n1730), .Y(po004));
  nand_5 g1569(.A(new_n435), .B(new_n435), .Y(new_n1955));
  or_6       g1570(.A(new_n572), .B(new_n492), .Y(new_n1956));
  nand_5 g1571(.A(new_n1309), .B(new_n1309), .Y(new_n1957));
  nand_5 g1572(.A(new_n1590), .B(new_n1590), .Y(new_n1958));
  nand_5     g1573(.A(new_n1514), .B(new_n1320), .Y(new_n1959));
  nand_5     g1574(.A(new_n1959), .B(new_n1683), .Y(new_n1960));
  nand_5     g1575(.A(new_n1960), .B(new_n1958), .Y(new_n1961));
  nand_5     g1576(.A(new_n1961), .B(new_n1256), .Y(new_n1962));
  nand_5 g1577(.A(new_n1475), .B(new_n1475), .Y(new_n1963));
  nand_5 g1578(.A(new_n1943), .B(new_n1943), .Y(new_n1964));
  nand_5 g1579(.A(new_n547), .B(new_n547), .Y(new_n1965));
  nor_5      g1580(.A(new_n1965), .B(new_n524), .Y(new_n1966));
  nor_5      g1581(.A(new_n1966), .B(new_n489), .Y(new_n1967));
  nor_5      g1582(.A(new_n1967), .B(new_n1964), .Y(new_n1968));
  nand_5 g1583(.A(new_n1968), .B(new_n1968), .Y(new_n1969));
  nand_5 g1584(.A(new_n1933), .B(new_n1933), .Y(new_n1970));
  nand_5     g1585(.A(new_n557), .B(new_n483), .Y(new_n1971));
  nor_5      g1586(.A(new_n1971), .B(new_n1970), .Y(new_n1972));
  nand_5     g1587(.A(new_n1972), .B(new_n1225), .Y(new_n1973));
  and_6      g1588(.A(new_n1973), .B(new_n1969), .Y(new_n1974));
  nor_5      g1589(.A(new_n1974), .B(new_n1963), .Y(new_n1975));
  nand_5     g1590(.A(new_n1975), .B(new_n1962), .Y(new_n1976));
  nor_5      g1591(.A(new_n1976), .B(new_n1957), .Y(new_n1977));
  nand_5     g1592(.A(new_n1902), .B(new_n1886), .Y(new_n1978));
  nand_5     g1593(.A(new_n1978), .B(new_n397), .Y(new_n1979));
  nand_5 g1594(.A(new_n1979), .B(new_n1979), .Y(new_n1980));
  nor_5      g1595(.A(new_n1980), .B(new_n1485), .Y(new_n1981));
  nand_5     g1596(.A(new_n1326), .B(new_n422), .Y(new_n1982));
  nor_5      g1597(.A(new_n1982), .B(new_n1981), .Y(new_n1983));
  nand_5     g1598(.A(new_n1983), .B(new_n1466), .Y(new_n1984));
  nand_5 g1599(.A(new_n1251), .B(new_n1251), .Y(new_n1985));
  nand_5     g1600(.A(new_n1340), .B(new_n420), .Y(new_n1986));
  nand_5     g1601(.A(new_n1986), .B(new_n1432), .Y(new_n1987));
  nand_5 g1602(.A(new_n1987), .B(new_n1987), .Y(new_n1988));
  nand_5     g1603(.A(new_n1988), .B(new_n1985), .Y(new_n1989));
  nand_5 g1604(.A(new_n1989), .B(new_n1989), .Y(new_n1990));
  nand_5     g1605(.A(new_n1349), .B(new_n1483), .Y(new_n1991));
  nand_5 g1606(.A(new_n1991), .B(new_n1991), .Y(new_n1992));
  nand_5     g1607(.A(new_n1992), .B(new_n1353), .Y(new_n1993));
  nor_5      g1608(.A(new_n1993), .B(new_n1920), .Y(new_n1994));
  nand_5 g1609(.A(new_n1994), .B(new_n1994), .Y(new_n1995));
  nand_5     g1610(.A(new_n1995), .B(new_n1983), .Y(new_n1996));
  nand_5     g1611(.A(new_n1996), .B(new_n1990), .Y(new_n1997));
  nand_5 g1612(.A(new_n1997), .B(new_n1997), .Y(new_n1998));
  and_6      g1613(.A(new_n1998), .B(new_n1984), .Y(new_n1999));
  nand_5     g1614(.A(new_n1999), .B(new_n1256), .Y(new_n2000));
  nand_5     g1615(.A(new_n2000), .B(new_n1977), .Y(new_n2001));
  nand_5     g1616(.A(new_n2001), .B(new_n1956), .Y(new_n2002));
  nor_5      g1617(.A(new_n2002), .B(new_n441), .Y(new_n2003));
  nor_5      g1618(.A(new_n2003), .B(new_n1955), .Y(new_n2004));
  nand_5 g1619(.A(new_n444), .B(new_n444), .Y(new_n2005));
  nand_5     g1620(.A(new_n2005), .B(pi030), .Y(new_n2006));
  nor_5      g1621(.A(new_n2006), .B(new_n2004), .Y(po005));
  nand_5 g1622(.A(pi206), .B(pi206), .Y(new_n2008));
  nand_5     g1623(.A(new_n1364), .B(new_n1406), .Y(new_n2009));
  nand_5     g1624(.A(new_n2009), .B(new_n1418), .Y(new_n2010));
  nand_5     g1625(.A(new_n2010), .B(new_n1275), .Y(new_n2011));
  nand_5     g1626(.A(new_n2011), .B(new_n1267), .Y(new_n2012));
  nor_5      g1627(.A(new_n2012), .B(new_n2008), .Y(po006));
  nand_5     g1628(.A(new_n594), .B(pi189), .Y(new_n2014));
  nand_5     g1629(.A(new_n1714), .B(new_n593), .Y(new_n2015));
  nand_5 g1630(.A(new_n647), .B(new_n647), .Y(new_n2016));
  nand_5 g1631(.A(new_n1003), .B(new_n1003), .Y(new_n2017));
  nand_5     g1632(.A(new_n2017), .B(new_n2016), .Y(new_n2018));
  nand_5     g1633(.A(new_n547), .B(new_n497), .Y(new_n2019));
  nor_5      g1634(.A(new_n2019), .B(new_n1790), .Y(new_n2020));
  nand_5     g1635(.A(new_n2020), .B(new_n2018), .Y(new_n2021));
  nand_5 g1636(.A(new_n2021), .B(new_n2021), .Y(new_n2022));
  nand_5     g1637(.A(new_n2022), .B(new_n2015), .Y(new_n2023));
  nor_5      g1638(.A(new_n1232), .B(new_n533), .Y(new_n2024));
  nand_5     g1639(.A(new_n1930), .B(new_n1459), .Y(new_n2025));
  nand_5     g1640(.A(new_n490), .B(new_n464), .Y(new_n2026));
  nor_5      g1641(.A(new_n2026), .B(new_n2025), .Y(new_n2027));
  nand_5 g1642(.A(new_n2027), .B(new_n2027), .Y(new_n2028));
  nor_5      g1643(.A(new_n2028), .B(new_n2024), .Y(new_n2029));
  nand_5     g1644(.A(new_n2029), .B(new_n1873), .Y(new_n2030));
  nand_5 g1645(.A(new_n2030), .B(new_n2030), .Y(new_n2031));
  nand_5     g1646(.A(new_n2031), .B(new_n2023), .Y(new_n2032));
  nand_5     g1647(.A(new_n2032), .B(new_n1878), .Y(new_n2033));
  nand_5 g1648(.A(new_n1674), .B(new_n1674), .Y(new_n2034));
  nand_5 g1649(.A(new_n1596), .B(new_n1596), .Y(new_n2035));
  nand_5     g1650(.A(new_n2035), .B(new_n1100), .Y(new_n2036));
  nand_5     g1651(.A(new_n2036), .B(new_n2034), .Y(new_n2037));
  nand_5 g1652(.A(new_n2037), .B(new_n2037), .Y(new_n2038));
  nand_5     g1653(.A(new_n2038), .B(new_n2033), .Y(new_n2039));
  nand_5 g1654(.A(new_n1673), .B(new_n1673), .Y(new_n2040));
  nand_5     g1655(.A(new_n1104), .B(new_n1028), .Y(new_n2041));
  nor_5      g1656(.A(new_n2041), .B(new_n2040), .Y(new_n2042));
  nor_5      g1657(.A(new_n2042), .B(new_n1670), .Y(new_n2043));
  nand_5 g1658(.A(new_n2043), .B(new_n2043), .Y(new_n2044));
  nor_5      g1659(.A(new_n2044), .B(new_n1221), .Y(new_n2045));
  nand_5     g1660(.A(new_n2045), .B(new_n2039), .Y(new_n2046));
  nor_5      g1661(.A(new_n1619), .B(new_n1221), .Y(new_n2047));
  nor_5      g1662(.A(new_n2047), .B(new_n1214), .Y(new_n2048));
  nand_5 g1663(.A(new_n2048), .B(new_n2048), .Y(new_n2049));
  nand_5 g1664(.A(new_n1378), .B(new_n1378), .Y(new_n2050));
  nand_5     g1665(.A(new_n1645), .B(new_n2050), .Y(new_n2051));
  nor_5      g1666(.A(new_n2051), .B(new_n2049), .Y(new_n2052));
  nand_5     g1667(.A(new_n2052), .B(new_n2046), .Y(new_n2053));
  nand_5     g1668(.A(new_n2053), .B(new_n1648), .Y(new_n2054));
  nand_5     g1669(.A(new_n2054), .B(new_n2014), .Y(new_n2055));
  nor_5      g1670(.A(new_n2055), .B(pi129), .Y(new_n2056));
  nor_5      g1671(.A(new_n2056), .B(pi057), .Y(new_n2057));
  nor_5      g1672(.A(new_n2057), .B(new_n667), .Y(po007));
  nand_5 g1673(.A(new_n1532), .B(new_n1532), .Y(new_n2059));
  nand_5     g1674(.A(new_n1820), .B(new_n1621), .Y(new_n2060));
  nand_5     g1675(.A(new_n2060), .B(new_n2059), .Y(new_n2061));
  nand_5 g1676(.A(new_n1759), .B(new_n1759), .Y(new_n2062));
  nand_5     g1677(.A(new_n2062), .B(new_n1449), .Y(new_n2063));
  nand_5 g1678(.A(new_n2063), .B(new_n2063), .Y(new_n2064));
  nand_5     g1679(.A(new_n2064), .B(new_n989), .Y(new_n2065));
  nor_5      g1680(.A(new_n2065), .B(new_n1659), .Y(new_n2066));
  nand_5     g1681(.A(new_n2066), .B(new_n2061), .Y(new_n2067));
  nand_5 g1682(.A(new_n1745), .B(new_n1745), .Y(new_n2068));
  nand_5     g1683(.A(new_n1795), .B(new_n1740), .Y(new_n2069));
  nand_5 g1684(.A(new_n2069), .B(new_n2069), .Y(new_n2070));
  nand_5 g1685(.A(new_n1769), .B(new_n1769), .Y(new_n2071));
  nand_5     g1686(.A(new_n988), .B(new_n620), .Y(new_n2072));
  nand_5     g1687(.A(new_n2072), .B(new_n2071), .Y(new_n2073));
  nand_5     g1688(.A(new_n2073), .B(new_n2070), .Y(new_n2074));
  nand_5     g1689(.A(new_n2074), .B(new_n1760), .Y(new_n2075));
  nand_5 g1690(.A(new_n2075), .B(new_n2075), .Y(new_n2076));
  nand_5     g1691(.A(new_n2076), .B(new_n2068), .Y(new_n2077));
  nand_5 g1692(.A(new_n2077), .B(new_n2077), .Y(new_n2078));
  nand_5     g1693(.A(new_n493), .B(new_n508), .Y(new_n2079));
  nor_5      g1694(.A(new_n514), .B(new_n499), .Y(new_n2080));
  nor_5      g1695(.A(new_n2080), .B(new_n2079), .Y(new_n2081));
  nand_5 g1696(.A(new_n2081), .B(new_n2081), .Y(new_n2082));
  nand_5     g1697(.A(new_n545), .B(new_n530), .Y(new_n2083));
  nor_5      g1698(.A(new_n2083), .B(new_n2082), .Y(new_n2084));
  nand_5     g1699(.A(new_n498), .B(new_n1015), .Y(new_n2085));
  nand_5     g1700(.A(new_n704), .B(new_n1758), .Y(new_n2086));
  nor_5      g1701(.A(new_n2086), .B(new_n698), .Y(new_n2087));
  nor_5      g1702(.A(new_n2087), .B(new_n2085), .Y(new_n2088));
  nand_5     g1703(.A(new_n2088), .B(new_n2084), .Y(new_n2089));
  nor_5      g1704(.A(new_n2089), .B(new_n2078), .Y(new_n2090));
  nand_5     g1705(.A(new_n2090), .B(new_n2067), .Y(new_n2091));
  nand_5     g1706(.A(new_n1922), .B(new_n1567), .Y(new_n2092));
  nand_5 g1707(.A(new_n2092), .B(new_n2092), .Y(new_n2093));
  nand_5     g1708(.A(new_n480), .B(new_n1453), .Y(new_n2094));
  nand_5     g1709(.A(new_n2094), .B(new_n1457), .Y(new_n2095));
  nand_5     g1710(.A(new_n2095), .B(new_n2093), .Y(new_n2096));
  nand_5 g1711(.A(new_n2096), .B(new_n2096), .Y(new_n2097));
  nand_5 g1712(.A(new_n1570), .B(new_n1570), .Y(new_n2098));
  nand_5     g1713(.A(new_n1889), .B(new_n1567), .Y(new_n2099));
  nand_5     g1714(.A(new_n2099), .B(new_n2098), .Y(new_n2100));
  nor_5      g1715(.A(new_n2100), .B(new_n2097), .Y(new_n2101));
  nand_5     g1716(.A(new_n512), .B(new_n541), .Y(new_n2102));
  nand_5     g1717(.A(new_n2102), .B(new_n516), .Y(new_n2103));
  nand_5     g1718(.A(new_n537), .B(new_n530), .Y(new_n2104));
  nand_5 g1719(.A(new_n2104), .B(new_n2104), .Y(new_n2105));
  nand_5     g1720(.A(new_n2105), .B(new_n2103), .Y(new_n2106));
  nand_5 g1721(.A(new_n2106), .B(new_n2106), .Y(new_n2107));
  nand_5     g1722(.A(new_n498), .B(pi043), .Y(new_n2108));
  nand_5     g1723(.A(new_n2108), .B(new_n1008), .Y(new_n2109));
  nand_5     g1724(.A(new_n2109), .B(new_n2084), .Y(new_n2110));
  nand_5 g1725(.A(new_n2110), .B(new_n2110), .Y(new_n2111));
  nor_5      g1726(.A(new_n2111), .B(new_n2025), .Y(new_n2112));
  nand_5     g1727(.A(new_n2112), .B(new_n1946), .Y(new_n2113));
  nor_5      g1728(.A(new_n2113), .B(new_n2107), .Y(new_n2114));
  nand_5     g1729(.A(new_n2114), .B(new_n2101), .Y(new_n2115));
  nand_5 g1730(.A(new_n2115), .B(new_n2115), .Y(new_n2116));
  nand_5     g1731(.A(new_n2116), .B(new_n2091), .Y(new_n2117));
  nand_5 g1732(.A(new_n2117), .B(new_n2117), .Y(new_n2118));
  nand_5 g1733(.A(new_n1934), .B(new_n1934), .Y(new_n2119));
  nand_5     g1734(.A(new_n466), .B(new_n549), .Y(new_n2120));
  nor_5      g1735(.A(new_n2120), .B(new_n550), .Y(new_n2121));
  nand_5     g1736(.A(new_n2121), .B(new_n2119), .Y(new_n2122));
  nand_5 g1737(.A(new_n2122), .B(new_n2122), .Y(new_n2123));
  nor_5      g1738(.A(new_n1971), .B(pi067), .Y(new_n2124));
  nand_5     g1739(.A(new_n2124), .B(new_n2123), .Y(new_n2125));
  nand_5 g1740(.A(new_n2125), .B(new_n2125), .Y(new_n2126));
  nand_5     g1741(.A(new_n2126), .B(new_n1900), .Y(new_n2127));
  nor_5      g1742(.A(new_n1313), .B(new_n472), .Y(new_n2128));
  nand_5     g1743(.A(new_n2128), .B(new_n1312), .Y(new_n2129));
  nand_5     g1744(.A(new_n2129), .B(new_n2127), .Y(new_n2130));
  nand_5     g1745(.A(new_n2130), .B(new_n478), .Y(new_n2131));
  nor_5      g1746(.A(new_n2131), .B(new_n2092), .Y(new_n2132));
  nand_5 g1747(.A(new_n2132), .B(new_n2132), .Y(new_n2133));
  and_6      g1748(.A(new_n2133), .B(new_n2101), .Y(new_n2134));
  nand_5 g1749(.A(new_n2134), .B(new_n2134), .Y(new_n2135));
  nand_5     g1750(.A(new_n1565), .B(new_n1411), .Y(new_n2136));
  nand_5 g1751(.A(new_n2136), .B(new_n2136), .Y(new_n2137));
  nand_5     g1752(.A(new_n2137), .B(new_n2135), .Y(new_n2138));
  nor_5      g1753(.A(new_n2138), .B(new_n2118), .Y(new_n2139));
  nand_5 g1754(.A(new_n2139), .B(new_n2139), .Y(new_n2140));
  nand_5     g1755(.A(new_n1422), .B(new_n1869), .Y(new_n2141));
  nand_5     g1756(.A(new_n1156), .B(new_n1036), .Y(new_n2142));
  nor_5      g1757(.A(new_n2142), .B(new_n2141), .Y(new_n2143));
  nand_5     g1758(.A(new_n2143), .B(new_n2140), .Y(new_n2144));
  nor_5      g1759(.A(new_n1836), .B(new_n1558), .Y(new_n2145));
  nor_5      g1760(.A(new_n2145), .B(new_n1827), .Y(new_n2146));
  nor_5      g1761(.A(new_n2146), .B(new_n1165), .Y(new_n2147));
  nor_5      g1762(.A(new_n1074), .B(new_n1033), .Y(new_n2148));
  nand_5 g1763(.A(new_n2148), .B(new_n2148), .Y(new_n2149));
  nor_5      g1764(.A(new_n2149), .B(new_n2147), .Y(new_n2150));
  nand_5     g1765(.A(new_n2150), .B(new_n2144), .Y(new_n2151));
  and_6      g1766(.A(new_n1075), .B(pi084), .Y(new_n2152));
  and_6      g1767(.A(new_n2152), .B(new_n2151), .Y(po008));
  nand_5 g1768(.A(new_n1161), .B(new_n1161), .Y(new_n2154));
  nor_5      g1769(.A(new_n2109), .B(new_n2088), .Y(new_n2155));
  nand_5 g1770(.A(new_n2155), .B(new_n2155), .Y(new_n2156));
  nand_5 g1771(.A(new_n1009), .B(new_n1009), .Y(new_n2157));
  nand_5     g1772(.A(new_n1770), .B(new_n1655), .Y(new_n2158));
  nand_5     g1773(.A(new_n2158), .B(new_n1745), .Y(new_n2159));
  nand_5     g1774(.A(new_n2159), .B(new_n2157), .Y(new_n2160));
  nor_5      g1775(.A(new_n2160), .B(new_n2075), .Y(new_n2161));
  nand_5 g1776(.A(new_n2161), .B(new_n2161), .Y(new_n2162));
  nand_5     g1777(.A(new_n2162), .B(new_n2156), .Y(new_n2163));
  nand_5     g1778(.A(new_n522), .B(new_n561), .Y(new_n2164));
  nor_5      g1779(.A(new_n2164), .B(new_n1497), .Y(new_n2165));
  nand_5     g1780(.A(new_n2165), .B(new_n2102), .Y(new_n2166));
  nand_5 g1781(.A(new_n2166), .B(new_n2166), .Y(new_n2167));
  nand_5     g1782(.A(new_n2167), .B(new_n2163), .Y(new_n2168));
  nand_5     g1783(.A(new_n1645), .B(new_n1386), .Y(new_n2169));
  nand_5 g1784(.A(new_n2169), .B(new_n2169), .Y(new_n2170));
  nand_5     g1785(.A(new_n2170), .B(new_n1818), .Y(new_n2171));
  nand_5     g1786(.A(new_n2171), .B(new_n1733), .Y(new_n2172));
  nand_5     g1787(.A(new_n974), .B(new_n669), .Y(new_n2173));
  nor_5      g1788(.A(new_n2173), .B(new_n1711), .Y(new_n2174));
  nand_5     g1789(.A(new_n2174), .B(new_n892), .Y(new_n2175));
  nand_5 g1790(.A(new_n2175), .B(new_n2175), .Y(new_n2176));
  nand_5     g1791(.A(new_n2176), .B(new_n2172), .Y(new_n2177));
  nand_5     g1792(.A(new_n1773), .B(new_n1738), .Y(new_n2178));
  nand_5 g1793(.A(new_n2178), .B(new_n2178), .Y(new_n2179));
  nand_5     g1794(.A(new_n2179), .B(new_n2177), .Y(new_n2180));
  nand_5 g1795(.A(new_n1195), .B(new_n1195), .Y(new_n2181));
  nand_5     g1796(.A(new_n2181), .B(new_n1177), .Y(new_n2182));
  nand_5 g1797(.A(new_n705), .B(new_n705), .Y(new_n2183));
  nand_5     g1798(.A(new_n1742), .B(new_n1789), .Y(new_n2184));
  nor_5      g1799(.A(new_n2184), .B(new_n2183), .Y(new_n2185));
  nand_5     g1800(.A(new_n2185), .B(new_n2182), .Y(new_n2186));
  nor_5      g1801(.A(new_n2186), .B(new_n2180), .Y(new_n2187));
  nor_5      g1802(.A(new_n2187), .B(new_n2168), .Y(new_n2188));
  nand_5 g1803(.A(pi226), .B(pi226), .Y(new_n2189));
  nand_5     g1804(.A(new_n1910), .B(new_n1903), .Y(new_n2190));
  nand_5     g1805(.A(new_n2190), .B(new_n1886), .Y(new_n2191));
  nand_5     g1806(.A(new_n2191), .B(new_n393), .Y(new_n2192));
  nand_5     g1807(.A(new_n2192), .B(new_n2189), .Y(new_n2193));
  nand_5 g1808(.A(new_n1915), .B(new_n1915), .Y(new_n2194));
  nor_5      g1809(.A(new_n1895), .B(pi207), .Y(new_n2195));
  nor_5      g1810(.A(new_n431), .B(pi126), .Y(new_n2196));
  nand_5 g1811(.A(new_n2196), .B(new_n2196), .Y(new_n2197));
  nand_5     g1812(.A(new_n2197), .B(new_n2195), .Y(new_n2198));
  nand_5     g1813(.A(new_n2198), .B(new_n2194), .Y(new_n2199));
  nor_5      g1814(.A(new_n2199), .B(new_n2193), .Y(new_n2200));
  nand_5 g1815(.A(new_n2200), .B(new_n2200), .Y(new_n2201));
  nand_5     g1816(.A(new_n413), .B(pi171), .Y(new_n2202));
  nand_5     g1817(.A(new_n2202), .B(new_n1329), .Y(new_n2203));
  nor_5      g1818(.A(new_n2203), .B(new_n1486), .Y(new_n2204));
  nand_5     g1819(.A(new_n445), .B(new_n447), .Y(new_n2205));
  nand_5 g1820(.A(new_n2205), .B(new_n2205), .Y(new_n2206));
  nand_5     g1821(.A(new_n2206), .B(new_n2204), .Y(new_n2207));
  nor_5      g1822(.A(new_n2207), .B(new_n2201), .Y(new_n2208));
  nand_5 g1823(.A(new_n565), .B(new_n565), .Y(new_n2209));
  nand_5     g1824(.A(new_n571), .B(new_n2209), .Y(new_n2210));
  nand_5     g1825(.A(new_n2210), .B(new_n1468), .Y(new_n2211));
  nand_5     g1826(.A(new_n2211), .B(new_n435), .Y(new_n2212));
  nand_5     g1827(.A(new_n1496), .B(new_n486), .Y(new_n2213));
  nand_5 g1828(.A(new_n2213), .B(new_n2213), .Y(new_n2214));
  nand_5     g1829(.A(new_n2214), .B(new_n529), .Y(new_n2215));
  nand_5     g1830(.A(new_n2215), .B(new_n1937), .Y(new_n2216));
  nand_5     g1831(.A(new_n2216), .B(new_n2212), .Y(new_n2217));
  nand_5 g1832(.A(new_n2217), .B(new_n2217), .Y(new_n2218));
  nand_5     g1833(.A(new_n2218), .B(new_n2208), .Y(new_n2219));
  nand_5 g1834(.A(pi240), .B(pi240), .Y(new_n2220));
  nand_5     g1835(.A(new_n2220), .B(pi147), .Y(new_n2221));
  nand_5     g1836(.A(new_n2221), .B(new_n1013), .Y(new_n2222));
  nor_5      g1837(.A(new_n2222), .B(new_n1759), .Y(new_n2223));
  nand_5 g1838(.A(new_n2223), .B(new_n2223), .Y(new_n2224));
  nand_5     g1839(.A(new_n2070), .B(new_n2220), .Y(new_n2225));
  nand_5 g1840(.A(new_n2225), .B(new_n2225), .Y(new_n2226));
  nand_5     g1841(.A(new_n2226), .B(new_n1769), .Y(new_n2227));
  nand_5     g1842(.A(new_n516), .B(new_n517), .Y(new_n2228));
  nand_5 g1843(.A(new_n2228), .B(new_n2228), .Y(new_n2229));
  nand_5     g1844(.A(new_n2229), .B(new_n2227), .Y(new_n2230));
  nor_5      g1845(.A(new_n2230), .B(new_n2224), .Y(new_n2231));
  nand_5 g1846(.A(new_n2231), .B(new_n2231), .Y(new_n2232));
  nor_5      g1847(.A(new_n2232), .B(new_n2219), .Y(new_n2233));
  nand_5     g1848(.A(new_n2233), .B(new_n2188), .Y(new_n2234));
  nor_5      g1849(.A(new_n697), .B(new_n500), .Y(new_n2235));
  nand_5     g1850(.A(new_n1792), .B(new_n1751), .Y(new_n2236));
  nor_5      g1851(.A(new_n2236), .B(new_n2235), .Y(new_n2237));
  nor_5      g1852(.A(new_n2237), .B(new_n2079), .Y(new_n2238));
  nor_5      g1853(.A(new_n2238), .B(new_n2166), .Y(new_n2239));
  nand_5     g1854(.A(new_n2123), .B(new_n1945), .Y(new_n2240));
  nand_5     g1855(.A(new_n2126), .B(new_n2105), .Y(new_n2241));
  nand_5     g1856(.A(new_n2241), .B(new_n2240), .Y(new_n2242));
  nand_5     g1857(.A(new_n2081), .B(new_n541), .Y(new_n2243));
  nand_5 g1858(.A(new_n2243), .B(new_n2243), .Y(new_n2244));
  nor_5      g1859(.A(new_n2244), .B(new_n2166), .Y(new_n2245));
  nor_5      g1860(.A(new_n2245), .B(new_n1906), .Y(new_n2246));
  nand_5     g1861(.A(new_n2246), .B(new_n2242), .Y(new_n2247));
  nor_5      g1862(.A(new_n2247), .B(new_n2239), .Y(new_n2248));
  nor_5      g1863(.A(new_n2248), .B(new_n2219), .Y(new_n2249));
  nand_5 g1864(.A(new_n2203), .B(new_n2203), .Y(new_n2250));
  nand_5 g1865(.A(pi128), .B(pi128), .Y(new_n2251));
  nand_5     g1866(.A(new_n1903), .B(new_n2251), .Y(new_n2252));
  nor_5      g1867(.A(new_n2252), .B(new_n1917), .Y(new_n2253));
  nor_5      g1868(.A(new_n2253), .B(new_n2193), .Y(new_n2254));
  nand_5     g1869(.A(new_n2189), .B(pi094), .Y(new_n2255));
  nand_5     g1870(.A(new_n2255), .B(new_n390), .Y(new_n2256));
  nor_5      g1871(.A(new_n2256), .B(new_n1325), .Y(new_n2257));
  nand_5 g1872(.A(new_n2257), .B(new_n2257), .Y(new_n2258));
  nor_5      g1873(.A(new_n2258), .B(new_n2254), .Y(new_n2259));
  nand_5     g1874(.A(new_n447), .B(pi156), .Y(new_n2260));
  and_6      g1875(.A(new_n2260), .B(new_n427), .Y(new_n2261));
  nand_5     g1876(.A(new_n2261), .B(new_n2195), .Y(new_n2262));
  nand_5     g1877(.A(new_n2262), .B(new_n2200), .Y(new_n2263));
  nand_5     g1878(.A(new_n2263), .B(new_n2259), .Y(new_n2264));
  nand_5     g1879(.A(new_n2264), .B(new_n2250), .Y(new_n2265));
  nand_5     g1880(.A(new_n2265), .B(new_n422), .Y(new_n2266));
  nand_5     g1881(.A(new_n2266), .B(new_n1986), .Y(new_n2267));
  nand_5 g1882(.A(new_n2267), .B(new_n2267), .Y(new_n2268));
  nor_5      g1883(.A(new_n2268), .B(new_n2249), .Y(new_n2269));
  nor_5      g1884(.A(new_n1424), .B(new_n1414), .Y(new_n2270));
  nand_5     g1885(.A(new_n2270), .B(new_n2269), .Y(new_n2271));
  nand_5 g1886(.A(new_n2271), .B(new_n2271), .Y(new_n2272));
  nand_5     g1887(.A(new_n2272), .B(new_n2234), .Y(new_n2273));
  nand_5 g1888(.A(new_n1854), .B(new_n1854), .Y(new_n2274));
  nand_5 g1889(.A(new_n1125), .B(new_n1125), .Y(new_n2275));
  nand_5     g1890(.A(new_n1805), .B(new_n806), .Y(new_n2276));
  nand_5     g1891(.A(new_n2276), .B(new_n2275), .Y(new_n2277));
  nand_5     g1892(.A(new_n2277), .B(new_n2274), .Y(new_n2278));
  nand_5     g1893(.A(new_n862), .B(new_n875), .Y(new_n2279));
  nand_5 g1894(.A(new_n2279), .B(new_n2279), .Y(new_n2280));
  nand_5     g1895(.A(new_n2280), .B(new_n2278), .Y(new_n2281));
  nand_5     g1896(.A(new_n2281), .B(new_n1133), .Y(new_n2282));
  nor_5      g1897(.A(new_n909), .B(new_n852), .Y(new_n2283));
  nand_5     g1898(.A(new_n2283), .B(new_n2176), .Y(new_n2284));
  nand_5 g1899(.A(new_n2284), .B(new_n2284), .Y(new_n2285));
  nand_5     g1900(.A(new_n2285), .B(new_n2233), .Y(new_n2286));
  nor_5      g1901(.A(new_n2286), .B(new_n2282), .Y(new_n2287));
  nor_5      g1902(.A(new_n2287), .B(new_n2273), .Y(new_n2288));
  nor_5      g1903(.A(new_n2288), .B(new_n1435), .Y(new_n2289));
  nor_5      g1904(.A(new_n2289), .B(new_n2154), .Y(new_n2290));
  nand_5     g1905(.A(new_n1148), .B(pi080), .Y(new_n2291));
  nor_5      g1906(.A(new_n2291), .B(new_n2290), .Y(po009));
  nand_5 g1907(.A(new_n1836), .B(new_n1836), .Y(new_n2293));
  nand_5     g1908(.A(new_n2137), .B(new_n2100), .Y(new_n2294));
  nand_5     g1909(.A(new_n2294), .B(new_n1422), .Y(new_n2295));
  nor_5      g1910(.A(new_n2295), .B(new_n1270), .Y(new_n2296));
  nand_5 g1911(.A(new_n921), .B(new_n921), .Y(new_n2297));
  nand_5     g1912(.A(new_n539), .B(new_n532), .Y(new_n2298));
  nand_5     g1913(.A(new_n2298), .B(new_n2214), .Y(new_n2299));
  nand_5     g1914(.A(new_n1927), .B(new_n565), .Y(new_n2300));
  nor_5      g1915(.A(new_n2300), .B(new_n2299), .Y(new_n2301));
  and_6      g1916(.A(new_n2301), .B(new_n1757), .Y(new_n2302));
  nor_5      g1917(.A(new_n1970), .B(new_n1800), .Y(new_n2303));
  nand_5 g1918(.A(new_n2303), .B(new_n2303), .Y(new_n2304));
  nand_5     g1919(.A(new_n2304), .B(new_n2301), .Y(new_n2305));
  nand_5 g1920(.A(new_n1937), .B(new_n1937), .Y(new_n2306));
  nand_5     g1921(.A(new_n2212), .B(new_n2306), .Y(new_n2307));
  nand_5     g1922(.A(new_n2307), .B(new_n551), .Y(new_n2308));
  nand_5 g1923(.A(new_n2308), .B(new_n2308), .Y(new_n2309));
  nand_5     g1924(.A(new_n2251), .B(new_n391), .Y(new_n2310));
  nor_5      g1925(.A(new_n2310), .B(new_n389), .Y(new_n2311));
  nand_5     g1926(.A(new_n2311), .B(new_n1896), .Y(new_n2312));
  nor_5      g1927(.A(new_n2312), .B(new_n1906), .Y(new_n2313));
  nand_5     g1928(.A(new_n2313), .B(new_n2309), .Y(new_n2314));
  nand_5 g1929(.A(new_n2314), .B(new_n2314), .Y(new_n2315));
  nand_5     g1930(.A(new_n2315), .B(new_n2305), .Y(new_n2316));
  nor_5      g1931(.A(new_n2316), .B(new_n2302), .Y(new_n2317));
  nand_5     g1932(.A(new_n1471), .B(new_n553), .Y(new_n2318));
  nand_5 g1933(.A(new_n445), .B(new_n445), .Y(new_n2319));
  nand_5     g1934(.A(new_n551), .B(new_n2319), .Y(new_n2320));
  nand_5 g1935(.A(new_n2320), .B(new_n2320), .Y(new_n2321));
  nor_5      g1936(.A(new_n2321), .B(new_n1893), .Y(new_n2322));
  nand_5     g1937(.A(new_n2322), .B(new_n2318), .Y(new_n2323));
  nand_5     g1938(.A(new_n2323), .B(new_n1896), .Y(new_n2324));
  nand_5     g1939(.A(new_n2324), .B(new_n462), .Y(new_n2325));
  nor_5      g1940(.A(new_n1904), .B(new_n470), .Y(new_n2326));
  nand_5     g1941(.A(new_n2326), .B(new_n2325), .Y(new_n2327));
  nand_5     g1942(.A(new_n2327), .B(new_n1994), .Y(new_n2328));
  nor_5      g1943(.A(new_n2328), .B(new_n2317), .Y(new_n2329));
  nor_5      g1944(.A(new_n2329), .B(new_n1981), .Y(new_n2330));
  nand_5 g1945(.A(new_n2330), .B(new_n2330), .Y(new_n2331));
  nand_5     g1946(.A(new_n2161), .B(new_n1737), .Y(new_n2332));
  nor_5      g1947(.A(new_n2332), .B(new_n1830), .Y(new_n2333));
  nand_5     g1948(.A(new_n2333), .B(new_n2331), .Y(new_n2334));
  nor_5      g1949(.A(new_n2334), .B(new_n2297), .Y(new_n2335));
  nand_5 g1950(.A(new_n2335), .B(new_n2335), .Y(new_n2336));
  nand_5     g1951(.A(new_n2336), .B(new_n2139), .Y(new_n2337));
  nand_5     g1952(.A(new_n2337), .B(new_n2296), .Y(new_n2338));
  nand_5     g1953(.A(new_n2338), .B(new_n1558), .Y(new_n2339));
  nand_5     g1954(.A(new_n2339), .B(new_n2293), .Y(new_n2340));
  nor_5      g1955(.A(new_n1068), .B(new_n1054), .Y(new_n2341));
  nand_5     g1956(.A(new_n2341), .B(new_n2340), .Y(new_n2342));
  nand_5 g1957(.A(new_n2342), .B(new_n2342), .Y(new_n2343));
  nand_5     g1958(.A(pi157), .B(new_n1052), .Y(new_n2344));
  nand_5     g1959(.A(new_n2344), .B(pi233), .Y(new_n2345));
  nor_5      g1960(.A(new_n2345), .B(new_n2343), .Y(po010));
  nor_5      g1961(.A(new_n2269), .B(new_n1318), .Y(new_n2347));
  nand_5 g1962(.A(new_n2186), .B(new_n2186), .Y(new_n2348));
  nand_5 g1963(.A(new_n1507), .B(new_n1507), .Y(new_n2349));
  nand_5     g1964(.A(new_n1990), .B(new_n2349), .Y(new_n2350));
  nand_5     g1965(.A(new_n1429), .B(new_n1161), .Y(new_n2351));
  nand_5     g1966(.A(new_n2351), .B(new_n1985), .Y(new_n2352));
  nand_5 g1967(.A(new_n1092), .B(new_n1092), .Y(new_n2353));
  nand_5 g1968(.A(new_n884), .B(new_n884), .Y(new_n2354));
  nand_5     g1969(.A(new_n2354), .B(new_n819), .Y(new_n2355));
  nor_5      g1970(.A(new_n2355), .B(new_n2353), .Y(new_n2356));
  nand_5     g1971(.A(new_n2356), .B(new_n2352), .Y(new_n2357));
  nand_5 g1972(.A(new_n2357), .B(new_n2357), .Y(new_n2358));
  nand_5     g1973(.A(new_n2358), .B(new_n2350), .Y(new_n2359));
  nand_5 g1974(.A(new_n867), .B(new_n867), .Y(new_n2360));
  nand_5 g1975(.A(new_n802), .B(new_n802), .Y(new_n2361));
  nor_5      g1976(.A(new_n1082), .B(new_n2361), .Y(new_n2362));
  nor_5      g1977(.A(new_n2362), .B(new_n2355), .Y(new_n2363));
  nor_5      g1978(.A(new_n2363), .B(new_n2360), .Y(new_n2364));
  nand_5     g1979(.A(new_n1175), .B(new_n1182), .Y(new_n2365));
  nand_5 g1980(.A(new_n2365), .B(new_n2365), .Y(new_n2366));
  nand_5     g1981(.A(new_n2366), .B(new_n2364), .Y(new_n2367));
  nand_5 g1982(.A(new_n2367), .B(new_n2367), .Y(new_n2368));
  nand_5     g1983(.A(new_n2368), .B(new_n2359), .Y(new_n2369));
  nand_5     g1984(.A(new_n2369), .B(new_n2348), .Y(new_n2370));
  nand_5 g1985(.A(new_n1790), .B(new_n1790), .Y(new_n2371));
  nand_5     g1986(.A(new_n2371), .B(new_n1003), .Y(new_n2372));
  nor_5      g1987(.A(new_n2236), .B(new_n505), .Y(new_n2373));
  nand_5     g1988(.A(new_n2373), .B(new_n2372), .Y(new_n2374));
  nand_5 g1989(.A(new_n2374), .B(new_n2374), .Y(new_n2375));
  nand_5     g1990(.A(new_n2375), .B(new_n2370), .Y(new_n2376));
  nand_5     g1991(.A(new_n2233), .B(new_n1317), .Y(new_n2377));
  nor_5      g1992(.A(new_n2377), .B(new_n2376), .Y(new_n2378));
  nor_5      g1993(.A(new_n2378), .B(new_n2347), .Y(new_n2379));
  nor_5      g1994(.A(new_n2379), .B(new_n1487), .Y(po011));
  nand_5 g1995(.A(new_n1747), .B(new_n1747), .Y(new_n2381));
  nor_5      g1996(.A(new_n1578), .B(new_n1562), .Y(new_n2382));
  nor_5      g1997(.A(new_n2382), .B(new_n1838), .Y(new_n2383));
  nand_5 g1998(.A(new_n2191), .B(new_n2191), .Y(new_n2384));
  nand_5     g1999(.A(new_n1905), .B(pi016), .Y(new_n2385));
  nand_5     g2000(.A(new_n2385), .B(new_n2384), .Y(new_n2386));
  nand_5 g2001(.A(new_n2386), .B(new_n2386), .Y(new_n2387));
  nand_5     g2002(.A(new_n2387), .B(new_n1881), .Y(new_n2388));
  nand_5 g2003(.A(new_n2388), .B(new_n2388), .Y(new_n2389));
  nand_5     g2004(.A(new_n2389), .B(new_n2240), .Y(new_n2390));
  nor_5      g2005(.A(new_n2390), .B(new_n2325), .Y(new_n2391));
  nand_5     g2006(.A(new_n2391), .B(new_n2383), .Y(new_n2392));
  nor_5      g2007(.A(new_n2392), .B(new_n2103), .Y(new_n2393));
  nand_5     g2008(.A(new_n2393), .B(new_n2161), .Y(new_n2394));
  nand_5 g2009(.A(new_n2394), .B(new_n2394), .Y(new_n2395));
  nand_5     g2010(.A(new_n2395), .B(new_n2381), .Y(new_n2396));
  nand_5     g2011(.A(new_n2244), .B(new_n2156), .Y(new_n2397));
  nand_5     g2012(.A(new_n2397), .B(new_n2393), .Y(new_n2398));
  nand_5 g2013(.A(new_n2241), .B(new_n2241), .Y(new_n2399));
  nor_5      g2014(.A(new_n2392), .B(new_n2399), .Y(new_n2400));
  nand_5 g2015(.A(new_n2193), .B(new_n2193), .Y(new_n2401));
  nand_5     g2016(.A(new_n2401), .B(new_n1456), .Y(new_n2402));
  nand_5     g2017(.A(new_n2402), .B(new_n2259), .Y(new_n2403));
  nand_5     g2018(.A(new_n2403), .B(new_n2204), .Y(new_n2404));
  nand_5     g2019(.A(new_n2404), .B(new_n1585), .Y(new_n2405));
  nand_5     g2020(.A(new_n2405), .B(new_n2383), .Y(new_n2406));
  nand_5 g2021(.A(new_n2406), .B(new_n2406), .Y(new_n2407));
  nor_5      g2022(.A(new_n2407), .B(new_n1831), .Y(new_n2408));
  nand_5 g2023(.A(new_n2408), .B(new_n2408), .Y(new_n2409));
  nor_5      g2024(.A(new_n2409), .B(new_n2400), .Y(new_n2410));
  nand_5     g2025(.A(new_n2410), .B(new_n2398), .Y(new_n2411));
  nor_5      g2026(.A(new_n2411), .B(new_n1820), .Y(new_n2412));
  nand_5     g2027(.A(new_n2412), .B(new_n2396), .Y(new_n2413));
  nand_5     g2028(.A(new_n1860), .B(new_n1847), .Y(new_n2414));
  nor_5      g2029(.A(new_n2414), .B(new_n1858), .Y(new_n2415));
  nand_5     g2030(.A(new_n2415), .B(new_n2413), .Y(new_n2416));
  nand_5     g2031(.A(new_n2416), .B(new_n1733), .Y(new_n2417));
  and_6      g2032(.A(new_n609), .B(pi108), .Y(new_n2418));
  nand_5     g2033(.A(new_n2418), .B(new_n2417), .Y(new_n2419));
  nand_5 g2034(.A(new_n2419), .B(new_n2419), .Y(po012));
  nand_5 g2035(.A(new_n2129), .B(new_n2129), .Y(new_n2421));
  nor_5      g2036(.A(new_n2421), .B(new_n1977), .Y(new_n2422));
  nand_5     g2037(.A(new_n1350), .B(new_n481), .Y(new_n2423));
  nor_5      g2038(.A(new_n2423), .B(new_n575), .Y(new_n2424));
  nand_5 g2039(.A(new_n2424), .B(new_n2424), .Y(new_n2425));
  nand_5 g2040(.A(new_n1882), .B(new_n1882), .Y(new_n2426));
  nor_5      g2041(.A(new_n2426), .B(pi117), .Y(new_n2427));
  nand_5     g2042(.A(new_n2427), .B(new_n2425), .Y(new_n2428));
  nor_5      g2043(.A(new_n2428), .B(new_n2422), .Y(new_n2429));
  nor_5      g2044(.A(new_n2429), .B(new_n1926), .Y(new_n2430));
  nor_5      g2045(.A(new_n2430), .B(new_n1566), .Y(new_n2431));
  nand_5     g2046(.A(new_n1569), .B(pi218), .Y(new_n2432));
  nor_5      g2047(.A(new_n2432), .B(new_n2431), .Y(po013));
  nand_5 g2048(.A(new_n960), .B(new_n960), .Y(new_n2434));
  nand_5     g2049(.A(new_n643), .B(new_n633), .Y(new_n2435));
  nand_5     g2050(.A(new_n2435), .B(new_n2017), .Y(new_n2436));
  nand_5     g2051(.A(new_n2436), .B(new_n1441), .Y(new_n2437));
  nand_5     g2052(.A(new_n2437), .B(new_n1502), .Y(new_n2438));
  nand_5 g2053(.A(new_n2438), .B(new_n2438), .Y(new_n2439));
  nand_5     g2054(.A(new_n1137), .B(new_n944), .Y(new_n2440));
  nand_5     g2055(.A(new_n2440), .B(new_n1398), .Y(new_n2441));
  nand_5 g2056(.A(new_n2441), .B(new_n2441), .Y(new_n2442));
  nor_5      g2057(.A(new_n2442), .B(new_n942), .Y(new_n2443));
  nor_5      g2058(.A(new_n2443), .B(new_n1393), .Y(new_n2444));
  nand_5 g2059(.A(new_n2444), .B(new_n2444), .Y(new_n2445));
  nand_5     g2060(.A(new_n2445), .B(new_n709), .Y(new_n2446));
  nand_5     g2061(.A(new_n2446), .B(new_n2439), .Y(new_n2447));
  nand_5     g2062(.A(new_n2447), .B(new_n1521), .Y(new_n2448));
  nand_5     g2063(.A(new_n2448), .B(new_n1556), .Y(new_n2449));
  nand_5     g2064(.A(new_n2449), .B(new_n2434), .Y(new_n2450));
  nand_5     g2065(.A(new_n2450), .B(new_n947), .Y(new_n2451));
  nor_5      g2066(.A(new_n2451), .B(new_n945), .Y(po014));
  nand_5 g2067(.A(new_n2247), .B(new_n2247), .Y(new_n2453));
  nand_5 g2068(.A(new_n2168), .B(new_n2168), .Y(new_n2454));
  nand_5     g2069(.A(new_n2049), .B(new_n1381), .Y(new_n2455));
  nand_5     g2070(.A(new_n599), .B(new_n578), .Y(new_n2456));
  nor_5      g2071(.A(new_n2456), .B(new_n2169), .Y(new_n2457));
  nand_5     g2072(.A(new_n2457), .B(new_n2455), .Y(new_n2458));
  nand_5 g2073(.A(new_n2458), .B(new_n2458), .Y(new_n2459));
  nand_5     g2074(.A(new_n1958), .B(new_n1258), .Y(new_n2460));
  nand_5     g2075(.A(new_n2460), .B(new_n2034), .Y(new_n2461));
  nor_5      g2076(.A(new_n2461), .B(new_n2035), .Y(new_n2462));
  nand_5     g2077(.A(new_n2462), .B(new_n2459), .Y(new_n2463));
  nand_5 g2078(.A(new_n2463), .B(new_n2463), .Y(new_n2464));
  nand_5     g2079(.A(new_n2464), .B(new_n1961), .Y(new_n2465));
  nand_5     g2080(.A(new_n2034), .B(new_n1101), .Y(new_n2466));
  nand_5     g2081(.A(new_n2466), .B(new_n1220), .Y(new_n2467));
  nor_5      g2082(.A(new_n2467), .B(new_n1670), .Y(new_n2468));
  nand_5     g2083(.A(new_n2468), .B(new_n1389), .Y(new_n2469));
  nand_5     g2084(.A(new_n2469), .B(new_n2459), .Y(new_n2470));
  nand_5     g2085(.A(new_n1645), .B(pi195), .Y(new_n2471));
  nand_5     g2086(.A(new_n2471), .B(new_n1639), .Y(new_n2472));
  nand_5     g2087(.A(new_n2472), .B(new_n1737), .Y(new_n2473));
  nand_5     g2088(.A(new_n2473), .B(new_n1747), .Y(new_n2474));
  nand_5 g2089(.A(new_n2474), .B(new_n2474), .Y(new_n2475));
  nor_5      g2090(.A(new_n2085), .B(new_n704), .Y(new_n2476));
  nand_5     g2091(.A(new_n2476), .B(new_n2475), .Y(new_n2477));
  nand_5 g2092(.A(new_n2477), .B(new_n2477), .Y(new_n2478));
  nand_5     g2093(.A(new_n2478), .B(new_n2470), .Y(new_n2479));
  nand_5 g2094(.A(new_n2479), .B(new_n2479), .Y(new_n2480));
  nand_5     g2095(.A(new_n2480), .B(new_n2465), .Y(new_n2481));
  nand_5 g2096(.A(new_n2481), .B(new_n2481), .Y(new_n2482));
  nor_5      g2097(.A(new_n1344), .B(new_n424), .Y(new_n2483));
  nand_5 g2098(.A(new_n2483), .B(new_n2483), .Y(new_n2484));
  nor_5      g2099(.A(new_n2484), .B(new_n1682), .Y(new_n2485));
  nand_5     g2100(.A(new_n2485), .B(new_n2464), .Y(new_n2486));
  nand_5     g2101(.A(new_n2486), .B(new_n2482), .Y(new_n2487));
  nand_5     g2102(.A(new_n2487), .B(new_n2454), .Y(new_n2488));
  nand_5     g2103(.A(new_n2488), .B(new_n2453), .Y(new_n2489));
  nand_5     g2104(.A(new_n2387), .B(new_n2327), .Y(new_n2490));
  nand_5 g2105(.A(new_n2490), .B(new_n2490), .Y(new_n2491));
  nand_5     g2106(.A(new_n2491), .B(new_n2489), .Y(new_n2492));
  nand_5 g2107(.A(new_n2492), .B(new_n2492), .Y(new_n2493));
  nor_5      g2108(.A(new_n2493), .B(new_n2426), .Y(new_n2494));
  nand_5     g2109(.A(new_n1879), .B(pi022), .Y(new_n2495));
  nor_5      g2110(.A(new_n2495), .B(new_n2494), .Y(po015));
  nand_5     g2111(.A(new_n1806), .B(new_n1128), .Y(new_n2497));
  nand_5     g2112(.A(new_n2497), .B(new_n1857), .Y(new_n2498));
  nand_5 g2113(.A(new_n2498), .B(new_n2498), .Y(new_n2499));
  nand_5 g2114(.A(new_n1721), .B(new_n1721), .Y(new_n2500));
  nand_5 g2115(.A(new_n2188), .B(new_n2188), .Y(new_n2501));
  nand_5     g2116(.A(new_n2501), .B(new_n1695), .Y(new_n2502));
  nand_5     g2117(.A(new_n2502), .B(new_n2500), .Y(new_n2503));
  nand_5     g2118(.A(new_n2503), .B(new_n1128), .Y(new_n2504));
  nand_5     g2119(.A(new_n2504), .B(new_n2499), .Y(new_n2505));
  nor_5      g2120(.A(new_n2505), .B(new_n830), .Y(new_n2506));
  nor_5      g2121(.A(new_n2506), .B(pi135), .Y(new_n2507));
  nor_5      g2122(.A(new_n2507), .B(new_n727), .Y(po016));
  nand_5 g2123(.A(new_n1477), .B(new_n1477), .Y(new_n2509));
  nand_5     g2124(.A(new_n2407), .B(new_n1855), .Y(new_n2510));
  nand_5     g2125(.A(new_n2510), .B(new_n2282), .Y(new_n2511));
  nand_5     g2126(.A(new_n2511), .B(new_n2285), .Y(new_n2512));
  nand_5     g2127(.A(new_n2512), .B(new_n2187), .Y(new_n2513));
  nand_5     g2128(.A(new_n2513), .B(new_n2454), .Y(new_n2514));
  nand_5     g2129(.A(new_n2514), .B(new_n1975), .Y(new_n2515));
  nand_5     g2130(.A(new_n2515), .B(new_n2509), .Y(new_n2516));
  nand_5     g2131(.A(new_n2516), .B(new_n437), .Y(new_n2517));
  nand_5     g2132(.A(new_n2517), .B(new_n1463), .Y(new_n2518));
  nor_5      g2133(.A(new_n2518), .B(pi159), .Y(new_n2519));
  nor_5      g2134(.A(new_n2519), .B(pi098), .Y(new_n2520));
  nor_5      g2135(.A(new_n2520), .B(new_n448), .Y(po017));
  nand_5     g2136(.A(new_n2492), .B(new_n397), .Y(new_n2522));
  nand_5     g2137(.A(new_n2522), .B(new_n1484), .Y(new_n2523));
  nor_5      g2138(.A(new_n2523), .B(pi081), .Y(new_n2524));
  nor_5      g2139(.A(new_n2524), .B(pi103), .Y(new_n2525));
  nor_5      g2140(.A(new_n2525), .B(new_n1321), .Y(po018));
  nand_5 g2141(.A(new_n1779), .B(new_n1779), .Y(new_n2527));
  nand_5 g2142(.A(new_n2238), .B(new_n2238), .Y(new_n2528));
  nand_5     g2143(.A(new_n2167), .B(new_n1932), .Y(new_n2529));
  nor_5      g2144(.A(new_n2529), .B(new_n1863), .Y(new_n2530));
  nand_5     g2145(.A(new_n2530), .B(new_n2528), .Y(new_n2531));
  nand_5     g2146(.A(new_n2322), .B(new_n2308), .Y(new_n2532));
  nand_5 g2147(.A(new_n2313), .B(new_n2313), .Y(new_n2533));
  nor_5      g2148(.A(new_n2533), .B(new_n1982), .Y(new_n2534));
  nand_5     g2149(.A(new_n2534), .B(new_n2532), .Y(new_n2535));
  nor_5      g2150(.A(new_n2535), .B(new_n2424), .Y(new_n2536));
  nor_5      g2151(.A(new_n2536), .B(new_n1997), .Y(new_n2537));
  nor_5      g2152(.A(new_n2537), .B(new_n2357), .Y(new_n2538));
  nor_5      g2153(.A(new_n2538), .B(new_n2367), .Y(new_n2539));
  nor_5      g2154(.A(new_n2539), .B(new_n2180), .Y(new_n2540));
  nand_5     g2155(.A(new_n2540), .B(new_n2531), .Y(new_n2541));
  nand_5     g2156(.A(new_n2541), .B(new_n2527), .Y(new_n2542));
  nand_5     g2157(.A(new_n2542), .B(new_n2226), .Y(new_n2543));
  nand_5     g2158(.A(new_n2543), .B(new_n2221), .Y(new_n2544));
  nor_5      g2159(.A(new_n2544), .B(pi070), .Y(new_n2545));
  nor_5      g2160(.A(new_n2545), .B(pi074), .Y(new_n2546));
  nor_5      g2161(.A(new_n2546), .B(new_n688), .Y(po019));
  nand_5     g2162(.A(new_n1745), .B(new_n1661), .Y(new_n2548));
  nand_5     g2163(.A(new_n2074), .B(pi147), .Y(new_n2549));
  nand_5 g2164(.A(new_n2549), .B(new_n2549), .Y(new_n2550));
  nand_5     g2165(.A(new_n2550), .B(new_n2548), .Y(new_n2551));
  nand_5 g2166(.A(new_n2551), .B(new_n2551), .Y(po020));
  nand_5     g2167(.A(new_n2492), .B(new_n395), .Y(new_n2553));
  nor_5      g2168(.A(new_n2553), .B(pi200), .Y(new_n2554));
  nand_5     g2169(.A(new_n404), .B(pi171), .Y(new_n2555));
  nor_5      g2170(.A(new_n2555), .B(new_n2554), .Y(po021));
  nand_5 g2171(.A(pi070), .B(pi070), .Y(new_n2557));
  nor_5      g2172(.A(new_n2544), .B(new_n2557), .Y(po022));
  nand_5 g2173(.A(new_n2090), .B(new_n2090), .Y(new_n2559));
  nand_5 g2174(.A(new_n2066), .B(new_n2066), .Y(new_n2560));
  nor_5      g2175(.A(new_n2560), .B(new_n1636), .Y(new_n2561));
  nor_5      g2176(.A(new_n2561), .B(new_n2559), .Y(new_n2562));
  nand_5 g2177(.A(new_n2114), .B(new_n2114), .Y(new_n2563));
  nor_5      g2178(.A(new_n2563), .B(new_n1458), .Y(new_n2564));
  nand_5 g2179(.A(new_n2564), .B(new_n2564), .Y(new_n2565));
  nor_5      g2180(.A(new_n2565), .B(new_n2562), .Y(new_n2566));
  nor_5      g2181(.A(new_n2566), .B(new_n2316), .Y(new_n2567));
  nor_5      g2182(.A(new_n2567), .B(new_n2330), .Y(new_n2568));
  nor_5      g2183(.A(new_n2568), .B(new_n1325), .Y(new_n2569));
  nand_5     g2184(.A(pi022), .B(new_n411), .Y(new_n2570));
  nand_5     g2185(.A(new_n2570), .B(pi075), .Y(new_n2571));
  nor_5      g2186(.A(new_n2571), .B(new_n2569), .Y(po023));
  nand_5     g2187(.A(new_n1873), .B(new_n1025), .Y(new_n2573));
  nor_5      g2188(.A(new_n1539), .B(new_n1306), .Y(new_n2574));
  nand_5     g2189(.A(new_n2574), .B(new_n2573), .Y(new_n2575));
  nand_5     g2190(.A(new_n2575), .B(new_n1534), .Y(new_n2576));
  nor_5      g2191(.A(new_n2576), .B(pi170), .Y(new_n2577));
  nor_5      g2192(.A(new_n2577), .B(pi023), .Y(new_n2578));
  nor_5      g2193(.A(new_n2578), .B(new_n957), .Y(po024));
  nand_5 g2194(.A(new_n497), .B(new_n497), .Y(new_n2580));
  nor_5      g2195(.A(new_n2539), .B(new_n2186), .Y(new_n2581));
  nor_5      g2196(.A(new_n2581), .B(new_n2374), .Y(new_n2582));
  nor_5      g2197(.A(new_n2582), .B(new_n2580), .Y(new_n2583));
  nand_5     g2198(.A(new_n509), .B(pi066), .Y(new_n2584));
  nor_5      g2199(.A(new_n2584), .B(new_n2583), .Y(po025));
  nor_5      g2200(.A(new_n941), .B(new_n866), .Y(new_n2586));
  nor_5      g2201(.A(new_n2586), .B(new_n684), .Y(new_n2587));
  nand_5     g2202(.A(new_n1191), .B(new_n918), .Y(new_n2588));
  nand_5     g2203(.A(new_n2588), .B(new_n1714), .Y(new_n2589));
  nor_5      g2204(.A(new_n2589), .B(new_n2587), .Y(new_n2590));
  nor_5      g2205(.A(new_n2590), .B(new_n2021), .Y(new_n2591));
  nand_5     g2206(.A(new_n778), .B(new_n824), .Y(new_n2592));
  nor_5      g2207(.A(new_n2592), .B(new_n2589), .Y(new_n2593));
  nand_5     g2208(.A(new_n2593), .B(new_n2044), .Y(new_n2594));
  nand_5     g2209(.A(new_n2594), .B(new_n2591), .Y(new_n2595));
  nand_5     g2210(.A(new_n2595), .B(new_n2031), .Y(new_n2596));
  nand_5     g2211(.A(new_n2596), .B(new_n1878), .Y(new_n2597));
  nand_5     g2212(.A(new_n2597), .B(new_n2036), .Y(new_n2598));
  and_6      g2213(.A(new_n2598), .B(new_n1099), .Y(new_n2599));
  nand_5     g2214(.A(new_n1110), .B(pi053), .Y(new_n2600));
  nor_5      g2215(.A(new_n2600), .B(new_n2599), .Y(po026));
  nand_5     g2216(.A(new_n1398), .B(new_n1164), .Y(new_n2602));
  nand_5 g2217(.A(new_n2602), .B(new_n2602), .Y(new_n2603));
  nand_5 g2218(.A(new_n742), .B(new_n742), .Y(new_n2604));
  nand_5     g2219(.A(new_n2352), .B(new_n1989), .Y(new_n2605));
  nand_5     g2220(.A(new_n2605), .B(new_n1237), .Y(new_n2606));
  nor_5      g2221(.A(new_n2606), .B(new_n2604), .Y(new_n2607));
  nor_5      g2222(.A(new_n2607), .B(new_n2603), .Y(new_n2608));
  nand_5     g2223(.A(new_n753), .B(new_n735), .Y(new_n2609));
  nor_5      g2224(.A(new_n2609), .B(new_n2608), .Y(new_n2610));
  nand_5 g2225(.A(new_n800), .B(new_n800), .Y(new_n2611));
  nor_5      g2226(.A(new_n1878), .B(new_n2611), .Y(new_n2612));
  nand_5     g2227(.A(new_n2612), .B(new_n2610), .Y(new_n2613));
  nand_5     g2228(.A(new_n2613), .B(new_n937), .Y(new_n2614));
  nand_5     g2229(.A(new_n2614), .B(new_n2593), .Y(new_n2615));
  nand_5     g2230(.A(new_n2615), .B(new_n2591), .Y(new_n2616));
  nand_5 g2231(.A(new_n484), .B(new_n484), .Y(new_n2617));
  nor_5      g2232(.A(new_n2024), .B(new_n2617), .Y(new_n2618));
  nand_5     g2233(.A(new_n2618), .B(new_n2616), .Y(new_n2619));
  nor_5      g2234(.A(new_n2619), .B(pi251), .Y(new_n2620));
  nor_5      g2235(.A(new_n2620), .B(pi242), .Y(new_n2621));
  nor_5      g2236(.A(new_n2621), .B(pi125), .Y(new_n2622));
  nor_5      g2237(.A(new_n2622), .B(pi210), .Y(new_n2623));
  nor_5      g2238(.A(new_n2623), .B(new_n561), .Y(po027));
  nand_5     g2239(.A(new_n2281), .B(new_n1129), .Y(new_n2625));
  nor_5      g2240(.A(new_n2625), .B(new_n2286), .Y(new_n2626));
  nor_5      g2241(.A(new_n2626), .B(new_n2273), .Y(new_n2627));
  nor_5      g2242(.A(new_n2627), .B(new_n1438), .Y(new_n2628));
  nand_5     g2243(.A(new_n2602), .B(new_n931), .Y(new_n2629));
  nor_5      g2244(.A(new_n2629), .B(new_n2628), .Y(new_n2630));
  nand_5 g2245(.A(new_n2630), .B(new_n2630), .Y(new_n2631));
  nand_5     g2246(.A(new_n2631), .B(new_n1367), .Y(new_n2632));
  nand_5     g2247(.A(new_n2632), .B(new_n922), .Y(new_n2633));
  nand_5     g2248(.A(new_n2633), .B(new_n798), .Y(new_n2634));
  nand_5     g2249(.A(new_n2634), .B(new_n803), .Y(new_n2635));
  nand_5     g2250(.A(new_n2635), .B(new_n806), .Y(new_n2636));
  nor_5      g2251(.A(new_n2636), .B(new_n1600), .Y(po028));
  nand_5 g2252(.A(pi127), .B(pi127), .Y(new_n2638));
  nor_5      g2253(.A(new_n2012), .B(pi206), .Y(new_n2639));
  nor_5      g2254(.A(new_n2639), .B(pi018), .Y(new_n2640));
  nor_5      g2255(.A(new_n2640), .B(pi020), .Y(new_n2641));
  nor_5      g2256(.A(new_n2641), .B(pi212), .Y(new_n2642));
  nor_5      g2257(.A(new_n2642), .B(new_n2638), .Y(po029));
  nand_5     g2258(.A(new_n2543), .B(new_n1002), .Y(new_n2644));
  nand_5     g2259(.A(new_n2644), .B(new_n707), .Y(new_n2645));
  and_6      g2260(.A(new_n1016), .B(pi043), .Y(new_n2646));
  nand_5     g2261(.A(new_n2646), .B(new_n2645), .Y(new_n2647));
  nand_5 g2262(.A(new_n2647), .B(new_n2647), .Y(po030));
  nor_5      g2263(.A(new_n2576), .B(new_n1536), .Y(po031));
  nand_5     g2264(.A(new_n1521), .B(new_n1235), .Y(new_n2650));
  nand_5     g2265(.A(new_n2650), .B(new_n1706), .Y(new_n2651));
  nand_5     g2266(.A(new_n2651), .B(new_n1693), .Y(new_n2652));
  nand_5     g2267(.A(new_n2652), .B(new_n1675), .Y(new_n2653));
  nand_5     g2268(.A(new_n1615), .B(pi112), .Y(new_n2654));
  nor_5      g2269(.A(new_n2654), .B(new_n2653), .Y(po032));
  nand_5     g2270(.A(new_n2634), .B(new_n1606), .Y(new_n2656));
  nand_5     g2271(.A(new_n2656), .B(pi008), .Y(new_n2657));
  nand_5 g2272(.A(new_n2657), .B(new_n2657), .Y(po033));
  nand_5 g2273(.A(new_n2010), .B(new_n2010), .Y(new_n2659));
  nor_5      g2274(.A(new_n2659), .B(pi032), .Y(new_n2660));
  nor_5      g2275(.A(new_n2660), .B(new_n1572), .Y(po034));
  nand_5 g2276(.A(new_n2174), .B(new_n2174), .Y(new_n2662));
  nand_5     g2277(.A(new_n1930), .B(new_n1645), .Y(new_n2663));
  nor_5      g2278(.A(new_n2663), .B(new_n1870), .Y(new_n2664));
  nand_5     g2279(.A(new_n2664), .B(new_n1376), .Y(new_n2665));
  nor_5      g2280(.A(new_n2665), .B(new_n2662), .Y(new_n2666));
  nand_5     g2281(.A(new_n1992), .B(new_n1461), .Y(new_n2667));
  nor_5      g2282(.A(new_n2063), .B(new_n1867), .Y(new_n2668));
  and_6      g2283(.A(new_n2668), .B(new_n2165), .Y(new_n2669));
  nand_5 g2284(.A(pi244), .B(pi244), .Y(new_n2670));
  nor_5      g2285(.A(pi110), .B(pi055), .Y(new_n2671));
  nand_5     g2286(.A(new_n2671), .B(new_n2670), .Y(new_n2672));
  nor_5      g2287(.A(new_n769), .B(new_n715), .Y(new_n2673));
  nand_5     g2288(.A(new_n2673), .B(new_n753), .Y(new_n2674));
  nor_5      g2289(.A(new_n2674), .B(new_n2672), .Y(new_n2675));
  and_6      g2290(.A(new_n1491), .B(new_n1013), .Y(new_n2676));
  nand_5     g2291(.A(new_n2676), .B(new_n2675), .Y(new_n2677));
  nand_5     g2292(.A(new_n1688), .B(new_n1673), .Y(new_n2678));
  nor_5      g2293(.A(new_n2678), .B(new_n2677), .Y(new_n2679));
  nand_5     g2294(.A(new_n2679), .B(new_n2669), .Y(new_n2680));
  nor_5      g2295(.A(new_n2680), .B(new_n2667), .Y(new_n2681));
  nand_5     g2296(.A(new_n2681), .B(new_n2666), .Y(po035));
  nor_5      g2297(.A(new_n2582), .B(new_n2243), .Y(new_n2683));
  nand_5     g2298(.A(new_n2102), .B(pi041), .Y(new_n2684));
  nor_5      g2299(.A(new_n2684), .B(new_n2683), .Y(po036));
  nor_5      g2300(.A(new_n2480), .B(new_n2438), .Y(new_n2686));
  nor_5      g2301(.A(new_n2686), .B(new_n1520), .Y(new_n2687));
  nor_5      g2302(.A(new_n2687), .B(new_n1557), .Y(new_n2688));
  nor_5      g2303(.A(new_n2688), .B(new_n971), .Y(new_n2689));
  nand_5     g2304(.A(new_n1593), .B(pi052), .Y(new_n2690));
  nor_5      g2305(.A(new_n2690), .B(new_n2689), .Y(po037));
  nand_5 g2306(.A(new_n2535), .B(new_n2535), .Y(new_n2692));
  nand_5     g2307(.A(new_n1787), .B(new_n648), .Y(new_n2693));
  nor_5      g2308(.A(new_n2304), .B(new_n1798), .Y(new_n2694));
  nand_5     g2309(.A(new_n2694), .B(new_n2693), .Y(new_n2695));
  and_6      g2310(.A(new_n2322), .B(new_n2301), .Y(new_n2696));
  nand_5     g2311(.A(new_n2696), .B(new_n2695), .Y(new_n2697));
  nand_5     g2312(.A(new_n2697), .B(new_n2692), .Y(new_n2698));
  nand_5     g2313(.A(new_n2698), .B(new_n1998), .Y(new_n2699));
  nand_5     g2314(.A(new_n2699), .B(new_n2358), .Y(new_n2700));
  and_6      g2315(.A(new_n910), .B(new_n913), .Y(new_n2701));
  and_6      g2316(.A(new_n2701), .B(new_n2364), .Y(new_n2702));
  nand_5     g2317(.A(new_n2702), .B(new_n2700), .Y(new_n2703));
  nand_5     g2318(.A(pi247), .B(new_n913), .Y(new_n2704));
  and_6      g2319(.A(new_n2704), .B(new_n652), .Y(new_n2705));
  nand_5     g2320(.A(new_n2705), .B(new_n2703), .Y(new_n2706));
  nand_5     g2321(.A(new_n2706), .B(new_n651), .Y(new_n2707));
  nand_5     g2322(.A(new_n2707), .B(new_n650), .Y(new_n2708));
  nand_5     g2323(.A(new_n2708), .B(pi221), .Y(new_n2709));
  nand_5 g2324(.A(new_n2709), .B(new_n2709), .Y(po038));
  nand_5 g2325(.A(pi017), .B(pi017), .Y(new_n2711));
  nand_5     g2326(.A(new_n1764), .B(new_n1665), .Y(new_n2712));
  nand_5     g2327(.A(new_n2712), .B(new_n2711), .Y(new_n2713));
  nand_5     g2328(.A(new_n2713), .B(pi005), .Y(new_n2714));
  nand_5 g2329(.A(new_n2714), .B(new_n2714), .Y(po039));
  nand_5 g2330(.A(new_n912), .B(new_n912), .Y(new_n2716));
  nand_5     g2331(.A(new_n2417), .B(new_n2716), .Y(new_n2717));
  nand_5     g2332(.A(new_n2717), .B(new_n600), .Y(new_n2718));
  nand_5     g2333(.A(new_n2718), .B(pi189), .Y(new_n2719));
  nand_5 g2334(.A(new_n2719), .B(new_n2719), .Y(po040));
  nor_5      g2335(.A(new_n2653), .B(new_n769), .Y(new_n2721));
  nor_5      g2336(.A(new_n2721), .B(new_n873), .Y(new_n2722));
  nand_5     g2337(.A(new_n711), .B(pi035), .Y(new_n2723));
  nor_5      g2338(.A(new_n2723), .B(new_n2722), .Y(po041));
  nand_5 g2339(.A(new_n1832), .B(new_n1832), .Y(new_n2725));
  nor_5      g2340(.A(new_n2316), .B(new_n1794), .Y(new_n2726));
  nor_5      g2341(.A(new_n2726), .B(new_n2330), .Y(new_n2727));
  nor_5      g2342(.A(new_n2727), .B(new_n1982), .Y(new_n2728));
  nor_5      g2343(.A(new_n2728), .B(new_n1987), .Y(new_n2729));
  nor_5      g2344(.A(new_n2729), .B(new_n1961), .Y(new_n2730));
  nor_5      g2345(.A(new_n2730), .B(new_n1255), .Y(new_n2731));
  nor_5      g2346(.A(new_n2731), .B(new_n2725), .Y(new_n2732));
  nor_5      g2347(.A(new_n2732), .B(new_n2297), .Y(new_n2733));
  nor_5      g2348(.A(new_n2733), .B(new_n1196), .Y(new_n2734));
  nor_5      g2349(.A(new_n2734), .B(new_n1178), .Y(new_n2735));
  nor_5      g2350(.A(new_n2735), .B(new_n623), .Y(new_n2736));
  nand_5     g2351(.A(new_n995), .B(pi037), .Y(new_n2737));
  nor_5      g2352(.A(new_n2737), .B(new_n2736), .Y(po042));
  nor_5      g2353(.A(new_n2653), .B(new_n1620), .Y(new_n2739));
  nor_5      g2354(.A(new_n2739), .B(new_n1219), .Y(new_n2740));
  nand_5     g2355(.A(new_n1208), .B(pi132), .Y(new_n2741));
  nor_5      g2356(.A(new_n2741), .B(new_n2740), .Y(po043));
  and_6      g2357(.A(new_n1723), .B(pi083), .Y(po044));
  nand_5 g2358(.A(new_n596), .B(new_n596), .Y(new_n2744));
  nand_5 g2359(.A(new_n2351), .B(new_n2351), .Y(new_n2745));
  nand_5 g2360(.A(new_n1233), .B(new_n1233), .Y(new_n2746));
  nor_5      g2361(.A(new_n1938), .B(new_n2746), .Y(new_n2747));
  nand_5     g2362(.A(new_n2299), .B(new_n1937), .Y(new_n2748));
  nand_5     g2363(.A(new_n2748), .B(new_n2212), .Y(new_n2749));
  nand_5 g2364(.A(new_n2749), .B(new_n2749), .Y(new_n2750));
  nor_5      g2365(.A(new_n2667), .B(new_n2319), .Y(new_n2751));
  nand_5     g2366(.A(new_n2751), .B(new_n2750), .Y(new_n2752));
  nor_5      g2367(.A(new_n2752), .B(new_n2747), .Y(new_n2753));
  nor_5      g2368(.A(new_n2753), .B(new_n2266), .Y(new_n2754));
  nand_5     g2369(.A(new_n2754), .B(new_n2745), .Y(new_n2755));
  nand_5     g2370(.A(new_n1780), .B(new_n2016), .Y(new_n2756));
  nor_5      g2371(.A(new_n2756), .B(new_n2330), .Y(new_n2757));
  nor_5      g2372(.A(new_n2757), .B(new_n2755), .Y(new_n2758));
  nor_5      g2373(.A(new_n2758), .B(new_n2606), .Y(new_n2759));
  nand_5 g2374(.A(new_n888), .B(new_n888), .Y(new_n2760));
  nand_5     g2375(.A(new_n2282), .B(new_n2760), .Y(new_n2761));
  nor_5      g2376(.A(new_n2761), .B(new_n2759), .Y(new_n2762));
  nor_5      g2377(.A(new_n2762), .B(new_n2297), .Y(new_n2763));
  nor_5      g2378(.A(new_n2763), .B(new_n2744), .Y(new_n2764));
  nor_5      g2379(.A(new_n2764), .B(new_n588), .Y(new_n2765));
  nor_5      g2380(.A(new_n2765), .B(pi102), .Y(new_n2766));
  nor_5      g2381(.A(new_n2766), .B(new_n637), .Y(po045));
  nand_5 g2382(.A(new_n1787), .B(new_n1787), .Y(new_n2768));
  nand_5     g2383(.A(new_n1404), .B(new_n1405), .Y(new_n2769));
  and_6      g2384(.A(new_n571), .B(new_n435), .Y(new_n2770));
  nor_5      g2385(.A(new_n2770), .B(new_n453), .Y(new_n2771));
  nand_5     g2386(.A(new_n2771), .B(new_n2208), .Y(new_n2772));
  and_6      g2387(.A(new_n2772), .B(new_n2270), .Y(new_n2773));
  nand_5     g2388(.A(new_n2773), .B(new_n2267), .Y(new_n2774));
  nor_5      g2389(.A(new_n2774), .B(new_n2769), .Y(new_n2775));
  nor_5      g2390(.A(new_n2775), .B(new_n2768), .Y(new_n2776));
  nand_5     g2391(.A(new_n2776), .B(new_n1440), .Y(new_n2777));
  nor_5      g2392(.A(new_n2695), .B(new_n1971), .Y(new_n2778));
  nand_5     g2393(.A(new_n2778), .B(new_n2777), .Y(new_n2779));
  nand_5     g2394(.A(new_n2779), .B(new_n1969), .Y(new_n2780));
  nand_5     g2395(.A(new_n2780), .B(new_n1473), .Y(new_n2781));
  nand_5     g2396(.A(pi253), .B(new_n1473), .Y(new_n2782));
  and_6      g2397(.A(new_n2782), .B(pi227), .Y(new_n2783));
  and_6      g2398(.A(new_n2783), .B(new_n1946), .Y(new_n2784));
  nand_5     g2399(.A(new_n2784), .B(new_n2781), .Y(new_n2785));
  nand_5 g2400(.A(new_n2785), .B(new_n2785), .Y(po046));
  nand_5     g2401(.A(new_n2151), .B(new_n1040), .Y(new_n2787));
  nand_5     g2402(.A(new_n2787), .B(new_n1137), .Y(new_n2788));
  nor_5      g2403(.A(new_n738), .B(new_n739), .Y(new_n2789));
  nand_5     g2404(.A(new_n2789), .B(new_n2788), .Y(new_n2790));
  nand_5 g2405(.A(new_n2790), .B(new_n2790), .Y(po047));
  nor_5      g2406(.A(new_n2640), .B(new_n1260), .Y(po048));
  nand_5 g2407(.A(new_n2233), .B(new_n2233), .Y(new_n2793));
  nor_5      g2408(.A(new_n993), .B(new_n633), .Y(new_n2794));
  nand_5     g2409(.A(new_n1742), .B(new_n2220), .Y(new_n2795));
  nor_5      g2410(.A(new_n2795), .B(new_n2794), .Y(new_n2796));
  nor_5      g2411(.A(new_n2796), .B(new_n2793), .Y(new_n2797));
  nor_5      g2412(.A(new_n2797), .B(new_n2769), .Y(new_n2798));
  nand_5     g2413(.A(new_n2798), .B(new_n2272), .Y(new_n2799));
  nand_5     g2414(.A(new_n2799), .B(new_n1440), .Y(new_n2800));
  nand_5     g2415(.A(new_n2800), .B(new_n1193), .Y(new_n2801));
  nand_5     g2416(.A(new_n2801), .B(new_n642), .Y(new_n2802));
  nand_5     g2417(.A(new_n2802), .B(new_n1525), .Y(new_n2803));
  nand_5     g2418(.A(new_n2803), .B(new_n1770), .Y(new_n2804));
  nor_5      g2419(.A(new_n2804), .B(new_n580), .Y(po049));
  nor_5      g2420(.A(new_n2523), .B(new_n1327), .Y(po050));
  nor_5      g2421(.A(new_n2546), .B(pi013), .Y(new_n2807));
  nor_5      g2422(.A(new_n2807), .B(pi051), .Y(new_n2808));
  nor_5      g2423(.A(new_n2808), .B(pi168), .Y(new_n2809));
  nor_5      g2424(.A(new_n2809), .B(pi179), .Y(new_n2810));
  nor_5      g2425(.A(new_n2810), .B(pi106), .Y(new_n2811));
  nor_5      g2426(.A(new_n2811), .B(new_n2085), .Y(new_n2812));
  nor_5      g2427(.A(new_n2812), .B(new_n2109), .Y(new_n2813));
  nor_5      g2428(.A(new_n2813), .B(new_n2080), .Y(new_n2814));
  nor_5      g2429(.A(new_n2814), .B(new_n504), .Y(po051));
  nand_5     g2430(.A(new_n2631), .B(new_n928), .Y(new_n2816));
  nand_5 g2431(.A(new_n2752), .B(new_n2752), .Y(new_n2817));
  nand_5 g2432(.A(new_n2414), .B(new_n2414), .Y(new_n2818));
  nand_5 g2433(.A(new_n813), .B(new_n813), .Y(new_n2819));
  nand_5     g2434(.A(new_n1784), .B(new_n2819), .Y(new_n2820));
  nor_5      g2435(.A(new_n2820), .B(new_n2224), .Y(new_n2821));
  nand_5     g2436(.A(new_n2821), .B(new_n2818), .Y(new_n2822));
  nor_5      g2437(.A(new_n2822), .B(new_n1779), .Y(new_n2823));
  nand_5     g2438(.A(new_n2823), .B(new_n2817), .Y(new_n2824));
  nor_5      g2439(.A(new_n2824), .B(new_n2498), .Y(new_n2825));
  nand_5     g2440(.A(new_n2825), .B(new_n2610), .Y(new_n2826));
  nand_5     g2441(.A(new_n2826), .B(new_n2816), .Y(new_n2827));
  nor_5      g2442(.A(new_n2827), .B(new_n1810), .Y(new_n2828));
  nand_5     g2443(.A(new_n1112), .B(pi124), .Y(new_n2829));
  nor_5      g2444(.A(new_n2829), .B(new_n2828), .Y(po052));
  nand_5     g2445(.A(new_n2376), .B(new_n497), .Y(new_n2831));
  nand_5     g2446(.A(new_n2831), .B(new_n2564), .Y(new_n2832));
  nand_5     g2447(.A(new_n2832), .B(new_n2425), .Y(new_n2833));
  nand_5     g2448(.A(new_n2833), .B(new_n1351), .Y(new_n2834));
  nand_5     g2449(.A(new_n2834), .B(new_n1883), .Y(new_n2835));
  nand_5     g2450(.A(new_n2835), .B(pi246), .Y(new_n2836));
  nand_5 g2451(.A(new_n2836), .B(new_n2836), .Y(po053));
  and_6      g2452(.A(new_n2702), .B(new_n2597), .Y(new_n2838));
  nor_5      g2453(.A(new_n2838), .B(new_n2706), .Y(new_n2839));
  nor_5      g2454(.A(new_n2839), .B(new_n651), .Y(po054));
  nor_5      g2455(.A(new_n2342), .B(pi202), .Y(new_n2841));
  nand_5     g2456(.A(new_n1046), .B(pi085), .Y(new_n2842));
  nor_5      g2457(.A(new_n2842), .B(new_n2841), .Y(po055));
  nor_5      g2458(.A(new_n1953), .B(pi215), .Y(new_n2844));
  nor_5      g2459(.A(new_n2844), .B(pi105), .Y(new_n2845));
  nor_5      g2460(.A(new_n2845), .B(new_n517), .Y(po056));
  nand_5 g2461(.A(new_n570), .B(new_n570), .Y(new_n2847));
  nand_5     g2462(.A(new_n2781), .B(new_n565), .Y(new_n2848));
  nand_5     g2463(.A(new_n2848), .B(new_n2847), .Y(new_n2849));
  nand_5     g2464(.A(new_n2849), .B(pi010), .Y(new_n2850));
  nand_5 g2465(.A(new_n2850), .B(new_n2850), .Y(po057));
  nand_5     g2466(.A(new_n2755), .B(new_n2530), .Y(new_n2852));
  nand_5     g2467(.A(new_n2852), .B(new_n2734), .Y(new_n2853));
  nand_5     g2468(.A(new_n2853), .B(new_n1177), .Y(new_n2854));
  nor_5      g2469(.A(new_n2854), .B(new_n991), .Y(new_n2855));
  nor_5      g2470(.A(new_n2855), .B(pi217), .Y(new_n2856));
  nor_5      g2471(.A(new_n2856), .B(new_n1447), .Y(po058));
  nand_5 g2472(.A(pi191), .B(pi191), .Y(new_n2858));
  nand_5 g2473(.A(new_n855), .B(new_n855), .Y(new_n2859));
  nor_5      g2474(.A(new_n856), .B(new_n2859), .Y(new_n2860));
  nand_5     g2475(.A(new_n2860), .B(new_n851), .Y(new_n2861));
  nand_5 g2476(.A(new_n2861), .B(new_n2861), .Y(new_n2862));
  nand_5     g2477(.A(new_n1381), .B(new_n1200), .Y(new_n2863));
  nor_5      g2478(.A(new_n2863), .B(new_n2862), .Y(new_n2864));
  nand_5     g2479(.A(new_n2170), .B(new_n1737), .Y(new_n2865));
  nor_5      g2480(.A(new_n2865), .B(new_n2864), .Y(new_n2866));
  nor_5      g2481(.A(new_n2866), .B(new_n2474), .Y(new_n2867));
  nor_5      g2482(.A(new_n2867), .B(new_n2394), .Y(new_n2868));
  nor_5      g2483(.A(new_n2868), .B(new_n2411), .Y(new_n2869));
  nand_5     g2484(.A(new_n2459), .B(new_n2395), .Y(new_n2870));
  and_6      g2485(.A(new_n2870), .B(new_n1120), .Y(new_n2871));
  nand_5     g2486(.A(new_n2871), .B(new_n2869), .Y(new_n2872));
  nand_5     g2487(.A(new_n2872), .B(new_n2858), .Y(new_n2873));
  nand_5     g2488(.A(new_n2873), .B(new_n756), .Y(new_n2874));
  nand_5     g2489(.A(new_n2869), .B(new_n1126), .Y(new_n2875));
  nand_5     g2490(.A(new_n2875), .B(new_n2874), .Y(new_n2876));
  nand_5     g2491(.A(new_n2876), .B(new_n757), .Y(new_n2877));
  and_6      g2492(.A(new_n762), .B(pi046), .Y(new_n2878));
  nand_5     g2493(.A(new_n2878), .B(new_n2877), .Y(new_n2879));
  nand_5 g2494(.A(new_n2879), .B(new_n2879), .Y(po059));
  nand_5 g2495(.A(pi107), .B(pi107), .Y(new_n2881));
  nor_5      g2496(.A(new_n986), .B(new_n2881), .Y(new_n2882));
  and_6      g2497(.A(new_n2882), .B(new_n984), .Y(new_n2883));
  nand_5     g2498(.A(new_n2883), .B(new_n990), .Y(new_n2884));
  nor_5      g2499(.A(new_n2884), .B(new_n2854), .Y(po060));
  nand_5     g2500(.A(new_n829), .B(pi208), .Y(new_n2886));
  nor_5      g2501(.A(new_n2886), .B(new_n2505), .Y(po061));
  nand_5 g2502(.A(new_n2812), .B(new_n2812), .Y(new_n2888));
  nand_5     g2503(.A(new_n2888), .B(new_n2108), .Y(new_n2889));
  nor_5      g2504(.A(new_n2889), .B(new_n1006), .Y(po062));
  nand_5 g2505(.A(new_n2339), .B(new_n2339), .Y(new_n2891));
  nor_5      g2506(.A(new_n2891), .B(pi000), .Y(new_n2892));
  nor_5      g2507(.A(new_n2892), .B(pi161), .Y(new_n2893));
  nand_5     g2508(.A(new_n1252), .B(pi231), .Y(new_n2894));
  nor_5      g2509(.A(new_n2894), .B(new_n2893), .Y(po063));
  nand_5     g2510(.A(new_n1725), .B(pi145), .Y(new_n2896));
  nand_5 g2511(.A(new_n2896), .B(new_n2896), .Y(po064));
  nor_5      g2512(.A(new_n2463), .B(new_n2141), .Y(new_n2898));
  nand_5     g2513(.A(new_n2898), .B(new_n2134), .Y(new_n2899));
  nand_5     g2514(.A(new_n2899), .B(new_n2482), .Y(new_n2900));
  nand_5     g2515(.A(new_n2900), .B(new_n2163), .Y(new_n2901));
  nand_5     g2516(.A(new_n2901), .B(new_n2084), .Y(new_n2902));
  nand_5     g2517(.A(new_n530), .B(pi050), .Y(new_n2903));
  nand_5     g2518(.A(new_n2903), .B(new_n2106), .Y(new_n2904));
  nand_5 g2519(.A(new_n2904), .B(new_n2904), .Y(new_n2905));
  nand_5     g2520(.A(new_n2905), .B(new_n2902), .Y(new_n2906));
  nand_5 g2521(.A(new_n2906), .B(new_n2906), .Y(new_n2907));
  nor_5      g2522(.A(new_n2907), .B(pi067), .Y(new_n2908));
  nand_5     g2523(.A(new_n529), .B(pi252), .Y(new_n2909));
  nor_5      g2524(.A(new_n2909), .B(new_n2908), .Y(po065));
  nor_5      g2525(.A(new_n2906), .B(new_n518), .Y(po066));
  nor_5      g2526(.A(new_n2662), .B(new_n1639), .Y(new_n2912));
  nand_5     g2527(.A(new_n2912), .B(new_n2161), .Y(new_n2913));
  nor_5      g2528(.A(new_n2913), .B(new_n2529), .Y(new_n2914));
  nor_5      g2529(.A(new_n2914), .B(new_n2413), .Y(new_n2915));
  nand_5     g2530(.A(new_n1859), .B(new_n903), .Y(new_n2916));
  nor_5      g2531(.A(new_n2916), .B(new_n2915), .Y(new_n2917));
  nor_5      g2532(.A(new_n2917), .B(new_n1642), .Y(new_n2918));
  nor_5      g2533(.A(new_n2918), .B(new_n661), .Y(po067));
  nand_5     g2534(.A(new_n587), .B(pi166), .Y(new_n2920));
  nor_5      g2535(.A(new_n2920), .B(new_n2764), .Y(po068));
  and_6      g2536(.A(new_n796), .B(pi229), .Y(new_n2922));
  and_6      g2537(.A(new_n2922), .B(new_n2633), .Y(po069));
  nor_5      g2538(.A(new_n2641), .B(new_n1289), .Y(new_n2924));
  nand_5     g2539(.A(new_n1287), .B(pi028), .Y(new_n2925));
  nor_5      g2540(.A(new_n2925), .B(new_n2924), .Y(po070));
  nand_5 g2541(.A(new_n2259), .B(new_n2259), .Y(new_n2927));
  nand_5     g2542(.A(new_n2296), .B(new_n2927), .Y(new_n2928));
  nand_5     g2543(.A(new_n2928), .B(new_n1866), .Y(new_n2929));
  nand_5     g2544(.A(new_n2929), .B(new_n1864), .Y(new_n2930));
  nor_5      g2545(.A(new_n1938), .B(new_n1802), .Y(new_n2931));
  nand_5     g2546(.A(new_n2931), .B(new_n2930), .Y(new_n2932));
  nand_5     g2547(.A(new_n2932), .B(new_n2750), .Y(new_n2933));
  nand_5     g2548(.A(new_n2933), .B(new_n551), .Y(new_n2934));
  nand_5     g2549(.A(new_n2934), .B(new_n2322), .Y(new_n2935));
  nand_5     g2550(.A(new_n2935), .B(new_n2195), .Y(new_n2936));
  nand_5     g2551(.A(new_n2936), .B(new_n1914), .Y(new_n2937));
  nand_5     g2552(.A(new_n2937), .B(new_n468), .Y(new_n2938));
  nand_5     g2553(.A(new_n2938), .B(pi016), .Y(new_n2939));
  nand_5 g2554(.A(new_n2939), .B(new_n2939), .Y(po071));
  nor_5      g2555(.A(new_n2598), .B(new_n1107), .Y(new_n2941));
  nor_5      g2556(.A(new_n2941), .B(pi031), .Y(new_n2942));
  nor_5      g2557(.A(new_n2942), .B(new_n2670), .Y(po072));
  nand_5 g2558(.A(pi097), .B(pi097), .Y(new_n2944));
  nand_5     g2559(.A(new_n2817), .B(new_n1236), .Y(new_n2945));
  nand_5     g2560(.A(new_n2945), .B(new_n2754), .Y(new_n2946));
  nand_5     g2561(.A(new_n2946), .B(new_n1988), .Y(new_n2947));
  nand_5     g2562(.A(new_n2947), .B(new_n1429), .Y(new_n2948));
  nand_5     g2563(.A(new_n2948), .B(new_n1271), .Y(new_n2949));
  nor_5      g2564(.A(new_n1297), .B(pi036), .Y(new_n2950));
  nand_5     g2565(.A(new_n2950), .B(new_n2949), .Y(new_n2951));
  nand_5     g2566(.A(new_n2951), .B(new_n1243), .Y(new_n2952));
  nand_5     g2567(.A(new_n2952), .B(new_n2944), .Y(new_n2953));
  nand_5     g2568(.A(new_n2953), .B(pi027), .Y(new_n2954));
  nand_5 g2569(.A(new_n2954), .B(new_n2954), .Y(po073));
  nand_5 g2570(.A(new_n493), .B(new_n493), .Y(new_n2956));
  nor_5      g2571(.A(new_n2814), .B(pi143), .Y(new_n2957));
  nor_5      g2572(.A(new_n2957), .B(new_n2956), .Y(new_n2958));
  nand_5 g2573(.A(new_n495), .B(new_n495), .Y(new_n2959));
  nand_5     g2574(.A(new_n2959), .B(pi199), .Y(new_n2960));
  nor_5      g2575(.A(new_n2960), .B(new_n2958), .Y(po074));
  nand_5     g2576(.A(new_n2951), .B(pi236), .Y(new_n2962));
  nand_5 g2577(.A(new_n2962), .B(new_n2962), .Y(po075));
  nand_5 g2578(.A(new_n859), .B(new_n859), .Y(new_n2964));
  nand_5     g2579(.A(new_n1373), .B(new_n2964), .Y(new_n2965));
  and_6      g2580(.A(new_n2965), .B(pi151), .Y(new_n2966));
  and_6      g2581(.A(new_n2966), .B(new_n2875), .Y(po076));
  nor_5      g2582(.A(new_n1699), .B(new_n850), .Y(new_n2968));
  nor_5      g2583(.A(new_n2968), .B(new_n1818), .Y(new_n2969));
  nand_5     g2584(.A(new_n1843), .B(pi158), .Y(new_n2970));
  nor_5      g2585(.A(new_n2970), .B(new_n2969), .Y(po077));
  nor_5      g2586(.A(new_n2430), .B(new_n1335), .Y(new_n2972));
  nor_5      g2587(.A(new_n2972), .B(new_n1332), .Y(po078));
  nor_5      g2588(.A(new_n2918), .B(pi201), .Y(new_n2974));
  nor_5      g2589(.A(new_n2974), .B(pi078), .Y(new_n2975));
  nor_5      g2590(.A(new_n2975), .B(pi196), .Y(new_n2976));
  nor_5      g2591(.A(new_n2976), .B(pi247), .Y(new_n2977));
  nor_5      g2592(.A(new_n2977), .B(new_n913), .Y(po079));
  nor_5      g2593(.A(new_n2855), .B(new_n621), .Y(new_n2979));
  nand_5     g2594(.A(new_n619), .B(pi019), .Y(new_n2980));
  nor_5      g2595(.A(new_n2980), .B(new_n2979), .Y(po080));
  nor_5      g2596(.A(new_n2802), .B(new_n579), .Y(po081));
  nor_5      g2597(.A(new_n2889), .B(pi198), .Y(new_n2983));
  nor_5      g2598(.A(new_n2983), .B(pi047), .Y(new_n2984));
  nor_5      g2599(.A(new_n2984), .B(new_n513), .Y(po082));
  nor_5      g2600(.A(new_n2957), .B(pi025), .Y(new_n2986));
  nor_5      g2601(.A(new_n2986), .B(new_n494), .Y(po083));
  and_6      g2602(.A(new_n790), .B(pi110), .Y(new_n2988));
  and_6      g2603(.A(new_n2988), .B(new_n2827), .Y(po084));
  and_6      g2604(.A(new_n1912), .B(pi139), .Y(new_n2990));
  nand_5     g2605(.A(new_n2990), .B(new_n2936), .Y(new_n2991));
  nand_5 g2606(.A(new_n2991), .B(new_n2991), .Y(po085));
  nor_5      g2607(.A(new_n2636), .B(pi150), .Y(new_n2993));
  nor_5      g2608(.A(new_n2993), .B(pi004), .Y(new_n2994));
  nor_5      g2609(.A(new_n2994), .B(new_n773), .Y(po086));
  nor_5      g2610(.A(new_n2520), .B(pi220), .Y(new_n2996));
  nor_5      g2611(.A(new_n2996), .B(pi069), .Y(new_n2997));
  nor_5      g2612(.A(new_n2997), .B(new_n428), .Y(po087));
  nor_5      g2613(.A(new_n2290), .B(new_n1682), .Y(new_n2999));
  nor_5      g2614(.A(new_n2999), .B(new_n1301), .Y(new_n3000));
  nand_5     g2615(.A(new_n1141), .B(pi065), .Y(new_n3001));
  nor_5      g2616(.A(new_n3001), .B(new_n3000), .Y(po088));
  nand_5     g2617(.A(new_n440), .B(pi239), .Y(new_n3003));
  nor_5      g2618(.A(new_n3003), .B(new_n2002), .Y(po089));
  and_6      g2619(.A(new_n2449), .B(new_n962), .Y(new_n3005));
  nand_5     g2620(.A(new_n954), .B(pi116), .Y(new_n3006));
  nor_5      g2621(.A(new_n3006), .B(new_n3005), .Y(po090));
  nand_5 g2622(.A(pi064), .B(pi064), .Y(new_n3008));
  nor_5      g2623(.A(new_n2876), .B(new_n3008), .Y(po091));
  nand_5     g2624(.A(new_n2938), .B(new_n455), .Y(new_n3010));
  nand_5     g2625(.A(new_n3010), .B(new_n476), .Y(new_n3011));
  nand_5     g2626(.A(new_n3011), .B(pi056), .Y(new_n3012));
  nand_5 g2627(.A(new_n3012), .B(new_n3012), .Y(po092));
  nand_5 g2628(.A(pi180), .B(pi180), .Y(new_n3014));
  nor_5      g2629(.A(new_n2804), .B(pi248), .Y(new_n3015));
  nor_5      g2630(.A(new_n3015), .B(pi100), .Y(new_n3016));
  nor_5      g2631(.A(new_n3016), .B(pi063), .Y(new_n3017));
  nor_5      g2632(.A(new_n3017), .B(pi113), .Y(new_n3018));
  nor_5      g2633(.A(new_n3018), .B(new_n3014), .Y(po093));
  nand_5     g2634(.A(new_n2518), .B(new_n2121), .Y(new_n3020));
  and_6      g2635(.A(new_n1897), .B(pi232), .Y(new_n3021));
  nand_5     g2636(.A(new_n3021), .B(new_n3020), .Y(new_n3022));
  nand_5 g2637(.A(new_n3022), .B(new_n3022), .Y(po094));
  nor_5      g2638(.A(new_n2621), .B(new_n485), .Y(po095));
  nand_5     g2639(.A(new_n2835), .B(new_n398), .Y(new_n3025));
  nand_5     g2640(.A(new_n3025), .B(new_n2251), .Y(new_n3026));
  nand_5     g2641(.A(new_n3026), .B(pi146), .Y(new_n3027));
  nand_5 g2642(.A(new_n3027), .B(new_n3027), .Y(po096));
  nand_5 g2643(.A(new_n554), .B(new_n554), .Y(new_n3029));
  nand_5     g2644(.A(new_n2516), .B(new_n3029), .Y(new_n3030));
  and_6      g2645(.A(new_n454), .B(pi126), .Y(new_n3031));
  nand_5     g2646(.A(new_n3031), .B(new_n3030), .Y(new_n3032));
  nand_5 g2647(.A(new_n3032), .B(new_n3032), .Y(po097));
  nor_5      g2648(.A(new_n2003), .B(pi076), .Y(new_n3034));
  nor_5      g2649(.A(new_n3034), .B(new_n443), .Y(po098));
  nand_5 g2650(.A(new_n1381), .B(new_n1381), .Y(new_n3036));
  nor_5      g2651(.A(new_n1848), .B(new_n1699), .Y(new_n3037));
  nor_5      g2652(.A(new_n3037), .B(new_n3036), .Y(new_n3038));
  nand_5     g2653(.A(new_n1382), .B(pi104), .Y(new_n3039));
  nor_5      g2654(.A(new_n3039), .B(new_n3038), .Y(po099));
  nor_5      g2655(.A(new_n2518), .B(new_n447), .Y(po100));
  nand_5     g2656(.A(new_n844), .B(pi243), .Y(new_n3042));
  nor_5      g2657(.A(new_n3042), .B(new_n1726), .Y(po101));
  nand_5     g2658(.A(new_n2689), .B(new_n743), .Y(new_n3044));
  nand_5     g2659(.A(new_n3044), .B(new_n747), .Y(new_n3045));
  nor_5      g2660(.A(new_n3045), .B(new_n735), .Y(po102));
  nand_5     g2661(.A(new_n2869), .B(new_n1402), .Y(new_n3047));
  and_6      g2662(.A(new_n1374), .B(new_n725), .Y(new_n3048));
  nand_5     g2663(.A(new_n3048), .B(new_n3047), .Y(new_n3049));
  nand_5 g2664(.A(new_n860), .B(new_n860), .Y(new_n3050));
  nor_5      g2665(.A(new_n3050), .B(pi140), .Y(new_n3051));
  nand_5     g2666(.A(new_n3051), .B(new_n3049), .Y(new_n3052));
  nand_5     g2667(.A(new_n3052), .B(pi001), .Y(new_n3053));
  nand_5 g2668(.A(new_n3053), .B(new_n3053), .Y(po103));
  nor_5      g2669(.A(new_n3045), .B(pi148), .Y(new_n3055));
  nor_5      g2670(.A(new_n3055), .B(pi086), .Y(new_n3056));
  nor_5      g2671(.A(new_n3056), .B(new_n751), .Y(po104));
  nor_5      g2672(.A(new_n1241), .B(new_n1242), .Y(new_n3058));
  and_6      g2673(.A(new_n3058), .B(new_n2948), .Y(po105));
  nor_5      g2674(.A(new_n2833), .B(new_n2337), .Y(new_n3060));
  nor_5      g2675(.A(new_n3060), .B(new_n2295), .Y(new_n3061));
  nor_5      g2676(.A(new_n3061), .B(new_n1293), .Y(new_n3062));
  nor_5      g2677(.A(new_n3062), .B(new_n1269), .Y(po106));
  nand_5     g2678(.A(new_n563), .B(pi253), .Y(new_n3064));
  nor_5      g2679(.A(new_n3064), .B(new_n2780), .Y(po107));
  nor_5      g2680(.A(new_n386), .B(pi131), .Y(new_n3066));
  nor_5      g2681(.A(new_n3066), .B(new_n1276), .Y(new_n3067));
  and_6      g2682(.A(new_n3067), .B(new_n2009), .Y(po108));
  nor_5      g2683(.A(new_n2721), .B(new_n871), .Y(new_n3069));
  nor_5      g2684(.A(new_n3069), .B(new_n1617), .Y(po109));
  nand_5     g2685(.A(new_n834), .B(pi173), .Y(new_n3071));
  nor_5      g2686(.A(new_n3071), .B(new_n1699), .Y(po110));
  nor_5      g2687(.A(new_n2765), .B(new_n636), .Y(new_n3073));
  nand_5     g2688(.A(new_n639), .B(pi219), .Y(new_n3074));
  nor_5      g2689(.A(new_n3074), .B(new_n3073), .Y(po111));
  nand_5     g2690(.A(new_n2708), .B(new_n649), .Y(new_n3076));
  nand_5     g2691(.A(new_n3076), .B(new_n606), .Y(new_n3077));
  nand_5     g2692(.A(new_n3077), .B(pi185), .Y(new_n3078));
  nand_5 g2693(.A(new_n3078), .B(new_n3078), .Y(po112));
  nor_5      g2694(.A(new_n3016), .B(new_n1653), .Y(po113));
  nor_5      g2695(.A(new_n2937), .B(new_n457), .Y(new_n3081));
  nor_5      g2696(.A(new_n3081), .B(new_n2131), .Y(new_n3082));
  nor_5      g2697(.A(new_n3082), .B(new_n1457), .Y(po114));
  and_6      g2698(.A(new_n2290), .B(new_n1511), .Y(new_n3084));
  and_6      g2699(.A(new_n1257), .B(pi157), .Y(new_n3085));
  nand_5     g2700(.A(new_n3085), .B(new_n1543), .Y(new_n3086));
  nor_5      g2701(.A(new_n3086), .B(new_n3084), .Y(po115));
  nor_5      g2702(.A(new_n2834), .B(new_n399), .Y(new_n3088));
  nor_5      g2703(.A(new_n3088), .B(new_n2553), .Y(new_n3089));
  nor_5      g2704(.A(new_n3089), .B(new_n2189), .Y(po116));
  and_6      g2705(.A(new_n2833), .B(pi121), .Y(po117));
  nand_5     g2706(.A(new_n1835), .B(pi000), .Y(new_n3092));
  nor_5      g2707(.A(new_n3092), .B(new_n2891), .Y(po118));
  nor_5      g2708(.A(new_n2808), .B(new_n689), .Y(po119));
  nor_5      g2709(.A(new_n2451), .B(pi002), .Y(new_n3095));
  nor_5      g2710(.A(new_n3095), .B(pi096), .Y(new_n3096));
  nor_5      g2711(.A(new_n3096), .B(new_n950), .Y(po120));
  nand_5 g2712(.A(pi129), .B(pi129), .Y(new_n3098));
  nor_5      g2713(.A(new_n2055), .B(new_n3098), .Y(po121));
  nor_5      g2714(.A(new_n2975), .B(new_n659), .Y(po122));
  nor_5      g2715(.A(new_n2578), .B(pi245), .Y(new_n3101));
  nor_5      g2716(.A(new_n3101), .B(pi101), .Y(new_n3102));
  nor_5      g2717(.A(new_n3102), .B(new_n1034), .Y(po123));
  nor_5      g2718(.A(new_n2619), .B(new_n486), .Y(po124));
  nor_5      g2719(.A(new_n2810), .B(new_n1758), .Y(po125));
  nand_5     g2720(.A(new_n1106), .B(pi091), .Y(new_n3106));
  nor_5      g2721(.A(new_n3106), .B(new_n2598), .Y(po126));
  nor_5      g2722(.A(new_n2993), .B(new_n1119), .Y(new_n3108));
  nand_5     g2723(.A(new_n1118), .B(pi191), .Y(new_n3109));
  nor_5      g2724(.A(new_n3109), .B(new_n3108), .Y(po127));
  or_6       g2725(.A(new_n1135), .B(new_n951), .Y(new_n3111));
  nor_5      g2726(.A(new_n1155), .B(pi044), .Y(new_n3112));
  nand_5     g2727(.A(new_n3112), .B(new_n2575), .Y(new_n3113));
  nand_5     g2728(.A(new_n3113), .B(new_n3111), .Y(new_n3114));
  nand_5     g2729(.A(new_n3114), .B(pi205), .Y(new_n3115));
  nand_5 g2730(.A(new_n3115), .B(new_n3115), .Y(po128));
endmodule


