// Benchmark "top_809568696_809776567_809698999_863110837_1234615" written by ABC on Mon Aug 19 01:01:33 2024

module top_809568696_809776567_809698999_863110837_1234615 ( 
    c, d,
    o  );
  input  c, d;
  output o;
  assign o = c & d;
endmodule


