module top_1598227639_809568180_776209382_1234615 (a, b, c, d, e, f, g, h, o);
 input a, b, c, d, e, f, g, h;
 output o;
 and_1 g0(a,b,y1); // 1
 and_1 g1(y1,y1,y2); // 2
 // and_1 g2(d,y2,y3); // 3
 // and_1 g3(y1,y3,y4); // 3
 // and_1 g4(y2,y2,y5);
 // and_1 g5(y3,y4,y6);
 // and_1 g6(y5,y6,o);
endmodule
