// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Mon Aug 12 17:42:23 2024

module top_810026173_826291639_946996917_1246901 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83,
    pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81,
    pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181;
  wire new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n501, new_n504, new_n505, new_n507, new_n508,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n781, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n831, new_n832, new_n833,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1099,
    new_n1102, new_n1103, new_n1105, new_n1107, new_n1109, new_n1110,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1139, new_n1141,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1155, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1353, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1398, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1433, new_n1434, new_n1435, new_n1436, new_n1437, new_n1438,
    new_n1439, new_n1440, new_n1441, new_n1442, new_n1443, new_n1444,
    new_n1445, new_n1446, new_n1447, new_n1448, new_n1449, new_n1450,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1459, new_n1460,
    new_n1461, new_n1466, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1480, new_n1481, new_n1482, new_n1483, new_n1485,
    new_n1488, new_n1489, new_n1490, new_n1494, new_n1495, new_n1497,
    new_n1498, new_n1501, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1516,
    new_n1517, new_n1521, new_n1522, new_n1523, new_n1524, new_n1527,
    new_n1528, new_n1531, new_n1532, new_n1533, new_n1540, new_n1543,
    new_n1552, new_n1555, new_n1557, new_n1558, new_n1570, new_n1573,
    new_n1575, new_n1576, new_n1580, new_n1581, new_n1587, new_n1589,
    new_n1590;
  nor_5  g0000(.A(pi60), .B(pi59), .Y(new_n276));
  not_8  g0001(.A(pi60), .Y(new_n277));
  nor_5  g0002(.A(new_n277), .B(pi32), .Y(new_n278));
  nor_5  g0003(.A(new_n278), .B(new_n276), .Y(new_n279));
  nor_5  g0004(.A(new_n277), .B(pi51), .Y(new_n280));
  nor_5  g0005(.A(pi60), .B(pi06), .Y(new_n281));
  nor_5  g0006(.A(new_n281), .B(new_n280), .Y(new_n282));
  nor_5  g0007(.A(new_n282), .B(new_n279), .Y(new_n283));
  not_8  g0008(.A(new_n283), .Y(new_n284));
  nor_5  g0009(.A(pi75), .B(pi60), .Y(new_n285));
  nor_5  g0010(.A(new_n277), .B(pi08), .Y(new_n286));
  nor_5  g0011(.A(new_n286), .B(new_n285), .Y(new_n287));
  xor_4  g0012(.A(new_n287), .B(new_n284), .Y(new_n288));
  not_8  g0013(.A(pi41), .Y(new_n289));
  xor_4  g0014(.A(new_n282), .B(new_n279), .Y(new_n290));
  nor_5  g0015(.A(new_n290), .B(new_n289), .Y(new_n291));
  xor_4  g0016(.A(new_n290), .B(new_n289), .Y(new_n292));
  not_8  g0017(.A(new_n292), .Y(new_n293));
  not_8  g0018(.A(pi91), .Y(new_n294));
  nand_5 g0019(.A(new_n279), .B(new_n294), .Y(new_n295));
  or_6   g0020(.A(new_n279), .B(new_n294), .Y(new_n296));
  nor_5  g0021(.A(pi76), .B(new_n277), .Y(new_n297));
  nor_5  g0022(.A(pi60), .B(pi18), .Y(new_n298));
  nor_5  g0023(.A(new_n298), .B(new_n297), .Y(new_n299));
  nand_5 g0024(.A(new_n299), .B(pi79), .Y(new_n300));
  nand_5 g0025(.A(new_n300), .B(new_n296), .Y(new_n301));
  nand_5 g0026(.A(new_n301), .B(new_n295), .Y(new_n302));
  nor_5  g0027(.A(new_n302), .B(new_n293), .Y(new_n303));
  nor_5  g0028(.A(new_n303), .B(new_n291), .Y(new_n304));
  or_6   g0029(.A(new_n304), .B(new_n288), .Y(new_n305));
  nor_5  g0030(.A(new_n287), .B(new_n284), .Y(new_n306));
  nor_5  g0031(.A(pi86), .B(new_n277), .Y(new_n307));
  nor_5  g0032(.A(pi60), .B(pi39), .Y(new_n308));
  nor_5  g0033(.A(new_n308), .B(new_n307), .Y(new_n309));
  xor_4  g0034(.A(new_n309), .B(new_n306), .Y(new_n310));
  or_6   g0035(.A(new_n310), .B(new_n305), .Y(new_n311));
  nand_5 g0036(.A(new_n309), .B(new_n306), .Y(new_n312));
  xor_4  g0037(.A(pi86), .B(pi34), .Y(new_n313));
  nor_5  g0038(.A(new_n313), .B(new_n277), .Y(new_n314));
  nor_5  g0039(.A(pi82), .B(pi39), .Y(new_n315));
  nand_5 g0040(.A(pi82), .B(pi39), .Y(new_n316));
  nand_5 g0041(.A(new_n316), .B(new_n277), .Y(new_n317));
  nor_5  g0042(.A(new_n317), .B(new_n315), .Y(new_n318));
  nor_5  g0043(.A(new_n318), .B(new_n314), .Y(new_n319));
  xor_4  g0044(.A(new_n319), .B(new_n312), .Y(new_n320));
  or_6   g0045(.A(new_n320), .B(new_n311), .Y(new_n321));
  or_6   g0046(.A(new_n319), .B(new_n312), .Y(new_n322));
  xor_4  g0047(.A(new_n315), .B(pi04), .Y(new_n323));
  nand_5 g0048(.A(new_n323), .B(new_n277), .Y(new_n324));
  not_8  g0049(.A(pi02), .Y(new_n325));
  nand_5 g0050(.A(pi86), .B(pi34), .Y(new_n326));
  nand_5 g0051(.A(new_n326), .B(new_n325), .Y(new_n327));
  nor_5  g0052(.A(new_n326), .B(new_n325), .Y(new_n328));
  nor_5  g0053(.A(new_n328), .B(new_n277), .Y(new_n329));
  nand_5 g0054(.A(new_n329), .B(new_n327), .Y(new_n330));
  nand_5 g0055(.A(new_n330), .B(new_n324), .Y(new_n331));
  xor_4  g0056(.A(new_n331), .B(new_n322), .Y(new_n332));
  xor_4  g0057(.A(new_n332), .B(new_n321), .Y(new_n333));
  not_8  g0058(.A(pi25), .Y(new_n334));
  nand_5 g0059(.A(pi85), .B(pi03), .Y(new_n335));
  xor_4  g0060(.A(pi85), .B(pi03), .Y(new_n336));
  nand_5 g0061(.A(pi47), .B(pi30), .Y(new_n337));
  nand_5 g0062(.A(pi45), .B(pi19), .Y(new_n338));
  xor_4  g0063(.A(pi45), .B(pi19), .Y(new_n339));
  or_6   g0064(.A(pi56), .B(pi17), .Y(new_n340));
  nand_5 g0065(.A(pi63), .B(pi55), .Y(new_n341));
  xor_4  g0066(.A(pi56), .B(pi17), .Y(new_n342));
  nand_5 g0067(.A(new_n342), .B(new_n341), .Y(new_n343));
  nand_5 g0068(.A(new_n343), .B(new_n340), .Y(new_n344));
  not_8  g0069(.A(new_n344), .Y(new_n345));
  nand_5 g0070(.A(new_n345), .B(new_n339), .Y(new_n346));
  nand_5 g0071(.A(new_n346), .B(new_n338), .Y(new_n347));
  xor_4  g0072(.A(pi47), .B(pi30), .Y(new_n348));
  nand_5 g0073(.A(new_n348), .B(new_n347), .Y(new_n349));
  nand_5 g0074(.A(new_n349), .B(new_n337), .Y(new_n350));
  nand_5 g0075(.A(new_n350), .B(new_n336), .Y(new_n351));
  nand_5 g0076(.A(new_n351), .B(new_n335), .Y(new_n352));
  nand_5 g0077(.A(new_n352), .B(pi77), .Y(new_n353));
  xor_4  g0078(.A(new_n353), .B(new_n334), .Y(new_n354));
  xor_4  g0079(.A(new_n354), .B(new_n333), .Y(new_n355));
  xor_4  g0080(.A(new_n320), .B(new_n311), .Y(new_n356));
  xor_4  g0081(.A(new_n352), .B(pi77), .Y(new_n357));
  nand_5 g0082(.A(new_n357), .B(new_n356), .Y(new_n358));
  xor_4  g0083(.A(new_n357), .B(new_n356), .Y(new_n359));
  xor_4  g0084(.A(new_n310), .B(new_n305), .Y(new_n360));
  xor_4  g0085(.A(new_n350), .B(new_n336), .Y(new_n361));
  nand_5 g0086(.A(new_n361), .B(new_n360), .Y(new_n362));
  xor_4  g0087(.A(new_n304), .B(new_n288), .Y(new_n363));
  xor_4  g0088(.A(new_n348), .B(new_n347), .Y(new_n364));
  nand_5 g0089(.A(new_n364), .B(new_n363), .Y(new_n365));
  not_8  g0090(.A(new_n364), .Y(new_n366));
  xor_4  g0091(.A(new_n366), .B(new_n363), .Y(new_n367));
  xor_4  g0092(.A(new_n302), .B(new_n293), .Y(new_n368));
  not_8  g0093(.A(new_n368), .Y(new_n369));
  xor_4  g0094(.A(new_n345), .B(new_n339), .Y(new_n370));
  not_8  g0095(.A(new_n370), .Y(new_n371));
  nand_5 g0096(.A(new_n371), .B(new_n369), .Y(new_n372));
  xor_4  g0097(.A(new_n370), .B(new_n368), .Y(new_n373));
  not_8  g0098(.A(new_n342), .Y(new_n374));
  xor_4  g0099(.A(new_n299), .B(pi79), .Y(new_n375));
  xor_4  g0100(.A(pi63), .B(pi55), .Y(new_n376));
  nand_5 g0101(.A(new_n376), .B(new_n375), .Y(new_n377));
  nor_5  g0102(.A(new_n377), .B(new_n374), .Y(new_n378));
  xor_4  g0103(.A(new_n342), .B(new_n341), .Y(new_n379));
  and_6  g0104(.A(new_n379), .B(new_n377), .Y(new_n380));
  or_6   g0105(.A(new_n380), .B(new_n378), .Y(new_n381));
  nand_5 g0106(.A(new_n296), .B(new_n295), .Y(new_n382));
  xnor_4 g0107(.A(new_n382), .B(new_n300), .Y(new_n383));
  nor_5  g0108(.A(new_n383), .B(new_n381), .Y(new_n384));
  nor_5  g0109(.A(new_n384), .B(new_n378), .Y(new_n385));
  nand_5 g0110(.A(new_n385), .B(new_n373), .Y(new_n386));
  nand_5 g0111(.A(new_n386), .B(new_n372), .Y(new_n387));
  or_6   g0112(.A(new_n387), .B(new_n367), .Y(new_n388));
  nand_5 g0113(.A(new_n388), .B(new_n365), .Y(new_n389));
  xor_4  g0114(.A(new_n361), .B(new_n360), .Y(new_n390));
  nand_5 g0115(.A(new_n390), .B(new_n389), .Y(new_n391));
  nand_5 g0116(.A(new_n391), .B(new_n362), .Y(new_n392));
  nand_5 g0117(.A(new_n392), .B(new_n359), .Y(new_n393));
  nand_5 g0118(.A(new_n393), .B(new_n358), .Y(new_n394));
  xor_4  g0119(.A(new_n394), .B(new_n355), .Y(po000));
  not_8  g0120(.A(pi73), .Y(new_n396));
  nand_5 g0121(.A(new_n396), .B(pi22), .Y(new_n397));
  nand_5 g0122(.A(new_n397), .B(pi51), .Y(new_n398));
  not_8  g0123(.A(new_n397), .Y(new_n399));
  nand_5 g0124(.A(new_n399), .B(pi06), .Y(new_n400));
  nand_5 g0125(.A(new_n400), .B(new_n398), .Y(new_n401));
  xor_4  g0126(.A(new_n401), .B(pi07), .Y(new_n402));
  nand_5 g0127(.A(new_n397), .B(pi32), .Y(new_n403));
  nand_5 g0128(.A(new_n399), .B(pi59), .Y(new_n404));
  nand_5 g0129(.A(new_n404), .B(new_n403), .Y(new_n405));
  nor_5  g0130(.A(new_n405), .B(pi57), .Y(new_n406));
  nand_5 g0131(.A(new_n397), .B(pi76), .Y(new_n407));
  nand_5 g0132(.A(new_n399), .B(pi18), .Y(new_n408));
  nand_5 g0133(.A(new_n408), .B(new_n407), .Y(new_n409));
  nand_5 g0134(.A(new_n409), .B(pi16), .Y(new_n410));
  xor_4  g0135(.A(new_n405), .B(pi57), .Y(new_n411));
  and_6  g0136(.A(new_n411), .B(new_n410), .Y(new_n412));
  nor_5  g0137(.A(new_n412), .B(new_n406), .Y(new_n413));
  xor_4  g0138(.A(new_n413), .B(new_n402), .Y(new_n414));
  xor_4  g0139(.A(new_n409), .B(pi16), .Y(new_n415));
  nand_5 g0140(.A(new_n415), .B(new_n376), .Y(new_n416));
  or_6   g0141(.A(new_n416), .B(new_n374), .Y(new_n417));
  xor_4  g0142(.A(new_n411), .B(new_n410), .Y(new_n418));
  nand_5 g0143(.A(new_n416), .B(new_n379), .Y(new_n419));
  nand_5 g0144(.A(new_n419), .B(new_n417), .Y(new_n420));
  or_6   g0145(.A(new_n420), .B(new_n418), .Y(new_n421));
  nand_5 g0146(.A(new_n421), .B(new_n417), .Y(new_n422));
  xor_4  g0147(.A(new_n422), .B(new_n414), .Y(new_n423));
  xor_4  g0148(.A(new_n423), .B(new_n370), .Y(po001));
  nand_5 g0149(.A(new_n397), .B(pi86), .Y(new_n425));
  nand_5 g0150(.A(new_n399), .B(pi39), .Y(new_n426));
  nand_5 g0151(.A(new_n426), .B(new_n425), .Y(new_n427));
  nand_5 g0152(.A(new_n427), .B(pi85), .Y(new_n428));
  xor_4  g0153(.A(new_n427), .B(pi85), .Y(new_n429));
  nand_5 g0154(.A(new_n397), .B(pi08), .Y(new_n430));
  nand_5 g0155(.A(new_n399), .B(pi75), .Y(new_n431));
  nand_5 g0156(.A(new_n431), .B(new_n430), .Y(new_n432));
  nand_5 g0157(.A(new_n432), .B(pi30), .Y(new_n433));
  nand_5 g0158(.A(new_n401), .B(pi19), .Y(new_n434));
  xor_4  g0159(.A(new_n401), .B(pi19), .Y(new_n435));
  nor_5  g0160(.A(new_n405), .B(pi56), .Y(new_n436));
  nand_5 g0161(.A(new_n409), .B(pi63), .Y(new_n437));
  not_8  g0162(.A(new_n437), .Y(new_n438));
  not_8  g0163(.A(pi56), .Y(new_n439));
  xor_4  g0164(.A(new_n405), .B(new_n439), .Y(new_n440));
  nor_5  g0165(.A(new_n440), .B(new_n438), .Y(new_n441));
  nor_5  g0166(.A(new_n441), .B(new_n436), .Y(new_n442));
  nand_5 g0167(.A(new_n442), .B(new_n435), .Y(new_n443));
  nand_5 g0168(.A(new_n443), .B(new_n434), .Y(new_n444));
  xor_4  g0169(.A(new_n432), .B(pi30), .Y(new_n445));
  nand_5 g0170(.A(new_n445), .B(new_n444), .Y(new_n446));
  nand_5 g0171(.A(new_n446), .B(new_n433), .Y(new_n447));
  nand_5 g0172(.A(new_n447), .B(new_n429), .Y(new_n448));
  nand_5 g0173(.A(new_n448), .B(new_n428), .Y(new_n449));
  not_8  g0174(.A(pi22), .Y(new_n450));
  nand_5 g0175(.A(pi34), .B(new_n450), .Y(new_n451));
  nand_5 g0176(.A(pi82), .B(pi22), .Y(new_n452));
  nand_5 g0177(.A(new_n452), .B(new_n451), .Y(new_n453));
  nand_5 g0178(.A(new_n453), .B(new_n396), .Y(new_n454));
  not_8  g0179(.A(pi34), .Y(new_n455));
  nand_5 g0180(.A(pi73), .B(new_n455), .Y(new_n456));
  nand_5 g0181(.A(new_n456), .B(new_n454), .Y(new_n457));
  and_6  g0182(.A(new_n457), .B(new_n449), .Y(new_n458));
  xor_4  g0183(.A(pi34), .B(new_n325), .Y(new_n459));
  nand_5 g0184(.A(new_n459), .B(pi73), .Y(new_n460));
  nand_5 g0185(.A(pi22), .B(pi04), .Y(new_n461));
  nor_5  g0186(.A(pi22), .B(pi02), .Y(new_n462));
  nor_5  g0187(.A(new_n462), .B(pi73), .Y(new_n463));
  nand_5 g0188(.A(new_n463), .B(new_n461), .Y(new_n464));
  nand_5 g0189(.A(new_n464), .B(new_n460), .Y(new_n465));
  nand_5 g0190(.A(new_n465), .B(new_n458), .Y(new_n466));
  not_8  g0191(.A(new_n466), .Y(new_n467));
  not_8  g0192(.A(pi13), .Y(new_n468));
  nand_5 g0193(.A(new_n455), .B(new_n325), .Y(new_n469));
  xor_4  g0194(.A(new_n469), .B(new_n468), .Y(new_n470));
  nand_5 g0195(.A(new_n470), .B(pi73), .Y(new_n471));
  nand_5 g0196(.A(pi78), .B(pi04), .Y(new_n472));
  not_8  g0197(.A(pi04), .Y(new_n473));
  not_8  g0198(.A(pi78), .Y(new_n474));
  nand_5 g0199(.A(new_n474), .B(new_n473), .Y(new_n475));
  not_8  g0200(.A(new_n475), .Y(new_n476));
  nor_5  g0201(.A(new_n476), .B(new_n450), .Y(new_n477));
  nand_5 g0202(.A(new_n477), .B(new_n472), .Y(new_n478));
  nor_5  g0203(.A(pi22), .B(pi13), .Y(new_n479));
  nor_5  g0204(.A(new_n479), .B(pi73), .Y(new_n480));
  nand_5 g0205(.A(new_n480), .B(new_n478), .Y(new_n481));
  nand_5 g0206(.A(new_n481), .B(new_n471), .Y(new_n482));
  nand_5 g0207(.A(new_n482), .B(new_n467), .Y(new_n483));
  or_6   g0208(.A(new_n469), .B(pi13), .Y(new_n484));
  xor_4  g0209(.A(new_n484), .B(pi84), .Y(new_n485));
  nor_5  g0210(.A(new_n485), .B(new_n396), .Y(new_n486));
  not_8  g0211(.A(pi20), .Y(new_n487));
  nor_5  g0212(.A(new_n476), .B(new_n487), .Y(new_n488));
  nand_5 g0213(.A(new_n476), .B(new_n487), .Y(new_n489));
  nand_5 g0214(.A(new_n489), .B(pi22), .Y(new_n490));
  nor_5  g0215(.A(new_n490), .B(new_n488), .Y(new_n491));
  not_8  g0216(.A(pi84), .Y(new_n492));
  nand_5 g0217(.A(new_n492), .B(new_n450), .Y(new_n493));
  nand_5 g0218(.A(new_n493), .B(new_n396), .Y(new_n494));
  nor_5  g0219(.A(new_n494), .B(new_n491), .Y(new_n495));
  nor_5  g0220(.A(new_n495), .B(new_n486), .Y(new_n496));
  xor_4  g0221(.A(new_n496), .B(new_n483), .Y(po179));
  xor_4  g0222(.A(new_n482), .B(new_n467), .Y(po109));
  xor_4  g0223(.A(new_n457), .B(new_n449), .Y(po177));
  xor_4  g0224(.A(new_n440), .B(new_n437), .Y(po148));
  or_6   g0225(.A(new_n409), .B(pi63), .Y(new_n501));
  nand_5 g0226(.A(new_n501), .B(new_n437), .Y(po123));
  not_8  g0227(.A(po123), .Y(po115));
  nor_5  g0228(.A(po115), .B(po148), .Y(new_n504));
  not_8  g0229(.A(new_n504), .Y(new_n505));
  xor_4  g0230(.A(new_n442), .B(new_n435), .Y(po029));
  nor_5  g0231(.A(po029), .B(new_n505), .Y(new_n507));
  not_8  g0232(.A(new_n507), .Y(new_n508));
  xor_4  g0233(.A(new_n445), .B(new_n444), .Y(po176));
  or_6   g0234(.A(po176), .B(new_n508), .Y(new_n510));
  xor_4  g0235(.A(new_n447), .B(new_n429), .Y(po064));
  and_6  g0236(.A(po064), .B(new_n510), .Y(new_n512));
  and_6  g0237(.A(new_n512), .B(po177), .Y(new_n513));
  nand_5 g0238(.A(new_n513), .B(new_n465), .Y(new_n514));
  not_8  g0239(.A(new_n514), .Y(new_n515));
  nand_5 g0240(.A(new_n515), .B(po109), .Y(new_n516));
  not_8  g0241(.A(new_n516), .Y(new_n517));
  nor_5  g0242(.A(new_n517), .B(po179), .Y(new_n518));
  nor_5  g0243(.A(new_n516), .B(new_n496), .Y(new_n519));
  nor_5  g0244(.A(new_n519), .B(new_n518), .Y(po002));
  xor_4  g0245(.A(new_n376), .B(new_n375), .Y(po003));
  not_8  g0246(.A(pi14), .Y(new_n522));
  nor_5  g0247(.A(pi51), .B(new_n522), .Y(new_n523));
  nor_5  g0248(.A(pi14), .B(pi06), .Y(new_n524));
  nor_5  g0249(.A(new_n524), .B(new_n523), .Y(new_n525));
  not_8  g0250(.A(new_n525), .Y(new_n526));
  nor_5  g0251(.A(pi75), .B(pi14), .Y(new_n527));
  nor_5  g0252(.A(new_n522), .B(pi08), .Y(new_n528));
  nor_5  g0253(.A(new_n528), .B(new_n527), .Y(new_n529));
  not_8  g0254(.A(new_n529), .Y(new_n530));
  nand_5 g0255(.A(new_n530), .B(new_n526), .Y(new_n531));
  nor_5  g0256(.A(pi86), .B(new_n522), .Y(new_n532));
  nor_5  g0257(.A(pi39), .B(pi14), .Y(new_n533));
  nor_5  g0258(.A(new_n533), .B(new_n532), .Y(new_n534));
  xor_4  g0259(.A(new_n534), .B(new_n531), .Y(new_n535));
  not_8  g0260(.A(new_n535), .Y(new_n536));
  not_8  g0261(.A(pi12), .Y(new_n537));
  xor_4  g0262(.A(new_n529), .B(new_n525), .Y(new_n538));
  or_6   g0263(.A(new_n538), .B(new_n537), .Y(new_n539));
  nand_5 g0264(.A(new_n526), .B(pi26), .Y(new_n540));
  xor_4  g0265(.A(new_n526), .B(pi26), .Y(new_n541));
  not_8  g0266(.A(new_n541), .Y(new_n542));
  nor_5  g0267(.A(pi59), .B(pi14), .Y(new_n543));
  nor_5  g0268(.A(pi32), .B(new_n522), .Y(new_n544));
  nor_5  g0269(.A(new_n544), .B(new_n543), .Y(new_n545));
  or_6   g0270(.A(new_n545), .B(pi28), .Y(new_n546));
  nor_5  g0271(.A(pi76), .B(new_n522), .Y(new_n547));
  nor_5  g0272(.A(pi18), .B(pi14), .Y(new_n548));
  nor_5  g0273(.A(new_n548), .B(new_n547), .Y(new_n549));
  nand_5 g0274(.A(new_n549), .B(pi48), .Y(new_n550));
  xor_4  g0275(.A(new_n545), .B(pi28), .Y(new_n551));
  nand_5 g0276(.A(new_n551), .B(new_n550), .Y(new_n552));
  nand_5 g0277(.A(new_n552), .B(new_n546), .Y(new_n553));
  or_6   g0278(.A(new_n553), .B(new_n542), .Y(new_n554));
  nand_5 g0279(.A(new_n554), .B(new_n540), .Y(new_n555));
  xor_4  g0280(.A(new_n538), .B(new_n537), .Y(new_n556));
  nand_5 g0281(.A(new_n556), .B(new_n555), .Y(new_n557));
  nand_5 g0282(.A(new_n557), .B(new_n539), .Y(new_n558));
  nand_5 g0283(.A(new_n558), .B(new_n536), .Y(new_n559));
  or_6   g0284(.A(new_n534), .B(new_n531), .Y(new_n560));
  not_8  g0285(.A(pi82), .Y(new_n561));
  nand_5 g0286(.A(new_n561), .B(new_n522), .Y(new_n562));
  nand_5 g0287(.A(pi34), .B(pi14), .Y(new_n563));
  nand_5 g0288(.A(new_n563), .B(new_n562), .Y(new_n564));
  xor_4  g0289(.A(new_n564), .B(new_n560), .Y(new_n565));
  or_6   g0290(.A(new_n565), .B(new_n559), .Y(new_n566));
  nor_5  g0291(.A(new_n564), .B(new_n560), .Y(new_n567));
  xor_4  g0292(.A(pi82), .B(pi04), .Y(new_n568));
  nor_5  g0293(.A(new_n568), .B(pi14), .Y(new_n569));
  nand_5 g0294(.A(pi14), .B(pi02), .Y(new_n570));
  not_8  g0295(.A(new_n570), .Y(new_n571));
  nor_5  g0296(.A(new_n571), .B(new_n569), .Y(new_n572));
  xor_4  g0297(.A(new_n572), .B(new_n567), .Y(new_n573));
  or_6   g0298(.A(new_n573), .B(new_n566), .Y(new_n574));
  nand_5 g0299(.A(new_n572), .B(new_n567), .Y(new_n575));
  nand_5 g0300(.A(new_n561), .B(new_n473), .Y(new_n576));
  xor_4  g0301(.A(new_n576), .B(new_n474), .Y(new_n577));
  nand_5 g0302(.A(new_n577), .B(new_n522), .Y(new_n578));
  nand_5 g0303(.A(pi14), .B(pi13), .Y(new_n579));
  nand_5 g0304(.A(new_n579), .B(new_n578), .Y(new_n580));
  xor_4  g0305(.A(new_n580), .B(new_n575), .Y(new_n581));
  xor_4  g0306(.A(new_n581), .B(new_n574), .Y(new_n582));
  not_8  g0307(.A(pi21), .Y(new_n583));
  nand_5 g0308(.A(pi87), .B(pi85), .Y(new_n584));
  xor_4  g0309(.A(pi87), .B(pi85), .Y(new_n585));
  nand_5 g0310(.A(pi62), .B(pi30), .Y(new_n586));
  nand_5 g0311(.A(pi71), .B(pi19), .Y(new_n587));
  xor_4  g0312(.A(pi71), .B(pi19), .Y(new_n588));
  or_6   g0313(.A(pi56), .B(pi43), .Y(new_n589));
  nand_5 g0314(.A(pi63), .B(pi40), .Y(new_n590));
  xor_4  g0315(.A(pi56), .B(pi43), .Y(new_n591));
  nand_5 g0316(.A(new_n591), .B(new_n590), .Y(new_n592));
  nand_5 g0317(.A(new_n592), .B(new_n589), .Y(new_n593));
  not_8  g0318(.A(new_n593), .Y(new_n594));
  nand_5 g0319(.A(new_n594), .B(new_n588), .Y(new_n595));
  nand_5 g0320(.A(new_n595), .B(new_n587), .Y(new_n596));
  xor_4  g0321(.A(pi62), .B(pi30), .Y(new_n597));
  nand_5 g0322(.A(new_n597), .B(new_n596), .Y(new_n598));
  nand_5 g0323(.A(new_n598), .B(new_n586), .Y(new_n599));
  nand_5 g0324(.A(new_n599), .B(new_n585), .Y(new_n600));
  nand_5 g0325(.A(new_n600), .B(new_n584), .Y(new_n601));
  nand_5 g0326(.A(new_n601), .B(pi69), .Y(new_n602));
  nor_5  g0327(.A(new_n602), .B(new_n583), .Y(new_n603));
  xor_4  g0328(.A(new_n603), .B(pi81), .Y(new_n604));
  xor_4  g0329(.A(new_n604), .B(new_n582), .Y(new_n605));
  xor_4  g0330(.A(new_n573), .B(new_n566), .Y(new_n606));
  xor_4  g0331(.A(new_n602), .B(new_n583), .Y(new_n607));
  nand_5 g0332(.A(new_n607), .B(new_n606), .Y(new_n608));
  xor_4  g0333(.A(new_n607), .B(new_n606), .Y(new_n609));
  xor_4  g0334(.A(new_n565), .B(new_n559), .Y(new_n610));
  xor_4  g0335(.A(new_n601), .B(pi69), .Y(new_n611));
  nand_5 g0336(.A(new_n611), .B(new_n610), .Y(new_n612));
  xor_4  g0337(.A(new_n558), .B(new_n536), .Y(new_n613));
  xor_4  g0338(.A(new_n599), .B(new_n585), .Y(new_n614));
  nand_5 g0339(.A(new_n614), .B(new_n613), .Y(new_n615));
  xor_4  g0340(.A(new_n614), .B(new_n613), .Y(new_n616));
  xor_4  g0341(.A(new_n597), .B(new_n596), .Y(new_n617));
  xor_4  g0342(.A(new_n553), .B(new_n542), .Y(new_n618));
  not_8  g0343(.A(new_n618), .Y(new_n619));
  not_8  g0344(.A(new_n591), .Y(new_n620));
  xor_4  g0345(.A(new_n549), .B(pi48), .Y(new_n621));
  xor_4  g0346(.A(pi63), .B(pi40), .Y(new_n622));
  nand_5 g0347(.A(new_n622), .B(new_n621), .Y(new_n623));
  nor_5  g0348(.A(new_n623), .B(new_n620), .Y(new_n624));
  xor_4  g0349(.A(new_n551), .B(new_n550), .Y(new_n625));
  xor_4  g0350(.A(new_n591), .B(new_n590), .Y(new_n626));
  and_6  g0351(.A(new_n626), .B(new_n623), .Y(new_n627));
  or_6   g0352(.A(new_n627), .B(new_n624), .Y(new_n628));
  nor_5  g0353(.A(new_n628), .B(new_n625), .Y(new_n629));
  nor_5  g0354(.A(new_n629), .B(new_n624), .Y(new_n630));
  nand_5 g0355(.A(new_n630), .B(new_n619), .Y(new_n631));
  xor_4  g0356(.A(new_n594), .B(new_n588), .Y(new_n632));
  not_8  g0357(.A(new_n632), .Y(new_n633));
  xor_4  g0358(.A(new_n630), .B(new_n619), .Y(new_n634));
  nand_5 g0359(.A(new_n634), .B(new_n633), .Y(new_n635));
  nand_5 g0360(.A(new_n635), .B(new_n631), .Y(new_n636));
  not_8  g0361(.A(new_n636), .Y(new_n637));
  nor_5  g0362(.A(new_n637), .B(new_n617), .Y(new_n638));
  xor_4  g0363(.A(new_n556), .B(new_n555), .Y(new_n639));
  xor_4  g0364(.A(new_n637), .B(new_n617), .Y(new_n640));
  not_8  g0365(.A(new_n640), .Y(new_n641));
  nor_5  g0366(.A(new_n641), .B(new_n639), .Y(new_n642));
  nor_5  g0367(.A(new_n642), .B(new_n638), .Y(new_n643));
  nand_5 g0368(.A(new_n643), .B(new_n616), .Y(new_n644));
  nand_5 g0369(.A(new_n644), .B(new_n615), .Y(new_n645));
  xor_4  g0370(.A(new_n611), .B(new_n610), .Y(new_n646));
  nand_5 g0371(.A(new_n646), .B(new_n645), .Y(new_n647));
  nand_5 g0372(.A(new_n647), .B(new_n612), .Y(new_n648));
  nand_5 g0373(.A(new_n648), .B(new_n609), .Y(new_n649));
  nand_5 g0374(.A(new_n649), .B(new_n608), .Y(new_n650));
  xor_4  g0375(.A(new_n650), .B(new_n605), .Y(po004));
  or_6   g0376(.A(new_n581), .B(new_n574), .Y(new_n652));
  or_6   g0377(.A(new_n580), .B(new_n575), .Y(new_n653));
  or_6   g0378(.A(new_n576), .B(pi78), .Y(new_n654));
  nand_5 g0379(.A(new_n654), .B(pi20), .Y(new_n655));
  not_8  g0380(.A(new_n489), .Y(new_n656));
  nand_5 g0381(.A(new_n656), .B(new_n561), .Y(new_n657));
  nand_5 g0382(.A(new_n657), .B(new_n655), .Y(new_n658));
  nand_5 g0383(.A(new_n658), .B(new_n522), .Y(new_n659));
  nand_5 g0384(.A(pi84), .B(pi14), .Y(new_n660));
  nand_5 g0385(.A(new_n660), .B(new_n659), .Y(new_n661));
  xor_4  g0386(.A(new_n661), .B(new_n653), .Y(new_n662));
  nor_5  g0387(.A(new_n662), .B(new_n652), .Y(new_n663));
  not_8  g0388(.A(new_n663), .Y(new_n664));
  nor_5  g0389(.A(new_n661), .B(new_n653), .Y(new_n665));
  not_8  g0390(.A(pi09), .Y(new_n666));
  nand_5 g0391(.A(pi14), .B(new_n666), .Y(new_n667));
  nand_5 g0392(.A(new_n657), .B(pi66), .Y(new_n668));
  nand_5 g0393(.A(new_n668), .B(new_n522), .Y(new_n669));
  not_8  g0394(.A(new_n669), .Y(new_n670));
  or_6   g0395(.A(new_n657), .B(pi66), .Y(new_n671));
  nand_5 g0396(.A(new_n671), .B(new_n670), .Y(new_n672));
  nand_5 g0397(.A(new_n672), .B(new_n667), .Y(new_n673));
  xor_4  g0398(.A(new_n673), .B(new_n665), .Y(new_n674));
  nor_5  g0399(.A(new_n674), .B(new_n664), .Y(new_n675));
  not_8  g0400(.A(new_n675), .Y(new_n676));
  nand_5 g0401(.A(new_n673), .B(new_n665), .Y(new_n677));
  nand_5 g0402(.A(new_n671), .B(pi74), .Y(new_n678));
  not_8  g0403(.A(pi74), .Y(new_n679));
  not_8  g0404(.A(pi66), .Y(new_n680));
  nand_5 g0405(.A(new_n656), .B(new_n680), .Y(new_n681));
  not_8  g0406(.A(new_n681), .Y(new_n682));
  nand_5 g0407(.A(new_n682), .B(new_n679), .Y(new_n683));
  not_8  g0408(.A(new_n683), .Y(new_n684));
  nand_5 g0409(.A(new_n684), .B(new_n561), .Y(new_n685));
  nand_5 g0410(.A(new_n685), .B(new_n678), .Y(new_n686));
  nand_5 g0411(.A(new_n686), .B(new_n522), .Y(new_n687));
  nand_5 g0412(.A(pi31), .B(pi14), .Y(new_n688));
  nand_5 g0413(.A(new_n688), .B(new_n687), .Y(new_n689));
  xor_4  g0414(.A(new_n689), .B(new_n677), .Y(new_n690));
  xor_4  g0415(.A(new_n690), .B(new_n676), .Y(new_n691));
  xor_4  g0416(.A(new_n674), .B(new_n664), .Y(new_n692));
  not_8  g0417(.A(pi35), .Y(new_n693));
  nand_5 g0418(.A(new_n603), .B(pi81), .Y(new_n694));
  nor_5  g0419(.A(new_n694), .B(new_n693), .Y(new_n695));
  nand_5 g0420(.A(new_n695), .B(new_n692), .Y(new_n696));
  xor_4  g0421(.A(new_n662), .B(new_n652), .Y(new_n697));
  xor_4  g0422(.A(new_n694), .B(new_n693), .Y(new_n698));
  nand_5 g0423(.A(new_n698), .B(new_n697), .Y(new_n699));
  xor_4  g0424(.A(new_n698), .B(new_n697), .Y(new_n700));
  nand_5 g0425(.A(new_n604), .B(new_n582), .Y(new_n701));
  nand_5 g0426(.A(new_n650), .B(new_n605), .Y(new_n702));
  nand_5 g0427(.A(new_n702), .B(new_n701), .Y(new_n703));
  nand_5 g0428(.A(new_n703), .B(new_n700), .Y(new_n704));
  nand_5 g0429(.A(new_n704), .B(new_n699), .Y(new_n705));
  xor_4  g0430(.A(new_n695), .B(new_n692), .Y(new_n706));
  nand_5 g0431(.A(new_n706), .B(new_n705), .Y(new_n707));
  nand_5 g0432(.A(new_n707), .B(new_n696), .Y(new_n708));
  xor_4  g0433(.A(new_n708), .B(new_n691), .Y(po005));
  xor_4  g0434(.A(pi85), .B(pi27), .Y(new_n710));
  nand_5 g0435(.A(pi54), .B(pi30), .Y(new_n711));
  nand_5 g0436(.A(pi37), .B(pi19), .Y(new_n712));
  xor_4  g0437(.A(pi37), .B(pi19), .Y(new_n713));
  or_6   g0438(.A(pi56), .B(pi36), .Y(new_n714));
  nand_5 g0439(.A(pi92), .B(pi63), .Y(new_n715));
  xor_4  g0440(.A(pi56), .B(pi36), .Y(new_n716));
  nand_5 g0441(.A(new_n716), .B(new_n715), .Y(new_n717));
  nand_5 g0442(.A(new_n717), .B(new_n714), .Y(new_n718));
  not_8  g0443(.A(new_n718), .Y(new_n719));
  nand_5 g0444(.A(new_n719), .B(new_n713), .Y(new_n720));
  nand_5 g0445(.A(new_n720), .B(new_n712), .Y(new_n721));
  xor_4  g0446(.A(pi54), .B(pi30), .Y(new_n722));
  nand_5 g0447(.A(new_n722), .B(new_n721), .Y(new_n723));
  nand_5 g0448(.A(new_n723), .B(new_n711), .Y(new_n724));
  xor_4  g0449(.A(new_n724), .B(new_n710), .Y(new_n725));
  xor_4  g0450(.A(new_n725), .B(new_n360), .Y(new_n726));
  xor_4  g0451(.A(new_n722), .B(new_n721), .Y(new_n727));
  nand_5 g0452(.A(new_n727), .B(new_n363), .Y(new_n728));
  xnor_4 g0453(.A(new_n727), .B(new_n363), .Y(new_n729));
  xor_4  g0454(.A(new_n718), .B(new_n713), .Y(new_n730));
  not_8  g0455(.A(new_n716), .Y(new_n731));
  xor_4  g0456(.A(pi92), .B(pi63), .Y(new_n732));
  nand_5 g0457(.A(new_n732), .B(new_n375), .Y(new_n733));
  nor_5  g0458(.A(new_n733), .B(new_n731), .Y(new_n734));
  xor_4  g0459(.A(new_n716), .B(new_n715), .Y(new_n735));
  and_6  g0460(.A(new_n735), .B(new_n733), .Y(new_n736));
  or_6   g0461(.A(new_n736), .B(new_n734), .Y(new_n737));
  nor_5  g0462(.A(new_n737), .B(new_n383), .Y(new_n738));
  nor_5  g0463(.A(new_n738), .B(new_n734), .Y(new_n739));
  nand_5 g0464(.A(new_n739), .B(new_n730), .Y(new_n740));
  xor_4  g0465(.A(new_n739), .B(new_n730), .Y(new_n741));
  nand_5 g0466(.A(new_n741), .B(new_n369), .Y(new_n742));
  nand_5 g0467(.A(new_n742), .B(new_n740), .Y(new_n743));
  or_6   g0468(.A(new_n743), .B(new_n729), .Y(new_n744));
  nand_5 g0469(.A(new_n744), .B(new_n728), .Y(new_n745));
  xor_4  g0470(.A(new_n745), .B(new_n726), .Y(po006));
  nor_5  g0471(.A(new_n496), .B(new_n483), .Y(new_n747));
  nor_5  g0472(.A(new_n484), .B(pi84), .Y(new_n748));
  xor_4  g0473(.A(new_n748), .B(pi09), .Y(new_n749));
  nand_5 g0474(.A(new_n749), .B(pi73), .Y(new_n750));
  nand_5 g0475(.A(new_n489), .B(pi66), .Y(new_n751));
  nor_5  g0476(.A(new_n682), .B(new_n450), .Y(new_n752));
  nand_5 g0477(.A(new_n752), .B(new_n751), .Y(new_n753));
  nor_5  g0478(.A(pi22), .B(pi09), .Y(new_n754));
  nor_5  g0479(.A(new_n754), .B(pi73), .Y(new_n755));
  nand_5 g0480(.A(new_n755), .B(new_n753), .Y(new_n756));
  nand_5 g0481(.A(new_n756), .B(new_n750), .Y(new_n757));
  xor_4  g0482(.A(new_n757), .B(new_n747), .Y(po111));
  nand_5 g0483(.A(po111), .B(new_n519), .Y(new_n759));
  not_8  g0484(.A(new_n759), .Y(new_n760));
  nand_5 g0485(.A(new_n757), .B(new_n747), .Y(new_n761));
  nand_5 g0486(.A(new_n748), .B(new_n666), .Y(new_n762));
  xor_4  g0487(.A(new_n762), .B(pi31), .Y(new_n763));
  nor_5  g0488(.A(new_n763), .B(new_n396), .Y(new_n764));
  nand_5 g0489(.A(new_n681), .B(pi74), .Y(new_n765));
  not_8  g0490(.A(new_n765), .Y(new_n766));
  nand_5 g0491(.A(new_n683), .B(pi22), .Y(new_n767));
  nor_5  g0492(.A(new_n767), .B(new_n766), .Y(new_n768));
  not_8  g0493(.A(pi31), .Y(new_n769));
  nand_5 g0494(.A(new_n769), .B(new_n450), .Y(new_n770));
  nand_5 g0495(.A(new_n770), .B(new_n396), .Y(new_n771));
  nor_5  g0496(.A(new_n771), .B(new_n768), .Y(new_n772));
  nor_5  g0497(.A(new_n772), .B(new_n764), .Y(new_n773));
  xor_4  g0498(.A(new_n773), .B(new_n761), .Y(po011));
  nor_5  g0499(.A(po011), .B(new_n760), .Y(new_n775));
  not_8  g0500(.A(new_n773), .Y(new_n776));
  nand_5 g0501(.A(new_n776), .B(new_n760), .Y(new_n777));
  not_8  g0502(.A(new_n777), .Y(new_n778));
  nor_5  g0503(.A(new_n778), .B(new_n775), .Y(po007));
  xor_4  g0504(.A(new_n465), .B(new_n458), .Y(po140));
  nor_5  g0505(.A(po140), .B(new_n513), .Y(new_n781));
  nor_5  g0506(.A(new_n781), .B(new_n515), .Y(po008));
  xor_4  g0507(.A(new_n643), .B(new_n616), .Y(po009));
  nand_5 g0508(.A(new_n534), .B(pi85), .Y(new_n784));
  xor_4  g0509(.A(new_n534), .B(pi85), .Y(new_n785));
  nand_5 g0510(.A(new_n529), .B(pi30), .Y(new_n786));
  nand_5 g0511(.A(new_n525), .B(pi19), .Y(new_n787));
  xor_4  g0512(.A(new_n526), .B(pi19), .Y(new_n788));
  or_6   g0513(.A(new_n545), .B(pi56), .Y(new_n789));
  nand_5 g0514(.A(new_n549), .B(pi63), .Y(new_n790));
  xor_4  g0515(.A(new_n545), .B(pi56), .Y(new_n791));
  nand_5 g0516(.A(new_n791), .B(new_n790), .Y(new_n792));
  nand_5 g0517(.A(new_n792), .B(new_n789), .Y(new_n793));
  or_6   g0518(.A(new_n793), .B(new_n788), .Y(new_n794));
  nand_5 g0519(.A(new_n794), .B(new_n787), .Y(new_n795));
  xor_4  g0520(.A(new_n529), .B(pi30), .Y(new_n796));
  nand_5 g0521(.A(new_n796), .B(new_n795), .Y(new_n797));
  nand_5 g0522(.A(new_n797), .B(new_n786), .Y(new_n798));
  nand_5 g0523(.A(new_n798), .B(new_n785), .Y(new_n799));
  nand_5 g0524(.A(new_n799), .B(new_n784), .Y(new_n800));
  nand_5 g0525(.A(new_n800), .B(new_n564), .Y(new_n801));
  xor_4  g0526(.A(new_n801), .B(new_n572), .Y(po010));
  xor_4  g0527(.A(new_n376), .B(pi18), .Y(po012));
  not_8  g0528(.A(pi75), .Y(new_n804));
  not_8  g0529(.A(pi06), .Y(new_n805));
  not_8  g0530(.A(pi59), .Y(new_n806));
  nand_5 g0531(.A(new_n376), .B(pi18), .Y(new_n807));
  nor_5  g0532(.A(new_n807), .B(new_n806), .Y(new_n808));
  not_8  g0533(.A(new_n379), .Y(new_n809));
  xor_4  g0534(.A(new_n807), .B(new_n806), .Y(new_n810));
  and_6  g0535(.A(new_n810), .B(new_n809), .Y(new_n811));
  nor_5  g0536(.A(new_n811), .B(new_n808), .Y(new_n812));
  nand_5 g0537(.A(new_n812), .B(new_n805), .Y(new_n813));
  xor_4  g0538(.A(new_n812), .B(new_n805), .Y(new_n814));
  nand_5 g0539(.A(new_n814), .B(new_n371), .Y(new_n815));
  nand_5 g0540(.A(new_n815), .B(new_n813), .Y(new_n816));
  nand_5 g0541(.A(new_n816), .B(new_n804), .Y(new_n817));
  xor_4  g0542(.A(new_n816), .B(new_n804), .Y(new_n818));
  nand_5 g0543(.A(new_n818), .B(new_n366), .Y(new_n819));
  and_6  g0544(.A(new_n819), .B(new_n817), .Y(new_n820));
  or_6   g0545(.A(new_n820), .B(new_n361), .Y(new_n821));
  not_8  g0546(.A(pi39), .Y(new_n822));
  xor_4  g0547(.A(new_n820), .B(new_n361), .Y(new_n823));
  nand_5 g0548(.A(new_n823), .B(new_n822), .Y(new_n824));
  nand_5 g0549(.A(new_n824), .B(new_n821), .Y(new_n825));
  xor_4  g0550(.A(new_n357), .B(pi82), .Y(new_n826));
  xor_4  g0551(.A(new_n826), .B(new_n825), .Y(new_n827));
  xor_4  g0552(.A(new_n814), .B(new_n371), .Y(po047));
  xor_4  g0553(.A(new_n823), .B(new_n822), .Y(new_n829));
  xor_4  g0554(.A(new_n818), .B(new_n366), .Y(po162));
  nand_5 g0555(.A(po162), .B(new_n829), .Y(new_n831));
  not_8  g0556(.A(new_n831), .Y(new_n832));
  nand_5 g0557(.A(new_n832), .B(po047), .Y(new_n833));
  xor_4  g0558(.A(new_n833), .B(new_n827), .Y(po013));
  xnor_4 g0559(.A(new_n385), .B(new_n373), .Y(po014));
  nand_5 g0560(.A(pi85), .B(pi24), .Y(new_n836));
  xor_4  g0561(.A(pi85), .B(pi24), .Y(new_n837));
  nand_5 g0562(.A(pi72), .B(pi30), .Y(new_n838));
  nand_5 g0563(.A(pi29), .B(pi19), .Y(new_n839));
  xor_4  g0564(.A(pi29), .B(pi19), .Y(new_n840));
  or_6   g0565(.A(pi56), .B(pi23), .Y(new_n841));
  nand_5 g0566(.A(pi63), .B(pi10), .Y(new_n842));
  xor_4  g0567(.A(pi56), .B(pi23), .Y(new_n843));
  nand_5 g0568(.A(new_n843), .B(new_n842), .Y(new_n844));
  nand_5 g0569(.A(new_n844), .B(new_n841), .Y(new_n845));
  not_8  g0570(.A(new_n845), .Y(new_n846));
  nand_5 g0571(.A(new_n846), .B(new_n840), .Y(new_n847));
  nand_5 g0572(.A(new_n847), .B(new_n839), .Y(new_n848));
  xor_4  g0573(.A(pi72), .B(pi30), .Y(new_n849));
  nand_5 g0574(.A(new_n849), .B(new_n848), .Y(new_n850));
  nand_5 g0575(.A(new_n850), .B(new_n838), .Y(new_n851));
  nand_5 g0576(.A(new_n851), .B(new_n837), .Y(new_n852));
  nand_5 g0577(.A(new_n852), .B(new_n836), .Y(new_n853));
  xor_4  g0578(.A(new_n853), .B(pi01), .Y(new_n854));
  not_8  g0579(.A(new_n534), .Y(new_n855));
  nand_5 g0580(.A(new_n525), .B(pi11), .Y(new_n856));
  not_8  g0581(.A(new_n856), .Y(new_n857));
  xor_4  g0582(.A(new_n525), .B(pi11), .Y(new_n858));
  not_8  g0583(.A(new_n858), .Y(new_n859));
  or_6   g0584(.A(new_n545), .B(pi88), .Y(new_n860));
  nand_5 g0585(.A(new_n549), .B(pi33), .Y(new_n861));
  xor_4  g0586(.A(new_n545), .B(pi88), .Y(new_n862));
  nand_5 g0587(.A(new_n862), .B(new_n861), .Y(new_n863));
  nand_5 g0588(.A(new_n863), .B(new_n860), .Y(new_n864));
  nor_5  g0589(.A(new_n864), .B(new_n859), .Y(new_n865));
  nor_5  g0590(.A(new_n865), .B(new_n857), .Y(new_n866));
  not_8  g0591(.A(new_n866), .Y(new_n867));
  nand_5 g0592(.A(new_n867), .B(new_n529), .Y(new_n868));
  or_6   g0593(.A(new_n868), .B(new_n855), .Y(new_n869));
  not_8  g0594(.A(new_n869), .Y(new_n870));
  xor_4  g0595(.A(new_n870), .B(new_n564), .Y(new_n871));
  xor_4  g0596(.A(new_n871), .B(new_n854), .Y(new_n872));
  xor_4  g0597(.A(new_n868), .B(new_n855), .Y(new_n873));
  xor_4  g0598(.A(new_n851), .B(new_n837), .Y(new_n874));
  nand_5 g0599(.A(new_n874), .B(new_n873), .Y(new_n875));
  xor_4  g0600(.A(new_n874), .B(new_n873), .Y(new_n876));
  xor_4  g0601(.A(new_n866), .B(new_n530), .Y(new_n877));
  xor_4  g0602(.A(new_n849), .B(new_n848), .Y(new_n878));
  nand_5 g0603(.A(new_n878), .B(new_n877), .Y(new_n879));
  not_8  g0604(.A(new_n879), .Y(new_n880));
  xnor_4 g0605(.A(new_n878), .B(new_n877), .Y(new_n881));
  xor_4  g0606(.A(new_n864), .B(new_n859), .Y(new_n882));
  not_8  g0607(.A(new_n882), .Y(new_n883));
  xor_4  g0608(.A(new_n845), .B(new_n840), .Y(new_n884));
  nor_5  g0609(.A(new_n884), .B(new_n883), .Y(new_n885));
  not_8  g0610(.A(new_n843), .Y(new_n886));
  xor_4  g0611(.A(new_n549), .B(pi33), .Y(new_n887));
  xor_4  g0612(.A(pi63), .B(pi10), .Y(new_n888));
  nand_5 g0613(.A(new_n888), .B(new_n887), .Y(new_n889));
  nor_5  g0614(.A(new_n889), .B(new_n886), .Y(new_n890));
  xor_4  g0615(.A(new_n862), .B(new_n861), .Y(new_n891));
  xor_4  g0616(.A(new_n843), .B(new_n842), .Y(new_n892));
  and_6  g0617(.A(new_n892), .B(new_n889), .Y(new_n893));
  or_6   g0618(.A(new_n893), .B(new_n890), .Y(new_n894));
  nor_5  g0619(.A(new_n894), .B(new_n891), .Y(new_n895));
  nor_5  g0620(.A(new_n895), .B(new_n890), .Y(new_n896));
  not_8  g0621(.A(new_n896), .Y(new_n897));
  xor_4  g0622(.A(new_n884), .B(new_n883), .Y(new_n898));
  and_6  g0623(.A(new_n898), .B(new_n897), .Y(new_n899));
  nor_5  g0624(.A(new_n899), .B(new_n885), .Y(new_n900));
  nor_5  g0625(.A(new_n900), .B(new_n881), .Y(new_n901));
  nor_5  g0626(.A(new_n901), .B(new_n880), .Y(new_n902));
  not_8  g0627(.A(new_n902), .Y(new_n903));
  nand_5 g0628(.A(new_n903), .B(new_n876), .Y(new_n904));
  nand_5 g0629(.A(new_n904), .B(new_n875), .Y(new_n905));
  xor_4  g0630(.A(new_n905), .B(new_n872), .Y(po015));
  xor_4  g0631(.A(new_n898), .B(new_n897), .Y(po016));
  xor_4  g0632(.A(new_n706), .B(new_n705), .Y(po017));
  not_8  g0633(.A(new_n661), .Y(new_n909));
  not_8  g0634(.A(new_n572), .Y(new_n910));
  nand_5 g0635(.A(new_n870), .B(new_n564), .Y(new_n911));
  not_8  g0636(.A(new_n911), .Y(new_n912));
  nand_5 g0637(.A(new_n912), .B(new_n910), .Y(new_n913));
  not_8  g0638(.A(new_n913), .Y(new_n914));
  nand_5 g0639(.A(new_n914), .B(new_n580), .Y(new_n915));
  xor_4  g0640(.A(new_n915), .B(new_n909), .Y(new_n916));
  not_8  g0641(.A(pi89), .Y(new_n917));
  not_8  g0642(.A(pi58), .Y(new_n918));
  nand_5 g0643(.A(new_n853), .B(pi01), .Y(new_n919));
  nor_5  g0644(.A(new_n919), .B(new_n918), .Y(new_n920));
  nand_5 g0645(.A(new_n920), .B(pi44), .Y(new_n921));
  xor_4  g0646(.A(new_n921), .B(new_n917), .Y(new_n922));
  xnor_4 g0647(.A(new_n922), .B(new_n916), .Y(new_n923));
  not_8  g0648(.A(new_n580), .Y(new_n924));
  xor_4  g0649(.A(new_n913), .B(new_n924), .Y(new_n925));
  xor_4  g0650(.A(new_n920), .B(pi44), .Y(new_n926));
  and_6  g0651(.A(new_n926), .B(new_n925), .Y(new_n927));
  xnor_4 g0652(.A(new_n926), .B(new_n925), .Y(new_n928));
  xor_4  g0653(.A(new_n911), .B(new_n572), .Y(new_n929));
  xor_4  g0654(.A(new_n919), .B(new_n918), .Y(new_n930));
  or_6   g0655(.A(new_n930), .B(new_n929), .Y(new_n931));
  nand_5 g0656(.A(new_n871), .B(new_n854), .Y(new_n932));
  nand_5 g0657(.A(new_n905), .B(new_n872), .Y(new_n933));
  nand_5 g0658(.A(new_n933), .B(new_n932), .Y(new_n934));
  not_8  g0659(.A(new_n934), .Y(new_n935));
  xor_4  g0660(.A(new_n930), .B(new_n929), .Y(new_n936));
  nand_5 g0661(.A(new_n936), .B(new_n935), .Y(new_n937));
  nand_5 g0662(.A(new_n937), .B(new_n931), .Y(new_n938));
  nor_5  g0663(.A(new_n938), .B(new_n928), .Y(new_n939));
  nor_5  g0664(.A(new_n939), .B(new_n927), .Y(new_n940));
  xor_4  g0665(.A(new_n940), .B(new_n923), .Y(po018));
  not_8  g0666(.A(pi38), .Y(new_n942));
  nor_5  g0667(.A(new_n353), .B(new_n334), .Y(new_n943));
  nand_5 g0668(.A(new_n943), .B(pi80), .Y(new_n944));
  nor_5  g0669(.A(new_n944), .B(new_n942), .Y(new_n945));
  xor_4  g0670(.A(new_n945), .B(pi66), .Y(new_n946));
  xor_4  g0671(.A(new_n944), .B(new_n942), .Y(new_n947));
  not_8  g0672(.A(new_n947), .Y(new_n948));
  nand_5 g0673(.A(new_n948), .B(new_n487), .Y(new_n949));
  xor_4  g0674(.A(new_n943), .B(pi80), .Y(new_n950));
  or_6   g0675(.A(new_n950), .B(pi78), .Y(new_n951));
  xor_4  g0676(.A(new_n950), .B(pi78), .Y(new_n952));
  or_6   g0677(.A(new_n354), .B(pi04), .Y(new_n953));
  not_8  g0678(.A(new_n357), .Y(new_n954));
  nand_5 g0679(.A(new_n954), .B(new_n561), .Y(new_n955));
  nand_5 g0680(.A(new_n826), .B(new_n825), .Y(new_n956));
  nand_5 g0681(.A(new_n956), .B(new_n955), .Y(new_n957));
  xor_4  g0682(.A(new_n354), .B(pi04), .Y(new_n958));
  nand_5 g0683(.A(new_n958), .B(new_n957), .Y(new_n959));
  nand_5 g0684(.A(new_n959), .B(new_n953), .Y(new_n960));
  nand_5 g0685(.A(new_n960), .B(new_n952), .Y(new_n961));
  nand_5 g0686(.A(new_n961), .B(new_n951), .Y(new_n962));
  xor_4  g0687(.A(new_n947), .B(pi20), .Y(new_n963));
  nand_5 g0688(.A(new_n963), .B(new_n962), .Y(new_n964));
  nand_5 g0689(.A(new_n964), .B(new_n949), .Y(new_n965));
  xor_4  g0690(.A(new_n965), .B(new_n946), .Y(new_n966));
  xor_4  g0691(.A(new_n963), .B(new_n962), .Y(new_n967));
  xor_4  g0692(.A(new_n960), .B(new_n952), .Y(new_n968));
  nand_5 g0693(.A(new_n832), .B(new_n827), .Y(new_n969));
  xor_4  g0694(.A(new_n958), .B(new_n957), .Y(new_n970));
  not_8  g0695(.A(new_n970), .Y(new_n971));
  nor_5  g0696(.A(new_n971), .B(new_n969), .Y(new_n972));
  nand_5 g0697(.A(new_n972), .B(new_n968), .Y(new_n973));
  not_8  g0698(.A(new_n973), .Y(new_n974));
  nand_5 g0699(.A(new_n974), .B(new_n967), .Y(new_n975));
  not_8  g0700(.A(new_n975), .Y(new_n976));
  nand_5 g0701(.A(new_n976), .B(po047), .Y(new_n977));
  xor_4  g0702(.A(new_n977), .B(new_n966), .Y(po019));
  xnor_4 g0703(.A(new_n613), .B(new_n361), .Y(new_n979));
  nand_5 g0704(.A(new_n621), .B(new_n376), .Y(new_n980));
  or_6   g0705(.A(new_n980), .B(new_n374), .Y(new_n981));
  nand_5 g0706(.A(new_n980), .B(new_n379), .Y(new_n982));
  nand_5 g0707(.A(new_n982), .B(new_n981), .Y(new_n983));
  or_6   g0708(.A(new_n983), .B(new_n625), .Y(new_n984));
  nand_5 g0709(.A(new_n984), .B(new_n981), .Y(new_n985));
  nor_5  g0710(.A(new_n985), .B(new_n618), .Y(new_n986));
  xor_4  g0711(.A(new_n985), .B(new_n618), .Y(new_n987));
  and_6  g0712(.A(new_n987), .B(new_n371), .Y(new_n988));
  nor_5  g0713(.A(new_n988), .B(new_n986), .Y(new_n989));
  or_6   g0714(.A(new_n989), .B(new_n639), .Y(new_n990));
  xor_4  g0715(.A(new_n989), .B(new_n639), .Y(new_n991));
  nand_5 g0716(.A(new_n991), .B(new_n366), .Y(new_n992));
  nand_5 g0717(.A(new_n992), .B(new_n990), .Y(new_n993));
  xor_4  g0718(.A(new_n993), .B(new_n979), .Y(po020));
  xor_4  g0719(.A(new_n732), .B(new_n375), .Y(po021));
  xor_4  g0720(.A(new_n810), .B(new_n809), .Y(po022));
  or_6   g0721(.A(new_n915), .B(new_n909), .Y(new_n997));
  nor_5  g0722(.A(new_n997), .B(new_n673), .Y(new_n998));
  xor_4  g0723(.A(new_n998), .B(new_n689), .Y(new_n999));
  nor_5  g0724(.A(new_n921), .B(new_n917), .Y(new_n1000));
  xor_4  g0725(.A(new_n997), .B(new_n673), .Y(new_n1001));
  nor_5  g0726(.A(new_n1001), .B(new_n1000), .Y(new_n1002));
  nand_5 g0727(.A(new_n1001), .B(new_n1000), .Y(new_n1003));
  nand_5 g0728(.A(new_n922), .B(new_n916), .Y(new_n1004));
  not_8  g0729(.A(new_n1004), .Y(new_n1005));
  nor_5  g0730(.A(new_n940), .B(new_n923), .Y(new_n1006));
  nor_5  g0731(.A(new_n1006), .B(new_n1005), .Y(new_n1007));
  nand_5 g0732(.A(new_n1007), .B(new_n1003), .Y(new_n1008));
  not_8  g0733(.A(new_n1008), .Y(new_n1009));
  nor_5  g0734(.A(new_n1009), .B(new_n1002), .Y(new_n1010));
  nand_5 g0735(.A(new_n1010), .B(new_n999), .Y(new_n1011));
  not_8  g0736(.A(new_n1011), .Y(new_n1012));
  nor_5  g0737(.A(new_n685), .B(new_n669), .Y(new_n1013));
  not_8  g0738(.A(new_n1013), .Y(new_n1014));
  or_6   g0739(.A(new_n1014), .B(new_n998), .Y(new_n1015));
  nor_5  g0740(.A(new_n1015), .B(new_n1012), .Y(po023));
  nand_5 g0741(.A(new_n432), .B(pi70), .Y(new_n1017));
  nand_5 g0742(.A(new_n401), .B(pi07), .Y(new_n1018));
  nand_5 g0743(.A(new_n413), .B(new_n402), .Y(new_n1019));
  nand_5 g0744(.A(new_n1019), .B(new_n1018), .Y(new_n1020));
  xor_4  g0745(.A(new_n432), .B(pi70), .Y(new_n1021));
  nand_5 g0746(.A(new_n1021), .B(new_n1020), .Y(new_n1022));
  nand_5 g0747(.A(new_n1022), .B(new_n1017), .Y(new_n1023));
  nand_5 g0748(.A(new_n1023), .B(new_n427), .Y(new_n1024));
  not_8  g0749(.A(new_n1024), .Y(new_n1025));
  nand_5 g0750(.A(new_n1025), .B(new_n457), .Y(new_n1026));
  not_8  g0751(.A(new_n1026), .Y(new_n1027));
  xor_4  g0752(.A(new_n1027), .B(new_n465), .Y(new_n1028));
  not_8  g0753(.A(pi65), .Y(new_n1029));
  nand_5 g0754(.A(pi85), .B(pi46), .Y(new_n1030));
  xor_4  g0755(.A(pi85), .B(pi46), .Y(new_n1031));
  nand_5 g0756(.A(pi64), .B(pi30), .Y(new_n1032));
  nand_5 g0757(.A(pi42), .B(pi19), .Y(new_n1033));
  xor_4  g0758(.A(pi42), .B(pi19), .Y(new_n1034));
  nor_5  g0759(.A(pi67), .B(pi56), .Y(new_n1035));
  nand_5 g0760(.A(pi63), .B(pi61), .Y(new_n1036));
  xor_4  g0761(.A(pi67), .B(pi56), .Y(new_n1037));
  nand_5 g0762(.A(new_n1037), .B(new_n1036), .Y(new_n1038));
  not_8  g0763(.A(new_n1038), .Y(new_n1039));
  nor_5  g0764(.A(new_n1039), .B(new_n1035), .Y(new_n1040));
  nand_5 g0765(.A(new_n1040), .B(new_n1034), .Y(new_n1041));
  nand_5 g0766(.A(new_n1041), .B(new_n1033), .Y(new_n1042));
  xor_4  g0767(.A(pi64), .B(pi30), .Y(new_n1043));
  nand_5 g0768(.A(new_n1043), .B(new_n1042), .Y(new_n1044));
  nand_5 g0769(.A(new_n1044), .B(new_n1032), .Y(new_n1045));
  nand_5 g0770(.A(new_n1045), .B(new_n1031), .Y(new_n1046));
  nand_5 g0771(.A(new_n1046), .B(new_n1030), .Y(new_n1047));
  nand_5 g0772(.A(new_n1047), .B(pi50), .Y(new_n1048));
  xor_4  g0773(.A(new_n1048), .B(new_n1029), .Y(new_n1049));
  xor_4  g0774(.A(new_n1049), .B(new_n1028), .Y(new_n1050));
  xor_4  g0775(.A(new_n1024), .B(new_n457), .Y(new_n1051));
  xor_4  g0776(.A(new_n1047), .B(pi50), .Y(new_n1052));
  not_8  g0777(.A(new_n1052), .Y(new_n1053));
  nor_5  g0778(.A(new_n1053), .B(new_n1051), .Y(new_n1054));
  xor_4  g0779(.A(new_n1053), .B(new_n1051), .Y(new_n1055));
  xor_4  g0780(.A(new_n1023), .B(new_n427), .Y(new_n1056));
  xor_4  g0781(.A(new_n1045), .B(new_n1031), .Y(new_n1057));
  nand_5 g0782(.A(new_n1057), .B(new_n1056), .Y(new_n1058));
  xor_4  g0783(.A(new_n1057), .B(new_n1056), .Y(new_n1059));
  xor_4  g0784(.A(new_n1021), .B(new_n1020), .Y(new_n1060));
  xor_4  g0785(.A(new_n1043), .B(new_n1042), .Y(new_n1061));
  nand_5 g0786(.A(new_n1061), .B(new_n1060), .Y(new_n1062));
  not_8  g0787(.A(new_n1060), .Y(new_n1063));
  xor_4  g0788(.A(new_n1061), .B(new_n1063), .Y(new_n1064));
  xnor_4 g0789(.A(new_n1040), .B(new_n1034), .Y(new_n1065));
  not_8  g0790(.A(new_n1037), .Y(new_n1066));
  xor_4  g0791(.A(pi63), .B(pi61), .Y(new_n1067));
  nand_5 g0792(.A(new_n1067), .B(new_n415), .Y(new_n1068));
  nor_5  g0793(.A(new_n1068), .B(new_n1066), .Y(new_n1069));
  xor_4  g0794(.A(new_n1037), .B(new_n1036), .Y(new_n1070));
  and_6  g0795(.A(new_n1070), .B(new_n1068), .Y(new_n1071));
  or_6   g0796(.A(new_n1071), .B(new_n1069), .Y(new_n1072));
  nor_5  g0797(.A(new_n1072), .B(new_n418), .Y(new_n1073));
  nor_5  g0798(.A(new_n1073), .B(new_n1069), .Y(new_n1074));
  nand_5 g0799(.A(new_n1074), .B(new_n1065), .Y(new_n1075));
  not_8  g0800(.A(new_n414), .Y(new_n1076));
  xor_4  g0801(.A(new_n1074), .B(new_n1065), .Y(new_n1077));
  nand_5 g0802(.A(new_n1077), .B(new_n1076), .Y(new_n1078));
  nand_5 g0803(.A(new_n1078), .B(new_n1075), .Y(new_n1079));
  or_6   g0804(.A(new_n1079), .B(new_n1064), .Y(new_n1080));
  nand_5 g0805(.A(new_n1080), .B(new_n1062), .Y(new_n1081));
  nand_5 g0806(.A(new_n1081), .B(new_n1059), .Y(new_n1082));
  nand_5 g0807(.A(new_n1082), .B(new_n1058), .Y(new_n1083));
  nand_5 g0808(.A(new_n1083), .B(new_n1055), .Y(new_n1084));
  not_8  g0809(.A(new_n1084), .Y(new_n1085));
  nor_5  g0810(.A(new_n1085), .B(new_n1054), .Y(new_n1086));
  not_8  g0811(.A(new_n1086), .Y(new_n1087));
  xor_4  g0812(.A(new_n1087), .B(new_n1050), .Y(po024));
  xor_4  g0813(.A(new_n1067), .B(new_n415), .Y(po025));
  xor_4  g0814(.A(new_n743), .B(new_n729), .Y(po026));
  or_6   g0815(.A(new_n801), .B(new_n572), .Y(new_n1091));
  nor_5  g0816(.A(new_n1091), .B(new_n924), .Y(new_n1092));
  nand_5 g0817(.A(new_n1092), .B(new_n661), .Y(new_n1093));
  nor_5  g0818(.A(new_n1093), .B(new_n673), .Y(new_n1094));
  nand_5 g0819(.A(new_n1094), .B(new_n689), .Y(new_n1095));
  xor_4  g0820(.A(new_n1095), .B(new_n1013), .Y(new_n1096));
  xor_4  g0821(.A(new_n1093), .B(new_n673), .Y(po124));
  xnor_4 g0822(.A(new_n791), .B(new_n790), .Y(po057));
  or_6   g0823(.A(new_n549), .B(pi63), .Y(new_n1099));
  nand_5 g0824(.A(new_n1099), .B(new_n790), .Y(po125));
  not_8  g0825(.A(po125), .Y(po058));
  nor_5  g0826(.A(po058), .B(po057), .Y(new_n1102));
  not_8  g0827(.A(new_n1102), .Y(new_n1103));
  xor_4  g0828(.A(new_n793), .B(new_n788), .Y(po100));
  or_6   g0829(.A(po100), .B(new_n1103), .Y(new_n1105));
  xor_4  g0830(.A(new_n796), .B(new_n795), .Y(po172));
  and_6  g0831(.A(po172), .B(new_n1105), .Y(new_n1107));
  xor_4  g0832(.A(new_n798), .B(new_n785), .Y(po050));
  nand_5 g0833(.A(po050), .B(new_n1107), .Y(new_n1109));
  not_8  g0834(.A(new_n1109), .Y(new_n1110));
  xor_4  g0835(.A(new_n800), .B(new_n564), .Y(po071));
  nand_5 g0836(.A(po071), .B(new_n1110), .Y(new_n1112));
  not_8  g0837(.A(new_n1112), .Y(new_n1113));
  nand_5 g0838(.A(new_n1113), .B(new_n910), .Y(new_n1114));
  not_8  g0839(.A(new_n1114), .Y(new_n1115));
  xor_4  g0840(.A(new_n1091), .B(new_n924), .Y(po107));
  nand_5 g0841(.A(po107), .B(new_n1115), .Y(new_n1117));
  not_8  g0842(.A(new_n1117), .Y(new_n1118));
  nand_5 g0843(.A(new_n1118), .B(new_n661), .Y(new_n1119));
  not_8  g0844(.A(new_n1119), .Y(new_n1120));
  and_6  g0845(.A(new_n1120), .B(po124), .Y(new_n1121));
  nand_5 g0846(.A(new_n1121), .B(new_n689), .Y(new_n1122));
  xor_4  g0847(.A(new_n1122), .B(new_n1096), .Y(po027));
  and_6  g0848(.A(new_n1027), .B(new_n465), .Y(new_n1124));
  xor_4  g0849(.A(new_n1124), .B(new_n482), .Y(new_n1125));
  nor_5  g0850(.A(new_n1048), .B(new_n1029), .Y(new_n1126));
  xor_4  g0851(.A(new_n1126), .B(pi90), .Y(new_n1127));
  xor_4  g0852(.A(new_n1127), .B(new_n1125), .Y(new_n1128));
  nand_5 g0853(.A(new_n1049), .B(new_n1028), .Y(new_n1129));
  nand_5 g0854(.A(new_n1087), .B(new_n1050), .Y(new_n1130));
  nand_5 g0855(.A(new_n1130), .B(new_n1129), .Y(new_n1131));
  xor_4  g0856(.A(new_n1131), .B(new_n1128), .Y(po028));
  xor_4  g0857(.A(new_n741), .B(new_n368), .Y(po030));
  or_6   g0858(.A(new_n422), .B(new_n414), .Y(new_n1134));
  nand_5 g0859(.A(new_n423), .B(new_n371), .Y(new_n1135));
  nand_5 g0860(.A(new_n1135), .B(new_n1134), .Y(new_n1136));
  xor_4  g0861(.A(new_n1136), .B(new_n1063), .Y(new_n1137));
  xor_4  g0862(.A(new_n1137), .B(new_n364), .Y(po031));
  not_8  g0863(.A(new_n1122), .Y(new_n1139));
  xor_4  g0864(.A(new_n1094), .B(new_n689), .Y(po040));
  nor_5  g0865(.A(po040), .B(new_n1121), .Y(new_n1141));
  nor_5  g0866(.A(new_n1141), .B(new_n1139), .Y(po032));
  xor_4  g0867(.A(po071), .B(new_n1110), .Y(po033));
  xor_4  g0868(.A(new_n1056), .B(new_n361), .Y(new_n1144));
  nand_5 g0869(.A(new_n1136), .B(new_n1063), .Y(new_n1145));
  nand_5 g0870(.A(new_n1137), .B(new_n366), .Y(new_n1146));
  nand_5 g0871(.A(new_n1146), .B(new_n1145), .Y(new_n1147));
  not_8  g0872(.A(new_n1147), .Y(new_n1148));
  xor_4  g0873(.A(new_n1148), .B(new_n1144), .Y(po034));
  not_8  g0874(.A(new_n827), .Y(new_n1150));
  or_6   g0875(.A(new_n833), .B(new_n1150), .Y(new_n1151));
  nand_5 g0876(.A(new_n971), .B(new_n1151), .Y(new_n1152));
  nand_5 g0877(.A(new_n972), .B(po047), .Y(new_n1153));
  nand_5 g0878(.A(new_n1153), .B(new_n1152), .Y(po035));
  xnor_4 g0879(.A(new_n1001), .B(new_n1000), .Y(new_n1155));
  xor_4  g0880(.A(new_n1155), .B(new_n1007), .Y(po036));
  xor_4  g0881(.A(new_n622), .B(new_n621), .Y(po037));
  xor_4  g0882(.A(new_n387), .B(new_n367), .Y(po038));
  nand_5 g0883(.A(new_n1124), .B(new_n482), .Y(new_n1159));
  xor_4  g0884(.A(new_n1159), .B(new_n496), .Y(new_n1160));
  nand_5 g0885(.A(new_n1160), .B(new_n947), .Y(new_n1161));
  xor_4  g0886(.A(new_n1160), .B(new_n947), .Y(new_n1162));
  nand_5 g0887(.A(new_n1125), .B(new_n950), .Y(new_n1163));
  xor_4  g0888(.A(new_n1125), .B(new_n950), .Y(new_n1164));
  nand_5 g0889(.A(new_n1028), .B(new_n354), .Y(new_n1165));
  xor_4  g0890(.A(new_n1028), .B(new_n354), .Y(new_n1166));
  nor_5  g0891(.A(new_n1051), .B(new_n954), .Y(new_n1167));
  xor_4  g0892(.A(new_n1051), .B(new_n954), .Y(new_n1168));
  nand_5 g0893(.A(new_n1056), .B(new_n361), .Y(new_n1169));
  nand_5 g0894(.A(new_n1148), .B(new_n1144), .Y(new_n1170));
  nand_5 g0895(.A(new_n1170), .B(new_n1169), .Y(new_n1171));
  nand_5 g0896(.A(new_n1171), .B(new_n1168), .Y(new_n1172));
  not_8  g0897(.A(new_n1172), .Y(new_n1173));
  nor_5  g0898(.A(new_n1173), .B(new_n1167), .Y(new_n1174));
  not_8  g0899(.A(new_n1174), .Y(new_n1175));
  nand_5 g0900(.A(new_n1175), .B(new_n1166), .Y(new_n1176));
  nand_5 g0901(.A(new_n1176), .B(new_n1165), .Y(new_n1177));
  nand_5 g0902(.A(new_n1177), .B(new_n1164), .Y(new_n1178));
  nand_5 g0903(.A(new_n1178), .B(new_n1163), .Y(new_n1179));
  nand_5 g0904(.A(new_n1179), .B(new_n1162), .Y(new_n1180));
  nand_5 g0905(.A(new_n1180), .B(new_n1161), .Y(new_n1181));
  nor_5  g0906(.A(new_n1159), .B(new_n496), .Y(new_n1182));
  xor_4  g0907(.A(new_n1182), .B(new_n757), .Y(new_n1183));
  xor_4  g0908(.A(new_n1183), .B(new_n945), .Y(new_n1184));
  xor_4  g0909(.A(new_n1184), .B(new_n1181), .Y(po041));
  xor_4  g0910(.A(new_n947), .B(new_n916), .Y(new_n1186));
  nand_5 g0911(.A(new_n950), .B(new_n925), .Y(new_n1187));
  xor_4  g0912(.A(new_n950), .B(new_n925), .Y(new_n1188));
  nand_5 g0913(.A(new_n929), .B(new_n354), .Y(new_n1189));
  xor_4  g0914(.A(new_n929), .B(new_n354), .Y(new_n1190));
  nand_5 g0915(.A(new_n871), .B(new_n357), .Y(new_n1191));
  xor_4  g0916(.A(new_n871), .B(new_n357), .Y(new_n1192));
  nand_5 g0917(.A(new_n873), .B(new_n361), .Y(new_n1193));
  nand_5 g0918(.A(new_n877), .B(new_n364), .Y(new_n1194));
  xor_4  g0919(.A(new_n877), .B(new_n364), .Y(new_n1195));
  nand_5 g0920(.A(new_n887), .B(new_n376), .Y(new_n1196));
  or_6   g0921(.A(new_n1196), .B(new_n374), .Y(new_n1197));
  nand_5 g0922(.A(new_n1196), .B(new_n379), .Y(new_n1198));
  nand_5 g0923(.A(new_n1198), .B(new_n1197), .Y(new_n1199));
  or_6   g0924(.A(new_n1199), .B(new_n891), .Y(new_n1200));
  nand_5 g0925(.A(new_n1200), .B(new_n1197), .Y(new_n1201));
  nor_5  g0926(.A(new_n1201), .B(new_n882), .Y(new_n1202));
  xor_4  g0927(.A(new_n1201), .B(new_n882), .Y(new_n1203));
  nand_5 g0928(.A(new_n1203), .B(new_n371), .Y(new_n1204));
  not_8  g0929(.A(new_n1204), .Y(new_n1205));
  nor_5  g0930(.A(new_n1205), .B(new_n1202), .Y(new_n1206));
  nand_5 g0931(.A(new_n1206), .B(new_n1195), .Y(new_n1207));
  nand_5 g0932(.A(new_n1207), .B(new_n1194), .Y(new_n1208));
  xor_4  g0933(.A(new_n873), .B(new_n361), .Y(new_n1209));
  nand_5 g0934(.A(new_n1209), .B(new_n1208), .Y(new_n1210));
  nand_5 g0935(.A(new_n1210), .B(new_n1193), .Y(new_n1211));
  nand_5 g0936(.A(new_n1211), .B(new_n1192), .Y(new_n1212));
  nand_5 g0937(.A(new_n1212), .B(new_n1191), .Y(new_n1213));
  nand_5 g0938(.A(new_n1213), .B(new_n1190), .Y(new_n1214));
  nand_5 g0939(.A(new_n1214), .B(new_n1189), .Y(new_n1215));
  nand_5 g0940(.A(new_n1215), .B(new_n1188), .Y(new_n1216));
  nand_5 g0941(.A(new_n1216), .B(new_n1187), .Y(new_n1217));
  xor_4  g0942(.A(new_n1217), .B(new_n1186), .Y(po042));
  xor_4  g0943(.A(new_n947), .B(new_n697), .Y(new_n1219));
  nand_5 g0944(.A(new_n950), .B(new_n582), .Y(new_n1220));
  xor_4  g0945(.A(new_n950), .B(new_n582), .Y(new_n1221));
  nand_5 g0946(.A(new_n606), .B(new_n354), .Y(new_n1222));
  xor_4  g0947(.A(new_n606), .B(new_n354), .Y(new_n1223));
  nand_5 g0948(.A(new_n610), .B(new_n357), .Y(new_n1224));
  xor_4  g0949(.A(new_n610), .B(new_n357), .Y(new_n1225));
  nand_5 g0950(.A(new_n613), .B(new_n361), .Y(new_n1226));
  not_8  g0951(.A(new_n1226), .Y(new_n1227));
  nor_5  g0952(.A(new_n993), .B(new_n979), .Y(new_n1228));
  nor_5  g0953(.A(new_n1228), .B(new_n1227), .Y(new_n1229));
  not_8  g0954(.A(new_n1229), .Y(new_n1230));
  nand_5 g0955(.A(new_n1230), .B(new_n1225), .Y(new_n1231));
  nand_5 g0956(.A(new_n1231), .B(new_n1224), .Y(new_n1232));
  nand_5 g0957(.A(new_n1232), .B(new_n1223), .Y(new_n1233));
  nand_5 g0958(.A(new_n1233), .B(new_n1222), .Y(new_n1234));
  nand_5 g0959(.A(new_n1234), .B(new_n1221), .Y(new_n1235));
  nand_5 g0960(.A(new_n1235), .B(new_n1220), .Y(new_n1236));
  xor_4  g0961(.A(new_n1236), .B(new_n1219), .Y(po043));
  xor_4  g0962(.A(new_n973), .B(new_n967), .Y(po044));
  or_6   g0963(.A(new_n332), .B(new_n321), .Y(new_n1239));
  nor_5  g0964(.A(new_n331), .B(new_n322), .Y(new_n1240));
  xor_4  g0965(.A(new_n328), .B(new_n468), .Y(new_n1241));
  nand_5 g0966(.A(new_n1241), .B(pi60), .Y(new_n1242));
  nor_5  g0967(.A(new_n654), .B(pi39), .Y(new_n1243));
  nand_5 g0968(.A(new_n315), .B(new_n473), .Y(new_n1244));
  nand_5 g0969(.A(new_n1244), .B(pi78), .Y(new_n1245));
  nand_5 g0970(.A(new_n1245), .B(new_n277), .Y(new_n1246));
  or_6   g0971(.A(new_n1246), .B(new_n1243), .Y(new_n1247));
  nand_5 g0972(.A(new_n1247), .B(new_n1242), .Y(new_n1248));
  xor_4  g0973(.A(new_n1248), .B(new_n1240), .Y(new_n1249));
  or_6   g0974(.A(new_n1249), .B(new_n1239), .Y(new_n1250));
  nand_5 g0975(.A(new_n1248), .B(new_n1240), .Y(new_n1251));
  xor_4  g0976(.A(new_n1243), .B(pi20), .Y(new_n1252));
  nand_5 g0977(.A(new_n1252), .B(new_n277), .Y(new_n1253));
  nand_5 g0978(.A(new_n328), .B(pi13), .Y(new_n1254));
  nor_5  g0979(.A(new_n1254), .B(new_n492), .Y(new_n1255));
  nand_5 g0980(.A(new_n1254), .B(new_n492), .Y(new_n1256));
  nand_5 g0981(.A(new_n1256), .B(pi60), .Y(new_n1257));
  or_6   g0982(.A(new_n1257), .B(new_n1255), .Y(new_n1258));
  nand_5 g0983(.A(new_n1258), .B(new_n1253), .Y(new_n1259));
  xor_4  g0984(.A(new_n1259), .B(new_n1251), .Y(new_n1260));
  or_6   g0985(.A(new_n1260), .B(new_n1250), .Y(new_n1261));
  nor_5  g0986(.A(new_n1259), .B(new_n1251), .Y(new_n1262));
  xor_4  g0987(.A(new_n1255), .B(new_n666), .Y(new_n1263));
  nand_5 g0988(.A(new_n1263), .B(pi60), .Y(new_n1264));
  nand_5 g0989(.A(new_n1243), .B(new_n487), .Y(new_n1265));
  nand_5 g0990(.A(new_n1265), .B(pi66), .Y(new_n1266));
  nor_5  g0991(.A(new_n1265), .B(pi66), .Y(new_n1267));
  nor_5  g0992(.A(new_n1267), .B(pi60), .Y(new_n1268));
  nand_5 g0993(.A(new_n1268), .B(new_n1266), .Y(new_n1269));
  nand_5 g0994(.A(new_n1269), .B(new_n1264), .Y(new_n1270));
  xor_4  g0995(.A(new_n1270), .B(new_n1262), .Y(new_n1271));
  or_6   g0996(.A(new_n1271), .B(new_n1261), .Y(new_n1272));
  nand_5 g0997(.A(new_n1270), .B(new_n1262), .Y(new_n1273));
  xor_4  g0998(.A(new_n1267), .B(pi74), .Y(new_n1274));
  nand_5 g0999(.A(new_n1274), .B(new_n277), .Y(new_n1275));
  nand_5 g1000(.A(new_n1255), .B(pi09), .Y(new_n1276));
  nand_5 g1001(.A(new_n1276), .B(new_n769), .Y(new_n1277));
  nor_5  g1002(.A(new_n1276), .B(new_n769), .Y(new_n1278));
  nor_5  g1003(.A(new_n1278), .B(new_n277), .Y(new_n1279));
  nand_5 g1004(.A(new_n1279), .B(new_n1277), .Y(new_n1280));
  nand_5 g1005(.A(new_n1280), .B(new_n1275), .Y(new_n1281));
  xor_4  g1006(.A(new_n1281), .B(new_n1273), .Y(new_n1282));
  nor_5  g1007(.A(new_n1282), .B(new_n1272), .Y(new_n1283));
  not_8  g1008(.A(new_n1283), .Y(new_n1284));
  nand_5 g1009(.A(new_n1267), .B(new_n679), .Y(new_n1285));
  nor_5  g1010(.A(new_n1285), .B(pi60), .Y(new_n1286));
  not_8  g1011(.A(new_n1286), .Y(new_n1287));
  nor_5  g1012(.A(new_n1281), .B(new_n1273), .Y(new_n1288));
  nand_5 g1013(.A(new_n1278), .B(pi60), .Y(new_n1289));
  nand_5 g1014(.A(new_n1289), .B(new_n1287), .Y(new_n1290));
  not_8  g1015(.A(new_n1290), .Y(new_n1291));
  nand_5 g1016(.A(new_n1291), .B(new_n1288), .Y(new_n1292));
  nand_5 g1017(.A(new_n1292), .B(new_n1287), .Y(new_n1293));
  nand_5 g1018(.A(new_n1293), .B(new_n1284), .Y(new_n1294));
  xor_4  g1019(.A(new_n1282), .B(new_n1272), .Y(new_n1295));
  xor_4  g1020(.A(new_n1271), .B(new_n1261), .Y(new_n1296));
  not_8  g1021(.A(pi15), .Y(new_n1297));
  not_8  g1022(.A(pi83), .Y(new_n1298));
  nand_5 g1023(.A(pi85), .B(pi27), .Y(new_n1299));
  nand_5 g1024(.A(new_n724), .B(new_n710), .Y(new_n1300));
  nand_5 g1025(.A(new_n1300), .B(new_n1299), .Y(new_n1301));
  nand_5 g1026(.A(new_n1301), .B(pi05), .Y(new_n1302));
  nor_5  g1027(.A(new_n1302), .B(new_n1298), .Y(new_n1303));
  nand_5 g1028(.A(new_n1303), .B(pi53), .Y(new_n1304));
  nor_5  g1029(.A(new_n1304), .B(new_n1297), .Y(new_n1305));
  nand_5 g1030(.A(new_n1305), .B(new_n1296), .Y(new_n1306));
  xor_4  g1031(.A(new_n1260), .B(new_n1250), .Y(new_n1307));
  xor_4  g1032(.A(new_n1304), .B(new_n1297), .Y(new_n1308));
  nand_5 g1033(.A(new_n1308), .B(new_n1307), .Y(new_n1309));
  xor_4  g1034(.A(new_n1308), .B(new_n1307), .Y(new_n1310));
  xor_4  g1035(.A(new_n1249), .B(new_n1239), .Y(new_n1311));
  xor_4  g1036(.A(new_n1303), .B(pi53), .Y(new_n1312));
  nand_5 g1037(.A(new_n1312), .B(new_n1311), .Y(new_n1313));
  xor_4  g1038(.A(new_n1312), .B(new_n1311), .Y(new_n1314));
  xor_4  g1039(.A(new_n1302), .B(new_n1298), .Y(new_n1315));
  nand_5 g1040(.A(new_n1315), .B(new_n333), .Y(new_n1316));
  xor_4  g1041(.A(new_n1315), .B(new_n333), .Y(new_n1317));
  xor_4  g1042(.A(new_n1301), .B(pi05), .Y(new_n1318));
  nand_5 g1043(.A(new_n1318), .B(new_n356), .Y(new_n1319));
  xor_4  g1044(.A(new_n1318), .B(new_n356), .Y(new_n1320));
  nand_5 g1045(.A(new_n725), .B(new_n360), .Y(new_n1321));
  nand_5 g1046(.A(new_n745), .B(new_n726), .Y(new_n1322));
  nand_5 g1047(.A(new_n1322), .B(new_n1321), .Y(new_n1323));
  nand_5 g1048(.A(new_n1323), .B(new_n1320), .Y(new_n1324));
  nand_5 g1049(.A(new_n1324), .B(new_n1319), .Y(new_n1325));
  nand_5 g1050(.A(new_n1325), .B(new_n1317), .Y(new_n1326));
  nand_5 g1051(.A(new_n1326), .B(new_n1316), .Y(new_n1327));
  nand_5 g1052(.A(new_n1327), .B(new_n1314), .Y(new_n1328));
  nand_5 g1053(.A(new_n1328), .B(new_n1313), .Y(new_n1329));
  nand_5 g1054(.A(new_n1329), .B(new_n1310), .Y(new_n1330));
  nand_5 g1055(.A(new_n1330), .B(new_n1309), .Y(new_n1331));
  xor_4  g1056(.A(new_n1305), .B(new_n1296), .Y(new_n1332));
  nand_5 g1057(.A(new_n1332), .B(new_n1331), .Y(new_n1333));
  nand_5 g1058(.A(new_n1333), .B(new_n1306), .Y(new_n1334));
  nand_5 g1059(.A(new_n1334), .B(new_n1295), .Y(new_n1335));
  not_8  g1060(.A(new_n1335), .Y(new_n1336));
  nor_5  g1061(.A(new_n1336), .B(new_n1294), .Y(po045));
  xor_4  g1062(.A(po176), .B(new_n507), .Y(po046));
  nand_5 g1063(.A(new_n1001), .B(new_n945), .Y(new_n1339));
  nand_5 g1064(.A(new_n947), .B(new_n916), .Y(new_n1340));
  nand_5 g1065(.A(new_n1217), .B(new_n1186), .Y(new_n1341));
  nand_5 g1066(.A(new_n1341), .B(new_n1340), .Y(new_n1342));
  xor_4  g1067(.A(new_n1001), .B(new_n945), .Y(new_n1343));
  nand_5 g1068(.A(new_n1343), .B(new_n1342), .Y(new_n1344));
  nand_5 g1069(.A(new_n1344), .B(new_n1339), .Y(new_n1345));
  nand_5 g1070(.A(new_n1345), .B(new_n999), .Y(new_n1346));
  not_8  g1071(.A(new_n1346), .Y(new_n1347));
  nor_5  g1072(.A(new_n1347), .B(new_n1015), .Y(po048));
  xor_4  g1073(.A(new_n1232), .B(new_n1223), .Y(po049));
  xor_4  g1074(.A(new_n1209), .B(new_n1208), .Y(po051));
  xor_4  g1075(.A(new_n1343), .B(new_n1342), .Y(po052));
  xor_4  g1076(.A(po029), .B(new_n504), .Y(po053));
  nand_5 g1077(.A(new_n1095), .B(new_n1013), .Y(new_n1353));
  nor_5  g1078(.A(new_n1139), .B(new_n1353), .Y(po054));
  xor_4  g1079(.A(new_n1010), .B(new_n999), .Y(po055));
  nor_5  g1080(.A(new_n773), .B(new_n761), .Y(new_n1356));
  not_8  g1081(.A(new_n1356), .Y(new_n1357));
  or_6   g1082(.A(new_n762), .B(pi31), .Y(new_n1358));
  nor_5  g1083(.A(new_n1358), .B(new_n396), .Y(new_n1359));
  nand_5 g1084(.A(new_n684), .B(new_n399), .Y(new_n1360));
  not_8  g1085(.A(new_n1360), .Y(new_n1361));
  nor_5  g1086(.A(new_n1361), .B(new_n1359), .Y(new_n1362));
  not_8  g1087(.A(new_n1362), .Y(new_n1363));
  nand_5 g1088(.A(new_n1363), .B(new_n1357), .Y(new_n1364));
  not_8  g1089(.A(new_n1364), .Y(po056));
  xor_4  g1090(.A(new_n1323), .B(new_n1320), .Y(po059));
  xor_4  g1091(.A(new_n646), .B(new_n645), .Y(po060));
  xor_4  g1092(.A(new_n938), .B(new_n928), .Y(po061));
  not_8  g1093(.A(new_n945), .Y(new_n1369));
  nand_5 g1094(.A(new_n1294), .B(new_n1369), .Y(new_n1370));
  xor_4  g1095(.A(new_n1291), .B(new_n1288), .Y(new_n1371));
  xor_4  g1096(.A(new_n1371), .B(new_n1283), .Y(new_n1372));
  xor_4  g1097(.A(new_n1295), .B(new_n1369), .Y(new_n1373));
  nor_5  g1098(.A(new_n1296), .B(new_n945), .Y(new_n1374));
  and_6  g1099(.A(new_n1296), .B(new_n945), .Y(new_n1375));
  nand_5 g1100(.A(new_n1307), .B(new_n947), .Y(new_n1376));
  xor_4  g1101(.A(new_n1307), .B(new_n947), .Y(new_n1377));
  nand_5 g1102(.A(new_n1311), .B(new_n950), .Y(new_n1378));
  xor_4  g1103(.A(new_n1311), .B(new_n950), .Y(new_n1379));
  nand_5 g1104(.A(new_n354), .B(new_n333), .Y(new_n1380));
  nand_5 g1105(.A(new_n394), .B(new_n355), .Y(new_n1381));
  nand_5 g1106(.A(new_n1381), .B(new_n1380), .Y(new_n1382));
  nand_5 g1107(.A(new_n1382), .B(new_n1379), .Y(new_n1383));
  nand_5 g1108(.A(new_n1383), .B(new_n1378), .Y(new_n1384));
  nand_5 g1109(.A(new_n1384), .B(new_n1377), .Y(new_n1385));
  nand_5 g1110(.A(new_n1385), .B(new_n1376), .Y(new_n1386));
  nor_5  g1111(.A(new_n1386), .B(new_n1375), .Y(new_n1387));
  or_6   g1112(.A(new_n1387), .B(new_n1374), .Y(new_n1388));
  nor_5  g1113(.A(new_n1388), .B(new_n1373), .Y(new_n1389));
  or_6   g1114(.A(new_n1295), .B(new_n1369), .Y(new_n1390));
  or_6   g1115(.A(new_n1390), .B(new_n1389), .Y(new_n1391));
  nand_5 g1116(.A(new_n1389), .B(new_n1369), .Y(new_n1392));
  nand_5 g1117(.A(new_n1392), .B(new_n1391), .Y(new_n1393));
  xor_4  g1118(.A(new_n1393), .B(new_n1372), .Y(new_n1394));
  not_8  g1119(.A(new_n1394), .Y(po112));
  and_6  g1120(.A(po112), .B(new_n1370), .Y(po062));
  xor_4  g1121(.A(new_n737), .B(new_n383), .Y(po063));
  nor_5  g1122(.A(new_n1113), .B(po010), .Y(new_n1398));
  nor_5  g1123(.A(new_n1398), .B(new_n1115), .Y(po065));
  xor_4  g1124(.A(po100), .B(new_n1102), .Y(po066));
  xor_4  g1125(.A(new_n1234), .B(new_n1221), .Y(po067));
  xor_4  g1126(.A(new_n1382), .B(new_n1379), .Y(po068));
  xor_4  g1127(.A(new_n1177), .B(new_n1164), .Y(po069));
  nand_5 g1128(.A(new_n976), .B(new_n966), .Y(new_n1404));
  nand_5 g1129(.A(new_n1369), .B(new_n680), .Y(new_n1405));
  nand_5 g1130(.A(new_n965), .B(new_n946), .Y(new_n1406));
  nand_5 g1131(.A(new_n1406), .B(new_n1405), .Y(new_n1407));
  nand_5 g1132(.A(new_n1407), .B(new_n679), .Y(new_n1408));
  nor_5  g1133(.A(new_n1408), .B(new_n1404), .Y(po070));
  xor_4  g1134(.A(new_n1211), .B(new_n1192), .Y(po072));
  xor_4  g1135(.A(new_n945), .B(new_n692), .Y(new_n1411));
  or_6   g1136(.A(new_n947), .B(new_n697), .Y(new_n1412));
  not_8  g1137(.A(new_n1412), .Y(new_n1413));
  not_8  g1138(.A(new_n1219), .Y(new_n1414));
  nor_5  g1139(.A(new_n1236), .B(new_n1414), .Y(new_n1415));
  nor_5  g1140(.A(new_n1415), .B(new_n1413), .Y(new_n1416));
  xor_4  g1141(.A(new_n1416), .B(new_n1411), .Y(po073));
  xor_4  g1142(.A(new_n903), .B(new_n876), .Y(po074));
  xor_4  g1143(.A(new_n1077), .B(new_n414), .Y(po075));
  not_8  g1144(.A(new_n1353), .Y(po076));
  xor_4  g1145(.A(new_n420), .B(new_n418), .Y(po077));
  xor_4  g1146(.A(new_n1384), .B(new_n1377), .Y(po078));
  xor_4  g1147(.A(new_n1083), .B(new_n1055), .Y(po079));
  xor_4  g1148(.A(new_n1092), .B(new_n661), .Y(po080));
  xor_4  g1149(.A(new_n1215), .B(new_n1188), .Y(po081));
  nand_5 g1150(.A(new_n1182), .B(new_n757), .Y(new_n1426));
  xor_4  g1151(.A(new_n1426), .B(new_n773), .Y(new_n1427));
  nand_5 g1152(.A(new_n1183), .B(new_n945), .Y(new_n1428));
  nand_5 g1153(.A(new_n1184), .B(new_n1181), .Y(new_n1429));
  nand_5 g1154(.A(new_n1429), .B(new_n1428), .Y(new_n1430));
  xor_4  g1155(.A(new_n1430), .B(new_n1427), .Y(po082));
  xor_4  g1156(.A(new_n648), .B(new_n609), .Y(po083));
  not_8  g1157(.A(pi49), .Y(new_n1433));
  nand_5 g1158(.A(new_n1126), .B(pi90), .Y(new_n1434));
  nor_5  g1159(.A(new_n1434), .B(new_n1433), .Y(new_n1435));
  nor_5  g1160(.A(new_n1435), .B(new_n1183), .Y(new_n1436));
  nand_5 g1161(.A(new_n1435), .B(new_n1183), .Y(new_n1437));
  xor_4  g1162(.A(new_n1434), .B(new_n1433), .Y(new_n1438));
  nand_5 g1163(.A(new_n1438), .B(new_n1160), .Y(new_n1439));
  not_8  g1164(.A(new_n1439), .Y(new_n1440));
  xnor_4 g1165(.A(new_n1438), .B(new_n1160), .Y(new_n1441));
  or_6   g1166(.A(new_n1127), .B(new_n1125), .Y(new_n1442));
  not_8  g1167(.A(new_n1131), .Y(new_n1443));
  nand_5 g1168(.A(new_n1443), .B(new_n1128), .Y(new_n1444));
  nand_5 g1169(.A(new_n1444), .B(new_n1442), .Y(new_n1445));
  nor_5  g1170(.A(new_n1445), .B(new_n1441), .Y(new_n1446));
  nor_5  g1171(.A(new_n1446), .B(new_n1440), .Y(new_n1447));
  nand_5 g1172(.A(new_n1447), .B(new_n1437), .Y(new_n1448));
  not_8  g1173(.A(new_n1448), .Y(new_n1449));
  nor_5  g1174(.A(new_n1449), .B(new_n1436), .Y(new_n1450));
  xor_4  g1175(.A(new_n1450), .B(new_n1427), .Y(po084));
  nand_5 g1176(.A(new_n1450), .B(new_n1427), .Y(new_n1452));
  not_8  g1177(.A(new_n1452), .Y(new_n1453));
  or_6   g1178(.A(new_n1426), .B(new_n773), .Y(new_n1454));
  nand_5 g1179(.A(new_n1454), .B(new_n1363), .Y(new_n1455));
  nor_5  g1180(.A(new_n1455), .B(new_n1453), .Y(po085));
  xor_4  g1181(.A(new_n888), .B(new_n887), .Y(po086));
  xor_4  g1182(.A(new_n991), .B(new_n364), .Y(po087));
  nand_5 g1183(.A(new_n974), .B(po047), .Y(new_n1459));
  not_8  g1184(.A(new_n968), .Y(new_n1460));
  nand_5 g1185(.A(new_n1153), .B(new_n1460), .Y(new_n1461));
  nand_5 g1186(.A(new_n1461), .B(new_n1459), .Y(po088));
  xor_4  g1187(.A(po111), .B(new_n519), .Y(po089));
  xor_4  g1188(.A(po107), .B(new_n1115), .Y(po090));
  xor_4  g1189(.A(new_n936), .B(new_n934), .Y(po091));
  nand_5 g1190(.A(po070), .B(po047), .Y(new_n1466));
  not_8  g1191(.A(new_n1466), .Y(po092));
  xor_4  g1192(.A(new_n392), .B(new_n359), .Y(po093));
  nand_5 g1193(.A(new_n708), .B(new_n691), .Y(new_n1469));
  nor_5  g1194(.A(new_n690), .B(new_n676), .Y(new_n1470));
  nor_5  g1195(.A(new_n689), .B(new_n677), .Y(new_n1471));
  nor_5  g1196(.A(new_n1013), .B(new_n1471), .Y(new_n1472));
  nor_5  g1197(.A(new_n1472), .B(new_n1470), .Y(new_n1473));
  and_6  g1198(.A(new_n1473), .B(new_n1469), .Y(po094));
  xor_4  g1199(.A(new_n1213), .B(new_n1190), .Y(po095));
  xor_4  g1200(.A(new_n1388), .B(new_n1373), .Y(po096));
  xor_4  g1201(.A(new_n1445), .B(new_n1441), .Y(po097));
  xor_4  g1202(.A(new_n1179), .B(new_n1162), .Y(po098));
  xor_4  g1203(.A(new_n831), .B(new_n827), .Y(po099));
  not_8  g1204(.A(new_n1469), .Y(new_n1480));
  xor_4  g1205(.A(new_n1472), .B(new_n1470), .Y(new_n1481));
  or_6   g1206(.A(new_n1481), .B(new_n1480), .Y(new_n1482));
  nand_5 g1207(.A(new_n1472), .B(new_n1480), .Y(new_n1483));
  nand_5 g1208(.A(new_n1483), .B(new_n1482), .Y(po101));
  xnor_4 g1209(.A(new_n1435), .B(new_n1183), .Y(new_n1485));
  xor_4  g1210(.A(new_n1485), .B(new_n1447), .Y(po102));
  xor_4  g1211(.A(new_n703), .B(new_n700), .Y(po103));
  nor_5  g1212(.A(new_n1452), .B(new_n1362), .Y(new_n1488));
  xor_4  g1213(.A(new_n1454), .B(new_n1362), .Y(new_n1489));
  nor_5  g1214(.A(new_n1489), .B(new_n1453), .Y(new_n1490));
  nor_5  g1215(.A(new_n1490), .B(new_n1488), .Y(po104));
  xor_4  g1216(.A(po064), .B(new_n510), .Y(po105));
  xor_4  g1217(.A(new_n415), .B(new_n376), .Y(po106));
  nor_5  g1218(.A(new_n1407), .B(new_n679), .Y(new_n1494));
  and_6  g1219(.A(new_n1494), .B(new_n1404), .Y(new_n1495));
  or_6   g1220(.A(new_n1495), .B(po070), .Y(po108));
  nor_5  g1221(.A(new_n1371), .B(new_n1335), .Y(new_n1497));
  and_6  g1222(.A(new_n1372), .B(new_n1335), .Y(new_n1498));
  nor_5  g1223(.A(new_n1498), .B(new_n1497), .Y(po110));
  xor_4  g1224(.A(new_n970), .B(new_n969), .Y(po113));
  nor_5  g1225(.A(po080), .B(new_n1118), .Y(new_n1501));
  nor_5  g1226(.A(new_n1501), .B(new_n1120), .Y(po114));
  nand_5 g1227(.A(new_n945), .B(new_n692), .Y(new_n1503));
  nand_5 g1228(.A(new_n1416), .B(new_n1411), .Y(new_n1504));
  nand_5 g1229(.A(new_n1504), .B(new_n1503), .Y(new_n1505));
  not_8  g1230(.A(new_n1505), .Y(new_n1506));
  or_6   g1231(.A(new_n1369), .B(new_n691), .Y(new_n1507));
  nand_5 g1232(.A(new_n1507), .B(new_n1506), .Y(new_n1508));
  nand_5 g1233(.A(new_n1369), .B(new_n691), .Y(new_n1509));
  nand_5 g1234(.A(new_n1509), .B(new_n1505), .Y(new_n1510));
  nand_5 g1235(.A(new_n1510), .B(new_n1508), .Y(new_n1511));
  xor_4  g1236(.A(new_n1511), .B(new_n1481), .Y(po116));
  xor_4  g1237(.A(new_n972), .B(new_n1460), .Y(po117));
  xor_4  g1238(.A(new_n390), .B(new_n389), .Y(po118));
  xor_4  g1239(.A(new_n1203), .B(new_n370), .Y(po119));
  not_8  g1240(.A(new_n792), .Y(new_n1516));
  nand_5 g1241(.A(new_n1099), .B(new_n1516), .Y(new_n1517));
  nand_5 g1242(.A(new_n1517), .B(new_n1103), .Y(po120));
  xor_4  g1243(.A(po050), .B(new_n1107), .Y(po121));
  xor_4  g1244(.A(new_n975), .B(new_n966), .Y(po122));
  nand_5 g1245(.A(new_n998), .B(new_n689), .Y(new_n1521));
  xor_4  g1246(.A(new_n1014), .B(new_n1521), .Y(new_n1522));
  nor_5  g1247(.A(new_n1522), .B(new_n1012), .Y(new_n1523));
  nor_5  g1248(.A(new_n1014), .B(new_n1011), .Y(new_n1524));
  nor_5  g1249(.A(new_n1524), .B(new_n1523), .Y(po126));
  xor_4  g1250(.A(new_n1120), .B(po124), .Y(po127));
  nand_5 g1251(.A(new_n1430), .B(new_n1427), .Y(new_n1527));
  not_8  g1252(.A(new_n1527), .Y(new_n1528));
  nor_5  g1253(.A(new_n1455), .B(new_n1528), .Y(po128));
  xor_4  g1254(.A(new_n383), .B(new_n381), .Y(po129));
  not_8  g1255(.A(new_n977), .Y(new_n1531));
  nand_5 g1256(.A(new_n1531), .B(new_n966), .Y(new_n1532));
  nand_5 g1257(.A(new_n1494), .B(new_n1532), .Y(new_n1533));
  nand_5 g1258(.A(new_n1533), .B(new_n1466), .Y(po130));
  xor_4  g1259(.A(new_n512), .B(po177), .Y(po131));
  xor_4  g1260(.A(new_n1329), .B(new_n1310), .Y(po132));
  xor_4  g1261(.A(new_n1230), .B(new_n1225), .Y(po133));
  xor_4  g1262(.A(new_n628), .B(new_n625), .Y(po134));
  xor_4  g1263(.A(new_n1334), .B(new_n1295), .Y(po135));
  xor_4  g1264(.A(new_n1362), .B(new_n1356), .Y(new_n1540));
  not_8  g1265(.A(new_n1540), .Y(po136));
  xor_4  g1266(.A(new_n1081), .B(new_n1059), .Y(po137));
  xor_4  g1267(.A(new_n1407), .B(new_n679), .Y(new_n1543));
  xnor_4 g1268(.A(new_n1543), .B(new_n1404), .Y(po138));
  xnor_4 g1269(.A(new_n1543), .B(new_n1532), .Y(po139));
  xor_4  g1270(.A(new_n1325), .B(new_n1317), .Y(po141));
  xor_4  g1271(.A(new_n1199), .B(new_n891), .Y(po142));
  xor_4  g1272(.A(new_n987), .B(new_n370), .Y(po143));
  not_8  g1273(.A(new_n1096), .Y(po144));
  not_8  g1274(.A(po047), .Y(po145));
  nor_5  g1275(.A(new_n1364), .B(new_n778), .Y(po146));
  not_8  g1276(.A(new_n829), .Y(new_n1552));
  xor_4  g1277(.A(po162), .B(new_n1552), .Y(po147));
  xor_4  g1278(.A(new_n983), .B(new_n625), .Y(po149));
  nand_5 g1279(.A(new_n1509), .B(new_n1507), .Y(new_n1555));
  xor_4  g1280(.A(new_n1555), .B(new_n1505), .Y(po150));
  not_8  g1281(.A(new_n967), .Y(new_n1557));
  nand_5 g1282(.A(new_n1459), .B(new_n1557), .Y(new_n1558));
  nand_5 g1283(.A(new_n1558), .B(new_n977), .Y(po151));
  xor_4  g1284(.A(new_n887), .B(new_n376), .Y(po152));
  xor_4  g1285(.A(new_n634), .B(new_n632), .Y(po153));
  xor_4  g1286(.A(new_n900), .B(new_n881), .Y(po154));
  xor_4  g1287(.A(new_n1327), .B(new_n1314), .Y(po155));
  xor_4  g1288(.A(new_n1079), .B(new_n1064), .Y(po156));
  xor_4  g1289(.A(po172), .B(new_n1105), .Y(po157));
  xor_4  g1290(.A(new_n640), .B(new_n639), .Y(po158));
  xor_4  g1291(.A(po162), .B(po145), .Y(po159));
  xor_4  g1292(.A(new_n1540), .B(new_n777), .Y(po160));
  xor_4  g1293(.A(new_n1206), .B(new_n1195), .Y(po161));
  nand_5 g1294(.A(new_n501), .B(new_n441), .Y(new_n1570));
  nand_5 g1295(.A(new_n1570), .B(new_n505), .Y(po163));
  xor_4  g1296(.A(new_n1072), .B(new_n418), .Y(po164));
  or_6   g1297(.A(new_n1473), .B(new_n945), .Y(new_n1573));
  and_6  g1298(.A(new_n1573), .B(po116), .Y(po165));
  nand_5 g1299(.A(po162), .B(po047), .Y(new_n1575));
  nand_5 g1300(.A(new_n1575), .B(new_n1552), .Y(new_n1576));
  nand_5 g1301(.A(new_n1576), .B(new_n833), .Y(po166));
  xor_4  g1302(.A(new_n1175), .B(new_n1166), .Y(po167));
  xor_4  g1303(.A(new_n515), .B(po109), .Y(po168));
  nor_5  g1304(.A(new_n1527), .B(new_n1362), .Y(new_n1580));
  nor_5  g1305(.A(new_n1489), .B(new_n1528), .Y(new_n1581));
  nor_5  g1306(.A(new_n1581), .B(new_n1580), .Y(po169));
  xor_4  g1307(.A(new_n894), .B(new_n891), .Y(po170));
  xor_4  g1308(.A(new_n1345), .B(new_n999), .Y(po173));
  xor_4  g1309(.A(new_n621), .B(new_n376), .Y(po174));
  xor_4  g1310(.A(new_n1332), .B(new_n1331), .Y(po175));
  nor_5  g1311(.A(new_n1375), .B(new_n1374), .Y(new_n1587));
  xor_4  g1312(.A(new_n1587), .B(new_n1386), .Y(po178));
  nor_5  g1313(.A(new_n1522), .B(new_n1347), .Y(new_n1589));
  nor_5  g1314(.A(new_n1346), .B(new_n1014), .Y(new_n1590));
  nor_5  g1315(.A(new_n1590), .B(new_n1589), .Y(po180));
  xor_4  g1316(.A(new_n1171), .B(new_n1168), .Y(po181));
  buf_8  g1317(.A(po012), .Y(po039));
  buf_8  g1318(.A(po022), .Y(po171));
endmodule


