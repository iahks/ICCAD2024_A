 module top_809960632_810038711_1598227639_893650103 (a, o);

      input a, b; output o; buf_12 g0(a,o); endmodule